magic
tech sky130l
timestamp 1731220586
<< m2 >>
rect 134 3659 140 3660
rect 134 3655 135 3659
rect 139 3655 140 3659
rect 134 3654 140 3655
rect 222 3659 228 3660
rect 222 3655 223 3659
rect 227 3655 228 3659
rect 222 3654 228 3655
rect 110 3649 116 3650
rect 110 3645 111 3649
rect 115 3645 116 3649
rect 110 3644 116 3645
rect 1822 3649 1828 3650
rect 1822 3645 1823 3649
rect 1827 3645 1828 3649
rect 1822 3644 1828 3645
rect 110 3632 116 3633
rect 110 3628 111 3632
rect 115 3628 116 3632
rect 110 3627 116 3628
rect 1822 3632 1828 3633
rect 1822 3628 1823 3632
rect 1827 3628 1828 3632
rect 1822 3627 1828 3628
rect 142 3619 148 3620
rect 142 3615 143 3619
rect 147 3615 148 3619
rect 142 3614 148 3615
rect 230 3619 236 3620
rect 230 3615 231 3619
rect 235 3615 236 3619
rect 230 3614 236 3615
rect 142 3585 148 3586
rect 142 3581 143 3585
rect 147 3581 148 3585
rect 142 3580 148 3581
rect 230 3585 236 3586
rect 230 3581 231 3585
rect 235 3581 236 3585
rect 230 3580 236 3581
rect 318 3585 324 3586
rect 318 3581 319 3585
rect 323 3581 324 3585
rect 318 3580 324 3581
rect 406 3585 412 3586
rect 406 3581 407 3585
rect 411 3581 412 3585
rect 406 3580 412 3581
rect 494 3585 500 3586
rect 494 3581 495 3585
rect 499 3581 500 3585
rect 494 3580 500 3581
rect 1886 3583 1892 3584
rect 1886 3579 1887 3583
rect 1891 3579 1892 3583
rect 1886 3578 1892 3579
rect 1974 3583 1980 3584
rect 1974 3579 1975 3583
rect 1979 3579 1980 3583
rect 1974 3578 1980 3579
rect 2062 3583 2068 3584
rect 2062 3579 2063 3583
rect 2067 3579 2068 3583
rect 2062 3578 2068 3579
rect 2150 3583 2156 3584
rect 2150 3579 2151 3583
rect 2155 3579 2156 3583
rect 2150 3578 2156 3579
rect 2238 3583 2244 3584
rect 2238 3579 2239 3583
rect 2243 3579 2244 3583
rect 2238 3578 2244 3579
rect 2326 3583 2332 3584
rect 2326 3579 2327 3583
rect 2331 3579 2332 3583
rect 2326 3578 2332 3579
rect 2430 3583 2436 3584
rect 2430 3579 2431 3583
rect 2435 3579 2436 3583
rect 2430 3578 2436 3579
rect 2534 3583 2540 3584
rect 2534 3579 2535 3583
rect 2539 3579 2540 3583
rect 2534 3578 2540 3579
rect 2630 3583 2636 3584
rect 2630 3579 2631 3583
rect 2635 3579 2636 3583
rect 2630 3578 2636 3579
rect 2726 3583 2732 3584
rect 2726 3579 2727 3583
rect 2731 3579 2732 3583
rect 2726 3578 2732 3579
rect 2822 3583 2828 3584
rect 2822 3579 2823 3583
rect 2827 3579 2828 3583
rect 2822 3578 2828 3579
rect 2918 3583 2924 3584
rect 2918 3579 2919 3583
rect 2923 3579 2924 3583
rect 2918 3578 2924 3579
rect 3014 3583 3020 3584
rect 3014 3579 3015 3583
rect 3019 3579 3020 3583
rect 3014 3578 3020 3579
rect 3118 3583 3124 3584
rect 3118 3579 3119 3583
rect 3123 3579 3124 3583
rect 3118 3578 3124 3579
rect 3222 3583 3228 3584
rect 3222 3579 3223 3583
rect 3227 3579 3228 3583
rect 3222 3578 3228 3579
rect 1862 3573 1868 3574
rect 110 3572 116 3573
rect 110 3568 111 3572
rect 115 3568 116 3572
rect 110 3567 116 3568
rect 1822 3572 1828 3573
rect 1822 3568 1823 3572
rect 1827 3568 1828 3572
rect 1862 3569 1863 3573
rect 1867 3569 1868 3573
rect 1862 3568 1868 3569
rect 3574 3573 3580 3574
rect 3574 3569 3575 3573
rect 3579 3569 3580 3573
rect 3574 3568 3580 3569
rect 1822 3567 1828 3568
rect 1862 3556 1868 3557
rect 110 3555 116 3556
rect 110 3551 111 3555
rect 115 3551 116 3555
rect 110 3550 116 3551
rect 1822 3555 1828 3556
rect 1822 3551 1823 3555
rect 1827 3551 1828 3555
rect 1862 3552 1863 3556
rect 1867 3552 1868 3556
rect 1862 3551 1868 3552
rect 3574 3556 3580 3557
rect 3574 3552 3575 3556
rect 3579 3552 3580 3556
rect 3574 3551 3580 3552
rect 1822 3550 1828 3551
rect 134 3545 140 3546
rect 134 3541 135 3545
rect 139 3541 140 3545
rect 134 3540 140 3541
rect 222 3545 228 3546
rect 222 3541 223 3545
rect 227 3541 228 3545
rect 222 3540 228 3541
rect 310 3545 316 3546
rect 310 3541 311 3545
rect 315 3541 316 3545
rect 310 3540 316 3541
rect 398 3545 404 3546
rect 398 3541 399 3545
rect 403 3541 404 3545
rect 398 3540 404 3541
rect 486 3545 492 3546
rect 486 3541 487 3545
rect 491 3541 492 3545
rect 486 3540 492 3541
rect 1894 3543 1900 3544
rect 1894 3539 1895 3543
rect 1899 3539 1900 3543
rect 1894 3538 1900 3539
rect 1982 3543 1988 3544
rect 1982 3539 1983 3543
rect 1987 3539 1988 3543
rect 1982 3538 1988 3539
rect 2070 3543 2076 3544
rect 2070 3539 2071 3543
rect 2075 3539 2076 3543
rect 2070 3538 2076 3539
rect 2158 3543 2164 3544
rect 2158 3539 2159 3543
rect 2163 3539 2164 3543
rect 2158 3538 2164 3539
rect 2246 3543 2252 3544
rect 2246 3539 2247 3543
rect 2251 3539 2252 3543
rect 2246 3538 2252 3539
rect 2334 3543 2340 3544
rect 2334 3539 2335 3543
rect 2339 3539 2340 3543
rect 2334 3538 2340 3539
rect 2438 3543 2444 3544
rect 2438 3539 2439 3543
rect 2443 3539 2444 3543
rect 2438 3538 2444 3539
rect 2542 3543 2548 3544
rect 2542 3539 2543 3543
rect 2547 3539 2548 3543
rect 2542 3538 2548 3539
rect 2638 3543 2644 3544
rect 2638 3539 2639 3543
rect 2643 3539 2644 3543
rect 2638 3538 2644 3539
rect 2734 3543 2740 3544
rect 2734 3539 2735 3543
rect 2739 3539 2740 3543
rect 2734 3538 2740 3539
rect 2830 3543 2836 3544
rect 2830 3539 2831 3543
rect 2835 3539 2836 3543
rect 2830 3538 2836 3539
rect 2926 3543 2932 3544
rect 2926 3539 2927 3543
rect 2931 3539 2932 3543
rect 2926 3538 2932 3539
rect 3022 3543 3028 3544
rect 3022 3539 3023 3543
rect 3027 3539 3028 3543
rect 3022 3538 3028 3539
rect 3126 3543 3132 3544
rect 3126 3539 3127 3543
rect 3131 3539 3132 3543
rect 3126 3538 3132 3539
rect 3230 3543 3236 3544
rect 3230 3539 3231 3543
rect 3235 3539 3236 3543
rect 3230 3538 3236 3539
rect 246 3523 252 3524
rect 246 3519 247 3523
rect 251 3519 252 3523
rect 246 3518 252 3519
rect 374 3523 380 3524
rect 374 3519 375 3523
rect 379 3519 380 3523
rect 374 3518 380 3519
rect 502 3523 508 3524
rect 502 3519 503 3523
rect 507 3519 508 3523
rect 502 3518 508 3519
rect 622 3523 628 3524
rect 622 3519 623 3523
rect 627 3519 628 3523
rect 622 3518 628 3519
rect 742 3523 748 3524
rect 742 3519 743 3523
rect 747 3519 748 3523
rect 742 3518 748 3519
rect 862 3523 868 3524
rect 862 3519 863 3523
rect 867 3519 868 3523
rect 862 3518 868 3519
rect 974 3523 980 3524
rect 974 3519 975 3523
rect 979 3519 980 3523
rect 974 3518 980 3519
rect 1078 3523 1084 3524
rect 1078 3519 1079 3523
rect 1083 3519 1084 3523
rect 1078 3518 1084 3519
rect 1174 3523 1180 3524
rect 1174 3519 1175 3523
rect 1179 3519 1180 3523
rect 1174 3518 1180 3519
rect 1270 3523 1276 3524
rect 1270 3519 1271 3523
rect 1275 3519 1276 3523
rect 1270 3518 1276 3519
rect 1366 3523 1372 3524
rect 1366 3519 1367 3523
rect 1371 3519 1372 3523
rect 1366 3518 1372 3519
rect 1470 3523 1476 3524
rect 1470 3519 1471 3523
rect 1475 3519 1476 3523
rect 1470 3518 1476 3519
rect 1574 3523 1580 3524
rect 1574 3519 1575 3523
rect 1579 3519 1580 3523
rect 1574 3518 1580 3519
rect 110 3513 116 3514
rect 110 3509 111 3513
rect 115 3509 116 3513
rect 110 3508 116 3509
rect 1822 3513 1828 3514
rect 1822 3509 1823 3513
rect 1827 3509 1828 3513
rect 1822 3508 1828 3509
rect 1894 3509 1900 3510
rect 1894 3505 1895 3509
rect 1899 3505 1900 3509
rect 1894 3504 1900 3505
rect 1982 3509 1988 3510
rect 1982 3505 1983 3509
rect 1987 3505 1988 3509
rect 1982 3504 1988 3505
rect 2102 3509 2108 3510
rect 2102 3505 2103 3509
rect 2107 3505 2108 3509
rect 2102 3504 2108 3505
rect 2230 3509 2236 3510
rect 2230 3505 2231 3509
rect 2235 3505 2236 3509
rect 2230 3504 2236 3505
rect 2366 3509 2372 3510
rect 2366 3505 2367 3509
rect 2371 3505 2372 3509
rect 2366 3504 2372 3505
rect 2510 3509 2516 3510
rect 2510 3505 2511 3509
rect 2515 3505 2516 3509
rect 2510 3504 2516 3505
rect 2654 3509 2660 3510
rect 2654 3505 2655 3509
rect 2659 3505 2660 3509
rect 2654 3504 2660 3505
rect 2790 3509 2796 3510
rect 2790 3505 2791 3509
rect 2795 3505 2796 3509
rect 2790 3504 2796 3505
rect 2934 3509 2940 3510
rect 2934 3505 2935 3509
rect 2939 3505 2940 3509
rect 2934 3504 2940 3505
rect 3078 3509 3084 3510
rect 3078 3505 3079 3509
rect 3083 3505 3084 3509
rect 3078 3504 3084 3505
rect 3222 3509 3228 3510
rect 3222 3505 3223 3509
rect 3227 3505 3228 3509
rect 3222 3504 3228 3505
rect 110 3496 116 3497
rect 110 3492 111 3496
rect 115 3492 116 3496
rect 110 3491 116 3492
rect 1822 3496 1828 3497
rect 1822 3492 1823 3496
rect 1827 3492 1828 3496
rect 1822 3491 1828 3492
rect 1862 3496 1868 3497
rect 1862 3492 1863 3496
rect 1867 3492 1868 3496
rect 1862 3491 1868 3492
rect 3574 3496 3580 3497
rect 3574 3492 3575 3496
rect 3579 3492 3580 3496
rect 3574 3491 3580 3492
rect 254 3483 260 3484
rect 254 3479 255 3483
rect 259 3479 260 3483
rect 254 3478 260 3479
rect 382 3483 388 3484
rect 382 3479 383 3483
rect 387 3479 388 3483
rect 382 3478 388 3479
rect 510 3483 516 3484
rect 510 3479 511 3483
rect 515 3479 516 3483
rect 510 3478 516 3479
rect 630 3483 636 3484
rect 630 3479 631 3483
rect 635 3479 636 3483
rect 630 3478 636 3479
rect 750 3483 756 3484
rect 750 3479 751 3483
rect 755 3479 756 3483
rect 750 3478 756 3479
rect 870 3483 876 3484
rect 870 3479 871 3483
rect 875 3479 876 3483
rect 870 3478 876 3479
rect 982 3483 988 3484
rect 982 3479 983 3483
rect 987 3479 988 3483
rect 982 3478 988 3479
rect 1086 3483 1092 3484
rect 1086 3479 1087 3483
rect 1091 3479 1092 3483
rect 1086 3478 1092 3479
rect 1182 3483 1188 3484
rect 1182 3479 1183 3483
rect 1187 3479 1188 3483
rect 1182 3478 1188 3479
rect 1278 3483 1284 3484
rect 1278 3479 1279 3483
rect 1283 3479 1284 3483
rect 1278 3478 1284 3479
rect 1374 3483 1380 3484
rect 1374 3479 1375 3483
rect 1379 3479 1380 3483
rect 1374 3478 1380 3479
rect 1478 3483 1484 3484
rect 1478 3479 1479 3483
rect 1483 3479 1484 3483
rect 1478 3478 1484 3479
rect 1582 3483 1588 3484
rect 1582 3479 1583 3483
rect 1587 3479 1588 3483
rect 1582 3478 1588 3479
rect 1862 3479 1868 3480
rect 1862 3475 1863 3479
rect 1867 3475 1868 3479
rect 1862 3474 1868 3475
rect 3574 3479 3580 3480
rect 3574 3475 3575 3479
rect 3579 3475 3580 3479
rect 3574 3474 3580 3475
rect 1886 3469 1892 3470
rect 1886 3465 1887 3469
rect 1891 3465 1892 3469
rect 1886 3464 1892 3465
rect 1974 3469 1980 3470
rect 1974 3465 1975 3469
rect 1979 3465 1980 3469
rect 1974 3464 1980 3465
rect 2094 3469 2100 3470
rect 2094 3465 2095 3469
rect 2099 3465 2100 3469
rect 2094 3464 2100 3465
rect 2222 3469 2228 3470
rect 2222 3465 2223 3469
rect 2227 3465 2228 3469
rect 2222 3464 2228 3465
rect 2358 3469 2364 3470
rect 2358 3465 2359 3469
rect 2363 3465 2364 3469
rect 2358 3464 2364 3465
rect 2502 3469 2508 3470
rect 2502 3465 2503 3469
rect 2507 3465 2508 3469
rect 2502 3464 2508 3465
rect 2646 3469 2652 3470
rect 2646 3465 2647 3469
rect 2651 3465 2652 3469
rect 2646 3464 2652 3465
rect 2782 3469 2788 3470
rect 2782 3465 2783 3469
rect 2787 3465 2788 3469
rect 2782 3464 2788 3465
rect 2926 3469 2932 3470
rect 2926 3465 2927 3469
rect 2931 3465 2932 3469
rect 2926 3464 2932 3465
rect 3070 3469 3076 3470
rect 3070 3465 3071 3469
rect 3075 3465 3076 3469
rect 3070 3464 3076 3465
rect 3214 3469 3220 3470
rect 3214 3465 3215 3469
rect 3219 3465 3220 3469
rect 3214 3464 3220 3465
rect 174 3449 180 3450
rect 174 3445 175 3449
rect 179 3445 180 3449
rect 174 3444 180 3445
rect 302 3449 308 3450
rect 302 3445 303 3449
rect 307 3445 308 3449
rect 302 3444 308 3445
rect 446 3449 452 3450
rect 446 3445 447 3449
rect 451 3445 452 3449
rect 446 3444 452 3445
rect 590 3449 596 3450
rect 590 3445 591 3449
rect 595 3445 596 3449
rect 590 3444 596 3445
rect 742 3449 748 3450
rect 742 3445 743 3449
rect 747 3445 748 3449
rect 742 3444 748 3445
rect 894 3449 900 3450
rect 894 3445 895 3449
rect 899 3445 900 3449
rect 894 3444 900 3445
rect 1038 3449 1044 3450
rect 1038 3445 1039 3449
rect 1043 3445 1044 3449
rect 1038 3444 1044 3445
rect 1182 3449 1188 3450
rect 1182 3445 1183 3449
rect 1187 3445 1188 3449
rect 1182 3444 1188 3445
rect 1326 3449 1332 3450
rect 1326 3445 1327 3449
rect 1331 3445 1332 3449
rect 1326 3444 1332 3445
rect 1478 3449 1484 3450
rect 1478 3445 1479 3449
rect 1483 3445 1484 3449
rect 1478 3444 1484 3445
rect 1886 3439 1892 3440
rect 110 3436 116 3437
rect 110 3432 111 3436
rect 115 3432 116 3436
rect 110 3431 116 3432
rect 1822 3436 1828 3437
rect 1822 3432 1823 3436
rect 1827 3432 1828 3436
rect 1886 3435 1887 3439
rect 1891 3435 1892 3439
rect 1886 3434 1892 3435
rect 2022 3439 2028 3440
rect 2022 3435 2023 3439
rect 2027 3435 2028 3439
rect 2022 3434 2028 3435
rect 2190 3439 2196 3440
rect 2190 3435 2191 3439
rect 2195 3435 2196 3439
rect 2190 3434 2196 3435
rect 2366 3439 2372 3440
rect 2366 3435 2367 3439
rect 2371 3435 2372 3439
rect 2366 3434 2372 3435
rect 2542 3439 2548 3440
rect 2542 3435 2543 3439
rect 2547 3435 2548 3439
rect 2542 3434 2548 3435
rect 2710 3439 2716 3440
rect 2710 3435 2711 3439
rect 2715 3435 2716 3439
rect 2710 3434 2716 3435
rect 2870 3439 2876 3440
rect 2870 3435 2871 3439
rect 2875 3435 2876 3439
rect 2870 3434 2876 3435
rect 3030 3439 3036 3440
rect 3030 3435 3031 3439
rect 3035 3435 3036 3439
rect 3030 3434 3036 3435
rect 3190 3439 3196 3440
rect 3190 3435 3191 3439
rect 3195 3435 3196 3439
rect 3190 3434 3196 3435
rect 3358 3439 3364 3440
rect 3358 3435 3359 3439
rect 3363 3435 3364 3439
rect 3358 3434 3364 3435
rect 1822 3431 1828 3432
rect 1862 3429 1868 3430
rect 1862 3425 1863 3429
rect 1867 3425 1868 3429
rect 1862 3424 1868 3425
rect 3574 3429 3580 3430
rect 3574 3425 3575 3429
rect 3579 3425 3580 3429
rect 3574 3424 3580 3425
rect 110 3419 116 3420
rect 110 3415 111 3419
rect 115 3415 116 3419
rect 110 3414 116 3415
rect 1822 3419 1828 3420
rect 1822 3415 1823 3419
rect 1827 3415 1828 3419
rect 1822 3414 1828 3415
rect 1862 3412 1868 3413
rect 166 3409 172 3410
rect 166 3405 167 3409
rect 171 3405 172 3409
rect 166 3404 172 3405
rect 294 3409 300 3410
rect 294 3405 295 3409
rect 299 3405 300 3409
rect 294 3404 300 3405
rect 438 3409 444 3410
rect 438 3405 439 3409
rect 443 3405 444 3409
rect 438 3404 444 3405
rect 582 3409 588 3410
rect 582 3405 583 3409
rect 587 3405 588 3409
rect 582 3404 588 3405
rect 734 3409 740 3410
rect 734 3405 735 3409
rect 739 3405 740 3409
rect 734 3404 740 3405
rect 886 3409 892 3410
rect 886 3405 887 3409
rect 891 3405 892 3409
rect 886 3404 892 3405
rect 1030 3409 1036 3410
rect 1030 3405 1031 3409
rect 1035 3405 1036 3409
rect 1030 3404 1036 3405
rect 1174 3409 1180 3410
rect 1174 3405 1175 3409
rect 1179 3405 1180 3409
rect 1174 3404 1180 3405
rect 1318 3409 1324 3410
rect 1318 3405 1319 3409
rect 1323 3405 1324 3409
rect 1318 3404 1324 3405
rect 1470 3409 1476 3410
rect 1470 3405 1471 3409
rect 1475 3405 1476 3409
rect 1862 3408 1863 3412
rect 1867 3408 1868 3412
rect 1862 3407 1868 3408
rect 3574 3412 3580 3413
rect 3574 3408 3575 3412
rect 3579 3408 3580 3412
rect 3574 3407 3580 3408
rect 1470 3404 1476 3405
rect 1894 3399 1900 3400
rect 1894 3395 1895 3399
rect 1899 3395 1900 3399
rect 1894 3394 1900 3395
rect 2030 3399 2036 3400
rect 2030 3395 2031 3399
rect 2035 3395 2036 3399
rect 2030 3394 2036 3395
rect 2198 3399 2204 3400
rect 2198 3395 2199 3399
rect 2203 3395 2204 3399
rect 2198 3394 2204 3395
rect 2374 3399 2380 3400
rect 2374 3395 2375 3399
rect 2379 3395 2380 3399
rect 2374 3394 2380 3395
rect 2550 3399 2556 3400
rect 2550 3395 2551 3399
rect 2555 3395 2556 3399
rect 2550 3394 2556 3395
rect 2718 3399 2724 3400
rect 2718 3395 2719 3399
rect 2723 3395 2724 3399
rect 2718 3394 2724 3395
rect 2878 3399 2884 3400
rect 2878 3395 2879 3399
rect 2883 3395 2884 3399
rect 2878 3394 2884 3395
rect 3038 3399 3044 3400
rect 3038 3395 3039 3399
rect 3043 3395 3044 3399
rect 3038 3394 3044 3395
rect 3198 3399 3204 3400
rect 3198 3395 3199 3399
rect 3203 3395 3204 3399
rect 3198 3394 3204 3395
rect 3366 3399 3372 3400
rect 3366 3395 3367 3399
rect 3371 3395 3372 3399
rect 3366 3394 3372 3395
rect 134 3387 140 3388
rect 134 3383 135 3387
rect 139 3383 140 3387
rect 134 3382 140 3383
rect 262 3387 268 3388
rect 262 3383 263 3387
rect 267 3383 268 3387
rect 262 3382 268 3383
rect 406 3387 412 3388
rect 406 3383 407 3387
rect 411 3383 412 3387
rect 406 3382 412 3383
rect 566 3387 572 3388
rect 566 3383 567 3387
rect 571 3383 572 3387
rect 566 3382 572 3383
rect 726 3387 732 3388
rect 726 3383 727 3387
rect 731 3383 732 3387
rect 726 3382 732 3383
rect 886 3387 892 3388
rect 886 3383 887 3387
rect 891 3383 892 3387
rect 886 3382 892 3383
rect 1046 3387 1052 3388
rect 1046 3383 1047 3387
rect 1051 3383 1052 3387
rect 1046 3382 1052 3383
rect 1206 3387 1212 3388
rect 1206 3383 1207 3387
rect 1211 3383 1212 3387
rect 1206 3382 1212 3383
rect 1366 3387 1372 3388
rect 1366 3383 1367 3387
rect 1371 3383 1372 3387
rect 1366 3382 1372 3383
rect 1526 3387 1532 3388
rect 1526 3383 1527 3387
rect 1531 3383 1532 3387
rect 1526 3382 1532 3383
rect 110 3377 116 3378
rect 110 3373 111 3377
rect 115 3373 116 3377
rect 110 3372 116 3373
rect 1822 3377 1828 3378
rect 1822 3373 1823 3377
rect 1827 3373 1828 3377
rect 1822 3372 1828 3373
rect 110 3360 116 3361
rect 110 3356 111 3360
rect 115 3356 116 3360
rect 110 3355 116 3356
rect 1822 3360 1828 3361
rect 1822 3356 1823 3360
rect 1827 3356 1828 3360
rect 1822 3355 1828 3356
rect 1894 3357 1900 3358
rect 1894 3353 1895 3357
rect 1899 3353 1900 3357
rect 1894 3352 1900 3353
rect 2030 3357 2036 3358
rect 2030 3353 2031 3357
rect 2035 3353 2036 3357
rect 2030 3352 2036 3353
rect 2198 3357 2204 3358
rect 2198 3353 2199 3357
rect 2203 3353 2204 3357
rect 2198 3352 2204 3353
rect 2374 3357 2380 3358
rect 2374 3353 2375 3357
rect 2379 3353 2380 3357
rect 2374 3352 2380 3353
rect 2550 3357 2556 3358
rect 2550 3353 2551 3357
rect 2555 3353 2556 3357
rect 2550 3352 2556 3353
rect 2718 3357 2724 3358
rect 2718 3353 2719 3357
rect 2723 3353 2724 3357
rect 2718 3352 2724 3353
rect 2878 3357 2884 3358
rect 2878 3353 2879 3357
rect 2883 3353 2884 3357
rect 2878 3352 2884 3353
rect 3038 3357 3044 3358
rect 3038 3353 3039 3357
rect 3043 3353 3044 3357
rect 3038 3352 3044 3353
rect 3190 3357 3196 3358
rect 3190 3353 3191 3357
rect 3195 3353 3196 3357
rect 3190 3352 3196 3353
rect 3342 3357 3348 3358
rect 3342 3353 3343 3357
rect 3347 3353 3348 3357
rect 3342 3352 3348 3353
rect 3486 3357 3492 3358
rect 3486 3353 3487 3357
rect 3491 3353 3492 3357
rect 3486 3352 3492 3353
rect 142 3347 148 3348
rect 142 3343 143 3347
rect 147 3343 148 3347
rect 142 3342 148 3343
rect 270 3347 276 3348
rect 270 3343 271 3347
rect 275 3343 276 3347
rect 270 3342 276 3343
rect 414 3347 420 3348
rect 414 3343 415 3347
rect 419 3343 420 3347
rect 414 3342 420 3343
rect 574 3347 580 3348
rect 574 3343 575 3347
rect 579 3343 580 3347
rect 574 3342 580 3343
rect 734 3347 740 3348
rect 734 3343 735 3347
rect 739 3343 740 3347
rect 734 3342 740 3343
rect 894 3347 900 3348
rect 894 3343 895 3347
rect 899 3343 900 3347
rect 894 3342 900 3343
rect 1054 3347 1060 3348
rect 1054 3343 1055 3347
rect 1059 3343 1060 3347
rect 1054 3342 1060 3343
rect 1214 3347 1220 3348
rect 1214 3343 1215 3347
rect 1219 3343 1220 3347
rect 1214 3342 1220 3343
rect 1374 3347 1380 3348
rect 1374 3343 1375 3347
rect 1379 3343 1380 3347
rect 1374 3342 1380 3343
rect 1534 3347 1540 3348
rect 1534 3343 1535 3347
rect 1539 3343 1540 3347
rect 1534 3342 1540 3343
rect 1862 3344 1868 3345
rect 1862 3340 1863 3344
rect 1867 3340 1868 3344
rect 1862 3339 1868 3340
rect 3574 3344 3580 3345
rect 3574 3340 3575 3344
rect 3579 3340 3580 3344
rect 3574 3339 3580 3340
rect 1862 3327 1868 3328
rect 1862 3323 1863 3327
rect 1867 3323 1868 3327
rect 1862 3322 1868 3323
rect 3574 3327 3580 3328
rect 3574 3323 3575 3327
rect 3579 3323 3580 3327
rect 3574 3322 3580 3323
rect 1886 3317 1892 3318
rect 1886 3313 1887 3317
rect 1891 3313 1892 3317
rect 1886 3312 1892 3313
rect 2022 3317 2028 3318
rect 2022 3313 2023 3317
rect 2027 3313 2028 3317
rect 2022 3312 2028 3313
rect 2190 3317 2196 3318
rect 2190 3313 2191 3317
rect 2195 3313 2196 3317
rect 2190 3312 2196 3313
rect 2366 3317 2372 3318
rect 2366 3313 2367 3317
rect 2371 3313 2372 3317
rect 2366 3312 2372 3313
rect 2542 3317 2548 3318
rect 2542 3313 2543 3317
rect 2547 3313 2548 3317
rect 2542 3312 2548 3313
rect 2710 3317 2716 3318
rect 2710 3313 2711 3317
rect 2715 3313 2716 3317
rect 2710 3312 2716 3313
rect 2870 3317 2876 3318
rect 2870 3313 2871 3317
rect 2875 3313 2876 3317
rect 2870 3312 2876 3313
rect 3030 3317 3036 3318
rect 3030 3313 3031 3317
rect 3035 3313 3036 3317
rect 3030 3312 3036 3313
rect 3182 3317 3188 3318
rect 3182 3313 3183 3317
rect 3187 3313 3188 3317
rect 3182 3312 3188 3313
rect 3334 3317 3340 3318
rect 3334 3313 3335 3317
rect 3339 3313 3340 3317
rect 3334 3312 3340 3313
rect 3478 3317 3484 3318
rect 3478 3313 3479 3317
rect 3483 3313 3484 3317
rect 3478 3312 3484 3313
rect 206 3309 212 3310
rect 206 3305 207 3309
rect 211 3305 212 3309
rect 206 3304 212 3305
rect 334 3309 340 3310
rect 334 3305 335 3309
rect 339 3305 340 3309
rect 334 3304 340 3305
rect 478 3309 484 3310
rect 478 3305 479 3309
rect 483 3305 484 3309
rect 478 3304 484 3305
rect 638 3309 644 3310
rect 638 3305 639 3309
rect 643 3305 644 3309
rect 638 3304 644 3305
rect 806 3309 812 3310
rect 806 3305 807 3309
rect 811 3305 812 3309
rect 806 3304 812 3305
rect 982 3309 988 3310
rect 982 3305 983 3309
rect 987 3305 988 3309
rect 982 3304 988 3305
rect 1166 3309 1172 3310
rect 1166 3305 1167 3309
rect 1171 3305 1172 3309
rect 1166 3304 1172 3305
rect 1350 3309 1356 3310
rect 1350 3305 1351 3309
rect 1355 3305 1356 3309
rect 1350 3304 1356 3305
rect 1542 3309 1548 3310
rect 1542 3305 1543 3309
rect 1547 3305 1548 3309
rect 1542 3304 1548 3305
rect 110 3296 116 3297
rect 110 3292 111 3296
rect 115 3292 116 3296
rect 110 3291 116 3292
rect 1822 3296 1828 3297
rect 1822 3292 1823 3296
rect 1827 3292 1828 3296
rect 1822 3291 1828 3292
rect 1886 3295 1892 3296
rect 1886 3291 1887 3295
rect 1891 3291 1892 3295
rect 1886 3290 1892 3291
rect 2006 3295 2012 3296
rect 2006 3291 2007 3295
rect 2011 3291 2012 3295
rect 2006 3290 2012 3291
rect 2150 3295 2156 3296
rect 2150 3291 2151 3295
rect 2155 3291 2156 3295
rect 2150 3290 2156 3291
rect 2302 3295 2308 3296
rect 2302 3291 2303 3295
rect 2307 3291 2308 3295
rect 2302 3290 2308 3291
rect 2462 3295 2468 3296
rect 2462 3291 2463 3295
rect 2467 3291 2468 3295
rect 2462 3290 2468 3291
rect 2630 3295 2636 3296
rect 2630 3291 2631 3295
rect 2635 3291 2636 3295
rect 2630 3290 2636 3291
rect 2798 3295 2804 3296
rect 2798 3291 2799 3295
rect 2803 3291 2804 3295
rect 2798 3290 2804 3291
rect 2966 3295 2972 3296
rect 2966 3291 2967 3295
rect 2971 3291 2972 3295
rect 2966 3290 2972 3291
rect 3134 3295 3140 3296
rect 3134 3291 3135 3295
rect 3139 3291 3140 3295
rect 3134 3290 3140 3291
rect 3310 3295 3316 3296
rect 3310 3291 3311 3295
rect 3315 3291 3316 3295
rect 3310 3290 3316 3291
rect 3478 3295 3484 3296
rect 3478 3291 3479 3295
rect 3483 3291 3484 3295
rect 3478 3290 3484 3291
rect 1862 3285 1868 3286
rect 1862 3281 1863 3285
rect 1867 3281 1868 3285
rect 1862 3280 1868 3281
rect 3574 3285 3580 3286
rect 3574 3281 3575 3285
rect 3579 3281 3580 3285
rect 3574 3280 3580 3281
rect 110 3279 116 3280
rect 110 3275 111 3279
rect 115 3275 116 3279
rect 110 3274 116 3275
rect 1822 3279 1828 3280
rect 1822 3275 1823 3279
rect 1827 3275 1828 3279
rect 1822 3274 1828 3275
rect 198 3269 204 3270
rect 198 3265 199 3269
rect 203 3265 204 3269
rect 198 3264 204 3265
rect 326 3269 332 3270
rect 326 3265 327 3269
rect 331 3265 332 3269
rect 326 3264 332 3265
rect 470 3269 476 3270
rect 470 3265 471 3269
rect 475 3265 476 3269
rect 470 3264 476 3265
rect 630 3269 636 3270
rect 630 3265 631 3269
rect 635 3265 636 3269
rect 630 3264 636 3265
rect 798 3269 804 3270
rect 798 3265 799 3269
rect 803 3265 804 3269
rect 798 3264 804 3265
rect 974 3269 980 3270
rect 974 3265 975 3269
rect 979 3265 980 3269
rect 974 3264 980 3265
rect 1158 3269 1164 3270
rect 1158 3265 1159 3269
rect 1163 3265 1164 3269
rect 1158 3264 1164 3265
rect 1342 3269 1348 3270
rect 1342 3265 1343 3269
rect 1347 3265 1348 3269
rect 1342 3264 1348 3265
rect 1534 3269 1540 3270
rect 1534 3265 1535 3269
rect 1539 3265 1540 3269
rect 1534 3264 1540 3265
rect 1862 3268 1868 3269
rect 1862 3264 1863 3268
rect 1867 3264 1868 3268
rect 1862 3263 1868 3264
rect 3574 3268 3580 3269
rect 3574 3264 3575 3268
rect 3579 3264 3580 3268
rect 3574 3263 3580 3264
rect 1894 3255 1900 3256
rect 1894 3251 1895 3255
rect 1899 3251 1900 3255
rect 1894 3250 1900 3251
rect 2014 3255 2020 3256
rect 2014 3251 2015 3255
rect 2019 3251 2020 3255
rect 2014 3250 2020 3251
rect 2158 3255 2164 3256
rect 2158 3251 2159 3255
rect 2163 3251 2164 3255
rect 2158 3250 2164 3251
rect 2310 3255 2316 3256
rect 2310 3251 2311 3255
rect 2315 3251 2316 3255
rect 2310 3250 2316 3251
rect 2470 3255 2476 3256
rect 2470 3251 2471 3255
rect 2475 3251 2476 3255
rect 2470 3250 2476 3251
rect 2638 3255 2644 3256
rect 2638 3251 2639 3255
rect 2643 3251 2644 3255
rect 2638 3250 2644 3251
rect 2806 3255 2812 3256
rect 2806 3251 2807 3255
rect 2811 3251 2812 3255
rect 2806 3250 2812 3251
rect 2974 3255 2980 3256
rect 2974 3251 2975 3255
rect 2979 3251 2980 3255
rect 2974 3250 2980 3251
rect 3142 3255 3148 3256
rect 3142 3251 3143 3255
rect 3147 3251 3148 3255
rect 3142 3250 3148 3251
rect 3318 3255 3324 3256
rect 3318 3251 3319 3255
rect 3323 3251 3324 3255
rect 3318 3250 3324 3251
rect 3486 3255 3492 3256
rect 3486 3251 3487 3255
rect 3491 3251 3492 3255
rect 3486 3250 3492 3251
rect 366 3243 372 3244
rect 366 3239 367 3243
rect 371 3239 372 3243
rect 366 3238 372 3239
rect 502 3243 508 3244
rect 502 3239 503 3243
rect 507 3239 508 3243
rect 502 3238 508 3239
rect 638 3243 644 3244
rect 638 3239 639 3243
rect 643 3239 644 3243
rect 638 3238 644 3239
rect 782 3243 788 3244
rect 782 3239 783 3243
rect 787 3239 788 3243
rect 782 3238 788 3239
rect 934 3243 940 3244
rect 934 3239 935 3243
rect 939 3239 940 3243
rect 934 3238 940 3239
rect 1094 3243 1100 3244
rect 1094 3239 1095 3243
rect 1099 3239 1100 3243
rect 1094 3238 1100 3239
rect 1254 3243 1260 3244
rect 1254 3239 1255 3243
rect 1259 3239 1260 3243
rect 1254 3238 1260 3239
rect 1414 3243 1420 3244
rect 1414 3239 1415 3243
rect 1419 3239 1420 3243
rect 1414 3238 1420 3239
rect 1574 3243 1580 3244
rect 1574 3239 1575 3243
rect 1579 3239 1580 3243
rect 1574 3238 1580 3239
rect 110 3233 116 3234
rect 110 3229 111 3233
rect 115 3229 116 3233
rect 110 3228 116 3229
rect 1822 3233 1828 3234
rect 1822 3229 1823 3233
rect 1827 3229 1828 3233
rect 1822 3228 1828 3229
rect 110 3216 116 3217
rect 110 3212 111 3216
rect 115 3212 116 3216
rect 110 3211 116 3212
rect 1822 3216 1828 3217
rect 1822 3212 1823 3216
rect 1827 3212 1828 3216
rect 1822 3211 1828 3212
rect 1894 3213 1900 3214
rect 1894 3209 1895 3213
rect 1899 3209 1900 3213
rect 1894 3208 1900 3209
rect 2022 3213 2028 3214
rect 2022 3209 2023 3213
rect 2027 3209 2028 3213
rect 2022 3208 2028 3209
rect 2174 3213 2180 3214
rect 2174 3209 2175 3213
rect 2179 3209 2180 3213
rect 2174 3208 2180 3209
rect 2326 3213 2332 3214
rect 2326 3209 2327 3213
rect 2331 3209 2332 3213
rect 2326 3208 2332 3209
rect 2462 3213 2468 3214
rect 2462 3209 2463 3213
rect 2467 3209 2468 3213
rect 2462 3208 2468 3209
rect 2598 3213 2604 3214
rect 2598 3209 2599 3213
rect 2603 3209 2604 3213
rect 2598 3208 2604 3209
rect 2734 3213 2740 3214
rect 2734 3209 2735 3213
rect 2739 3209 2740 3213
rect 2734 3208 2740 3209
rect 2870 3213 2876 3214
rect 2870 3209 2871 3213
rect 2875 3209 2876 3213
rect 2870 3208 2876 3209
rect 3014 3213 3020 3214
rect 3014 3209 3015 3213
rect 3019 3209 3020 3213
rect 3014 3208 3020 3209
rect 3166 3213 3172 3214
rect 3166 3209 3167 3213
rect 3171 3209 3172 3213
rect 3166 3208 3172 3209
rect 3326 3213 3332 3214
rect 3326 3209 3327 3213
rect 3331 3209 3332 3213
rect 3326 3208 3332 3209
rect 3486 3213 3492 3214
rect 3486 3209 3487 3213
rect 3491 3209 3492 3213
rect 3486 3208 3492 3209
rect 374 3203 380 3204
rect 374 3199 375 3203
rect 379 3199 380 3203
rect 374 3198 380 3199
rect 510 3203 516 3204
rect 510 3199 511 3203
rect 515 3199 516 3203
rect 510 3198 516 3199
rect 646 3203 652 3204
rect 646 3199 647 3203
rect 651 3199 652 3203
rect 646 3198 652 3199
rect 790 3203 796 3204
rect 790 3199 791 3203
rect 795 3199 796 3203
rect 790 3198 796 3199
rect 942 3203 948 3204
rect 942 3199 943 3203
rect 947 3199 948 3203
rect 942 3198 948 3199
rect 1102 3203 1108 3204
rect 1102 3199 1103 3203
rect 1107 3199 1108 3203
rect 1102 3198 1108 3199
rect 1262 3203 1268 3204
rect 1262 3199 1263 3203
rect 1267 3199 1268 3203
rect 1262 3198 1268 3199
rect 1422 3203 1428 3204
rect 1422 3199 1423 3203
rect 1427 3199 1428 3203
rect 1422 3198 1428 3199
rect 1582 3203 1588 3204
rect 1582 3199 1583 3203
rect 1587 3199 1588 3203
rect 1582 3198 1588 3199
rect 1862 3200 1868 3201
rect 1862 3196 1863 3200
rect 1867 3196 1868 3200
rect 1862 3195 1868 3196
rect 3574 3200 3580 3201
rect 3574 3196 3575 3200
rect 3579 3196 3580 3200
rect 3574 3195 3580 3196
rect 1862 3183 1868 3184
rect 1862 3179 1863 3183
rect 1867 3179 1868 3183
rect 1862 3178 1868 3179
rect 3574 3183 3580 3184
rect 3574 3179 3575 3183
rect 3579 3179 3580 3183
rect 3574 3178 3580 3179
rect 1886 3173 1892 3174
rect 1886 3169 1887 3173
rect 1891 3169 1892 3173
rect 1886 3168 1892 3169
rect 2014 3173 2020 3174
rect 2014 3169 2015 3173
rect 2019 3169 2020 3173
rect 2014 3168 2020 3169
rect 2166 3173 2172 3174
rect 2166 3169 2167 3173
rect 2171 3169 2172 3173
rect 2166 3168 2172 3169
rect 2318 3173 2324 3174
rect 2318 3169 2319 3173
rect 2323 3169 2324 3173
rect 2318 3168 2324 3169
rect 2454 3173 2460 3174
rect 2454 3169 2455 3173
rect 2459 3169 2460 3173
rect 2454 3168 2460 3169
rect 2590 3173 2596 3174
rect 2590 3169 2591 3173
rect 2595 3169 2596 3173
rect 2590 3168 2596 3169
rect 2726 3173 2732 3174
rect 2726 3169 2727 3173
rect 2731 3169 2732 3173
rect 2726 3168 2732 3169
rect 2862 3173 2868 3174
rect 2862 3169 2863 3173
rect 2867 3169 2868 3173
rect 2862 3168 2868 3169
rect 3006 3173 3012 3174
rect 3006 3169 3007 3173
rect 3011 3169 3012 3173
rect 3006 3168 3012 3169
rect 3158 3173 3164 3174
rect 3158 3169 3159 3173
rect 3163 3169 3164 3173
rect 3158 3168 3164 3169
rect 3318 3173 3324 3174
rect 3318 3169 3319 3173
rect 3323 3169 3324 3173
rect 3318 3168 3324 3169
rect 3478 3173 3484 3174
rect 3478 3169 3479 3173
rect 3483 3169 3484 3173
rect 3478 3168 3484 3169
rect 446 3161 452 3162
rect 446 3157 447 3161
rect 451 3157 452 3161
rect 446 3156 452 3157
rect 558 3161 564 3162
rect 558 3157 559 3161
rect 563 3157 564 3161
rect 558 3156 564 3157
rect 686 3161 692 3162
rect 686 3157 687 3161
rect 691 3157 692 3161
rect 686 3156 692 3157
rect 822 3161 828 3162
rect 822 3157 823 3161
rect 827 3157 828 3161
rect 822 3156 828 3157
rect 974 3161 980 3162
rect 974 3157 975 3161
rect 979 3157 980 3161
rect 974 3156 980 3157
rect 1134 3161 1140 3162
rect 1134 3157 1135 3161
rect 1139 3157 1140 3161
rect 1134 3156 1140 3157
rect 1294 3161 1300 3162
rect 1294 3157 1295 3161
rect 1299 3157 1300 3161
rect 1294 3156 1300 3157
rect 1462 3161 1468 3162
rect 1462 3157 1463 3161
rect 1467 3157 1468 3161
rect 1462 3156 1468 3157
rect 1638 3161 1644 3162
rect 1638 3157 1639 3161
rect 1643 3157 1644 3161
rect 1638 3156 1644 3157
rect 110 3148 116 3149
rect 110 3144 111 3148
rect 115 3144 116 3148
rect 110 3143 116 3144
rect 1822 3148 1828 3149
rect 1822 3144 1823 3148
rect 1827 3144 1828 3148
rect 1822 3143 1828 3144
rect 1886 3147 1892 3148
rect 1886 3143 1887 3147
rect 1891 3143 1892 3147
rect 1886 3142 1892 3143
rect 2046 3147 2052 3148
rect 2046 3143 2047 3147
rect 2051 3143 2052 3147
rect 2046 3142 2052 3143
rect 2198 3147 2204 3148
rect 2198 3143 2199 3147
rect 2203 3143 2204 3147
rect 2198 3142 2204 3143
rect 2350 3147 2356 3148
rect 2350 3143 2351 3147
rect 2355 3143 2356 3147
rect 2350 3142 2356 3143
rect 2510 3147 2516 3148
rect 2510 3143 2511 3147
rect 2515 3143 2516 3147
rect 2510 3142 2516 3143
rect 2678 3147 2684 3148
rect 2678 3143 2679 3147
rect 2683 3143 2684 3147
rect 2678 3142 2684 3143
rect 2870 3147 2876 3148
rect 2870 3143 2871 3147
rect 2875 3143 2876 3147
rect 2870 3142 2876 3143
rect 3070 3147 3076 3148
rect 3070 3143 3071 3147
rect 3075 3143 3076 3147
rect 3070 3142 3076 3143
rect 3286 3147 3292 3148
rect 3286 3143 3287 3147
rect 3291 3143 3292 3147
rect 3286 3142 3292 3143
rect 3478 3147 3484 3148
rect 3478 3143 3479 3147
rect 3483 3143 3484 3147
rect 3478 3142 3484 3143
rect 1862 3137 1868 3138
rect 1862 3133 1863 3137
rect 1867 3133 1868 3137
rect 1862 3132 1868 3133
rect 3574 3137 3580 3138
rect 3574 3133 3575 3137
rect 3579 3133 3580 3137
rect 3574 3132 3580 3133
rect 110 3131 116 3132
rect 110 3127 111 3131
rect 115 3127 116 3131
rect 110 3126 116 3127
rect 1822 3131 1828 3132
rect 1822 3127 1823 3131
rect 1827 3127 1828 3131
rect 1822 3126 1828 3127
rect 438 3121 444 3122
rect 438 3117 439 3121
rect 443 3117 444 3121
rect 438 3116 444 3117
rect 550 3121 556 3122
rect 550 3117 551 3121
rect 555 3117 556 3121
rect 550 3116 556 3117
rect 678 3121 684 3122
rect 678 3117 679 3121
rect 683 3117 684 3121
rect 678 3116 684 3117
rect 814 3121 820 3122
rect 814 3117 815 3121
rect 819 3117 820 3121
rect 814 3116 820 3117
rect 966 3121 972 3122
rect 966 3117 967 3121
rect 971 3117 972 3121
rect 966 3116 972 3117
rect 1126 3121 1132 3122
rect 1126 3117 1127 3121
rect 1131 3117 1132 3121
rect 1126 3116 1132 3117
rect 1286 3121 1292 3122
rect 1286 3117 1287 3121
rect 1291 3117 1292 3121
rect 1286 3116 1292 3117
rect 1454 3121 1460 3122
rect 1454 3117 1455 3121
rect 1459 3117 1460 3121
rect 1454 3116 1460 3117
rect 1630 3121 1636 3122
rect 1630 3117 1631 3121
rect 1635 3117 1636 3121
rect 1630 3116 1636 3117
rect 1862 3120 1868 3121
rect 1862 3116 1863 3120
rect 1867 3116 1868 3120
rect 1862 3115 1868 3116
rect 3574 3120 3580 3121
rect 3574 3116 3575 3120
rect 3579 3116 3580 3120
rect 3574 3115 3580 3116
rect 1894 3107 1900 3108
rect 1894 3103 1895 3107
rect 1899 3103 1900 3107
rect 1894 3102 1900 3103
rect 2054 3107 2060 3108
rect 2054 3103 2055 3107
rect 2059 3103 2060 3107
rect 2054 3102 2060 3103
rect 2206 3107 2212 3108
rect 2206 3103 2207 3107
rect 2211 3103 2212 3107
rect 2206 3102 2212 3103
rect 2358 3107 2364 3108
rect 2358 3103 2359 3107
rect 2363 3103 2364 3107
rect 2358 3102 2364 3103
rect 2518 3107 2524 3108
rect 2518 3103 2519 3107
rect 2523 3103 2524 3107
rect 2518 3102 2524 3103
rect 2686 3107 2692 3108
rect 2686 3103 2687 3107
rect 2691 3103 2692 3107
rect 2686 3102 2692 3103
rect 2878 3107 2884 3108
rect 2878 3103 2879 3107
rect 2883 3103 2884 3107
rect 2878 3102 2884 3103
rect 3078 3107 3084 3108
rect 3078 3103 3079 3107
rect 3083 3103 3084 3107
rect 3078 3102 3084 3103
rect 3294 3107 3300 3108
rect 3294 3103 3295 3107
rect 3299 3103 3300 3107
rect 3294 3102 3300 3103
rect 3486 3107 3492 3108
rect 3486 3103 3487 3107
rect 3491 3103 3492 3107
rect 3486 3102 3492 3103
rect 550 3091 556 3092
rect 550 3087 551 3091
rect 555 3087 556 3091
rect 550 3086 556 3087
rect 662 3091 668 3092
rect 662 3087 663 3091
rect 667 3087 668 3091
rect 662 3086 668 3087
rect 782 3091 788 3092
rect 782 3087 783 3091
rect 787 3087 788 3091
rect 782 3086 788 3087
rect 902 3091 908 3092
rect 902 3087 903 3091
rect 907 3087 908 3091
rect 902 3086 908 3087
rect 1030 3091 1036 3092
rect 1030 3087 1031 3091
rect 1035 3087 1036 3091
rect 1030 3086 1036 3087
rect 1158 3091 1164 3092
rect 1158 3087 1159 3091
rect 1163 3087 1164 3091
rect 1158 3086 1164 3087
rect 1286 3091 1292 3092
rect 1286 3087 1287 3091
rect 1291 3087 1292 3091
rect 1286 3086 1292 3087
rect 1422 3091 1428 3092
rect 1422 3087 1423 3091
rect 1427 3087 1428 3091
rect 1422 3086 1428 3087
rect 1558 3091 1564 3092
rect 1558 3087 1559 3091
rect 1563 3087 1564 3091
rect 1558 3086 1564 3087
rect 1694 3091 1700 3092
rect 1694 3087 1695 3091
rect 1699 3087 1700 3091
rect 1694 3086 1700 3087
rect 110 3081 116 3082
rect 110 3077 111 3081
rect 115 3077 116 3081
rect 110 3076 116 3077
rect 1822 3081 1828 3082
rect 1822 3077 1823 3081
rect 1827 3077 1828 3081
rect 1822 3076 1828 3077
rect 1918 3065 1924 3066
rect 110 3064 116 3065
rect 110 3060 111 3064
rect 115 3060 116 3064
rect 110 3059 116 3060
rect 1822 3064 1828 3065
rect 1822 3060 1823 3064
rect 1827 3060 1828 3064
rect 1918 3061 1919 3065
rect 1923 3061 1924 3065
rect 1918 3060 1924 3061
rect 2086 3065 2092 3066
rect 2086 3061 2087 3065
rect 2091 3061 2092 3065
rect 2086 3060 2092 3061
rect 2278 3065 2284 3066
rect 2278 3061 2279 3065
rect 2283 3061 2284 3065
rect 2278 3060 2284 3061
rect 2486 3065 2492 3066
rect 2486 3061 2487 3065
rect 2491 3061 2492 3065
rect 2486 3060 2492 3061
rect 2718 3065 2724 3066
rect 2718 3061 2719 3065
rect 2723 3061 2724 3065
rect 2718 3060 2724 3061
rect 2974 3065 2980 3066
rect 2974 3061 2975 3065
rect 2979 3061 2980 3065
rect 2974 3060 2980 3061
rect 3238 3065 3244 3066
rect 3238 3061 3239 3065
rect 3243 3061 3244 3065
rect 3238 3060 3244 3061
rect 3486 3065 3492 3066
rect 3486 3061 3487 3065
rect 3491 3061 3492 3065
rect 3486 3060 3492 3061
rect 1822 3059 1828 3060
rect 1862 3052 1868 3053
rect 558 3051 564 3052
rect 558 3047 559 3051
rect 563 3047 564 3051
rect 558 3046 564 3047
rect 670 3051 676 3052
rect 670 3047 671 3051
rect 675 3047 676 3051
rect 670 3046 676 3047
rect 790 3051 796 3052
rect 790 3047 791 3051
rect 795 3047 796 3051
rect 790 3046 796 3047
rect 910 3051 916 3052
rect 910 3047 911 3051
rect 915 3047 916 3051
rect 910 3046 916 3047
rect 1038 3051 1044 3052
rect 1038 3047 1039 3051
rect 1043 3047 1044 3051
rect 1038 3046 1044 3047
rect 1166 3051 1172 3052
rect 1166 3047 1167 3051
rect 1171 3047 1172 3051
rect 1166 3046 1172 3047
rect 1294 3051 1300 3052
rect 1294 3047 1295 3051
rect 1299 3047 1300 3051
rect 1294 3046 1300 3047
rect 1430 3051 1436 3052
rect 1430 3047 1431 3051
rect 1435 3047 1436 3051
rect 1430 3046 1436 3047
rect 1566 3051 1572 3052
rect 1566 3047 1567 3051
rect 1571 3047 1572 3051
rect 1566 3046 1572 3047
rect 1702 3051 1708 3052
rect 1702 3047 1703 3051
rect 1707 3047 1708 3051
rect 1862 3048 1863 3052
rect 1867 3048 1868 3052
rect 1862 3047 1868 3048
rect 3574 3052 3580 3053
rect 3574 3048 3575 3052
rect 3579 3048 3580 3052
rect 3574 3047 3580 3048
rect 1702 3046 1708 3047
rect 1862 3035 1868 3036
rect 1862 3031 1863 3035
rect 1867 3031 1868 3035
rect 1862 3030 1868 3031
rect 3574 3035 3580 3036
rect 3574 3031 3575 3035
rect 3579 3031 3580 3035
rect 3574 3030 3580 3031
rect 1910 3025 1916 3026
rect 1910 3021 1911 3025
rect 1915 3021 1916 3025
rect 1910 3020 1916 3021
rect 2078 3025 2084 3026
rect 2078 3021 2079 3025
rect 2083 3021 2084 3025
rect 2078 3020 2084 3021
rect 2270 3025 2276 3026
rect 2270 3021 2271 3025
rect 2275 3021 2276 3025
rect 2270 3020 2276 3021
rect 2478 3025 2484 3026
rect 2478 3021 2479 3025
rect 2483 3021 2484 3025
rect 2478 3020 2484 3021
rect 2710 3025 2716 3026
rect 2710 3021 2711 3025
rect 2715 3021 2716 3025
rect 2710 3020 2716 3021
rect 2966 3025 2972 3026
rect 2966 3021 2967 3025
rect 2971 3021 2972 3025
rect 2966 3020 2972 3021
rect 3230 3025 3236 3026
rect 3230 3021 3231 3025
rect 3235 3021 3236 3025
rect 3230 3020 3236 3021
rect 3478 3025 3484 3026
rect 3478 3021 3479 3025
rect 3483 3021 3484 3025
rect 3478 3020 3484 3021
rect 574 3013 580 3014
rect 574 3009 575 3013
rect 579 3009 580 3013
rect 574 3008 580 3009
rect 702 3013 708 3014
rect 702 3009 703 3013
rect 707 3009 708 3013
rect 702 3008 708 3009
rect 830 3013 836 3014
rect 830 3009 831 3013
rect 835 3009 836 3013
rect 830 3008 836 3009
rect 966 3013 972 3014
rect 966 3009 967 3013
rect 971 3009 972 3013
rect 966 3008 972 3009
rect 1102 3013 1108 3014
rect 1102 3009 1103 3013
rect 1107 3009 1108 3013
rect 1102 3008 1108 3009
rect 1238 3013 1244 3014
rect 1238 3009 1239 3013
rect 1243 3009 1244 3013
rect 1238 3008 1244 3009
rect 1366 3013 1372 3014
rect 1366 3009 1367 3013
rect 1371 3009 1372 3013
rect 1366 3008 1372 3009
rect 1494 3013 1500 3014
rect 1494 3009 1495 3013
rect 1499 3009 1500 3013
rect 1494 3008 1500 3009
rect 1622 3013 1628 3014
rect 1622 3009 1623 3013
rect 1627 3009 1628 3013
rect 1622 3008 1628 3009
rect 1734 3013 1740 3014
rect 1734 3009 1735 3013
rect 1739 3009 1740 3013
rect 1734 3008 1740 3009
rect 110 3000 116 3001
rect 110 2996 111 3000
rect 115 2996 116 3000
rect 110 2995 116 2996
rect 1822 3000 1828 3001
rect 1822 2996 1823 3000
rect 1827 2996 1828 3000
rect 1822 2995 1828 2996
rect 2022 2999 2028 3000
rect 2022 2995 2023 2999
rect 2027 2995 2028 2999
rect 2022 2994 2028 2995
rect 2158 2999 2164 3000
rect 2158 2995 2159 2999
rect 2163 2995 2164 2999
rect 2158 2994 2164 2995
rect 2286 2999 2292 3000
rect 2286 2995 2287 2999
rect 2291 2995 2292 2999
rect 2286 2994 2292 2995
rect 2414 2999 2420 3000
rect 2414 2995 2415 2999
rect 2419 2995 2420 2999
rect 2414 2994 2420 2995
rect 2534 2999 2540 3000
rect 2534 2995 2535 2999
rect 2539 2995 2540 2999
rect 2534 2994 2540 2995
rect 2662 2999 2668 3000
rect 2662 2995 2663 2999
rect 2667 2995 2668 2999
rect 2662 2994 2668 2995
rect 2806 2999 2812 3000
rect 2806 2995 2807 2999
rect 2811 2995 2812 2999
rect 2806 2994 2812 2995
rect 2966 2999 2972 3000
rect 2966 2995 2967 2999
rect 2971 2995 2972 2999
rect 2966 2994 2972 2995
rect 3142 2999 3148 3000
rect 3142 2995 3143 2999
rect 3147 2995 3148 2999
rect 3142 2994 3148 2995
rect 3318 2999 3324 3000
rect 3318 2995 3319 2999
rect 3323 2995 3324 2999
rect 3318 2994 3324 2995
rect 3478 2999 3484 3000
rect 3478 2995 3479 2999
rect 3483 2995 3484 2999
rect 3478 2994 3484 2995
rect 1862 2989 1868 2990
rect 1862 2985 1863 2989
rect 1867 2985 1868 2989
rect 1862 2984 1868 2985
rect 3574 2989 3580 2990
rect 3574 2985 3575 2989
rect 3579 2985 3580 2989
rect 3574 2984 3580 2985
rect 110 2983 116 2984
rect 110 2979 111 2983
rect 115 2979 116 2983
rect 110 2978 116 2979
rect 1822 2983 1828 2984
rect 1822 2979 1823 2983
rect 1827 2979 1828 2983
rect 1822 2978 1828 2979
rect 566 2973 572 2974
rect 566 2969 567 2973
rect 571 2969 572 2973
rect 566 2968 572 2969
rect 694 2973 700 2974
rect 694 2969 695 2973
rect 699 2969 700 2973
rect 694 2968 700 2969
rect 822 2973 828 2974
rect 822 2969 823 2973
rect 827 2969 828 2973
rect 822 2968 828 2969
rect 958 2973 964 2974
rect 958 2969 959 2973
rect 963 2969 964 2973
rect 958 2968 964 2969
rect 1094 2973 1100 2974
rect 1094 2969 1095 2973
rect 1099 2969 1100 2973
rect 1094 2968 1100 2969
rect 1230 2973 1236 2974
rect 1230 2969 1231 2973
rect 1235 2969 1236 2973
rect 1230 2968 1236 2969
rect 1358 2973 1364 2974
rect 1358 2969 1359 2973
rect 1363 2969 1364 2973
rect 1358 2968 1364 2969
rect 1486 2973 1492 2974
rect 1486 2969 1487 2973
rect 1491 2969 1492 2973
rect 1486 2968 1492 2969
rect 1614 2973 1620 2974
rect 1614 2969 1615 2973
rect 1619 2969 1620 2973
rect 1614 2968 1620 2969
rect 1726 2973 1732 2974
rect 1726 2969 1727 2973
rect 1731 2969 1732 2973
rect 1726 2968 1732 2969
rect 1862 2972 1868 2973
rect 1862 2968 1863 2972
rect 1867 2968 1868 2972
rect 1862 2967 1868 2968
rect 3574 2972 3580 2973
rect 3574 2968 3575 2972
rect 3579 2968 3580 2972
rect 3574 2967 3580 2968
rect 2030 2959 2036 2960
rect 2030 2955 2031 2959
rect 2035 2955 2036 2959
rect 2030 2954 2036 2955
rect 2166 2959 2172 2960
rect 2166 2955 2167 2959
rect 2171 2955 2172 2959
rect 2166 2954 2172 2955
rect 2294 2959 2300 2960
rect 2294 2955 2295 2959
rect 2299 2955 2300 2959
rect 2294 2954 2300 2955
rect 2422 2959 2428 2960
rect 2422 2955 2423 2959
rect 2427 2955 2428 2959
rect 2422 2954 2428 2955
rect 2542 2959 2548 2960
rect 2542 2955 2543 2959
rect 2547 2955 2548 2959
rect 2542 2954 2548 2955
rect 2670 2959 2676 2960
rect 2670 2955 2671 2959
rect 2675 2955 2676 2959
rect 2670 2954 2676 2955
rect 2814 2959 2820 2960
rect 2814 2955 2815 2959
rect 2819 2955 2820 2959
rect 2814 2954 2820 2955
rect 2974 2959 2980 2960
rect 2974 2955 2975 2959
rect 2979 2955 2980 2959
rect 2974 2954 2980 2955
rect 3150 2959 3156 2960
rect 3150 2955 3151 2959
rect 3155 2955 3156 2959
rect 3150 2954 3156 2955
rect 3326 2959 3332 2960
rect 3326 2955 3327 2959
rect 3331 2955 3332 2959
rect 3326 2954 3332 2955
rect 3486 2959 3492 2960
rect 3486 2955 3487 2959
rect 3491 2955 3492 2959
rect 3486 2954 3492 2955
rect 494 2951 500 2952
rect 494 2947 495 2951
rect 499 2947 500 2951
rect 494 2946 500 2947
rect 638 2951 644 2952
rect 638 2947 639 2951
rect 643 2947 644 2951
rect 638 2946 644 2947
rect 782 2951 788 2952
rect 782 2947 783 2951
rect 787 2947 788 2951
rect 782 2946 788 2947
rect 918 2951 924 2952
rect 918 2947 919 2951
rect 923 2947 924 2951
rect 918 2946 924 2947
rect 1054 2951 1060 2952
rect 1054 2947 1055 2951
rect 1059 2947 1060 2951
rect 1054 2946 1060 2947
rect 1182 2951 1188 2952
rect 1182 2947 1183 2951
rect 1187 2947 1188 2951
rect 1182 2946 1188 2947
rect 1302 2951 1308 2952
rect 1302 2947 1303 2951
rect 1307 2947 1308 2951
rect 1302 2946 1308 2947
rect 1414 2951 1420 2952
rect 1414 2947 1415 2951
rect 1419 2947 1420 2951
rect 1414 2946 1420 2947
rect 1526 2951 1532 2952
rect 1526 2947 1527 2951
rect 1531 2947 1532 2951
rect 1526 2946 1532 2947
rect 1638 2951 1644 2952
rect 1638 2947 1639 2951
rect 1643 2947 1644 2951
rect 1638 2946 1644 2947
rect 1726 2951 1732 2952
rect 1726 2947 1727 2951
rect 1731 2947 1732 2951
rect 1726 2946 1732 2947
rect 110 2941 116 2942
rect 110 2937 111 2941
rect 115 2937 116 2941
rect 110 2936 116 2937
rect 1822 2941 1828 2942
rect 1822 2937 1823 2941
rect 1827 2937 1828 2941
rect 1822 2936 1828 2937
rect 110 2924 116 2925
rect 110 2920 111 2924
rect 115 2920 116 2924
rect 110 2919 116 2920
rect 1822 2924 1828 2925
rect 1822 2920 1823 2924
rect 1827 2920 1828 2924
rect 1822 2919 1828 2920
rect 1894 2917 1900 2918
rect 1894 2913 1895 2917
rect 1899 2913 1900 2917
rect 1894 2912 1900 2913
rect 2174 2917 2180 2918
rect 2174 2913 2175 2917
rect 2179 2913 2180 2917
rect 2174 2912 2180 2913
rect 2494 2917 2500 2918
rect 2494 2913 2495 2917
rect 2499 2913 2500 2917
rect 2494 2912 2500 2913
rect 2822 2917 2828 2918
rect 2822 2913 2823 2917
rect 2827 2913 2828 2917
rect 2822 2912 2828 2913
rect 3166 2917 3172 2918
rect 3166 2913 3167 2917
rect 3171 2913 3172 2917
rect 3166 2912 3172 2913
rect 3486 2917 3492 2918
rect 3486 2913 3487 2917
rect 3491 2913 3492 2917
rect 3486 2912 3492 2913
rect 502 2911 508 2912
rect 502 2907 503 2911
rect 507 2907 508 2911
rect 502 2906 508 2907
rect 646 2911 652 2912
rect 646 2907 647 2911
rect 651 2907 652 2911
rect 646 2906 652 2907
rect 790 2911 796 2912
rect 790 2907 791 2911
rect 795 2907 796 2911
rect 790 2906 796 2907
rect 926 2911 932 2912
rect 926 2907 927 2911
rect 931 2907 932 2911
rect 926 2906 932 2907
rect 1062 2911 1068 2912
rect 1062 2907 1063 2911
rect 1067 2907 1068 2911
rect 1062 2906 1068 2907
rect 1190 2911 1196 2912
rect 1190 2907 1191 2911
rect 1195 2907 1196 2911
rect 1190 2906 1196 2907
rect 1310 2911 1316 2912
rect 1310 2907 1311 2911
rect 1315 2907 1316 2911
rect 1310 2906 1316 2907
rect 1422 2911 1428 2912
rect 1422 2907 1423 2911
rect 1427 2907 1428 2911
rect 1422 2906 1428 2907
rect 1534 2911 1540 2912
rect 1534 2907 1535 2911
rect 1539 2907 1540 2911
rect 1534 2906 1540 2907
rect 1646 2911 1652 2912
rect 1646 2907 1647 2911
rect 1651 2907 1652 2911
rect 1646 2906 1652 2907
rect 1734 2911 1740 2912
rect 1734 2907 1735 2911
rect 1739 2907 1740 2911
rect 1734 2906 1740 2907
rect 1862 2904 1868 2905
rect 1862 2900 1863 2904
rect 1867 2900 1868 2904
rect 1862 2899 1868 2900
rect 3574 2904 3580 2905
rect 3574 2900 3575 2904
rect 3579 2900 3580 2904
rect 3574 2899 3580 2900
rect 1862 2887 1868 2888
rect 1862 2883 1863 2887
rect 1867 2883 1868 2887
rect 1862 2882 1868 2883
rect 3574 2887 3580 2888
rect 3574 2883 3575 2887
rect 3579 2883 3580 2887
rect 3574 2882 3580 2883
rect 1886 2877 1892 2878
rect 326 2873 332 2874
rect 326 2869 327 2873
rect 331 2869 332 2873
rect 326 2868 332 2869
rect 454 2873 460 2874
rect 454 2869 455 2873
rect 459 2869 460 2873
rect 454 2868 460 2869
rect 590 2873 596 2874
rect 590 2869 591 2873
rect 595 2869 596 2873
rect 590 2868 596 2869
rect 726 2873 732 2874
rect 726 2869 727 2873
rect 731 2869 732 2873
rect 726 2868 732 2869
rect 870 2873 876 2874
rect 870 2869 871 2873
rect 875 2869 876 2873
rect 870 2868 876 2869
rect 1006 2873 1012 2874
rect 1006 2869 1007 2873
rect 1011 2869 1012 2873
rect 1006 2868 1012 2869
rect 1142 2873 1148 2874
rect 1142 2869 1143 2873
rect 1147 2869 1148 2873
rect 1142 2868 1148 2869
rect 1278 2873 1284 2874
rect 1278 2869 1279 2873
rect 1283 2869 1284 2873
rect 1278 2868 1284 2869
rect 1414 2873 1420 2874
rect 1414 2869 1415 2873
rect 1419 2869 1420 2873
rect 1414 2868 1420 2869
rect 1550 2873 1556 2874
rect 1550 2869 1551 2873
rect 1555 2869 1556 2873
rect 1886 2873 1887 2877
rect 1891 2873 1892 2877
rect 1886 2872 1892 2873
rect 2166 2877 2172 2878
rect 2166 2873 2167 2877
rect 2171 2873 2172 2877
rect 2166 2872 2172 2873
rect 2486 2877 2492 2878
rect 2486 2873 2487 2877
rect 2491 2873 2492 2877
rect 2486 2872 2492 2873
rect 2814 2877 2820 2878
rect 2814 2873 2815 2877
rect 2819 2873 2820 2877
rect 2814 2872 2820 2873
rect 3158 2877 3164 2878
rect 3158 2873 3159 2877
rect 3163 2873 3164 2877
rect 3158 2872 3164 2873
rect 3478 2877 3484 2878
rect 3478 2873 3479 2877
rect 3483 2873 3484 2877
rect 3478 2872 3484 2873
rect 1550 2868 1556 2869
rect 110 2860 116 2861
rect 110 2856 111 2860
rect 115 2856 116 2860
rect 110 2855 116 2856
rect 1822 2860 1828 2861
rect 1822 2856 1823 2860
rect 1827 2856 1828 2860
rect 1822 2855 1828 2856
rect 1886 2855 1892 2856
rect 1886 2851 1887 2855
rect 1891 2851 1892 2855
rect 1886 2850 1892 2851
rect 2022 2855 2028 2856
rect 2022 2851 2023 2855
rect 2027 2851 2028 2855
rect 2022 2850 2028 2851
rect 2190 2855 2196 2856
rect 2190 2851 2191 2855
rect 2195 2851 2196 2855
rect 2190 2850 2196 2851
rect 2358 2855 2364 2856
rect 2358 2851 2359 2855
rect 2363 2851 2364 2855
rect 2358 2850 2364 2851
rect 2518 2855 2524 2856
rect 2518 2851 2519 2855
rect 2523 2851 2524 2855
rect 2518 2850 2524 2851
rect 2670 2855 2676 2856
rect 2670 2851 2671 2855
rect 2675 2851 2676 2855
rect 2670 2850 2676 2851
rect 2806 2855 2812 2856
rect 2806 2851 2807 2855
rect 2811 2851 2812 2855
rect 2806 2850 2812 2851
rect 2934 2855 2940 2856
rect 2934 2851 2935 2855
rect 2939 2851 2940 2855
rect 2934 2850 2940 2851
rect 3054 2855 3060 2856
rect 3054 2851 3055 2855
rect 3059 2851 3060 2855
rect 3054 2850 3060 2851
rect 3166 2855 3172 2856
rect 3166 2851 3167 2855
rect 3171 2851 3172 2855
rect 3166 2850 3172 2851
rect 3278 2855 3284 2856
rect 3278 2851 3279 2855
rect 3283 2851 3284 2855
rect 3278 2850 3284 2851
rect 3390 2855 3396 2856
rect 3390 2851 3391 2855
rect 3395 2851 3396 2855
rect 3390 2850 3396 2851
rect 3478 2855 3484 2856
rect 3478 2851 3479 2855
rect 3483 2851 3484 2855
rect 3478 2850 3484 2851
rect 1862 2845 1868 2846
rect 110 2843 116 2844
rect 110 2839 111 2843
rect 115 2839 116 2843
rect 110 2838 116 2839
rect 1822 2843 1828 2844
rect 1822 2839 1823 2843
rect 1827 2839 1828 2843
rect 1862 2841 1863 2845
rect 1867 2841 1868 2845
rect 1862 2840 1868 2841
rect 3574 2845 3580 2846
rect 3574 2841 3575 2845
rect 3579 2841 3580 2845
rect 3574 2840 3580 2841
rect 1822 2838 1828 2839
rect 318 2833 324 2834
rect 318 2829 319 2833
rect 323 2829 324 2833
rect 318 2828 324 2829
rect 446 2833 452 2834
rect 446 2829 447 2833
rect 451 2829 452 2833
rect 446 2828 452 2829
rect 582 2833 588 2834
rect 582 2829 583 2833
rect 587 2829 588 2833
rect 582 2828 588 2829
rect 718 2833 724 2834
rect 718 2829 719 2833
rect 723 2829 724 2833
rect 718 2828 724 2829
rect 862 2833 868 2834
rect 862 2829 863 2833
rect 867 2829 868 2833
rect 862 2828 868 2829
rect 998 2833 1004 2834
rect 998 2829 999 2833
rect 1003 2829 1004 2833
rect 998 2828 1004 2829
rect 1134 2833 1140 2834
rect 1134 2829 1135 2833
rect 1139 2829 1140 2833
rect 1134 2828 1140 2829
rect 1270 2833 1276 2834
rect 1270 2829 1271 2833
rect 1275 2829 1276 2833
rect 1270 2828 1276 2829
rect 1406 2833 1412 2834
rect 1406 2829 1407 2833
rect 1411 2829 1412 2833
rect 1406 2828 1412 2829
rect 1542 2833 1548 2834
rect 1542 2829 1543 2833
rect 1547 2829 1548 2833
rect 1542 2828 1548 2829
rect 1862 2828 1868 2829
rect 1862 2824 1863 2828
rect 1867 2824 1868 2828
rect 1862 2823 1868 2824
rect 3574 2828 3580 2829
rect 3574 2824 3575 2828
rect 3579 2824 3580 2828
rect 3574 2823 3580 2824
rect 1894 2815 1900 2816
rect 1894 2811 1895 2815
rect 1899 2811 1900 2815
rect 1894 2810 1900 2811
rect 2030 2815 2036 2816
rect 2030 2811 2031 2815
rect 2035 2811 2036 2815
rect 2030 2810 2036 2811
rect 2198 2815 2204 2816
rect 2198 2811 2199 2815
rect 2203 2811 2204 2815
rect 2198 2810 2204 2811
rect 2366 2815 2372 2816
rect 2366 2811 2367 2815
rect 2371 2811 2372 2815
rect 2366 2810 2372 2811
rect 2526 2815 2532 2816
rect 2526 2811 2527 2815
rect 2531 2811 2532 2815
rect 2526 2810 2532 2811
rect 2678 2815 2684 2816
rect 2678 2811 2679 2815
rect 2683 2811 2684 2815
rect 2678 2810 2684 2811
rect 2814 2815 2820 2816
rect 2814 2811 2815 2815
rect 2819 2811 2820 2815
rect 2814 2810 2820 2811
rect 2942 2815 2948 2816
rect 2942 2811 2943 2815
rect 2947 2811 2948 2815
rect 2942 2810 2948 2811
rect 3062 2815 3068 2816
rect 3062 2811 3063 2815
rect 3067 2811 3068 2815
rect 3062 2810 3068 2811
rect 3174 2815 3180 2816
rect 3174 2811 3175 2815
rect 3179 2811 3180 2815
rect 3174 2810 3180 2811
rect 3286 2815 3292 2816
rect 3286 2811 3287 2815
rect 3291 2811 3292 2815
rect 3286 2810 3292 2811
rect 3398 2815 3404 2816
rect 3398 2811 3399 2815
rect 3403 2811 3404 2815
rect 3398 2810 3404 2811
rect 3486 2815 3492 2816
rect 3486 2811 3487 2815
rect 3491 2811 3492 2815
rect 3486 2810 3492 2811
rect 166 2803 172 2804
rect 166 2799 167 2803
rect 171 2799 172 2803
rect 166 2798 172 2799
rect 294 2803 300 2804
rect 294 2799 295 2803
rect 299 2799 300 2803
rect 294 2798 300 2799
rect 422 2803 428 2804
rect 422 2799 423 2803
rect 427 2799 428 2803
rect 422 2798 428 2799
rect 558 2803 564 2804
rect 558 2799 559 2803
rect 563 2799 564 2803
rect 558 2798 564 2799
rect 694 2803 700 2804
rect 694 2799 695 2803
rect 699 2799 700 2803
rect 694 2798 700 2799
rect 822 2803 828 2804
rect 822 2799 823 2803
rect 827 2799 828 2803
rect 822 2798 828 2799
rect 950 2803 956 2804
rect 950 2799 951 2803
rect 955 2799 956 2803
rect 950 2798 956 2799
rect 1078 2803 1084 2804
rect 1078 2799 1079 2803
rect 1083 2799 1084 2803
rect 1078 2798 1084 2799
rect 1206 2803 1212 2804
rect 1206 2799 1207 2803
rect 1211 2799 1212 2803
rect 1206 2798 1212 2799
rect 1342 2803 1348 2804
rect 1342 2799 1343 2803
rect 1347 2799 1348 2803
rect 1342 2798 1348 2799
rect 110 2793 116 2794
rect 110 2789 111 2793
rect 115 2789 116 2793
rect 110 2788 116 2789
rect 1822 2793 1828 2794
rect 1822 2789 1823 2793
rect 1827 2789 1828 2793
rect 1822 2788 1828 2789
rect 1894 2781 1900 2782
rect 1894 2777 1895 2781
rect 1899 2777 1900 2781
rect 110 2776 116 2777
rect 110 2772 111 2776
rect 115 2772 116 2776
rect 110 2771 116 2772
rect 1822 2776 1828 2777
rect 1894 2776 1900 2777
rect 2062 2781 2068 2782
rect 2062 2777 2063 2781
rect 2067 2777 2068 2781
rect 2062 2776 2068 2777
rect 2254 2781 2260 2782
rect 2254 2777 2255 2781
rect 2259 2777 2260 2781
rect 2254 2776 2260 2777
rect 2438 2781 2444 2782
rect 2438 2777 2439 2781
rect 2443 2777 2444 2781
rect 2438 2776 2444 2777
rect 2614 2781 2620 2782
rect 2614 2777 2615 2781
rect 2619 2777 2620 2781
rect 2614 2776 2620 2777
rect 2782 2781 2788 2782
rect 2782 2777 2783 2781
rect 2787 2777 2788 2781
rect 2782 2776 2788 2777
rect 2934 2781 2940 2782
rect 2934 2777 2935 2781
rect 2939 2777 2940 2781
rect 2934 2776 2940 2777
rect 3078 2781 3084 2782
rect 3078 2777 3079 2781
rect 3083 2777 3084 2781
rect 3078 2776 3084 2777
rect 3222 2781 3228 2782
rect 3222 2777 3223 2781
rect 3227 2777 3228 2781
rect 3222 2776 3228 2777
rect 3366 2781 3372 2782
rect 3366 2777 3367 2781
rect 3371 2777 3372 2781
rect 3366 2776 3372 2777
rect 3486 2781 3492 2782
rect 3486 2777 3487 2781
rect 3491 2777 3492 2781
rect 3486 2776 3492 2777
rect 1822 2772 1823 2776
rect 1827 2772 1828 2776
rect 1822 2771 1828 2772
rect 1862 2768 1868 2769
rect 1862 2764 1863 2768
rect 1867 2764 1868 2768
rect 174 2763 180 2764
rect 174 2759 175 2763
rect 179 2759 180 2763
rect 174 2758 180 2759
rect 302 2763 308 2764
rect 302 2759 303 2763
rect 307 2759 308 2763
rect 302 2758 308 2759
rect 430 2763 436 2764
rect 430 2759 431 2763
rect 435 2759 436 2763
rect 430 2758 436 2759
rect 566 2763 572 2764
rect 566 2759 567 2763
rect 571 2759 572 2763
rect 566 2758 572 2759
rect 702 2763 708 2764
rect 702 2759 703 2763
rect 707 2759 708 2763
rect 702 2758 708 2759
rect 830 2763 836 2764
rect 830 2759 831 2763
rect 835 2759 836 2763
rect 830 2758 836 2759
rect 958 2763 964 2764
rect 958 2759 959 2763
rect 963 2759 964 2763
rect 958 2758 964 2759
rect 1086 2763 1092 2764
rect 1086 2759 1087 2763
rect 1091 2759 1092 2763
rect 1086 2758 1092 2759
rect 1214 2763 1220 2764
rect 1214 2759 1215 2763
rect 1219 2759 1220 2763
rect 1214 2758 1220 2759
rect 1350 2763 1356 2764
rect 1862 2763 1868 2764
rect 3574 2768 3580 2769
rect 3574 2764 3575 2768
rect 3579 2764 3580 2768
rect 3574 2763 3580 2764
rect 1350 2759 1351 2763
rect 1355 2759 1356 2763
rect 1350 2758 1356 2759
rect 1862 2751 1868 2752
rect 1862 2747 1863 2751
rect 1867 2747 1868 2751
rect 1862 2746 1868 2747
rect 3574 2751 3580 2752
rect 3574 2747 3575 2751
rect 3579 2747 3580 2751
rect 3574 2746 3580 2747
rect 1886 2741 1892 2742
rect 1886 2737 1887 2741
rect 1891 2737 1892 2741
rect 1886 2736 1892 2737
rect 2054 2741 2060 2742
rect 2054 2737 2055 2741
rect 2059 2737 2060 2741
rect 2054 2736 2060 2737
rect 2246 2741 2252 2742
rect 2246 2737 2247 2741
rect 2251 2737 2252 2741
rect 2246 2736 2252 2737
rect 2430 2741 2436 2742
rect 2430 2737 2431 2741
rect 2435 2737 2436 2741
rect 2430 2736 2436 2737
rect 2606 2741 2612 2742
rect 2606 2737 2607 2741
rect 2611 2737 2612 2741
rect 2606 2736 2612 2737
rect 2774 2741 2780 2742
rect 2774 2737 2775 2741
rect 2779 2737 2780 2741
rect 2774 2736 2780 2737
rect 2926 2741 2932 2742
rect 2926 2737 2927 2741
rect 2931 2737 2932 2741
rect 2926 2736 2932 2737
rect 3070 2741 3076 2742
rect 3070 2737 3071 2741
rect 3075 2737 3076 2741
rect 3070 2736 3076 2737
rect 3214 2741 3220 2742
rect 3214 2737 3215 2741
rect 3219 2737 3220 2741
rect 3214 2736 3220 2737
rect 3358 2741 3364 2742
rect 3358 2737 3359 2741
rect 3363 2737 3364 2741
rect 3358 2736 3364 2737
rect 3478 2741 3484 2742
rect 3478 2737 3479 2741
rect 3483 2737 3484 2741
rect 3478 2736 3484 2737
rect 142 2721 148 2722
rect 142 2717 143 2721
rect 147 2717 148 2721
rect 142 2716 148 2717
rect 230 2721 236 2722
rect 230 2717 231 2721
rect 235 2717 236 2721
rect 230 2716 236 2717
rect 350 2721 356 2722
rect 350 2717 351 2721
rect 355 2717 356 2721
rect 350 2716 356 2717
rect 478 2721 484 2722
rect 478 2717 479 2721
rect 483 2717 484 2721
rect 478 2716 484 2717
rect 614 2721 620 2722
rect 614 2717 615 2721
rect 619 2717 620 2721
rect 614 2716 620 2717
rect 758 2721 764 2722
rect 758 2717 759 2721
rect 763 2717 764 2721
rect 758 2716 764 2717
rect 902 2721 908 2722
rect 902 2717 903 2721
rect 907 2717 908 2721
rect 902 2716 908 2717
rect 1046 2721 1052 2722
rect 1046 2717 1047 2721
rect 1051 2717 1052 2721
rect 1046 2716 1052 2717
rect 1886 2715 1892 2716
rect 1886 2711 1887 2715
rect 1891 2711 1892 2715
rect 1886 2710 1892 2711
rect 2046 2715 2052 2716
rect 2046 2711 2047 2715
rect 2051 2711 2052 2715
rect 2046 2710 2052 2711
rect 2206 2715 2212 2716
rect 2206 2711 2207 2715
rect 2211 2711 2212 2715
rect 2206 2710 2212 2711
rect 2358 2715 2364 2716
rect 2358 2711 2359 2715
rect 2363 2711 2364 2715
rect 2358 2710 2364 2711
rect 2494 2715 2500 2716
rect 2494 2711 2495 2715
rect 2499 2711 2500 2715
rect 2494 2710 2500 2711
rect 2622 2715 2628 2716
rect 2622 2711 2623 2715
rect 2627 2711 2628 2715
rect 2622 2710 2628 2711
rect 2742 2715 2748 2716
rect 2742 2711 2743 2715
rect 2747 2711 2748 2715
rect 2742 2710 2748 2711
rect 2862 2715 2868 2716
rect 2862 2711 2863 2715
rect 2867 2711 2868 2715
rect 2862 2710 2868 2711
rect 2982 2715 2988 2716
rect 2982 2711 2983 2715
rect 2987 2711 2988 2715
rect 2982 2710 2988 2711
rect 3102 2715 3108 2716
rect 3102 2711 3103 2715
rect 3107 2711 3108 2715
rect 3102 2710 3108 2711
rect 110 2708 116 2709
rect 110 2704 111 2708
rect 115 2704 116 2708
rect 110 2703 116 2704
rect 1822 2708 1828 2709
rect 1822 2704 1823 2708
rect 1827 2704 1828 2708
rect 1822 2703 1828 2704
rect 1862 2705 1868 2706
rect 1862 2701 1863 2705
rect 1867 2701 1868 2705
rect 1862 2700 1868 2701
rect 3574 2705 3580 2706
rect 3574 2701 3575 2705
rect 3579 2701 3580 2705
rect 3574 2700 3580 2701
rect 110 2691 116 2692
rect 110 2687 111 2691
rect 115 2687 116 2691
rect 110 2686 116 2687
rect 1822 2691 1828 2692
rect 1822 2687 1823 2691
rect 1827 2687 1828 2691
rect 1822 2686 1828 2687
rect 1862 2688 1868 2689
rect 1862 2684 1863 2688
rect 1867 2684 1868 2688
rect 1862 2683 1868 2684
rect 3574 2688 3580 2689
rect 3574 2684 3575 2688
rect 3579 2684 3580 2688
rect 3574 2683 3580 2684
rect 134 2681 140 2682
rect 134 2677 135 2681
rect 139 2677 140 2681
rect 134 2676 140 2677
rect 222 2681 228 2682
rect 222 2677 223 2681
rect 227 2677 228 2681
rect 222 2676 228 2677
rect 342 2681 348 2682
rect 342 2677 343 2681
rect 347 2677 348 2681
rect 342 2676 348 2677
rect 470 2681 476 2682
rect 470 2677 471 2681
rect 475 2677 476 2681
rect 470 2676 476 2677
rect 606 2681 612 2682
rect 606 2677 607 2681
rect 611 2677 612 2681
rect 606 2676 612 2677
rect 750 2681 756 2682
rect 750 2677 751 2681
rect 755 2677 756 2681
rect 750 2676 756 2677
rect 894 2681 900 2682
rect 894 2677 895 2681
rect 899 2677 900 2681
rect 894 2676 900 2677
rect 1038 2681 1044 2682
rect 1038 2677 1039 2681
rect 1043 2677 1044 2681
rect 1038 2676 1044 2677
rect 1894 2675 1900 2676
rect 1894 2671 1895 2675
rect 1899 2671 1900 2675
rect 1894 2670 1900 2671
rect 2054 2675 2060 2676
rect 2054 2671 2055 2675
rect 2059 2671 2060 2675
rect 2054 2670 2060 2671
rect 2214 2675 2220 2676
rect 2214 2671 2215 2675
rect 2219 2671 2220 2675
rect 2214 2670 2220 2671
rect 2366 2675 2372 2676
rect 2366 2671 2367 2675
rect 2371 2671 2372 2675
rect 2366 2670 2372 2671
rect 2502 2675 2508 2676
rect 2502 2671 2503 2675
rect 2507 2671 2508 2675
rect 2502 2670 2508 2671
rect 2630 2675 2636 2676
rect 2630 2671 2631 2675
rect 2635 2671 2636 2675
rect 2630 2670 2636 2671
rect 2750 2675 2756 2676
rect 2750 2671 2751 2675
rect 2755 2671 2756 2675
rect 2750 2670 2756 2671
rect 2870 2675 2876 2676
rect 2870 2671 2871 2675
rect 2875 2671 2876 2675
rect 2870 2670 2876 2671
rect 2990 2675 2996 2676
rect 2990 2671 2991 2675
rect 2995 2671 2996 2675
rect 2990 2670 2996 2671
rect 3110 2675 3116 2676
rect 3110 2671 3111 2675
rect 3115 2671 3116 2675
rect 3110 2670 3116 2671
rect 134 2655 140 2656
rect 134 2651 135 2655
rect 139 2651 140 2655
rect 134 2650 140 2651
rect 230 2655 236 2656
rect 230 2651 231 2655
rect 235 2651 236 2655
rect 230 2650 236 2651
rect 350 2655 356 2656
rect 350 2651 351 2655
rect 355 2651 356 2655
rect 350 2650 356 2651
rect 470 2655 476 2656
rect 470 2651 471 2655
rect 475 2651 476 2655
rect 470 2650 476 2651
rect 582 2655 588 2656
rect 582 2651 583 2655
rect 587 2651 588 2655
rect 582 2650 588 2651
rect 694 2655 700 2656
rect 694 2651 695 2655
rect 699 2651 700 2655
rect 694 2650 700 2651
rect 798 2655 804 2656
rect 798 2651 799 2655
rect 803 2651 804 2655
rect 798 2650 804 2651
rect 902 2655 908 2656
rect 902 2651 903 2655
rect 907 2651 908 2655
rect 902 2650 908 2651
rect 998 2655 1004 2656
rect 998 2651 999 2655
rect 1003 2651 1004 2655
rect 998 2650 1004 2651
rect 1102 2655 1108 2656
rect 1102 2651 1103 2655
rect 1107 2651 1108 2655
rect 1102 2650 1108 2651
rect 1206 2655 1212 2656
rect 1206 2651 1207 2655
rect 1211 2651 1212 2655
rect 1206 2650 1212 2651
rect 1310 2655 1316 2656
rect 1310 2651 1311 2655
rect 1315 2651 1316 2655
rect 1310 2650 1316 2651
rect 110 2645 116 2646
rect 110 2641 111 2645
rect 115 2641 116 2645
rect 110 2640 116 2641
rect 1822 2645 1828 2646
rect 1822 2641 1823 2645
rect 1827 2641 1828 2645
rect 1822 2640 1828 2641
rect 1894 2633 1900 2634
rect 1894 2629 1895 2633
rect 1899 2629 1900 2633
rect 110 2628 116 2629
rect 110 2624 111 2628
rect 115 2624 116 2628
rect 110 2623 116 2624
rect 1822 2628 1828 2629
rect 1894 2628 1900 2629
rect 1998 2633 2004 2634
rect 1998 2629 1999 2633
rect 2003 2629 2004 2633
rect 1998 2628 2004 2629
rect 2118 2633 2124 2634
rect 2118 2629 2119 2633
rect 2123 2629 2124 2633
rect 2118 2628 2124 2629
rect 2238 2633 2244 2634
rect 2238 2629 2239 2633
rect 2243 2629 2244 2633
rect 2238 2628 2244 2629
rect 2350 2633 2356 2634
rect 2350 2629 2351 2633
rect 2355 2629 2356 2633
rect 2350 2628 2356 2629
rect 2454 2633 2460 2634
rect 2454 2629 2455 2633
rect 2459 2629 2460 2633
rect 2454 2628 2460 2629
rect 2550 2633 2556 2634
rect 2550 2629 2551 2633
rect 2555 2629 2556 2633
rect 2550 2628 2556 2629
rect 2654 2633 2660 2634
rect 2654 2629 2655 2633
rect 2659 2629 2660 2633
rect 2654 2628 2660 2629
rect 2758 2633 2764 2634
rect 2758 2629 2759 2633
rect 2763 2629 2764 2633
rect 2758 2628 2764 2629
rect 2862 2633 2868 2634
rect 2862 2629 2863 2633
rect 2867 2629 2868 2633
rect 2862 2628 2868 2629
rect 1822 2624 1823 2628
rect 1827 2624 1828 2628
rect 1822 2623 1828 2624
rect 1862 2620 1868 2621
rect 1862 2616 1863 2620
rect 1867 2616 1868 2620
rect 142 2615 148 2616
rect 142 2611 143 2615
rect 147 2611 148 2615
rect 142 2610 148 2611
rect 238 2615 244 2616
rect 238 2611 239 2615
rect 243 2611 244 2615
rect 238 2610 244 2611
rect 358 2615 364 2616
rect 358 2611 359 2615
rect 363 2611 364 2615
rect 358 2610 364 2611
rect 478 2615 484 2616
rect 478 2611 479 2615
rect 483 2611 484 2615
rect 478 2610 484 2611
rect 590 2615 596 2616
rect 590 2611 591 2615
rect 595 2611 596 2615
rect 590 2610 596 2611
rect 702 2615 708 2616
rect 702 2611 703 2615
rect 707 2611 708 2615
rect 702 2610 708 2611
rect 806 2615 812 2616
rect 806 2611 807 2615
rect 811 2611 812 2615
rect 806 2610 812 2611
rect 910 2615 916 2616
rect 910 2611 911 2615
rect 915 2611 916 2615
rect 910 2610 916 2611
rect 1006 2615 1012 2616
rect 1006 2611 1007 2615
rect 1011 2611 1012 2615
rect 1006 2610 1012 2611
rect 1110 2615 1116 2616
rect 1110 2611 1111 2615
rect 1115 2611 1116 2615
rect 1110 2610 1116 2611
rect 1214 2615 1220 2616
rect 1214 2611 1215 2615
rect 1219 2611 1220 2615
rect 1214 2610 1220 2611
rect 1318 2615 1324 2616
rect 1862 2615 1868 2616
rect 3574 2620 3580 2621
rect 3574 2616 3575 2620
rect 3579 2616 3580 2620
rect 3574 2615 3580 2616
rect 1318 2611 1319 2615
rect 1323 2611 1324 2615
rect 1318 2610 1324 2611
rect 1862 2603 1868 2604
rect 1862 2599 1863 2603
rect 1867 2599 1868 2603
rect 1862 2598 1868 2599
rect 3574 2603 3580 2604
rect 3574 2599 3575 2603
rect 3579 2599 3580 2603
rect 3574 2598 3580 2599
rect 1886 2593 1892 2594
rect 1886 2589 1887 2593
rect 1891 2589 1892 2593
rect 1886 2588 1892 2589
rect 1990 2593 1996 2594
rect 1990 2589 1991 2593
rect 1995 2589 1996 2593
rect 1990 2588 1996 2589
rect 2110 2593 2116 2594
rect 2110 2589 2111 2593
rect 2115 2589 2116 2593
rect 2110 2588 2116 2589
rect 2230 2593 2236 2594
rect 2230 2589 2231 2593
rect 2235 2589 2236 2593
rect 2230 2588 2236 2589
rect 2342 2593 2348 2594
rect 2342 2589 2343 2593
rect 2347 2589 2348 2593
rect 2342 2588 2348 2589
rect 2446 2593 2452 2594
rect 2446 2589 2447 2593
rect 2451 2589 2452 2593
rect 2446 2588 2452 2589
rect 2542 2593 2548 2594
rect 2542 2589 2543 2593
rect 2547 2589 2548 2593
rect 2542 2588 2548 2589
rect 2646 2593 2652 2594
rect 2646 2589 2647 2593
rect 2651 2589 2652 2593
rect 2646 2588 2652 2589
rect 2750 2593 2756 2594
rect 2750 2589 2751 2593
rect 2755 2589 2756 2593
rect 2750 2588 2756 2589
rect 2854 2593 2860 2594
rect 2854 2589 2855 2593
rect 2859 2589 2860 2593
rect 2854 2588 2860 2589
rect 142 2577 148 2578
rect 142 2573 143 2577
rect 147 2573 148 2577
rect 142 2572 148 2573
rect 270 2577 276 2578
rect 270 2573 271 2577
rect 275 2573 276 2577
rect 270 2572 276 2573
rect 414 2577 420 2578
rect 414 2573 415 2577
rect 419 2573 420 2577
rect 414 2572 420 2573
rect 550 2577 556 2578
rect 550 2573 551 2577
rect 555 2573 556 2577
rect 550 2572 556 2573
rect 678 2577 684 2578
rect 678 2573 679 2577
rect 683 2573 684 2577
rect 678 2572 684 2573
rect 806 2577 812 2578
rect 806 2573 807 2577
rect 811 2573 812 2577
rect 806 2572 812 2573
rect 926 2577 932 2578
rect 926 2573 927 2577
rect 931 2573 932 2577
rect 926 2572 932 2573
rect 1046 2577 1052 2578
rect 1046 2573 1047 2577
rect 1051 2573 1052 2577
rect 1046 2572 1052 2573
rect 1174 2577 1180 2578
rect 1174 2573 1175 2577
rect 1179 2573 1180 2577
rect 1174 2572 1180 2573
rect 1886 2567 1892 2568
rect 110 2564 116 2565
rect 110 2560 111 2564
rect 115 2560 116 2564
rect 110 2559 116 2560
rect 1822 2564 1828 2565
rect 1822 2560 1823 2564
rect 1827 2560 1828 2564
rect 1886 2563 1887 2567
rect 1891 2563 1892 2567
rect 1886 2562 1892 2563
rect 1990 2567 1996 2568
rect 1990 2563 1991 2567
rect 1995 2563 1996 2567
rect 1990 2562 1996 2563
rect 2110 2567 2116 2568
rect 2110 2563 2111 2567
rect 2115 2563 2116 2567
rect 2110 2562 2116 2563
rect 2230 2567 2236 2568
rect 2230 2563 2231 2567
rect 2235 2563 2236 2567
rect 2230 2562 2236 2563
rect 2350 2567 2356 2568
rect 2350 2563 2351 2567
rect 2355 2563 2356 2567
rect 2350 2562 2356 2563
rect 2470 2567 2476 2568
rect 2470 2563 2471 2567
rect 2475 2563 2476 2567
rect 2470 2562 2476 2563
rect 2590 2567 2596 2568
rect 2590 2563 2591 2567
rect 2595 2563 2596 2567
rect 2590 2562 2596 2563
rect 2710 2567 2716 2568
rect 2710 2563 2711 2567
rect 2715 2563 2716 2567
rect 2710 2562 2716 2563
rect 2830 2567 2836 2568
rect 2830 2563 2831 2567
rect 2835 2563 2836 2567
rect 2830 2562 2836 2563
rect 1822 2559 1828 2560
rect 1862 2557 1868 2558
rect 1862 2553 1863 2557
rect 1867 2553 1868 2557
rect 1862 2552 1868 2553
rect 3574 2557 3580 2558
rect 3574 2553 3575 2557
rect 3579 2553 3580 2557
rect 3574 2552 3580 2553
rect 110 2547 116 2548
rect 110 2543 111 2547
rect 115 2543 116 2547
rect 110 2542 116 2543
rect 1822 2547 1828 2548
rect 1822 2543 1823 2547
rect 1827 2543 1828 2547
rect 1822 2542 1828 2543
rect 1862 2540 1868 2541
rect 134 2537 140 2538
rect 134 2533 135 2537
rect 139 2533 140 2537
rect 134 2532 140 2533
rect 262 2537 268 2538
rect 262 2533 263 2537
rect 267 2533 268 2537
rect 262 2532 268 2533
rect 406 2537 412 2538
rect 406 2533 407 2537
rect 411 2533 412 2537
rect 406 2532 412 2533
rect 542 2537 548 2538
rect 542 2533 543 2537
rect 547 2533 548 2537
rect 542 2532 548 2533
rect 670 2537 676 2538
rect 670 2533 671 2537
rect 675 2533 676 2537
rect 670 2532 676 2533
rect 798 2537 804 2538
rect 798 2533 799 2537
rect 803 2533 804 2537
rect 798 2532 804 2533
rect 918 2537 924 2538
rect 918 2533 919 2537
rect 923 2533 924 2537
rect 918 2532 924 2533
rect 1038 2537 1044 2538
rect 1038 2533 1039 2537
rect 1043 2533 1044 2537
rect 1038 2532 1044 2533
rect 1166 2537 1172 2538
rect 1166 2533 1167 2537
rect 1171 2533 1172 2537
rect 1862 2536 1863 2540
rect 1867 2536 1868 2540
rect 1862 2535 1868 2536
rect 3574 2540 3580 2541
rect 3574 2536 3575 2540
rect 3579 2536 3580 2540
rect 3574 2535 3580 2536
rect 1166 2532 1172 2533
rect 1894 2527 1900 2528
rect 1894 2523 1895 2527
rect 1899 2523 1900 2527
rect 1894 2522 1900 2523
rect 1998 2527 2004 2528
rect 1998 2523 1999 2527
rect 2003 2523 2004 2527
rect 1998 2522 2004 2523
rect 2118 2527 2124 2528
rect 2118 2523 2119 2527
rect 2123 2523 2124 2527
rect 2118 2522 2124 2523
rect 2238 2527 2244 2528
rect 2238 2523 2239 2527
rect 2243 2523 2244 2527
rect 2238 2522 2244 2523
rect 2358 2527 2364 2528
rect 2358 2523 2359 2527
rect 2363 2523 2364 2527
rect 2358 2522 2364 2523
rect 2478 2527 2484 2528
rect 2478 2523 2479 2527
rect 2483 2523 2484 2527
rect 2478 2522 2484 2523
rect 2598 2527 2604 2528
rect 2598 2523 2599 2527
rect 2603 2523 2604 2527
rect 2598 2522 2604 2523
rect 2718 2527 2724 2528
rect 2718 2523 2719 2527
rect 2723 2523 2724 2527
rect 2718 2522 2724 2523
rect 2838 2527 2844 2528
rect 2838 2523 2839 2527
rect 2843 2523 2844 2527
rect 2838 2522 2844 2523
rect 134 2515 140 2516
rect 134 2511 135 2515
rect 139 2511 140 2515
rect 134 2510 140 2511
rect 278 2515 284 2516
rect 278 2511 279 2515
rect 283 2511 284 2515
rect 278 2510 284 2511
rect 438 2515 444 2516
rect 438 2511 439 2515
rect 443 2511 444 2515
rect 438 2510 444 2511
rect 590 2515 596 2516
rect 590 2511 591 2515
rect 595 2511 596 2515
rect 590 2510 596 2511
rect 734 2515 740 2516
rect 734 2511 735 2515
rect 739 2511 740 2515
rect 734 2510 740 2511
rect 870 2515 876 2516
rect 870 2511 871 2515
rect 875 2511 876 2515
rect 870 2510 876 2511
rect 1006 2515 1012 2516
rect 1006 2511 1007 2515
rect 1011 2511 1012 2515
rect 1006 2510 1012 2511
rect 1142 2515 1148 2516
rect 1142 2511 1143 2515
rect 1147 2511 1148 2515
rect 1142 2510 1148 2511
rect 1278 2515 1284 2516
rect 1278 2511 1279 2515
rect 1283 2511 1284 2515
rect 1278 2510 1284 2511
rect 110 2505 116 2506
rect 110 2501 111 2505
rect 115 2501 116 2505
rect 110 2500 116 2501
rect 1822 2505 1828 2506
rect 1822 2501 1823 2505
rect 1827 2501 1828 2505
rect 1822 2500 1828 2501
rect 1894 2489 1900 2490
rect 110 2488 116 2489
rect 110 2484 111 2488
rect 115 2484 116 2488
rect 110 2483 116 2484
rect 1822 2488 1828 2489
rect 1822 2484 1823 2488
rect 1827 2484 1828 2488
rect 1894 2485 1895 2489
rect 1899 2485 1900 2489
rect 1894 2484 1900 2485
rect 2030 2489 2036 2490
rect 2030 2485 2031 2489
rect 2035 2485 2036 2489
rect 2030 2484 2036 2485
rect 2190 2489 2196 2490
rect 2190 2485 2191 2489
rect 2195 2485 2196 2489
rect 2190 2484 2196 2485
rect 2342 2489 2348 2490
rect 2342 2485 2343 2489
rect 2347 2485 2348 2489
rect 2342 2484 2348 2485
rect 2486 2489 2492 2490
rect 2486 2485 2487 2489
rect 2491 2485 2492 2489
rect 2486 2484 2492 2485
rect 2622 2489 2628 2490
rect 2622 2485 2623 2489
rect 2627 2485 2628 2489
rect 2622 2484 2628 2485
rect 2750 2489 2756 2490
rect 2750 2485 2751 2489
rect 2755 2485 2756 2489
rect 2750 2484 2756 2485
rect 2878 2489 2884 2490
rect 2878 2485 2879 2489
rect 2883 2485 2884 2489
rect 2878 2484 2884 2485
rect 3014 2489 3020 2490
rect 3014 2485 3015 2489
rect 3019 2485 3020 2489
rect 3014 2484 3020 2485
rect 1822 2483 1828 2484
rect 1862 2476 1868 2477
rect 142 2475 148 2476
rect 142 2471 143 2475
rect 147 2471 148 2475
rect 142 2470 148 2471
rect 286 2475 292 2476
rect 286 2471 287 2475
rect 291 2471 292 2475
rect 286 2470 292 2471
rect 446 2475 452 2476
rect 446 2471 447 2475
rect 451 2471 452 2475
rect 446 2470 452 2471
rect 598 2475 604 2476
rect 598 2471 599 2475
rect 603 2471 604 2475
rect 598 2470 604 2471
rect 742 2475 748 2476
rect 742 2471 743 2475
rect 747 2471 748 2475
rect 742 2470 748 2471
rect 878 2475 884 2476
rect 878 2471 879 2475
rect 883 2471 884 2475
rect 878 2470 884 2471
rect 1014 2475 1020 2476
rect 1014 2471 1015 2475
rect 1019 2471 1020 2475
rect 1014 2470 1020 2471
rect 1150 2475 1156 2476
rect 1150 2471 1151 2475
rect 1155 2471 1156 2475
rect 1150 2470 1156 2471
rect 1286 2475 1292 2476
rect 1286 2471 1287 2475
rect 1291 2471 1292 2475
rect 1862 2472 1863 2476
rect 1867 2472 1868 2476
rect 1862 2471 1868 2472
rect 3574 2476 3580 2477
rect 3574 2472 3575 2476
rect 3579 2472 3580 2476
rect 3574 2471 3580 2472
rect 1286 2470 1292 2471
rect 1862 2459 1868 2460
rect 1862 2455 1863 2459
rect 1867 2455 1868 2459
rect 1862 2454 1868 2455
rect 3574 2459 3580 2460
rect 3574 2455 3575 2459
rect 3579 2455 3580 2459
rect 3574 2454 3580 2455
rect 1886 2449 1892 2450
rect 1886 2445 1887 2449
rect 1891 2445 1892 2449
rect 1886 2444 1892 2445
rect 2022 2449 2028 2450
rect 2022 2445 2023 2449
rect 2027 2445 2028 2449
rect 2022 2444 2028 2445
rect 2182 2449 2188 2450
rect 2182 2445 2183 2449
rect 2187 2445 2188 2449
rect 2182 2444 2188 2445
rect 2334 2449 2340 2450
rect 2334 2445 2335 2449
rect 2339 2445 2340 2449
rect 2334 2444 2340 2445
rect 2478 2449 2484 2450
rect 2478 2445 2479 2449
rect 2483 2445 2484 2449
rect 2478 2444 2484 2445
rect 2614 2449 2620 2450
rect 2614 2445 2615 2449
rect 2619 2445 2620 2449
rect 2614 2444 2620 2445
rect 2742 2449 2748 2450
rect 2742 2445 2743 2449
rect 2747 2445 2748 2449
rect 2742 2444 2748 2445
rect 2870 2449 2876 2450
rect 2870 2445 2871 2449
rect 2875 2445 2876 2449
rect 2870 2444 2876 2445
rect 3006 2449 3012 2450
rect 3006 2445 3007 2449
rect 3011 2445 3012 2449
rect 3006 2444 3012 2445
rect 190 2441 196 2442
rect 190 2437 191 2441
rect 195 2437 196 2441
rect 190 2436 196 2437
rect 318 2441 324 2442
rect 318 2437 319 2441
rect 323 2437 324 2441
rect 318 2436 324 2437
rect 454 2441 460 2442
rect 454 2437 455 2441
rect 459 2437 460 2441
rect 454 2436 460 2437
rect 590 2441 596 2442
rect 590 2437 591 2441
rect 595 2437 596 2441
rect 590 2436 596 2437
rect 726 2441 732 2442
rect 726 2437 727 2441
rect 731 2437 732 2441
rect 726 2436 732 2437
rect 862 2441 868 2442
rect 862 2437 863 2441
rect 867 2437 868 2441
rect 862 2436 868 2437
rect 998 2441 1004 2442
rect 998 2437 999 2441
rect 1003 2437 1004 2441
rect 998 2436 1004 2437
rect 1134 2441 1140 2442
rect 1134 2437 1135 2441
rect 1139 2437 1140 2441
rect 1134 2436 1140 2437
rect 1270 2441 1276 2442
rect 1270 2437 1271 2441
rect 1275 2437 1276 2441
rect 1270 2436 1276 2437
rect 1406 2441 1412 2442
rect 1406 2437 1407 2441
rect 1411 2437 1412 2441
rect 1406 2436 1412 2437
rect 110 2428 116 2429
rect 110 2424 111 2428
rect 115 2424 116 2428
rect 110 2423 116 2424
rect 1822 2428 1828 2429
rect 1822 2424 1823 2428
rect 1827 2424 1828 2428
rect 1822 2423 1828 2424
rect 1886 2427 1892 2428
rect 1886 2423 1887 2427
rect 1891 2423 1892 2427
rect 1886 2422 1892 2423
rect 2014 2427 2020 2428
rect 2014 2423 2015 2427
rect 2019 2423 2020 2427
rect 2014 2422 2020 2423
rect 2174 2427 2180 2428
rect 2174 2423 2175 2427
rect 2179 2423 2180 2427
rect 2174 2422 2180 2423
rect 2334 2427 2340 2428
rect 2334 2423 2335 2427
rect 2339 2423 2340 2427
rect 2334 2422 2340 2423
rect 2494 2427 2500 2428
rect 2494 2423 2495 2427
rect 2499 2423 2500 2427
rect 2494 2422 2500 2423
rect 2646 2427 2652 2428
rect 2646 2423 2647 2427
rect 2651 2423 2652 2427
rect 2646 2422 2652 2423
rect 2798 2427 2804 2428
rect 2798 2423 2799 2427
rect 2803 2423 2804 2427
rect 2798 2422 2804 2423
rect 2950 2427 2956 2428
rect 2950 2423 2951 2427
rect 2955 2423 2956 2427
rect 2950 2422 2956 2423
rect 3110 2427 3116 2428
rect 3110 2423 3111 2427
rect 3115 2423 3116 2427
rect 3110 2422 3116 2423
rect 1862 2417 1868 2418
rect 1862 2413 1863 2417
rect 1867 2413 1868 2417
rect 1862 2412 1868 2413
rect 3574 2417 3580 2418
rect 3574 2413 3575 2417
rect 3579 2413 3580 2417
rect 3574 2412 3580 2413
rect 110 2411 116 2412
rect 110 2407 111 2411
rect 115 2407 116 2411
rect 110 2406 116 2407
rect 1822 2411 1828 2412
rect 1822 2407 1823 2411
rect 1827 2407 1828 2411
rect 1822 2406 1828 2407
rect 182 2401 188 2402
rect 182 2397 183 2401
rect 187 2397 188 2401
rect 182 2396 188 2397
rect 310 2401 316 2402
rect 310 2397 311 2401
rect 315 2397 316 2401
rect 310 2396 316 2397
rect 446 2401 452 2402
rect 446 2397 447 2401
rect 451 2397 452 2401
rect 446 2396 452 2397
rect 582 2401 588 2402
rect 582 2397 583 2401
rect 587 2397 588 2401
rect 582 2396 588 2397
rect 718 2401 724 2402
rect 718 2397 719 2401
rect 723 2397 724 2401
rect 718 2396 724 2397
rect 854 2401 860 2402
rect 854 2397 855 2401
rect 859 2397 860 2401
rect 854 2396 860 2397
rect 990 2401 996 2402
rect 990 2397 991 2401
rect 995 2397 996 2401
rect 990 2396 996 2397
rect 1126 2401 1132 2402
rect 1126 2397 1127 2401
rect 1131 2397 1132 2401
rect 1126 2396 1132 2397
rect 1262 2401 1268 2402
rect 1262 2397 1263 2401
rect 1267 2397 1268 2401
rect 1262 2396 1268 2397
rect 1398 2401 1404 2402
rect 1398 2397 1399 2401
rect 1403 2397 1404 2401
rect 1398 2396 1404 2397
rect 1862 2400 1868 2401
rect 1862 2396 1863 2400
rect 1867 2396 1868 2400
rect 1862 2395 1868 2396
rect 3574 2400 3580 2401
rect 3574 2396 3575 2400
rect 3579 2396 3580 2400
rect 3574 2395 3580 2396
rect 1894 2387 1900 2388
rect 1894 2383 1895 2387
rect 1899 2383 1900 2387
rect 1894 2382 1900 2383
rect 2022 2387 2028 2388
rect 2022 2383 2023 2387
rect 2027 2383 2028 2387
rect 2022 2382 2028 2383
rect 2182 2387 2188 2388
rect 2182 2383 2183 2387
rect 2187 2383 2188 2387
rect 2182 2382 2188 2383
rect 2342 2387 2348 2388
rect 2342 2383 2343 2387
rect 2347 2383 2348 2387
rect 2342 2382 2348 2383
rect 2502 2387 2508 2388
rect 2502 2383 2503 2387
rect 2507 2383 2508 2387
rect 2502 2382 2508 2383
rect 2654 2387 2660 2388
rect 2654 2383 2655 2387
rect 2659 2383 2660 2387
rect 2654 2382 2660 2383
rect 2806 2387 2812 2388
rect 2806 2383 2807 2387
rect 2811 2383 2812 2387
rect 2806 2382 2812 2383
rect 2958 2387 2964 2388
rect 2958 2383 2959 2387
rect 2963 2383 2964 2387
rect 2958 2382 2964 2383
rect 3118 2387 3124 2388
rect 3118 2383 3119 2387
rect 3123 2383 3124 2387
rect 3118 2382 3124 2383
rect 158 2367 164 2368
rect 158 2363 159 2367
rect 163 2363 164 2367
rect 158 2362 164 2363
rect 246 2367 252 2368
rect 246 2363 247 2367
rect 251 2363 252 2367
rect 246 2362 252 2363
rect 334 2367 340 2368
rect 334 2363 335 2367
rect 339 2363 340 2367
rect 334 2362 340 2363
rect 438 2367 444 2368
rect 438 2363 439 2367
rect 443 2363 444 2367
rect 438 2362 444 2363
rect 558 2367 564 2368
rect 558 2363 559 2367
rect 563 2363 564 2367
rect 558 2362 564 2363
rect 686 2367 692 2368
rect 686 2363 687 2367
rect 691 2363 692 2367
rect 686 2362 692 2363
rect 814 2367 820 2368
rect 814 2363 815 2367
rect 819 2363 820 2367
rect 814 2362 820 2363
rect 950 2367 956 2368
rect 950 2363 951 2367
rect 955 2363 956 2367
rect 950 2362 956 2363
rect 1078 2367 1084 2368
rect 1078 2363 1079 2367
rect 1083 2363 1084 2367
rect 1078 2362 1084 2363
rect 1206 2367 1212 2368
rect 1206 2363 1207 2367
rect 1211 2363 1212 2367
rect 1206 2362 1212 2363
rect 1326 2367 1332 2368
rect 1326 2363 1327 2367
rect 1331 2363 1332 2367
rect 1326 2362 1332 2363
rect 1454 2367 1460 2368
rect 1454 2363 1455 2367
rect 1459 2363 1460 2367
rect 1454 2362 1460 2363
rect 1582 2367 1588 2368
rect 1582 2363 1583 2367
rect 1587 2363 1588 2367
rect 1582 2362 1588 2363
rect 110 2357 116 2358
rect 110 2353 111 2357
rect 115 2353 116 2357
rect 110 2352 116 2353
rect 1822 2357 1828 2358
rect 1822 2353 1823 2357
rect 1827 2353 1828 2357
rect 1822 2352 1828 2353
rect 1926 2349 1932 2350
rect 1926 2345 1927 2349
rect 1931 2345 1932 2349
rect 1926 2344 1932 2345
rect 2086 2349 2092 2350
rect 2086 2345 2087 2349
rect 2091 2345 2092 2349
rect 2086 2344 2092 2345
rect 2246 2349 2252 2350
rect 2246 2345 2247 2349
rect 2251 2345 2252 2349
rect 2246 2344 2252 2345
rect 2406 2349 2412 2350
rect 2406 2345 2407 2349
rect 2411 2345 2412 2349
rect 2406 2344 2412 2345
rect 2558 2349 2564 2350
rect 2558 2345 2559 2349
rect 2563 2345 2564 2349
rect 2558 2344 2564 2345
rect 2702 2349 2708 2350
rect 2702 2345 2703 2349
rect 2707 2345 2708 2349
rect 2702 2344 2708 2345
rect 2830 2349 2836 2350
rect 2830 2345 2831 2349
rect 2835 2345 2836 2349
rect 2830 2344 2836 2345
rect 2950 2349 2956 2350
rect 2950 2345 2951 2349
rect 2955 2345 2956 2349
rect 2950 2344 2956 2345
rect 3070 2349 3076 2350
rect 3070 2345 3071 2349
rect 3075 2345 3076 2349
rect 3070 2344 3076 2345
rect 3182 2349 3188 2350
rect 3182 2345 3183 2349
rect 3187 2345 3188 2349
rect 3182 2344 3188 2345
rect 3286 2349 3292 2350
rect 3286 2345 3287 2349
rect 3291 2345 3292 2349
rect 3286 2344 3292 2345
rect 3398 2349 3404 2350
rect 3398 2345 3399 2349
rect 3403 2345 3404 2349
rect 3398 2344 3404 2345
rect 3486 2349 3492 2350
rect 3486 2345 3487 2349
rect 3491 2345 3492 2349
rect 3486 2344 3492 2345
rect 110 2340 116 2341
rect 110 2336 111 2340
rect 115 2336 116 2340
rect 110 2335 116 2336
rect 1822 2340 1828 2341
rect 1822 2336 1823 2340
rect 1827 2336 1828 2340
rect 1822 2335 1828 2336
rect 1862 2336 1868 2337
rect 1862 2332 1863 2336
rect 1867 2332 1868 2336
rect 1862 2331 1868 2332
rect 3574 2336 3580 2337
rect 3574 2332 3575 2336
rect 3579 2332 3580 2336
rect 3574 2331 3580 2332
rect 166 2327 172 2328
rect 166 2323 167 2327
rect 171 2323 172 2327
rect 166 2322 172 2323
rect 254 2327 260 2328
rect 254 2323 255 2327
rect 259 2323 260 2327
rect 254 2322 260 2323
rect 342 2327 348 2328
rect 342 2323 343 2327
rect 347 2323 348 2327
rect 342 2322 348 2323
rect 446 2327 452 2328
rect 446 2323 447 2327
rect 451 2323 452 2327
rect 446 2322 452 2323
rect 566 2327 572 2328
rect 566 2323 567 2327
rect 571 2323 572 2327
rect 566 2322 572 2323
rect 694 2327 700 2328
rect 694 2323 695 2327
rect 699 2323 700 2327
rect 694 2322 700 2323
rect 822 2327 828 2328
rect 822 2323 823 2327
rect 827 2323 828 2327
rect 822 2322 828 2323
rect 958 2327 964 2328
rect 958 2323 959 2327
rect 963 2323 964 2327
rect 958 2322 964 2323
rect 1086 2327 1092 2328
rect 1086 2323 1087 2327
rect 1091 2323 1092 2327
rect 1086 2322 1092 2323
rect 1214 2327 1220 2328
rect 1214 2323 1215 2327
rect 1219 2323 1220 2327
rect 1214 2322 1220 2323
rect 1334 2327 1340 2328
rect 1334 2323 1335 2327
rect 1339 2323 1340 2327
rect 1334 2322 1340 2323
rect 1462 2327 1468 2328
rect 1462 2323 1463 2327
rect 1467 2323 1468 2327
rect 1462 2322 1468 2323
rect 1590 2327 1596 2328
rect 1590 2323 1591 2327
rect 1595 2323 1596 2327
rect 1590 2322 1596 2323
rect 1862 2319 1868 2320
rect 1862 2315 1863 2319
rect 1867 2315 1868 2319
rect 1862 2314 1868 2315
rect 3574 2319 3580 2320
rect 3574 2315 3575 2319
rect 3579 2315 3580 2319
rect 3574 2314 3580 2315
rect 1918 2309 1924 2310
rect 1918 2305 1919 2309
rect 1923 2305 1924 2309
rect 1918 2304 1924 2305
rect 2078 2309 2084 2310
rect 2078 2305 2079 2309
rect 2083 2305 2084 2309
rect 2078 2304 2084 2305
rect 2238 2309 2244 2310
rect 2238 2305 2239 2309
rect 2243 2305 2244 2309
rect 2238 2304 2244 2305
rect 2398 2309 2404 2310
rect 2398 2305 2399 2309
rect 2403 2305 2404 2309
rect 2398 2304 2404 2305
rect 2550 2309 2556 2310
rect 2550 2305 2551 2309
rect 2555 2305 2556 2309
rect 2550 2304 2556 2305
rect 2694 2309 2700 2310
rect 2694 2305 2695 2309
rect 2699 2305 2700 2309
rect 2694 2304 2700 2305
rect 2822 2309 2828 2310
rect 2822 2305 2823 2309
rect 2827 2305 2828 2309
rect 2822 2304 2828 2305
rect 2942 2309 2948 2310
rect 2942 2305 2943 2309
rect 2947 2305 2948 2309
rect 2942 2304 2948 2305
rect 3062 2309 3068 2310
rect 3062 2305 3063 2309
rect 3067 2305 3068 2309
rect 3062 2304 3068 2305
rect 3174 2309 3180 2310
rect 3174 2305 3175 2309
rect 3179 2305 3180 2309
rect 3174 2304 3180 2305
rect 3278 2309 3284 2310
rect 3278 2305 3279 2309
rect 3283 2305 3284 2309
rect 3278 2304 3284 2305
rect 3390 2309 3396 2310
rect 3390 2305 3391 2309
rect 3395 2305 3396 2309
rect 3390 2304 3396 2305
rect 3478 2309 3484 2310
rect 3478 2305 3479 2309
rect 3483 2305 3484 2309
rect 3478 2304 3484 2305
rect 694 2285 700 2286
rect 694 2281 695 2285
rect 699 2281 700 2285
rect 694 2280 700 2281
rect 862 2285 868 2286
rect 862 2281 863 2285
rect 867 2281 868 2285
rect 862 2280 868 2281
rect 1022 2285 1028 2286
rect 1022 2281 1023 2285
rect 1027 2281 1028 2285
rect 1022 2280 1028 2281
rect 1174 2285 1180 2286
rect 1174 2281 1175 2285
rect 1179 2281 1180 2285
rect 1174 2280 1180 2281
rect 1318 2285 1324 2286
rect 1318 2281 1319 2285
rect 1323 2281 1324 2285
rect 1318 2280 1324 2281
rect 1462 2285 1468 2286
rect 1462 2281 1463 2285
rect 1467 2281 1468 2285
rect 1462 2280 1468 2281
rect 1598 2285 1604 2286
rect 1598 2281 1599 2285
rect 1603 2281 1604 2285
rect 1598 2280 1604 2281
rect 1734 2285 1740 2286
rect 1734 2281 1735 2285
rect 1739 2281 1740 2285
rect 1734 2280 1740 2281
rect 1974 2283 1980 2284
rect 1974 2279 1975 2283
rect 1979 2279 1980 2283
rect 1974 2278 1980 2279
rect 2142 2283 2148 2284
rect 2142 2279 2143 2283
rect 2147 2279 2148 2283
rect 2142 2278 2148 2279
rect 2310 2283 2316 2284
rect 2310 2279 2311 2283
rect 2315 2279 2316 2283
rect 2310 2278 2316 2279
rect 2478 2283 2484 2284
rect 2478 2279 2479 2283
rect 2483 2279 2484 2283
rect 2478 2278 2484 2279
rect 2638 2283 2644 2284
rect 2638 2279 2639 2283
rect 2643 2279 2644 2283
rect 2638 2278 2644 2279
rect 2782 2283 2788 2284
rect 2782 2279 2783 2283
rect 2787 2279 2788 2283
rect 2782 2278 2788 2279
rect 2918 2283 2924 2284
rect 2918 2279 2919 2283
rect 2923 2279 2924 2283
rect 2918 2278 2924 2279
rect 3038 2283 3044 2284
rect 3038 2279 3039 2283
rect 3043 2279 3044 2283
rect 3038 2278 3044 2279
rect 3158 2283 3164 2284
rect 3158 2279 3159 2283
rect 3163 2279 3164 2283
rect 3158 2278 3164 2279
rect 3270 2283 3276 2284
rect 3270 2279 3271 2283
rect 3275 2279 3276 2283
rect 3270 2278 3276 2279
rect 3382 2283 3388 2284
rect 3382 2279 3383 2283
rect 3387 2279 3388 2283
rect 3382 2278 3388 2279
rect 3478 2283 3484 2284
rect 3478 2279 3479 2283
rect 3483 2279 3484 2283
rect 3478 2278 3484 2279
rect 1862 2273 1868 2274
rect 110 2272 116 2273
rect 110 2268 111 2272
rect 115 2268 116 2272
rect 110 2267 116 2268
rect 1822 2272 1828 2273
rect 1822 2268 1823 2272
rect 1827 2268 1828 2272
rect 1862 2269 1863 2273
rect 1867 2269 1868 2273
rect 1862 2268 1868 2269
rect 3574 2273 3580 2274
rect 3574 2269 3575 2273
rect 3579 2269 3580 2273
rect 3574 2268 3580 2269
rect 1822 2267 1828 2268
rect 1862 2256 1868 2257
rect 110 2255 116 2256
rect 110 2251 111 2255
rect 115 2251 116 2255
rect 110 2250 116 2251
rect 1822 2255 1828 2256
rect 1822 2251 1823 2255
rect 1827 2251 1828 2255
rect 1862 2252 1863 2256
rect 1867 2252 1868 2256
rect 1862 2251 1868 2252
rect 3574 2256 3580 2257
rect 3574 2252 3575 2256
rect 3579 2252 3580 2256
rect 3574 2251 3580 2252
rect 1822 2250 1828 2251
rect 686 2245 692 2246
rect 686 2241 687 2245
rect 691 2241 692 2245
rect 686 2240 692 2241
rect 854 2245 860 2246
rect 854 2241 855 2245
rect 859 2241 860 2245
rect 854 2240 860 2241
rect 1014 2245 1020 2246
rect 1014 2241 1015 2245
rect 1019 2241 1020 2245
rect 1014 2240 1020 2241
rect 1166 2245 1172 2246
rect 1166 2241 1167 2245
rect 1171 2241 1172 2245
rect 1166 2240 1172 2241
rect 1310 2245 1316 2246
rect 1310 2241 1311 2245
rect 1315 2241 1316 2245
rect 1310 2240 1316 2241
rect 1454 2245 1460 2246
rect 1454 2241 1455 2245
rect 1459 2241 1460 2245
rect 1454 2240 1460 2241
rect 1590 2245 1596 2246
rect 1590 2241 1591 2245
rect 1595 2241 1596 2245
rect 1590 2240 1596 2241
rect 1726 2245 1732 2246
rect 1726 2241 1727 2245
rect 1731 2241 1732 2245
rect 1726 2240 1732 2241
rect 1982 2243 1988 2244
rect 1982 2239 1983 2243
rect 1987 2239 1988 2243
rect 1982 2238 1988 2239
rect 2150 2243 2156 2244
rect 2150 2239 2151 2243
rect 2155 2239 2156 2243
rect 2150 2238 2156 2239
rect 2318 2243 2324 2244
rect 2318 2239 2319 2243
rect 2323 2239 2324 2243
rect 2318 2238 2324 2239
rect 2486 2243 2492 2244
rect 2486 2239 2487 2243
rect 2491 2239 2492 2243
rect 2486 2238 2492 2239
rect 2646 2243 2652 2244
rect 2646 2239 2647 2243
rect 2651 2239 2652 2243
rect 2646 2238 2652 2239
rect 2790 2243 2796 2244
rect 2790 2239 2791 2243
rect 2795 2239 2796 2243
rect 2790 2238 2796 2239
rect 2926 2243 2932 2244
rect 2926 2239 2927 2243
rect 2931 2239 2932 2243
rect 2926 2238 2932 2239
rect 3046 2243 3052 2244
rect 3046 2239 3047 2243
rect 3051 2239 3052 2243
rect 3046 2238 3052 2239
rect 3166 2243 3172 2244
rect 3166 2239 3167 2243
rect 3171 2239 3172 2243
rect 3166 2238 3172 2239
rect 3278 2243 3284 2244
rect 3278 2239 3279 2243
rect 3283 2239 3284 2243
rect 3278 2238 3284 2239
rect 3390 2243 3396 2244
rect 3390 2239 3391 2243
rect 3395 2239 3396 2243
rect 3390 2238 3396 2239
rect 3486 2243 3492 2244
rect 3486 2239 3487 2243
rect 3491 2239 3492 2243
rect 3486 2238 3492 2239
rect 534 2215 540 2216
rect 534 2211 535 2215
rect 539 2211 540 2215
rect 534 2210 540 2211
rect 718 2215 724 2216
rect 718 2211 719 2215
rect 723 2211 724 2215
rect 718 2210 724 2211
rect 894 2215 900 2216
rect 894 2211 895 2215
rect 899 2211 900 2215
rect 894 2210 900 2211
rect 1070 2215 1076 2216
rect 1070 2211 1071 2215
rect 1075 2211 1076 2215
rect 1070 2210 1076 2211
rect 1238 2215 1244 2216
rect 1238 2211 1239 2215
rect 1243 2211 1244 2215
rect 1238 2210 1244 2211
rect 1406 2215 1412 2216
rect 1406 2211 1407 2215
rect 1411 2211 1412 2215
rect 1406 2210 1412 2211
rect 1574 2215 1580 2216
rect 1574 2211 1575 2215
rect 1579 2211 1580 2215
rect 1574 2210 1580 2211
rect 1726 2215 1732 2216
rect 1726 2211 1727 2215
rect 1731 2211 1732 2215
rect 1726 2210 1732 2211
rect 2006 2209 2012 2210
rect 110 2205 116 2206
rect 110 2201 111 2205
rect 115 2201 116 2205
rect 110 2200 116 2201
rect 1822 2205 1828 2206
rect 1822 2201 1823 2205
rect 1827 2201 1828 2205
rect 2006 2205 2007 2209
rect 2011 2205 2012 2209
rect 2006 2204 2012 2205
rect 2166 2209 2172 2210
rect 2166 2205 2167 2209
rect 2171 2205 2172 2209
rect 2166 2204 2172 2205
rect 2334 2209 2340 2210
rect 2334 2205 2335 2209
rect 2339 2205 2340 2209
rect 2334 2204 2340 2205
rect 2518 2209 2524 2210
rect 2518 2205 2519 2209
rect 2523 2205 2524 2209
rect 2518 2204 2524 2205
rect 2710 2209 2716 2210
rect 2710 2205 2711 2209
rect 2715 2205 2716 2209
rect 2710 2204 2716 2205
rect 2902 2209 2908 2210
rect 2902 2205 2903 2209
rect 2907 2205 2908 2209
rect 2902 2204 2908 2205
rect 3102 2209 3108 2210
rect 3102 2205 3103 2209
rect 3107 2205 3108 2209
rect 3102 2204 3108 2205
rect 3302 2209 3308 2210
rect 3302 2205 3303 2209
rect 3307 2205 3308 2209
rect 3302 2204 3308 2205
rect 3486 2209 3492 2210
rect 3486 2205 3487 2209
rect 3491 2205 3492 2209
rect 3486 2204 3492 2205
rect 1822 2200 1828 2201
rect 1862 2196 1868 2197
rect 1862 2192 1863 2196
rect 1867 2192 1868 2196
rect 1862 2191 1868 2192
rect 3574 2196 3580 2197
rect 3574 2192 3575 2196
rect 3579 2192 3580 2196
rect 3574 2191 3580 2192
rect 110 2188 116 2189
rect 110 2184 111 2188
rect 115 2184 116 2188
rect 110 2183 116 2184
rect 1822 2188 1828 2189
rect 1822 2184 1823 2188
rect 1827 2184 1828 2188
rect 1822 2183 1828 2184
rect 1862 2179 1868 2180
rect 542 2175 548 2176
rect 542 2171 543 2175
rect 547 2171 548 2175
rect 542 2170 548 2171
rect 726 2175 732 2176
rect 726 2171 727 2175
rect 731 2171 732 2175
rect 726 2170 732 2171
rect 902 2175 908 2176
rect 902 2171 903 2175
rect 907 2171 908 2175
rect 902 2170 908 2171
rect 1078 2175 1084 2176
rect 1078 2171 1079 2175
rect 1083 2171 1084 2175
rect 1078 2170 1084 2171
rect 1246 2175 1252 2176
rect 1246 2171 1247 2175
rect 1251 2171 1252 2175
rect 1246 2170 1252 2171
rect 1414 2175 1420 2176
rect 1414 2171 1415 2175
rect 1419 2171 1420 2175
rect 1414 2170 1420 2171
rect 1582 2175 1588 2176
rect 1582 2171 1583 2175
rect 1587 2171 1588 2175
rect 1582 2170 1588 2171
rect 1734 2175 1740 2176
rect 1734 2171 1735 2175
rect 1739 2171 1740 2175
rect 1862 2175 1863 2179
rect 1867 2175 1868 2179
rect 1862 2174 1868 2175
rect 3574 2179 3580 2180
rect 3574 2175 3575 2179
rect 3579 2175 3580 2179
rect 3574 2174 3580 2175
rect 1734 2170 1740 2171
rect 1998 2169 2004 2170
rect 1998 2165 1999 2169
rect 2003 2165 2004 2169
rect 1998 2164 2004 2165
rect 2158 2169 2164 2170
rect 2158 2165 2159 2169
rect 2163 2165 2164 2169
rect 2158 2164 2164 2165
rect 2326 2169 2332 2170
rect 2326 2165 2327 2169
rect 2331 2165 2332 2169
rect 2326 2164 2332 2165
rect 2510 2169 2516 2170
rect 2510 2165 2511 2169
rect 2515 2165 2516 2169
rect 2510 2164 2516 2165
rect 2702 2169 2708 2170
rect 2702 2165 2703 2169
rect 2707 2165 2708 2169
rect 2702 2164 2708 2165
rect 2894 2169 2900 2170
rect 2894 2165 2895 2169
rect 2899 2165 2900 2169
rect 2894 2164 2900 2165
rect 3094 2169 3100 2170
rect 3094 2165 3095 2169
rect 3099 2165 3100 2169
rect 3094 2164 3100 2165
rect 3294 2169 3300 2170
rect 3294 2165 3295 2169
rect 3299 2165 3300 2169
rect 3294 2164 3300 2165
rect 3478 2169 3484 2170
rect 3478 2165 3479 2169
rect 3483 2165 3484 2169
rect 3478 2164 3484 2165
rect 494 2141 500 2142
rect 494 2137 495 2141
rect 499 2137 500 2141
rect 494 2136 500 2137
rect 622 2141 628 2142
rect 622 2137 623 2141
rect 627 2137 628 2141
rect 622 2136 628 2137
rect 758 2141 764 2142
rect 758 2137 759 2141
rect 763 2137 764 2141
rect 758 2136 764 2137
rect 894 2141 900 2142
rect 894 2137 895 2141
rect 899 2137 900 2141
rect 894 2136 900 2137
rect 1038 2141 1044 2142
rect 1038 2137 1039 2141
rect 1043 2137 1044 2141
rect 1038 2136 1044 2137
rect 1182 2141 1188 2142
rect 1182 2137 1183 2141
rect 1187 2137 1188 2141
rect 1182 2136 1188 2137
rect 1326 2141 1332 2142
rect 1326 2137 1327 2141
rect 1331 2137 1332 2141
rect 1326 2136 1332 2137
rect 1470 2141 1476 2142
rect 1470 2137 1471 2141
rect 1475 2137 1476 2141
rect 1470 2136 1476 2137
rect 1622 2141 1628 2142
rect 1622 2137 1623 2141
rect 1627 2137 1628 2141
rect 1622 2136 1628 2137
rect 2022 2139 2028 2140
rect 2022 2135 2023 2139
rect 2027 2135 2028 2139
rect 2022 2134 2028 2135
rect 2166 2139 2172 2140
rect 2166 2135 2167 2139
rect 2171 2135 2172 2139
rect 2166 2134 2172 2135
rect 2318 2139 2324 2140
rect 2318 2135 2319 2139
rect 2323 2135 2324 2139
rect 2318 2134 2324 2135
rect 2470 2139 2476 2140
rect 2470 2135 2471 2139
rect 2475 2135 2476 2139
rect 2470 2134 2476 2135
rect 2614 2139 2620 2140
rect 2614 2135 2615 2139
rect 2619 2135 2620 2139
rect 2614 2134 2620 2135
rect 2758 2139 2764 2140
rect 2758 2135 2759 2139
rect 2763 2135 2764 2139
rect 2758 2134 2764 2135
rect 2894 2139 2900 2140
rect 2894 2135 2895 2139
rect 2899 2135 2900 2139
rect 2894 2134 2900 2135
rect 3022 2139 3028 2140
rect 3022 2135 3023 2139
rect 3027 2135 3028 2139
rect 3022 2134 3028 2135
rect 3142 2139 3148 2140
rect 3142 2135 3143 2139
rect 3147 2135 3148 2139
rect 3142 2134 3148 2135
rect 3262 2139 3268 2140
rect 3262 2135 3263 2139
rect 3267 2135 3268 2139
rect 3262 2134 3268 2135
rect 3382 2139 3388 2140
rect 3382 2135 3383 2139
rect 3387 2135 3388 2139
rect 3382 2134 3388 2135
rect 3478 2139 3484 2140
rect 3478 2135 3479 2139
rect 3483 2135 3484 2139
rect 3478 2134 3484 2135
rect 1862 2129 1868 2130
rect 110 2128 116 2129
rect 110 2124 111 2128
rect 115 2124 116 2128
rect 110 2123 116 2124
rect 1822 2128 1828 2129
rect 1822 2124 1823 2128
rect 1827 2124 1828 2128
rect 1862 2125 1863 2129
rect 1867 2125 1868 2129
rect 1862 2124 1868 2125
rect 3574 2129 3580 2130
rect 3574 2125 3575 2129
rect 3579 2125 3580 2129
rect 3574 2124 3580 2125
rect 1822 2123 1828 2124
rect 1862 2112 1868 2113
rect 110 2111 116 2112
rect 110 2107 111 2111
rect 115 2107 116 2111
rect 110 2106 116 2107
rect 1822 2111 1828 2112
rect 1822 2107 1823 2111
rect 1827 2107 1828 2111
rect 1862 2108 1863 2112
rect 1867 2108 1868 2112
rect 1862 2107 1868 2108
rect 3574 2112 3580 2113
rect 3574 2108 3575 2112
rect 3579 2108 3580 2112
rect 3574 2107 3580 2108
rect 1822 2106 1828 2107
rect 486 2101 492 2102
rect 486 2097 487 2101
rect 491 2097 492 2101
rect 486 2096 492 2097
rect 614 2101 620 2102
rect 614 2097 615 2101
rect 619 2097 620 2101
rect 614 2096 620 2097
rect 750 2101 756 2102
rect 750 2097 751 2101
rect 755 2097 756 2101
rect 750 2096 756 2097
rect 886 2101 892 2102
rect 886 2097 887 2101
rect 891 2097 892 2101
rect 886 2096 892 2097
rect 1030 2101 1036 2102
rect 1030 2097 1031 2101
rect 1035 2097 1036 2101
rect 1030 2096 1036 2097
rect 1174 2101 1180 2102
rect 1174 2097 1175 2101
rect 1179 2097 1180 2101
rect 1174 2096 1180 2097
rect 1318 2101 1324 2102
rect 1318 2097 1319 2101
rect 1323 2097 1324 2101
rect 1318 2096 1324 2097
rect 1462 2101 1468 2102
rect 1462 2097 1463 2101
rect 1467 2097 1468 2101
rect 1462 2096 1468 2097
rect 1614 2101 1620 2102
rect 1614 2097 1615 2101
rect 1619 2097 1620 2101
rect 1614 2096 1620 2097
rect 2030 2099 2036 2100
rect 2030 2095 2031 2099
rect 2035 2095 2036 2099
rect 2030 2094 2036 2095
rect 2174 2099 2180 2100
rect 2174 2095 2175 2099
rect 2179 2095 2180 2099
rect 2174 2094 2180 2095
rect 2326 2099 2332 2100
rect 2326 2095 2327 2099
rect 2331 2095 2332 2099
rect 2326 2094 2332 2095
rect 2478 2099 2484 2100
rect 2478 2095 2479 2099
rect 2483 2095 2484 2099
rect 2478 2094 2484 2095
rect 2622 2099 2628 2100
rect 2622 2095 2623 2099
rect 2627 2095 2628 2099
rect 2622 2094 2628 2095
rect 2766 2099 2772 2100
rect 2766 2095 2767 2099
rect 2771 2095 2772 2099
rect 2766 2094 2772 2095
rect 2902 2099 2908 2100
rect 2902 2095 2903 2099
rect 2907 2095 2908 2099
rect 2902 2094 2908 2095
rect 3030 2099 3036 2100
rect 3030 2095 3031 2099
rect 3035 2095 3036 2099
rect 3030 2094 3036 2095
rect 3150 2099 3156 2100
rect 3150 2095 3151 2099
rect 3155 2095 3156 2099
rect 3150 2094 3156 2095
rect 3270 2099 3276 2100
rect 3270 2095 3271 2099
rect 3275 2095 3276 2099
rect 3270 2094 3276 2095
rect 3390 2099 3396 2100
rect 3390 2095 3391 2099
rect 3395 2095 3396 2099
rect 3390 2094 3396 2095
rect 3486 2099 3492 2100
rect 3486 2095 3487 2099
rect 3491 2095 3492 2099
rect 3486 2094 3492 2095
rect 318 2075 324 2076
rect 318 2071 319 2075
rect 323 2071 324 2075
rect 318 2070 324 2071
rect 430 2075 436 2076
rect 430 2071 431 2075
rect 435 2071 436 2075
rect 430 2070 436 2071
rect 550 2075 556 2076
rect 550 2071 551 2075
rect 555 2071 556 2075
rect 550 2070 556 2071
rect 678 2075 684 2076
rect 678 2071 679 2075
rect 683 2071 684 2075
rect 678 2070 684 2071
rect 798 2075 804 2076
rect 798 2071 799 2075
rect 803 2071 804 2075
rect 798 2070 804 2071
rect 918 2075 924 2076
rect 918 2071 919 2075
rect 923 2071 924 2075
rect 918 2070 924 2071
rect 1038 2075 1044 2076
rect 1038 2071 1039 2075
rect 1043 2071 1044 2075
rect 1038 2070 1044 2071
rect 1158 2075 1164 2076
rect 1158 2071 1159 2075
rect 1163 2071 1164 2075
rect 1158 2070 1164 2071
rect 1278 2075 1284 2076
rect 1278 2071 1279 2075
rect 1283 2071 1284 2075
rect 1278 2070 1284 2071
rect 1406 2075 1412 2076
rect 1406 2071 1407 2075
rect 1411 2071 1412 2075
rect 1406 2070 1412 2071
rect 110 2065 116 2066
rect 110 2061 111 2065
rect 115 2061 116 2065
rect 110 2060 116 2061
rect 1822 2065 1828 2066
rect 1822 2061 1823 2065
rect 1827 2061 1828 2065
rect 1822 2060 1828 2061
rect 1982 2061 1988 2062
rect 1982 2057 1983 2061
rect 1987 2057 1988 2061
rect 1982 2056 1988 2057
rect 2142 2061 2148 2062
rect 2142 2057 2143 2061
rect 2147 2057 2148 2061
rect 2142 2056 2148 2057
rect 2310 2061 2316 2062
rect 2310 2057 2311 2061
rect 2315 2057 2316 2061
rect 2310 2056 2316 2057
rect 2470 2061 2476 2062
rect 2470 2057 2471 2061
rect 2475 2057 2476 2061
rect 2470 2056 2476 2057
rect 2630 2061 2636 2062
rect 2630 2057 2631 2061
rect 2635 2057 2636 2061
rect 2630 2056 2636 2057
rect 2774 2061 2780 2062
rect 2774 2057 2775 2061
rect 2779 2057 2780 2061
rect 2774 2056 2780 2057
rect 2910 2061 2916 2062
rect 2910 2057 2911 2061
rect 2915 2057 2916 2061
rect 2910 2056 2916 2057
rect 3038 2061 3044 2062
rect 3038 2057 3039 2061
rect 3043 2057 3044 2061
rect 3038 2056 3044 2057
rect 3158 2061 3164 2062
rect 3158 2057 3159 2061
rect 3163 2057 3164 2061
rect 3158 2056 3164 2057
rect 3278 2061 3284 2062
rect 3278 2057 3279 2061
rect 3283 2057 3284 2061
rect 3278 2056 3284 2057
rect 3390 2061 3396 2062
rect 3390 2057 3391 2061
rect 3395 2057 3396 2061
rect 3390 2056 3396 2057
rect 3486 2061 3492 2062
rect 3486 2057 3487 2061
rect 3491 2057 3492 2061
rect 3486 2056 3492 2057
rect 110 2048 116 2049
rect 110 2044 111 2048
rect 115 2044 116 2048
rect 110 2043 116 2044
rect 1822 2048 1828 2049
rect 1822 2044 1823 2048
rect 1827 2044 1828 2048
rect 1822 2043 1828 2044
rect 1862 2048 1868 2049
rect 1862 2044 1863 2048
rect 1867 2044 1868 2048
rect 1862 2043 1868 2044
rect 3574 2048 3580 2049
rect 3574 2044 3575 2048
rect 3579 2044 3580 2048
rect 3574 2043 3580 2044
rect 326 2035 332 2036
rect 326 2031 327 2035
rect 331 2031 332 2035
rect 326 2030 332 2031
rect 438 2035 444 2036
rect 438 2031 439 2035
rect 443 2031 444 2035
rect 438 2030 444 2031
rect 558 2035 564 2036
rect 558 2031 559 2035
rect 563 2031 564 2035
rect 558 2030 564 2031
rect 686 2035 692 2036
rect 686 2031 687 2035
rect 691 2031 692 2035
rect 686 2030 692 2031
rect 806 2035 812 2036
rect 806 2031 807 2035
rect 811 2031 812 2035
rect 806 2030 812 2031
rect 926 2035 932 2036
rect 926 2031 927 2035
rect 931 2031 932 2035
rect 926 2030 932 2031
rect 1046 2035 1052 2036
rect 1046 2031 1047 2035
rect 1051 2031 1052 2035
rect 1046 2030 1052 2031
rect 1166 2035 1172 2036
rect 1166 2031 1167 2035
rect 1171 2031 1172 2035
rect 1166 2030 1172 2031
rect 1286 2035 1292 2036
rect 1286 2031 1287 2035
rect 1291 2031 1292 2035
rect 1286 2030 1292 2031
rect 1414 2035 1420 2036
rect 1414 2031 1415 2035
rect 1419 2031 1420 2035
rect 1414 2030 1420 2031
rect 1862 2031 1868 2032
rect 1862 2027 1863 2031
rect 1867 2027 1868 2031
rect 1862 2026 1868 2027
rect 3574 2031 3580 2032
rect 3574 2027 3575 2031
rect 3579 2027 3580 2031
rect 3574 2026 3580 2027
rect 1974 2021 1980 2022
rect 1974 2017 1975 2021
rect 1979 2017 1980 2021
rect 1974 2016 1980 2017
rect 2134 2021 2140 2022
rect 2134 2017 2135 2021
rect 2139 2017 2140 2021
rect 2134 2016 2140 2017
rect 2302 2021 2308 2022
rect 2302 2017 2303 2021
rect 2307 2017 2308 2021
rect 2302 2016 2308 2017
rect 2462 2021 2468 2022
rect 2462 2017 2463 2021
rect 2467 2017 2468 2021
rect 2462 2016 2468 2017
rect 2622 2021 2628 2022
rect 2622 2017 2623 2021
rect 2627 2017 2628 2021
rect 2622 2016 2628 2017
rect 2766 2021 2772 2022
rect 2766 2017 2767 2021
rect 2771 2017 2772 2021
rect 2766 2016 2772 2017
rect 2902 2021 2908 2022
rect 2902 2017 2903 2021
rect 2907 2017 2908 2021
rect 2902 2016 2908 2017
rect 3030 2021 3036 2022
rect 3030 2017 3031 2021
rect 3035 2017 3036 2021
rect 3030 2016 3036 2017
rect 3150 2021 3156 2022
rect 3150 2017 3151 2021
rect 3155 2017 3156 2021
rect 3150 2016 3156 2017
rect 3270 2021 3276 2022
rect 3270 2017 3271 2021
rect 3275 2017 3276 2021
rect 3270 2016 3276 2017
rect 3382 2021 3388 2022
rect 3382 2017 3383 2021
rect 3387 2017 3388 2021
rect 3382 2016 3388 2017
rect 3478 2021 3484 2022
rect 3478 2017 3479 2021
rect 3483 2017 3484 2021
rect 3478 2016 3484 2017
rect 1886 1999 1892 2000
rect 182 1997 188 1998
rect 182 1993 183 1997
rect 187 1993 188 1997
rect 182 1992 188 1993
rect 294 1997 300 1998
rect 294 1993 295 1997
rect 299 1993 300 1997
rect 294 1992 300 1993
rect 414 1997 420 1998
rect 414 1993 415 1997
rect 419 1993 420 1997
rect 414 1992 420 1993
rect 534 1997 540 1998
rect 534 1993 535 1997
rect 539 1993 540 1997
rect 534 1992 540 1993
rect 654 1997 660 1998
rect 654 1993 655 1997
rect 659 1993 660 1997
rect 654 1992 660 1993
rect 774 1997 780 1998
rect 774 1993 775 1997
rect 779 1993 780 1997
rect 774 1992 780 1993
rect 894 1997 900 1998
rect 894 1993 895 1997
rect 899 1993 900 1997
rect 894 1992 900 1993
rect 1014 1997 1020 1998
rect 1014 1993 1015 1997
rect 1019 1993 1020 1997
rect 1014 1992 1020 1993
rect 1134 1997 1140 1998
rect 1134 1993 1135 1997
rect 1139 1993 1140 1997
rect 1134 1992 1140 1993
rect 1254 1997 1260 1998
rect 1254 1993 1255 1997
rect 1259 1993 1260 1997
rect 1886 1995 1887 1999
rect 1891 1995 1892 1999
rect 1886 1994 1892 1995
rect 2030 1999 2036 2000
rect 2030 1995 2031 1999
rect 2035 1995 2036 1999
rect 2030 1994 2036 1995
rect 2198 1999 2204 2000
rect 2198 1995 2199 1999
rect 2203 1995 2204 1999
rect 2198 1994 2204 1995
rect 2374 1999 2380 2000
rect 2374 1995 2375 1999
rect 2379 1995 2380 1999
rect 2374 1994 2380 1995
rect 2542 1999 2548 2000
rect 2542 1995 2543 1999
rect 2547 1995 2548 1999
rect 2542 1994 2548 1995
rect 2710 1999 2716 2000
rect 2710 1995 2711 1999
rect 2715 1995 2716 1999
rect 2710 1994 2716 1995
rect 2870 1999 2876 2000
rect 2870 1995 2871 1999
rect 2875 1995 2876 1999
rect 2870 1994 2876 1995
rect 3038 1999 3044 2000
rect 3038 1995 3039 1999
rect 3043 1995 3044 1999
rect 3038 1994 3044 1995
rect 3206 1999 3212 2000
rect 3206 1995 3207 1999
rect 3211 1995 3212 1999
rect 3206 1994 3212 1995
rect 1254 1992 1260 1993
rect 1862 1989 1868 1990
rect 1862 1985 1863 1989
rect 1867 1985 1868 1989
rect 110 1984 116 1985
rect 110 1980 111 1984
rect 115 1980 116 1984
rect 110 1979 116 1980
rect 1822 1984 1828 1985
rect 1862 1984 1868 1985
rect 3574 1989 3580 1990
rect 3574 1985 3575 1989
rect 3579 1985 3580 1989
rect 3574 1984 3580 1985
rect 1822 1980 1823 1984
rect 1827 1980 1828 1984
rect 1822 1979 1828 1980
rect 1862 1972 1868 1973
rect 1862 1968 1863 1972
rect 1867 1968 1868 1972
rect 110 1967 116 1968
rect 110 1963 111 1967
rect 115 1963 116 1967
rect 110 1962 116 1963
rect 1822 1967 1828 1968
rect 1862 1967 1868 1968
rect 3574 1972 3580 1973
rect 3574 1968 3575 1972
rect 3579 1968 3580 1972
rect 3574 1967 3580 1968
rect 1822 1963 1823 1967
rect 1827 1963 1828 1967
rect 1822 1962 1828 1963
rect 1894 1959 1900 1960
rect 174 1957 180 1958
rect 174 1953 175 1957
rect 179 1953 180 1957
rect 174 1952 180 1953
rect 286 1957 292 1958
rect 286 1953 287 1957
rect 291 1953 292 1957
rect 286 1952 292 1953
rect 406 1957 412 1958
rect 406 1953 407 1957
rect 411 1953 412 1957
rect 406 1952 412 1953
rect 526 1957 532 1958
rect 526 1953 527 1957
rect 531 1953 532 1957
rect 526 1952 532 1953
rect 646 1957 652 1958
rect 646 1953 647 1957
rect 651 1953 652 1957
rect 646 1952 652 1953
rect 766 1957 772 1958
rect 766 1953 767 1957
rect 771 1953 772 1957
rect 766 1952 772 1953
rect 886 1957 892 1958
rect 886 1953 887 1957
rect 891 1953 892 1957
rect 886 1952 892 1953
rect 1006 1957 1012 1958
rect 1006 1953 1007 1957
rect 1011 1953 1012 1957
rect 1006 1952 1012 1953
rect 1126 1957 1132 1958
rect 1126 1953 1127 1957
rect 1131 1953 1132 1957
rect 1126 1952 1132 1953
rect 1246 1957 1252 1958
rect 1246 1953 1247 1957
rect 1251 1953 1252 1957
rect 1894 1955 1895 1959
rect 1899 1955 1900 1959
rect 1894 1954 1900 1955
rect 2038 1959 2044 1960
rect 2038 1955 2039 1959
rect 2043 1955 2044 1959
rect 2038 1954 2044 1955
rect 2206 1959 2212 1960
rect 2206 1955 2207 1959
rect 2211 1955 2212 1959
rect 2206 1954 2212 1955
rect 2382 1959 2388 1960
rect 2382 1955 2383 1959
rect 2387 1955 2388 1959
rect 2382 1954 2388 1955
rect 2550 1959 2556 1960
rect 2550 1955 2551 1959
rect 2555 1955 2556 1959
rect 2550 1954 2556 1955
rect 2718 1959 2724 1960
rect 2718 1955 2719 1959
rect 2723 1955 2724 1959
rect 2718 1954 2724 1955
rect 2878 1959 2884 1960
rect 2878 1955 2879 1959
rect 2883 1955 2884 1959
rect 2878 1954 2884 1955
rect 3046 1959 3052 1960
rect 3046 1955 3047 1959
rect 3051 1955 3052 1959
rect 3046 1954 3052 1955
rect 3214 1959 3220 1960
rect 3214 1955 3215 1959
rect 3219 1955 3220 1959
rect 3214 1954 3220 1955
rect 1246 1952 1252 1953
rect 134 1931 140 1932
rect 134 1927 135 1931
rect 139 1927 140 1931
rect 134 1926 140 1927
rect 222 1931 228 1932
rect 222 1927 223 1931
rect 227 1927 228 1931
rect 222 1926 228 1927
rect 350 1931 356 1932
rect 350 1927 351 1931
rect 355 1927 356 1931
rect 350 1926 356 1927
rect 494 1931 500 1932
rect 494 1927 495 1931
rect 499 1927 500 1931
rect 494 1926 500 1927
rect 654 1931 660 1932
rect 654 1927 655 1931
rect 659 1927 660 1931
rect 654 1926 660 1927
rect 838 1931 844 1932
rect 838 1927 839 1931
rect 843 1927 844 1931
rect 838 1926 844 1927
rect 1038 1931 1044 1932
rect 1038 1927 1039 1931
rect 1043 1927 1044 1931
rect 1038 1926 1044 1927
rect 1246 1931 1252 1932
rect 1246 1927 1247 1931
rect 1251 1927 1252 1931
rect 1246 1926 1252 1927
rect 1462 1931 1468 1932
rect 1462 1927 1463 1931
rect 1467 1927 1468 1931
rect 1462 1926 1468 1927
rect 110 1921 116 1922
rect 110 1917 111 1921
rect 115 1917 116 1921
rect 110 1916 116 1917
rect 1822 1921 1828 1922
rect 1822 1917 1823 1921
rect 1827 1917 1828 1921
rect 1822 1916 1828 1917
rect 1894 1917 1900 1918
rect 1894 1913 1895 1917
rect 1899 1913 1900 1917
rect 1894 1912 1900 1913
rect 1990 1917 1996 1918
rect 1990 1913 1991 1917
rect 1995 1913 1996 1917
rect 1990 1912 1996 1913
rect 2118 1917 2124 1918
rect 2118 1913 2119 1917
rect 2123 1913 2124 1917
rect 2118 1912 2124 1913
rect 2254 1917 2260 1918
rect 2254 1913 2255 1917
rect 2259 1913 2260 1917
rect 2254 1912 2260 1913
rect 2382 1917 2388 1918
rect 2382 1913 2383 1917
rect 2387 1913 2388 1917
rect 2382 1912 2388 1913
rect 2510 1917 2516 1918
rect 2510 1913 2511 1917
rect 2515 1913 2516 1917
rect 2510 1912 2516 1913
rect 2630 1917 2636 1918
rect 2630 1913 2631 1917
rect 2635 1913 2636 1917
rect 2630 1912 2636 1913
rect 2750 1917 2756 1918
rect 2750 1913 2751 1917
rect 2755 1913 2756 1917
rect 2750 1912 2756 1913
rect 2878 1917 2884 1918
rect 2878 1913 2879 1917
rect 2883 1913 2884 1917
rect 2878 1912 2884 1913
rect 3006 1917 3012 1918
rect 3006 1913 3007 1917
rect 3011 1913 3012 1917
rect 3006 1912 3012 1913
rect 110 1904 116 1905
rect 110 1900 111 1904
rect 115 1900 116 1904
rect 110 1899 116 1900
rect 1822 1904 1828 1905
rect 1822 1900 1823 1904
rect 1827 1900 1828 1904
rect 1822 1899 1828 1900
rect 1862 1904 1868 1905
rect 1862 1900 1863 1904
rect 1867 1900 1868 1904
rect 1862 1899 1868 1900
rect 3574 1904 3580 1905
rect 3574 1900 3575 1904
rect 3579 1900 3580 1904
rect 3574 1899 3580 1900
rect 142 1891 148 1892
rect 142 1887 143 1891
rect 147 1887 148 1891
rect 142 1886 148 1887
rect 230 1891 236 1892
rect 230 1887 231 1891
rect 235 1887 236 1891
rect 230 1886 236 1887
rect 358 1891 364 1892
rect 358 1887 359 1891
rect 363 1887 364 1891
rect 358 1886 364 1887
rect 502 1891 508 1892
rect 502 1887 503 1891
rect 507 1887 508 1891
rect 502 1886 508 1887
rect 662 1891 668 1892
rect 662 1887 663 1891
rect 667 1887 668 1891
rect 662 1886 668 1887
rect 846 1891 852 1892
rect 846 1887 847 1891
rect 851 1887 852 1891
rect 846 1886 852 1887
rect 1046 1891 1052 1892
rect 1046 1887 1047 1891
rect 1051 1887 1052 1891
rect 1046 1886 1052 1887
rect 1254 1891 1260 1892
rect 1254 1887 1255 1891
rect 1259 1887 1260 1891
rect 1254 1886 1260 1887
rect 1470 1891 1476 1892
rect 1470 1887 1471 1891
rect 1475 1887 1476 1891
rect 1470 1886 1476 1887
rect 1862 1887 1868 1888
rect 1862 1883 1863 1887
rect 1867 1883 1868 1887
rect 1862 1882 1868 1883
rect 3574 1887 3580 1888
rect 3574 1883 3575 1887
rect 3579 1883 3580 1887
rect 3574 1882 3580 1883
rect 1886 1877 1892 1878
rect 1886 1873 1887 1877
rect 1891 1873 1892 1877
rect 1886 1872 1892 1873
rect 1982 1877 1988 1878
rect 1982 1873 1983 1877
rect 1987 1873 1988 1877
rect 1982 1872 1988 1873
rect 2110 1877 2116 1878
rect 2110 1873 2111 1877
rect 2115 1873 2116 1877
rect 2110 1872 2116 1873
rect 2246 1877 2252 1878
rect 2246 1873 2247 1877
rect 2251 1873 2252 1877
rect 2246 1872 2252 1873
rect 2374 1877 2380 1878
rect 2374 1873 2375 1877
rect 2379 1873 2380 1877
rect 2374 1872 2380 1873
rect 2502 1877 2508 1878
rect 2502 1873 2503 1877
rect 2507 1873 2508 1877
rect 2502 1872 2508 1873
rect 2622 1877 2628 1878
rect 2622 1873 2623 1877
rect 2627 1873 2628 1877
rect 2622 1872 2628 1873
rect 2742 1877 2748 1878
rect 2742 1873 2743 1877
rect 2747 1873 2748 1877
rect 2742 1872 2748 1873
rect 2870 1877 2876 1878
rect 2870 1873 2871 1877
rect 2875 1873 2876 1877
rect 2870 1872 2876 1873
rect 2998 1877 3004 1878
rect 2998 1873 2999 1877
rect 3003 1873 3004 1877
rect 2998 1872 3004 1873
rect 142 1849 148 1850
rect 142 1845 143 1849
rect 147 1845 148 1849
rect 142 1844 148 1845
rect 270 1849 276 1850
rect 270 1845 271 1849
rect 275 1845 276 1849
rect 270 1844 276 1845
rect 414 1849 420 1850
rect 414 1845 415 1849
rect 419 1845 420 1849
rect 414 1844 420 1845
rect 558 1849 564 1850
rect 558 1845 559 1849
rect 563 1845 564 1849
rect 558 1844 564 1845
rect 694 1849 700 1850
rect 694 1845 695 1849
rect 699 1845 700 1849
rect 694 1844 700 1845
rect 822 1849 828 1850
rect 822 1845 823 1849
rect 827 1845 828 1849
rect 822 1844 828 1845
rect 942 1849 948 1850
rect 942 1845 943 1849
rect 947 1845 948 1849
rect 942 1844 948 1845
rect 1054 1849 1060 1850
rect 1054 1845 1055 1849
rect 1059 1845 1060 1849
rect 1054 1844 1060 1845
rect 1158 1849 1164 1850
rect 1158 1845 1159 1849
rect 1163 1845 1164 1849
rect 1158 1844 1164 1845
rect 1262 1849 1268 1850
rect 1262 1845 1263 1849
rect 1267 1845 1268 1849
rect 1262 1844 1268 1845
rect 1358 1849 1364 1850
rect 1358 1845 1359 1849
rect 1363 1845 1364 1849
rect 1358 1844 1364 1845
rect 1454 1849 1460 1850
rect 1454 1845 1455 1849
rect 1459 1845 1460 1849
rect 1454 1844 1460 1845
rect 1550 1849 1556 1850
rect 1550 1845 1551 1849
rect 1555 1845 1556 1849
rect 1550 1844 1556 1845
rect 1646 1849 1652 1850
rect 1646 1845 1647 1849
rect 1651 1845 1652 1849
rect 1646 1844 1652 1845
rect 1734 1849 1740 1850
rect 1734 1845 1735 1849
rect 1739 1845 1740 1849
rect 1734 1844 1740 1845
rect 2222 1847 2228 1848
rect 2222 1843 2223 1847
rect 2227 1843 2228 1847
rect 2222 1842 2228 1843
rect 2358 1847 2364 1848
rect 2358 1843 2359 1847
rect 2363 1843 2364 1847
rect 2358 1842 2364 1843
rect 2494 1847 2500 1848
rect 2494 1843 2495 1847
rect 2499 1843 2500 1847
rect 2494 1842 2500 1843
rect 2622 1847 2628 1848
rect 2622 1843 2623 1847
rect 2627 1843 2628 1847
rect 2622 1842 2628 1843
rect 2742 1847 2748 1848
rect 2742 1843 2743 1847
rect 2747 1843 2748 1847
rect 2742 1842 2748 1843
rect 2862 1847 2868 1848
rect 2862 1843 2863 1847
rect 2867 1843 2868 1847
rect 2862 1842 2868 1843
rect 2990 1847 2996 1848
rect 2990 1843 2991 1847
rect 2995 1843 2996 1847
rect 2990 1842 2996 1843
rect 1862 1837 1868 1838
rect 110 1836 116 1837
rect 110 1832 111 1836
rect 115 1832 116 1836
rect 110 1831 116 1832
rect 1822 1836 1828 1837
rect 1822 1832 1823 1836
rect 1827 1832 1828 1836
rect 1862 1833 1863 1837
rect 1867 1833 1868 1837
rect 1862 1832 1868 1833
rect 3574 1837 3580 1838
rect 3574 1833 3575 1837
rect 3579 1833 3580 1837
rect 3574 1832 3580 1833
rect 1822 1831 1828 1832
rect 1862 1820 1868 1821
rect 110 1819 116 1820
rect 110 1815 111 1819
rect 115 1815 116 1819
rect 110 1814 116 1815
rect 1822 1819 1828 1820
rect 1822 1815 1823 1819
rect 1827 1815 1828 1819
rect 1862 1816 1863 1820
rect 1867 1816 1868 1820
rect 1862 1815 1868 1816
rect 3574 1820 3580 1821
rect 3574 1816 3575 1820
rect 3579 1816 3580 1820
rect 3574 1815 3580 1816
rect 1822 1814 1828 1815
rect 134 1809 140 1810
rect 134 1805 135 1809
rect 139 1805 140 1809
rect 134 1804 140 1805
rect 262 1809 268 1810
rect 262 1805 263 1809
rect 267 1805 268 1809
rect 262 1804 268 1805
rect 406 1809 412 1810
rect 406 1805 407 1809
rect 411 1805 412 1809
rect 406 1804 412 1805
rect 550 1809 556 1810
rect 550 1805 551 1809
rect 555 1805 556 1809
rect 550 1804 556 1805
rect 686 1809 692 1810
rect 686 1805 687 1809
rect 691 1805 692 1809
rect 686 1804 692 1805
rect 814 1809 820 1810
rect 814 1805 815 1809
rect 819 1805 820 1809
rect 814 1804 820 1805
rect 934 1809 940 1810
rect 934 1805 935 1809
rect 939 1805 940 1809
rect 934 1804 940 1805
rect 1046 1809 1052 1810
rect 1046 1805 1047 1809
rect 1051 1805 1052 1809
rect 1046 1804 1052 1805
rect 1150 1809 1156 1810
rect 1150 1805 1151 1809
rect 1155 1805 1156 1809
rect 1150 1804 1156 1805
rect 1254 1809 1260 1810
rect 1254 1805 1255 1809
rect 1259 1805 1260 1809
rect 1254 1804 1260 1805
rect 1350 1809 1356 1810
rect 1350 1805 1351 1809
rect 1355 1805 1356 1809
rect 1350 1804 1356 1805
rect 1446 1809 1452 1810
rect 1446 1805 1447 1809
rect 1451 1805 1452 1809
rect 1446 1804 1452 1805
rect 1542 1809 1548 1810
rect 1542 1805 1543 1809
rect 1547 1805 1548 1809
rect 1542 1804 1548 1805
rect 1638 1809 1644 1810
rect 1638 1805 1639 1809
rect 1643 1805 1644 1809
rect 1638 1804 1644 1805
rect 1726 1809 1732 1810
rect 1726 1805 1727 1809
rect 1731 1805 1732 1809
rect 1726 1804 1732 1805
rect 2230 1807 2236 1808
rect 2230 1803 2231 1807
rect 2235 1803 2236 1807
rect 2230 1802 2236 1803
rect 2366 1807 2372 1808
rect 2366 1803 2367 1807
rect 2371 1803 2372 1807
rect 2366 1802 2372 1803
rect 2502 1807 2508 1808
rect 2502 1803 2503 1807
rect 2507 1803 2508 1807
rect 2502 1802 2508 1803
rect 2630 1807 2636 1808
rect 2630 1803 2631 1807
rect 2635 1803 2636 1807
rect 2630 1802 2636 1803
rect 2750 1807 2756 1808
rect 2750 1803 2751 1807
rect 2755 1803 2756 1807
rect 2750 1802 2756 1803
rect 2870 1807 2876 1808
rect 2870 1803 2871 1807
rect 2875 1803 2876 1807
rect 2870 1802 2876 1803
rect 2998 1807 3004 1808
rect 2998 1803 2999 1807
rect 3003 1803 3004 1807
rect 2998 1802 3004 1803
rect 134 1775 140 1776
rect 134 1771 135 1775
rect 139 1771 140 1775
rect 134 1770 140 1771
rect 302 1775 308 1776
rect 302 1771 303 1775
rect 307 1771 308 1775
rect 302 1770 308 1771
rect 494 1775 500 1776
rect 494 1771 495 1775
rect 499 1771 500 1775
rect 494 1770 500 1771
rect 686 1775 692 1776
rect 686 1771 687 1775
rect 691 1771 692 1775
rect 686 1770 692 1771
rect 870 1775 876 1776
rect 870 1771 871 1775
rect 875 1771 876 1775
rect 870 1770 876 1771
rect 1046 1775 1052 1776
rect 1046 1771 1047 1775
rect 1051 1771 1052 1775
rect 1046 1770 1052 1771
rect 1214 1775 1220 1776
rect 1214 1771 1215 1775
rect 1219 1771 1220 1775
rect 1214 1770 1220 1771
rect 1374 1775 1380 1776
rect 1374 1771 1375 1775
rect 1379 1771 1380 1775
rect 1374 1770 1380 1771
rect 1534 1775 1540 1776
rect 1534 1771 1535 1775
rect 1539 1771 1540 1775
rect 1534 1770 1540 1771
rect 1702 1775 1708 1776
rect 1702 1771 1703 1775
rect 1707 1771 1708 1775
rect 1702 1770 1708 1771
rect 2270 1769 2276 1770
rect 110 1765 116 1766
rect 110 1761 111 1765
rect 115 1761 116 1765
rect 110 1760 116 1761
rect 1822 1765 1828 1766
rect 1822 1761 1823 1765
rect 1827 1761 1828 1765
rect 2270 1765 2271 1769
rect 2275 1765 2276 1769
rect 2270 1764 2276 1765
rect 2358 1769 2364 1770
rect 2358 1765 2359 1769
rect 2363 1765 2364 1769
rect 2358 1764 2364 1765
rect 2454 1769 2460 1770
rect 2454 1765 2455 1769
rect 2459 1765 2460 1769
rect 2454 1764 2460 1765
rect 2558 1769 2564 1770
rect 2558 1765 2559 1769
rect 2563 1765 2564 1769
rect 2558 1764 2564 1765
rect 2662 1769 2668 1770
rect 2662 1765 2663 1769
rect 2667 1765 2668 1769
rect 2662 1764 2668 1765
rect 2758 1769 2764 1770
rect 2758 1765 2759 1769
rect 2763 1765 2764 1769
rect 2758 1764 2764 1765
rect 2862 1769 2868 1770
rect 2862 1765 2863 1769
rect 2867 1765 2868 1769
rect 2862 1764 2868 1765
rect 2966 1769 2972 1770
rect 2966 1765 2967 1769
rect 2971 1765 2972 1769
rect 2966 1764 2972 1765
rect 3070 1769 3076 1770
rect 3070 1765 3071 1769
rect 3075 1765 3076 1769
rect 3070 1764 3076 1765
rect 3174 1769 3180 1770
rect 3174 1765 3175 1769
rect 3179 1765 3180 1769
rect 3174 1764 3180 1765
rect 1822 1760 1828 1761
rect 1862 1756 1868 1757
rect 1862 1752 1863 1756
rect 1867 1752 1868 1756
rect 1862 1751 1868 1752
rect 3574 1756 3580 1757
rect 3574 1752 3575 1756
rect 3579 1752 3580 1756
rect 3574 1751 3580 1752
rect 110 1748 116 1749
rect 110 1744 111 1748
rect 115 1744 116 1748
rect 110 1743 116 1744
rect 1822 1748 1828 1749
rect 1822 1744 1823 1748
rect 1827 1744 1828 1748
rect 1822 1743 1828 1744
rect 1862 1739 1868 1740
rect 142 1735 148 1736
rect 142 1731 143 1735
rect 147 1731 148 1735
rect 142 1730 148 1731
rect 310 1735 316 1736
rect 310 1731 311 1735
rect 315 1731 316 1735
rect 310 1730 316 1731
rect 502 1735 508 1736
rect 502 1731 503 1735
rect 507 1731 508 1735
rect 502 1730 508 1731
rect 694 1735 700 1736
rect 694 1731 695 1735
rect 699 1731 700 1735
rect 694 1730 700 1731
rect 878 1735 884 1736
rect 878 1731 879 1735
rect 883 1731 884 1735
rect 878 1730 884 1731
rect 1054 1735 1060 1736
rect 1054 1731 1055 1735
rect 1059 1731 1060 1735
rect 1054 1730 1060 1731
rect 1222 1735 1228 1736
rect 1222 1731 1223 1735
rect 1227 1731 1228 1735
rect 1222 1730 1228 1731
rect 1382 1735 1388 1736
rect 1382 1731 1383 1735
rect 1387 1731 1388 1735
rect 1382 1730 1388 1731
rect 1542 1735 1548 1736
rect 1542 1731 1543 1735
rect 1547 1731 1548 1735
rect 1542 1730 1548 1731
rect 1710 1735 1716 1736
rect 1710 1731 1711 1735
rect 1715 1731 1716 1735
rect 1862 1735 1863 1739
rect 1867 1735 1868 1739
rect 1862 1734 1868 1735
rect 3574 1739 3580 1740
rect 3574 1735 3575 1739
rect 3579 1735 3580 1739
rect 3574 1734 3580 1735
rect 1710 1730 1716 1731
rect 2262 1729 2268 1730
rect 2262 1725 2263 1729
rect 2267 1725 2268 1729
rect 2262 1724 2268 1725
rect 2350 1729 2356 1730
rect 2350 1725 2351 1729
rect 2355 1725 2356 1729
rect 2350 1724 2356 1725
rect 2446 1729 2452 1730
rect 2446 1725 2447 1729
rect 2451 1725 2452 1729
rect 2446 1724 2452 1725
rect 2550 1729 2556 1730
rect 2550 1725 2551 1729
rect 2555 1725 2556 1729
rect 2550 1724 2556 1725
rect 2654 1729 2660 1730
rect 2654 1725 2655 1729
rect 2659 1725 2660 1729
rect 2654 1724 2660 1725
rect 2750 1729 2756 1730
rect 2750 1725 2751 1729
rect 2755 1725 2756 1729
rect 2750 1724 2756 1725
rect 2854 1729 2860 1730
rect 2854 1725 2855 1729
rect 2859 1725 2860 1729
rect 2854 1724 2860 1725
rect 2958 1729 2964 1730
rect 2958 1725 2959 1729
rect 2963 1725 2964 1729
rect 2958 1724 2964 1725
rect 3062 1729 3068 1730
rect 3062 1725 3063 1729
rect 3067 1725 3068 1729
rect 3062 1724 3068 1725
rect 3166 1729 3172 1730
rect 3166 1725 3167 1729
rect 3171 1725 3172 1729
rect 3166 1724 3172 1725
rect 2246 1703 2252 1704
rect 2246 1699 2247 1703
rect 2251 1699 2252 1703
rect 2246 1698 2252 1699
rect 2366 1703 2372 1704
rect 2366 1699 2367 1703
rect 2371 1699 2372 1703
rect 2366 1698 2372 1699
rect 2494 1703 2500 1704
rect 2494 1699 2495 1703
rect 2499 1699 2500 1703
rect 2494 1698 2500 1699
rect 2622 1703 2628 1704
rect 2622 1699 2623 1703
rect 2627 1699 2628 1703
rect 2622 1698 2628 1699
rect 2758 1703 2764 1704
rect 2758 1699 2759 1703
rect 2763 1699 2764 1703
rect 2758 1698 2764 1699
rect 2886 1703 2892 1704
rect 2886 1699 2887 1703
rect 2891 1699 2892 1703
rect 2886 1698 2892 1699
rect 3014 1703 3020 1704
rect 3014 1699 3015 1703
rect 3019 1699 3020 1703
rect 3014 1698 3020 1699
rect 3134 1703 3140 1704
rect 3134 1699 3135 1703
rect 3139 1699 3140 1703
rect 3134 1698 3140 1699
rect 3246 1703 3252 1704
rect 3246 1699 3247 1703
rect 3251 1699 3252 1703
rect 3246 1698 3252 1699
rect 3366 1703 3372 1704
rect 3366 1699 3367 1703
rect 3371 1699 3372 1703
rect 3366 1698 3372 1699
rect 3478 1703 3484 1704
rect 3478 1699 3479 1703
rect 3483 1699 3484 1703
rect 3478 1698 3484 1699
rect 142 1697 148 1698
rect 142 1693 143 1697
rect 147 1693 148 1697
rect 142 1692 148 1693
rect 286 1697 292 1698
rect 286 1693 287 1697
rect 291 1693 292 1697
rect 286 1692 292 1693
rect 470 1697 476 1698
rect 470 1693 471 1697
rect 475 1693 476 1697
rect 470 1692 476 1693
rect 654 1697 660 1698
rect 654 1693 655 1697
rect 659 1693 660 1697
rect 654 1692 660 1693
rect 838 1697 844 1698
rect 838 1693 839 1697
rect 843 1693 844 1697
rect 838 1692 844 1693
rect 1022 1697 1028 1698
rect 1022 1693 1023 1697
rect 1027 1693 1028 1697
rect 1022 1692 1028 1693
rect 1190 1697 1196 1698
rect 1190 1693 1191 1697
rect 1195 1693 1196 1697
rect 1190 1692 1196 1693
rect 1358 1697 1364 1698
rect 1358 1693 1359 1697
rect 1363 1693 1364 1697
rect 1358 1692 1364 1693
rect 1526 1697 1532 1698
rect 1526 1693 1527 1697
rect 1531 1693 1532 1697
rect 1526 1692 1532 1693
rect 1694 1697 1700 1698
rect 1694 1693 1695 1697
rect 1699 1693 1700 1697
rect 1694 1692 1700 1693
rect 1862 1693 1868 1694
rect 1862 1689 1863 1693
rect 1867 1689 1868 1693
rect 1862 1688 1868 1689
rect 3574 1693 3580 1694
rect 3574 1689 3575 1693
rect 3579 1689 3580 1693
rect 3574 1688 3580 1689
rect 110 1684 116 1685
rect 110 1680 111 1684
rect 115 1680 116 1684
rect 110 1679 116 1680
rect 1822 1684 1828 1685
rect 1822 1680 1823 1684
rect 1827 1680 1828 1684
rect 1822 1679 1828 1680
rect 1862 1676 1868 1677
rect 1862 1672 1863 1676
rect 1867 1672 1868 1676
rect 1862 1671 1868 1672
rect 3574 1676 3580 1677
rect 3574 1672 3575 1676
rect 3579 1672 3580 1676
rect 3574 1671 3580 1672
rect 110 1667 116 1668
rect 110 1663 111 1667
rect 115 1663 116 1667
rect 110 1662 116 1663
rect 1822 1667 1828 1668
rect 1822 1663 1823 1667
rect 1827 1663 1828 1667
rect 1822 1662 1828 1663
rect 2254 1663 2260 1664
rect 2254 1659 2255 1663
rect 2259 1659 2260 1663
rect 2254 1658 2260 1659
rect 2374 1663 2380 1664
rect 2374 1659 2375 1663
rect 2379 1659 2380 1663
rect 2374 1658 2380 1659
rect 2502 1663 2508 1664
rect 2502 1659 2503 1663
rect 2507 1659 2508 1663
rect 2502 1658 2508 1659
rect 2630 1663 2636 1664
rect 2630 1659 2631 1663
rect 2635 1659 2636 1663
rect 2630 1658 2636 1659
rect 2766 1663 2772 1664
rect 2766 1659 2767 1663
rect 2771 1659 2772 1663
rect 2766 1658 2772 1659
rect 2894 1663 2900 1664
rect 2894 1659 2895 1663
rect 2899 1659 2900 1663
rect 2894 1658 2900 1659
rect 3022 1663 3028 1664
rect 3022 1659 3023 1663
rect 3027 1659 3028 1663
rect 3022 1658 3028 1659
rect 3142 1663 3148 1664
rect 3142 1659 3143 1663
rect 3147 1659 3148 1663
rect 3142 1658 3148 1659
rect 3254 1663 3260 1664
rect 3254 1659 3255 1663
rect 3259 1659 3260 1663
rect 3254 1658 3260 1659
rect 3374 1663 3380 1664
rect 3374 1659 3375 1663
rect 3379 1659 3380 1663
rect 3374 1658 3380 1659
rect 3486 1663 3492 1664
rect 3486 1659 3487 1663
rect 3491 1659 3492 1663
rect 3486 1658 3492 1659
rect 134 1657 140 1658
rect 134 1653 135 1657
rect 139 1653 140 1657
rect 134 1652 140 1653
rect 278 1657 284 1658
rect 278 1653 279 1657
rect 283 1653 284 1657
rect 278 1652 284 1653
rect 462 1657 468 1658
rect 462 1653 463 1657
rect 467 1653 468 1657
rect 462 1652 468 1653
rect 646 1657 652 1658
rect 646 1653 647 1657
rect 651 1653 652 1657
rect 646 1652 652 1653
rect 830 1657 836 1658
rect 830 1653 831 1657
rect 835 1653 836 1657
rect 830 1652 836 1653
rect 1014 1657 1020 1658
rect 1014 1653 1015 1657
rect 1019 1653 1020 1657
rect 1014 1652 1020 1653
rect 1182 1657 1188 1658
rect 1182 1653 1183 1657
rect 1187 1653 1188 1657
rect 1182 1652 1188 1653
rect 1350 1657 1356 1658
rect 1350 1653 1351 1657
rect 1355 1653 1356 1657
rect 1350 1652 1356 1653
rect 1518 1657 1524 1658
rect 1518 1653 1519 1657
rect 1523 1653 1524 1657
rect 1518 1652 1524 1653
rect 1686 1657 1692 1658
rect 1686 1653 1687 1657
rect 1691 1653 1692 1657
rect 1686 1652 1692 1653
rect 134 1627 140 1628
rect 134 1623 135 1627
rect 139 1623 140 1627
rect 134 1622 140 1623
rect 270 1627 276 1628
rect 270 1623 271 1627
rect 275 1623 276 1627
rect 270 1622 276 1623
rect 446 1627 452 1628
rect 446 1623 447 1627
rect 451 1623 452 1627
rect 446 1622 452 1623
rect 630 1627 636 1628
rect 630 1623 631 1627
rect 635 1623 636 1627
rect 630 1622 636 1623
rect 814 1627 820 1628
rect 814 1623 815 1627
rect 819 1623 820 1627
rect 814 1622 820 1623
rect 990 1627 996 1628
rect 990 1623 991 1627
rect 995 1623 996 1627
rect 990 1622 996 1623
rect 1150 1627 1156 1628
rect 1150 1623 1151 1627
rect 1155 1623 1156 1627
rect 1150 1622 1156 1623
rect 1302 1627 1308 1628
rect 1302 1623 1303 1627
rect 1307 1623 1308 1627
rect 1302 1622 1308 1623
rect 1454 1627 1460 1628
rect 1454 1623 1455 1627
rect 1459 1623 1460 1627
rect 1454 1622 1460 1623
rect 1598 1627 1604 1628
rect 1598 1623 1599 1627
rect 1603 1623 1604 1627
rect 1598 1622 1604 1623
rect 1726 1627 1732 1628
rect 1726 1623 1727 1627
rect 1731 1623 1732 1627
rect 1726 1622 1732 1623
rect 2150 1625 2156 1626
rect 2150 1621 2151 1625
rect 2155 1621 2156 1625
rect 2150 1620 2156 1621
rect 2342 1625 2348 1626
rect 2342 1621 2343 1625
rect 2347 1621 2348 1625
rect 2342 1620 2348 1621
rect 2526 1625 2532 1626
rect 2526 1621 2527 1625
rect 2531 1621 2532 1625
rect 2526 1620 2532 1621
rect 2702 1625 2708 1626
rect 2702 1621 2703 1625
rect 2707 1621 2708 1625
rect 2702 1620 2708 1621
rect 2870 1625 2876 1626
rect 2870 1621 2871 1625
rect 2875 1621 2876 1625
rect 2870 1620 2876 1621
rect 3030 1625 3036 1626
rect 3030 1621 3031 1625
rect 3035 1621 3036 1625
rect 3030 1620 3036 1621
rect 3190 1625 3196 1626
rect 3190 1621 3191 1625
rect 3195 1621 3196 1625
rect 3190 1620 3196 1621
rect 3350 1625 3356 1626
rect 3350 1621 3351 1625
rect 3355 1621 3356 1625
rect 3350 1620 3356 1621
rect 3486 1625 3492 1626
rect 3486 1621 3487 1625
rect 3491 1621 3492 1625
rect 3486 1620 3492 1621
rect 110 1617 116 1618
rect 110 1613 111 1617
rect 115 1613 116 1617
rect 110 1612 116 1613
rect 1822 1617 1828 1618
rect 1822 1613 1823 1617
rect 1827 1613 1828 1617
rect 1822 1612 1828 1613
rect 1862 1612 1868 1613
rect 1862 1608 1863 1612
rect 1867 1608 1868 1612
rect 1862 1607 1868 1608
rect 3574 1612 3580 1613
rect 3574 1608 3575 1612
rect 3579 1608 3580 1612
rect 3574 1607 3580 1608
rect 110 1600 116 1601
rect 110 1596 111 1600
rect 115 1596 116 1600
rect 110 1595 116 1596
rect 1822 1600 1828 1601
rect 1822 1596 1823 1600
rect 1827 1596 1828 1600
rect 1822 1595 1828 1596
rect 1862 1595 1868 1596
rect 1862 1591 1863 1595
rect 1867 1591 1868 1595
rect 1862 1590 1868 1591
rect 3574 1595 3580 1596
rect 3574 1591 3575 1595
rect 3579 1591 3580 1595
rect 3574 1590 3580 1591
rect 142 1587 148 1588
rect 142 1583 143 1587
rect 147 1583 148 1587
rect 142 1582 148 1583
rect 278 1587 284 1588
rect 278 1583 279 1587
rect 283 1583 284 1587
rect 278 1582 284 1583
rect 454 1587 460 1588
rect 454 1583 455 1587
rect 459 1583 460 1587
rect 454 1582 460 1583
rect 638 1587 644 1588
rect 638 1583 639 1587
rect 643 1583 644 1587
rect 638 1582 644 1583
rect 822 1587 828 1588
rect 822 1583 823 1587
rect 827 1583 828 1587
rect 822 1582 828 1583
rect 998 1587 1004 1588
rect 998 1583 999 1587
rect 1003 1583 1004 1587
rect 998 1582 1004 1583
rect 1158 1587 1164 1588
rect 1158 1583 1159 1587
rect 1163 1583 1164 1587
rect 1158 1582 1164 1583
rect 1310 1587 1316 1588
rect 1310 1583 1311 1587
rect 1315 1583 1316 1587
rect 1310 1582 1316 1583
rect 1462 1587 1468 1588
rect 1462 1583 1463 1587
rect 1467 1583 1468 1587
rect 1462 1582 1468 1583
rect 1606 1587 1612 1588
rect 1606 1583 1607 1587
rect 1611 1583 1612 1587
rect 1606 1582 1612 1583
rect 1734 1587 1740 1588
rect 1734 1583 1735 1587
rect 1739 1583 1740 1587
rect 1734 1582 1740 1583
rect 2142 1585 2148 1586
rect 2142 1581 2143 1585
rect 2147 1581 2148 1585
rect 2142 1580 2148 1581
rect 2334 1585 2340 1586
rect 2334 1581 2335 1585
rect 2339 1581 2340 1585
rect 2334 1580 2340 1581
rect 2518 1585 2524 1586
rect 2518 1581 2519 1585
rect 2523 1581 2524 1585
rect 2518 1580 2524 1581
rect 2694 1585 2700 1586
rect 2694 1581 2695 1585
rect 2699 1581 2700 1585
rect 2694 1580 2700 1581
rect 2862 1585 2868 1586
rect 2862 1581 2863 1585
rect 2867 1581 2868 1585
rect 2862 1580 2868 1581
rect 3022 1585 3028 1586
rect 3022 1581 3023 1585
rect 3027 1581 3028 1585
rect 3022 1580 3028 1581
rect 3182 1585 3188 1586
rect 3182 1581 3183 1585
rect 3187 1581 3188 1585
rect 3182 1580 3188 1581
rect 3342 1585 3348 1586
rect 3342 1581 3343 1585
rect 3347 1581 3348 1585
rect 3342 1580 3348 1581
rect 3478 1585 3484 1586
rect 3478 1581 3479 1585
rect 3483 1581 3484 1585
rect 3478 1580 3484 1581
rect 2086 1563 2092 1564
rect 2086 1559 2087 1563
rect 2091 1559 2092 1563
rect 2086 1558 2092 1559
rect 2278 1563 2284 1564
rect 2278 1559 2279 1563
rect 2283 1559 2284 1563
rect 2278 1558 2284 1559
rect 2454 1563 2460 1564
rect 2454 1559 2455 1563
rect 2459 1559 2460 1563
rect 2454 1558 2460 1559
rect 2622 1563 2628 1564
rect 2622 1559 2623 1563
rect 2627 1559 2628 1563
rect 2622 1558 2628 1559
rect 2790 1563 2796 1564
rect 2790 1559 2791 1563
rect 2795 1559 2796 1563
rect 2790 1558 2796 1559
rect 2950 1563 2956 1564
rect 2950 1559 2951 1563
rect 2955 1559 2956 1563
rect 2950 1558 2956 1559
rect 3110 1563 3116 1564
rect 3110 1559 3111 1563
rect 3115 1559 3116 1563
rect 3110 1558 3116 1559
rect 3270 1563 3276 1564
rect 3270 1559 3271 1563
rect 3275 1559 3276 1563
rect 3270 1558 3276 1559
rect 3430 1563 3436 1564
rect 3430 1559 3431 1563
rect 3435 1559 3436 1563
rect 3430 1558 3436 1559
rect 142 1553 148 1554
rect 142 1549 143 1553
rect 147 1549 148 1553
rect 142 1548 148 1549
rect 270 1553 276 1554
rect 270 1549 271 1553
rect 275 1549 276 1553
rect 270 1548 276 1549
rect 430 1553 436 1554
rect 430 1549 431 1553
rect 435 1549 436 1553
rect 430 1548 436 1549
rect 598 1553 604 1554
rect 598 1549 599 1553
rect 603 1549 604 1553
rect 598 1548 604 1549
rect 766 1553 772 1554
rect 766 1549 767 1553
rect 771 1549 772 1553
rect 766 1548 772 1549
rect 934 1553 940 1554
rect 934 1549 935 1553
rect 939 1549 940 1553
rect 934 1548 940 1549
rect 1102 1553 1108 1554
rect 1102 1549 1103 1553
rect 1107 1549 1108 1553
rect 1102 1548 1108 1549
rect 1262 1553 1268 1554
rect 1262 1549 1263 1553
rect 1267 1549 1268 1553
rect 1262 1548 1268 1549
rect 1422 1553 1428 1554
rect 1422 1549 1423 1553
rect 1427 1549 1428 1553
rect 1422 1548 1428 1549
rect 1590 1553 1596 1554
rect 1590 1549 1591 1553
rect 1595 1549 1596 1553
rect 1590 1548 1596 1549
rect 1734 1553 1740 1554
rect 1734 1549 1735 1553
rect 1739 1549 1740 1553
rect 1734 1548 1740 1549
rect 1862 1553 1868 1554
rect 1862 1549 1863 1553
rect 1867 1549 1868 1553
rect 1862 1548 1868 1549
rect 3574 1553 3580 1554
rect 3574 1549 3575 1553
rect 3579 1549 3580 1553
rect 3574 1548 3580 1549
rect 110 1540 116 1541
rect 110 1536 111 1540
rect 115 1536 116 1540
rect 110 1535 116 1536
rect 1822 1540 1828 1541
rect 1822 1536 1823 1540
rect 1827 1536 1828 1540
rect 1822 1535 1828 1536
rect 1862 1536 1868 1537
rect 1862 1532 1863 1536
rect 1867 1532 1868 1536
rect 1862 1531 1868 1532
rect 3574 1536 3580 1537
rect 3574 1532 3575 1536
rect 3579 1532 3580 1536
rect 3574 1531 3580 1532
rect 110 1523 116 1524
rect 110 1519 111 1523
rect 115 1519 116 1523
rect 110 1518 116 1519
rect 1822 1523 1828 1524
rect 1822 1519 1823 1523
rect 1827 1519 1828 1523
rect 1822 1518 1828 1519
rect 2094 1523 2100 1524
rect 2094 1519 2095 1523
rect 2099 1519 2100 1523
rect 2094 1518 2100 1519
rect 2286 1523 2292 1524
rect 2286 1519 2287 1523
rect 2291 1519 2292 1523
rect 2286 1518 2292 1519
rect 2462 1523 2468 1524
rect 2462 1519 2463 1523
rect 2467 1519 2468 1523
rect 2462 1518 2468 1519
rect 2630 1523 2636 1524
rect 2630 1519 2631 1523
rect 2635 1519 2636 1523
rect 2630 1518 2636 1519
rect 2798 1523 2804 1524
rect 2798 1519 2799 1523
rect 2803 1519 2804 1523
rect 2798 1518 2804 1519
rect 2958 1523 2964 1524
rect 2958 1519 2959 1523
rect 2963 1519 2964 1523
rect 2958 1518 2964 1519
rect 3118 1523 3124 1524
rect 3118 1519 3119 1523
rect 3123 1519 3124 1523
rect 3118 1518 3124 1519
rect 3278 1523 3284 1524
rect 3278 1519 3279 1523
rect 3283 1519 3284 1523
rect 3278 1518 3284 1519
rect 3438 1523 3444 1524
rect 3438 1519 3439 1523
rect 3443 1519 3444 1523
rect 3438 1518 3444 1519
rect 134 1513 140 1514
rect 134 1509 135 1513
rect 139 1509 140 1513
rect 134 1508 140 1509
rect 262 1513 268 1514
rect 262 1509 263 1513
rect 267 1509 268 1513
rect 262 1508 268 1509
rect 422 1513 428 1514
rect 422 1509 423 1513
rect 427 1509 428 1513
rect 422 1508 428 1509
rect 590 1513 596 1514
rect 590 1509 591 1513
rect 595 1509 596 1513
rect 590 1508 596 1509
rect 758 1513 764 1514
rect 758 1509 759 1513
rect 763 1509 764 1513
rect 758 1508 764 1509
rect 926 1513 932 1514
rect 926 1509 927 1513
rect 931 1509 932 1513
rect 926 1508 932 1509
rect 1094 1513 1100 1514
rect 1094 1509 1095 1513
rect 1099 1509 1100 1513
rect 1094 1508 1100 1509
rect 1254 1513 1260 1514
rect 1254 1509 1255 1513
rect 1259 1509 1260 1513
rect 1254 1508 1260 1509
rect 1414 1513 1420 1514
rect 1414 1509 1415 1513
rect 1419 1509 1420 1513
rect 1414 1508 1420 1509
rect 1582 1513 1588 1514
rect 1582 1509 1583 1513
rect 1587 1509 1588 1513
rect 1582 1508 1588 1509
rect 1726 1513 1732 1514
rect 1726 1509 1727 1513
rect 1731 1509 1732 1513
rect 1726 1508 1732 1509
rect 182 1487 188 1488
rect 182 1483 183 1487
rect 187 1483 188 1487
rect 182 1482 188 1483
rect 326 1487 332 1488
rect 326 1483 327 1487
rect 331 1483 332 1487
rect 326 1482 332 1483
rect 470 1487 476 1488
rect 470 1483 471 1487
rect 475 1483 476 1487
rect 470 1482 476 1483
rect 606 1487 612 1488
rect 606 1483 607 1487
rect 611 1483 612 1487
rect 606 1482 612 1483
rect 742 1487 748 1488
rect 742 1483 743 1487
rect 747 1483 748 1487
rect 742 1482 748 1483
rect 870 1487 876 1488
rect 870 1483 871 1487
rect 875 1483 876 1487
rect 870 1482 876 1483
rect 990 1487 996 1488
rect 990 1483 991 1487
rect 995 1483 996 1487
rect 990 1482 996 1483
rect 1118 1487 1124 1488
rect 1118 1483 1119 1487
rect 1123 1483 1124 1487
rect 1118 1482 1124 1483
rect 1246 1487 1252 1488
rect 1246 1483 1247 1487
rect 1251 1483 1252 1487
rect 1246 1482 1252 1483
rect 1374 1487 1380 1488
rect 1374 1483 1375 1487
rect 1379 1483 1380 1487
rect 1374 1482 1380 1483
rect 1894 1481 1900 1482
rect 110 1477 116 1478
rect 110 1473 111 1477
rect 115 1473 116 1477
rect 110 1472 116 1473
rect 1822 1477 1828 1478
rect 1822 1473 1823 1477
rect 1827 1473 1828 1477
rect 1894 1477 1895 1481
rect 1899 1477 1900 1481
rect 1894 1476 1900 1477
rect 1990 1481 1996 1482
rect 1990 1477 1991 1481
rect 1995 1477 1996 1481
rect 1990 1476 1996 1477
rect 2118 1481 2124 1482
rect 2118 1477 2119 1481
rect 2123 1477 2124 1481
rect 2118 1476 2124 1477
rect 2246 1481 2252 1482
rect 2246 1477 2247 1481
rect 2251 1477 2252 1481
rect 2246 1476 2252 1477
rect 2382 1481 2388 1482
rect 2382 1477 2383 1481
rect 2387 1477 2388 1481
rect 2382 1476 2388 1477
rect 2534 1481 2540 1482
rect 2534 1477 2535 1481
rect 2539 1477 2540 1481
rect 2534 1476 2540 1477
rect 2702 1481 2708 1482
rect 2702 1477 2703 1481
rect 2707 1477 2708 1481
rect 2702 1476 2708 1477
rect 2886 1481 2892 1482
rect 2886 1477 2887 1481
rect 2891 1477 2892 1481
rect 2886 1476 2892 1477
rect 3086 1481 3092 1482
rect 3086 1477 3087 1481
rect 3091 1477 3092 1481
rect 3086 1476 3092 1477
rect 3294 1481 3300 1482
rect 3294 1477 3295 1481
rect 3299 1477 3300 1481
rect 3294 1476 3300 1477
rect 3486 1481 3492 1482
rect 3486 1477 3487 1481
rect 3491 1477 3492 1481
rect 3486 1476 3492 1477
rect 1822 1472 1828 1473
rect 1862 1468 1868 1469
rect 1862 1464 1863 1468
rect 1867 1464 1868 1468
rect 1862 1463 1868 1464
rect 3574 1468 3580 1469
rect 3574 1464 3575 1468
rect 3579 1464 3580 1468
rect 3574 1463 3580 1464
rect 110 1460 116 1461
rect 110 1456 111 1460
rect 115 1456 116 1460
rect 110 1455 116 1456
rect 1822 1460 1828 1461
rect 1822 1456 1823 1460
rect 1827 1456 1828 1460
rect 1822 1455 1828 1456
rect 1862 1451 1868 1452
rect 190 1447 196 1448
rect 190 1443 191 1447
rect 195 1443 196 1447
rect 190 1442 196 1443
rect 334 1447 340 1448
rect 334 1443 335 1447
rect 339 1443 340 1447
rect 334 1442 340 1443
rect 478 1447 484 1448
rect 478 1443 479 1447
rect 483 1443 484 1447
rect 478 1442 484 1443
rect 614 1447 620 1448
rect 614 1443 615 1447
rect 619 1443 620 1447
rect 614 1442 620 1443
rect 750 1447 756 1448
rect 750 1443 751 1447
rect 755 1443 756 1447
rect 750 1442 756 1443
rect 878 1447 884 1448
rect 878 1443 879 1447
rect 883 1443 884 1447
rect 878 1442 884 1443
rect 998 1447 1004 1448
rect 998 1443 999 1447
rect 1003 1443 1004 1447
rect 998 1442 1004 1443
rect 1126 1447 1132 1448
rect 1126 1443 1127 1447
rect 1131 1443 1132 1447
rect 1126 1442 1132 1443
rect 1254 1447 1260 1448
rect 1254 1443 1255 1447
rect 1259 1443 1260 1447
rect 1254 1442 1260 1443
rect 1382 1447 1388 1448
rect 1382 1443 1383 1447
rect 1387 1443 1388 1447
rect 1862 1447 1863 1451
rect 1867 1447 1868 1451
rect 1862 1446 1868 1447
rect 3574 1451 3580 1452
rect 3574 1447 3575 1451
rect 3579 1447 3580 1451
rect 3574 1446 3580 1447
rect 1382 1442 1388 1443
rect 1886 1441 1892 1442
rect 1886 1437 1887 1441
rect 1891 1437 1892 1441
rect 1886 1436 1892 1437
rect 1982 1441 1988 1442
rect 1982 1437 1983 1441
rect 1987 1437 1988 1441
rect 1982 1436 1988 1437
rect 2110 1441 2116 1442
rect 2110 1437 2111 1441
rect 2115 1437 2116 1441
rect 2110 1436 2116 1437
rect 2238 1441 2244 1442
rect 2238 1437 2239 1441
rect 2243 1437 2244 1441
rect 2238 1436 2244 1437
rect 2374 1441 2380 1442
rect 2374 1437 2375 1441
rect 2379 1437 2380 1441
rect 2374 1436 2380 1437
rect 2526 1441 2532 1442
rect 2526 1437 2527 1441
rect 2531 1437 2532 1441
rect 2526 1436 2532 1437
rect 2694 1441 2700 1442
rect 2694 1437 2695 1441
rect 2699 1437 2700 1441
rect 2694 1436 2700 1437
rect 2878 1441 2884 1442
rect 2878 1437 2879 1441
rect 2883 1437 2884 1441
rect 2878 1436 2884 1437
rect 3078 1441 3084 1442
rect 3078 1437 3079 1441
rect 3083 1437 3084 1441
rect 3078 1436 3084 1437
rect 3286 1441 3292 1442
rect 3286 1437 3287 1441
rect 3291 1437 3292 1441
rect 3286 1436 3292 1437
rect 3478 1441 3484 1442
rect 3478 1437 3479 1441
rect 3483 1437 3484 1441
rect 3478 1436 3484 1437
rect 1886 1415 1892 1416
rect 1886 1411 1887 1415
rect 1891 1411 1892 1415
rect 1886 1410 1892 1411
rect 1974 1415 1980 1416
rect 1974 1411 1975 1415
rect 1979 1411 1980 1415
rect 1974 1410 1980 1411
rect 2070 1415 2076 1416
rect 2070 1411 2071 1415
rect 2075 1411 2076 1415
rect 2070 1410 2076 1411
rect 2182 1415 2188 1416
rect 2182 1411 2183 1415
rect 2187 1411 2188 1415
rect 2182 1410 2188 1411
rect 2302 1415 2308 1416
rect 2302 1411 2303 1415
rect 2307 1411 2308 1415
rect 2302 1410 2308 1411
rect 2438 1415 2444 1416
rect 2438 1411 2439 1415
rect 2443 1411 2444 1415
rect 2438 1410 2444 1411
rect 2606 1415 2612 1416
rect 2606 1411 2607 1415
rect 2611 1411 2612 1415
rect 2606 1410 2612 1411
rect 2806 1415 2812 1416
rect 2806 1411 2807 1415
rect 2811 1411 2812 1415
rect 2806 1410 2812 1411
rect 3030 1415 3036 1416
rect 3030 1411 3031 1415
rect 3035 1411 3036 1415
rect 3030 1410 3036 1411
rect 3262 1415 3268 1416
rect 3262 1411 3263 1415
rect 3267 1411 3268 1415
rect 3262 1410 3268 1411
rect 3478 1415 3484 1416
rect 3478 1411 3479 1415
rect 3483 1411 3484 1415
rect 3478 1410 3484 1411
rect 198 1405 204 1406
rect 198 1401 199 1405
rect 203 1401 204 1405
rect 198 1400 204 1401
rect 334 1405 340 1406
rect 334 1401 335 1405
rect 339 1401 340 1405
rect 334 1400 340 1401
rect 462 1405 468 1406
rect 462 1401 463 1405
rect 467 1401 468 1405
rect 462 1400 468 1401
rect 582 1405 588 1406
rect 582 1401 583 1405
rect 587 1401 588 1405
rect 582 1400 588 1401
rect 702 1405 708 1406
rect 702 1401 703 1405
rect 707 1401 708 1405
rect 702 1400 708 1401
rect 814 1405 820 1406
rect 814 1401 815 1405
rect 819 1401 820 1405
rect 814 1400 820 1401
rect 918 1405 924 1406
rect 918 1401 919 1405
rect 923 1401 924 1405
rect 918 1400 924 1401
rect 1014 1405 1020 1406
rect 1014 1401 1015 1405
rect 1019 1401 1020 1405
rect 1014 1400 1020 1401
rect 1118 1405 1124 1406
rect 1118 1401 1119 1405
rect 1123 1401 1124 1405
rect 1118 1400 1124 1401
rect 1222 1405 1228 1406
rect 1222 1401 1223 1405
rect 1227 1401 1228 1405
rect 1222 1400 1228 1401
rect 1326 1405 1332 1406
rect 1326 1401 1327 1405
rect 1331 1401 1332 1405
rect 1326 1400 1332 1401
rect 1862 1405 1868 1406
rect 1862 1401 1863 1405
rect 1867 1401 1868 1405
rect 1862 1400 1868 1401
rect 3574 1405 3580 1406
rect 3574 1401 3575 1405
rect 3579 1401 3580 1405
rect 3574 1400 3580 1401
rect 110 1392 116 1393
rect 110 1388 111 1392
rect 115 1388 116 1392
rect 110 1387 116 1388
rect 1822 1392 1828 1393
rect 1822 1388 1823 1392
rect 1827 1388 1828 1392
rect 1822 1387 1828 1388
rect 1862 1388 1868 1389
rect 1862 1384 1863 1388
rect 1867 1384 1868 1388
rect 1862 1383 1868 1384
rect 3574 1388 3580 1389
rect 3574 1384 3575 1388
rect 3579 1384 3580 1388
rect 3574 1383 3580 1384
rect 110 1375 116 1376
rect 110 1371 111 1375
rect 115 1371 116 1375
rect 110 1370 116 1371
rect 1822 1375 1828 1376
rect 1822 1371 1823 1375
rect 1827 1371 1828 1375
rect 1822 1370 1828 1371
rect 1894 1375 1900 1376
rect 1894 1371 1895 1375
rect 1899 1371 1900 1375
rect 1894 1370 1900 1371
rect 1982 1375 1988 1376
rect 1982 1371 1983 1375
rect 1987 1371 1988 1375
rect 1982 1370 1988 1371
rect 2078 1375 2084 1376
rect 2078 1371 2079 1375
rect 2083 1371 2084 1375
rect 2078 1370 2084 1371
rect 2190 1375 2196 1376
rect 2190 1371 2191 1375
rect 2195 1371 2196 1375
rect 2190 1370 2196 1371
rect 2310 1375 2316 1376
rect 2310 1371 2311 1375
rect 2315 1371 2316 1375
rect 2310 1370 2316 1371
rect 2446 1375 2452 1376
rect 2446 1371 2447 1375
rect 2451 1371 2452 1375
rect 2446 1370 2452 1371
rect 2614 1375 2620 1376
rect 2614 1371 2615 1375
rect 2619 1371 2620 1375
rect 2614 1370 2620 1371
rect 2814 1375 2820 1376
rect 2814 1371 2815 1375
rect 2819 1371 2820 1375
rect 2814 1370 2820 1371
rect 3038 1375 3044 1376
rect 3038 1371 3039 1375
rect 3043 1371 3044 1375
rect 3038 1370 3044 1371
rect 3270 1375 3276 1376
rect 3270 1371 3271 1375
rect 3275 1371 3276 1375
rect 3270 1370 3276 1371
rect 3486 1375 3492 1376
rect 3486 1371 3487 1375
rect 3491 1371 3492 1375
rect 3486 1370 3492 1371
rect 190 1365 196 1366
rect 190 1361 191 1365
rect 195 1361 196 1365
rect 190 1360 196 1361
rect 326 1365 332 1366
rect 326 1361 327 1365
rect 331 1361 332 1365
rect 326 1360 332 1361
rect 454 1365 460 1366
rect 454 1361 455 1365
rect 459 1361 460 1365
rect 454 1360 460 1361
rect 574 1365 580 1366
rect 574 1361 575 1365
rect 579 1361 580 1365
rect 574 1360 580 1361
rect 694 1365 700 1366
rect 694 1361 695 1365
rect 699 1361 700 1365
rect 694 1360 700 1361
rect 806 1365 812 1366
rect 806 1361 807 1365
rect 811 1361 812 1365
rect 806 1360 812 1361
rect 910 1365 916 1366
rect 910 1361 911 1365
rect 915 1361 916 1365
rect 910 1360 916 1361
rect 1006 1365 1012 1366
rect 1006 1361 1007 1365
rect 1011 1361 1012 1365
rect 1006 1360 1012 1361
rect 1110 1365 1116 1366
rect 1110 1361 1111 1365
rect 1115 1361 1116 1365
rect 1110 1360 1116 1361
rect 1214 1365 1220 1366
rect 1214 1361 1215 1365
rect 1219 1361 1220 1365
rect 1214 1360 1220 1361
rect 1318 1365 1324 1366
rect 1318 1361 1319 1365
rect 1323 1361 1324 1365
rect 1318 1360 1324 1361
rect 230 1339 236 1340
rect 230 1335 231 1339
rect 235 1335 236 1339
rect 230 1334 236 1335
rect 382 1339 388 1340
rect 382 1335 383 1339
rect 387 1335 388 1339
rect 382 1334 388 1335
rect 542 1339 548 1340
rect 542 1335 543 1339
rect 547 1335 548 1339
rect 542 1334 548 1335
rect 702 1339 708 1340
rect 702 1335 703 1339
rect 707 1335 708 1339
rect 702 1334 708 1335
rect 870 1339 876 1340
rect 870 1335 871 1339
rect 875 1335 876 1339
rect 870 1334 876 1335
rect 1038 1339 1044 1340
rect 1038 1335 1039 1339
rect 1043 1335 1044 1339
rect 1038 1334 1044 1335
rect 1206 1339 1212 1340
rect 1206 1335 1207 1339
rect 1211 1335 1212 1339
rect 1206 1334 1212 1335
rect 1374 1339 1380 1340
rect 1374 1335 1375 1339
rect 1379 1335 1380 1339
rect 1374 1334 1380 1335
rect 1894 1337 1900 1338
rect 1894 1333 1895 1337
rect 1899 1333 1900 1337
rect 1894 1332 1900 1333
rect 1982 1337 1988 1338
rect 1982 1333 1983 1337
rect 1987 1333 1988 1337
rect 1982 1332 1988 1333
rect 2102 1337 2108 1338
rect 2102 1333 2103 1337
rect 2107 1333 2108 1337
rect 2102 1332 2108 1333
rect 2222 1337 2228 1338
rect 2222 1333 2223 1337
rect 2227 1333 2228 1337
rect 2222 1332 2228 1333
rect 2358 1337 2364 1338
rect 2358 1333 2359 1337
rect 2363 1333 2364 1337
rect 2358 1332 2364 1333
rect 2510 1337 2516 1338
rect 2510 1333 2511 1337
rect 2515 1333 2516 1337
rect 2510 1332 2516 1333
rect 2686 1337 2692 1338
rect 2686 1333 2687 1337
rect 2691 1333 2692 1337
rect 2686 1332 2692 1333
rect 2870 1337 2876 1338
rect 2870 1333 2871 1337
rect 2875 1333 2876 1337
rect 2870 1332 2876 1333
rect 3070 1337 3076 1338
rect 3070 1333 3071 1337
rect 3075 1333 3076 1337
rect 3070 1332 3076 1333
rect 3278 1337 3284 1338
rect 3278 1333 3279 1337
rect 3283 1333 3284 1337
rect 3278 1332 3284 1333
rect 3486 1337 3492 1338
rect 3486 1333 3487 1337
rect 3491 1333 3492 1337
rect 3486 1332 3492 1333
rect 110 1329 116 1330
rect 110 1325 111 1329
rect 115 1325 116 1329
rect 110 1324 116 1325
rect 1822 1329 1828 1330
rect 1822 1325 1823 1329
rect 1827 1325 1828 1329
rect 1822 1324 1828 1325
rect 1862 1324 1868 1325
rect 1862 1320 1863 1324
rect 1867 1320 1868 1324
rect 1862 1319 1868 1320
rect 3574 1324 3580 1325
rect 3574 1320 3575 1324
rect 3579 1320 3580 1324
rect 3574 1319 3580 1320
rect 110 1312 116 1313
rect 110 1308 111 1312
rect 115 1308 116 1312
rect 110 1307 116 1308
rect 1822 1312 1828 1313
rect 1822 1308 1823 1312
rect 1827 1308 1828 1312
rect 1822 1307 1828 1308
rect 1862 1307 1868 1308
rect 1862 1303 1863 1307
rect 1867 1303 1868 1307
rect 1862 1302 1868 1303
rect 3574 1307 3580 1308
rect 3574 1303 3575 1307
rect 3579 1303 3580 1307
rect 3574 1302 3580 1303
rect 238 1299 244 1300
rect 238 1295 239 1299
rect 243 1295 244 1299
rect 238 1294 244 1295
rect 390 1299 396 1300
rect 390 1295 391 1299
rect 395 1295 396 1299
rect 390 1294 396 1295
rect 550 1299 556 1300
rect 550 1295 551 1299
rect 555 1295 556 1299
rect 550 1294 556 1295
rect 710 1299 716 1300
rect 710 1295 711 1299
rect 715 1295 716 1299
rect 710 1294 716 1295
rect 878 1299 884 1300
rect 878 1295 879 1299
rect 883 1295 884 1299
rect 878 1294 884 1295
rect 1046 1299 1052 1300
rect 1046 1295 1047 1299
rect 1051 1295 1052 1299
rect 1046 1294 1052 1295
rect 1214 1299 1220 1300
rect 1214 1295 1215 1299
rect 1219 1295 1220 1299
rect 1214 1294 1220 1295
rect 1382 1299 1388 1300
rect 1382 1295 1383 1299
rect 1387 1295 1388 1299
rect 1382 1294 1388 1295
rect 1886 1297 1892 1298
rect 1886 1293 1887 1297
rect 1891 1293 1892 1297
rect 1886 1292 1892 1293
rect 1974 1297 1980 1298
rect 1974 1293 1975 1297
rect 1979 1293 1980 1297
rect 1974 1292 1980 1293
rect 2094 1297 2100 1298
rect 2094 1293 2095 1297
rect 2099 1293 2100 1297
rect 2094 1292 2100 1293
rect 2214 1297 2220 1298
rect 2214 1293 2215 1297
rect 2219 1293 2220 1297
rect 2214 1292 2220 1293
rect 2350 1297 2356 1298
rect 2350 1293 2351 1297
rect 2355 1293 2356 1297
rect 2350 1292 2356 1293
rect 2502 1297 2508 1298
rect 2502 1293 2503 1297
rect 2507 1293 2508 1297
rect 2502 1292 2508 1293
rect 2678 1297 2684 1298
rect 2678 1293 2679 1297
rect 2683 1293 2684 1297
rect 2678 1292 2684 1293
rect 2862 1297 2868 1298
rect 2862 1293 2863 1297
rect 2867 1293 2868 1297
rect 2862 1292 2868 1293
rect 3062 1297 3068 1298
rect 3062 1293 3063 1297
rect 3067 1293 3068 1297
rect 3062 1292 3068 1293
rect 3270 1297 3276 1298
rect 3270 1293 3271 1297
rect 3275 1293 3276 1297
rect 3270 1292 3276 1293
rect 3478 1297 3484 1298
rect 3478 1293 3479 1297
rect 3483 1293 3484 1297
rect 3478 1292 3484 1293
rect 214 1265 220 1266
rect 214 1261 215 1265
rect 219 1261 220 1265
rect 214 1260 220 1261
rect 358 1265 364 1266
rect 358 1261 359 1265
rect 363 1261 364 1265
rect 358 1260 364 1261
rect 518 1265 524 1266
rect 518 1261 519 1265
rect 523 1261 524 1265
rect 518 1260 524 1261
rect 678 1265 684 1266
rect 678 1261 679 1265
rect 683 1261 684 1265
rect 678 1260 684 1261
rect 838 1265 844 1266
rect 838 1261 839 1265
rect 843 1261 844 1265
rect 838 1260 844 1261
rect 998 1265 1004 1266
rect 998 1261 999 1265
rect 1003 1261 1004 1265
rect 998 1260 1004 1261
rect 1150 1265 1156 1266
rect 1150 1261 1151 1265
rect 1155 1261 1156 1265
rect 1150 1260 1156 1261
rect 1294 1265 1300 1266
rect 1294 1261 1295 1265
rect 1299 1261 1300 1265
rect 1294 1260 1300 1261
rect 1438 1265 1444 1266
rect 1438 1261 1439 1265
rect 1443 1261 1444 1265
rect 1438 1260 1444 1261
rect 1590 1265 1596 1266
rect 1590 1261 1591 1265
rect 1595 1261 1596 1265
rect 1590 1260 1596 1261
rect 2054 1263 2060 1264
rect 2054 1259 2055 1263
rect 2059 1259 2060 1263
rect 2054 1258 2060 1259
rect 2142 1263 2148 1264
rect 2142 1259 2143 1263
rect 2147 1259 2148 1263
rect 2142 1258 2148 1259
rect 2238 1263 2244 1264
rect 2238 1259 2239 1263
rect 2243 1259 2244 1263
rect 2238 1258 2244 1259
rect 2334 1263 2340 1264
rect 2334 1259 2335 1263
rect 2339 1259 2340 1263
rect 2334 1258 2340 1259
rect 2430 1263 2436 1264
rect 2430 1259 2431 1263
rect 2435 1259 2436 1263
rect 2430 1258 2436 1259
rect 2550 1263 2556 1264
rect 2550 1259 2551 1263
rect 2555 1259 2556 1263
rect 2550 1258 2556 1259
rect 2686 1263 2692 1264
rect 2686 1259 2687 1263
rect 2691 1259 2692 1263
rect 2686 1258 2692 1259
rect 2854 1263 2860 1264
rect 2854 1259 2855 1263
rect 2859 1259 2860 1263
rect 2854 1258 2860 1259
rect 3038 1263 3044 1264
rect 3038 1259 3039 1263
rect 3043 1259 3044 1263
rect 3038 1258 3044 1259
rect 3230 1263 3236 1264
rect 3230 1259 3231 1263
rect 3235 1259 3236 1263
rect 3230 1258 3236 1259
rect 3430 1263 3436 1264
rect 3430 1259 3431 1263
rect 3435 1259 3436 1263
rect 3430 1258 3436 1259
rect 1862 1253 1868 1254
rect 110 1252 116 1253
rect 110 1248 111 1252
rect 115 1248 116 1252
rect 110 1247 116 1248
rect 1822 1252 1828 1253
rect 1822 1248 1823 1252
rect 1827 1248 1828 1252
rect 1862 1249 1863 1253
rect 1867 1249 1868 1253
rect 1862 1248 1868 1249
rect 3574 1253 3580 1254
rect 3574 1249 3575 1253
rect 3579 1249 3580 1253
rect 3574 1248 3580 1249
rect 1822 1247 1828 1248
rect 1862 1236 1868 1237
rect 110 1235 116 1236
rect 110 1231 111 1235
rect 115 1231 116 1235
rect 110 1230 116 1231
rect 1822 1235 1828 1236
rect 1822 1231 1823 1235
rect 1827 1231 1828 1235
rect 1862 1232 1863 1236
rect 1867 1232 1868 1236
rect 1862 1231 1868 1232
rect 3574 1236 3580 1237
rect 3574 1232 3575 1236
rect 3579 1232 3580 1236
rect 3574 1231 3580 1232
rect 1822 1230 1828 1231
rect 206 1225 212 1226
rect 206 1221 207 1225
rect 211 1221 212 1225
rect 206 1220 212 1221
rect 350 1225 356 1226
rect 350 1221 351 1225
rect 355 1221 356 1225
rect 350 1220 356 1221
rect 510 1225 516 1226
rect 510 1221 511 1225
rect 515 1221 516 1225
rect 510 1220 516 1221
rect 670 1225 676 1226
rect 670 1221 671 1225
rect 675 1221 676 1225
rect 670 1220 676 1221
rect 830 1225 836 1226
rect 830 1221 831 1225
rect 835 1221 836 1225
rect 830 1220 836 1221
rect 990 1225 996 1226
rect 990 1221 991 1225
rect 995 1221 996 1225
rect 990 1220 996 1221
rect 1142 1225 1148 1226
rect 1142 1221 1143 1225
rect 1147 1221 1148 1225
rect 1142 1220 1148 1221
rect 1286 1225 1292 1226
rect 1286 1221 1287 1225
rect 1291 1221 1292 1225
rect 1286 1220 1292 1221
rect 1430 1225 1436 1226
rect 1430 1221 1431 1225
rect 1435 1221 1436 1225
rect 1430 1220 1436 1221
rect 1582 1225 1588 1226
rect 1582 1221 1583 1225
rect 1587 1221 1588 1225
rect 1582 1220 1588 1221
rect 2062 1223 2068 1224
rect 2062 1219 2063 1223
rect 2067 1219 2068 1223
rect 2062 1218 2068 1219
rect 2150 1223 2156 1224
rect 2150 1219 2151 1223
rect 2155 1219 2156 1223
rect 2150 1218 2156 1219
rect 2246 1223 2252 1224
rect 2246 1219 2247 1223
rect 2251 1219 2252 1223
rect 2246 1218 2252 1219
rect 2342 1223 2348 1224
rect 2342 1219 2343 1223
rect 2347 1219 2348 1223
rect 2342 1218 2348 1219
rect 2438 1223 2444 1224
rect 2438 1219 2439 1223
rect 2443 1219 2444 1223
rect 2438 1218 2444 1219
rect 2558 1223 2564 1224
rect 2558 1219 2559 1223
rect 2563 1219 2564 1223
rect 2558 1218 2564 1219
rect 2694 1223 2700 1224
rect 2694 1219 2695 1223
rect 2699 1219 2700 1223
rect 2694 1218 2700 1219
rect 2862 1223 2868 1224
rect 2862 1219 2863 1223
rect 2867 1219 2868 1223
rect 2862 1218 2868 1219
rect 3046 1223 3052 1224
rect 3046 1219 3047 1223
rect 3051 1219 3052 1223
rect 3046 1218 3052 1219
rect 3238 1223 3244 1224
rect 3238 1219 3239 1223
rect 3243 1219 3244 1223
rect 3238 1218 3244 1219
rect 3438 1223 3444 1224
rect 3438 1219 3439 1223
rect 3443 1219 3444 1223
rect 3438 1218 3444 1219
rect 134 1195 140 1196
rect 134 1191 135 1195
rect 139 1191 140 1195
rect 134 1190 140 1191
rect 270 1195 276 1196
rect 270 1191 271 1195
rect 275 1191 276 1195
rect 270 1190 276 1191
rect 422 1195 428 1196
rect 422 1191 423 1195
rect 427 1191 428 1195
rect 422 1190 428 1191
rect 574 1195 580 1196
rect 574 1191 575 1195
rect 579 1191 580 1195
rect 574 1190 580 1191
rect 726 1195 732 1196
rect 726 1191 727 1195
rect 731 1191 732 1195
rect 726 1190 732 1191
rect 886 1195 892 1196
rect 886 1191 887 1195
rect 891 1191 892 1195
rect 886 1190 892 1191
rect 1054 1195 1060 1196
rect 1054 1191 1055 1195
rect 1059 1191 1060 1195
rect 1054 1190 1060 1191
rect 1230 1195 1236 1196
rect 1230 1191 1231 1195
rect 1235 1191 1236 1195
rect 1230 1190 1236 1191
rect 1414 1195 1420 1196
rect 1414 1191 1415 1195
rect 1419 1191 1420 1195
rect 1414 1190 1420 1191
rect 1598 1195 1604 1196
rect 1598 1191 1599 1195
rect 1603 1191 1604 1195
rect 1598 1190 1604 1191
rect 110 1185 116 1186
rect 110 1181 111 1185
rect 115 1181 116 1185
rect 110 1180 116 1181
rect 1822 1185 1828 1186
rect 1822 1181 1823 1185
rect 1827 1181 1828 1185
rect 1822 1180 1828 1181
rect 2038 1185 2044 1186
rect 2038 1181 2039 1185
rect 2043 1181 2044 1185
rect 2038 1180 2044 1181
rect 2150 1185 2156 1186
rect 2150 1181 2151 1185
rect 2155 1181 2156 1185
rect 2150 1180 2156 1181
rect 2278 1185 2284 1186
rect 2278 1181 2279 1185
rect 2283 1181 2284 1185
rect 2278 1180 2284 1181
rect 2414 1185 2420 1186
rect 2414 1181 2415 1185
rect 2419 1181 2420 1185
rect 2414 1180 2420 1181
rect 2558 1185 2564 1186
rect 2558 1181 2559 1185
rect 2563 1181 2564 1185
rect 2558 1180 2564 1181
rect 2710 1185 2716 1186
rect 2710 1181 2711 1185
rect 2715 1181 2716 1185
rect 2710 1180 2716 1181
rect 2862 1185 2868 1186
rect 2862 1181 2863 1185
rect 2867 1181 2868 1185
rect 2862 1180 2868 1181
rect 3014 1185 3020 1186
rect 3014 1181 3015 1185
rect 3019 1181 3020 1185
rect 3014 1180 3020 1181
rect 3166 1185 3172 1186
rect 3166 1181 3167 1185
rect 3171 1181 3172 1185
rect 3166 1180 3172 1181
rect 3326 1185 3332 1186
rect 3326 1181 3327 1185
rect 3331 1181 3332 1185
rect 3326 1180 3332 1181
rect 3486 1185 3492 1186
rect 3486 1181 3487 1185
rect 3491 1181 3492 1185
rect 3486 1180 3492 1181
rect 1862 1172 1868 1173
rect 110 1168 116 1169
rect 110 1164 111 1168
rect 115 1164 116 1168
rect 110 1163 116 1164
rect 1822 1168 1828 1169
rect 1822 1164 1823 1168
rect 1827 1164 1828 1168
rect 1862 1168 1863 1172
rect 1867 1168 1868 1172
rect 1862 1167 1868 1168
rect 3574 1172 3580 1173
rect 3574 1168 3575 1172
rect 3579 1168 3580 1172
rect 3574 1167 3580 1168
rect 1822 1163 1828 1164
rect 142 1155 148 1156
rect 142 1151 143 1155
rect 147 1151 148 1155
rect 142 1150 148 1151
rect 278 1155 284 1156
rect 278 1151 279 1155
rect 283 1151 284 1155
rect 278 1150 284 1151
rect 430 1155 436 1156
rect 430 1151 431 1155
rect 435 1151 436 1155
rect 430 1150 436 1151
rect 582 1155 588 1156
rect 582 1151 583 1155
rect 587 1151 588 1155
rect 582 1150 588 1151
rect 734 1155 740 1156
rect 734 1151 735 1155
rect 739 1151 740 1155
rect 734 1150 740 1151
rect 894 1155 900 1156
rect 894 1151 895 1155
rect 899 1151 900 1155
rect 894 1150 900 1151
rect 1062 1155 1068 1156
rect 1062 1151 1063 1155
rect 1067 1151 1068 1155
rect 1062 1150 1068 1151
rect 1238 1155 1244 1156
rect 1238 1151 1239 1155
rect 1243 1151 1244 1155
rect 1238 1150 1244 1151
rect 1422 1155 1428 1156
rect 1422 1151 1423 1155
rect 1427 1151 1428 1155
rect 1422 1150 1428 1151
rect 1606 1155 1612 1156
rect 1606 1151 1607 1155
rect 1611 1151 1612 1155
rect 1606 1150 1612 1151
rect 1862 1155 1868 1156
rect 1862 1151 1863 1155
rect 1867 1151 1868 1155
rect 1862 1150 1868 1151
rect 3574 1155 3580 1156
rect 3574 1151 3575 1155
rect 3579 1151 3580 1155
rect 3574 1150 3580 1151
rect 2030 1145 2036 1146
rect 2030 1141 2031 1145
rect 2035 1141 2036 1145
rect 2030 1140 2036 1141
rect 2142 1145 2148 1146
rect 2142 1141 2143 1145
rect 2147 1141 2148 1145
rect 2142 1140 2148 1141
rect 2270 1145 2276 1146
rect 2270 1141 2271 1145
rect 2275 1141 2276 1145
rect 2270 1140 2276 1141
rect 2406 1145 2412 1146
rect 2406 1141 2407 1145
rect 2411 1141 2412 1145
rect 2406 1140 2412 1141
rect 2550 1145 2556 1146
rect 2550 1141 2551 1145
rect 2555 1141 2556 1145
rect 2550 1140 2556 1141
rect 2702 1145 2708 1146
rect 2702 1141 2703 1145
rect 2707 1141 2708 1145
rect 2702 1140 2708 1141
rect 2854 1145 2860 1146
rect 2854 1141 2855 1145
rect 2859 1141 2860 1145
rect 2854 1140 2860 1141
rect 3006 1145 3012 1146
rect 3006 1141 3007 1145
rect 3011 1141 3012 1145
rect 3006 1140 3012 1141
rect 3158 1145 3164 1146
rect 3158 1141 3159 1145
rect 3163 1141 3164 1145
rect 3158 1140 3164 1141
rect 3318 1145 3324 1146
rect 3318 1141 3319 1145
rect 3323 1141 3324 1145
rect 3318 1140 3324 1141
rect 3478 1145 3484 1146
rect 3478 1141 3479 1145
rect 3483 1141 3484 1145
rect 3478 1140 3484 1141
rect 142 1121 148 1122
rect 142 1117 143 1121
rect 147 1117 148 1121
rect 142 1116 148 1117
rect 294 1121 300 1122
rect 294 1117 295 1121
rect 299 1117 300 1121
rect 294 1116 300 1117
rect 478 1121 484 1122
rect 478 1117 479 1121
rect 483 1117 484 1121
rect 478 1116 484 1117
rect 662 1121 668 1122
rect 662 1117 663 1121
rect 667 1117 668 1121
rect 662 1116 668 1117
rect 846 1121 852 1122
rect 846 1117 847 1121
rect 851 1117 852 1121
rect 846 1116 852 1117
rect 1030 1121 1036 1122
rect 1030 1117 1031 1121
rect 1035 1117 1036 1121
rect 1030 1116 1036 1117
rect 1206 1121 1212 1122
rect 1206 1117 1207 1121
rect 1211 1117 1212 1121
rect 1206 1116 1212 1117
rect 1390 1121 1396 1122
rect 1390 1117 1391 1121
rect 1395 1117 1396 1121
rect 1390 1116 1396 1117
rect 1574 1121 1580 1122
rect 1574 1117 1575 1121
rect 1579 1117 1580 1121
rect 1574 1116 1580 1117
rect 1734 1121 1740 1122
rect 1734 1117 1735 1121
rect 1739 1117 1740 1121
rect 1734 1116 1740 1117
rect 1942 1111 1948 1112
rect 110 1108 116 1109
rect 110 1104 111 1108
rect 115 1104 116 1108
rect 110 1103 116 1104
rect 1822 1108 1828 1109
rect 1822 1104 1823 1108
rect 1827 1104 1828 1108
rect 1942 1107 1943 1111
rect 1947 1107 1948 1111
rect 1942 1106 1948 1107
rect 2086 1111 2092 1112
rect 2086 1107 2087 1111
rect 2091 1107 2092 1111
rect 2086 1106 2092 1107
rect 2230 1111 2236 1112
rect 2230 1107 2231 1111
rect 2235 1107 2236 1111
rect 2230 1106 2236 1107
rect 2382 1111 2388 1112
rect 2382 1107 2383 1111
rect 2387 1107 2388 1111
rect 2382 1106 2388 1107
rect 2534 1111 2540 1112
rect 2534 1107 2535 1111
rect 2539 1107 2540 1111
rect 2534 1106 2540 1107
rect 2686 1111 2692 1112
rect 2686 1107 2687 1111
rect 2691 1107 2692 1111
rect 2686 1106 2692 1107
rect 2838 1111 2844 1112
rect 2838 1107 2839 1111
rect 2843 1107 2844 1111
rect 2838 1106 2844 1107
rect 2990 1111 2996 1112
rect 2990 1107 2991 1111
rect 2995 1107 2996 1111
rect 2990 1106 2996 1107
rect 3150 1111 3156 1112
rect 3150 1107 3151 1111
rect 3155 1107 3156 1111
rect 3150 1106 3156 1107
rect 3318 1111 3324 1112
rect 3318 1107 3319 1111
rect 3323 1107 3324 1111
rect 3318 1106 3324 1107
rect 3478 1111 3484 1112
rect 3478 1107 3479 1111
rect 3483 1107 3484 1111
rect 3478 1106 3484 1107
rect 1822 1103 1828 1104
rect 1862 1101 1868 1102
rect 1862 1097 1863 1101
rect 1867 1097 1868 1101
rect 1862 1096 1868 1097
rect 3574 1101 3580 1102
rect 3574 1097 3575 1101
rect 3579 1097 3580 1101
rect 3574 1096 3580 1097
rect 110 1091 116 1092
rect 110 1087 111 1091
rect 115 1087 116 1091
rect 110 1086 116 1087
rect 1822 1091 1828 1092
rect 1822 1087 1823 1091
rect 1827 1087 1828 1091
rect 1822 1086 1828 1087
rect 1862 1084 1868 1085
rect 134 1081 140 1082
rect 134 1077 135 1081
rect 139 1077 140 1081
rect 134 1076 140 1077
rect 286 1081 292 1082
rect 286 1077 287 1081
rect 291 1077 292 1081
rect 286 1076 292 1077
rect 470 1081 476 1082
rect 470 1077 471 1081
rect 475 1077 476 1081
rect 470 1076 476 1077
rect 654 1081 660 1082
rect 654 1077 655 1081
rect 659 1077 660 1081
rect 654 1076 660 1077
rect 838 1081 844 1082
rect 838 1077 839 1081
rect 843 1077 844 1081
rect 838 1076 844 1077
rect 1022 1081 1028 1082
rect 1022 1077 1023 1081
rect 1027 1077 1028 1081
rect 1022 1076 1028 1077
rect 1198 1081 1204 1082
rect 1198 1077 1199 1081
rect 1203 1077 1204 1081
rect 1198 1076 1204 1077
rect 1382 1081 1388 1082
rect 1382 1077 1383 1081
rect 1387 1077 1388 1081
rect 1382 1076 1388 1077
rect 1566 1081 1572 1082
rect 1566 1077 1567 1081
rect 1571 1077 1572 1081
rect 1566 1076 1572 1077
rect 1726 1081 1732 1082
rect 1726 1077 1727 1081
rect 1731 1077 1732 1081
rect 1862 1080 1863 1084
rect 1867 1080 1868 1084
rect 1862 1079 1868 1080
rect 3574 1084 3580 1085
rect 3574 1080 3575 1084
rect 3579 1080 3580 1084
rect 3574 1079 3580 1080
rect 1726 1076 1732 1077
rect 1950 1071 1956 1072
rect 1950 1067 1951 1071
rect 1955 1067 1956 1071
rect 1950 1066 1956 1067
rect 2094 1071 2100 1072
rect 2094 1067 2095 1071
rect 2099 1067 2100 1071
rect 2094 1066 2100 1067
rect 2238 1071 2244 1072
rect 2238 1067 2239 1071
rect 2243 1067 2244 1071
rect 2238 1066 2244 1067
rect 2390 1071 2396 1072
rect 2390 1067 2391 1071
rect 2395 1067 2396 1071
rect 2390 1066 2396 1067
rect 2542 1071 2548 1072
rect 2542 1067 2543 1071
rect 2547 1067 2548 1071
rect 2542 1066 2548 1067
rect 2694 1071 2700 1072
rect 2694 1067 2695 1071
rect 2699 1067 2700 1071
rect 2694 1066 2700 1067
rect 2846 1071 2852 1072
rect 2846 1067 2847 1071
rect 2851 1067 2852 1071
rect 2846 1066 2852 1067
rect 2998 1071 3004 1072
rect 2998 1067 2999 1071
rect 3003 1067 3004 1071
rect 2998 1066 3004 1067
rect 3158 1071 3164 1072
rect 3158 1067 3159 1071
rect 3163 1067 3164 1071
rect 3158 1066 3164 1067
rect 3326 1071 3332 1072
rect 3326 1067 3327 1071
rect 3331 1067 3332 1071
rect 3326 1066 3332 1067
rect 3486 1071 3492 1072
rect 3486 1067 3487 1071
rect 3491 1067 3492 1071
rect 3486 1066 3492 1067
rect 134 1059 140 1060
rect 134 1055 135 1059
rect 139 1055 140 1059
rect 134 1054 140 1055
rect 270 1059 276 1060
rect 270 1055 271 1059
rect 275 1055 276 1059
rect 270 1054 276 1055
rect 430 1059 436 1060
rect 430 1055 431 1059
rect 435 1055 436 1059
rect 430 1054 436 1055
rect 582 1059 588 1060
rect 582 1055 583 1059
rect 587 1055 588 1059
rect 582 1054 588 1055
rect 734 1059 740 1060
rect 734 1055 735 1059
rect 739 1055 740 1059
rect 734 1054 740 1055
rect 886 1059 892 1060
rect 886 1055 887 1059
rect 891 1055 892 1059
rect 886 1054 892 1055
rect 1046 1059 1052 1060
rect 1046 1055 1047 1059
rect 1051 1055 1052 1059
rect 1046 1054 1052 1055
rect 1214 1059 1220 1060
rect 1214 1055 1215 1059
rect 1219 1055 1220 1059
rect 1214 1054 1220 1055
rect 1382 1059 1388 1060
rect 1382 1055 1383 1059
rect 1387 1055 1388 1059
rect 1382 1054 1388 1055
rect 1558 1059 1564 1060
rect 1558 1055 1559 1059
rect 1563 1055 1564 1059
rect 1558 1054 1564 1055
rect 1726 1059 1732 1060
rect 1726 1055 1727 1059
rect 1731 1055 1732 1059
rect 1726 1054 1732 1055
rect 110 1049 116 1050
rect 110 1045 111 1049
rect 115 1045 116 1049
rect 110 1044 116 1045
rect 1822 1049 1828 1050
rect 1822 1045 1823 1049
rect 1827 1045 1828 1049
rect 1822 1044 1828 1045
rect 110 1032 116 1033
rect 110 1028 111 1032
rect 115 1028 116 1032
rect 110 1027 116 1028
rect 1822 1032 1828 1033
rect 1822 1028 1823 1032
rect 1827 1028 1828 1032
rect 1822 1027 1828 1028
rect 1918 1025 1924 1026
rect 1918 1021 1919 1025
rect 1923 1021 1924 1025
rect 1918 1020 1924 1021
rect 2126 1025 2132 1026
rect 2126 1021 2127 1025
rect 2131 1021 2132 1025
rect 2126 1020 2132 1021
rect 2326 1025 2332 1026
rect 2326 1021 2327 1025
rect 2331 1021 2332 1025
rect 2326 1020 2332 1021
rect 2518 1025 2524 1026
rect 2518 1021 2519 1025
rect 2523 1021 2524 1025
rect 2518 1020 2524 1021
rect 2694 1025 2700 1026
rect 2694 1021 2695 1025
rect 2699 1021 2700 1025
rect 2694 1020 2700 1021
rect 2862 1025 2868 1026
rect 2862 1021 2863 1025
rect 2867 1021 2868 1025
rect 2862 1020 2868 1021
rect 3022 1025 3028 1026
rect 3022 1021 3023 1025
rect 3027 1021 3028 1025
rect 3022 1020 3028 1021
rect 3182 1025 3188 1026
rect 3182 1021 3183 1025
rect 3187 1021 3188 1025
rect 3182 1020 3188 1021
rect 3342 1025 3348 1026
rect 3342 1021 3343 1025
rect 3347 1021 3348 1025
rect 3342 1020 3348 1021
rect 3486 1025 3492 1026
rect 3486 1021 3487 1025
rect 3491 1021 3492 1025
rect 3486 1020 3492 1021
rect 142 1019 148 1020
rect 142 1015 143 1019
rect 147 1015 148 1019
rect 142 1014 148 1015
rect 278 1019 284 1020
rect 278 1015 279 1019
rect 283 1015 284 1019
rect 278 1014 284 1015
rect 438 1019 444 1020
rect 438 1015 439 1019
rect 443 1015 444 1019
rect 438 1014 444 1015
rect 590 1019 596 1020
rect 590 1015 591 1019
rect 595 1015 596 1019
rect 590 1014 596 1015
rect 742 1019 748 1020
rect 742 1015 743 1019
rect 747 1015 748 1019
rect 742 1014 748 1015
rect 894 1019 900 1020
rect 894 1015 895 1019
rect 899 1015 900 1019
rect 894 1014 900 1015
rect 1054 1019 1060 1020
rect 1054 1015 1055 1019
rect 1059 1015 1060 1019
rect 1054 1014 1060 1015
rect 1222 1019 1228 1020
rect 1222 1015 1223 1019
rect 1227 1015 1228 1019
rect 1222 1014 1228 1015
rect 1390 1019 1396 1020
rect 1390 1015 1391 1019
rect 1395 1015 1396 1019
rect 1390 1014 1396 1015
rect 1566 1019 1572 1020
rect 1566 1015 1567 1019
rect 1571 1015 1572 1019
rect 1566 1014 1572 1015
rect 1734 1019 1740 1020
rect 1734 1015 1735 1019
rect 1739 1015 1740 1019
rect 1734 1014 1740 1015
rect 1862 1012 1868 1013
rect 1862 1008 1863 1012
rect 1867 1008 1868 1012
rect 1862 1007 1868 1008
rect 3574 1012 3580 1013
rect 3574 1008 3575 1012
rect 3579 1008 3580 1012
rect 3574 1007 3580 1008
rect 1862 995 1868 996
rect 1862 991 1863 995
rect 1867 991 1868 995
rect 1862 990 1868 991
rect 3574 995 3580 996
rect 3574 991 3575 995
rect 3579 991 3580 995
rect 3574 990 3580 991
rect 1910 985 1916 986
rect 142 981 148 982
rect 142 977 143 981
rect 147 977 148 981
rect 142 976 148 977
rect 286 981 292 982
rect 286 977 287 981
rect 291 977 292 981
rect 286 976 292 977
rect 462 981 468 982
rect 462 977 463 981
rect 467 977 468 981
rect 462 976 468 977
rect 646 981 652 982
rect 646 977 647 981
rect 651 977 652 981
rect 646 976 652 977
rect 822 981 828 982
rect 822 977 823 981
rect 827 977 828 981
rect 822 976 828 977
rect 998 981 1004 982
rect 998 977 999 981
rect 1003 977 1004 981
rect 998 976 1004 977
rect 1166 981 1172 982
rect 1166 977 1167 981
rect 1171 977 1172 981
rect 1166 976 1172 977
rect 1326 981 1332 982
rect 1326 977 1327 981
rect 1331 977 1332 981
rect 1326 976 1332 977
rect 1486 981 1492 982
rect 1486 977 1487 981
rect 1491 977 1492 981
rect 1486 976 1492 977
rect 1654 981 1660 982
rect 1654 977 1655 981
rect 1659 977 1660 981
rect 1910 981 1911 985
rect 1915 981 1916 985
rect 1910 980 1916 981
rect 2118 985 2124 986
rect 2118 981 2119 985
rect 2123 981 2124 985
rect 2118 980 2124 981
rect 2318 985 2324 986
rect 2318 981 2319 985
rect 2323 981 2324 985
rect 2318 980 2324 981
rect 2510 985 2516 986
rect 2510 981 2511 985
rect 2515 981 2516 985
rect 2510 980 2516 981
rect 2686 985 2692 986
rect 2686 981 2687 985
rect 2691 981 2692 985
rect 2686 980 2692 981
rect 2854 985 2860 986
rect 2854 981 2855 985
rect 2859 981 2860 985
rect 2854 980 2860 981
rect 3014 985 3020 986
rect 3014 981 3015 985
rect 3019 981 3020 985
rect 3014 980 3020 981
rect 3174 985 3180 986
rect 3174 981 3175 985
rect 3179 981 3180 985
rect 3174 980 3180 981
rect 3334 985 3340 986
rect 3334 981 3335 985
rect 3339 981 3340 985
rect 3334 980 3340 981
rect 3478 985 3484 986
rect 3478 981 3479 985
rect 3483 981 3484 985
rect 3478 980 3484 981
rect 1654 976 1660 977
rect 110 968 116 969
rect 110 964 111 968
rect 115 964 116 968
rect 110 963 116 964
rect 1822 968 1828 969
rect 1822 964 1823 968
rect 1827 964 1828 968
rect 1822 963 1828 964
rect 1886 959 1892 960
rect 1886 955 1887 959
rect 1891 955 1892 959
rect 1886 954 1892 955
rect 2070 959 2076 960
rect 2070 955 2071 959
rect 2075 955 2076 959
rect 2070 954 2076 955
rect 2262 959 2268 960
rect 2262 955 2263 959
rect 2267 955 2268 959
rect 2262 954 2268 955
rect 2454 959 2460 960
rect 2454 955 2455 959
rect 2459 955 2460 959
rect 2454 954 2460 955
rect 2630 959 2636 960
rect 2630 955 2631 959
rect 2635 955 2636 959
rect 2630 954 2636 955
rect 2798 959 2804 960
rect 2798 955 2799 959
rect 2803 955 2804 959
rect 2798 954 2804 955
rect 2950 959 2956 960
rect 2950 955 2951 959
rect 2955 955 2956 959
rect 2950 954 2956 955
rect 3094 959 3100 960
rect 3094 955 3095 959
rect 3099 955 3100 959
rect 3094 954 3100 955
rect 3230 959 3236 960
rect 3230 955 3231 959
rect 3235 955 3236 959
rect 3230 954 3236 955
rect 3366 959 3372 960
rect 3366 955 3367 959
rect 3371 955 3372 959
rect 3366 954 3372 955
rect 3478 959 3484 960
rect 3478 955 3479 959
rect 3483 955 3484 959
rect 3478 954 3484 955
rect 110 951 116 952
rect 110 947 111 951
rect 115 947 116 951
rect 110 946 116 947
rect 1822 951 1828 952
rect 1822 947 1823 951
rect 1827 947 1828 951
rect 1822 946 1828 947
rect 1862 949 1868 950
rect 1862 945 1863 949
rect 1867 945 1868 949
rect 1862 944 1868 945
rect 3574 949 3580 950
rect 3574 945 3575 949
rect 3579 945 3580 949
rect 3574 944 3580 945
rect 134 941 140 942
rect 134 937 135 941
rect 139 937 140 941
rect 134 936 140 937
rect 278 941 284 942
rect 278 937 279 941
rect 283 937 284 941
rect 278 936 284 937
rect 454 941 460 942
rect 454 937 455 941
rect 459 937 460 941
rect 454 936 460 937
rect 638 941 644 942
rect 638 937 639 941
rect 643 937 644 941
rect 638 936 644 937
rect 814 941 820 942
rect 814 937 815 941
rect 819 937 820 941
rect 814 936 820 937
rect 990 941 996 942
rect 990 937 991 941
rect 995 937 996 941
rect 990 936 996 937
rect 1158 941 1164 942
rect 1158 937 1159 941
rect 1163 937 1164 941
rect 1158 936 1164 937
rect 1318 941 1324 942
rect 1318 937 1319 941
rect 1323 937 1324 941
rect 1318 936 1324 937
rect 1478 941 1484 942
rect 1478 937 1479 941
rect 1483 937 1484 941
rect 1478 936 1484 937
rect 1646 941 1652 942
rect 1646 937 1647 941
rect 1651 937 1652 941
rect 1646 936 1652 937
rect 1862 932 1868 933
rect 1862 928 1863 932
rect 1867 928 1868 932
rect 1862 927 1868 928
rect 3574 932 3580 933
rect 3574 928 3575 932
rect 3579 928 3580 932
rect 3574 927 3580 928
rect 1894 919 1900 920
rect 1894 915 1895 919
rect 1899 915 1900 919
rect 1894 914 1900 915
rect 2078 919 2084 920
rect 2078 915 2079 919
rect 2083 915 2084 919
rect 2078 914 2084 915
rect 2270 919 2276 920
rect 2270 915 2271 919
rect 2275 915 2276 919
rect 2270 914 2276 915
rect 2462 919 2468 920
rect 2462 915 2463 919
rect 2467 915 2468 919
rect 2462 914 2468 915
rect 2638 919 2644 920
rect 2638 915 2639 919
rect 2643 915 2644 919
rect 2638 914 2644 915
rect 2806 919 2812 920
rect 2806 915 2807 919
rect 2811 915 2812 919
rect 2806 914 2812 915
rect 2958 919 2964 920
rect 2958 915 2959 919
rect 2963 915 2964 919
rect 2958 914 2964 915
rect 3102 919 3108 920
rect 3102 915 3103 919
rect 3107 915 3108 919
rect 3102 914 3108 915
rect 3238 919 3244 920
rect 3238 915 3239 919
rect 3243 915 3244 919
rect 3238 914 3244 915
rect 3374 919 3380 920
rect 3374 915 3375 919
rect 3379 915 3380 919
rect 3374 914 3380 915
rect 3486 919 3492 920
rect 3486 915 3487 919
rect 3491 915 3492 919
rect 3486 914 3492 915
rect 134 911 140 912
rect 134 907 135 911
rect 139 907 140 911
rect 134 906 140 907
rect 270 911 276 912
rect 270 907 271 911
rect 275 907 276 911
rect 270 906 276 907
rect 438 911 444 912
rect 438 907 439 911
rect 443 907 444 911
rect 438 906 444 907
rect 606 911 612 912
rect 606 907 607 911
rect 611 907 612 911
rect 606 906 612 907
rect 774 911 780 912
rect 774 907 775 911
rect 779 907 780 911
rect 774 906 780 907
rect 934 911 940 912
rect 934 907 935 911
rect 939 907 940 911
rect 934 906 940 907
rect 1094 911 1100 912
rect 1094 907 1095 911
rect 1099 907 1100 911
rect 1094 906 1100 907
rect 1246 911 1252 912
rect 1246 907 1247 911
rect 1251 907 1252 911
rect 1246 906 1252 907
rect 1398 911 1404 912
rect 1398 907 1399 911
rect 1403 907 1404 911
rect 1398 906 1404 907
rect 1550 911 1556 912
rect 1550 907 1551 911
rect 1555 907 1556 911
rect 1550 906 1556 907
rect 110 901 116 902
rect 110 897 111 901
rect 115 897 116 901
rect 110 896 116 897
rect 1822 901 1828 902
rect 1822 897 1823 901
rect 1827 897 1828 901
rect 1822 896 1828 897
rect 110 884 116 885
rect 110 880 111 884
rect 115 880 116 884
rect 110 879 116 880
rect 1822 884 1828 885
rect 1822 880 1823 884
rect 1827 880 1828 884
rect 1822 879 1828 880
rect 1894 877 1900 878
rect 1894 873 1895 877
rect 1899 873 1900 877
rect 1894 872 1900 873
rect 2022 877 2028 878
rect 2022 873 2023 877
rect 2027 873 2028 877
rect 2022 872 2028 873
rect 2182 877 2188 878
rect 2182 873 2183 877
rect 2187 873 2188 877
rect 2182 872 2188 873
rect 2350 877 2356 878
rect 2350 873 2351 877
rect 2355 873 2356 877
rect 2350 872 2356 873
rect 2518 877 2524 878
rect 2518 873 2519 877
rect 2523 873 2524 877
rect 2518 872 2524 873
rect 2686 877 2692 878
rect 2686 873 2687 877
rect 2691 873 2692 877
rect 2686 872 2692 873
rect 2838 877 2844 878
rect 2838 873 2839 877
rect 2843 873 2844 877
rect 2838 872 2844 873
rect 2982 877 2988 878
rect 2982 873 2983 877
rect 2987 873 2988 877
rect 2982 872 2988 873
rect 3118 877 3124 878
rect 3118 873 3119 877
rect 3123 873 3124 877
rect 3118 872 3124 873
rect 3246 877 3252 878
rect 3246 873 3247 877
rect 3251 873 3252 877
rect 3246 872 3252 873
rect 3374 877 3380 878
rect 3374 873 3375 877
rect 3379 873 3380 877
rect 3374 872 3380 873
rect 3486 877 3492 878
rect 3486 873 3487 877
rect 3491 873 3492 877
rect 3486 872 3492 873
rect 142 871 148 872
rect 142 867 143 871
rect 147 867 148 871
rect 142 866 148 867
rect 278 871 284 872
rect 278 867 279 871
rect 283 867 284 871
rect 278 866 284 867
rect 446 871 452 872
rect 446 867 447 871
rect 451 867 452 871
rect 446 866 452 867
rect 614 871 620 872
rect 614 867 615 871
rect 619 867 620 871
rect 614 866 620 867
rect 782 871 788 872
rect 782 867 783 871
rect 787 867 788 871
rect 782 866 788 867
rect 942 871 948 872
rect 942 867 943 871
rect 947 867 948 871
rect 942 866 948 867
rect 1102 871 1108 872
rect 1102 867 1103 871
rect 1107 867 1108 871
rect 1102 866 1108 867
rect 1254 871 1260 872
rect 1254 867 1255 871
rect 1259 867 1260 871
rect 1254 866 1260 867
rect 1406 871 1412 872
rect 1406 867 1407 871
rect 1411 867 1412 871
rect 1406 866 1412 867
rect 1558 871 1564 872
rect 1558 867 1559 871
rect 1563 867 1564 871
rect 1558 866 1564 867
rect 1862 864 1868 865
rect 1862 860 1863 864
rect 1867 860 1868 864
rect 1862 859 1868 860
rect 3574 864 3580 865
rect 3574 860 3575 864
rect 3579 860 3580 864
rect 3574 859 3580 860
rect 1862 847 1868 848
rect 1862 843 1863 847
rect 1867 843 1868 847
rect 1862 842 1868 843
rect 3574 847 3580 848
rect 3574 843 3575 847
rect 3579 843 3580 847
rect 3574 842 3580 843
rect 142 837 148 838
rect 142 833 143 837
rect 147 833 148 837
rect 142 832 148 833
rect 286 837 292 838
rect 286 833 287 837
rect 291 833 292 837
rect 286 832 292 833
rect 462 837 468 838
rect 462 833 463 837
rect 467 833 468 837
rect 462 832 468 833
rect 638 837 644 838
rect 638 833 639 837
rect 643 833 644 837
rect 638 832 644 833
rect 806 837 812 838
rect 806 833 807 837
rect 811 833 812 837
rect 806 832 812 833
rect 982 837 988 838
rect 982 833 983 837
rect 987 833 988 837
rect 982 832 988 833
rect 1158 837 1164 838
rect 1158 833 1159 837
rect 1163 833 1164 837
rect 1158 832 1164 833
rect 1334 837 1340 838
rect 1334 833 1335 837
rect 1339 833 1340 837
rect 1334 832 1340 833
rect 1510 837 1516 838
rect 1510 833 1511 837
rect 1515 833 1516 837
rect 1510 832 1516 833
rect 1886 837 1892 838
rect 1886 833 1887 837
rect 1891 833 1892 837
rect 1886 832 1892 833
rect 2014 837 2020 838
rect 2014 833 2015 837
rect 2019 833 2020 837
rect 2014 832 2020 833
rect 2174 837 2180 838
rect 2174 833 2175 837
rect 2179 833 2180 837
rect 2174 832 2180 833
rect 2342 837 2348 838
rect 2342 833 2343 837
rect 2347 833 2348 837
rect 2342 832 2348 833
rect 2510 837 2516 838
rect 2510 833 2511 837
rect 2515 833 2516 837
rect 2510 832 2516 833
rect 2678 837 2684 838
rect 2678 833 2679 837
rect 2683 833 2684 837
rect 2678 832 2684 833
rect 2830 837 2836 838
rect 2830 833 2831 837
rect 2835 833 2836 837
rect 2830 832 2836 833
rect 2974 837 2980 838
rect 2974 833 2975 837
rect 2979 833 2980 837
rect 2974 832 2980 833
rect 3110 837 3116 838
rect 3110 833 3111 837
rect 3115 833 3116 837
rect 3110 832 3116 833
rect 3238 837 3244 838
rect 3238 833 3239 837
rect 3243 833 3244 837
rect 3238 832 3244 833
rect 3366 837 3372 838
rect 3366 833 3367 837
rect 3371 833 3372 837
rect 3366 832 3372 833
rect 3478 837 3484 838
rect 3478 833 3479 837
rect 3483 833 3484 837
rect 3478 832 3484 833
rect 110 824 116 825
rect 110 820 111 824
rect 115 820 116 824
rect 110 819 116 820
rect 1822 824 1828 825
rect 1822 820 1823 824
rect 1827 820 1828 824
rect 1822 819 1828 820
rect 110 807 116 808
rect 110 803 111 807
rect 115 803 116 807
rect 110 802 116 803
rect 1822 807 1828 808
rect 1822 803 1823 807
rect 1827 803 1828 807
rect 1822 802 1828 803
rect 1886 807 1892 808
rect 1886 803 1887 807
rect 1891 803 1892 807
rect 1886 802 1892 803
rect 2070 807 2076 808
rect 2070 803 2071 807
rect 2075 803 2076 807
rect 2070 802 2076 803
rect 2262 807 2268 808
rect 2262 803 2263 807
rect 2267 803 2268 807
rect 2262 802 2268 803
rect 2446 807 2452 808
rect 2446 803 2447 807
rect 2451 803 2452 807
rect 2446 802 2452 803
rect 2622 807 2628 808
rect 2622 803 2623 807
rect 2627 803 2628 807
rect 2622 802 2628 803
rect 2790 807 2796 808
rect 2790 803 2791 807
rect 2795 803 2796 807
rect 2790 802 2796 803
rect 2942 807 2948 808
rect 2942 803 2943 807
rect 2947 803 2948 807
rect 2942 802 2948 803
rect 3086 807 3092 808
rect 3086 803 3087 807
rect 3091 803 3092 807
rect 3086 802 3092 803
rect 3222 807 3228 808
rect 3222 803 3223 807
rect 3227 803 3228 807
rect 3222 802 3228 803
rect 3358 807 3364 808
rect 3358 803 3359 807
rect 3363 803 3364 807
rect 3358 802 3364 803
rect 3478 807 3484 808
rect 3478 803 3479 807
rect 3483 803 3484 807
rect 3478 802 3484 803
rect 134 797 140 798
rect 134 793 135 797
rect 139 793 140 797
rect 134 792 140 793
rect 278 797 284 798
rect 278 793 279 797
rect 283 793 284 797
rect 278 792 284 793
rect 454 797 460 798
rect 454 793 455 797
rect 459 793 460 797
rect 454 792 460 793
rect 630 797 636 798
rect 630 793 631 797
rect 635 793 636 797
rect 630 792 636 793
rect 798 797 804 798
rect 798 793 799 797
rect 803 793 804 797
rect 798 792 804 793
rect 974 797 980 798
rect 974 793 975 797
rect 979 793 980 797
rect 974 792 980 793
rect 1150 797 1156 798
rect 1150 793 1151 797
rect 1155 793 1156 797
rect 1150 792 1156 793
rect 1326 797 1332 798
rect 1326 793 1327 797
rect 1331 793 1332 797
rect 1326 792 1332 793
rect 1502 797 1508 798
rect 1502 793 1503 797
rect 1507 793 1508 797
rect 1502 792 1508 793
rect 1862 797 1868 798
rect 1862 793 1863 797
rect 1867 793 1868 797
rect 1862 792 1868 793
rect 3574 797 3580 798
rect 3574 793 3575 797
rect 3579 793 3580 797
rect 3574 792 3580 793
rect 1862 780 1868 781
rect 1862 776 1863 780
rect 1867 776 1868 780
rect 1862 775 1868 776
rect 3574 780 3580 781
rect 3574 776 3575 780
rect 3579 776 3580 780
rect 3574 775 3580 776
rect 134 771 140 772
rect 134 767 135 771
rect 139 767 140 771
rect 134 766 140 767
rect 270 771 276 772
rect 270 767 271 771
rect 275 767 276 771
rect 270 766 276 767
rect 438 771 444 772
rect 438 767 439 771
rect 443 767 444 771
rect 438 766 444 767
rect 606 771 612 772
rect 606 767 607 771
rect 611 767 612 771
rect 606 766 612 767
rect 774 771 780 772
rect 774 767 775 771
rect 779 767 780 771
rect 774 766 780 767
rect 934 771 940 772
rect 934 767 935 771
rect 939 767 940 771
rect 934 766 940 767
rect 1086 771 1092 772
rect 1086 767 1087 771
rect 1091 767 1092 771
rect 1086 766 1092 767
rect 1238 771 1244 772
rect 1238 767 1239 771
rect 1243 767 1244 771
rect 1238 766 1244 767
rect 1390 771 1396 772
rect 1390 767 1391 771
rect 1395 767 1396 771
rect 1390 766 1396 767
rect 1550 771 1556 772
rect 1550 767 1551 771
rect 1555 767 1556 771
rect 1550 766 1556 767
rect 1894 767 1900 768
rect 1894 763 1895 767
rect 1899 763 1900 767
rect 1894 762 1900 763
rect 2078 767 2084 768
rect 2078 763 2079 767
rect 2083 763 2084 767
rect 2078 762 2084 763
rect 2270 767 2276 768
rect 2270 763 2271 767
rect 2275 763 2276 767
rect 2270 762 2276 763
rect 2454 767 2460 768
rect 2454 763 2455 767
rect 2459 763 2460 767
rect 2454 762 2460 763
rect 2630 767 2636 768
rect 2630 763 2631 767
rect 2635 763 2636 767
rect 2630 762 2636 763
rect 2798 767 2804 768
rect 2798 763 2799 767
rect 2803 763 2804 767
rect 2798 762 2804 763
rect 2950 767 2956 768
rect 2950 763 2951 767
rect 2955 763 2956 767
rect 2950 762 2956 763
rect 3094 767 3100 768
rect 3094 763 3095 767
rect 3099 763 3100 767
rect 3094 762 3100 763
rect 3230 767 3236 768
rect 3230 763 3231 767
rect 3235 763 3236 767
rect 3230 762 3236 763
rect 3366 767 3372 768
rect 3366 763 3367 767
rect 3371 763 3372 767
rect 3366 762 3372 763
rect 3486 767 3492 768
rect 3486 763 3487 767
rect 3491 763 3492 767
rect 3486 762 3492 763
rect 110 761 116 762
rect 110 757 111 761
rect 115 757 116 761
rect 110 756 116 757
rect 1822 761 1828 762
rect 1822 757 1823 761
rect 1827 757 1828 761
rect 1822 756 1828 757
rect 110 744 116 745
rect 110 740 111 744
rect 115 740 116 744
rect 110 739 116 740
rect 1822 744 1828 745
rect 1822 740 1823 744
rect 1827 740 1828 744
rect 1822 739 1828 740
rect 1894 733 1900 734
rect 142 731 148 732
rect 142 727 143 731
rect 147 727 148 731
rect 142 726 148 727
rect 278 731 284 732
rect 278 727 279 731
rect 283 727 284 731
rect 278 726 284 727
rect 446 731 452 732
rect 446 727 447 731
rect 451 727 452 731
rect 446 726 452 727
rect 614 731 620 732
rect 614 727 615 731
rect 619 727 620 731
rect 614 726 620 727
rect 782 731 788 732
rect 782 727 783 731
rect 787 727 788 731
rect 782 726 788 727
rect 942 731 948 732
rect 942 727 943 731
rect 947 727 948 731
rect 942 726 948 727
rect 1094 731 1100 732
rect 1094 727 1095 731
rect 1099 727 1100 731
rect 1094 726 1100 727
rect 1246 731 1252 732
rect 1246 727 1247 731
rect 1251 727 1252 731
rect 1246 726 1252 727
rect 1398 731 1404 732
rect 1398 727 1399 731
rect 1403 727 1404 731
rect 1398 726 1404 727
rect 1558 731 1564 732
rect 1558 727 1559 731
rect 1563 727 1564 731
rect 1894 729 1895 733
rect 1899 729 1900 733
rect 1894 728 1900 729
rect 2070 733 2076 734
rect 2070 729 2071 733
rect 2075 729 2076 733
rect 2070 728 2076 729
rect 2262 733 2268 734
rect 2262 729 2263 733
rect 2267 729 2268 733
rect 2262 728 2268 729
rect 2446 733 2452 734
rect 2446 729 2447 733
rect 2451 729 2452 733
rect 2446 728 2452 729
rect 2622 733 2628 734
rect 2622 729 2623 733
rect 2627 729 2628 733
rect 2622 728 2628 729
rect 2798 733 2804 734
rect 2798 729 2799 733
rect 2803 729 2804 733
rect 2798 728 2804 729
rect 2974 733 2980 734
rect 2974 729 2975 733
rect 2979 729 2980 733
rect 2974 728 2980 729
rect 3150 733 3156 734
rect 3150 729 3151 733
rect 3155 729 3156 733
rect 3150 728 3156 729
rect 3326 733 3332 734
rect 3326 729 3327 733
rect 3331 729 3332 733
rect 3326 728 3332 729
rect 3486 733 3492 734
rect 3486 729 3487 733
rect 3491 729 3492 733
rect 3486 728 3492 729
rect 1558 726 1564 727
rect 1862 720 1868 721
rect 1862 716 1863 720
rect 1867 716 1868 720
rect 1862 715 1868 716
rect 3574 720 3580 721
rect 3574 716 3575 720
rect 3579 716 3580 720
rect 3574 715 3580 716
rect 1862 703 1868 704
rect 1862 699 1863 703
rect 1867 699 1868 703
rect 1862 698 1868 699
rect 3574 703 3580 704
rect 3574 699 3575 703
rect 3579 699 3580 703
rect 3574 698 3580 699
rect 142 693 148 694
rect 142 689 143 693
rect 147 689 148 693
rect 142 688 148 689
rect 286 693 292 694
rect 286 689 287 693
rect 291 689 292 693
rect 286 688 292 689
rect 454 693 460 694
rect 454 689 455 693
rect 459 689 460 693
rect 454 688 460 689
rect 622 693 628 694
rect 622 689 623 693
rect 627 689 628 693
rect 622 688 628 689
rect 790 693 796 694
rect 790 689 791 693
rect 795 689 796 693
rect 790 688 796 689
rect 958 693 964 694
rect 958 689 959 693
rect 963 689 964 693
rect 958 688 964 689
rect 1118 693 1124 694
rect 1118 689 1119 693
rect 1123 689 1124 693
rect 1118 688 1124 689
rect 1278 693 1284 694
rect 1278 689 1279 693
rect 1283 689 1284 693
rect 1278 688 1284 689
rect 1438 693 1444 694
rect 1438 689 1439 693
rect 1443 689 1444 693
rect 1438 688 1444 689
rect 1598 693 1604 694
rect 1598 689 1599 693
rect 1603 689 1604 693
rect 1598 688 1604 689
rect 1886 693 1892 694
rect 1886 689 1887 693
rect 1891 689 1892 693
rect 1886 688 1892 689
rect 2062 693 2068 694
rect 2062 689 2063 693
rect 2067 689 2068 693
rect 2062 688 2068 689
rect 2254 693 2260 694
rect 2254 689 2255 693
rect 2259 689 2260 693
rect 2254 688 2260 689
rect 2438 693 2444 694
rect 2438 689 2439 693
rect 2443 689 2444 693
rect 2438 688 2444 689
rect 2614 693 2620 694
rect 2614 689 2615 693
rect 2619 689 2620 693
rect 2614 688 2620 689
rect 2790 693 2796 694
rect 2790 689 2791 693
rect 2795 689 2796 693
rect 2790 688 2796 689
rect 2966 693 2972 694
rect 2966 689 2967 693
rect 2971 689 2972 693
rect 2966 688 2972 689
rect 3142 693 3148 694
rect 3142 689 3143 693
rect 3147 689 3148 693
rect 3142 688 3148 689
rect 3318 693 3324 694
rect 3318 689 3319 693
rect 3323 689 3324 693
rect 3318 688 3324 689
rect 3478 693 3484 694
rect 3478 689 3479 693
rect 3483 689 3484 693
rect 3478 688 3484 689
rect 110 680 116 681
rect 110 676 111 680
rect 115 676 116 680
rect 110 675 116 676
rect 1822 680 1828 681
rect 1822 676 1823 680
rect 1827 676 1828 680
rect 1822 675 1828 676
rect 1886 667 1892 668
rect 110 663 116 664
rect 110 659 111 663
rect 115 659 116 663
rect 110 658 116 659
rect 1822 663 1828 664
rect 1822 659 1823 663
rect 1827 659 1828 663
rect 1886 663 1887 667
rect 1891 663 1892 667
rect 1886 662 1892 663
rect 1974 667 1980 668
rect 1974 663 1975 667
rect 1979 663 1980 667
rect 1974 662 1980 663
rect 2094 667 2100 668
rect 2094 663 2095 667
rect 2099 663 2100 667
rect 2094 662 2100 663
rect 2222 667 2228 668
rect 2222 663 2223 667
rect 2227 663 2228 667
rect 2222 662 2228 663
rect 2350 667 2356 668
rect 2350 663 2351 667
rect 2355 663 2356 667
rect 2350 662 2356 663
rect 2478 667 2484 668
rect 2478 663 2479 667
rect 2483 663 2484 667
rect 2478 662 2484 663
rect 2614 667 2620 668
rect 2614 663 2615 667
rect 2619 663 2620 667
rect 2614 662 2620 663
rect 2766 667 2772 668
rect 2766 663 2767 667
rect 2771 663 2772 667
rect 2766 662 2772 663
rect 2934 667 2940 668
rect 2934 663 2935 667
rect 2939 663 2940 667
rect 2934 662 2940 663
rect 3118 667 3124 668
rect 3118 663 3119 667
rect 3123 663 3124 667
rect 3118 662 3124 663
rect 3310 667 3316 668
rect 3310 663 3311 667
rect 3315 663 3316 667
rect 3310 662 3316 663
rect 3478 667 3484 668
rect 3478 663 3479 667
rect 3483 663 3484 667
rect 3478 662 3484 663
rect 1822 658 1828 659
rect 1862 657 1868 658
rect 134 653 140 654
rect 134 649 135 653
rect 139 649 140 653
rect 134 648 140 649
rect 278 653 284 654
rect 278 649 279 653
rect 283 649 284 653
rect 278 648 284 649
rect 446 653 452 654
rect 446 649 447 653
rect 451 649 452 653
rect 446 648 452 649
rect 614 653 620 654
rect 614 649 615 653
rect 619 649 620 653
rect 614 648 620 649
rect 782 653 788 654
rect 782 649 783 653
rect 787 649 788 653
rect 782 648 788 649
rect 950 653 956 654
rect 950 649 951 653
rect 955 649 956 653
rect 950 648 956 649
rect 1110 653 1116 654
rect 1110 649 1111 653
rect 1115 649 1116 653
rect 1110 648 1116 649
rect 1270 653 1276 654
rect 1270 649 1271 653
rect 1275 649 1276 653
rect 1270 648 1276 649
rect 1430 653 1436 654
rect 1430 649 1431 653
rect 1435 649 1436 653
rect 1430 648 1436 649
rect 1590 653 1596 654
rect 1590 649 1591 653
rect 1595 649 1596 653
rect 1862 653 1863 657
rect 1867 653 1868 657
rect 1862 652 1868 653
rect 3574 657 3580 658
rect 3574 653 3575 657
rect 3579 653 3580 657
rect 3574 652 3580 653
rect 1590 648 1596 649
rect 1862 640 1868 641
rect 1862 636 1863 640
rect 1867 636 1868 640
rect 1862 635 1868 636
rect 3574 640 3580 641
rect 3574 636 3575 640
rect 3579 636 3580 640
rect 3574 635 3580 636
rect 1894 627 1900 628
rect 134 623 140 624
rect 134 619 135 623
rect 139 619 140 623
rect 134 618 140 619
rect 286 623 292 624
rect 286 619 287 623
rect 291 619 292 623
rect 286 618 292 619
rect 454 623 460 624
rect 454 619 455 623
rect 459 619 460 623
rect 454 618 460 619
rect 630 623 636 624
rect 630 619 631 623
rect 635 619 636 623
rect 630 618 636 619
rect 798 623 804 624
rect 798 619 799 623
rect 803 619 804 623
rect 798 618 804 619
rect 966 623 972 624
rect 966 619 967 623
rect 971 619 972 623
rect 966 618 972 619
rect 1118 623 1124 624
rect 1118 619 1119 623
rect 1123 619 1124 623
rect 1118 618 1124 619
rect 1270 623 1276 624
rect 1270 619 1271 623
rect 1275 619 1276 623
rect 1270 618 1276 619
rect 1414 623 1420 624
rect 1414 619 1415 623
rect 1419 619 1420 623
rect 1414 618 1420 619
rect 1558 623 1564 624
rect 1558 619 1559 623
rect 1563 619 1564 623
rect 1558 618 1564 619
rect 1710 623 1716 624
rect 1710 619 1711 623
rect 1715 619 1716 623
rect 1894 623 1895 627
rect 1899 623 1900 627
rect 1894 622 1900 623
rect 1982 627 1988 628
rect 1982 623 1983 627
rect 1987 623 1988 627
rect 1982 622 1988 623
rect 2102 627 2108 628
rect 2102 623 2103 627
rect 2107 623 2108 627
rect 2102 622 2108 623
rect 2230 627 2236 628
rect 2230 623 2231 627
rect 2235 623 2236 627
rect 2230 622 2236 623
rect 2358 627 2364 628
rect 2358 623 2359 627
rect 2363 623 2364 627
rect 2358 622 2364 623
rect 2486 627 2492 628
rect 2486 623 2487 627
rect 2491 623 2492 627
rect 2486 622 2492 623
rect 2622 627 2628 628
rect 2622 623 2623 627
rect 2627 623 2628 627
rect 2622 622 2628 623
rect 2774 627 2780 628
rect 2774 623 2775 627
rect 2779 623 2780 627
rect 2774 622 2780 623
rect 2942 627 2948 628
rect 2942 623 2943 627
rect 2947 623 2948 627
rect 2942 622 2948 623
rect 3126 627 3132 628
rect 3126 623 3127 627
rect 3131 623 3132 627
rect 3126 622 3132 623
rect 3318 627 3324 628
rect 3318 623 3319 627
rect 3323 623 3324 627
rect 3318 622 3324 623
rect 3486 627 3492 628
rect 3486 623 3487 627
rect 3491 623 3492 627
rect 3486 622 3492 623
rect 1710 618 1716 619
rect 110 613 116 614
rect 110 609 111 613
rect 115 609 116 613
rect 110 608 116 609
rect 1822 613 1828 614
rect 1822 609 1823 613
rect 1827 609 1828 613
rect 1822 608 1828 609
rect 110 596 116 597
rect 110 592 111 596
rect 115 592 116 596
rect 110 591 116 592
rect 1822 596 1828 597
rect 1822 592 1823 596
rect 1827 592 1828 596
rect 1822 591 1828 592
rect 1894 589 1900 590
rect 1894 585 1895 589
rect 1899 585 1900 589
rect 1894 584 1900 585
rect 2046 589 2052 590
rect 2046 585 2047 589
rect 2051 585 2052 589
rect 2046 584 2052 585
rect 2214 589 2220 590
rect 2214 585 2215 589
rect 2219 585 2220 589
rect 2214 584 2220 585
rect 2390 589 2396 590
rect 2390 585 2391 589
rect 2395 585 2396 589
rect 2390 584 2396 585
rect 2582 589 2588 590
rect 2582 585 2583 589
rect 2587 585 2588 589
rect 2582 584 2588 585
rect 2798 589 2804 590
rect 2798 585 2799 589
rect 2803 585 2804 589
rect 2798 584 2804 585
rect 3022 589 3028 590
rect 3022 585 3023 589
rect 3027 585 3028 589
rect 3022 584 3028 585
rect 3254 589 3260 590
rect 3254 585 3255 589
rect 3259 585 3260 589
rect 3254 584 3260 585
rect 3486 589 3492 590
rect 3486 585 3487 589
rect 3491 585 3492 589
rect 3486 584 3492 585
rect 142 583 148 584
rect 142 579 143 583
rect 147 579 148 583
rect 142 578 148 579
rect 294 583 300 584
rect 294 579 295 583
rect 299 579 300 583
rect 294 578 300 579
rect 462 583 468 584
rect 462 579 463 583
rect 467 579 468 583
rect 462 578 468 579
rect 638 583 644 584
rect 638 579 639 583
rect 643 579 644 583
rect 638 578 644 579
rect 806 583 812 584
rect 806 579 807 583
rect 811 579 812 583
rect 806 578 812 579
rect 974 583 980 584
rect 974 579 975 583
rect 979 579 980 583
rect 974 578 980 579
rect 1126 583 1132 584
rect 1126 579 1127 583
rect 1131 579 1132 583
rect 1126 578 1132 579
rect 1278 583 1284 584
rect 1278 579 1279 583
rect 1283 579 1284 583
rect 1278 578 1284 579
rect 1422 583 1428 584
rect 1422 579 1423 583
rect 1427 579 1428 583
rect 1422 578 1428 579
rect 1566 583 1572 584
rect 1566 579 1567 583
rect 1571 579 1572 583
rect 1566 578 1572 579
rect 1718 583 1724 584
rect 1718 579 1719 583
rect 1723 579 1724 583
rect 1718 578 1724 579
rect 1862 576 1868 577
rect 1862 572 1863 576
rect 1867 572 1868 576
rect 1862 571 1868 572
rect 3574 576 3580 577
rect 3574 572 3575 576
rect 3579 572 3580 576
rect 3574 571 3580 572
rect 1862 559 1868 560
rect 1862 555 1863 559
rect 1867 555 1868 559
rect 1862 554 1868 555
rect 3574 559 3580 560
rect 3574 555 3575 559
rect 3579 555 3580 559
rect 3574 554 3580 555
rect 1886 549 1892 550
rect 150 545 156 546
rect 150 541 151 545
rect 155 541 156 545
rect 150 540 156 541
rect 310 545 316 546
rect 310 541 311 545
rect 315 541 316 545
rect 310 540 316 541
rect 470 545 476 546
rect 470 541 471 545
rect 475 541 476 545
rect 470 540 476 541
rect 630 545 636 546
rect 630 541 631 545
rect 635 541 636 545
rect 630 540 636 541
rect 782 545 788 546
rect 782 541 783 545
rect 787 541 788 545
rect 782 540 788 541
rect 926 545 932 546
rect 926 541 927 545
rect 931 541 932 545
rect 926 540 932 541
rect 1062 545 1068 546
rect 1062 541 1063 545
rect 1067 541 1068 545
rect 1062 540 1068 541
rect 1190 545 1196 546
rect 1190 541 1191 545
rect 1195 541 1196 545
rect 1190 540 1196 541
rect 1310 545 1316 546
rect 1310 541 1311 545
rect 1315 541 1316 545
rect 1310 540 1316 541
rect 1422 545 1428 546
rect 1422 541 1423 545
rect 1427 541 1428 545
rect 1422 540 1428 541
rect 1534 545 1540 546
rect 1534 541 1535 545
rect 1539 541 1540 545
rect 1534 540 1540 541
rect 1646 545 1652 546
rect 1646 541 1647 545
rect 1651 541 1652 545
rect 1646 540 1652 541
rect 1734 545 1740 546
rect 1734 541 1735 545
rect 1739 541 1740 545
rect 1886 545 1887 549
rect 1891 545 1892 549
rect 1886 544 1892 545
rect 2038 549 2044 550
rect 2038 545 2039 549
rect 2043 545 2044 549
rect 2038 544 2044 545
rect 2206 549 2212 550
rect 2206 545 2207 549
rect 2211 545 2212 549
rect 2206 544 2212 545
rect 2382 549 2388 550
rect 2382 545 2383 549
rect 2387 545 2388 549
rect 2382 544 2388 545
rect 2574 549 2580 550
rect 2574 545 2575 549
rect 2579 545 2580 549
rect 2574 544 2580 545
rect 2790 549 2796 550
rect 2790 545 2791 549
rect 2795 545 2796 549
rect 2790 544 2796 545
rect 3014 549 3020 550
rect 3014 545 3015 549
rect 3019 545 3020 549
rect 3014 544 3020 545
rect 3246 549 3252 550
rect 3246 545 3247 549
rect 3251 545 3252 549
rect 3246 544 3252 545
rect 3478 549 3484 550
rect 3478 545 3479 549
rect 3483 545 3484 549
rect 3478 544 3484 545
rect 1734 540 1740 541
rect 110 532 116 533
rect 110 528 111 532
rect 115 528 116 532
rect 110 527 116 528
rect 1822 532 1828 533
rect 1822 528 1823 532
rect 1827 528 1828 532
rect 1822 527 1828 528
rect 2190 519 2196 520
rect 110 515 116 516
rect 110 511 111 515
rect 115 511 116 515
rect 110 510 116 511
rect 1822 515 1828 516
rect 1822 511 1823 515
rect 1827 511 1828 515
rect 2190 515 2191 519
rect 2195 515 2196 519
rect 2190 514 2196 515
rect 2278 519 2284 520
rect 2278 515 2279 519
rect 2283 515 2284 519
rect 2278 514 2284 515
rect 2374 519 2380 520
rect 2374 515 2375 519
rect 2379 515 2380 519
rect 2374 514 2380 515
rect 2486 519 2492 520
rect 2486 515 2487 519
rect 2491 515 2492 519
rect 2486 514 2492 515
rect 2630 519 2636 520
rect 2630 515 2631 519
rect 2635 515 2636 519
rect 2630 514 2636 515
rect 2806 519 2812 520
rect 2806 515 2807 519
rect 2811 515 2812 519
rect 2806 514 2812 515
rect 3006 519 3012 520
rect 3006 515 3007 519
rect 3011 515 3012 519
rect 3006 514 3012 515
rect 3214 519 3220 520
rect 3214 515 3215 519
rect 3219 515 3220 519
rect 3214 514 3220 515
rect 3430 519 3436 520
rect 3430 515 3431 519
rect 3435 515 3436 519
rect 3430 514 3436 515
rect 1822 510 1828 511
rect 1862 509 1868 510
rect 142 505 148 506
rect 142 501 143 505
rect 147 501 148 505
rect 142 500 148 501
rect 302 505 308 506
rect 302 501 303 505
rect 307 501 308 505
rect 302 500 308 501
rect 462 505 468 506
rect 462 501 463 505
rect 467 501 468 505
rect 462 500 468 501
rect 622 505 628 506
rect 622 501 623 505
rect 627 501 628 505
rect 622 500 628 501
rect 774 505 780 506
rect 774 501 775 505
rect 779 501 780 505
rect 774 500 780 501
rect 918 505 924 506
rect 918 501 919 505
rect 923 501 924 505
rect 918 500 924 501
rect 1054 505 1060 506
rect 1054 501 1055 505
rect 1059 501 1060 505
rect 1054 500 1060 501
rect 1182 505 1188 506
rect 1182 501 1183 505
rect 1187 501 1188 505
rect 1182 500 1188 501
rect 1302 505 1308 506
rect 1302 501 1303 505
rect 1307 501 1308 505
rect 1302 500 1308 501
rect 1414 505 1420 506
rect 1414 501 1415 505
rect 1419 501 1420 505
rect 1414 500 1420 501
rect 1526 505 1532 506
rect 1526 501 1527 505
rect 1531 501 1532 505
rect 1526 500 1532 501
rect 1638 505 1644 506
rect 1638 501 1639 505
rect 1643 501 1644 505
rect 1638 500 1644 501
rect 1726 505 1732 506
rect 1726 501 1727 505
rect 1731 501 1732 505
rect 1862 505 1863 509
rect 1867 505 1868 509
rect 1862 504 1868 505
rect 3574 509 3580 510
rect 3574 505 3575 509
rect 3579 505 3580 509
rect 3574 504 3580 505
rect 1726 500 1732 501
rect 1862 492 1868 493
rect 1862 488 1863 492
rect 1867 488 1868 492
rect 1862 487 1868 488
rect 3574 492 3580 493
rect 3574 488 3575 492
rect 3579 488 3580 492
rect 3574 487 3580 488
rect 2198 479 2204 480
rect 158 475 164 476
rect 158 471 159 475
rect 163 471 164 475
rect 158 470 164 471
rect 310 475 316 476
rect 310 471 311 475
rect 315 471 316 475
rect 310 470 316 471
rect 462 475 468 476
rect 462 471 463 475
rect 467 471 468 475
rect 462 470 468 471
rect 614 475 620 476
rect 614 471 615 475
rect 619 471 620 475
rect 614 470 620 471
rect 758 475 764 476
rect 758 471 759 475
rect 763 471 764 475
rect 758 470 764 471
rect 886 475 892 476
rect 886 471 887 475
rect 891 471 892 475
rect 886 470 892 471
rect 1006 475 1012 476
rect 1006 471 1007 475
rect 1011 471 1012 475
rect 1006 470 1012 471
rect 1126 475 1132 476
rect 1126 471 1127 475
rect 1131 471 1132 475
rect 1126 470 1132 471
rect 1238 475 1244 476
rect 1238 471 1239 475
rect 1243 471 1244 475
rect 1238 470 1244 471
rect 1342 475 1348 476
rect 1342 471 1343 475
rect 1347 471 1348 475
rect 1342 470 1348 471
rect 1438 475 1444 476
rect 1438 471 1439 475
rect 1443 471 1444 475
rect 1438 470 1444 471
rect 1542 475 1548 476
rect 1542 471 1543 475
rect 1547 471 1548 475
rect 1542 470 1548 471
rect 1638 475 1644 476
rect 1638 471 1639 475
rect 1643 471 1644 475
rect 1638 470 1644 471
rect 1726 475 1732 476
rect 1726 471 1727 475
rect 1731 471 1732 475
rect 2198 475 2199 479
rect 2203 475 2204 479
rect 2198 474 2204 475
rect 2286 479 2292 480
rect 2286 475 2287 479
rect 2291 475 2292 479
rect 2286 474 2292 475
rect 2382 479 2388 480
rect 2382 475 2383 479
rect 2387 475 2388 479
rect 2382 474 2388 475
rect 2494 479 2500 480
rect 2494 475 2495 479
rect 2499 475 2500 479
rect 2494 474 2500 475
rect 2638 479 2644 480
rect 2638 475 2639 479
rect 2643 475 2644 479
rect 2638 474 2644 475
rect 2814 479 2820 480
rect 2814 475 2815 479
rect 2819 475 2820 479
rect 2814 474 2820 475
rect 3014 479 3020 480
rect 3014 475 3015 479
rect 3019 475 3020 479
rect 3014 474 3020 475
rect 3222 479 3228 480
rect 3222 475 3223 479
rect 3227 475 3228 479
rect 3222 474 3228 475
rect 3438 479 3444 480
rect 3438 475 3439 479
rect 3443 475 3444 479
rect 3438 474 3444 475
rect 1726 470 1732 471
rect 110 465 116 466
rect 110 461 111 465
rect 115 461 116 465
rect 110 460 116 461
rect 1822 465 1828 466
rect 1822 461 1823 465
rect 1827 461 1828 465
rect 1822 460 1828 461
rect 110 448 116 449
rect 110 444 111 448
rect 115 444 116 448
rect 110 443 116 444
rect 1822 448 1828 449
rect 1822 444 1823 448
rect 1827 444 1828 448
rect 1822 443 1828 444
rect 1894 437 1900 438
rect 166 435 172 436
rect 166 431 167 435
rect 171 431 172 435
rect 166 430 172 431
rect 318 435 324 436
rect 318 431 319 435
rect 323 431 324 435
rect 318 430 324 431
rect 470 435 476 436
rect 470 431 471 435
rect 475 431 476 435
rect 470 430 476 431
rect 622 435 628 436
rect 622 431 623 435
rect 627 431 628 435
rect 622 430 628 431
rect 766 435 772 436
rect 766 431 767 435
rect 771 431 772 435
rect 766 430 772 431
rect 894 435 900 436
rect 894 431 895 435
rect 899 431 900 435
rect 894 430 900 431
rect 1014 435 1020 436
rect 1014 431 1015 435
rect 1019 431 1020 435
rect 1014 430 1020 431
rect 1134 435 1140 436
rect 1134 431 1135 435
rect 1139 431 1140 435
rect 1134 430 1140 431
rect 1246 435 1252 436
rect 1246 431 1247 435
rect 1251 431 1252 435
rect 1246 430 1252 431
rect 1350 435 1356 436
rect 1350 431 1351 435
rect 1355 431 1356 435
rect 1350 430 1356 431
rect 1446 435 1452 436
rect 1446 431 1447 435
rect 1451 431 1452 435
rect 1446 430 1452 431
rect 1550 435 1556 436
rect 1550 431 1551 435
rect 1555 431 1556 435
rect 1550 430 1556 431
rect 1646 435 1652 436
rect 1646 431 1647 435
rect 1651 431 1652 435
rect 1646 430 1652 431
rect 1734 435 1740 436
rect 1734 431 1735 435
rect 1739 431 1740 435
rect 1894 433 1895 437
rect 1899 433 1900 437
rect 1894 432 1900 433
rect 2038 437 2044 438
rect 2038 433 2039 437
rect 2043 433 2044 437
rect 2038 432 2044 433
rect 2206 437 2212 438
rect 2206 433 2207 437
rect 2211 433 2212 437
rect 2206 432 2212 433
rect 2382 437 2388 438
rect 2382 433 2383 437
rect 2387 433 2388 437
rect 2382 432 2388 433
rect 2574 437 2580 438
rect 2574 433 2575 437
rect 2579 433 2580 437
rect 2574 432 2580 433
rect 2782 437 2788 438
rect 2782 433 2783 437
rect 2787 433 2788 437
rect 2782 432 2788 433
rect 3006 437 3012 438
rect 3006 433 3007 437
rect 3011 433 3012 437
rect 3006 432 3012 433
rect 3238 437 3244 438
rect 3238 433 3239 437
rect 3243 433 3244 437
rect 3238 432 3244 433
rect 3470 437 3476 438
rect 3470 433 3471 437
rect 3475 433 3476 437
rect 3470 432 3476 433
rect 1734 430 1740 431
rect 1862 424 1868 425
rect 1862 420 1863 424
rect 1867 420 1868 424
rect 1862 419 1868 420
rect 3574 424 3580 425
rect 3574 420 3575 424
rect 3579 420 3580 424
rect 3574 419 3580 420
rect 1862 407 1868 408
rect 1862 403 1863 407
rect 1867 403 1868 407
rect 1862 402 1868 403
rect 3574 407 3580 408
rect 3574 403 3575 407
rect 3579 403 3580 407
rect 3574 402 3580 403
rect 150 401 156 402
rect 150 397 151 401
rect 155 397 156 401
rect 150 396 156 397
rect 270 401 276 402
rect 270 397 271 401
rect 275 397 276 401
rect 270 396 276 397
rect 406 401 412 402
rect 406 397 407 401
rect 411 397 412 401
rect 406 396 412 397
rect 550 401 556 402
rect 550 397 551 401
rect 555 397 556 401
rect 550 396 556 397
rect 710 401 716 402
rect 710 397 711 401
rect 715 397 716 401
rect 710 396 716 397
rect 886 401 892 402
rect 886 397 887 401
rect 891 397 892 401
rect 886 396 892 397
rect 1062 401 1068 402
rect 1062 397 1063 401
rect 1067 397 1068 401
rect 1062 396 1068 397
rect 1246 401 1252 402
rect 1246 397 1247 401
rect 1251 397 1252 401
rect 1246 396 1252 397
rect 1438 401 1444 402
rect 1438 397 1439 401
rect 1443 397 1444 401
rect 1438 396 1444 397
rect 1638 401 1644 402
rect 1638 397 1639 401
rect 1643 397 1644 401
rect 1638 396 1644 397
rect 1886 397 1892 398
rect 1886 393 1887 397
rect 1891 393 1892 397
rect 1886 392 1892 393
rect 2030 397 2036 398
rect 2030 393 2031 397
rect 2035 393 2036 397
rect 2030 392 2036 393
rect 2198 397 2204 398
rect 2198 393 2199 397
rect 2203 393 2204 397
rect 2198 392 2204 393
rect 2374 397 2380 398
rect 2374 393 2375 397
rect 2379 393 2380 397
rect 2374 392 2380 393
rect 2566 397 2572 398
rect 2566 393 2567 397
rect 2571 393 2572 397
rect 2566 392 2572 393
rect 2774 397 2780 398
rect 2774 393 2775 397
rect 2779 393 2780 397
rect 2774 392 2780 393
rect 2998 397 3004 398
rect 2998 393 2999 397
rect 3003 393 3004 397
rect 2998 392 3004 393
rect 3230 397 3236 398
rect 3230 393 3231 397
rect 3235 393 3236 397
rect 3230 392 3236 393
rect 3462 397 3468 398
rect 3462 393 3463 397
rect 3467 393 3468 397
rect 3462 392 3468 393
rect 110 388 116 389
rect 110 384 111 388
rect 115 384 116 388
rect 110 383 116 384
rect 1822 388 1828 389
rect 1822 384 1823 388
rect 1827 384 1828 388
rect 1822 383 1828 384
rect 1886 375 1892 376
rect 110 371 116 372
rect 110 367 111 371
rect 115 367 116 371
rect 110 366 116 367
rect 1822 371 1828 372
rect 1822 367 1823 371
rect 1827 367 1828 371
rect 1886 371 1887 375
rect 1891 371 1892 375
rect 1886 370 1892 371
rect 1974 375 1980 376
rect 1974 371 1975 375
rect 1979 371 1980 375
rect 1974 370 1980 371
rect 2062 375 2068 376
rect 2062 371 2063 375
rect 2067 371 2068 375
rect 2062 370 2068 371
rect 2150 375 2156 376
rect 2150 371 2151 375
rect 2155 371 2156 375
rect 2150 370 2156 371
rect 2262 375 2268 376
rect 2262 371 2263 375
rect 2267 371 2268 375
rect 2262 370 2268 371
rect 2382 375 2388 376
rect 2382 371 2383 375
rect 2387 371 2388 375
rect 2382 370 2388 371
rect 2518 375 2524 376
rect 2518 371 2519 375
rect 2523 371 2524 375
rect 2518 370 2524 371
rect 2670 375 2676 376
rect 2670 371 2671 375
rect 2675 371 2676 375
rect 2670 370 2676 371
rect 2846 375 2852 376
rect 2846 371 2847 375
rect 2851 371 2852 375
rect 2846 370 2852 371
rect 3030 375 3036 376
rect 3030 371 3031 375
rect 3035 371 3036 375
rect 3030 370 3036 371
rect 3230 375 3236 376
rect 3230 371 3231 375
rect 3235 371 3236 375
rect 3230 370 3236 371
rect 3430 375 3436 376
rect 3430 371 3431 375
rect 3435 371 3436 375
rect 3430 370 3436 371
rect 1822 366 1828 367
rect 1862 365 1868 366
rect 142 361 148 362
rect 142 357 143 361
rect 147 357 148 361
rect 142 356 148 357
rect 262 361 268 362
rect 262 357 263 361
rect 267 357 268 361
rect 262 356 268 357
rect 398 361 404 362
rect 398 357 399 361
rect 403 357 404 361
rect 398 356 404 357
rect 542 361 548 362
rect 542 357 543 361
rect 547 357 548 361
rect 542 356 548 357
rect 702 361 708 362
rect 702 357 703 361
rect 707 357 708 361
rect 702 356 708 357
rect 878 361 884 362
rect 878 357 879 361
rect 883 357 884 361
rect 878 356 884 357
rect 1054 361 1060 362
rect 1054 357 1055 361
rect 1059 357 1060 361
rect 1054 356 1060 357
rect 1238 361 1244 362
rect 1238 357 1239 361
rect 1243 357 1244 361
rect 1238 356 1244 357
rect 1430 361 1436 362
rect 1430 357 1431 361
rect 1435 357 1436 361
rect 1430 356 1436 357
rect 1630 361 1636 362
rect 1630 357 1631 361
rect 1635 357 1636 361
rect 1862 361 1863 365
rect 1867 361 1868 365
rect 1862 360 1868 361
rect 3574 365 3580 366
rect 3574 361 3575 365
rect 3579 361 3580 365
rect 3574 360 3580 361
rect 1630 356 1636 357
rect 1862 348 1868 349
rect 1862 344 1863 348
rect 1867 344 1868 348
rect 1862 343 1868 344
rect 3574 348 3580 349
rect 3574 344 3575 348
rect 3579 344 3580 348
rect 3574 343 3580 344
rect 1894 335 1900 336
rect 1894 331 1895 335
rect 1899 331 1900 335
rect 1894 330 1900 331
rect 1982 335 1988 336
rect 1982 331 1983 335
rect 1987 331 1988 335
rect 1982 330 1988 331
rect 2070 335 2076 336
rect 2070 331 2071 335
rect 2075 331 2076 335
rect 2070 330 2076 331
rect 2158 335 2164 336
rect 2158 331 2159 335
rect 2163 331 2164 335
rect 2158 330 2164 331
rect 2270 335 2276 336
rect 2270 331 2271 335
rect 2275 331 2276 335
rect 2270 330 2276 331
rect 2390 335 2396 336
rect 2390 331 2391 335
rect 2395 331 2396 335
rect 2390 330 2396 331
rect 2526 335 2532 336
rect 2526 331 2527 335
rect 2531 331 2532 335
rect 2526 330 2532 331
rect 2678 335 2684 336
rect 2678 331 2679 335
rect 2683 331 2684 335
rect 2678 330 2684 331
rect 2854 335 2860 336
rect 2854 331 2855 335
rect 2859 331 2860 335
rect 2854 330 2860 331
rect 3038 335 3044 336
rect 3038 331 3039 335
rect 3043 331 3044 335
rect 3038 330 3044 331
rect 3238 335 3244 336
rect 3238 331 3239 335
rect 3243 331 3244 335
rect 3238 330 3244 331
rect 3438 335 3444 336
rect 3438 331 3439 335
rect 3443 331 3444 335
rect 3438 330 3444 331
rect 134 323 140 324
rect 134 319 135 323
rect 139 319 140 323
rect 134 318 140 319
rect 222 323 228 324
rect 222 319 223 323
rect 227 319 228 323
rect 222 318 228 319
rect 310 323 316 324
rect 310 319 311 323
rect 315 319 316 323
rect 310 318 316 319
rect 398 323 404 324
rect 398 319 399 323
rect 403 319 404 323
rect 398 318 404 319
rect 486 323 492 324
rect 486 319 487 323
rect 491 319 492 323
rect 486 318 492 319
rect 574 323 580 324
rect 574 319 575 323
rect 579 319 580 323
rect 574 318 580 319
rect 662 323 668 324
rect 662 319 663 323
rect 667 319 668 323
rect 662 318 668 319
rect 750 323 756 324
rect 750 319 751 323
rect 755 319 756 323
rect 750 318 756 319
rect 838 323 844 324
rect 838 319 839 323
rect 843 319 844 323
rect 838 318 844 319
rect 926 323 932 324
rect 926 319 927 323
rect 931 319 932 323
rect 926 318 932 319
rect 1014 323 1020 324
rect 1014 319 1015 323
rect 1019 319 1020 323
rect 1014 318 1020 319
rect 1102 323 1108 324
rect 1102 319 1103 323
rect 1107 319 1108 323
rect 1102 318 1108 319
rect 1190 323 1196 324
rect 1190 319 1191 323
rect 1195 319 1196 323
rect 1190 318 1196 319
rect 1286 323 1292 324
rect 1286 319 1287 323
rect 1291 319 1292 323
rect 1286 318 1292 319
rect 1382 323 1388 324
rect 1382 319 1383 323
rect 1387 319 1388 323
rect 1382 318 1388 319
rect 1478 323 1484 324
rect 1478 319 1479 323
rect 1483 319 1484 323
rect 1478 318 1484 319
rect 1574 323 1580 324
rect 1574 319 1575 323
rect 1579 319 1580 323
rect 1574 318 1580 319
rect 1670 323 1676 324
rect 1670 319 1671 323
rect 1675 319 1676 323
rect 1670 318 1676 319
rect 110 313 116 314
rect 110 309 111 313
rect 115 309 116 313
rect 110 308 116 309
rect 1822 313 1828 314
rect 1822 309 1823 313
rect 1827 309 1828 313
rect 1822 308 1828 309
rect 1894 301 1900 302
rect 1894 297 1895 301
rect 1899 297 1900 301
rect 110 296 116 297
rect 110 292 111 296
rect 115 292 116 296
rect 110 291 116 292
rect 1822 296 1828 297
rect 1894 296 1900 297
rect 1982 301 1988 302
rect 1982 297 1983 301
rect 1987 297 1988 301
rect 1982 296 1988 297
rect 2070 301 2076 302
rect 2070 297 2071 301
rect 2075 297 2076 301
rect 2070 296 2076 297
rect 2158 301 2164 302
rect 2158 297 2159 301
rect 2163 297 2164 301
rect 2158 296 2164 297
rect 2246 301 2252 302
rect 2246 297 2247 301
rect 2251 297 2252 301
rect 2246 296 2252 297
rect 2358 301 2364 302
rect 2358 297 2359 301
rect 2363 297 2364 301
rect 2358 296 2364 297
rect 2470 301 2476 302
rect 2470 297 2471 301
rect 2475 297 2476 301
rect 2470 296 2476 297
rect 2582 301 2588 302
rect 2582 297 2583 301
rect 2587 297 2588 301
rect 2582 296 2588 297
rect 2694 301 2700 302
rect 2694 297 2695 301
rect 2699 297 2700 301
rect 2694 296 2700 297
rect 2806 301 2812 302
rect 2806 297 2807 301
rect 2811 297 2812 301
rect 2806 296 2812 297
rect 2918 301 2924 302
rect 2918 297 2919 301
rect 2923 297 2924 301
rect 2918 296 2924 297
rect 3038 301 3044 302
rect 3038 297 3039 301
rect 3043 297 3044 301
rect 3038 296 3044 297
rect 3158 301 3164 302
rect 3158 297 3159 301
rect 3163 297 3164 301
rect 3158 296 3164 297
rect 1822 292 1823 296
rect 1827 292 1828 296
rect 1822 291 1828 292
rect 1862 288 1868 289
rect 1862 284 1863 288
rect 1867 284 1868 288
rect 142 283 148 284
rect 142 279 143 283
rect 147 279 148 283
rect 142 278 148 279
rect 230 283 236 284
rect 230 279 231 283
rect 235 279 236 283
rect 230 278 236 279
rect 318 283 324 284
rect 318 279 319 283
rect 323 279 324 283
rect 318 278 324 279
rect 406 283 412 284
rect 406 279 407 283
rect 411 279 412 283
rect 406 278 412 279
rect 494 283 500 284
rect 494 279 495 283
rect 499 279 500 283
rect 494 278 500 279
rect 582 283 588 284
rect 582 279 583 283
rect 587 279 588 283
rect 582 278 588 279
rect 670 283 676 284
rect 670 279 671 283
rect 675 279 676 283
rect 670 278 676 279
rect 758 283 764 284
rect 758 279 759 283
rect 763 279 764 283
rect 758 278 764 279
rect 846 283 852 284
rect 846 279 847 283
rect 851 279 852 283
rect 846 278 852 279
rect 934 283 940 284
rect 934 279 935 283
rect 939 279 940 283
rect 934 278 940 279
rect 1022 283 1028 284
rect 1022 279 1023 283
rect 1027 279 1028 283
rect 1022 278 1028 279
rect 1110 283 1116 284
rect 1110 279 1111 283
rect 1115 279 1116 283
rect 1110 278 1116 279
rect 1198 283 1204 284
rect 1198 279 1199 283
rect 1203 279 1204 283
rect 1198 278 1204 279
rect 1294 283 1300 284
rect 1294 279 1295 283
rect 1299 279 1300 283
rect 1294 278 1300 279
rect 1390 283 1396 284
rect 1390 279 1391 283
rect 1395 279 1396 283
rect 1390 278 1396 279
rect 1486 283 1492 284
rect 1486 279 1487 283
rect 1491 279 1492 283
rect 1486 278 1492 279
rect 1582 283 1588 284
rect 1582 279 1583 283
rect 1587 279 1588 283
rect 1582 278 1588 279
rect 1678 283 1684 284
rect 1862 283 1868 284
rect 3574 288 3580 289
rect 3574 284 3575 288
rect 3579 284 3580 288
rect 3574 283 3580 284
rect 1678 279 1679 283
rect 1683 279 1684 283
rect 1678 278 1684 279
rect 1862 271 1868 272
rect 1862 267 1863 271
rect 1867 267 1868 271
rect 1862 266 1868 267
rect 3574 271 3580 272
rect 3574 267 3575 271
rect 3579 267 3580 271
rect 3574 266 3580 267
rect 1886 261 1892 262
rect 1886 257 1887 261
rect 1891 257 1892 261
rect 1886 256 1892 257
rect 1974 261 1980 262
rect 1974 257 1975 261
rect 1979 257 1980 261
rect 1974 256 1980 257
rect 2062 261 2068 262
rect 2062 257 2063 261
rect 2067 257 2068 261
rect 2062 256 2068 257
rect 2150 261 2156 262
rect 2150 257 2151 261
rect 2155 257 2156 261
rect 2150 256 2156 257
rect 2238 261 2244 262
rect 2238 257 2239 261
rect 2243 257 2244 261
rect 2238 256 2244 257
rect 2350 261 2356 262
rect 2350 257 2351 261
rect 2355 257 2356 261
rect 2350 256 2356 257
rect 2462 261 2468 262
rect 2462 257 2463 261
rect 2467 257 2468 261
rect 2462 256 2468 257
rect 2574 261 2580 262
rect 2574 257 2575 261
rect 2579 257 2580 261
rect 2574 256 2580 257
rect 2686 261 2692 262
rect 2686 257 2687 261
rect 2691 257 2692 261
rect 2686 256 2692 257
rect 2798 261 2804 262
rect 2798 257 2799 261
rect 2803 257 2804 261
rect 2798 256 2804 257
rect 2910 261 2916 262
rect 2910 257 2911 261
rect 2915 257 2916 261
rect 2910 256 2916 257
rect 3030 261 3036 262
rect 3030 257 3031 261
rect 3035 257 3036 261
rect 3030 256 3036 257
rect 3150 261 3156 262
rect 3150 257 3151 261
rect 3155 257 3156 261
rect 3150 256 3156 257
rect 142 245 148 246
rect 142 241 143 245
rect 147 241 148 245
rect 142 240 148 241
rect 230 245 236 246
rect 230 241 231 245
rect 235 241 236 245
rect 230 240 236 241
rect 318 245 324 246
rect 318 241 319 245
rect 323 241 324 245
rect 318 240 324 241
rect 406 245 412 246
rect 406 241 407 245
rect 411 241 412 245
rect 406 240 412 241
rect 494 245 500 246
rect 494 241 495 245
rect 499 241 500 245
rect 494 240 500 241
rect 582 245 588 246
rect 582 241 583 245
rect 587 241 588 245
rect 582 240 588 241
rect 670 245 676 246
rect 670 241 671 245
rect 675 241 676 245
rect 670 240 676 241
rect 758 245 764 246
rect 758 241 759 245
rect 763 241 764 245
rect 758 240 764 241
rect 846 245 852 246
rect 846 241 847 245
rect 851 241 852 245
rect 846 240 852 241
rect 934 245 940 246
rect 934 241 935 245
rect 939 241 940 245
rect 934 240 940 241
rect 1022 245 1028 246
rect 1022 241 1023 245
rect 1027 241 1028 245
rect 1022 240 1028 241
rect 1110 245 1116 246
rect 1110 241 1111 245
rect 1115 241 1116 245
rect 1110 240 1116 241
rect 1198 245 1204 246
rect 1198 241 1199 245
rect 1203 241 1204 245
rect 1198 240 1204 241
rect 1286 245 1292 246
rect 1286 241 1287 245
rect 1291 241 1292 245
rect 1286 240 1292 241
rect 1374 245 1380 246
rect 1374 241 1375 245
rect 1379 241 1380 245
rect 1374 240 1380 241
rect 1462 245 1468 246
rect 1462 241 1463 245
rect 1467 241 1468 245
rect 1462 240 1468 241
rect 1550 245 1556 246
rect 1550 241 1551 245
rect 1555 241 1556 245
rect 1550 240 1556 241
rect 1638 245 1644 246
rect 1638 241 1639 245
rect 1643 241 1644 245
rect 1638 240 1644 241
rect 1726 245 1732 246
rect 1726 241 1727 245
rect 1731 241 1732 245
rect 1726 240 1732 241
rect 1886 239 1892 240
rect 1886 235 1887 239
rect 1891 235 1892 239
rect 1886 234 1892 235
rect 1974 239 1980 240
rect 1974 235 1975 239
rect 1979 235 1980 239
rect 1974 234 1980 235
rect 2062 239 2068 240
rect 2062 235 2063 239
rect 2067 235 2068 239
rect 2062 234 2068 235
rect 2150 239 2156 240
rect 2150 235 2151 239
rect 2155 235 2156 239
rect 2150 234 2156 235
rect 2262 239 2268 240
rect 2262 235 2263 239
rect 2267 235 2268 239
rect 2262 234 2268 235
rect 2398 239 2404 240
rect 2398 235 2399 239
rect 2403 235 2404 239
rect 2398 234 2404 235
rect 2534 239 2540 240
rect 2534 235 2535 239
rect 2539 235 2540 239
rect 2534 234 2540 235
rect 2678 239 2684 240
rect 2678 235 2679 239
rect 2683 235 2684 239
rect 2678 234 2684 235
rect 2814 239 2820 240
rect 2814 235 2815 239
rect 2819 235 2820 239
rect 2814 234 2820 235
rect 2950 239 2956 240
rect 2950 235 2951 239
rect 2955 235 2956 239
rect 2950 234 2956 235
rect 3086 239 3092 240
rect 3086 235 3087 239
rect 3091 235 3092 239
rect 3086 234 3092 235
rect 3222 239 3228 240
rect 3222 235 3223 239
rect 3227 235 3228 239
rect 3222 234 3228 235
rect 3358 239 3364 240
rect 3358 235 3359 239
rect 3363 235 3364 239
rect 3358 234 3364 235
rect 3478 239 3484 240
rect 3478 235 3479 239
rect 3483 235 3484 239
rect 3478 234 3484 235
rect 110 232 116 233
rect 110 228 111 232
rect 115 228 116 232
rect 110 227 116 228
rect 1822 232 1828 233
rect 1822 228 1823 232
rect 1827 228 1828 232
rect 1822 227 1828 228
rect 1862 229 1868 230
rect 1862 225 1863 229
rect 1867 225 1868 229
rect 1862 224 1868 225
rect 3574 229 3580 230
rect 3574 225 3575 229
rect 3579 225 3580 229
rect 3574 224 3580 225
rect 110 215 116 216
rect 110 211 111 215
rect 115 211 116 215
rect 110 210 116 211
rect 1822 215 1828 216
rect 1822 211 1823 215
rect 1827 211 1828 215
rect 1822 210 1828 211
rect 1862 212 1868 213
rect 1862 208 1863 212
rect 1867 208 1868 212
rect 1862 207 1868 208
rect 3574 212 3580 213
rect 3574 208 3575 212
rect 3579 208 3580 212
rect 3574 207 3580 208
rect 134 205 140 206
rect 134 201 135 205
rect 139 201 140 205
rect 134 200 140 201
rect 222 205 228 206
rect 222 201 223 205
rect 227 201 228 205
rect 222 200 228 201
rect 310 205 316 206
rect 310 201 311 205
rect 315 201 316 205
rect 310 200 316 201
rect 398 205 404 206
rect 398 201 399 205
rect 403 201 404 205
rect 398 200 404 201
rect 486 205 492 206
rect 486 201 487 205
rect 491 201 492 205
rect 486 200 492 201
rect 574 205 580 206
rect 574 201 575 205
rect 579 201 580 205
rect 574 200 580 201
rect 662 205 668 206
rect 662 201 663 205
rect 667 201 668 205
rect 662 200 668 201
rect 750 205 756 206
rect 750 201 751 205
rect 755 201 756 205
rect 750 200 756 201
rect 838 205 844 206
rect 838 201 839 205
rect 843 201 844 205
rect 838 200 844 201
rect 926 205 932 206
rect 926 201 927 205
rect 931 201 932 205
rect 926 200 932 201
rect 1014 205 1020 206
rect 1014 201 1015 205
rect 1019 201 1020 205
rect 1014 200 1020 201
rect 1102 205 1108 206
rect 1102 201 1103 205
rect 1107 201 1108 205
rect 1102 200 1108 201
rect 1190 205 1196 206
rect 1190 201 1191 205
rect 1195 201 1196 205
rect 1190 200 1196 201
rect 1278 205 1284 206
rect 1278 201 1279 205
rect 1283 201 1284 205
rect 1278 200 1284 201
rect 1366 205 1372 206
rect 1366 201 1367 205
rect 1371 201 1372 205
rect 1366 200 1372 201
rect 1454 205 1460 206
rect 1454 201 1455 205
rect 1459 201 1460 205
rect 1454 200 1460 201
rect 1542 205 1548 206
rect 1542 201 1543 205
rect 1547 201 1548 205
rect 1542 200 1548 201
rect 1630 205 1636 206
rect 1630 201 1631 205
rect 1635 201 1636 205
rect 1630 200 1636 201
rect 1718 205 1724 206
rect 1718 201 1719 205
rect 1723 201 1724 205
rect 1718 200 1724 201
rect 1894 199 1900 200
rect 1894 195 1895 199
rect 1899 195 1900 199
rect 1894 194 1900 195
rect 1982 199 1988 200
rect 1982 195 1983 199
rect 1987 195 1988 199
rect 1982 194 1988 195
rect 2070 199 2076 200
rect 2070 195 2071 199
rect 2075 195 2076 199
rect 2070 194 2076 195
rect 2158 199 2164 200
rect 2158 195 2159 199
rect 2163 195 2164 199
rect 2158 194 2164 195
rect 2270 199 2276 200
rect 2270 195 2271 199
rect 2275 195 2276 199
rect 2270 194 2276 195
rect 2406 199 2412 200
rect 2406 195 2407 199
rect 2411 195 2412 199
rect 2406 194 2412 195
rect 2542 199 2548 200
rect 2542 195 2543 199
rect 2547 195 2548 199
rect 2542 194 2548 195
rect 2686 199 2692 200
rect 2686 195 2687 199
rect 2691 195 2692 199
rect 2686 194 2692 195
rect 2822 199 2828 200
rect 2822 195 2823 199
rect 2827 195 2828 199
rect 2822 194 2828 195
rect 2958 199 2964 200
rect 2958 195 2959 199
rect 2963 195 2964 199
rect 2958 194 2964 195
rect 3094 199 3100 200
rect 3094 195 3095 199
rect 3099 195 3100 199
rect 3094 194 3100 195
rect 3230 199 3236 200
rect 3230 195 3231 199
rect 3235 195 3236 199
rect 3230 194 3236 195
rect 3366 199 3372 200
rect 3366 195 3367 199
rect 3371 195 3372 199
rect 3366 194 3372 195
rect 3486 199 3492 200
rect 3486 195 3487 199
rect 3491 195 3492 199
rect 3486 194 3492 195
rect 2782 133 2788 134
rect 2782 129 2783 133
rect 2787 129 2788 133
rect 2782 128 2788 129
rect 2870 133 2876 134
rect 2870 129 2871 133
rect 2875 129 2876 133
rect 2870 128 2876 129
rect 2958 133 2964 134
rect 2958 129 2959 133
rect 2963 129 2964 133
rect 2958 128 2964 129
rect 3046 133 3052 134
rect 3046 129 3047 133
rect 3051 129 3052 133
rect 3046 128 3052 129
rect 3134 133 3140 134
rect 3134 129 3135 133
rect 3139 129 3140 133
rect 3134 128 3140 129
rect 3222 133 3228 134
rect 3222 129 3223 133
rect 3227 129 3228 133
rect 3222 128 3228 129
rect 3310 133 3316 134
rect 3310 129 3311 133
rect 3315 129 3316 133
rect 3310 128 3316 129
rect 3398 133 3404 134
rect 3398 129 3399 133
rect 3403 129 3404 133
rect 3398 128 3404 129
rect 3486 133 3492 134
rect 3486 129 3487 133
rect 3491 129 3492 133
rect 3486 128 3492 129
rect 1862 120 1868 121
rect 1862 116 1863 120
rect 1867 116 1868 120
rect 1862 115 1868 116
rect 3574 120 3580 121
rect 3574 116 3575 120
rect 3579 116 3580 120
rect 3574 115 3580 116
rect 1862 103 1868 104
rect 1862 99 1863 103
rect 1867 99 1868 103
rect 1862 98 1868 99
rect 3574 103 3580 104
rect 3574 99 3575 103
rect 3579 99 3580 103
rect 3574 98 3580 99
rect 2774 93 2780 94
rect 2774 89 2775 93
rect 2779 89 2780 93
rect 2774 88 2780 89
rect 2862 93 2868 94
rect 2862 89 2863 93
rect 2867 89 2868 93
rect 2862 88 2868 89
rect 2950 93 2956 94
rect 2950 89 2951 93
rect 2955 89 2956 93
rect 2950 88 2956 89
rect 3038 93 3044 94
rect 3038 89 3039 93
rect 3043 89 3044 93
rect 3038 88 3044 89
rect 3126 93 3132 94
rect 3126 89 3127 93
rect 3131 89 3132 93
rect 3126 88 3132 89
rect 3214 93 3220 94
rect 3214 89 3215 93
rect 3219 89 3220 93
rect 3214 88 3220 89
rect 3302 93 3308 94
rect 3302 89 3303 93
rect 3307 89 3308 93
rect 3302 88 3308 89
rect 3390 93 3396 94
rect 3390 89 3391 93
rect 3395 89 3396 93
rect 3390 88 3396 89
rect 3478 93 3484 94
rect 3478 89 3479 93
rect 3483 89 3484 93
rect 3478 88 3484 89
<< m3c >>
rect 135 3655 139 3659
rect 223 3655 227 3659
rect 111 3645 115 3649
rect 1823 3645 1827 3649
rect 111 3628 115 3632
rect 1823 3628 1827 3632
rect 143 3615 147 3619
rect 231 3615 235 3619
rect 143 3581 147 3585
rect 231 3581 235 3585
rect 319 3581 323 3585
rect 407 3581 411 3585
rect 495 3581 499 3585
rect 1887 3579 1891 3583
rect 1975 3579 1979 3583
rect 2063 3579 2067 3583
rect 2151 3579 2155 3583
rect 2239 3579 2243 3583
rect 2327 3579 2331 3583
rect 2431 3579 2435 3583
rect 2535 3579 2539 3583
rect 2631 3579 2635 3583
rect 2727 3579 2731 3583
rect 2823 3579 2827 3583
rect 2919 3579 2923 3583
rect 3015 3579 3019 3583
rect 3119 3579 3123 3583
rect 3223 3579 3227 3583
rect 111 3568 115 3572
rect 1823 3568 1827 3572
rect 1863 3569 1867 3573
rect 3575 3569 3579 3573
rect 111 3551 115 3555
rect 1823 3551 1827 3555
rect 1863 3552 1867 3556
rect 3575 3552 3579 3556
rect 135 3541 139 3545
rect 223 3541 227 3545
rect 311 3541 315 3545
rect 399 3541 403 3545
rect 487 3541 491 3545
rect 1895 3539 1899 3543
rect 1983 3539 1987 3543
rect 2071 3539 2075 3543
rect 2159 3539 2163 3543
rect 2247 3539 2251 3543
rect 2335 3539 2339 3543
rect 2439 3539 2443 3543
rect 2543 3539 2547 3543
rect 2639 3539 2643 3543
rect 2735 3539 2739 3543
rect 2831 3539 2835 3543
rect 2927 3539 2931 3543
rect 3023 3539 3027 3543
rect 3127 3539 3131 3543
rect 3231 3539 3235 3543
rect 247 3519 251 3523
rect 375 3519 379 3523
rect 503 3519 507 3523
rect 623 3519 627 3523
rect 743 3519 747 3523
rect 863 3519 867 3523
rect 975 3519 979 3523
rect 1079 3519 1083 3523
rect 1175 3519 1179 3523
rect 1271 3519 1275 3523
rect 1367 3519 1371 3523
rect 1471 3519 1475 3523
rect 1575 3519 1579 3523
rect 111 3509 115 3513
rect 1823 3509 1827 3513
rect 1895 3505 1899 3509
rect 1983 3505 1987 3509
rect 2103 3505 2107 3509
rect 2231 3505 2235 3509
rect 2367 3505 2371 3509
rect 2511 3505 2515 3509
rect 2655 3505 2659 3509
rect 2791 3505 2795 3509
rect 2935 3505 2939 3509
rect 3079 3505 3083 3509
rect 3223 3505 3227 3509
rect 111 3492 115 3496
rect 1823 3492 1827 3496
rect 1863 3492 1867 3496
rect 3575 3492 3579 3496
rect 255 3479 259 3483
rect 383 3479 387 3483
rect 511 3479 515 3483
rect 631 3479 635 3483
rect 751 3479 755 3483
rect 871 3479 875 3483
rect 983 3479 987 3483
rect 1087 3479 1091 3483
rect 1183 3479 1187 3483
rect 1279 3479 1283 3483
rect 1375 3479 1379 3483
rect 1479 3479 1483 3483
rect 1583 3479 1587 3483
rect 1863 3475 1867 3479
rect 3575 3475 3579 3479
rect 1887 3465 1891 3469
rect 1975 3465 1979 3469
rect 2095 3465 2099 3469
rect 2223 3465 2227 3469
rect 2359 3465 2363 3469
rect 2503 3465 2507 3469
rect 2647 3465 2651 3469
rect 2783 3465 2787 3469
rect 2927 3465 2931 3469
rect 3071 3465 3075 3469
rect 3215 3465 3219 3469
rect 175 3445 179 3449
rect 303 3445 307 3449
rect 447 3445 451 3449
rect 591 3445 595 3449
rect 743 3445 747 3449
rect 895 3445 899 3449
rect 1039 3445 1043 3449
rect 1183 3445 1187 3449
rect 1327 3445 1331 3449
rect 1479 3445 1483 3449
rect 111 3432 115 3436
rect 1823 3432 1827 3436
rect 1887 3435 1891 3439
rect 2023 3435 2027 3439
rect 2191 3435 2195 3439
rect 2367 3435 2371 3439
rect 2543 3435 2547 3439
rect 2711 3435 2715 3439
rect 2871 3435 2875 3439
rect 3031 3435 3035 3439
rect 3191 3435 3195 3439
rect 3359 3435 3363 3439
rect 1863 3425 1867 3429
rect 3575 3425 3579 3429
rect 111 3415 115 3419
rect 1823 3415 1827 3419
rect 167 3405 171 3409
rect 295 3405 299 3409
rect 439 3405 443 3409
rect 583 3405 587 3409
rect 735 3405 739 3409
rect 887 3405 891 3409
rect 1031 3405 1035 3409
rect 1175 3405 1179 3409
rect 1319 3405 1323 3409
rect 1471 3405 1475 3409
rect 1863 3408 1867 3412
rect 3575 3408 3579 3412
rect 1895 3395 1899 3399
rect 2031 3395 2035 3399
rect 2199 3395 2203 3399
rect 2375 3395 2379 3399
rect 2551 3395 2555 3399
rect 2719 3395 2723 3399
rect 2879 3395 2883 3399
rect 3039 3395 3043 3399
rect 3199 3395 3203 3399
rect 3367 3395 3371 3399
rect 135 3383 139 3387
rect 263 3383 267 3387
rect 407 3383 411 3387
rect 567 3383 571 3387
rect 727 3383 731 3387
rect 887 3383 891 3387
rect 1047 3383 1051 3387
rect 1207 3383 1211 3387
rect 1367 3383 1371 3387
rect 1527 3383 1531 3387
rect 111 3373 115 3377
rect 1823 3373 1827 3377
rect 111 3356 115 3360
rect 1823 3356 1827 3360
rect 1895 3353 1899 3357
rect 2031 3353 2035 3357
rect 2199 3353 2203 3357
rect 2375 3353 2379 3357
rect 2551 3353 2555 3357
rect 2719 3353 2723 3357
rect 2879 3353 2883 3357
rect 3039 3353 3043 3357
rect 3191 3353 3195 3357
rect 3343 3353 3347 3357
rect 3487 3353 3491 3357
rect 143 3343 147 3347
rect 271 3343 275 3347
rect 415 3343 419 3347
rect 575 3343 579 3347
rect 735 3343 739 3347
rect 895 3343 899 3347
rect 1055 3343 1059 3347
rect 1215 3343 1219 3347
rect 1375 3343 1379 3347
rect 1535 3343 1539 3347
rect 1863 3340 1867 3344
rect 3575 3340 3579 3344
rect 1863 3323 1867 3327
rect 3575 3323 3579 3327
rect 1887 3313 1891 3317
rect 2023 3313 2027 3317
rect 2191 3313 2195 3317
rect 2367 3313 2371 3317
rect 2543 3313 2547 3317
rect 2711 3313 2715 3317
rect 2871 3313 2875 3317
rect 3031 3313 3035 3317
rect 3183 3313 3187 3317
rect 3335 3313 3339 3317
rect 3479 3313 3483 3317
rect 207 3305 211 3309
rect 335 3305 339 3309
rect 479 3305 483 3309
rect 639 3305 643 3309
rect 807 3305 811 3309
rect 983 3305 987 3309
rect 1167 3305 1171 3309
rect 1351 3305 1355 3309
rect 1543 3305 1547 3309
rect 111 3292 115 3296
rect 1823 3292 1827 3296
rect 1887 3291 1891 3295
rect 2007 3291 2011 3295
rect 2151 3291 2155 3295
rect 2303 3291 2307 3295
rect 2463 3291 2467 3295
rect 2631 3291 2635 3295
rect 2799 3291 2803 3295
rect 2967 3291 2971 3295
rect 3135 3291 3139 3295
rect 3311 3291 3315 3295
rect 3479 3291 3483 3295
rect 1863 3281 1867 3285
rect 3575 3281 3579 3285
rect 111 3275 115 3279
rect 1823 3275 1827 3279
rect 199 3265 203 3269
rect 327 3265 331 3269
rect 471 3265 475 3269
rect 631 3265 635 3269
rect 799 3265 803 3269
rect 975 3265 979 3269
rect 1159 3265 1163 3269
rect 1343 3265 1347 3269
rect 1535 3265 1539 3269
rect 1863 3264 1867 3268
rect 3575 3264 3579 3268
rect 1895 3251 1899 3255
rect 2015 3251 2019 3255
rect 2159 3251 2163 3255
rect 2311 3251 2315 3255
rect 2471 3251 2475 3255
rect 2639 3251 2643 3255
rect 2807 3251 2811 3255
rect 2975 3251 2979 3255
rect 3143 3251 3147 3255
rect 3319 3251 3323 3255
rect 3487 3251 3491 3255
rect 367 3239 371 3243
rect 503 3239 507 3243
rect 639 3239 643 3243
rect 783 3239 787 3243
rect 935 3239 939 3243
rect 1095 3239 1099 3243
rect 1255 3239 1259 3243
rect 1415 3239 1419 3243
rect 1575 3239 1579 3243
rect 111 3229 115 3233
rect 1823 3229 1827 3233
rect 111 3212 115 3216
rect 1823 3212 1827 3216
rect 1895 3209 1899 3213
rect 2023 3209 2027 3213
rect 2175 3209 2179 3213
rect 2327 3209 2331 3213
rect 2463 3209 2467 3213
rect 2599 3209 2603 3213
rect 2735 3209 2739 3213
rect 2871 3209 2875 3213
rect 3015 3209 3019 3213
rect 3167 3209 3171 3213
rect 3327 3209 3331 3213
rect 3487 3209 3491 3213
rect 375 3199 379 3203
rect 511 3199 515 3203
rect 647 3199 651 3203
rect 791 3199 795 3203
rect 943 3199 947 3203
rect 1103 3199 1107 3203
rect 1263 3199 1267 3203
rect 1423 3199 1427 3203
rect 1583 3199 1587 3203
rect 1863 3196 1867 3200
rect 3575 3196 3579 3200
rect 1863 3179 1867 3183
rect 3575 3179 3579 3183
rect 1887 3169 1891 3173
rect 2015 3169 2019 3173
rect 2167 3169 2171 3173
rect 2319 3169 2323 3173
rect 2455 3169 2459 3173
rect 2591 3169 2595 3173
rect 2727 3169 2731 3173
rect 2863 3169 2867 3173
rect 3007 3169 3011 3173
rect 3159 3169 3163 3173
rect 3319 3169 3323 3173
rect 3479 3169 3483 3173
rect 447 3157 451 3161
rect 559 3157 563 3161
rect 687 3157 691 3161
rect 823 3157 827 3161
rect 975 3157 979 3161
rect 1135 3157 1139 3161
rect 1295 3157 1299 3161
rect 1463 3157 1467 3161
rect 1639 3157 1643 3161
rect 111 3144 115 3148
rect 1823 3144 1827 3148
rect 1887 3143 1891 3147
rect 2047 3143 2051 3147
rect 2199 3143 2203 3147
rect 2351 3143 2355 3147
rect 2511 3143 2515 3147
rect 2679 3143 2683 3147
rect 2871 3143 2875 3147
rect 3071 3143 3075 3147
rect 3287 3143 3291 3147
rect 3479 3143 3483 3147
rect 1863 3133 1867 3137
rect 3575 3133 3579 3137
rect 111 3127 115 3131
rect 1823 3127 1827 3131
rect 439 3117 443 3121
rect 551 3117 555 3121
rect 679 3117 683 3121
rect 815 3117 819 3121
rect 967 3117 971 3121
rect 1127 3117 1131 3121
rect 1287 3117 1291 3121
rect 1455 3117 1459 3121
rect 1631 3117 1635 3121
rect 1863 3116 1867 3120
rect 3575 3116 3579 3120
rect 1895 3103 1899 3107
rect 2055 3103 2059 3107
rect 2207 3103 2211 3107
rect 2359 3103 2363 3107
rect 2519 3103 2523 3107
rect 2687 3103 2691 3107
rect 2879 3103 2883 3107
rect 3079 3103 3083 3107
rect 3295 3103 3299 3107
rect 3487 3103 3491 3107
rect 551 3087 555 3091
rect 663 3087 667 3091
rect 783 3087 787 3091
rect 903 3087 907 3091
rect 1031 3087 1035 3091
rect 1159 3087 1163 3091
rect 1287 3087 1291 3091
rect 1423 3087 1427 3091
rect 1559 3087 1563 3091
rect 1695 3087 1699 3091
rect 111 3077 115 3081
rect 1823 3077 1827 3081
rect 111 3060 115 3064
rect 1823 3060 1827 3064
rect 1919 3061 1923 3065
rect 2087 3061 2091 3065
rect 2279 3061 2283 3065
rect 2487 3061 2491 3065
rect 2719 3061 2723 3065
rect 2975 3061 2979 3065
rect 3239 3061 3243 3065
rect 3487 3061 3491 3065
rect 559 3047 563 3051
rect 671 3047 675 3051
rect 791 3047 795 3051
rect 911 3047 915 3051
rect 1039 3047 1043 3051
rect 1167 3047 1171 3051
rect 1295 3047 1299 3051
rect 1431 3047 1435 3051
rect 1567 3047 1571 3051
rect 1703 3047 1707 3051
rect 1863 3048 1867 3052
rect 3575 3048 3579 3052
rect 1863 3031 1867 3035
rect 3575 3031 3579 3035
rect 1911 3021 1915 3025
rect 2079 3021 2083 3025
rect 2271 3021 2275 3025
rect 2479 3021 2483 3025
rect 2711 3021 2715 3025
rect 2967 3021 2971 3025
rect 3231 3021 3235 3025
rect 3479 3021 3483 3025
rect 575 3009 579 3013
rect 703 3009 707 3013
rect 831 3009 835 3013
rect 967 3009 971 3013
rect 1103 3009 1107 3013
rect 1239 3009 1243 3013
rect 1367 3009 1371 3013
rect 1495 3009 1499 3013
rect 1623 3009 1627 3013
rect 1735 3009 1739 3013
rect 111 2996 115 3000
rect 1823 2996 1827 3000
rect 2023 2995 2027 2999
rect 2159 2995 2163 2999
rect 2287 2995 2291 2999
rect 2415 2995 2419 2999
rect 2535 2995 2539 2999
rect 2663 2995 2667 2999
rect 2807 2995 2811 2999
rect 2967 2995 2971 2999
rect 3143 2995 3147 2999
rect 3319 2995 3323 2999
rect 3479 2995 3483 2999
rect 1863 2985 1867 2989
rect 3575 2985 3579 2989
rect 111 2979 115 2983
rect 1823 2979 1827 2983
rect 567 2969 571 2973
rect 695 2969 699 2973
rect 823 2969 827 2973
rect 959 2969 963 2973
rect 1095 2969 1099 2973
rect 1231 2969 1235 2973
rect 1359 2969 1363 2973
rect 1487 2969 1491 2973
rect 1615 2969 1619 2973
rect 1727 2969 1731 2973
rect 1863 2968 1867 2972
rect 3575 2968 3579 2972
rect 2031 2955 2035 2959
rect 2167 2955 2171 2959
rect 2295 2955 2299 2959
rect 2423 2955 2427 2959
rect 2543 2955 2547 2959
rect 2671 2955 2675 2959
rect 2815 2955 2819 2959
rect 2975 2955 2979 2959
rect 3151 2955 3155 2959
rect 3327 2955 3331 2959
rect 3487 2955 3491 2959
rect 495 2947 499 2951
rect 639 2947 643 2951
rect 783 2947 787 2951
rect 919 2947 923 2951
rect 1055 2947 1059 2951
rect 1183 2947 1187 2951
rect 1303 2947 1307 2951
rect 1415 2947 1419 2951
rect 1527 2947 1531 2951
rect 1639 2947 1643 2951
rect 1727 2947 1731 2951
rect 111 2937 115 2941
rect 1823 2937 1827 2941
rect 111 2920 115 2924
rect 1823 2920 1827 2924
rect 1895 2913 1899 2917
rect 2175 2913 2179 2917
rect 2495 2913 2499 2917
rect 2823 2913 2827 2917
rect 3167 2913 3171 2917
rect 3487 2913 3491 2917
rect 503 2907 507 2911
rect 647 2907 651 2911
rect 791 2907 795 2911
rect 927 2907 931 2911
rect 1063 2907 1067 2911
rect 1191 2907 1195 2911
rect 1311 2907 1315 2911
rect 1423 2907 1427 2911
rect 1535 2907 1539 2911
rect 1647 2907 1651 2911
rect 1735 2907 1739 2911
rect 1863 2900 1867 2904
rect 3575 2900 3579 2904
rect 1863 2883 1867 2887
rect 3575 2883 3579 2887
rect 327 2869 331 2873
rect 455 2869 459 2873
rect 591 2869 595 2873
rect 727 2869 731 2873
rect 871 2869 875 2873
rect 1007 2869 1011 2873
rect 1143 2869 1147 2873
rect 1279 2869 1283 2873
rect 1415 2869 1419 2873
rect 1551 2869 1555 2873
rect 1887 2873 1891 2877
rect 2167 2873 2171 2877
rect 2487 2873 2491 2877
rect 2815 2873 2819 2877
rect 3159 2873 3163 2877
rect 3479 2873 3483 2877
rect 111 2856 115 2860
rect 1823 2856 1827 2860
rect 1887 2851 1891 2855
rect 2023 2851 2027 2855
rect 2191 2851 2195 2855
rect 2359 2851 2363 2855
rect 2519 2851 2523 2855
rect 2671 2851 2675 2855
rect 2807 2851 2811 2855
rect 2935 2851 2939 2855
rect 3055 2851 3059 2855
rect 3167 2851 3171 2855
rect 3279 2851 3283 2855
rect 3391 2851 3395 2855
rect 3479 2851 3483 2855
rect 111 2839 115 2843
rect 1823 2839 1827 2843
rect 1863 2841 1867 2845
rect 3575 2841 3579 2845
rect 319 2829 323 2833
rect 447 2829 451 2833
rect 583 2829 587 2833
rect 719 2829 723 2833
rect 863 2829 867 2833
rect 999 2829 1003 2833
rect 1135 2829 1139 2833
rect 1271 2829 1275 2833
rect 1407 2829 1411 2833
rect 1543 2829 1547 2833
rect 1863 2824 1867 2828
rect 3575 2824 3579 2828
rect 1895 2811 1899 2815
rect 2031 2811 2035 2815
rect 2199 2811 2203 2815
rect 2367 2811 2371 2815
rect 2527 2811 2531 2815
rect 2679 2811 2683 2815
rect 2815 2811 2819 2815
rect 2943 2811 2947 2815
rect 3063 2811 3067 2815
rect 3175 2811 3179 2815
rect 3287 2811 3291 2815
rect 3399 2811 3403 2815
rect 3487 2811 3491 2815
rect 167 2799 171 2803
rect 295 2799 299 2803
rect 423 2799 427 2803
rect 559 2799 563 2803
rect 695 2799 699 2803
rect 823 2799 827 2803
rect 951 2799 955 2803
rect 1079 2799 1083 2803
rect 1207 2799 1211 2803
rect 1343 2799 1347 2803
rect 111 2789 115 2793
rect 1823 2789 1827 2793
rect 1895 2777 1899 2781
rect 111 2772 115 2776
rect 2063 2777 2067 2781
rect 2255 2777 2259 2781
rect 2439 2777 2443 2781
rect 2615 2777 2619 2781
rect 2783 2777 2787 2781
rect 2935 2777 2939 2781
rect 3079 2777 3083 2781
rect 3223 2777 3227 2781
rect 3367 2777 3371 2781
rect 3487 2777 3491 2781
rect 1823 2772 1827 2776
rect 1863 2764 1867 2768
rect 175 2759 179 2763
rect 303 2759 307 2763
rect 431 2759 435 2763
rect 567 2759 571 2763
rect 703 2759 707 2763
rect 831 2759 835 2763
rect 959 2759 963 2763
rect 1087 2759 1091 2763
rect 1215 2759 1219 2763
rect 3575 2764 3579 2768
rect 1351 2759 1355 2763
rect 1863 2747 1867 2751
rect 3575 2747 3579 2751
rect 1887 2737 1891 2741
rect 2055 2737 2059 2741
rect 2247 2737 2251 2741
rect 2431 2737 2435 2741
rect 2607 2737 2611 2741
rect 2775 2737 2779 2741
rect 2927 2737 2931 2741
rect 3071 2737 3075 2741
rect 3215 2737 3219 2741
rect 3359 2737 3363 2741
rect 3479 2737 3483 2741
rect 143 2717 147 2721
rect 231 2717 235 2721
rect 351 2717 355 2721
rect 479 2717 483 2721
rect 615 2717 619 2721
rect 759 2717 763 2721
rect 903 2717 907 2721
rect 1047 2717 1051 2721
rect 1887 2711 1891 2715
rect 2047 2711 2051 2715
rect 2207 2711 2211 2715
rect 2359 2711 2363 2715
rect 2495 2711 2499 2715
rect 2623 2711 2627 2715
rect 2743 2711 2747 2715
rect 2863 2711 2867 2715
rect 2983 2711 2987 2715
rect 3103 2711 3107 2715
rect 111 2704 115 2708
rect 1823 2704 1827 2708
rect 1863 2701 1867 2705
rect 3575 2701 3579 2705
rect 111 2687 115 2691
rect 1823 2687 1827 2691
rect 1863 2684 1867 2688
rect 3575 2684 3579 2688
rect 135 2677 139 2681
rect 223 2677 227 2681
rect 343 2677 347 2681
rect 471 2677 475 2681
rect 607 2677 611 2681
rect 751 2677 755 2681
rect 895 2677 899 2681
rect 1039 2677 1043 2681
rect 1895 2671 1899 2675
rect 2055 2671 2059 2675
rect 2215 2671 2219 2675
rect 2367 2671 2371 2675
rect 2503 2671 2507 2675
rect 2631 2671 2635 2675
rect 2751 2671 2755 2675
rect 2871 2671 2875 2675
rect 2991 2671 2995 2675
rect 3111 2671 3115 2675
rect 135 2651 139 2655
rect 231 2651 235 2655
rect 351 2651 355 2655
rect 471 2651 475 2655
rect 583 2651 587 2655
rect 695 2651 699 2655
rect 799 2651 803 2655
rect 903 2651 907 2655
rect 999 2651 1003 2655
rect 1103 2651 1107 2655
rect 1207 2651 1211 2655
rect 1311 2651 1315 2655
rect 111 2641 115 2645
rect 1823 2641 1827 2645
rect 1895 2629 1899 2633
rect 111 2624 115 2628
rect 1999 2629 2003 2633
rect 2119 2629 2123 2633
rect 2239 2629 2243 2633
rect 2351 2629 2355 2633
rect 2455 2629 2459 2633
rect 2551 2629 2555 2633
rect 2655 2629 2659 2633
rect 2759 2629 2763 2633
rect 2863 2629 2867 2633
rect 1823 2624 1827 2628
rect 1863 2616 1867 2620
rect 143 2611 147 2615
rect 239 2611 243 2615
rect 359 2611 363 2615
rect 479 2611 483 2615
rect 591 2611 595 2615
rect 703 2611 707 2615
rect 807 2611 811 2615
rect 911 2611 915 2615
rect 1007 2611 1011 2615
rect 1111 2611 1115 2615
rect 1215 2611 1219 2615
rect 3575 2616 3579 2620
rect 1319 2611 1323 2615
rect 1863 2599 1867 2603
rect 3575 2599 3579 2603
rect 1887 2589 1891 2593
rect 1991 2589 1995 2593
rect 2111 2589 2115 2593
rect 2231 2589 2235 2593
rect 2343 2589 2347 2593
rect 2447 2589 2451 2593
rect 2543 2589 2547 2593
rect 2647 2589 2651 2593
rect 2751 2589 2755 2593
rect 2855 2589 2859 2593
rect 143 2573 147 2577
rect 271 2573 275 2577
rect 415 2573 419 2577
rect 551 2573 555 2577
rect 679 2573 683 2577
rect 807 2573 811 2577
rect 927 2573 931 2577
rect 1047 2573 1051 2577
rect 1175 2573 1179 2577
rect 111 2560 115 2564
rect 1823 2560 1827 2564
rect 1887 2563 1891 2567
rect 1991 2563 1995 2567
rect 2111 2563 2115 2567
rect 2231 2563 2235 2567
rect 2351 2563 2355 2567
rect 2471 2563 2475 2567
rect 2591 2563 2595 2567
rect 2711 2563 2715 2567
rect 2831 2563 2835 2567
rect 1863 2553 1867 2557
rect 3575 2553 3579 2557
rect 111 2543 115 2547
rect 1823 2543 1827 2547
rect 135 2533 139 2537
rect 263 2533 267 2537
rect 407 2533 411 2537
rect 543 2533 547 2537
rect 671 2533 675 2537
rect 799 2533 803 2537
rect 919 2533 923 2537
rect 1039 2533 1043 2537
rect 1167 2533 1171 2537
rect 1863 2536 1867 2540
rect 3575 2536 3579 2540
rect 1895 2523 1899 2527
rect 1999 2523 2003 2527
rect 2119 2523 2123 2527
rect 2239 2523 2243 2527
rect 2359 2523 2363 2527
rect 2479 2523 2483 2527
rect 2599 2523 2603 2527
rect 2719 2523 2723 2527
rect 2839 2523 2843 2527
rect 135 2511 139 2515
rect 279 2511 283 2515
rect 439 2511 443 2515
rect 591 2511 595 2515
rect 735 2511 739 2515
rect 871 2511 875 2515
rect 1007 2511 1011 2515
rect 1143 2511 1147 2515
rect 1279 2511 1283 2515
rect 111 2501 115 2505
rect 1823 2501 1827 2505
rect 111 2484 115 2488
rect 1823 2484 1827 2488
rect 1895 2485 1899 2489
rect 2031 2485 2035 2489
rect 2191 2485 2195 2489
rect 2343 2485 2347 2489
rect 2487 2485 2491 2489
rect 2623 2485 2627 2489
rect 2751 2485 2755 2489
rect 2879 2485 2883 2489
rect 3015 2485 3019 2489
rect 143 2471 147 2475
rect 287 2471 291 2475
rect 447 2471 451 2475
rect 599 2471 603 2475
rect 743 2471 747 2475
rect 879 2471 883 2475
rect 1015 2471 1019 2475
rect 1151 2471 1155 2475
rect 1287 2471 1291 2475
rect 1863 2472 1867 2476
rect 3575 2472 3579 2476
rect 1863 2455 1867 2459
rect 3575 2455 3579 2459
rect 1887 2445 1891 2449
rect 2023 2445 2027 2449
rect 2183 2445 2187 2449
rect 2335 2445 2339 2449
rect 2479 2445 2483 2449
rect 2615 2445 2619 2449
rect 2743 2445 2747 2449
rect 2871 2445 2875 2449
rect 3007 2445 3011 2449
rect 191 2437 195 2441
rect 319 2437 323 2441
rect 455 2437 459 2441
rect 591 2437 595 2441
rect 727 2437 731 2441
rect 863 2437 867 2441
rect 999 2437 1003 2441
rect 1135 2437 1139 2441
rect 1271 2437 1275 2441
rect 1407 2437 1411 2441
rect 111 2424 115 2428
rect 1823 2424 1827 2428
rect 1887 2423 1891 2427
rect 2015 2423 2019 2427
rect 2175 2423 2179 2427
rect 2335 2423 2339 2427
rect 2495 2423 2499 2427
rect 2647 2423 2651 2427
rect 2799 2423 2803 2427
rect 2951 2423 2955 2427
rect 3111 2423 3115 2427
rect 1863 2413 1867 2417
rect 3575 2413 3579 2417
rect 111 2407 115 2411
rect 1823 2407 1827 2411
rect 183 2397 187 2401
rect 311 2397 315 2401
rect 447 2397 451 2401
rect 583 2397 587 2401
rect 719 2397 723 2401
rect 855 2397 859 2401
rect 991 2397 995 2401
rect 1127 2397 1131 2401
rect 1263 2397 1267 2401
rect 1399 2397 1403 2401
rect 1863 2396 1867 2400
rect 3575 2396 3579 2400
rect 1895 2383 1899 2387
rect 2023 2383 2027 2387
rect 2183 2383 2187 2387
rect 2343 2383 2347 2387
rect 2503 2383 2507 2387
rect 2655 2383 2659 2387
rect 2807 2383 2811 2387
rect 2959 2383 2963 2387
rect 3119 2383 3123 2387
rect 159 2363 163 2367
rect 247 2363 251 2367
rect 335 2363 339 2367
rect 439 2363 443 2367
rect 559 2363 563 2367
rect 687 2363 691 2367
rect 815 2363 819 2367
rect 951 2363 955 2367
rect 1079 2363 1083 2367
rect 1207 2363 1211 2367
rect 1327 2363 1331 2367
rect 1455 2363 1459 2367
rect 1583 2363 1587 2367
rect 111 2353 115 2357
rect 1823 2353 1827 2357
rect 1927 2345 1931 2349
rect 2087 2345 2091 2349
rect 2247 2345 2251 2349
rect 2407 2345 2411 2349
rect 2559 2345 2563 2349
rect 2703 2345 2707 2349
rect 2831 2345 2835 2349
rect 2951 2345 2955 2349
rect 3071 2345 3075 2349
rect 3183 2345 3187 2349
rect 3287 2345 3291 2349
rect 3399 2345 3403 2349
rect 3487 2345 3491 2349
rect 111 2336 115 2340
rect 1823 2336 1827 2340
rect 1863 2332 1867 2336
rect 3575 2332 3579 2336
rect 167 2323 171 2327
rect 255 2323 259 2327
rect 343 2323 347 2327
rect 447 2323 451 2327
rect 567 2323 571 2327
rect 695 2323 699 2327
rect 823 2323 827 2327
rect 959 2323 963 2327
rect 1087 2323 1091 2327
rect 1215 2323 1219 2327
rect 1335 2323 1339 2327
rect 1463 2323 1467 2327
rect 1591 2323 1595 2327
rect 1863 2315 1867 2319
rect 3575 2315 3579 2319
rect 1919 2305 1923 2309
rect 2079 2305 2083 2309
rect 2239 2305 2243 2309
rect 2399 2305 2403 2309
rect 2551 2305 2555 2309
rect 2695 2305 2699 2309
rect 2823 2305 2827 2309
rect 2943 2305 2947 2309
rect 3063 2305 3067 2309
rect 3175 2305 3179 2309
rect 3279 2305 3283 2309
rect 3391 2305 3395 2309
rect 3479 2305 3483 2309
rect 695 2281 699 2285
rect 863 2281 867 2285
rect 1023 2281 1027 2285
rect 1175 2281 1179 2285
rect 1319 2281 1323 2285
rect 1463 2281 1467 2285
rect 1599 2281 1603 2285
rect 1735 2281 1739 2285
rect 1975 2279 1979 2283
rect 2143 2279 2147 2283
rect 2311 2279 2315 2283
rect 2479 2279 2483 2283
rect 2639 2279 2643 2283
rect 2783 2279 2787 2283
rect 2919 2279 2923 2283
rect 3039 2279 3043 2283
rect 3159 2279 3163 2283
rect 3271 2279 3275 2283
rect 3383 2279 3387 2283
rect 3479 2279 3483 2283
rect 111 2268 115 2272
rect 1823 2268 1827 2272
rect 1863 2269 1867 2273
rect 3575 2269 3579 2273
rect 111 2251 115 2255
rect 1823 2251 1827 2255
rect 1863 2252 1867 2256
rect 3575 2252 3579 2256
rect 687 2241 691 2245
rect 855 2241 859 2245
rect 1015 2241 1019 2245
rect 1167 2241 1171 2245
rect 1311 2241 1315 2245
rect 1455 2241 1459 2245
rect 1591 2241 1595 2245
rect 1727 2241 1731 2245
rect 1983 2239 1987 2243
rect 2151 2239 2155 2243
rect 2319 2239 2323 2243
rect 2487 2239 2491 2243
rect 2647 2239 2651 2243
rect 2791 2239 2795 2243
rect 2927 2239 2931 2243
rect 3047 2239 3051 2243
rect 3167 2239 3171 2243
rect 3279 2239 3283 2243
rect 3391 2239 3395 2243
rect 3487 2239 3491 2243
rect 535 2211 539 2215
rect 719 2211 723 2215
rect 895 2211 899 2215
rect 1071 2211 1075 2215
rect 1239 2211 1243 2215
rect 1407 2211 1411 2215
rect 1575 2211 1579 2215
rect 1727 2211 1731 2215
rect 111 2201 115 2205
rect 1823 2201 1827 2205
rect 2007 2205 2011 2209
rect 2167 2205 2171 2209
rect 2335 2205 2339 2209
rect 2519 2205 2523 2209
rect 2711 2205 2715 2209
rect 2903 2205 2907 2209
rect 3103 2205 3107 2209
rect 3303 2205 3307 2209
rect 3487 2205 3491 2209
rect 1863 2192 1867 2196
rect 3575 2192 3579 2196
rect 111 2184 115 2188
rect 1823 2184 1827 2188
rect 543 2171 547 2175
rect 727 2171 731 2175
rect 903 2171 907 2175
rect 1079 2171 1083 2175
rect 1247 2171 1251 2175
rect 1415 2171 1419 2175
rect 1583 2171 1587 2175
rect 1735 2171 1739 2175
rect 1863 2175 1867 2179
rect 3575 2175 3579 2179
rect 1999 2165 2003 2169
rect 2159 2165 2163 2169
rect 2327 2165 2331 2169
rect 2511 2165 2515 2169
rect 2703 2165 2707 2169
rect 2895 2165 2899 2169
rect 3095 2165 3099 2169
rect 3295 2165 3299 2169
rect 3479 2165 3483 2169
rect 495 2137 499 2141
rect 623 2137 627 2141
rect 759 2137 763 2141
rect 895 2137 899 2141
rect 1039 2137 1043 2141
rect 1183 2137 1187 2141
rect 1327 2137 1331 2141
rect 1471 2137 1475 2141
rect 1623 2137 1627 2141
rect 2023 2135 2027 2139
rect 2167 2135 2171 2139
rect 2319 2135 2323 2139
rect 2471 2135 2475 2139
rect 2615 2135 2619 2139
rect 2759 2135 2763 2139
rect 2895 2135 2899 2139
rect 3023 2135 3027 2139
rect 3143 2135 3147 2139
rect 3263 2135 3267 2139
rect 3383 2135 3387 2139
rect 3479 2135 3483 2139
rect 111 2124 115 2128
rect 1823 2124 1827 2128
rect 1863 2125 1867 2129
rect 3575 2125 3579 2129
rect 111 2107 115 2111
rect 1823 2107 1827 2111
rect 1863 2108 1867 2112
rect 3575 2108 3579 2112
rect 487 2097 491 2101
rect 615 2097 619 2101
rect 751 2097 755 2101
rect 887 2097 891 2101
rect 1031 2097 1035 2101
rect 1175 2097 1179 2101
rect 1319 2097 1323 2101
rect 1463 2097 1467 2101
rect 1615 2097 1619 2101
rect 2031 2095 2035 2099
rect 2175 2095 2179 2099
rect 2327 2095 2331 2099
rect 2479 2095 2483 2099
rect 2623 2095 2627 2099
rect 2767 2095 2771 2099
rect 2903 2095 2907 2099
rect 3031 2095 3035 2099
rect 3151 2095 3155 2099
rect 3271 2095 3275 2099
rect 3391 2095 3395 2099
rect 3487 2095 3491 2099
rect 319 2071 323 2075
rect 431 2071 435 2075
rect 551 2071 555 2075
rect 679 2071 683 2075
rect 799 2071 803 2075
rect 919 2071 923 2075
rect 1039 2071 1043 2075
rect 1159 2071 1163 2075
rect 1279 2071 1283 2075
rect 1407 2071 1411 2075
rect 111 2061 115 2065
rect 1823 2061 1827 2065
rect 1983 2057 1987 2061
rect 2143 2057 2147 2061
rect 2311 2057 2315 2061
rect 2471 2057 2475 2061
rect 2631 2057 2635 2061
rect 2775 2057 2779 2061
rect 2911 2057 2915 2061
rect 3039 2057 3043 2061
rect 3159 2057 3163 2061
rect 3279 2057 3283 2061
rect 3391 2057 3395 2061
rect 3487 2057 3491 2061
rect 111 2044 115 2048
rect 1823 2044 1827 2048
rect 1863 2044 1867 2048
rect 3575 2044 3579 2048
rect 327 2031 331 2035
rect 439 2031 443 2035
rect 559 2031 563 2035
rect 687 2031 691 2035
rect 807 2031 811 2035
rect 927 2031 931 2035
rect 1047 2031 1051 2035
rect 1167 2031 1171 2035
rect 1287 2031 1291 2035
rect 1415 2031 1419 2035
rect 1863 2027 1867 2031
rect 3575 2027 3579 2031
rect 1975 2017 1979 2021
rect 2135 2017 2139 2021
rect 2303 2017 2307 2021
rect 2463 2017 2467 2021
rect 2623 2017 2627 2021
rect 2767 2017 2771 2021
rect 2903 2017 2907 2021
rect 3031 2017 3035 2021
rect 3151 2017 3155 2021
rect 3271 2017 3275 2021
rect 3383 2017 3387 2021
rect 3479 2017 3483 2021
rect 183 1993 187 1997
rect 295 1993 299 1997
rect 415 1993 419 1997
rect 535 1993 539 1997
rect 655 1993 659 1997
rect 775 1993 779 1997
rect 895 1993 899 1997
rect 1015 1993 1019 1997
rect 1135 1993 1139 1997
rect 1255 1993 1259 1997
rect 1887 1995 1891 1999
rect 2031 1995 2035 1999
rect 2199 1995 2203 1999
rect 2375 1995 2379 1999
rect 2543 1995 2547 1999
rect 2711 1995 2715 1999
rect 2871 1995 2875 1999
rect 3039 1995 3043 1999
rect 3207 1995 3211 1999
rect 1863 1985 1867 1989
rect 111 1980 115 1984
rect 3575 1985 3579 1989
rect 1823 1980 1827 1984
rect 1863 1968 1867 1972
rect 111 1963 115 1967
rect 3575 1968 3579 1972
rect 1823 1963 1827 1967
rect 175 1953 179 1957
rect 287 1953 291 1957
rect 407 1953 411 1957
rect 527 1953 531 1957
rect 647 1953 651 1957
rect 767 1953 771 1957
rect 887 1953 891 1957
rect 1007 1953 1011 1957
rect 1127 1953 1131 1957
rect 1247 1953 1251 1957
rect 1895 1955 1899 1959
rect 2039 1955 2043 1959
rect 2207 1955 2211 1959
rect 2383 1955 2387 1959
rect 2551 1955 2555 1959
rect 2719 1955 2723 1959
rect 2879 1955 2883 1959
rect 3047 1955 3051 1959
rect 3215 1955 3219 1959
rect 135 1927 139 1931
rect 223 1927 227 1931
rect 351 1927 355 1931
rect 495 1927 499 1931
rect 655 1927 659 1931
rect 839 1927 843 1931
rect 1039 1927 1043 1931
rect 1247 1927 1251 1931
rect 1463 1927 1467 1931
rect 111 1917 115 1921
rect 1823 1917 1827 1921
rect 1895 1913 1899 1917
rect 1991 1913 1995 1917
rect 2119 1913 2123 1917
rect 2255 1913 2259 1917
rect 2383 1913 2387 1917
rect 2511 1913 2515 1917
rect 2631 1913 2635 1917
rect 2751 1913 2755 1917
rect 2879 1913 2883 1917
rect 3007 1913 3011 1917
rect 111 1900 115 1904
rect 1823 1900 1827 1904
rect 1863 1900 1867 1904
rect 3575 1900 3579 1904
rect 143 1887 147 1891
rect 231 1887 235 1891
rect 359 1887 363 1891
rect 503 1887 507 1891
rect 663 1887 667 1891
rect 847 1887 851 1891
rect 1047 1887 1051 1891
rect 1255 1887 1259 1891
rect 1471 1887 1475 1891
rect 1863 1883 1867 1887
rect 3575 1883 3579 1887
rect 1887 1873 1891 1877
rect 1983 1873 1987 1877
rect 2111 1873 2115 1877
rect 2247 1873 2251 1877
rect 2375 1873 2379 1877
rect 2503 1873 2507 1877
rect 2623 1873 2627 1877
rect 2743 1873 2747 1877
rect 2871 1873 2875 1877
rect 2999 1873 3003 1877
rect 143 1845 147 1849
rect 271 1845 275 1849
rect 415 1845 419 1849
rect 559 1845 563 1849
rect 695 1845 699 1849
rect 823 1845 827 1849
rect 943 1845 947 1849
rect 1055 1845 1059 1849
rect 1159 1845 1163 1849
rect 1263 1845 1267 1849
rect 1359 1845 1363 1849
rect 1455 1845 1459 1849
rect 1551 1845 1555 1849
rect 1647 1845 1651 1849
rect 1735 1845 1739 1849
rect 2223 1843 2227 1847
rect 2359 1843 2363 1847
rect 2495 1843 2499 1847
rect 2623 1843 2627 1847
rect 2743 1843 2747 1847
rect 2863 1843 2867 1847
rect 2991 1843 2995 1847
rect 111 1832 115 1836
rect 1823 1832 1827 1836
rect 1863 1833 1867 1837
rect 3575 1833 3579 1837
rect 111 1815 115 1819
rect 1823 1815 1827 1819
rect 1863 1816 1867 1820
rect 3575 1816 3579 1820
rect 135 1805 139 1809
rect 263 1805 267 1809
rect 407 1805 411 1809
rect 551 1805 555 1809
rect 687 1805 691 1809
rect 815 1805 819 1809
rect 935 1805 939 1809
rect 1047 1805 1051 1809
rect 1151 1805 1155 1809
rect 1255 1805 1259 1809
rect 1351 1805 1355 1809
rect 1447 1805 1451 1809
rect 1543 1805 1547 1809
rect 1639 1805 1643 1809
rect 1727 1805 1731 1809
rect 2231 1803 2235 1807
rect 2367 1803 2371 1807
rect 2503 1803 2507 1807
rect 2631 1803 2635 1807
rect 2751 1803 2755 1807
rect 2871 1803 2875 1807
rect 2999 1803 3003 1807
rect 135 1771 139 1775
rect 303 1771 307 1775
rect 495 1771 499 1775
rect 687 1771 691 1775
rect 871 1771 875 1775
rect 1047 1771 1051 1775
rect 1215 1771 1219 1775
rect 1375 1771 1379 1775
rect 1535 1771 1539 1775
rect 1703 1771 1707 1775
rect 111 1761 115 1765
rect 1823 1761 1827 1765
rect 2271 1765 2275 1769
rect 2359 1765 2363 1769
rect 2455 1765 2459 1769
rect 2559 1765 2563 1769
rect 2663 1765 2667 1769
rect 2759 1765 2763 1769
rect 2863 1765 2867 1769
rect 2967 1765 2971 1769
rect 3071 1765 3075 1769
rect 3175 1765 3179 1769
rect 1863 1752 1867 1756
rect 3575 1752 3579 1756
rect 111 1744 115 1748
rect 1823 1744 1827 1748
rect 143 1731 147 1735
rect 311 1731 315 1735
rect 503 1731 507 1735
rect 695 1731 699 1735
rect 879 1731 883 1735
rect 1055 1731 1059 1735
rect 1223 1731 1227 1735
rect 1383 1731 1387 1735
rect 1543 1731 1547 1735
rect 1711 1731 1715 1735
rect 1863 1735 1867 1739
rect 3575 1735 3579 1739
rect 2263 1725 2267 1729
rect 2351 1725 2355 1729
rect 2447 1725 2451 1729
rect 2551 1725 2555 1729
rect 2655 1725 2659 1729
rect 2751 1725 2755 1729
rect 2855 1725 2859 1729
rect 2959 1725 2963 1729
rect 3063 1725 3067 1729
rect 3167 1725 3171 1729
rect 2247 1699 2251 1703
rect 2367 1699 2371 1703
rect 2495 1699 2499 1703
rect 2623 1699 2627 1703
rect 2759 1699 2763 1703
rect 2887 1699 2891 1703
rect 3015 1699 3019 1703
rect 3135 1699 3139 1703
rect 3247 1699 3251 1703
rect 3367 1699 3371 1703
rect 3479 1699 3483 1703
rect 143 1693 147 1697
rect 287 1693 291 1697
rect 471 1693 475 1697
rect 655 1693 659 1697
rect 839 1693 843 1697
rect 1023 1693 1027 1697
rect 1191 1693 1195 1697
rect 1359 1693 1363 1697
rect 1527 1693 1531 1697
rect 1695 1693 1699 1697
rect 1863 1689 1867 1693
rect 3575 1689 3579 1693
rect 111 1680 115 1684
rect 1823 1680 1827 1684
rect 1863 1672 1867 1676
rect 3575 1672 3579 1676
rect 111 1663 115 1667
rect 1823 1663 1827 1667
rect 2255 1659 2259 1663
rect 2375 1659 2379 1663
rect 2503 1659 2507 1663
rect 2631 1659 2635 1663
rect 2767 1659 2771 1663
rect 2895 1659 2899 1663
rect 3023 1659 3027 1663
rect 3143 1659 3147 1663
rect 3255 1659 3259 1663
rect 3375 1659 3379 1663
rect 3487 1659 3491 1663
rect 135 1653 139 1657
rect 279 1653 283 1657
rect 463 1653 467 1657
rect 647 1653 651 1657
rect 831 1653 835 1657
rect 1015 1653 1019 1657
rect 1183 1653 1187 1657
rect 1351 1653 1355 1657
rect 1519 1653 1523 1657
rect 1687 1653 1691 1657
rect 135 1623 139 1627
rect 271 1623 275 1627
rect 447 1623 451 1627
rect 631 1623 635 1627
rect 815 1623 819 1627
rect 991 1623 995 1627
rect 1151 1623 1155 1627
rect 1303 1623 1307 1627
rect 1455 1623 1459 1627
rect 1599 1623 1603 1627
rect 1727 1623 1731 1627
rect 2151 1621 2155 1625
rect 2343 1621 2347 1625
rect 2527 1621 2531 1625
rect 2703 1621 2707 1625
rect 2871 1621 2875 1625
rect 3031 1621 3035 1625
rect 3191 1621 3195 1625
rect 3351 1621 3355 1625
rect 3487 1621 3491 1625
rect 111 1613 115 1617
rect 1823 1613 1827 1617
rect 1863 1608 1867 1612
rect 3575 1608 3579 1612
rect 111 1596 115 1600
rect 1823 1596 1827 1600
rect 1863 1591 1867 1595
rect 3575 1591 3579 1595
rect 143 1583 147 1587
rect 279 1583 283 1587
rect 455 1583 459 1587
rect 639 1583 643 1587
rect 823 1583 827 1587
rect 999 1583 1003 1587
rect 1159 1583 1163 1587
rect 1311 1583 1315 1587
rect 1463 1583 1467 1587
rect 1607 1583 1611 1587
rect 1735 1583 1739 1587
rect 2143 1581 2147 1585
rect 2335 1581 2339 1585
rect 2519 1581 2523 1585
rect 2695 1581 2699 1585
rect 2863 1581 2867 1585
rect 3023 1581 3027 1585
rect 3183 1581 3187 1585
rect 3343 1581 3347 1585
rect 3479 1581 3483 1585
rect 2087 1559 2091 1563
rect 2279 1559 2283 1563
rect 2455 1559 2459 1563
rect 2623 1559 2627 1563
rect 2791 1559 2795 1563
rect 2951 1559 2955 1563
rect 3111 1559 3115 1563
rect 3271 1559 3275 1563
rect 3431 1559 3435 1563
rect 143 1549 147 1553
rect 271 1549 275 1553
rect 431 1549 435 1553
rect 599 1549 603 1553
rect 767 1549 771 1553
rect 935 1549 939 1553
rect 1103 1549 1107 1553
rect 1263 1549 1267 1553
rect 1423 1549 1427 1553
rect 1591 1549 1595 1553
rect 1735 1549 1739 1553
rect 1863 1549 1867 1553
rect 3575 1549 3579 1553
rect 111 1536 115 1540
rect 1823 1536 1827 1540
rect 1863 1532 1867 1536
rect 3575 1532 3579 1536
rect 111 1519 115 1523
rect 1823 1519 1827 1523
rect 2095 1519 2099 1523
rect 2287 1519 2291 1523
rect 2463 1519 2467 1523
rect 2631 1519 2635 1523
rect 2799 1519 2803 1523
rect 2959 1519 2963 1523
rect 3119 1519 3123 1523
rect 3279 1519 3283 1523
rect 3439 1519 3443 1523
rect 135 1509 139 1513
rect 263 1509 267 1513
rect 423 1509 427 1513
rect 591 1509 595 1513
rect 759 1509 763 1513
rect 927 1509 931 1513
rect 1095 1509 1099 1513
rect 1255 1509 1259 1513
rect 1415 1509 1419 1513
rect 1583 1509 1587 1513
rect 1727 1509 1731 1513
rect 183 1483 187 1487
rect 327 1483 331 1487
rect 471 1483 475 1487
rect 607 1483 611 1487
rect 743 1483 747 1487
rect 871 1483 875 1487
rect 991 1483 995 1487
rect 1119 1483 1123 1487
rect 1247 1483 1251 1487
rect 1375 1483 1379 1487
rect 111 1473 115 1477
rect 1823 1473 1827 1477
rect 1895 1477 1899 1481
rect 1991 1477 1995 1481
rect 2119 1477 2123 1481
rect 2247 1477 2251 1481
rect 2383 1477 2387 1481
rect 2535 1477 2539 1481
rect 2703 1477 2707 1481
rect 2887 1477 2891 1481
rect 3087 1477 3091 1481
rect 3295 1477 3299 1481
rect 3487 1477 3491 1481
rect 1863 1464 1867 1468
rect 3575 1464 3579 1468
rect 111 1456 115 1460
rect 1823 1456 1827 1460
rect 191 1443 195 1447
rect 335 1443 339 1447
rect 479 1443 483 1447
rect 615 1443 619 1447
rect 751 1443 755 1447
rect 879 1443 883 1447
rect 999 1443 1003 1447
rect 1127 1443 1131 1447
rect 1255 1443 1259 1447
rect 1383 1443 1387 1447
rect 1863 1447 1867 1451
rect 3575 1447 3579 1451
rect 1887 1437 1891 1441
rect 1983 1437 1987 1441
rect 2111 1437 2115 1441
rect 2239 1437 2243 1441
rect 2375 1437 2379 1441
rect 2527 1437 2531 1441
rect 2695 1437 2699 1441
rect 2879 1437 2883 1441
rect 3079 1437 3083 1441
rect 3287 1437 3291 1441
rect 3479 1437 3483 1441
rect 1887 1411 1891 1415
rect 1975 1411 1979 1415
rect 2071 1411 2075 1415
rect 2183 1411 2187 1415
rect 2303 1411 2307 1415
rect 2439 1411 2443 1415
rect 2607 1411 2611 1415
rect 2807 1411 2811 1415
rect 3031 1411 3035 1415
rect 3263 1411 3267 1415
rect 3479 1411 3483 1415
rect 199 1401 203 1405
rect 335 1401 339 1405
rect 463 1401 467 1405
rect 583 1401 587 1405
rect 703 1401 707 1405
rect 815 1401 819 1405
rect 919 1401 923 1405
rect 1015 1401 1019 1405
rect 1119 1401 1123 1405
rect 1223 1401 1227 1405
rect 1327 1401 1331 1405
rect 1863 1401 1867 1405
rect 3575 1401 3579 1405
rect 111 1388 115 1392
rect 1823 1388 1827 1392
rect 1863 1384 1867 1388
rect 3575 1384 3579 1388
rect 111 1371 115 1375
rect 1823 1371 1827 1375
rect 1895 1371 1899 1375
rect 1983 1371 1987 1375
rect 2079 1371 2083 1375
rect 2191 1371 2195 1375
rect 2311 1371 2315 1375
rect 2447 1371 2451 1375
rect 2615 1371 2619 1375
rect 2815 1371 2819 1375
rect 3039 1371 3043 1375
rect 3271 1371 3275 1375
rect 3487 1371 3491 1375
rect 191 1361 195 1365
rect 327 1361 331 1365
rect 455 1361 459 1365
rect 575 1361 579 1365
rect 695 1361 699 1365
rect 807 1361 811 1365
rect 911 1361 915 1365
rect 1007 1361 1011 1365
rect 1111 1361 1115 1365
rect 1215 1361 1219 1365
rect 1319 1361 1323 1365
rect 231 1335 235 1339
rect 383 1335 387 1339
rect 543 1335 547 1339
rect 703 1335 707 1339
rect 871 1335 875 1339
rect 1039 1335 1043 1339
rect 1207 1335 1211 1339
rect 1375 1335 1379 1339
rect 1895 1333 1899 1337
rect 1983 1333 1987 1337
rect 2103 1333 2107 1337
rect 2223 1333 2227 1337
rect 2359 1333 2363 1337
rect 2511 1333 2515 1337
rect 2687 1333 2691 1337
rect 2871 1333 2875 1337
rect 3071 1333 3075 1337
rect 3279 1333 3283 1337
rect 3487 1333 3491 1337
rect 111 1325 115 1329
rect 1823 1325 1827 1329
rect 1863 1320 1867 1324
rect 3575 1320 3579 1324
rect 111 1308 115 1312
rect 1823 1308 1827 1312
rect 1863 1303 1867 1307
rect 3575 1303 3579 1307
rect 239 1295 243 1299
rect 391 1295 395 1299
rect 551 1295 555 1299
rect 711 1295 715 1299
rect 879 1295 883 1299
rect 1047 1295 1051 1299
rect 1215 1295 1219 1299
rect 1383 1295 1387 1299
rect 1887 1293 1891 1297
rect 1975 1293 1979 1297
rect 2095 1293 2099 1297
rect 2215 1293 2219 1297
rect 2351 1293 2355 1297
rect 2503 1293 2507 1297
rect 2679 1293 2683 1297
rect 2863 1293 2867 1297
rect 3063 1293 3067 1297
rect 3271 1293 3275 1297
rect 3479 1293 3483 1297
rect 215 1261 219 1265
rect 359 1261 363 1265
rect 519 1261 523 1265
rect 679 1261 683 1265
rect 839 1261 843 1265
rect 999 1261 1003 1265
rect 1151 1261 1155 1265
rect 1295 1261 1299 1265
rect 1439 1261 1443 1265
rect 1591 1261 1595 1265
rect 2055 1259 2059 1263
rect 2143 1259 2147 1263
rect 2239 1259 2243 1263
rect 2335 1259 2339 1263
rect 2431 1259 2435 1263
rect 2551 1259 2555 1263
rect 2687 1259 2691 1263
rect 2855 1259 2859 1263
rect 3039 1259 3043 1263
rect 3231 1259 3235 1263
rect 3431 1259 3435 1263
rect 111 1248 115 1252
rect 1823 1248 1827 1252
rect 1863 1249 1867 1253
rect 3575 1249 3579 1253
rect 111 1231 115 1235
rect 1823 1231 1827 1235
rect 1863 1232 1867 1236
rect 3575 1232 3579 1236
rect 207 1221 211 1225
rect 351 1221 355 1225
rect 511 1221 515 1225
rect 671 1221 675 1225
rect 831 1221 835 1225
rect 991 1221 995 1225
rect 1143 1221 1147 1225
rect 1287 1221 1291 1225
rect 1431 1221 1435 1225
rect 1583 1221 1587 1225
rect 2063 1219 2067 1223
rect 2151 1219 2155 1223
rect 2247 1219 2251 1223
rect 2343 1219 2347 1223
rect 2439 1219 2443 1223
rect 2559 1219 2563 1223
rect 2695 1219 2699 1223
rect 2863 1219 2867 1223
rect 3047 1219 3051 1223
rect 3239 1219 3243 1223
rect 3439 1219 3443 1223
rect 135 1191 139 1195
rect 271 1191 275 1195
rect 423 1191 427 1195
rect 575 1191 579 1195
rect 727 1191 731 1195
rect 887 1191 891 1195
rect 1055 1191 1059 1195
rect 1231 1191 1235 1195
rect 1415 1191 1419 1195
rect 1599 1191 1603 1195
rect 111 1181 115 1185
rect 1823 1181 1827 1185
rect 2039 1181 2043 1185
rect 2151 1181 2155 1185
rect 2279 1181 2283 1185
rect 2415 1181 2419 1185
rect 2559 1181 2563 1185
rect 2711 1181 2715 1185
rect 2863 1181 2867 1185
rect 3015 1181 3019 1185
rect 3167 1181 3171 1185
rect 3327 1181 3331 1185
rect 3487 1181 3491 1185
rect 111 1164 115 1168
rect 1823 1164 1827 1168
rect 1863 1168 1867 1172
rect 3575 1168 3579 1172
rect 143 1151 147 1155
rect 279 1151 283 1155
rect 431 1151 435 1155
rect 583 1151 587 1155
rect 735 1151 739 1155
rect 895 1151 899 1155
rect 1063 1151 1067 1155
rect 1239 1151 1243 1155
rect 1423 1151 1427 1155
rect 1607 1151 1611 1155
rect 1863 1151 1867 1155
rect 3575 1151 3579 1155
rect 2031 1141 2035 1145
rect 2143 1141 2147 1145
rect 2271 1141 2275 1145
rect 2407 1141 2411 1145
rect 2551 1141 2555 1145
rect 2703 1141 2707 1145
rect 2855 1141 2859 1145
rect 3007 1141 3011 1145
rect 3159 1141 3163 1145
rect 3319 1141 3323 1145
rect 3479 1141 3483 1145
rect 143 1117 147 1121
rect 295 1117 299 1121
rect 479 1117 483 1121
rect 663 1117 667 1121
rect 847 1117 851 1121
rect 1031 1117 1035 1121
rect 1207 1117 1211 1121
rect 1391 1117 1395 1121
rect 1575 1117 1579 1121
rect 1735 1117 1739 1121
rect 111 1104 115 1108
rect 1823 1104 1827 1108
rect 1943 1107 1947 1111
rect 2087 1107 2091 1111
rect 2231 1107 2235 1111
rect 2383 1107 2387 1111
rect 2535 1107 2539 1111
rect 2687 1107 2691 1111
rect 2839 1107 2843 1111
rect 2991 1107 2995 1111
rect 3151 1107 3155 1111
rect 3319 1107 3323 1111
rect 3479 1107 3483 1111
rect 1863 1097 1867 1101
rect 3575 1097 3579 1101
rect 111 1087 115 1091
rect 1823 1087 1827 1091
rect 135 1077 139 1081
rect 287 1077 291 1081
rect 471 1077 475 1081
rect 655 1077 659 1081
rect 839 1077 843 1081
rect 1023 1077 1027 1081
rect 1199 1077 1203 1081
rect 1383 1077 1387 1081
rect 1567 1077 1571 1081
rect 1727 1077 1731 1081
rect 1863 1080 1867 1084
rect 3575 1080 3579 1084
rect 1951 1067 1955 1071
rect 2095 1067 2099 1071
rect 2239 1067 2243 1071
rect 2391 1067 2395 1071
rect 2543 1067 2547 1071
rect 2695 1067 2699 1071
rect 2847 1067 2851 1071
rect 2999 1067 3003 1071
rect 3159 1067 3163 1071
rect 3327 1067 3331 1071
rect 3487 1067 3491 1071
rect 135 1055 139 1059
rect 271 1055 275 1059
rect 431 1055 435 1059
rect 583 1055 587 1059
rect 735 1055 739 1059
rect 887 1055 891 1059
rect 1047 1055 1051 1059
rect 1215 1055 1219 1059
rect 1383 1055 1387 1059
rect 1559 1055 1563 1059
rect 1727 1055 1731 1059
rect 111 1045 115 1049
rect 1823 1045 1827 1049
rect 111 1028 115 1032
rect 1823 1028 1827 1032
rect 1919 1021 1923 1025
rect 2127 1021 2131 1025
rect 2327 1021 2331 1025
rect 2519 1021 2523 1025
rect 2695 1021 2699 1025
rect 2863 1021 2867 1025
rect 3023 1021 3027 1025
rect 3183 1021 3187 1025
rect 3343 1021 3347 1025
rect 3487 1021 3491 1025
rect 143 1015 147 1019
rect 279 1015 283 1019
rect 439 1015 443 1019
rect 591 1015 595 1019
rect 743 1015 747 1019
rect 895 1015 899 1019
rect 1055 1015 1059 1019
rect 1223 1015 1227 1019
rect 1391 1015 1395 1019
rect 1567 1015 1571 1019
rect 1735 1015 1739 1019
rect 1863 1008 1867 1012
rect 3575 1008 3579 1012
rect 1863 991 1867 995
rect 3575 991 3579 995
rect 143 977 147 981
rect 287 977 291 981
rect 463 977 467 981
rect 647 977 651 981
rect 823 977 827 981
rect 999 977 1003 981
rect 1167 977 1171 981
rect 1327 977 1331 981
rect 1487 977 1491 981
rect 1655 977 1659 981
rect 1911 981 1915 985
rect 2119 981 2123 985
rect 2319 981 2323 985
rect 2511 981 2515 985
rect 2687 981 2691 985
rect 2855 981 2859 985
rect 3015 981 3019 985
rect 3175 981 3179 985
rect 3335 981 3339 985
rect 3479 981 3483 985
rect 111 964 115 968
rect 1823 964 1827 968
rect 1887 955 1891 959
rect 2071 955 2075 959
rect 2263 955 2267 959
rect 2455 955 2459 959
rect 2631 955 2635 959
rect 2799 955 2803 959
rect 2951 955 2955 959
rect 3095 955 3099 959
rect 3231 955 3235 959
rect 3367 955 3371 959
rect 3479 955 3483 959
rect 111 947 115 951
rect 1823 947 1827 951
rect 1863 945 1867 949
rect 3575 945 3579 949
rect 135 937 139 941
rect 279 937 283 941
rect 455 937 459 941
rect 639 937 643 941
rect 815 937 819 941
rect 991 937 995 941
rect 1159 937 1163 941
rect 1319 937 1323 941
rect 1479 937 1483 941
rect 1647 937 1651 941
rect 1863 928 1867 932
rect 3575 928 3579 932
rect 1895 915 1899 919
rect 2079 915 2083 919
rect 2271 915 2275 919
rect 2463 915 2467 919
rect 2639 915 2643 919
rect 2807 915 2811 919
rect 2959 915 2963 919
rect 3103 915 3107 919
rect 3239 915 3243 919
rect 3375 915 3379 919
rect 3487 915 3491 919
rect 135 907 139 911
rect 271 907 275 911
rect 439 907 443 911
rect 607 907 611 911
rect 775 907 779 911
rect 935 907 939 911
rect 1095 907 1099 911
rect 1247 907 1251 911
rect 1399 907 1403 911
rect 1551 907 1555 911
rect 111 897 115 901
rect 1823 897 1827 901
rect 111 880 115 884
rect 1823 880 1827 884
rect 1895 873 1899 877
rect 2023 873 2027 877
rect 2183 873 2187 877
rect 2351 873 2355 877
rect 2519 873 2523 877
rect 2687 873 2691 877
rect 2839 873 2843 877
rect 2983 873 2987 877
rect 3119 873 3123 877
rect 3247 873 3251 877
rect 3375 873 3379 877
rect 3487 873 3491 877
rect 143 867 147 871
rect 279 867 283 871
rect 447 867 451 871
rect 615 867 619 871
rect 783 867 787 871
rect 943 867 947 871
rect 1103 867 1107 871
rect 1255 867 1259 871
rect 1407 867 1411 871
rect 1559 867 1563 871
rect 1863 860 1867 864
rect 3575 860 3579 864
rect 1863 843 1867 847
rect 3575 843 3579 847
rect 143 833 147 837
rect 287 833 291 837
rect 463 833 467 837
rect 639 833 643 837
rect 807 833 811 837
rect 983 833 987 837
rect 1159 833 1163 837
rect 1335 833 1339 837
rect 1511 833 1515 837
rect 1887 833 1891 837
rect 2015 833 2019 837
rect 2175 833 2179 837
rect 2343 833 2347 837
rect 2511 833 2515 837
rect 2679 833 2683 837
rect 2831 833 2835 837
rect 2975 833 2979 837
rect 3111 833 3115 837
rect 3239 833 3243 837
rect 3367 833 3371 837
rect 3479 833 3483 837
rect 111 820 115 824
rect 1823 820 1827 824
rect 111 803 115 807
rect 1823 803 1827 807
rect 1887 803 1891 807
rect 2071 803 2075 807
rect 2263 803 2267 807
rect 2447 803 2451 807
rect 2623 803 2627 807
rect 2791 803 2795 807
rect 2943 803 2947 807
rect 3087 803 3091 807
rect 3223 803 3227 807
rect 3359 803 3363 807
rect 3479 803 3483 807
rect 135 793 139 797
rect 279 793 283 797
rect 455 793 459 797
rect 631 793 635 797
rect 799 793 803 797
rect 975 793 979 797
rect 1151 793 1155 797
rect 1327 793 1331 797
rect 1503 793 1507 797
rect 1863 793 1867 797
rect 3575 793 3579 797
rect 1863 776 1867 780
rect 3575 776 3579 780
rect 135 767 139 771
rect 271 767 275 771
rect 439 767 443 771
rect 607 767 611 771
rect 775 767 779 771
rect 935 767 939 771
rect 1087 767 1091 771
rect 1239 767 1243 771
rect 1391 767 1395 771
rect 1551 767 1555 771
rect 1895 763 1899 767
rect 2079 763 2083 767
rect 2271 763 2275 767
rect 2455 763 2459 767
rect 2631 763 2635 767
rect 2799 763 2803 767
rect 2951 763 2955 767
rect 3095 763 3099 767
rect 3231 763 3235 767
rect 3367 763 3371 767
rect 3487 763 3491 767
rect 111 757 115 761
rect 1823 757 1827 761
rect 111 740 115 744
rect 1823 740 1827 744
rect 143 727 147 731
rect 279 727 283 731
rect 447 727 451 731
rect 615 727 619 731
rect 783 727 787 731
rect 943 727 947 731
rect 1095 727 1099 731
rect 1247 727 1251 731
rect 1399 727 1403 731
rect 1559 727 1563 731
rect 1895 729 1899 733
rect 2071 729 2075 733
rect 2263 729 2267 733
rect 2447 729 2451 733
rect 2623 729 2627 733
rect 2799 729 2803 733
rect 2975 729 2979 733
rect 3151 729 3155 733
rect 3327 729 3331 733
rect 3487 729 3491 733
rect 1863 716 1867 720
rect 3575 716 3579 720
rect 1863 699 1867 703
rect 3575 699 3579 703
rect 143 689 147 693
rect 287 689 291 693
rect 455 689 459 693
rect 623 689 627 693
rect 791 689 795 693
rect 959 689 963 693
rect 1119 689 1123 693
rect 1279 689 1283 693
rect 1439 689 1443 693
rect 1599 689 1603 693
rect 1887 689 1891 693
rect 2063 689 2067 693
rect 2255 689 2259 693
rect 2439 689 2443 693
rect 2615 689 2619 693
rect 2791 689 2795 693
rect 2967 689 2971 693
rect 3143 689 3147 693
rect 3319 689 3323 693
rect 3479 689 3483 693
rect 111 676 115 680
rect 1823 676 1827 680
rect 111 659 115 663
rect 1823 659 1827 663
rect 1887 663 1891 667
rect 1975 663 1979 667
rect 2095 663 2099 667
rect 2223 663 2227 667
rect 2351 663 2355 667
rect 2479 663 2483 667
rect 2615 663 2619 667
rect 2767 663 2771 667
rect 2935 663 2939 667
rect 3119 663 3123 667
rect 3311 663 3315 667
rect 3479 663 3483 667
rect 135 649 139 653
rect 279 649 283 653
rect 447 649 451 653
rect 615 649 619 653
rect 783 649 787 653
rect 951 649 955 653
rect 1111 649 1115 653
rect 1271 649 1275 653
rect 1431 649 1435 653
rect 1591 649 1595 653
rect 1863 653 1867 657
rect 3575 653 3579 657
rect 1863 636 1867 640
rect 3575 636 3579 640
rect 135 619 139 623
rect 287 619 291 623
rect 455 619 459 623
rect 631 619 635 623
rect 799 619 803 623
rect 967 619 971 623
rect 1119 619 1123 623
rect 1271 619 1275 623
rect 1415 619 1419 623
rect 1559 619 1563 623
rect 1711 619 1715 623
rect 1895 623 1899 627
rect 1983 623 1987 627
rect 2103 623 2107 627
rect 2231 623 2235 627
rect 2359 623 2363 627
rect 2487 623 2491 627
rect 2623 623 2627 627
rect 2775 623 2779 627
rect 2943 623 2947 627
rect 3127 623 3131 627
rect 3319 623 3323 627
rect 3487 623 3491 627
rect 111 609 115 613
rect 1823 609 1827 613
rect 111 592 115 596
rect 1823 592 1827 596
rect 1895 585 1899 589
rect 2047 585 2051 589
rect 2215 585 2219 589
rect 2391 585 2395 589
rect 2583 585 2587 589
rect 2799 585 2803 589
rect 3023 585 3027 589
rect 3255 585 3259 589
rect 3487 585 3491 589
rect 143 579 147 583
rect 295 579 299 583
rect 463 579 467 583
rect 639 579 643 583
rect 807 579 811 583
rect 975 579 979 583
rect 1127 579 1131 583
rect 1279 579 1283 583
rect 1423 579 1427 583
rect 1567 579 1571 583
rect 1719 579 1723 583
rect 1863 572 1867 576
rect 3575 572 3579 576
rect 1863 555 1867 559
rect 3575 555 3579 559
rect 151 541 155 545
rect 311 541 315 545
rect 471 541 475 545
rect 631 541 635 545
rect 783 541 787 545
rect 927 541 931 545
rect 1063 541 1067 545
rect 1191 541 1195 545
rect 1311 541 1315 545
rect 1423 541 1427 545
rect 1535 541 1539 545
rect 1647 541 1651 545
rect 1735 541 1739 545
rect 1887 545 1891 549
rect 2039 545 2043 549
rect 2207 545 2211 549
rect 2383 545 2387 549
rect 2575 545 2579 549
rect 2791 545 2795 549
rect 3015 545 3019 549
rect 3247 545 3251 549
rect 3479 545 3483 549
rect 111 528 115 532
rect 1823 528 1827 532
rect 111 511 115 515
rect 1823 511 1827 515
rect 2191 515 2195 519
rect 2279 515 2283 519
rect 2375 515 2379 519
rect 2487 515 2491 519
rect 2631 515 2635 519
rect 2807 515 2811 519
rect 3007 515 3011 519
rect 3215 515 3219 519
rect 3431 515 3435 519
rect 143 501 147 505
rect 303 501 307 505
rect 463 501 467 505
rect 623 501 627 505
rect 775 501 779 505
rect 919 501 923 505
rect 1055 501 1059 505
rect 1183 501 1187 505
rect 1303 501 1307 505
rect 1415 501 1419 505
rect 1527 501 1531 505
rect 1639 501 1643 505
rect 1727 501 1731 505
rect 1863 505 1867 509
rect 3575 505 3579 509
rect 1863 488 1867 492
rect 3575 488 3579 492
rect 159 471 163 475
rect 311 471 315 475
rect 463 471 467 475
rect 615 471 619 475
rect 759 471 763 475
rect 887 471 891 475
rect 1007 471 1011 475
rect 1127 471 1131 475
rect 1239 471 1243 475
rect 1343 471 1347 475
rect 1439 471 1443 475
rect 1543 471 1547 475
rect 1639 471 1643 475
rect 1727 471 1731 475
rect 2199 475 2203 479
rect 2287 475 2291 479
rect 2383 475 2387 479
rect 2495 475 2499 479
rect 2639 475 2643 479
rect 2815 475 2819 479
rect 3015 475 3019 479
rect 3223 475 3227 479
rect 3439 475 3443 479
rect 111 461 115 465
rect 1823 461 1827 465
rect 111 444 115 448
rect 1823 444 1827 448
rect 167 431 171 435
rect 319 431 323 435
rect 471 431 475 435
rect 623 431 627 435
rect 767 431 771 435
rect 895 431 899 435
rect 1015 431 1019 435
rect 1135 431 1139 435
rect 1247 431 1251 435
rect 1351 431 1355 435
rect 1447 431 1451 435
rect 1551 431 1555 435
rect 1647 431 1651 435
rect 1735 431 1739 435
rect 1895 433 1899 437
rect 2039 433 2043 437
rect 2207 433 2211 437
rect 2383 433 2387 437
rect 2575 433 2579 437
rect 2783 433 2787 437
rect 3007 433 3011 437
rect 3239 433 3243 437
rect 3471 433 3475 437
rect 1863 420 1867 424
rect 3575 420 3579 424
rect 1863 403 1867 407
rect 3575 403 3579 407
rect 151 397 155 401
rect 271 397 275 401
rect 407 397 411 401
rect 551 397 555 401
rect 711 397 715 401
rect 887 397 891 401
rect 1063 397 1067 401
rect 1247 397 1251 401
rect 1439 397 1443 401
rect 1639 397 1643 401
rect 1887 393 1891 397
rect 2031 393 2035 397
rect 2199 393 2203 397
rect 2375 393 2379 397
rect 2567 393 2571 397
rect 2775 393 2779 397
rect 2999 393 3003 397
rect 3231 393 3235 397
rect 3463 393 3467 397
rect 111 384 115 388
rect 1823 384 1827 388
rect 111 367 115 371
rect 1823 367 1827 371
rect 1887 371 1891 375
rect 1975 371 1979 375
rect 2063 371 2067 375
rect 2151 371 2155 375
rect 2263 371 2267 375
rect 2383 371 2387 375
rect 2519 371 2523 375
rect 2671 371 2675 375
rect 2847 371 2851 375
rect 3031 371 3035 375
rect 3231 371 3235 375
rect 3431 371 3435 375
rect 143 357 147 361
rect 263 357 267 361
rect 399 357 403 361
rect 543 357 547 361
rect 703 357 707 361
rect 879 357 883 361
rect 1055 357 1059 361
rect 1239 357 1243 361
rect 1431 357 1435 361
rect 1631 357 1635 361
rect 1863 361 1867 365
rect 3575 361 3579 365
rect 1863 344 1867 348
rect 3575 344 3579 348
rect 1895 331 1899 335
rect 1983 331 1987 335
rect 2071 331 2075 335
rect 2159 331 2163 335
rect 2271 331 2275 335
rect 2391 331 2395 335
rect 2527 331 2531 335
rect 2679 331 2683 335
rect 2855 331 2859 335
rect 3039 331 3043 335
rect 3239 331 3243 335
rect 3439 331 3443 335
rect 135 319 139 323
rect 223 319 227 323
rect 311 319 315 323
rect 399 319 403 323
rect 487 319 491 323
rect 575 319 579 323
rect 663 319 667 323
rect 751 319 755 323
rect 839 319 843 323
rect 927 319 931 323
rect 1015 319 1019 323
rect 1103 319 1107 323
rect 1191 319 1195 323
rect 1287 319 1291 323
rect 1383 319 1387 323
rect 1479 319 1483 323
rect 1575 319 1579 323
rect 1671 319 1675 323
rect 111 309 115 313
rect 1823 309 1827 313
rect 1895 297 1899 301
rect 111 292 115 296
rect 1983 297 1987 301
rect 2071 297 2075 301
rect 2159 297 2163 301
rect 2247 297 2251 301
rect 2359 297 2363 301
rect 2471 297 2475 301
rect 2583 297 2587 301
rect 2695 297 2699 301
rect 2807 297 2811 301
rect 2919 297 2923 301
rect 3039 297 3043 301
rect 3159 297 3163 301
rect 1823 292 1827 296
rect 1863 284 1867 288
rect 143 279 147 283
rect 231 279 235 283
rect 319 279 323 283
rect 407 279 411 283
rect 495 279 499 283
rect 583 279 587 283
rect 671 279 675 283
rect 759 279 763 283
rect 847 279 851 283
rect 935 279 939 283
rect 1023 279 1027 283
rect 1111 279 1115 283
rect 1199 279 1203 283
rect 1295 279 1299 283
rect 1391 279 1395 283
rect 1487 279 1491 283
rect 1583 279 1587 283
rect 3575 284 3579 288
rect 1679 279 1683 283
rect 1863 267 1867 271
rect 3575 267 3579 271
rect 1887 257 1891 261
rect 1975 257 1979 261
rect 2063 257 2067 261
rect 2151 257 2155 261
rect 2239 257 2243 261
rect 2351 257 2355 261
rect 2463 257 2467 261
rect 2575 257 2579 261
rect 2687 257 2691 261
rect 2799 257 2803 261
rect 2911 257 2915 261
rect 3031 257 3035 261
rect 3151 257 3155 261
rect 143 241 147 245
rect 231 241 235 245
rect 319 241 323 245
rect 407 241 411 245
rect 495 241 499 245
rect 583 241 587 245
rect 671 241 675 245
rect 759 241 763 245
rect 847 241 851 245
rect 935 241 939 245
rect 1023 241 1027 245
rect 1111 241 1115 245
rect 1199 241 1203 245
rect 1287 241 1291 245
rect 1375 241 1379 245
rect 1463 241 1467 245
rect 1551 241 1555 245
rect 1639 241 1643 245
rect 1727 241 1731 245
rect 1887 235 1891 239
rect 1975 235 1979 239
rect 2063 235 2067 239
rect 2151 235 2155 239
rect 2263 235 2267 239
rect 2399 235 2403 239
rect 2535 235 2539 239
rect 2679 235 2683 239
rect 2815 235 2819 239
rect 2951 235 2955 239
rect 3087 235 3091 239
rect 3223 235 3227 239
rect 3359 235 3363 239
rect 3479 235 3483 239
rect 111 228 115 232
rect 1823 228 1827 232
rect 1863 225 1867 229
rect 3575 225 3579 229
rect 111 211 115 215
rect 1823 211 1827 215
rect 1863 208 1867 212
rect 3575 208 3579 212
rect 135 201 139 205
rect 223 201 227 205
rect 311 201 315 205
rect 399 201 403 205
rect 487 201 491 205
rect 575 201 579 205
rect 663 201 667 205
rect 751 201 755 205
rect 839 201 843 205
rect 927 201 931 205
rect 1015 201 1019 205
rect 1103 201 1107 205
rect 1191 201 1195 205
rect 1279 201 1283 205
rect 1367 201 1371 205
rect 1455 201 1459 205
rect 1543 201 1547 205
rect 1631 201 1635 205
rect 1719 201 1723 205
rect 1895 195 1899 199
rect 1983 195 1987 199
rect 2071 195 2075 199
rect 2159 195 2163 199
rect 2271 195 2275 199
rect 2407 195 2411 199
rect 2543 195 2547 199
rect 2687 195 2691 199
rect 2823 195 2827 199
rect 2959 195 2963 199
rect 3095 195 3099 199
rect 3231 195 3235 199
rect 3367 195 3371 199
rect 3487 195 3491 199
rect 2783 129 2787 133
rect 2871 129 2875 133
rect 2959 129 2963 133
rect 3047 129 3051 133
rect 3135 129 3139 133
rect 3223 129 3227 133
rect 3311 129 3315 133
rect 3399 129 3403 133
rect 3487 129 3491 133
rect 1863 116 1867 120
rect 3575 116 3579 120
rect 1863 99 1867 103
rect 3575 99 3579 103
rect 2775 89 2779 93
rect 2863 89 2867 93
rect 2951 89 2955 93
rect 3039 89 3043 93
rect 3127 89 3131 93
rect 3215 89 3219 93
rect 3303 89 3307 93
rect 3391 89 3395 93
rect 3479 89 3483 93
<< m3 >>
rect 111 3670 115 3671
rect 111 3665 115 3666
rect 135 3670 139 3671
rect 135 3665 139 3666
rect 223 3670 227 3671
rect 223 3665 227 3666
rect 1823 3670 1827 3671
rect 1823 3665 1827 3666
rect 112 3650 114 3665
rect 136 3660 138 3665
rect 224 3660 226 3665
rect 134 3659 140 3660
rect 134 3655 135 3659
rect 139 3655 140 3659
rect 134 3654 140 3655
rect 222 3659 228 3660
rect 222 3655 223 3659
rect 227 3655 228 3659
rect 222 3654 228 3655
rect 1824 3650 1826 3665
rect 110 3649 116 3650
rect 110 3645 111 3649
rect 115 3645 116 3649
rect 110 3644 116 3645
rect 1822 3649 1828 3650
rect 1822 3645 1823 3649
rect 1827 3645 1828 3649
rect 1822 3644 1828 3645
rect 110 3632 116 3633
rect 110 3628 111 3632
rect 115 3628 116 3632
rect 110 3627 116 3628
rect 1822 3632 1828 3633
rect 1822 3628 1823 3632
rect 1827 3628 1828 3632
rect 1822 3627 1828 3628
rect 112 3603 114 3627
rect 142 3619 148 3620
rect 142 3615 143 3619
rect 147 3615 148 3619
rect 142 3614 148 3615
rect 230 3619 236 3620
rect 230 3615 231 3619
rect 235 3615 236 3619
rect 230 3614 236 3615
rect 144 3603 146 3614
rect 232 3603 234 3614
rect 1824 3603 1826 3627
rect 111 3602 115 3603
rect 111 3597 115 3598
rect 143 3602 147 3603
rect 143 3597 147 3598
rect 231 3602 235 3603
rect 231 3597 235 3598
rect 319 3602 323 3603
rect 319 3597 323 3598
rect 407 3602 411 3603
rect 407 3597 411 3598
rect 495 3602 499 3603
rect 495 3597 499 3598
rect 1823 3602 1827 3603
rect 1823 3597 1827 3598
rect 112 3573 114 3597
rect 144 3586 146 3597
rect 232 3586 234 3597
rect 320 3586 322 3597
rect 408 3586 410 3597
rect 496 3586 498 3597
rect 142 3585 148 3586
rect 142 3581 143 3585
rect 147 3581 148 3585
rect 142 3580 148 3581
rect 230 3585 236 3586
rect 230 3581 231 3585
rect 235 3581 236 3585
rect 230 3580 236 3581
rect 318 3585 324 3586
rect 318 3581 319 3585
rect 323 3581 324 3585
rect 318 3580 324 3581
rect 406 3585 412 3586
rect 406 3581 407 3585
rect 411 3581 412 3585
rect 406 3580 412 3581
rect 494 3585 500 3586
rect 494 3581 495 3585
rect 499 3581 500 3585
rect 494 3580 500 3581
rect 1824 3573 1826 3597
rect 1863 3594 1867 3595
rect 1863 3589 1867 3590
rect 1887 3594 1891 3595
rect 1887 3589 1891 3590
rect 1975 3594 1979 3595
rect 1975 3589 1979 3590
rect 2063 3594 2067 3595
rect 2063 3589 2067 3590
rect 2151 3594 2155 3595
rect 2151 3589 2155 3590
rect 2239 3594 2243 3595
rect 2239 3589 2243 3590
rect 2327 3594 2331 3595
rect 2327 3589 2331 3590
rect 2431 3594 2435 3595
rect 2431 3589 2435 3590
rect 2535 3594 2539 3595
rect 2535 3589 2539 3590
rect 2631 3594 2635 3595
rect 2631 3589 2635 3590
rect 2727 3594 2731 3595
rect 2727 3589 2731 3590
rect 2823 3594 2827 3595
rect 2823 3589 2827 3590
rect 2919 3594 2923 3595
rect 2919 3589 2923 3590
rect 3015 3594 3019 3595
rect 3015 3589 3019 3590
rect 3119 3594 3123 3595
rect 3119 3589 3123 3590
rect 3223 3594 3227 3595
rect 3223 3589 3227 3590
rect 3575 3594 3579 3595
rect 3575 3589 3579 3590
rect 1864 3574 1866 3589
rect 1888 3584 1890 3589
rect 1976 3584 1978 3589
rect 2064 3584 2066 3589
rect 2152 3584 2154 3589
rect 2240 3584 2242 3589
rect 2328 3584 2330 3589
rect 2432 3584 2434 3589
rect 2536 3584 2538 3589
rect 2632 3584 2634 3589
rect 2728 3584 2730 3589
rect 2824 3584 2826 3589
rect 2920 3584 2922 3589
rect 3016 3584 3018 3589
rect 3120 3584 3122 3589
rect 3224 3584 3226 3589
rect 1886 3583 1892 3584
rect 1886 3579 1887 3583
rect 1891 3579 1892 3583
rect 1886 3578 1892 3579
rect 1974 3583 1980 3584
rect 1974 3579 1975 3583
rect 1979 3579 1980 3583
rect 1974 3578 1980 3579
rect 2062 3583 2068 3584
rect 2062 3579 2063 3583
rect 2067 3579 2068 3583
rect 2062 3578 2068 3579
rect 2150 3583 2156 3584
rect 2150 3579 2151 3583
rect 2155 3579 2156 3583
rect 2150 3578 2156 3579
rect 2238 3583 2244 3584
rect 2238 3579 2239 3583
rect 2243 3579 2244 3583
rect 2238 3578 2244 3579
rect 2326 3583 2332 3584
rect 2326 3579 2327 3583
rect 2331 3579 2332 3583
rect 2326 3578 2332 3579
rect 2430 3583 2436 3584
rect 2430 3579 2431 3583
rect 2435 3579 2436 3583
rect 2430 3578 2436 3579
rect 2534 3583 2540 3584
rect 2534 3579 2535 3583
rect 2539 3579 2540 3583
rect 2534 3578 2540 3579
rect 2630 3583 2636 3584
rect 2630 3579 2631 3583
rect 2635 3579 2636 3583
rect 2630 3578 2636 3579
rect 2726 3583 2732 3584
rect 2726 3579 2727 3583
rect 2731 3579 2732 3583
rect 2726 3578 2732 3579
rect 2822 3583 2828 3584
rect 2822 3579 2823 3583
rect 2827 3579 2828 3583
rect 2822 3578 2828 3579
rect 2918 3583 2924 3584
rect 2918 3579 2919 3583
rect 2923 3579 2924 3583
rect 2918 3578 2924 3579
rect 3014 3583 3020 3584
rect 3014 3579 3015 3583
rect 3019 3579 3020 3583
rect 3014 3578 3020 3579
rect 3118 3583 3124 3584
rect 3118 3579 3119 3583
rect 3123 3579 3124 3583
rect 3118 3578 3124 3579
rect 3222 3583 3228 3584
rect 3222 3579 3223 3583
rect 3227 3579 3228 3583
rect 3222 3578 3228 3579
rect 3576 3574 3578 3589
rect 1862 3573 1868 3574
rect 110 3572 116 3573
rect 110 3568 111 3572
rect 115 3568 116 3572
rect 110 3567 116 3568
rect 1822 3572 1828 3573
rect 1822 3568 1823 3572
rect 1827 3568 1828 3572
rect 1862 3569 1863 3573
rect 1867 3569 1868 3573
rect 1862 3568 1868 3569
rect 3574 3573 3580 3574
rect 3574 3569 3575 3573
rect 3579 3569 3580 3573
rect 3574 3568 3580 3569
rect 1822 3567 1828 3568
rect 1862 3556 1868 3557
rect 110 3555 116 3556
rect 110 3551 111 3555
rect 115 3551 116 3555
rect 110 3550 116 3551
rect 1822 3555 1828 3556
rect 1822 3551 1823 3555
rect 1827 3551 1828 3555
rect 1862 3552 1863 3556
rect 1867 3552 1868 3556
rect 1862 3551 1868 3552
rect 3574 3556 3580 3557
rect 3574 3552 3575 3556
rect 3579 3552 3580 3556
rect 3574 3551 3580 3552
rect 1822 3550 1828 3551
rect 112 3535 114 3550
rect 134 3545 140 3546
rect 134 3541 135 3545
rect 139 3541 140 3545
rect 134 3540 140 3541
rect 222 3545 228 3546
rect 222 3541 223 3545
rect 227 3541 228 3545
rect 222 3540 228 3541
rect 310 3545 316 3546
rect 310 3541 311 3545
rect 315 3541 316 3545
rect 310 3540 316 3541
rect 398 3545 404 3546
rect 398 3541 399 3545
rect 403 3541 404 3545
rect 398 3540 404 3541
rect 486 3545 492 3546
rect 486 3541 487 3545
rect 491 3541 492 3545
rect 486 3540 492 3541
rect 136 3535 138 3540
rect 224 3535 226 3540
rect 312 3535 314 3540
rect 400 3535 402 3540
rect 488 3535 490 3540
rect 1824 3535 1826 3550
rect 111 3534 115 3535
rect 111 3529 115 3530
rect 135 3534 139 3535
rect 135 3529 139 3530
rect 223 3534 227 3535
rect 223 3529 227 3530
rect 247 3534 251 3535
rect 247 3529 251 3530
rect 311 3534 315 3535
rect 311 3529 315 3530
rect 375 3534 379 3535
rect 375 3529 379 3530
rect 399 3534 403 3535
rect 399 3529 403 3530
rect 487 3534 491 3535
rect 487 3529 491 3530
rect 503 3534 507 3535
rect 503 3529 507 3530
rect 623 3534 627 3535
rect 623 3529 627 3530
rect 743 3534 747 3535
rect 743 3529 747 3530
rect 863 3534 867 3535
rect 863 3529 867 3530
rect 975 3534 979 3535
rect 975 3529 979 3530
rect 1079 3534 1083 3535
rect 1079 3529 1083 3530
rect 1175 3534 1179 3535
rect 1175 3529 1179 3530
rect 1271 3534 1275 3535
rect 1271 3529 1275 3530
rect 1367 3534 1371 3535
rect 1367 3529 1371 3530
rect 1471 3534 1475 3535
rect 1471 3529 1475 3530
rect 1575 3534 1579 3535
rect 1575 3529 1579 3530
rect 1823 3534 1827 3535
rect 1823 3529 1827 3530
rect 112 3514 114 3529
rect 248 3524 250 3529
rect 376 3524 378 3529
rect 504 3524 506 3529
rect 624 3524 626 3529
rect 744 3524 746 3529
rect 864 3524 866 3529
rect 976 3524 978 3529
rect 1080 3524 1082 3529
rect 1176 3524 1178 3529
rect 1272 3524 1274 3529
rect 1368 3524 1370 3529
rect 1472 3524 1474 3529
rect 1576 3524 1578 3529
rect 246 3523 252 3524
rect 246 3519 247 3523
rect 251 3519 252 3523
rect 246 3518 252 3519
rect 374 3523 380 3524
rect 374 3519 375 3523
rect 379 3519 380 3523
rect 374 3518 380 3519
rect 502 3523 508 3524
rect 502 3519 503 3523
rect 507 3519 508 3523
rect 502 3518 508 3519
rect 622 3523 628 3524
rect 622 3519 623 3523
rect 627 3519 628 3523
rect 622 3518 628 3519
rect 742 3523 748 3524
rect 742 3519 743 3523
rect 747 3519 748 3523
rect 742 3518 748 3519
rect 862 3523 868 3524
rect 862 3519 863 3523
rect 867 3519 868 3523
rect 862 3518 868 3519
rect 974 3523 980 3524
rect 974 3519 975 3523
rect 979 3519 980 3523
rect 974 3518 980 3519
rect 1078 3523 1084 3524
rect 1078 3519 1079 3523
rect 1083 3519 1084 3523
rect 1078 3518 1084 3519
rect 1174 3523 1180 3524
rect 1174 3519 1175 3523
rect 1179 3519 1180 3523
rect 1174 3518 1180 3519
rect 1270 3523 1276 3524
rect 1270 3519 1271 3523
rect 1275 3519 1276 3523
rect 1270 3518 1276 3519
rect 1366 3523 1372 3524
rect 1366 3519 1367 3523
rect 1371 3519 1372 3523
rect 1366 3518 1372 3519
rect 1470 3523 1476 3524
rect 1470 3519 1471 3523
rect 1475 3519 1476 3523
rect 1470 3518 1476 3519
rect 1574 3523 1580 3524
rect 1574 3519 1575 3523
rect 1579 3519 1580 3523
rect 1574 3518 1580 3519
rect 1824 3514 1826 3529
rect 1864 3527 1866 3551
rect 1894 3543 1900 3544
rect 1894 3539 1895 3543
rect 1899 3539 1900 3543
rect 1894 3538 1900 3539
rect 1982 3543 1988 3544
rect 1982 3539 1983 3543
rect 1987 3539 1988 3543
rect 1982 3538 1988 3539
rect 2070 3543 2076 3544
rect 2070 3539 2071 3543
rect 2075 3539 2076 3543
rect 2070 3538 2076 3539
rect 2158 3543 2164 3544
rect 2158 3539 2159 3543
rect 2163 3539 2164 3543
rect 2158 3538 2164 3539
rect 2246 3543 2252 3544
rect 2246 3539 2247 3543
rect 2251 3539 2252 3543
rect 2246 3538 2252 3539
rect 2334 3543 2340 3544
rect 2334 3539 2335 3543
rect 2339 3539 2340 3543
rect 2334 3538 2340 3539
rect 2438 3543 2444 3544
rect 2438 3539 2439 3543
rect 2443 3539 2444 3543
rect 2438 3538 2444 3539
rect 2542 3543 2548 3544
rect 2542 3539 2543 3543
rect 2547 3539 2548 3543
rect 2542 3538 2548 3539
rect 2638 3543 2644 3544
rect 2638 3539 2639 3543
rect 2643 3539 2644 3543
rect 2638 3538 2644 3539
rect 2734 3543 2740 3544
rect 2734 3539 2735 3543
rect 2739 3539 2740 3543
rect 2734 3538 2740 3539
rect 2830 3543 2836 3544
rect 2830 3539 2831 3543
rect 2835 3539 2836 3543
rect 2830 3538 2836 3539
rect 2926 3543 2932 3544
rect 2926 3539 2927 3543
rect 2931 3539 2932 3543
rect 2926 3538 2932 3539
rect 3022 3543 3028 3544
rect 3022 3539 3023 3543
rect 3027 3539 3028 3543
rect 3022 3538 3028 3539
rect 3126 3543 3132 3544
rect 3126 3539 3127 3543
rect 3131 3539 3132 3543
rect 3126 3538 3132 3539
rect 3230 3543 3236 3544
rect 3230 3539 3231 3543
rect 3235 3539 3236 3543
rect 3230 3538 3236 3539
rect 1896 3527 1898 3538
rect 1984 3527 1986 3538
rect 2072 3527 2074 3538
rect 2160 3527 2162 3538
rect 2248 3527 2250 3538
rect 2336 3527 2338 3538
rect 2440 3527 2442 3538
rect 2544 3527 2546 3538
rect 2640 3527 2642 3538
rect 2736 3527 2738 3538
rect 2832 3527 2834 3538
rect 2928 3527 2930 3538
rect 3024 3527 3026 3538
rect 3128 3527 3130 3538
rect 3232 3527 3234 3538
rect 3576 3527 3578 3551
rect 1863 3526 1867 3527
rect 1863 3521 1867 3522
rect 1895 3526 1899 3527
rect 1895 3521 1899 3522
rect 1983 3526 1987 3527
rect 1983 3521 1987 3522
rect 2071 3526 2075 3527
rect 2071 3521 2075 3522
rect 2103 3526 2107 3527
rect 2103 3521 2107 3522
rect 2159 3526 2163 3527
rect 2159 3521 2163 3522
rect 2231 3526 2235 3527
rect 2231 3521 2235 3522
rect 2247 3526 2251 3527
rect 2247 3521 2251 3522
rect 2335 3526 2339 3527
rect 2335 3521 2339 3522
rect 2367 3526 2371 3527
rect 2367 3521 2371 3522
rect 2439 3526 2443 3527
rect 2439 3521 2443 3522
rect 2511 3526 2515 3527
rect 2511 3521 2515 3522
rect 2543 3526 2547 3527
rect 2543 3521 2547 3522
rect 2639 3526 2643 3527
rect 2639 3521 2643 3522
rect 2655 3526 2659 3527
rect 2655 3521 2659 3522
rect 2735 3526 2739 3527
rect 2735 3521 2739 3522
rect 2791 3526 2795 3527
rect 2791 3521 2795 3522
rect 2831 3526 2835 3527
rect 2831 3521 2835 3522
rect 2927 3526 2931 3527
rect 2927 3521 2931 3522
rect 2935 3526 2939 3527
rect 2935 3521 2939 3522
rect 3023 3526 3027 3527
rect 3023 3521 3027 3522
rect 3079 3526 3083 3527
rect 3079 3521 3083 3522
rect 3127 3526 3131 3527
rect 3127 3521 3131 3522
rect 3223 3526 3227 3527
rect 3223 3521 3227 3522
rect 3231 3526 3235 3527
rect 3231 3521 3235 3522
rect 3575 3526 3579 3527
rect 3575 3521 3579 3522
rect 110 3513 116 3514
rect 110 3509 111 3513
rect 115 3509 116 3513
rect 110 3508 116 3509
rect 1822 3513 1828 3514
rect 1822 3509 1823 3513
rect 1827 3509 1828 3513
rect 1822 3508 1828 3509
rect 1864 3497 1866 3521
rect 1896 3510 1898 3521
rect 1984 3510 1986 3521
rect 2104 3510 2106 3521
rect 2232 3510 2234 3521
rect 2368 3510 2370 3521
rect 2512 3510 2514 3521
rect 2656 3510 2658 3521
rect 2792 3510 2794 3521
rect 2936 3510 2938 3521
rect 3080 3510 3082 3521
rect 3224 3510 3226 3521
rect 1894 3509 1900 3510
rect 1894 3505 1895 3509
rect 1899 3505 1900 3509
rect 1894 3504 1900 3505
rect 1982 3509 1988 3510
rect 1982 3505 1983 3509
rect 1987 3505 1988 3509
rect 1982 3504 1988 3505
rect 2102 3509 2108 3510
rect 2102 3505 2103 3509
rect 2107 3505 2108 3509
rect 2102 3504 2108 3505
rect 2230 3509 2236 3510
rect 2230 3505 2231 3509
rect 2235 3505 2236 3509
rect 2230 3504 2236 3505
rect 2366 3509 2372 3510
rect 2366 3505 2367 3509
rect 2371 3505 2372 3509
rect 2366 3504 2372 3505
rect 2510 3509 2516 3510
rect 2510 3505 2511 3509
rect 2515 3505 2516 3509
rect 2510 3504 2516 3505
rect 2654 3509 2660 3510
rect 2654 3505 2655 3509
rect 2659 3505 2660 3509
rect 2654 3504 2660 3505
rect 2790 3509 2796 3510
rect 2790 3505 2791 3509
rect 2795 3505 2796 3509
rect 2790 3504 2796 3505
rect 2934 3509 2940 3510
rect 2934 3505 2935 3509
rect 2939 3505 2940 3509
rect 2934 3504 2940 3505
rect 3078 3509 3084 3510
rect 3078 3505 3079 3509
rect 3083 3505 3084 3509
rect 3078 3504 3084 3505
rect 3222 3509 3228 3510
rect 3222 3505 3223 3509
rect 3227 3505 3228 3509
rect 3222 3504 3228 3505
rect 3576 3497 3578 3521
rect 110 3496 116 3497
rect 110 3492 111 3496
rect 115 3492 116 3496
rect 110 3491 116 3492
rect 1822 3496 1828 3497
rect 1822 3492 1823 3496
rect 1827 3492 1828 3496
rect 1822 3491 1828 3492
rect 1862 3496 1868 3497
rect 1862 3492 1863 3496
rect 1867 3492 1868 3496
rect 1862 3491 1868 3492
rect 3574 3496 3580 3497
rect 3574 3492 3575 3496
rect 3579 3492 3580 3496
rect 3574 3491 3580 3492
rect 112 3467 114 3491
rect 254 3483 260 3484
rect 254 3479 255 3483
rect 259 3479 260 3483
rect 254 3478 260 3479
rect 382 3483 388 3484
rect 382 3479 383 3483
rect 387 3479 388 3483
rect 382 3478 388 3479
rect 510 3483 516 3484
rect 510 3479 511 3483
rect 515 3479 516 3483
rect 510 3478 516 3479
rect 630 3483 636 3484
rect 630 3479 631 3483
rect 635 3479 636 3483
rect 630 3478 636 3479
rect 750 3483 756 3484
rect 750 3479 751 3483
rect 755 3479 756 3483
rect 750 3478 756 3479
rect 870 3483 876 3484
rect 870 3479 871 3483
rect 875 3479 876 3483
rect 870 3478 876 3479
rect 982 3483 988 3484
rect 982 3479 983 3483
rect 987 3479 988 3483
rect 982 3478 988 3479
rect 1086 3483 1092 3484
rect 1086 3479 1087 3483
rect 1091 3479 1092 3483
rect 1086 3478 1092 3479
rect 1182 3483 1188 3484
rect 1182 3479 1183 3483
rect 1187 3479 1188 3483
rect 1182 3478 1188 3479
rect 1278 3483 1284 3484
rect 1278 3479 1279 3483
rect 1283 3479 1284 3483
rect 1278 3478 1284 3479
rect 1374 3483 1380 3484
rect 1374 3479 1375 3483
rect 1379 3479 1380 3483
rect 1374 3478 1380 3479
rect 1478 3483 1484 3484
rect 1478 3479 1479 3483
rect 1483 3479 1484 3483
rect 1478 3478 1484 3479
rect 1582 3483 1588 3484
rect 1582 3479 1583 3483
rect 1587 3479 1588 3483
rect 1582 3478 1588 3479
rect 256 3467 258 3478
rect 384 3467 386 3478
rect 512 3467 514 3478
rect 632 3467 634 3478
rect 752 3467 754 3478
rect 872 3467 874 3478
rect 984 3467 986 3478
rect 1088 3467 1090 3478
rect 1184 3467 1186 3478
rect 1280 3467 1282 3478
rect 1376 3467 1378 3478
rect 1480 3467 1482 3478
rect 1584 3467 1586 3478
rect 1824 3467 1826 3491
rect 1862 3479 1868 3480
rect 1862 3475 1863 3479
rect 1867 3475 1868 3479
rect 1862 3474 1868 3475
rect 3574 3479 3580 3480
rect 3574 3475 3575 3479
rect 3579 3475 3580 3479
rect 3574 3474 3580 3475
rect 111 3466 115 3467
rect 111 3461 115 3462
rect 175 3466 179 3467
rect 175 3461 179 3462
rect 255 3466 259 3467
rect 255 3461 259 3462
rect 303 3466 307 3467
rect 303 3461 307 3462
rect 383 3466 387 3467
rect 383 3461 387 3462
rect 447 3466 451 3467
rect 447 3461 451 3462
rect 511 3466 515 3467
rect 511 3461 515 3462
rect 591 3466 595 3467
rect 591 3461 595 3462
rect 631 3466 635 3467
rect 631 3461 635 3462
rect 743 3466 747 3467
rect 743 3461 747 3462
rect 751 3466 755 3467
rect 751 3461 755 3462
rect 871 3466 875 3467
rect 871 3461 875 3462
rect 895 3466 899 3467
rect 895 3461 899 3462
rect 983 3466 987 3467
rect 983 3461 987 3462
rect 1039 3466 1043 3467
rect 1039 3461 1043 3462
rect 1087 3466 1091 3467
rect 1087 3461 1091 3462
rect 1183 3466 1187 3467
rect 1183 3461 1187 3462
rect 1279 3466 1283 3467
rect 1279 3461 1283 3462
rect 1327 3466 1331 3467
rect 1327 3461 1331 3462
rect 1375 3466 1379 3467
rect 1375 3461 1379 3462
rect 1479 3466 1483 3467
rect 1479 3461 1483 3462
rect 1583 3466 1587 3467
rect 1583 3461 1587 3462
rect 1823 3466 1827 3467
rect 1823 3461 1827 3462
rect 112 3437 114 3461
rect 176 3450 178 3461
rect 304 3450 306 3461
rect 448 3450 450 3461
rect 592 3450 594 3461
rect 744 3450 746 3461
rect 896 3450 898 3461
rect 1040 3450 1042 3461
rect 1184 3450 1186 3461
rect 1328 3450 1330 3461
rect 1480 3450 1482 3461
rect 174 3449 180 3450
rect 174 3445 175 3449
rect 179 3445 180 3449
rect 174 3444 180 3445
rect 302 3449 308 3450
rect 302 3445 303 3449
rect 307 3445 308 3449
rect 302 3444 308 3445
rect 446 3449 452 3450
rect 446 3445 447 3449
rect 451 3445 452 3449
rect 446 3444 452 3445
rect 590 3449 596 3450
rect 590 3445 591 3449
rect 595 3445 596 3449
rect 590 3444 596 3445
rect 742 3449 748 3450
rect 742 3445 743 3449
rect 747 3445 748 3449
rect 742 3444 748 3445
rect 894 3449 900 3450
rect 894 3445 895 3449
rect 899 3445 900 3449
rect 894 3444 900 3445
rect 1038 3449 1044 3450
rect 1038 3445 1039 3449
rect 1043 3445 1044 3449
rect 1038 3444 1044 3445
rect 1182 3449 1188 3450
rect 1182 3445 1183 3449
rect 1187 3445 1188 3449
rect 1182 3444 1188 3445
rect 1326 3449 1332 3450
rect 1326 3445 1327 3449
rect 1331 3445 1332 3449
rect 1326 3444 1332 3445
rect 1478 3449 1484 3450
rect 1478 3445 1479 3449
rect 1483 3445 1484 3449
rect 1478 3444 1484 3445
rect 1824 3437 1826 3461
rect 1864 3451 1866 3474
rect 1886 3469 1892 3470
rect 1886 3465 1887 3469
rect 1891 3465 1892 3469
rect 1886 3464 1892 3465
rect 1974 3469 1980 3470
rect 1974 3465 1975 3469
rect 1979 3465 1980 3469
rect 1974 3464 1980 3465
rect 2094 3469 2100 3470
rect 2094 3465 2095 3469
rect 2099 3465 2100 3469
rect 2094 3464 2100 3465
rect 2222 3469 2228 3470
rect 2222 3465 2223 3469
rect 2227 3465 2228 3469
rect 2222 3464 2228 3465
rect 2358 3469 2364 3470
rect 2358 3465 2359 3469
rect 2363 3465 2364 3469
rect 2358 3464 2364 3465
rect 2502 3469 2508 3470
rect 2502 3465 2503 3469
rect 2507 3465 2508 3469
rect 2502 3464 2508 3465
rect 2646 3469 2652 3470
rect 2646 3465 2647 3469
rect 2651 3465 2652 3469
rect 2646 3464 2652 3465
rect 2782 3469 2788 3470
rect 2782 3465 2783 3469
rect 2787 3465 2788 3469
rect 2782 3464 2788 3465
rect 2926 3469 2932 3470
rect 2926 3465 2927 3469
rect 2931 3465 2932 3469
rect 2926 3464 2932 3465
rect 3070 3469 3076 3470
rect 3070 3465 3071 3469
rect 3075 3465 3076 3469
rect 3070 3464 3076 3465
rect 3214 3469 3220 3470
rect 3214 3465 3215 3469
rect 3219 3465 3220 3469
rect 3214 3464 3220 3465
rect 1888 3451 1890 3464
rect 1976 3451 1978 3464
rect 2096 3451 2098 3464
rect 2224 3451 2226 3464
rect 2360 3451 2362 3464
rect 2504 3451 2506 3464
rect 2648 3451 2650 3464
rect 2784 3451 2786 3464
rect 2928 3451 2930 3464
rect 3072 3451 3074 3464
rect 3216 3451 3218 3464
rect 3576 3451 3578 3474
rect 1863 3450 1867 3451
rect 1863 3445 1867 3446
rect 1887 3450 1891 3451
rect 1887 3445 1891 3446
rect 1975 3450 1979 3451
rect 1975 3445 1979 3446
rect 2023 3450 2027 3451
rect 2023 3445 2027 3446
rect 2095 3450 2099 3451
rect 2095 3445 2099 3446
rect 2191 3450 2195 3451
rect 2191 3445 2195 3446
rect 2223 3450 2227 3451
rect 2223 3445 2227 3446
rect 2359 3450 2363 3451
rect 2359 3445 2363 3446
rect 2367 3450 2371 3451
rect 2367 3445 2371 3446
rect 2503 3450 2507 3451
rect 2503 3445 2507 3446
rect 2543 3450 2547 3451
rect 2543 3445 2547 3446
rect 2647 3450 2651 3451
rect 2647 3445 2651 3446
rect 2711 3450 2715 3451
rect 2711 3445 2715 3446
rect 2783 3450 2787 3451
rect 2783 3445 2787 3446
rect 2871 3450 2875 3451
rect 2871 3445 2875 3446
rect 2927 3450 2931 3451
rect 2927 3445 2931 3446
rect 3031 3450 3035 3451
rect 3031 3445 3035 3446
rect 3071 3450 3075 3451
rect 3071 3445 3075 3446
rect 3191 3450 3195 3451
rect 3191 3445 3195 3446
rect 3215 3450 3219 3451
rect 3215 3445 3219 3446
rect 3359 3450 3363 3451
rect 3359 3445 3363 3446
rect 3575 3450 3579 3451
rect 3575 3445 3579 3446
rect 110 3436 116 3437
rect 110 3432 111 3436
rect 115 3432 116 3436
rect 110 3431 116 3432
rect 1822 3436 1828 3437
rect 1822 3432 1823 3436
rect 1827 3432 1828 3436
rect 1822 3431 1828 3432
rect 1864 3430 1866 3445
rect 1888 3440 1890 3445
rect 2024 3440 2026 3445
rect 2192 3440 2194 3445
rect 2368 3440 2370 3445
rect 2544 3440 2546 3445
rect 2712 3440 2714 3445
rect 2872 3440 2874 3445
rect 3032 3440 3034 3445
rect 3192 3440 3194 3445
rect 3360 3440 3362 3445
rect 1886 3439 1892 3440
rect 1886 3435 1887 3439
rect 1891 3435 1892 3439
rect 1886 3434 1892 3435
rect 2022 3439 2028 3440
rect 2022 3435 2023 3439
rect 2027 3435 2028 3439
rect 2022 3434 2028 3435
rect 2190 3439 2196 3440
rect 2190 3435 2191 3439
rect 2195 3435 2196 3439
rect 2190 3434 2196 3435
rect 2366 3439 2372 3440
rect 2366 3435 2367 3439
rect 2371 3435 2372 3439
rect 2366 3434 2372 3435
rect 2542 3439 2548 3440
rect 2542 3435 2543 3439
rect 2547 3435 2548 3439
rect 2542 3434 2548 3435
rect 2710 3439 2716 3440
rect 2710 3435 2711 3439
rect 2715 3435 2716 3439
rect 2710 3434 2716 3435
rect 2870 3439 2876 3440
rect 2870 3435 2871 3439
rect 2875 3435 2876 3439
rect 2870 3434 2876 3435
rect 3030 3439 3036 3440
rect 3030 3435 3031 3439
rect 3035 3435 3036 3439
rect 3030 3434 3036 3435
rect 3190 3439 3196 3440
rect 3190 3435 3191 3439
rect 3195 3435 3196 3439
rect 3190 3434 3196 3435
rect 3358 3439 3364 3440
rect 3358 3435 3359 3439
rect 3363 3435 3364 3439
rect 3358 3434 3364 3435
rect 3576 3430 3578 3445
rect 1862 3429 1868 3430
rect 1862 3425 1863 3429
rect 1867 3425 1868 3429
rect 1862 3424 1868 3425
rect 3574 3429 3580 3430
rect 3574 3425 3575 3429
rect 3579 3425 3580 3429
rect 3574 3424 3580 3425
rect 110 3419 116 3420
rect 110 3415 111 3419
rect 115 3415 116 3419
rect 110 3414 116 3415
rect 1822 3419 1828 3420
rect 1822 3415 1823 3419
rect 1827 3415 1828 3419
rect 1822 3414 1828 3415
rect 112 3399 114 3414
rect 166 3409 172 3410
rect 166 3405 167 3409
rect 171 3405 172 3409
rect 166 3404 172 3405
rect 294 3409 300 3410
rect 294 3405 295 3409
rect 299 3405 300 3409
rect 294 3404 300 3405
rect 438 3409 444 3410
rect 438 3405 439 3409
rect 443 3405 444 3409
rect 438 3404 444 3405
rect 582 3409 588 3410
rect 582 3405 583 3409
rect 587 3405 588 3409
rect 582 3404 588 3405
rect 734 3409 740 3410
rect 734 3405 735 3409
rect 739 3405 740 3409
rect 734 3404 740 3405
rect 886 3409 892 3410
rect 886 3405 887 3409
rect 891 3405 892 3409
rect 886 3404 892 3405
rect 1030 3409 1036 3410
rect 1030 3405 1031 3409
rect 1035 3405 1036 3409
rect 1030 3404 1036 3405
rect 1174 3409 1180 3410
rect 1174 3405 1175 3409
rect 1179 3405 1180 3409
rect 1174 3404 1180 3405
rect 1318 3409 1324 3410
rect 1318 3405 1319 3409
rect 1323 3405 1324 3409
rect 1318 3404 1324 3405
rect 1470 3409 1476 3410
rect 1470 3405 1471 3409
rect 1475 3405 1476 3409
rect 1470 3404 1476 3405
rect 168 3399 170 3404
rect 296 3399 298 3404
rect 440 3399 442 3404
rect 584 3399 586 3404
rect 736 3399 738 3404
rect 888 3399 890 3404
rect 1032 3399 1034 3404
rect 1176 3399 1178 3404
rect 1320 3399 1322 3404
rect 1472 3399 1474 3404
rect 1824 3399 1826 3414
rect 1862 3412 1868 3413
rect 1862 3408 1863 3412
rect 1867 3408 1868 3412
rect 1862 3407 1868 3408
rect 3574 3412 3580 3413
rect 3574 3408 3575 3412
rect 3579 3408 3580 3412
rect 3574 3407 3580 3408
rect 111 3398 115 3399
rect 111 3393 115 3394
rect 135 3398 139 3399
rect 135 3393 139 3394
rect 167 3398 171 3399
rect 167 3393 171 3394
rect 263 3398 267 3399
rect 263 3393 267 3394
rect 295 3398 299 3399
rect 295 3393 299 3394
rect 407 3398 411 3399
rect 407 3393 411 3394
rect 439 3398 443 3399
rect 439 3393 443 3394
rect 567 3398 571 3399
rect 567 3393 571 3394
rect 583 3398 587 3399
rect 583 3393 587 3394
rect 727 3398 731 3399
rect 727 3393 731 3394
rect 735 3398 739 3399
rect 735 3393 739 3394
rect 887 3398 891 3399
rect 887 3393 891 3394
rect 1031 3398 1035 3399
rect 1031 3393 1035 3394
rect 1047 3398 1051 3399
rect 1047 3393 1051 3394
rect 1175 3398 1179 3399
rect 1175 3393 1179 3394
rect 1207 3398 1211 3399
rect 1207 3393 1211 3394
rect 1319 3398 1323 3399
rect 1319 3393 1323 3394
rect 1367 3398 1371 3399
rect 1367 3393 1371 3394
rect 1471 3398 1475 3399
rect 1471 3393 1475 3394
rect 1527 3398 1531 3399
rect 1527 3393 1531 3394
rect 1823 3398 1827 3399
rect 1823 3393 1827 3394
rect 112 3378 114 3393
rect 136 3388 138 3393
rect 264 3388 266 3393
rect 408 3388 410 3393
rect 568 3388 570 3393
rect 728 3388 730 3393
rect 888 3388 890 3393
rect 1048 3388 1050 3393
rect 1208 3388 1210 3393
rect 1368 3388 1370 3393
rect 1528 3388 1530 3393
rect 134 3387 140 3388
rect 134 3383 135 3387
rect 139 3383 140 3387
rect 134 3382 140 3383
rect 262 3387 268 3388
rect 262 3383 263 3387
rect 267 3383 268 3387
rect 262 3382 268 3383
rect 406 3387 412 3388
rect 406 3383 407 3387
rect 411 3383 412 3387
rect 406 3382 412 3383
rect 566 3387 572 3388
rect 566 3383 567 3387
rect 571 3383 572 3387
rect 566 3382 572 3383
rect 726 3387 732 3388
rect 726 3383 727 3387
rect 731 3383 732 3387
rect 726 3382 732 3383
rect 886 3387 892 3388
rect 886 3383 887 3387
rect 891 3383 892 3387
rect 886 3382 892 3383
rect 1046 3387 1052 3388
rect 1046 3383 1047 3387
rect 1051 3383 1052 3387
rect 1046 3382 1052 3383
rect 1206 3387 1212 3388
rect 1206 3383 1207 3387
rect 1211 3383 1212 3387
rect 1206 3382 1212 3383
rect 1366 3387 1372 3388
rect 1366 3383 1367 3387
rect 1371 3383 1372 3387
rect 1366 3382 1372 3383
rect 1526 3387 1532 3388
rect 1526 3383 1527 3387
rect 1531 3383 1532 3387
rect 1526 3382 1532 3383
rect 1824 3378 1826 3393
rect 110 3377 116 3378
rect 110 3373 111 3377
rect 115 3373 116 3377
rect 110 3372 116 3373
rect 1822 3377 1828 3378
rect 1822 3373 1823 3377
rect 1827 3373 1828 3377
rect 1864 3375 1866 3407
rect 1894 3399 1900 3400
rect 1894 3395 1895 3399
rect 1899 3395 1900 3399
rect 1894 3394 1900 3395
rect 2030 3399 2036 3400
rect 2030 3395 2031 3399
rect 2035 3395 2036 3399
rect 2030 3394 2036 3395
rect 2198 3399 2204 3400
rect 2198 3395 2199 3399
rect 2203 3395 2204 3399
rect 2198 3394 2204 3395
rect 2374 3399 2380 3400
rect 2374 3395 2375 3399
rect 2379 3395 2380 3399
rect 2374 3394 2380 3395
rect 2550 3399 2556 3400
rect 2550 3395 2551 3399
rect 2555 3395 2556 3399
rect 2550 3394 2556 3395
rect 2718 3399 2724 3400
rect 2718 3395 2719 3399
rect 2723 3395 2724 3399
rect 2718 3394 2724 3395
rect 2878 3399 2884 3400
rect 2878 3395 2879 3399
rect 2883 3395 2884 3399
rect 2878 3394 2884 3395
rect 3038 3399 3044 3400
rect 3038 3395 3039 3399
rect 3043 3395 3044 3399
rect 3038 3394 3044 3395
rect 3198 3399 3204 3400
rect 3198 3395 3199 3399
rect 3203 3395 3204 3399
rect 3198 3394 3204 3395
rect 3366 3399 3372 3400
rect 3366 3395 3367 3399
rect 3371 3395 3372 3399
rect 3366 3394 3372 3395
rect 1896 3375 1898 3394
rect 2032 3375 2034 3394
rect 2200 3375 2202 3394
rect 2376 3375 2378 3394
rect 2552 3375 2554 3394
rect 2720 3375 2722 3394
rect 2880 3375 2882 3394
rect 3040 3375 3042 3394
rect 3200 3375 3202 3394
rect 3368 3375 3370 3394
rect 3576 3375 3578 3407
rect 1822 3372 1828 3373
rect 1863 3374 1867 3375
rect 1863 3369 1867 3370
rect 1895 3374 1899 3375
rect 1895 3369 1899 3370
rect 2031 3374 2035 3375
rect 2031 3369 2035 3370
rect 2199 3374 2203 3375
rect 2199 3369 2203 3370
rect 2375 3374 2379 3375
rect 2375 3369 2379 3370
rect 2551 3374 2555 3375
rect 2551 3369 2555 3370
rect 2719 3374 2723 3375
rect 2719 3369 2723 3370
rect 2879 3374 2883 3375
rect 2879 3369 2883 3370
rect 3039 3374 3043 3375
rect 3039 3369 3043 3370
rect 3191 3374 3195 3375
rect 3191 3369 3195 3370
rect 3199 3374 3203 3375
rect 3199 3369 3203 3370
rect 3343 3374 3347 3375
rect 3343 3369 3347 3370
rect 3367 3374 3371 3375
rect 3367 3369 3371 3370
rect 3487 3374 3491 3375
rect 3487 3369 3491 3370
rect 3575 3374 3579 3375
rect 3575 3369 3579 3370
rect 110 3360 116 3361
rect 110 3356 111 3360
rect 115 3356 116 3360
rect 110 3355 116 3356
rect 1822 3360 1828 3361
rect 1822 3356 1823 3360
rect 1827 3356 1828 3360
rect 1822 3355 1828 3356
rect 112 3327 114 3355
rect 142 3347 148 3348
rect 142 3343 143 3347
rect 147 3343 148 3347
rect 142 3342 148 3343
rect 270 3347 276 3348
rect 270 3343 271 3347
rect 275 3343 276 3347
rect 270 3342 276 3343
rect 414 3347 420 3348
rect 414 3343 415 3347
rect 419 3343 420 3347
rect 414 3342 420 3343
rect 574 3347 580 3348
rect 574 3343 575 3347
rect 579 3343 580 3347
rect 574 3342 580 3343
rect 734 3347 740 3348
rect 734 3343 735 3347
rect 739 3343 740 3347
rect 734 3342 740 3343
rect 894 3347 900 3348
rect 894 3343 895 3347
rect 899 3343 900 3347
rect 894 3342 900 3343
rect 1054 3347 1060 3348
rect 1054 3343 1055 3347
rect 1059 3343 1060 3347
rect 1054 3342 1060 3343
rect 1214 3347 1220 3348
rect 1214 3343 1215 3347
rect 1219 3343 1220 3347
rect 1214 3342 1220 3343
rect 1374 3347 1380 3348
rect 1374 3343 1375 3347
rect 1379 3343 1380 3347
rect 1374 3342 1380 3343
rect 1534 3347 1540 3348
rect 1534 3343 1535 3347
rect 1539 3343 1540 3347
rect 1534 3342 1540 3343
rect 144 3327 146 3342
rect 272 3327 274 3342
rect 416 3327 418 3342
rect 576 3327 578 3342
rect 736 3327 738 3342
rect 896 3327 898 3342
rect 1056 3327 1058 3342
rect 1216 3327 1218 3342
rect 1376 3327 1378 3342
rect 1536 3327 1538 3342
rect 1824 3327 1826 3355
rect 1864 3345 1866 3369
rect 1896 3358 1898 3369
rect 2032 3358 2034 3369
rect 2200 3358 2202 3369
rect 2376 3358 2378 3369
rect 2552 3358 2554 3369
rect 2720 3358 2722 3369
rect 2880 3358 2882 3369
rect 3040 3358 3042 3369
rect 3192 3358 3194 3369
rect 3344 3358 3346 3369
rect 3488 3358 3490 3369
rect 1894 3357 1900 3358
rect 1894 3353 1895 3357
rect 1899 3353 1900 3357
rect 1894 3352 1900 3353
rect 2030 3357 2036 3358
rect 2030 3353 2031 3357
rect 2035 3353 2036 3357
rect 2030 3352 2036 3353
rect 2198 3357 2204 3358
rect 2198 3353 2199 3357
rect 2203 3353 2204 3357
rect 2198 3352 2204 3353
rect 2374 3357 2380 3358
rect 2374 3353 2375 3357
rect 2379 3353 2380 3357
rect 2374 3352 2380 3353
rect 2550 3357 2556 3358
rect 2550 3353 2551 3357
rect 2555 3353 2556 3357
rect 2550 3352 2556 3353
rect 2718 3357 2724 3358
rect 2718 3353 2719 3357
rect 2723 3353 2724 3357
rect 2718 3352 2724 3353
rect 2878 3357 2884 3358
rect 2878 3353 2879 3357
rect 2883 3353 2884 3357
rect 2878 3352 2884 3353
rect 3038 3357 3044 3358
rect 3038 3353 3039 3357
rect 3043 3353 3044 3357
rect 3038 3352 3044 3353
rect 3190 3357 3196 3358
rect 3190 3353 3191 3357
rect 3195 3353 3196 3357
rect 3190 3352 3196 3353
rect 3342 3357 3348 3358
rect 3342 3353 3343 3357
rect 3347 3353 3348 3357
rect 3342 3352 3348 3353
rect 3486 3357 3492 3358
rect 3486 3353 3487 3357
rect 3491 3353 3492 3357
rect 3486 3352 3492 3353
rect 3576 3345 3578 3369
rect 1862 3344 1868 3345
rect 1862 3340 1863 3344
rect 1867 3340 1868 3344
rect 1862 3339 1868 3340
rect 3574 3344 3580 3345
rect 3574 3340 3575 3344
rect 3579 3340 3580 3344
rect 3574 3339 3580 3340
rect 1862 3327 1868 3328
rect 111 3326 115 3327
rect 111 3321 115 3322
rect 143 3326 147 3327
rect 143 3321 147 3322
rect 207 3326 211 3327
rect 207 3321 211 3322
rect 271 3326 275 3327
rect 271 3321 275 3322
rect 335 3326 339 3327
rect 335 3321 339 3322
rect 415 3326 419 3327
rect 415 3321 419 3322
rect 479 3326 483 3327
rect 479 3321 483 3322
rect 575 3326 579 3327
rect 575 3321 579 3322
rect 639 3326 643 3327
rect 639 3321 643 3322
rect 735 3326 739 3327
rect 735 3321 739 3322
rect 807 3326 811 3327
rect 807 3321 811 3322
rect 895 3326 899 3327
rect 895 3321 899 3322
rect 983 3326 987 3327
rect 983 3321 987 3322
rect 1055 3326 1059 3327
rect 1055 3321 1059 3322
rect 1167 3326 1171 3327
rect 1167 3321 1171 3322
rect 1215 3326 1219 3327
rect 1215 3321 1219 3322
rect 1351 3326 1355 3327
rect 1351 3321 1355 3322
rect 1375 3326 1379 3327
rect 1375 3321 1379 3322
rect 1535 3326 1539 3327
rect 1535 3321 1539 3322
rect 1543 3326 1547 3327
rect 1543 3321 1547 3322
rect 1823 3326 1827 3327
rect 1862 3323 1863 3327
rect 1867 3323 1868 3327
rect 1862 3322 1868 3323
rect 3574 3327 3580 3328
rect 3574 3323 3575 3327
rect 3579 3323 3580 3327
rect 3574 3322 3580 3323
rect 1823 3321 1827 3322
rect 112 3297 114 3321
rect 208 3310 210 3321
rect 336 3310 338 3321
rect 480 3310 482 3321
rect 640 3310 642 3321
rect 808 3310 810 3321
rect 984 3310 986 3321
rect 1168 3310 1170 3321
rect 1352 3310 1354 3321
rect 1544 3310 1546 3321
rect 206 3309 212 3310
rect 206 3305 207 3309
rect 211 3305 212 3309
rect 206 3304 212 3305
rect 334 3309 340 3310
rect 334 3305 335 3309
rect 339 3305 340 3309
rect 334 3304 340 3305
rect 478 3309 484 3310
rect 478 3305 479 3309
rect 483 3305 484 3309
rect 478 3304 484 3305
rect 638 3309 644 3310
rect 638 3305 639 3309
rect 643 3305 644 3309
rect 638 3304 644 3305
rect 806 3309 812 3310
rect 806 3305 807 3309
rect 811 3305 812 3309
rect 806 3304 812 3305
rect 982 3309 988 3310
rect 982 3305 983 3309
rect 987 3305 988 3309
rect 982 3304 988 3305
rect 1166 3309 1172 3310
rect 1166 3305 1167 3309
rect 1171 3305 1172 3309
rect 1166 3304 1172 3305
rect 1350 3309 1356 3310
rect 1350 3305 1351 3309
rect 1355 3305 1356 3309
rect 1350 3304 1356 3305
rect 1542 3309 1548 3310
rect 1542 3305 1543 3309
rect 1547 3305 1548 3309
rect 1542 3304 1548 3305
rect 1824 3297 1826 3321
rect 1864 3307 1866 3322
rect 1886 3317 1892 3318
rect 1886 3313 1887 3317
rect 1891 3313 1892 3317
rect 1886 3312 1892 3313
rect 2022 3317 2028 3318
rect 2022 3313 2023 3317
rect 2027 3313 2028 3317
rect 2022 3312 2028 3313
rect 2190 3317 2196 3318
rect 2190 3313 2191 3317
rect 2195 3313 2196 3317
rect 2190 3312 2196 3313
rect 2366 3317 2372 3318
rect 2366 3313 2367 3317
rect 2371 3313 2372 3317
rect 2366 3312 2372 3313
rect 2542 3317 2548 3318
rect 2542 3313 2543 3317
rect 2547 3313 2548 3317
rect 2542 3312 2548 3313
rect 2710 3317 2716 3318
rect 2710 3313 2711 3317
rect 2715 3313 2716 3317
rect 2710 3312 2716 3313
rect 2870 3317 2876 3318
rect 2870 3313 2871 3317
rect 2875 3313 2876 3317
rect 2870 3312 2876 3313
rect 3030 3317 3036 3318
rect 3030 3313 3031 3317
rect 3035 3313 3036 3317
rect 3030 3312 3036 3313
rect 3182 3317 3188 3318
rect 3182 3313 3183 3317
rect 3187 3313 3188 3317
rect 3182 3312 3188 3313
rect 3334 3317 3340 3318
rect 3334 3313 3335 3317
rect 3339 3313 3340 3317
rect 3334 3312 3340 3313
rect 3478 3317 3484 3318
rect 3478 3313 3479 3317
rect 3483 3313 3484 3317
rect 3478 3312 3484 3313
rect 1888 3307 1890 3312
rect 2024 3307 2026 3312
rect 2192 3307 2194 3312
rect 2368 3307 2370 3312
rect 2544 3307 2546 3312
rect 2712 3307 2714 3312
rect 2872 3307 2874 3312
rect 3032 3307 3034 3312
rect 3184 3307 3186 3312
rect 3336 3307 3338 3312
rect 3480 3307 3482 3312
rect 3576 3307 3578 3322
rect 1863 3306 1867 3307
rect 1863 3301 1867 3302
rect 1887 3306 1891 3307
rect 1887 3301 1891 3302
rect 2007 3306 2011 3307
rect 2007 3301 2011 3302
rect 2023 3306 2027 3307
rect 2023 3301 2027 3302
rect 2151 3306 2155 3307
rect 2151 3301 2155 3302
rect 2191 3306 2195 3307
rect 2191 3301 2195 3302
rect 2303 3306 2307 3307
rect 2303 3301 2307 3302
rect 2367 3306 2371 3307
rect 2367 3301 2371 3302
rect 2463 3306 2467 3307
rect 2463 3301 2467 3302
rect 2543 3306 2547 3307
rect 2543 3301 2547 3302
rect 2631 3306 2635 3307
rect 2631 3301 2635 3302
rect 2711 3306 2715 3307
rect 2711 3301 2715 3302
rect 2799 3306 2803 3307
rect 2799 3301 2803 3302
rect 2871 3306 2875 3307
rect 2871 3301 2875 3302
rect 2967 3306 2971 3307
rect 2967 3301 2971 3302
rect 3031 3306 3035 3307
rect 3031 3301 3035 3302
rect 3135 3306 3139 3307
rect 3135 3301 3139 3302
rect 3183 3306 3187 3307
rect 3183 3301 3187 3302
rect 3311 3306 3315 3307
rect 3311 3301 3315 3302
rect 3335 3306 3339 3307
rect 3335 3301 3339 3302
rect 3479 3306 3483 3307
rect 3479 3301 3483 3302
rect 3575 3306 3579 3307
rect 3575 3301 3579 3302
rect 110 3296 116 3297
rect 110 3292 111 3296
rect 115 3292 116 3296
rect 110 3291 116 3292
rect 1822 3296 1828 3297
rect 1822 3292 1823 3296
rect 1827 3292 1828 3296
rect 1822 3291 1828 3292
rect 1864 3286 1866 3301
rect 1888 3296 1890 3301
rect 2008 3296 2010 3301
rect 2152 3296 2154 3301
rect 2304 3296 2306 3301
rect 2464 3296 2466 3301
rect 2632 3296 2634 3301
rect 2800 3296 2802 3301
rect 2968 3296 2970 3301
rect 3136 3296 3138 3301
rect 3312 3296 3314 3301
rect 3480 3296 3482 3301
rect 1886 3295 1892 3296
rect 1886 3291 1887 3295
rect 1891 3291 1892 3295
rect 1886 3290 1892 3291
rect 2006 3295 2012 3296
rect 2006 3291 2007 3295
rect 2011 3291 2012 3295
rect 2006 3290 2012 3291
rect 2150 3295 2156 3296
rect 2150 3291 2151 3295
rect 2155 3291 2156 3295
rect 2150 3290 2156 3291
rect 2302 3295 2308 3296
rect 2302 3291 2303 3295
rect 2307 3291 2308 3295
rect 2302 3290 2308 3291
rect 2462 3295 2468 3296
rect 2462 3291 2463 3295
rect 2467 3291 2468 3295
rect 2462 3290 2468 3291
rect 2630 3295 2636 3296
rect 2630 3291 2631 3295
rect 2635 3291 2636 3295
rect 2630 3290 2636 3291
rect 2798 3295 2804 3296
rect 2798 3291 2799 3295
rect 2803 3291 2804 3295
rect 2798 3290 2804 3291
rect 2966 3295 2972 3296
rect 2966 3291 2967 3295
rect 2971 3291 2972 3295
rect 2966 3290 2972 3291
rect 3134 3295 3140 3296
rect 3134 3291 3135 3295
rect 3139 3291 3140 3295
rect 3134 3290 3140 3291
rect 3310 3295 3316 3296
rect 3310 3291 3311 3295
rect 3315 3291 3316 3295
rect 3310 3290 3316 3291
rect 3478 3295 3484 3296
rect 3478 3291 3479 3295
rect 3483 3291 3484 3295
rect 3478 3290 3484 3291
rect 3576 3286 3578 3301
rect 1862 3285 1868 3286
rect 1862 3281 1863 3285
rect 1867 3281 1868 3285
rect 1862 3280 1868 3281
rect 3574 3285 3580 3286
rect 3574 3281 3575 3285
rect 3579 3281 3580 3285
rect 3574 3280 3580 3281
rect 110 3279 116 3280
rect 110 3275 111 3279
rect 115 3275 116 3279
rect 110 3274 116 3275
rect 1822 3279 1828 3280
rect 1822 3275 1823 3279
rect 1827 3275 1828 3279
rect 1822 3274 1828 3275
rect 112 3255 114 3274
rect 198 3269 204 3270
rect 198 3265 199 3269
rect 203 3265 204 3269
rect 198 3264 204 3265
rect 326 3269 332 3270
rect 326 3265 327 3269
rect 331 3265 332 3269
rect 326 3264 332 3265
rect 470 3269 476 3270
rect 470 3265 471 3269
rect 475 3265 476 3269
rect 470 3264 476 3265
rect 630 3269 636 3270
rect 630 3265 631 3269
rect 635 3265 636 3269
rect 630 3264 636 3265
rect 798 3269 804 3270
rect 798 3265 799 3269
rect 803 3265 804 3269
rect 798 3264 804 3265
rect 974 3269 980 3270
rect 974 3265 975 3269
rect 979 3265 980 3269
rect 974 3264 980 3265
rect 1158 3269 1164 3270
rect 1158 3265 1159 3269
rect 1163 3265 1164 3269
rect 1158 3264 1164 3265
rect 1342 3269 1348 3270
rect 1342 3265 1343 3269
rect 1347 3265 1348 3269
rect 1342 3264 1348 3265
rect 1534 3269 1540 3270
rect 1534 3265 1535 3269
rect 1539 3265 1540 3269
rect 1534 3264 1540 3265
rect 200 3255 202 3264
rect 328 3255 330 3264
rect 472 3255 474 3264
rect 632 3255 634 3264
rect 800 3255 802 3264
rect 976 3255 978 3264
rect 1160 3255 1162 3264
rect 1344 3255 1346 3264
rect 1536 3255 1538 3264
rect 1824 3255 1826 3274
rect 1862 3268 1868 3269
rect 1862 3264 1863 3268
rect 1867 3264 1868 3268
rect 1862 3263 1868 3264
rect 3574 3268 3580 3269
rect 3574 3264 3575 3268
rect 3579 3264 3580 3268
rect 3574 3263 3580 3264
rect 111 3254 115 3255
rect 111 3249 115 3250
rect 199 3254 203 3255
rect 199 3249 203 3250
rect 327 3254 331 3255
rect 327 3249 331 3250
rect 367 3254 371 3255
rect 367 3249 371 3250
rect 471 3254 475 3255
rect 471 3249 475 3250
rect 503 3254 507 3255
rect 503 3249 507 3250
rect 631 3254 635 3255
rect 631 3249 635 3250
rect 639 3254 643 3255
rect 639 3249 643 3250
rect 783 3254 787 3255
rect 783 3249 787 3250
rect 799 3254 803 3255
rect 799 3249 803 3250
rect 935 3254 939 3255
rect 935 3249 939 3250
rect 975 3254 979 3255
rect 975 3249 979 3250
rect 1095 3254 1099 3255
rect 1095 3249 1099 3250
rect 1159 3254 1163 3255
rect 1159 3249 1163 3250
rect 1255 3254 1259 3255
rect 1255 3249 1259 3250
rect 1343 3254 1347 3255
rect 1343 3249 1347 3250
rect 1415 3254 1419 3255
rect 1415 3249 1419 3250
rect 1535 3254 1539 3255
rect 1535 3249 1539 3250
rect 1575 3254 1579 3255
rect 1575 3249 1579 3250
rect 1823 3254 1827 3255
rect 1823 3249 1827 3250
rect 112 3234 114 3249
rect 368 3244 370 3249
rect 504 3244 506 3249
rect 640 3244 642 3249
rect 784 3244 786 3249
rect 936 3244 938 3249
rect 1096 3244 1098 3249
rect 1256 3244 1258 3249
rect 1416 3244 1418 3249
rect 1576 3244 1578 3249
rect 366 3243 372 3244
rect 366 3239 367 3243
rect 371 3239 372 3243
rect 366 3238 372 3239
rect 502 3243 508 3244
rect 502 3239 503 3243
rect 507 3239 508 3243
rect 502 3238 508 3239
rect 638 3243 644 3244
rect 638 3239 639 3243
rect 643 3239 644 3243
rect 638 3238 644 3239
rect 782 3243 788 3244
rect 782 3239 783 3243
rect 787 3239 788 3243
rect 782 3238 788 3239
rect 934 3243 940 3244
rect 934 3239 935 3243
rect 939 3239 940 3243
rect 934 3238 940 3239
rect 1094 3243 1100 3244
rect 1094 3239 1095 3243
rect 1099 3239 1100 3243
rect 1094 3238 1100 3239
rect 1254 3243 1260 3244
rect 1254 3239 1255 3243
rect 1259 3239 1260 3243
rect 1254 3238 1260 3239
rect 1414 3243 1420 3244
rect 1414 3239 1415 3243
rect 1419 3239 1420 3243
rect 1414 3238 1420 3239
rect 1574 3243 1580 3244
rect 1574 3239 1575 3243
rect 1579 3239 1580 3243
rect 1574 3238 1580 3239
rect 1824 3234 1826 3249
rect 110 3233 116 3234
rect 110 3229 111 3233
rect 115 3229 116 3233
rect 110 3228 116 3229
rect 1822 3233 1828 3234
rect 1822 3229 1823 3233
rect 1827 3229 1828 3233
rect 1864 3231 1866 3263
rect 1894 3255 1900 3256
rect 1894 3251 1895 3255
rect 1899 3251 1900 3255
rect 1894 3250 1900 3251
rect 2014 3255 2020 3256
rect 2014 3251 2015 3255
rect 2019 3251 2020 3255
rect 2014 3250 2020 3251
rect 2158 3255 2164 3256
rect 2158 3251 2159 3255
rect 2163 3251 2164 3255
rect 2158 3250 2164 3251
rect 2310 3255 2316 3256
rect 2310 3251 2311 3255
rect 2315 3251 2316 3255
rect 2310 3250 2316 3251
rect 2470 3255 2476 3256
rect 2470 3251 2471 3255
rect 2475 3251 2476 3255
rect 2470 3250 2476 3251
rect 2638 3255 2644 3256
rect 2638 3251 2639 3255
rect 2643 3251 2644 3255
rect 2638 3250 2644 3251
rect 2806 3255 2812 3256
rect 2806 3251 2807 3255
rect 2811 3251 2812 3255
rect 2806 3250 2812 3251
rect 2974 3255 2980 3256
rect 2974 3251 2975 3255
rect 2979 3251 2980 3255
rect 2974 3250 2980 3251
rect 3142 3255 3148 3256
rect 3142 3251 3143 3255
rect 3147 3251 3148 3255
rect 3142 3250 3148 3251
rect 3318 3255 3324 3256
rect 3318 3251 3319 3255
rect 3323 3251 3324 3255
rect 3318 3250 3324 3251
rect 3486 3255 3492 3256
rect 3486 3251 3487 3255
rect 3491 3251 3492 3255
rect 3486 3250 3492 3251
rect 1896 3231 1898 3250
rect 2016 3231 2018 3250
rect 2160 3231 2162 3250
rect 2312 3231 2314 3250
rect 2472 3231 2474 3250
rect 2640 3231 2642 3250
rect 2808 3231 2810 3250
rect 2976 3231 2978 3250
rect 3144 3231 3146 3250
rect 3320 3231 3322 3250
rect 3488 3231 3490 3250
rect 3576 3231 3578 3263
rect 1822 3228 1828 3229
rect 1863 3230 1867 3231
rect 1863 3225 1867 3226
rect 1895 3230 1899 3231
rect 1895 3225 1899 3226
rect 2015 3230 2019 3231
rect 2015 3225 2019 3226
rect 2023 3230 2027 3231
rect 2023 3225 2027 3226
rect 2159 3230 2163 3231
rect 2159 3225 2163 3226
rect 2175 3230 2179 3231
rect 2175 3225 2179 3226
rect 2311 3230 2315 3231
rect 2311 3225 2315 3226
rect 2327 3230 2331 3231
rect 2327 3225 2331 3226
rect 2463 3230 2467 3231
rect 2463 3225 2467 3226
rect 2471 3230 2475 3231
rect 2471 3225 2475 3226
rect 2599 3230 2603 3231
rect 2599 3225 2603 3226
rect 2639 3230 2643 3231
rect 2639 3225 2643 3226
rect 2735 3230 2739 3231
rect 2735 3225 2739 3226
rect 2807 3230 2811 3231
rect 2807 3225 2811 3226
rect 2871 3230 2875 3231
rect 2871 3225 2875 3226
rect 2975 3230 2979 3231
rect 2975 3225 2979 3226
rect 3015 3230 3019 3231
rect 3015 3225 3019 3226
rect 3143 3230 3147 3231
rect 3143 3225 3147 3226
rect 3167 3230 3171 3231
rect 3167 3225 3171 3226
rect 3319 3230 3323 3231
rect 3319 3225 3323 3226
rect 3327 3230 3331 3231
rect 3327 3225 3331 3226
rect 3487 3230 3491 3231
rect 3487 3225 3491 3226
rect 3575 3230 3579 3231
rect 3575 3225 3579 3226
rect 110 3216 116 3217
rect 110 3212 111 3216
rect 115 3212 116 3216
rect 110 3211 116 3212
rect 1822 3216 1828 3217
rect 1822 3212 1823 3216
rect 1827 3212 1828 3216
rect 1822 3211 1828 3212
rect 112 3179 114 3211
rect 374 3203 380 3204
rect 374 3199 375 3203
rect 379 3199 380 3203
rect 374 3198 380 3199
rect 510 3203 516 3204
rect 510 3199 511 3203
rect 515 3199 516 3203
rect 510 3198 516 3199
rect 646 3203 652 3204
rect 646 3199 647 3203
rect 651 3199 652 3203
rect 646 3198 652 3199
rect 790 3203 796 3204
rect 790 3199 791 3203
rect 795 3199 796 3203
rect 790 3198 796 3199
rect 942 3203 948 3204
rect 942 3199 943 3203
rect 947 3199 948 3203
rect 942 3198 948 3199
rect 1102 3203 1108 3204
rect 1102 3199 1103 3203
rect 1107 3199 1108 3203
rect 1102 3198 1108 3199
rect 1262 3203 1268 3204
rect 1262 3199 1263 3203
rect 1267 3199 1268 3203
rect 1262 3198 1268 3199
rect 1422 3203 1428 3204
rect 1422 3199 1423 3203
rect 1427 3199 1428 3203
rect 1422 3198 1428 3199
rect 1582 3203 1588 3204
rect 1582 3199 1583 3203
rect 1587 3199 1588 3203
rect 1582 3198 1588 3199
rect 376 3179 378 3198
rect 512 3179 514 3198
rect 648 3179 650 3198
rect 792 3179 794 3198
rect 944 3179 946 3198
rect 1104 3179 1106 3198
rect 1264 3179 1266 3198
rect 1424 3179 1426 3198
rect 1584 3179 1586 3198
rect 1824 3179 1826 3211
rect 1864 3201 1866 3225
rect 1896 3214 1898 3225
rect 2024 3214 2026 3225
rect 2176 3214 2178 3225
rect 2328 3214 2330 3225
rect 2464 3214 2466 3225
rect 2600 3214 2602 3225
rect 2736 3214 2738 3225
rect 2872 3214 2874 3225
rect 3016 3214 3018 3225
rect 3168 3214 3170 3225
rect 3328 3214 3330 3225
rect 3488 3214 3490 3225
rect 1894 3213 1900 3214
rect 1894 3209 1895 3213
rect 1899 3209 1900 3213
rect 1894 3208 1900 3209
rect 2022 3213 2028 3214
rect 2022 3209 2023 3213
rect 2027 3209 2028 3213
rect 2022 3208 2028 3209
rect 2174 3213 2180 3214
rect 2174 3209 2175 3213
rect 2179 3209 2180 3213
rect 2174 3208 2180 3209
rect 2326 3213 2332 3214
rect 2326 3209 2327 3213
rect 2331 3209 2332 3213
rect 2326 3208 2332 3209
rect 2462 3213 2468 3214
rect 2462 3209 2463 3213
rect 2467 3209 2468 3213
rect 2462 3208 2468 3209
rect 2598 3213 2604 3214
rect 2598 3209 2599 3213
rect 2603 3209 2604 3213
rect 2598 3208 2604 3209
rect 2734 3213 2740 3214
rect 2734 3209 2735 3213
rect 2739 3209 2740 3213
rect 2734 3208 2740 3209
rect 2870 3213 2876 3214
rect 2870 3209 2871 3213
rect 2875 3209 2876 3213
rect 2870 3208 2876 3209
rect 3014 3213 3020 3214
rect 3014 3209 3015 3213
rect 3019 3209 3020 3213
rect 3014 3208 3020 3209
rect 3166 3213 3172 3214
rect 3166 3209 3167 3213
rect 3171 3209 3172 3213
rect 3166 3208 3172 3209
rect 3326 3213 3332 3214
rect 3326 3209 3327 3213
rect 3331 3209 3332 3213
rect 3326 3208 3332 3209
rect 3486 3213 3492 3214
rect 3486 3209 3487 3213
rect 3491 3209 3492 3213
rect 3486 3208 3492 3209
rect 3576 3201 3578 3225
rect 1862 3200 1868 3201
rect 1862 3196 1863 3200
rect 1867 3196 1868 3200
rect 1862 3195 1868 3196
rect 3574 3200 3580 3201
rect 3574 3196 3575 3200
rect 3579 3196 3580 3200
rect 3574 3195 3580 3196
rect 1862 3183 1868 3184
rect 1862 3179 1863 3183
rect 1867 3179 1868 3183
rect 111 3178 115 3179
rect 111 3173 115 3174
rect 375 3178 379 3179
rect 375 3173 379 3174
rect 447 3178 451 3179
rect 447 3173 451 3174
rect 511 3178 515 3179
rect 511 3173 515 3174
rect 559 3178 563 3179
rect 559 3173 563 3174
rect 647 3178 651 3179
rect 647 3173 651 3174
rect 687 3178 691 3179
rect 687 3173 691 3174
rect 791 3178 795 3179
rect 791 3173 795 3174
rect 823 3178 827 3179
rect 823 3173 827 3174
rect 943 3178 947 3179
rect 943 3173 947 3174
rect 975 3178 979 3179
rect 975 3173 979 3174
rect 1103 3178 1107 3179
rect 1103 3173 1107 3174
rect 1135 3178 1139 3179
rect 1135 3173 1139 3174
rect 1263 3178 1267 3179
rect 1263 3173 1267 3174
rect 1295 3178 1299 3179
rect 1295 3173 1299 3174
rect 1423 3178 1427 3179
rect 1423 3173 1427 3174
rect 1463 3178 1467 3179
rect 1463 3173 1467 3174
rect 1583 3178 1587 3179
rect 1583 3173 1587 3174
rect 1639 3178 1643 3179
rect 1639 3173 1643 3174
rect 1823 3178 1827 3179
rect 1862 3178 1868 3179
rect 3574 3183 3580 3184
rect 3574 3179 3575 3183
rect 3579 3179 3580 3183
rect 3574 3178 3580 3179
rect 1823 3173 1827 3174
rect 112 3149 114 3173
rect 448 3162 450 3173
rect 560 3162 562 3173
rect 688 3162 690 3173
rect 824 3162 826 3173
rect 976 3162 978 3173
rect 1136 3162 1138 3173
rect 1296 3162 1298 3173
rect 1464 3162 1466 3173
rect 1640 3162 1642 3173
rect 446 3161 452 3162
rect 446 3157 447 3161
rect 451 3157 452 3161
rect 446 3156 452 3157
rect 558 3161 564 3162
rect 558 3157 559 3161
rect 563 3157 564 3161
rect 558 3156 564 3157
rect 686 3161 692 3162
rect 686 3157 687 3161
rect 691 3157 692 3161
rect 686 3156 692 3157
rect 822 3161 828 3162
rect 822 3157 823 3161
rect 827 3157 828 3161
rect 822 3156 828 3157
rect 974 3161 980 3162
rect 974 3157 975 3161
rect 979 3157 980 3161
rect 974 3156 980 3157
rect 1134 3161 1140 3162
rect 1134 3157 1135 3161
rect 1139 3157 1140 3161
rect 1134 3156 1140 3157
rect 1294 3161 1300 3162
rect 1294 3157 1295 3161
rect 1299 3157 1300 3161
rect 1294 3156 1300 3157
rect 1462 3161 1468 3162
rect 1462 3157 1463 3161
rect 1467 3157 1468 3161
rect 1462 3156 1468 3157
rect 1638 3161 1644 3162
rect 1638 3157 1639 3161
rect 1643 3157 1644 3161
rect 1638 3156 1644 3157
rect 1824 3149 1826 3173
rect 1864 3159 1866 3178
rect 1886 3173 1892 3174
rect 1886 3169 1887 3173
rect 1891 3169 1892 3173
rect 1886 3168 1892 3169
rect 2014 3173 2020 3174
rect 2014 3169 2015 3173
rect 2019 3169 2020 3173
rect 2014 3168 2020 3169
rect 2166 3173 2172 3174
rect 2166 3169 2167 3173
rect 2171 3169 2172 3173
rect 2166 3168 2172 3169
rect 2318 3173 2324 3174
rect 2318 3169 2319 3173
rect 2323 3169 2324 3173
rect 2318 3168 2324 3169
rect 2454 3173 2460 3174
rect 2454 3169 2455 3173
rect 2459 3169 2460 3173
rect 2454 3168 2460 3169
rect 2590 3173 2596 3174
rect 2590 3169 2591 3173
rect 2595 3169 2596 3173
rect 2590 3168 2596 3169
rect 2726 3173 2732 3174
rect 2726 3169 2727 3173
rect 2731 3169 2732 3173
rect 2726 3168 2732 3169
rect 2862 3173 2868 3174
rect 2862 3169 2863 3173
rect 2867 3169 2868 3173
rect 2862 3168 2868 3169
rect 3006 3173 3012 3174
rect 3006 3169 3007 3173
rect 3011 3169 3012 3173
rect 3006 3168 3012 3169
rect 3158 3173 3164 3174
rect 3158 3169 3159 3173
rect 3163 3169 3164 3173
rect 3158 3168 3164 3169
rect 3318 3173 3324 3174
rect 3318 3169 3319 3173
rect 3323 3169 3324 3173
rect 3318 3168 3324 3169
rect 3478 3173 3484 3174
rect 3478 3169 3479 3173
rect 3483 3169 3484 3173
rect 3478 3168 3484 3169
rect 1888 3159 1890 3168
rect 2016 3159 2018 3168
rect 2168 3159 2170 3168
rect 2320 3159 2322 3168
rect 2456 3159 2458 3168
rect 2592 3159 2594 3168
rect 2728 3159 2730 3168
rect 2864 3159 2866 3168
rect 3008 3159 3010 3168
rect 3160 3159 3162 3168
rect 3320 3159 3322 3168
rect 3480 3159 3482 3168
rect 3576 3159 3578 3178
rect 1863 3158 1867 3159
rect 1863 3153 1867 3154
rect 1887 3158 1891 3159
rect 1887 3153 1891 3154
rect 2015 3158 2019 3159
rect 2015 3153 2019 3154
rect 2047 3158 2051 3159
rect 2047 3153 2051 3154
rect 2167 3158 2171 3159
rect 2167 3153 2171 3154
rect 2199 3158 2203 3159
rect 2199 3153 2203 3154
rect 2319 3158 2323 3159
rect 2319 3153 2323 3154
rect 2351 3158 2355 3159
rect 2351 3153 2355 3154
rect 2455 3158 2459 3159
rect 2455 3153 2459 3154
rect 2511 3158 2515 3159
rect 2511 3153 2515 3154
rect 2591 3158 2595 3159
rect 2591 3153 2595 3154
rect 2679 3158 2683 3159
rect 2679 3153 2683 3154
rect 2727 3158 2731 3159
rect 2727 3153 2731 3154
rect 2863 3158 2867 3159
rect 2863 3153 2867 3154
rect 2871 3158 2875 3159
rect 2871 3153 2875 3154
rect 3007 3158 3011 3159
rect 3007 3153 3011 3154
rect 3071 3158 3075 3159
rect 3071 3153 3075 3154
rect 3159 3158 3163 3159
rect 3159 3153 3163 3154
rect 3287 3158 3291 3159
rect 3287 3153 3291 3154
rect 3319 3158 3323 3159
rect 3319 3153 3323 3154
rect 3479 3158 3483 3159
rect 3479 3153 3483 3154
rect 3575 3158 3579 3159
rect 3575 3153 3579 3154
rect 110 3148 116 3149
rect 110 3144 111 3148
rect 115 3144 116 3148
rect 110 3143 116 3144
rect 1822 3148 1828 3149
rect 1822 3144 1823 3148
rect 1827 3144 1828 3148
rect 1822 3143 1828 3144
rect 1864 3138 1866 3153
rect 1888 3148 1890 3153
rect 2048 3148 2050 3153
rect 2200 3148 2202 3153
rect 2352 3148 2354 3153
rect 2512 3148 2514 3153
rect 2680 3148 2682 3153
rect 2872 3148 2874 3153
rect 3072 3148 3074 3153
rect 3288 3148 3290 3153
rect 3480 3148 3482 3153
rect 1886 3147 1892 3148
rect 1886 3143 1887 3147
rect 1891 3143 1892 3147
rect 1886 3142 1892 3143
rect 2046 3147 2052 3148
rect 2046 3143 2047 3147
rect 2051 3143 2052 3147
rect 2046 3142 2052 3143
rect 2198 3147 2204 3148
rect 2198 3143 2199 3147
rect 2203 3143 2204 3147
rect 2198 3142 2204 3143
rect 2350 3147 2356 3148
rect 2350 3143 2351 3147
rect 2355 3143 2356 3147
rect 2350 3142 2356 3143
rect 2510 3147 2516 3148
rect 2510 3143 2511 3147
rect 2515 3143 2516 3147
rect 2510 3142 2516 3143
rect 2678 3147 2684 3148
rect 2678 3143 2679 3147
rect 2683 3143 2684 3147
rect 2678 3142 2684 3143
rect 2870 3147 2876 3148
rect 2870 3143 2871 3147
rect 2875 3143 2876 3147
rect 2870 3142 2876 3143
rect 3070 3147 3076 3148
rect 3070 3143 3071 3147
rect 3075 3143 3076 3147
rect 3070 3142 3076 3143
rect 3286 3147 3292 3148
rect 3286 3143 3287 3147
rect 3291 3143 3292 3147
rect 3286 3142 3292 3143
rect 3478 3147 3484 3148
rect 3478 3143 3479 3147
rect 3483 3143 3484 3147
rect 3478 3142 3484 3143
rect 3576 3138 3578 3153
rect 1862 3137 1868 3138
rect 1862 3133 1863 3137
rect 1867 3133 1868 3137
rect 1862 3132 1868 3133
rect 3574 3137 3580 3138
rect 3574 3133 3575 3137
rect 3579 3133 3580 3137
rect 3574 3132 3580 3133
rect 110 3131 116 3132
rect 110 3127 111 3131
rect 115 3127 116 3131
rect 110 3126 116 3127
rect 1822 3131 1828 3132
rect 1822 3127 1823 3131
rect 1827 3127 1828 3131
rect 1822 3126 1828 3127
rect 112 3103 114 3126
rect 438 3121 444 3122
rect 438 3117 439 3121
rect 443 3117 444 3121
rect 438 3116 444 3117
rect 550 3121 556 3122
rect 550 3117 551 3121
rect 555 3117 556 3121
rect 550 3116 556 3117
rect 678 3121 684 3122
rect 678 3117 679 3121
rect 683 3117 684 3121
rect 678 3116 684 3117
rect 814 3121 820 3122
rect 814 3117 815 3121
rect 819 3117 820 3121
rect 814 3116 820 3117
rect 966 3121 972 3122
rect 966 3117 967 3121
rect 971 3117 972 3121
rect 966 3116 972 3117
rect 1126 3121 1132 3122
rect 1126 3117 1127 3121
rect 1131 3117 1132 3121
rect 1126 3116 1132 3117
rect 1286 3121 1292 3122
rect 1286 3117 1287 3121
rect 1291 3117 1292 3121
rect 1286 3116 1292 3117
rect 1454 3121 1460 3122
rect 1454 3117 1455 3121
rect 1459 3117 1460 3121
rect 1454 3116 1460 3117
rect 1630 3121 1636 3122
rect 1630 3117 1631 3121
rect 1635 3117 1636 3121
rect 1630 3116 1636 3117
rect 440 3103 442 3116
rect 552 3103 554 3116
rect 680 3103 682 3116
rect 816 3103 818 3116
rect 968 3103 970 3116
rect 1128 3103 1130 3116
rect 1288 3103 1290 3116
rect 1456 3103 1458 3116
rect 1632 3103 1634 3116
rect 1824 3103 1826 3126
rect 1862 3120 1868 3121
rect 1862 3116 1863 3120
rect 1867 3116 1868 3120
rect 1862 3115 1868 3116
rect 3574 3120 3580 3121
rect 3574 3116 3575 3120
rect 3579 3116 3580 3120
rect 3574 3115 3580 3116
rect 111 3102 115 3103
rect 111 3097 115 3098
rect 439 3102 443 3103
rect 439 3097 443 3098
rect 551 3102 555 3103
rect 551 3097 555 3098
rect 663 3102 667 3103
rect 663 3097 667 3098
rect 679 3102 683 3103
rect 679 3097 683 3098
rect 783 3102 787 3103
rect 783 3097 787 3098
rect 815 3102 819 3103
rect 815 3097 819 3098
rect 903 3102 907 3103
rect 903 3097 907 3098
rect 967 3102 971 3103
rect 967 3097 971 3098
rect 1031 3102 1035 3103
rect 1031 3097 1035 3098
rect 1127 3102 1131 3103
rect 1127 3097 1131 3098
rect 1159 3102 1163 3103
rect 1159 3097 1163 3098
rect 1287 3102 1291 3103
rect 1287 3097 1291 3098
rect 1423 3102 1427 3103
rect 1423 3097 1427 3098
rect 1455 3102 1459 3103
rect 1455 3097 1459 3098
rect 1559 3102 1563 3103
rect 1559 3097 1563 3098
rect 1631 3102 1635 3103
rect 1631 3097 1635 3098
rect 1695 3102 1699 3103
rect 1695 3097 1699 3098
rect 1823 3102 1827 3103
rect 1823 3097 1827 3098
rect 112 3082 114 3097
rect 552 3092 554 3097
rect 664 3092 666 3097
rect 784 3092 786 3097
rect 904 3092 906 3097
rect 1032 3092 1034 3097
rect 1160 3092 1162 3097
rect 1288 3092 1290 3097
rect 1424 3092 1426 3097
rect 1560 3092 1562 3097
rect 1696 3092 1698 3097
rect 550 3091 556 3092
rect 550 3087 551 3091
rect 555 3087 556 3091
rect 550 3086 556 3087
rect 662 3091 668 3092
rect 662 3087 663 3091
rect 667 3087 668 3091
rect 662 3086 668 3087
rect 782 3091 788 3092
rect 782 3087 783 3091
rect 787 3087 788 3091
rect 782 3086 788 3087
rect 902 3091 908 3092
rect 902 3087 903 3091
rect 907 3087 908 3091
rect 902 3086 908 3087
rect 1030 3091 1036 3092
rect 1030 3087 1031 3091
rect 1035 3087 1036 3091
rect 1030 3086 1036 3087
rect 1158 3091 1164 3092
rect 1158 3087 1159 3091
rect 1163 3087 1164 3091
rect 1158 3086 1164 3087
rect 1286 3091 1292 3092
rect 1286 3087 1287 3091
rect 1291 3087 1292 3091
rect 1286 3086 1292 3087
rect 1422 3091 1428 3092
rect 1422 3087 1423 3091
rect 1427 3087 1428 3091
rect 1422 3086 1428 3087
rect 1558 3091 1564 3092
rect 1558 3087 1559 3091
rect 1563 3087 1564 3091
rect 1558 3086 1564 3087
rect 1694 3091 1700 3092
rect 1694 3087 1695 3091
rect 1699 3087 1700 3091
rect 1694 3086 1700 3087
rect 1824 3082 1826 3097
rect 1864 3083 1866 3115
rect 1894 3107 1900 3108
rect 1894 3103 1895 3107
rect 1899 3103 1900 3107
rect 1894 3102 1900 3103
rect 2054 3107 2060 3108
rect 2054 3103 2055 3107
rect 2059 3103 2060 3107
rect 2054 3102 2060 3103
rect 2206 3107 2212 3108
rect 2206 3103 2207 3107
rect 2211 3103 2212 3107
rect 2206 3102 2212 3103
rect 2358 3107 2364 3108
rect 2358 3103 2359 3107
rect 2363 3103 2364 3107
rect 2358 3102 2364 3103
rect 2518 3107 2524 3108
rect 2518 3103 2519 3107
rect 2523 3103 2524 3107
rect 2518 3102 2524 3103
rect 2686 3107 2692 3108
rect 2686 3103 2687 3107
rect 2691 3103 2692 3107
rect 2686 3102 2692 3103
rect 2878 3107 2884 3108
rect 2878 3103 2879 3107
rect 2883 3103 2884 3107
rect 2878 3102 2884 3103
rect 3078 3107 3084 3108
rect 3078 3103 3079 3107
rect 3083 3103 3084 3107
rect 3078 3102 3084 3103
rect 3294 3107 3300 3108
rect 3294 3103 3295 3107
rect 3299 3103 3300 3107
rect 3294 3102 3300 3103
rect 3486 3107 3492 3108
rect 3486 3103 3487 3107
rect 3491 3103 3492 3107
rect 3486 3102 3492 3103
rect 1896 3083 1898 3102
rect 2056 3083 2058 3102
rect 2208 3083 2210 3102
rect 2360 3083 2362 3102
rect 2520 3083 2522 3102
rect 2688 3083 2690 3102
rect 2880 3083 2882 3102
rect 3080 3083 3082 3102
rect 3296 3083 3298 3102
rect 3488 3083 3490 3102
rect 3576 3083 3578 3115
rect 1863 3082 1867 3083
rect 110 3081 116 3082
rect 110 3077 111 3081
rect 115 3077 116 3081
rect 110 3076 116 3077
rect 1822 3081 1828 3082
rect 1822 3077 1823 3081
rect 1827 3077 1828 3081
rect 1863 3077 1867 3078
rect 1895 3082 1899 3083
rect 1895 3077 1899 3078
rect 1919 3082 1923 3083
rect 1919 3077 1923 3078
rect 2055 3082 2059 3083
rect 2055 3077 2059 3078
rect 2087 3082 2091 3083
rect 2087 3077 2091 3078
rect 2207 3082 2211 3083
rect 2207 3077 2211 3078
rect 2279 3082 2283 3083
rect 2279 3077 2283 3078
rect 2359 3082 2363 3083
rect 2359 3077 2363 3078
rect 2487 3082 2491 3083
rect 2487 3077 2491 3078
rect 2519 3082 2523 3083
rect 2519 3077 2523 3078
rect 2687 3082 2691 3083
rect 2687 3077 2691 3078
rect 2719 3082 2723 3083
rect 2719 3077 2723 3078
rect 2879 3082 2883 3083
rect 2879 3077 2883 3078
rect 2975 3082 2979 3083
rect 2975 3077 2979 3078
rect 3079 3082 3083 3083
rect 3079 3077 3083 3078
rect 3239 3082 3243 3083
rect 3239 3077 3243 3078
rect 3295 3082 3299 3083
rect 3295 3077 3299 3078
rect 3487 3082 3491 3083
rect 3487 3077 3491 3078
rect 3575 3082 3579 3083
rect 3575 3077 3579 3078
rect 1822 3076 1828 3077
rect 110 3064 116 3065
rect 110 3060 111 3064
rect 115 3060 116 3064
rect 110 3059 116 3060
rect 1822 3064 1828 3065
rect 1822 3060 1823 3064
rect 1827 3060 1828 3064
rect 1822 3059 1828 3060
rect 112 3031 114 3059
rect 558 3051 564 3052
rect 558 3047 559 3051
rect 563 3047 564 3051
rect 558 3046 564 3047
rect 670 3051 676 3052
rect 670 3047 671 3051
rect 675 3047 676 3051
rect 670 3046 676 3047
rect 790 3051 796 3052
rect 790 3047 791 3051
rect 795 3047 796 3051
rect 790 3046 796 3047
rect 910 3051 916 3052
rect 910 3047 911 3051
rect 915 3047 916 3051
rect 910 3046 916 3047
rect 1038 3051 1044 3052
rect 1038 3047 1039 3051
rect 1043 3047 1044 3051
rect 1038 3046 1044 3047
rect 1166 3051 1172 3052
rect 1166 3047 1167 3051
rect 1171 3047 1172 3051
rect 1166 3046 1172 3047
rect 1294 3051 1300 3052
rect 1294 3047 1295 3051
rect 1299 3047 1300 3051
rect 1294 3046 1300 3047
rect 1430 3051 1436 3052
rect 1430 3047 1431 3051
rect 1435 3047 1436 3051
rect 1430 3046 1436 3047
rect 1566 3051 1572 3052
rect 1566 3047 1567 3051
rect 1571 3047 1572 3051
rect 1566 3046 1572 3047
rect 1702 3051 1708 3052
rect 1702 3047 1703 3051
rect 1707 3047 1708 3051
rect 1702 3046 1708 3047
rect 560 3031 562 3046
rect 672 3031 674 3046
rect 792 3031 794 3046
rect 912 3031 914 3046
rect 1040 3031 1042 3046
rect 1168 3031 1170 3046
rect 1296 3031 1298 3046
rect 1432 3031 1434 3046
rect 1568 3031 1570 3046
rect 1704 3031 1706 3046
rect 1824 3031 1826 3059
rect 1864 3053 1866 3077
rect 1920 3066 1922 3077
rect 2088 3066 2090 3077
rect 2280 3066 2282 3077
rect 2488 3066 2490 3077
rect 2720 3066 2722 3077
rect 2976 3066 2978 3077
rect 3240 3066 3242 3077
rect 3488 3066 3490 3077
rect 1918 3065 1924 3066
rect 1918 3061 1919 3065
rect 1923 3061 1924 3065
rect 1918 3060 1924 3061
rect 2086 3065 2092 3066
rect 2086 3061 2087 3065
rect 2091 3061 2092 3065
rect 2086 3060 2092 3061
rect 2278 3065 2284 3066
rect 2278 3061 2279 3065
rect 2283 3061 2284 3065
rect 2278 3060 2284 3061
rect 2486 3065 2492 3066
rect 2486 3061 2487 3065
rect 2491 3061 2492 3065
rect 2486 3060 2492 3061
rect 2718 3065 2724 3066
rect 2718 3061 2719 3065
rect 2723 3061 2724 3065
rect 2718 3060 2724 3061
rect 2974 3065 2980 3066
rect 2974 3061 2975 3065
rect 2979 3061 2980 3065
rect 2974 3060 2980 3061
rect 3238 3065 3244 3066
rect 3238 3061 3239 3065
rect 3243 3061 3244 3065
rect 3238 3060 3244 3061
rect 3486 3065 3492 3066
rect 3486 3061 3487 3065
rect 3491 3061 3492 3065
rect 3486 3060 3492 3061
rect 3576 3053 3578 3077
rect 1862 3052 1868 3053
rect 1862 3048 1863 3052
rect 1867 3048 1868 3052
rect 1862 3047 1868 3048
rect 3574 3052 3580 3053
rect 3574 3048 3575 3052
rect 3579 3048 3580 3052
rect 3574 3047 3580 3048
rect 1862 3035 1868 3036
rect 1862 3031 1863 3035
rect 1867 3031 1868 3035
rect 111 3030 115 3031
rect 111 3025 115 3026
rect 559 3030 563 3031
rect 559 3025 563 3026
rect 575 3030 579 3031
rect 575 3025 579 3026
rect 671 3030 675 3031
rect 671 3025 675 3026
rect 703 3030 707 3031
rect 703 3025 707 3026
rect 791 3030 795 3031
rect 791 3025 795 3026
rect 831 3030 835 3031
rect 831 3025 835 3026
rect 911 3030 915 3031
rect 911 3025 915 3026
rect 967 3030 971 3031
rect 967 3025 971 3026
rect 1039 3030 1043 3031
rect 1039 3025 1043 3026
rect 1103 3030 1107 3031
rect 1103 3025 1107 3026
rect 1167 3030 1171 3031
rect 1167 3025 1171 3026
rect 1239 3030 1243 3031
rect 1239 3025 1243 3026
rect 1295 3030 1299 3031
rect 1295 3025 1299 3026
rect 1367 3030 1371 3031
rect 1367 3025 1371 3026
rect 1431 3030 1435 3031
rect 1431 3025 1435 3026
rect 1495 3030 1499 3031
rect 1495 3025 1499 3026
rect 1567 3030 1571 3031
rect 1567 3025 1571 3026
rect 1623 3030 1627 3031
rect 1623 3025 1627 3026
rect 1703 3030 1707 3031
rect 1703 3025 1707 3026
rect 1735 3030 1739 3031
rect 1735 3025 1739 3026
rect 1823 3030 1827 3031
rect 1862 3030 1868 3031
rect 3574 3035 3580 3036
rect 3574 3031 3575 3035
rect 3579 3031 3580 3035
rect 3574 3030 3580 3031
rect 1823 3025 1827 3026
rect 112 3001 114 3025
rect 576 3014 578 3025
rect 704 3014 706 3025
rect 832 3014 834 3025
rect 968 3014 970 3025
rect 1104 3014 1106 3025
rect 1240 3014 1242 3025
rect 1368 3014 1370 3025
rect 1496 3014 1498 3025
rect 1624 3014 1626 3025
rect 1736 3014 1738 3025
rect 574 3013 580 3014
rect 574 3009 575 3013
rect 579 3009 580 3013
rect 574 3008 580 3009
rect 702 3013 708 3014
rect 702 3009 703 3013
rect 707 3009 708 3013
rect 702 3008 708 3009
rect 830 3013 836 3014
rect 830 3009 831 3013
rect 835 3009 836 3013
rect 830 3008 836 3009
rect 966 3013 972 3014
rect 966 3009 967 3013
rect 971 3009 972 3013
rect 966 3008 972 3009
rect 1102 3013 1108 3014
rect 1102 3009 1103 3013
rect 1107 3009 1108 3013
rect 1102 3008 1108 3009
rect 1238 3013 1244 3014
rect 1238 3009 1239 3013
rect 1243 3009 1244 3013
rect 1238 3008 1244 3009
rect 1366 3013 1372 3014
rect 1366 3009 1367 3013
rect 1371 3009 1372 3013
rect 1366 3008 1372 3009
rect 1494 3013 1500 3014
rect 1494 3009 1495 3013
rect 1499 3009 1500 3013
rect 1494 3008 1500 3009
rect 1622 3013 1628 3014
rect 1622 3009 1623 3013
rect 1627 3009 1628 3013
rect 1622 3008 1628 3009
rect 1734 3013 1740 3014
rect 1734 3009 1735 3013
rect 1739 3009 1740 3013
rect 1734 3008 1740 3009
rect 1824 3001 1826 3025
rect 1864 3011 1866 3030
rect 1910 3025 1916 3026
rect 1910 3021 1911 3025
rect 1915 3021 1916 3025
rect 1910 3020 1916 3021
rect 2078 3025 2084 3026
rect 2078 3021 2079 3025
rect 2083 3021 2084 3025
rect 2078 3020 2084 3021
rect 2270 3025 2276 3026
rect 2270 3021 2271 3025
rect 2275 3021 2276 3025
rect 2270 3020 2276 3021
rect 2478 3025 2484 3026
rect 2478 3021 2479 3025
rect 2483 3021 2484 3025
rect 2478 3020 2484 3021
rect 2710 3025 2716 3026
rect 2710 3021 2711 3025
rect 2715 3021 2716 3025
rect 2710 3020 2716 3021
rect 2966 3025 2972 3026
rect 2966 3021 2967 3025
rect 2971 3021 2972 3025
rect 2966 3020 2972 3021
rect 3230 3025 3236 3026
rect 3230 3021 3231 3025
rect 3235 3021 3236 3025
rect 3230 3020 3236 3021
rect 3478 3025 3484 3026
rect 3478 3021 3479 3025
rect 3483 3021 3484 3025
rect 3478 3020 3484 3021
rect 1912 3011 1914 3020
rect 2080 3011 2082 3020
rect 2272 3011 2274 3020
rect 2480 3011 2482 3020
rect 2712 3011 2714 3020
rect 2968 3011 2970 3020
rect 3232 3011 3234 3020
rect 3480 3011 3482 3020
rect 3576 3011 3578 3030
rect 1863 3010 1867 3011
rect 1863 3005 1867 3006
rect 1911 3010 1915 3011
rect 1911 3005 1915 3006
rect 2023 3010 2027 3011
rect 2023 3005 2027 3006
rect 2079 3010 2083 3011
rect 2079 3005 2083 3006
rect 2159 3010 2163 3011
rect 2159 3005 2163 3006
rect 2271 3010 2275 3011
rect 2271 3005 2275 3006
rect 2287 3010 2291 3011
rect 2287 3005 2291 3006
rect 2415 3010 2419 3011
rect 2415 3005 2419 3006
rect 2479 3010 2483 3011
rect 2479 3005 2483 3006
rect 2535 3010 2539 3011
rect 2535 3005 2539 3006
rect 2663 3010 2667 3011
rect 2663 3005 2667 3006
rect 2711 3010 2715 3011
rect 2711 3005 2715 3006
rect 2807 3010 2811 3011
rect 2807 3005 2811 3006
rect 2967 3010 2971 3011
rect 2967 3005 2971 3006
rect 3143 3010 3147 3011
rect 3143 3005 3147 3006
rect 3231 3010 3235 3011
rect 3231 3005 3235 3006
rect 3319 3010 3323 3011
rect 3319 3005 3323 3006
rect 3479 3010 3483 3011
rect 3479 3005 3483 3006
rect 3575 3010 3579 3011
rect 3575 3005 3579 3006
rect 110 3000 116 3001
rect 110 2996 111 3000
rect 115 2996 116 3000
rect 110 2995 116 2996
rect 1822 3000 1828 3001
rect 1822 2996 1823 3000
rect 1827 2996 1828 3000
rect 1822 2995 1828 2996
rect 1864 2990 1866 3005
rect 2024 3000 2026 3005
rect 2160 3000 2162 3005
rect 2288 3000 2290 3005
rect 2416 3000 2418 3005
rect 2536 3000 2538 3005
rect 2664 3000 2666 3005
rect 2808 3000 2810 3005
rect 2968 3000 2970 3005
rect 3144 3000 3146 3005
rect 3320 3000 3322 3005
rect 3480 3000 3482 3005
rect 2022 2999 2028 3000
rect 2022 2995 2023 2999
rect 2027 2995 2028 2999
rect 2022 2994 2028 2995
rect 2158 2999 2164 3000
rect 2158 2995 2159 2999
rect 2163 2995 2164 2999
rect 2158 2994 2164 2995
rect 2286 2999 2292 3000
rect 2286 2995 2287 2999
rect 2291 2995 2292 2999
rect 2286 2994 2292 2995
rect 2414 2999 2420 3000
rect 2414 2995 2415 2999
rect 2419 2995 2420 2999
rect 2414 2994 2420 2995
rect 2534 2999 2540 3000
rect 2534 2995 2535 2999
rect 2539 2995 2540 2999
rect 2534 2994 2540 2995
rect 2662 2999 2668 3000
rect 2662 2995 2663 2999
rect 2667 2995 2668 2999
rect 2662 2994 2668 2995
rect 2806 2999 2812 3000
rect 2806 2995 2807 2999
rect 2811 2995 2812 2999
rect 2806 2994 2812 2995
rect 2966 2999 2972 3000
rect 2966 2995 2967 2999
rect 2971 2995 2972 2999
rect 2966 2994 2972 2995
rect 3142 2999 3148 3000
rect 3142 2995 3143 2999
rect 3147 2995 3148 2999
rect 3142 2994 3148 2995
rect 3318 2999 3324 3000
rect 3318 2995 3319 2999
rect 3323 2995 3324 2999
rect 3318 2994 3324 2995
rect 3478 2999 3484 3000
rect 3478 2995 3479 2999
rect 3483 2995 3484 2999
rect 3478 2994 3484 2995
rect 3576 2990 3578 3005
rect 1862 2989 1868 2990
rect 1862 2985 1863 2989
rect 1867 2985 1868 2989
rect 1862 2984 1868 2985
rect 3574 2989 3580 2990
rect 3574 2985 3575 2989
rect 3579 2985 3580 2989
rect 3574 2984 3580 2985
rect 110 2983 116 2984
rect 110 2979 111 2983
rect 115 2979 116 2983
rect 110 2978 116 2979
rect 1822 2983 1828 2984
rect 1822 2979 1823 2983
rect 1827 2979 1828 2983
rect 1822 2978 1828 2979
rect 112 2963 114 2978
rect 566 2973 572 2974
rect 566 2969 567 2973
rect 571 2969 572 2973
rect 566 2968 572 2969
rect 694 2973 700 2974
rect 694 2969 695 2973
rect 699 2969 700 2973
rect 694 2968 700 2969
rect 822 2973 828 2974
rect 822 2969 823 2973
rect 827 2969 828 2973
rect 822 2968 828 2969
rect 958 2973 964 2974
rect 958 2969 959 2973
rect 963 2969 964 2973
rect 958 2968 964 2969
rect 1094 2973 1100 2974
rect 1094 2969 1095 2973
rect 1099 2969 1100 2973
rect 1094 2968 1100 2969
rect 1230 2973 1236 2974
rect 1230 2969 1231 2973
rect 1235 2969 1236 2973
rect 1230 2968 1236 2969
rect 1358 2973 1364 2974
rect 1358 2969 1359 2973
rect 1363 2969 1364 2973
rect 1358 2968 1364 2969
rect 1486 2973 1492 2974
rect 1486 2969 1487 2973
rect 1491 2969 1492 2973
rect 1486 2968 1492 2969
rect 1614 2973 1620 2974
rect 1614 2969 1615 2973
rect 1619 2969 1620 2973
rect 1614 2968 1620 2969
rect 1726 2973 1732 2974
rect 1726 2969 1727 2973
rect 1731 2969 1732 2973
rect 1726 2968 1732 2969
rect 568 2963 570 2968
rect 696 2963 698 2968
rect 824 2963 826 2968
rect 960 2963 962 2968
rect 1096 2963 1098 2968
rect 1232 2963 1234 2968
rect 1360 2963 1362 2968
rect 1488 2963 1490 2968
rect 1616 2963 1618 2968
rect 1728 2963 1730 2968
rect 1824 2963 1826 2978
rect 1862 2972 1868 2973
rect 1862 2968 1863 2972
rect 1867 2968 1868 2972
rect 1862 2967 1868 2968
rect 3574 2972 3580 2973
rect 3574 2968 3575 2972
rect 3579 2968 3580 2972
rect 3574 2967 3580 2968
rect 111 2962 115 2963
rect 111 2957 115 2958
rect 495 2962 499 2963
rect 495 2957 499 2958
rect 567 2962 571 2963
rect 567 2957 571 2958
rect 639 2962 643 2963
rect 639 2957 643 2958
rect 695 2962 699 2963
rect 695 2957 699 2958
rect 783 2962 787 2963
rect 783 2957 787 2958
rect 823 2962 827 2963
rect 823 2957 827 2958
rect 919 2962 923 2963
rect 919 2957 923 2958
rect 959 2962 963 2963
rect 959 2957 963 2958
rect 1055 2962 1059 2963
rect 1055 2957 1059 2958
rect 1095 2962 1099 2963
rect 1095 2957 1099 2958
rect 1183 2962 1187 2963
rect 1183 2957 1187 2958
rect 1231 2962 1235 2963
rect 1231 2957 1235 2958
rect 1303 2962 1307 2963
rect 1303 2957 1307 2958
rect 1359 2962 1363 2963
rect 1359 2957 1363 2958
rect 1415 2962 1419 2963
rect 1415 2957 1419 2958
rect 1487 2962 1491 2963
rect 1487 2957 1491 2958
rect 1527 2962 1531 2963
rect 1527 2957 1531 2958
rect 1615 2962 1619 2963
rect 1615 2957 1619 2958
rect 1639 2962 1643 2963
rect 1639 2957 1643 2958
rect 1727 2962 1731 2963
rect 1727 2957 1731 2958
rect 1823 2962 1827 2963
rect 1823 2957 1827 2958
rect 112 2942 114 2957
rect 496 2952 498 2957
rect 640 2952 642 2957
rect 784 2952 786 2957
rect 920 2952 922 2957
rect 1056 2952 1058 2957
rect 1184 2952 1186 2957
rect 1304 2952 1306 2957
rect 1416 2952 1418 2957
rect 1528 2952 1530 2957
rect 1640 2952 1642 2957
rect 1728 2952 1730 2957
rect 494 2951 500 2952
rect 494 2947 495 2951
rect 499 2947 500 2951
rect 494 2946 500 2947
rect 638 2951 644 2952
rect 638 2947 639 2951
rect 643 2947 644 2951
rect 638 2946 644 2947
rect 782 2951 788 2952
rect 782 2947 783 2951
rect 787 2947 788 2951
rect 782 2946 788 2947
rect 918 2951 924 2952
rect 918 2947 919 2951
rect 923 2947 924 2951
rect 918 2946 924 2947
rect 1054 2951 1060 2952
rect 1054 2947 1055 2951
rect 1059 2947 1060 2951
rect 1054 2946 1060 2947
rect 1182 2951 1188 2952
rect 1182 2947 1183 2951
rect 1187 2947 1188 2951
rect 1182 2946 1188 2947
rect 1302 2951 1308 2952
rect 1302 2947 1303 2951
rect 1307 2947 1308 2951
rect 1302 2946 1308 2947
rect 1414 2951 1420 2952
rect 1414 2947 1415 2951
rect 1419 2947 1420 2951
rect 1414 2946 1420 2947
rect 1526 2951 1532 2952
rect 1526 2947 1527 2951
rect 1531 2947 1532 2951
rect 1526 2946 1532 2947
rect 1638 2951 1644 2952
rect 1638 2947 1639 2951
rect 1643 2947 1644 2951
rect 1638 2946 1644 2947
rect 1726 2951 1732 2952
rect 1726 2947 1727 2951
rect 1731 2947 1732 2951
rect 1726 2946 1732 2947
rect 1824 2942 1826 2957
rect 110 2941 116 2942
rect 110 2937 111 2941
rect 115 2937 116 2941
rect 110 2936 116 2937
rect 1822 2941 1828 2942
rect 1822 2937 1823 2941
rect 1827 2937 1828 2941
rect 1822 2936 1828 2937
rect 1864 2935 1866 2967
rect 2030 2959 2036 2960
rect 2030 2955 2031 2959
rect 2035 2955 2036 2959
rect 2030 2954 2036 2955
rect 2166 2959 2172 2960
rect 2166 2955 2167 2959
rect 2171 2955 2172 2959
rect 2166 2954 2172 2955
rect 2294 2959 2300 2960
rect 2294 2955 2295 2959
rect 2299 2955 2300 2959
rect 2294 2954 2300 2955
rect 2422 2959 2428 2960
rect 2422 2955 2423 2959
rect 2427 2955 2428 2959
rect 2422 2954 2428 2955
rect 2542 2959 2548 2960
rect 2542 2955 2543 2959
rect 2547 2955 2548 2959
rect 2542 2954 2548 2955
rect 2670 2959 2676 2960
rect 2670 2955 2671 2959
rect 2675 2955 2676 2959
rect 2670 2954 2676 2955
rect 2814 2959 2820 2960
rect 2814 2955 2815 2959
rect 2819 2955 2820 2959
rect 2814 2954 2820 2955
rect 2974 2959 2980 2960
rect 2974 2955 2975 2959
rect 2979 2955 2980 2959
rect 2974 2954 2980 2955
rect 3150 2959 3156 2960
rect 3150 2955 3151 2959
rect 3155 2955 3156 2959
rect 3150 2954 3156 2955
rect 3326 2959 3332 2960
rect 3326 2955 3327 2959
rect 3331 2955 3332 2959
rect 3326 2954 3332 2955
rect 3486 2959 3492 2960
rect 3486 2955 3487 2959
rect 3491 2955 3492 2959
rect 3486 2954 3492 2955
rect 2032 2935 2034 2954
rect 2168 2935 2170 2954
rect 2296 2935 2298 2954
rect 2424 2935 2426 2954
rect 2544 2935 2546 2954
rect 2672 2935 2674 2954
rect 2816 2935 2818 2954
rect 2976 2935 2978 2954
rect 3152 2935 3154 2954
rect 3328 2935 3330 2954
rect 3488 2935 3490 2954
rect 3576 2935 3578 2967
rect 1863 2934 1867 2935
rect 1863 2929 1867 2930
rect 1895 2934 1899 2935
rect 1895 2929 1899 2930
rect 2031 2934 2035 2935
rect 2031 2929 2035 2930
rect 2167 2934 2171 2935
rect 2167 2929 2171 2930
rect 2175 2934 2179 2935
rect 2175 2929 2179 2930
rect 2295 2934 2299 2935
rect 2295 2929 2299 2930
rect 2423 2934 2427 2935
rect 2423 2929 2427 2930
rect 2495 2934 2499 2935
rect 2495 2929 2499 2930
rect 2543 2934 2547 2935
rect 2543 2929 2547 2930
rect 2671 2934 2675 2935
rect 2671 2929 2675 2930
rect 2815 2934 2819 2935
rect 2815 2929 2819 2930
rect 2823 2934 2827 2935
rect 2823 2929 2827 2930
rect 2975 2934 2979 2935
rect 2975 2929 2979 2930
rect 3151 2934 3155 2935
rect 3151 2929 3155 2930
rect 3167 2934 3171 2935
rect 3167 2929 3171 2930
rect 3327 2934 3331 2935
rect 3327 2929 3331 2930
rect 3487 2934 3491 2935
rect 3487 2929 3491 2930
rect 3575 2934 3579 2935
rect 3575 2929 3579 2930
rect 110 2924 116 2925
rect 110 2920 111 2924
rect 115 2920 116 2924
rect 110 2919 116 2920
rect 1822 2924 1828 2925
rect 1822 2920 1823 2924
rect 1827 2920 1828 2924
rect 1822 2919 1828 2920
rect 112 2891 114 2919
rect 502 2911 508 2912
rect 502 2907 503 2911
rect 507 2907 508 2911
rect 502 2906 508 2907
rect 646 2911 652 2912
rect 646 2907 647 2911
rect 651 2907 652 2911
rect 646 2906 652 2907
rect 790 2911 796 2912
rect 790 2907 791 2911
rect 795 2907 796 2911
rect 790 2906 796 2907
rect 926 2911 932 2912
rect 926 2907 927 2911
rect 931 2907 932 2911
rect 926 2906 932 2907
rect 1062 2911 1068 2912
rect 1062 2907 1063 2911
rect 1067 2907 1068 2911
rect 1062 2906 1068 2907
rect 1190 2911 1196 2912
rect 1190 2907 1191 2911
rect 1195 2907 1196 2911
rect 1190 2906 1196 2907
rect 1310 2911 1316 2912
rect 1310 2907 1311 2911
rect 1315 2907 1316 2911
rect 1310 2906 1316 2907
rect 1422 2911 1428 2912
rect 1422 2907 1423 2911
rect 1427 2907 1428 2911
rect 1422 2906 1428 2907
rect 1534 2911 1540 2912
rect 1534 2907 1535 2911
rect 1539 2907 1540 2911
rect 1534 2906 1540 2907
rect 1646 2911 1652 2912
rect 1646 2907 1647 2911
rect 1651 2907 1652 2911
rect 1646 2906 1652 2907
rect 1734 2911 1740 2912
rect 1734 2907 1735 2911
rect 1739 2907 1740 2911
rect 1734 2906 1740 2907
rect 504 2891 506 2906
rect 648 2891 650 2906
rect 792 2891 794 2906
rect 928 2891 930 2906
rect 1064 2891 1066 2906
rect 1192 2891 1194 2906
rect 1312 2891 1314 2906
rect 1424 2891 1426 2906
rect 1536 2891 1538 2906
rect 1648 2891 1650 2906
rect 1736 2891 1738 2906
rect 1824 2891 1826 2919
rect 1864 2905 1866 2929
rect 1896 2918 1898 2929
rect 2176 2918 2178 2929
rect 2496 2918 2498 2929
rect 2824 2918 2826 2929
rect 3168 2918 3170 2929
rect 3488 2918 3490 2929
rect 1894 2917 1900 2918
rect 1894 2913 1895 2917
rect 1899 2913 1900 2917
rect 1894 2912 1900 2913
rect 2174 2917 2180 2918
rect 2174 2913 2175 2917
rect 2179 2913 2180 2917
rect 2174 2912 2180 2913
rect 2494 2917 2500 2918
rect 2494 2913 2495 2917
rect 2499 2913 2500 2917
rect 2494 2912 2500 2913
rect 2822 2917 2828 2918
rect 2822 2913 2823 2917
rect 2827 2913 2828 2917
rect 2822 2912 2828 2913
rect 3166 2917 3172 2918
rect 3166 2913 3167 2917
rect 3171 2913 3172 2917
rect 3166 2912 3172 2913
rect 3486 2917 3492 2918
rect 3486 2913 3487 2917
rect 3491 2913 3492 2917
rect 3486 2912 3492 2913
rect 3576 2905 3578 2929
rect 1862 2904 1868 2905
rect 1862 2900 1863 2904
rect 1867 2900 1868 2904
rect 1862 2899 1868 2900
rect 3574 2904 3580 2905
rect 3574 2900 3575 2904
rect 3579 2900 3580 2904
rect 3574 2899 3580 2900
rect 111 2890 115 2891
rect 111 2885 115 2886
rect 327 2890 331 2891
rect 327 2885 331 2886
rect 455 2890 459 2891
rect 455 2885 459 2886
rect 503 2890 507 2891
rect 503 2885 507 2886
rect 591 2890 595 2891
rect 591 2885 595 2886
rect 647 2890 651 2891
rect 647 2885 651 2886
rect 727 2890 731 2891
rect 727 2885 731 2886
rect 791 2890 795 2891
rect 791 2885 795 2886
rect 871 2890 875 2891
rect 871 2885 875 2886
rect 927 2890 931 2891
rect 927 2885 931 2886
rect 1007 2890 1011 2891
rect 1007 2885 1011 2886
rect 1063 2890 1067 2891
rect 1063 2885 1067 2886
rect 1143 2890 1147 2891
rect 1143 2885 1147 2886
rect 1191 2890 1195 2891
rect 1191 2885 1195 2886
rect 1279 2890 1283 2891
rect 1279 2885 1283 2886
rect 1311 2890 1315 2891
rect 1311 2885 1315 2886
rect 1415 2890 1419 2891
rect 1415 2885 1419 2886
rect 1423 2890 1427 2891
rect 1423 2885 1427 2886
rect 1535 2890 1539 2891
rect 1535 2885 1539 2886
rect 1551 2890 1555 2891
rect 1551 2885 1555 2886
rect 1647 2890 1651 2891
rect 1647 2885 1651 2886
rect 1735 2890 1739 2891
rect 1735 2885 1739 2886
rect 1823 2890 1827 2891
rect 1823 2885 1827 2886
rect 1862 2887 1868 2888
rect 112 2861 114 2885
rect 328 2874 330 2885
rect 456 2874 458 2885
rect 592 2874 594 2885
rect 728 2874 730 2885
rect 872 2874 874 2885
rect 1008 2874 1010 2885
rect 1144 2874 1146 2885
rect 1280 2874 1282 2885
rect 1416 2874 1418 2885
rect 1552 2874 1554 2885
rect 326 2873 332 2874
rect 326 2869 327 2873
rect 331 2869 332 2873
rect 326 2868 332 2869
rect 454 2873 460 2874
rect 454 2869 455 2873
rect 459 2869 460 2873
rect 454 2868 460 2869
rect 590 2873 596 2874
rect 590 2869 591 2873
rect 595 2869 596 2873
rect 590 2868 596 2869
rect 726 2873 732 2874
rect 726 2869 727 2873
rect 731 2869 732 2873
rect 726 2868 732 2869
rect 870 2873 876 2874
rect 870 2869 871 2873
rect 875 2869 876 2873
rect 870 2868 876 2869
rect 1006 2873 1012 2874
rect 1006 2869 1007 2873
rect 1011 2869 1012 2873
rect 1006 2868 1012 2869
rect 1142 2873 1148 2874
rect 1142 2869 1143 2873
rect 1147 2869 1148 2873
rect 1142 2868 1148 2869
rect 1278 2873 1284 2874
rect 1278 2869 1279 2873
rect 1283 2869 1284 2873
rect 1278 2868 1284 2869
rect 1414 2873 1420 2874
rect 1414 2869 1415 2873
rect 1419 2869 1420 2873
rect 1414 2868 1420 2869
rect 1550 2873 1556 2874
rect 1550 2869 1551 2873
rect 1555 2869 1556 2873
rect 1550 2868 1556 2869
rect 1824 2861 1826 2885
rect 1862 2883 1863 2887
rect 1867 2883 1868 2887
rect 1862 2882 1868 2883
rect 3574 2887 3580 2888
rect 3574 2883 3575 2887
rect 3579 2883 3580 2887
rect 3574 2882 3580 2883
rect 1864 2867 1866 2882
rect 1886 2877 1892 2878
rect 1886 2873 1887 2877
rect 1891 2873 1892 2877
rect 1886 2872 1892 2873
rect 2166 2877 2172 2878
rect 2166 2873 2167 2877
rect 2171 2873 2172 2877
rect 2166 2872 2172 2873
rect 2486 2877 2492 2878
rect 2486 2873 2487 2877
rect 2491 2873 2492 2877
rect 2486 2872 2492 2873
rect 2814 2877 2820 2878
rect 2814 2873 2815 2877
rect 2819 2873 2820 2877
rect 2814 2872 2820 2873
rect 3158 2877 3164 2878
rect 3158 2873 3159 2877
rect 3163 2873 3164 2877
rect 3158 2872 3164 2873
rect 3478 2877 3484 2878
rect 3478 2873 3479 2877
rect 3483 2873 3484 2877
rect 3478 2872 3484 2873
rect 1888 2867 1890 2872
rect 2168 2867 2170 2872
rect 2488 2867 2490 2872
rect 2816 2867 2818 2872
rect 3160 2867 3162 2872
rect 3480 2867 3482 2872
rect 3576 2867 3578 2882
rect 1863 2866 1867 2867
rect 1863 2861 1867 2862
rect 1887 2866 1891 2867
rect 1887 2861 1891 2862
rect 2023 2866 2027 2867
rect 2023 2861 2027 2862
rect 2167 2866 2171 2867
rect 2167 2861 2171 2862
rect 2191 2866 2195 2867
rect 2191 2861 2195 2862
rect 2359 2866 2363 2867
rect 2359 2861 2363 2862
rect 2487 2866 2491 2867
rect 2487 2861 2491 2862
rect 2519 2866 2523 2867
rect 2519 2861 2523 2862
rect 2671 2866 2675 2867
rect 2671 2861 2675 2862
rect 2807 2866 2811 2867
rect 2807 2861 2811 2862
rect 2815 2866 2819 2867
rect 2815 2861 2819 2862
rect 2935 2866 2939 2867
rect 2935 2861 2939 2862
rect 3055 2866 3059 2867
rect 3055 2861 3059 2862
rect 3159 2866 3163 2867
rect 3159 2861 3163 2862
rect 3167 2866 3171 2867
rect 3167 2861 3171 2862
rect 3279 2866 3283 2867
rect 3279 2861 3283 2862
rect 3391 2866 3395 2867
rect 3391 2861 3395 2862
rect 3479 2866 3483 2867
rect 3479 2861 3483 2862
rect 3575 2866 3579 2867
rect 3575 2861 3579 2862
rect 110 2860 116 2861
rect 110 2856 111 2860
rect 115 2856 116 2860
rect 110 2855 116 2856
rect 1822 2860 1828 2861
rect 1822 2856 1823 2860
rect 1827 2856 1828 2860
rect 1822 2855 1828 2856
rect 1864 2846 1866 2861
rect 1888 2856 1890 2861
rect 2024 2856 2026 2861
rect 2192 2856 2194 2861
rect 2360 2856 2362 2861
rect 2520 2856 2522 2861
rect 2672 2856 2674 2861
rect 2808 2856 2810 2861
rect 2936 2856 2938 2861
rect 3056 2856 3058 2861
rect 3168 2856 3170 2861
rect 3280 2856 3282 2861
rect 3392 2856 3394 2861
rect 3480 2856 3482 2861
rect 1886 2855 1892 2856
rect 1886 2851 1887 2855
rect 1891 2851 1892 2855
rect 1886 2850 1892 2851
rect 2022 2855 2028 2856
rect 2022 2851 2023 2855
rect 2027 2851 2028 2855
rect 2022 2850 2028 2851
rect 2190 2855 2196 2856
rect 2190 2851 2191 2855
rect 2195 2851 2196 2855
rect 2190 2850 2196 2851
rect 2358 2855 2364 2856
rect 2358 2851 2359 2855
rect 2363 2851 2364 2855
rect 2358 2850 2364 2851
rect 2518 2855 2524 2856
rect 2518 2851 2519 2855
rect 2523 2851 2524 2855
rect 2518 2850 2524 2851
rect 2670 2855 2676 2856
rect 2670 2851 2671 2855
rect 2675 2851 2676 2855
rect 2670 2850 2676 2851
rect 2806 2855 2812 2856
rect 2806 2851 2807 2855
rect 2811 2851 2812 2855
rect 2806 2850 2812 2851
rect 2934 2855 2940 2856
rect 2934 2851 2935 2855
rect 2939 2851 2940 2855
rect 2934 2850 2940 2851
rect 3054 2855 3060 2856
rect 3054 2851 3055 2855
rect 3059 2851 3060 2855
rect 3054 2850 3060 2851
rect 3166 2855 3172 2856
rect 3166 2851 3167 2855
rect 3171 2851 3172 2855
rect 3166 2850 3172 2851
rect 3278 2855 3284 2856
rect 3278 2851 3279 2855
rect 3283 2851 3284 2855
rect 3278 2850 3284 2851
rect 3390 2855 3396 2856
rect 3390 2851 3391 2855
rect 3395 2851 3396 2855
rect 3390 2850 3396 2851
rect 3478 2855 3484 2856
rect 3478 2851 3479 2855
rect 3483 2851 3484 2855
rect 3478 2850 3484 2851
rect 3576 2846 3578 2861
rect 1862 2845 1868 2846
rect 110 2843 116 2844
rect 110 2839 111 2843
rect 115 2839 116 2843
rect 110 2838 116 2839
rect 1822 2843 1828 2844
rect 1822 2839 1823 2843
rect 1827 2839 1828 2843
rect 1862 2841 1863 2845
rect 1867 2841 1868 2845
rect 1862 2840 1868 2841
rect 3574 2845 3580 2846
rect 3574 2841 3575 2845
rect 3579 2841 3580 2845
rect 3574 2840 3580 2841
rect 1822 2838 1828 2839
rect 112 2815 114 2838
rect 318 2833 324 2834
rect 318 2829 319 2833
rect 323 2829 324 2833
rect 318 2828 324 2829
rect 446 2833 452 2834
rect 446 2829 447 2833
rect 451 2829 452 2833
rect 446 2828 452 2829
rect 582 2833 588 2834
rect 582 2829 583 2833
rect 587 2829 588 2833
rect 582 2828 588 2829
rect 718 2833 724 2834
rect 718 2829 719 2833
rect 723 2829 724 2833
rect 718 2828 724 2829
rect 862 2833 868 2834
rect 862 2829 863 2833
rect 867 2829 868 2833
rect 862 2828 868 2829
rect 998 2833 1004 2834
rect 998 2829 999 2833
rect 1003 2829 1004 2833
rect 998 2828 1004 2829
rect 1134 2833 1140 2834
rect 1134 2829 1135 2833
rect 1139 2829 1140 2833
rect 1134 2828 1140 2829
rect 1270 2833 1276 2834
rect 1270 2829 1271 2833
rect 1275 2829 1276 2833
rect 1270 2828 1276 2829
rect 1406 2833 1412 2834
rect 1406 2829 1407 2833
rect 1411 2829 1412 2833
rect 1406 2828 1412 2829
rect 1542 2833 1548 2834
rect 1542 2829 1543 2833
rect 1547 2829 1548 2833
rect 1542 2828 1548 2829
rect 320 2815 322 2828
rect 448 2815 450 2828
rect 584 2815 586 2828
rect 720 2815 722 2828
rect 864 2815 866 2828
rect 1000 2815 1002 2828
rect 1136 2815 1138 2828
rect 1272 2815 1274 2828
rect 1408 2815 1410 2828
rect 1544 2815 1546 2828
rect 1824 2815 1826 2838
rect 1862 2828 1868 2829
rect 1862 2824 1863 2828
rect 1867 2824 1868 2828
rect 1862 2823 1868 2824
rect 3574 2828 3580 2829
rect 3574 2824 3575 2828
rect 3579 2824 3580 2828
rect 3574 2823 3580 2824
rect 111 2814 115 2815
rect 111 2809 115 2810
rect 167 2814 171 2815
rect 167 2809 171 2810
rect 295 2814 299 2815
rect 295 2809 299 2810
rect 319 2814 323 2815
rect 319 2809 323 2810
rect 423 2814 427 2815
rect 423 2809 427 2810
rect 447 2814 451 2815
rect 447 2809 451 2810
rect 559 2814 563 2815
rect 559 2809 563 2810
rect 583 2814 587 2815
rect 583 2809 587 2810
rect 695 2814 699 2815
rect 695 2809 699 2810
rect 719 2814 723 2815
rect 719 2809 723 2810
rect 823 2814 827 2815
rect 823 2809 827 2810
rect 863 2814 867 2815
rect 863 2809 867 2810
rect 951 2814 955 2815
rect 951 2809 955 2810
rect 999 2814 1003 2815
rect 999 2809 1003 2810
rect 1079 2814 1083 2815
rect 1079 2809 1083 2810
rect 1135 2814 1139 2815
rect 1135 2809 1139 2810
rect 1207 2814 1211 2815
rect 1207 2809 1211 2810
rect 1271 2814 1275 2815
rect 1271 2809 1275 2810
rect 1343 2814 1347 2815
rect 1343 2809 1347 2810
rect 1407 2814 1411 2815
rect 1407 2809 1411 2810
rect 1543 2814 1547 2815
rect 1543 2809 1547 2810
rect 1823 2814 1827 2815
rect 1823 2809 1827 2810
rect 112 2794 114 2809
rect 168 2804 170 2809
rect 296 2804 298 2809
rect 424 2804 426 2809
rect 560 2804 562 2809
rect 696 2804 698 2809
rect 824 2804 826 2809
rect 952 2804 954 2809
rect 1080 2804 1082 2809
rect 1208 2804 1210 2809
rect 1344 2804 1346 2809
rect 166 2803 172 2804
rect 166 2799 167 2803
rect 171 2799 172 2803
rect 166 2798 172 2799
rect 294 2803 300 2804
rect 294 2799 295 2803
rect 299 2799 300 2803
rect 294 2798 300 2799
rect 422 2803 428 2804
rect 422 2799 423 2803
rect 427 2799 428 2803
rect 422 2798 428 2799
rect 558 2803 564 2804
rect 558 2799 559 2803
rect 563 2799 564 2803
rect 558 2798 564 2799
rect 694 2803 700 2804
rect 694 2799 695 2803
rect 699 2799 700 2803
rect 694 2798 700 2799
rect 822 2803 828 2804
rect 822 2799 823 2803
rect 827 2799 828 2803
rect 822 2798 828 2799
rect 950 2803 956 2804
rect 950 2799 951 2803
rect 955 2799 956 2803
rect 950 2798 956 2799
rect 1078 2803 1084 2804
rect 1078 2799 1079 2803
rect 1083 2799 1084 2803
rect 1078 2798 1084 2799
rect 1206 2803 1212 2804
rect 1206 2799 1207 2803
rect 1211 2799 1212 2803
rect 1206 2798 1212 2799
rect 1342 2803 1348 2804
rect 1342 2799 1343 2803
rect 1347 2799 1348 2803
rect 1342 2798 1348 2799
rect 1824 2794 1826 2809
rect 1864 2799 1866 2823
rect 1894 2815 1900 2816
rect 1894 2811 1895 2815
rect 1899 2811 1900 2815
rect 1894 2810 1900 2811
rect 2030 2815 2036 2816
rect 2030 2811 2031 2815
rect 2035 2811 2036 2815
rect 2030 2810 2036 2811
rect 2198 2815 2204 2816
rect 2198 2811 2199 2815
rect 2203 2811 2204 2815
rect 2198 2810 2204 2811
rect 2366 2815 2372 2816
rect 2366 2811 2367 2815
rect 2371 2811 2372 2815
rect 2366 2810 2372 2811
rect 2526 2815 2532 2816
rect 2526 2811 2527 2815
rect 2531 2811 2532 2815
rect 2526 2810 2532 2811
rect 2678 2815 2684 2816
rect 2678 2811 2679 2815
rect 2683 2811 2684 2815
rect 2678 2810 2684 2811
rect 2814 2815 2820 2816
rect 2814 2811 2815 2815
rect 2819 2811 2820 2815
rect 2814 2810 2820 2811
rect 2942 2815 2948 2816
rect 2942 2811 2943 2815
rect 2947 2811 2948 2815
rect 2942 2810 2948 2811
rect 3062 2815 3068 2816
rect 3062 2811 3063 2815
rect 3067 2811 3068 2815
rect 3062 2810 3068 2811
rect 3174 2815 3180 2816
rect 3174 2811 3175 2815
rect 3179 2811 3180 2815
rect 3174 2810 3180 2811
rect 3286 2815 3292 2816
rect 3286 2811 3287 2815
rect 3291 2811 3292 2815
rect 3286 2810 3292 2811
rect 3398 2815 3404 2816
rect 3398 2811 3399 2815
rect 3403 2811 3404 2815
rect 3398 2810 3404 2811
rect 3486 2815 3492 2816
rect 3486 2811 3487 2815
rect 3491 2811 3492 2815
rect 3486 2810 3492 2811
rect 1896 2799 1898 2810
rect 2032 2799 2034 2810
rect 2200 2799 2202 2810
rect 2368 2799 2370 2810
rect 2528 2799 2530 2810
rect 2680 2799 2682 2810
rect 2816 2799 2818 2810
rect 2944 2799 2946 2810
rect 3064 2799 3066 2810
rect 3176 2799 3178 2810
rect 3288 2799 3290 2810
rect 3400 2799 3402 2810
rect 3488 2799 3490 2810
rect 3576 2799 3578 2823
rect 1863 2798 1867 2799
rect 110 2793 116 2794
rect 110 2789 111 2793
rect 115 2789 116 2793
rect 110 2788 116 2789
rect 1822 2793 1828 2794
rect 1863 2793 1867 2794
rect 1895 2798 1899 2799
rect 1895 2793 1899 2794
rect 2031 2798 2035 2799
rect 2031 2793 2035 2794
rect 2063 2798 2067 2799
rect 2063 2793 2067 2794
rect 2199 2798 2203 2799
rect 2199 2793 2203 2794
rect 2255 2798 2259 2799
rect 2255 2793 2259 2794
rect 2367 2798 2371 2799
rect 2367 2793 2371 2794
rect 2439 2798 2443 2799
rect 2439 2793 2443 2794
rect 2527 2798 2531 2799
rect 2527 2793 2531 2794
rect 2615 2798 2619 2799
rect 2615 2793 2619 2794
rect 2679 2798 2683 2799
rect 2679 2793 2683 2794
rect 2783 2798 2787 2799
rect 2783 2793 2787 2794
rect 2815 2798 2819 2799
rect 2815 2793 2819 2794
rect 2935 2798 2939 2799
rect 2935 2793 2939 2794
rect 2943 2798 2947 2799
rect 2943 2793 2947 2794
rect 3063 2798 3067 2799
rect 3063 2793 3067 2794
rect 3079 2798 3083 2799
rect 3079 2793 3083 2794
rect 3175 2798 3179 2799
rect 3175 2793 3179 2794
rect 3223 2798 3227 2799
rect 3223 2793 3227 2794
rect 3287 2798 3291 2799
rect 3287 2793 3291 2794
rect 3367 2798 3371 2799
rect 3367 2793 3371 2794
rect 3399 2798 3403 2799
rect 3399 2793 3403 2794
rect 3487 2798 3491 2799
rect 3487 2793 3491 2794
rect 3575 2798 3579 2799
rect 3575 2793 3579 2794
rect 1822 2789 1823 2793
rect 1827 2789 1828 2793
rect 1822 2788 1828 2789
rect 110 2776 116 2777
rect 110 2772 111 2776
rect 115 2772 116 2776
rect 110 2771 116 2772
rect 1822 2776 1828 2777
rect 1822 2772 1823 2776
rect 1827 2772 1828 2776
rect 1822 2771 1828 2772
rect 112 2739 114 2771
rect 174 2763 180 2764
rect 174 2759 175 2763
rect 179 2759 180 2763
rect 174 2758 180 2759
rect 302 2763 308 2764
rect 302 2759 303 2763
rect 307 2759 308 2763
rect 302 2758 308 2759
rect 430 2763 436 2764
rect 430 2759 431 2763
rect 435 2759 436 2763
rect 430 2758 436 2759
rect 566 2763 572 2764
rect 566 2759 567 2763
rect 571 2759 572 2763
rect 566 2758 572 2759
rect 702 2763 708 2764
rect 702 2759 703 2763
rect 707 2759 708 2763
rect 702 2758 708 2759
rect 830 2763 836 2764
rect 830 2759 831 2763
rect 835 2759 836 2763
rect 830 2758 836 2759
rect 958 2763 964 2764
rect 958 2759 959 2763
rect 963 2759 964 2763
rect 958 2758 964 2759
rect 1086 2763 1092 2764
rect 1086 2759 1087 2763
rect 1091 2759 1092 2763
rect 1086 2758 1092 2759
rect 1214 2763 1220 2764
rect 1214 2759 1215 2763
rect 1219 2759 1220 2763
rect 1214 2758 1220 2759
rect 1350 2763 1356 2764
rect 1350 2759 1351 2763
rect 1355 2759 1356 2763
rect 1350 2758 1356 2759
rect 176 2739 178 2758
rect 304 2739 306 2758
rect 432 2739 434 2758
rect 568 2739 570 2758
rect 704 2739 706 2758
rect 832 2739 834 2758
rect 960 2739 962 2758
rect 1088 2739 1090 2758
rect 1216 2739 1218 2758
rect 1352 2739 1354 2758
rect 1824 2739 1826 2771
rect 1864 2769 1866 2793
rect 1896 2782 1898 2793
rect 2064 2782 2066 2793
rect 2256 2782 2258 2793
rect 2440 2782 2442 2793
rect 2616 2782 2618 2793
rect 2784 2782 2786 2793
rect 2936 2782 2938 2793
rect 3080 2782 3082 2793
rect 3224 2782 3226 2793
rect 3368 2782 3370 2793
rect 3488 2782 3490 2793
rect 1894 2781 1900 2782
rect 1894 2777 1895 2781
rect 1899 2777 1900 2781
rect 1894 2776 1900 2777
rect 2062 2781 2068 2782
rect 2062 2777 2063 2781
rect 2067 2777 2068 2781
rect 2062 2776 2068 2777
rect 2254 2781 2260 2782
rect 2254 2777 2255 2781
rect 2259 2777 2260 2781
rect 2254 2776 2260 2777
rect 2438 2781 2444 2782
rect 2438 2777 2439 2781
rect 2443 2777 2444 2781
rect 2438 2776 2444 2777
rect 2614 2781 2620 2782
rect 2614 2777 2615 2781
rect 2619 2777 2620 2781
rect 2614 2776 2620 2777
rect 2782 2781 2788 2782
rect 2782 2777 2783 2781
rect 2787 2777 2788 2781
rect 2782 2776 2788 2777
rect 2934 2781 2940 2782
rect 2934 2777 2935 2781
rect 2939 2777 2940 2781
rect 2934 2776 2940 2777
rect 3078 2781 3084 2782
rect 3078 2777 3079 2781
rect 3083 2777 3084 2781
rect 3078 2776 3084 2777
rect 3222 2781 3228 2782
rect 3222 2777 3223 2781
rect 3227 2777 3228 2781
rect 3222 2776 3228 2777
rect 3366 2781 3372 2782
rect 3366 2777 3367 2781
rect 3371 2777 3372 2781
rect 3366 2776 3372 2777
rect 3486 2781 3492 2782
rect 3486 2777 3487 2781
rect 3491 2777 3492 2781
rect 3486 2776 3492 2777
rect 3576 2769 3578 2793
rect 1862 2768 1868 2769
rect 1862 2764 1863 2768
rect 1867 2764 1868 2768
rect 1862 2763 1868 2764
rect 3574 2768 3580 2769
rect 3574 2764 3575 2768
rect 3579 2764 3580 2768
rect 3574 2763 3580 2764
rect 1862 2751 1868 2752
rect 1862 2747 1863 2751
rect 1867 2747 1868 2751
rect 1862 2746 1868 2747
rect 3574 2751 3580 2752
rect 3574 2747 3575 2751
rect 3579 2747 3580 2751
rect 3574 2746 3580 2747
rect 111 2738 115 2739
rect 111 2733 115 2734
rect 143 2738 147 2739
rect 143 2733 147 2734
rect 175 2738 179 2739
rect 175 2733 179 2734
rect 231 2738 235 2739
rect 231 2733 235 2734
rect 303 2738 307 2739
rect 303 2733 307 2734
rect 351 2738 355 2739
rect 351 2733 355 2734
rect 431 2738 435 2739
rect 431 2733 435 2734
rect 479 2738 483 2739
rect 479 2733 483 2734
rect 567 2738 571 2739
rect 567 2733 571 2734
rect 615 2738 619 2739
rect 615 2733 619 2734
rect 703 2738 707 2739
rect 703 2733 707 2734
rect 759 2738 763 2739
rect 759 2733 763 2734
rect 831 2738 835 2739
rect 831 2733 835 2734
rect 903 2738 907 2739
rect 903 2733 907 2734
rect 959 2738 963 2739
rect 959 2733 963 2734
rect 1047 2738 1051 2739
rect 1047 2733 1051 2734
rect 1087 2738 1091 2739
rect 1087 2733 1091 2734
rect 1215 2738 1219 2739
rect 1215 2733 1219 2734
rect 1351 2738 1355 2739
rect 1351 2733 1355 2734
rect 1823 2738 1827 2739
rect 1823 2733 1827 2734
rect 112 2709 114 2733
rect 144 2722 146 2733
rect 232 2722 234 2733
rect 352 2722 354 2733
rect 480 2722 482 2733
rect 616 2722 618 2733
rect 760 2722 762 2733
rect 904 2722 906 2733
rect 1048 2722 1050 2733
rect 142 2721 148 2722
rect 142 2717 143 2721
rect 147 2717 148 2721
rect 142 2716 148 2717
rect 230 2721 236 2722
rect 230 2717 231 2721
rect 235 2717 236 2721
rect 230 2716 236 2717
rect 350 2721 356 2722
rect 350 2717 351 2721
rect 355 2717 356 2721
rect 350 2716 356 2717
rect 478 2721 484 2722
rect 478 2717 479 2721
rect 483 2717 484 2721
rect 478 2716 484 2717
rect 614 2721 620 2722
rect 614 2717 615 2721
rect 619 2717 620 2721
rect 614 2716 620 2717
rect 758 2721 764 2722
rect 758 2717 759 2721
rect 763 2717 764 2721
rect 758 2716 764 2717
rect 902 2721 908 2722
rect 902 2717 903 2721
rect 907 2717 908 2721
rect 902 2716 908 2717
rect 1046 2721 1052 2722
rect 1046 2717 1047 2721
rect 1051 2717 1052 2721
rect 1046 2716 1052 2717
rect 1824 2709 1826 2733
rect 1864 2727 1866 2746
rect 1886 2741 1892 2742
rect 1886 2737 1887 2741
rect 1891 2737 1892 2741
rect 1886 2736 1892 2737
rect 2054 2741 2060 2742
rect 2054 2737 2055 2741
rect 2059 2737 2060 2741
rect 2054 2736 2060 2737
rect 2246 2741 2252 2742
rect 2246 2737 2247 2741
rect 2251 2737 2252 2741
rect 2246 2736 2252 2737
rect 2430 2741 2436 2742
rect 2430 2737 2431 2741
rect 2435 2737 2436 2741
rect 2430 2736 2436 2737
rect 2606 2741 2612 2742
rect 2606 2737 2607 2741
rect 2611 2737 2612 2741
rect 2606 2736 2612 2737
rect 2774 2741 2780 2742
rect 2774 2737 2775 2741
rect 2779 2737 2780 2741
rect 2774 2736 2780 2737
rect 2926 2741 2932 2742
rect 2926 2737 2927 2741
rect 2931 2737 2932 2741
rect 2926 2736 2932 2737
rect 3070 2741 3076 2742
rect 3070 2737 3071 2741
rect 3075 2737 3076 2741
rect 3070 2736 3076 2737
rect 3214 2741 3220 2742
rect 3214 2737 3215 2741
rect 3219 2737 3220 2741
rect 3214 2736 3220 2737
rect 3358 2741 3364 2742
rect 3358 2737 3359 2741
rect 3363 2737 3364 2741
rect 3358 2736 3364 2737
rect 3478 2741 3484 2742
rect 3478 2737 3479 2741
rect 3483 2737 3484 2741
rect 3478 2736 3484 2737
rect 1888 2727 1890 2736
rect 2056 2727 2058 2736
rect 2248 2727 2250 2736
rect 2432 2727 2434 2736
rect 2608 2727 2610 2736
rect 2776 2727 2778 2736
rect 2928 2727 2930 2736
rect 3072 2727 3074 2736
rect 3216 2727 3218 2736
rect 3360 2727 3362 2736
rect 3480 2727 3482 2736
rect 3576 2727 3578 2746
rect 1863 2726 1867 2727
rect 1863 2721 1867 2722
rect 1887 2726 1891 2727
rect 1887 2721 1891 2722
rect 2047 2726 2051 2727
rect 2047 2721 2051 2722
rect 2055 2726 2059 2727
rect 2055 2721 2059 2722
rect 2207 2726 2211 2727
rect 2207 2721 2211 2722
rect 2247 2726 2251 2727
rect 2247 2721 2251 2722
rect 2359 2726 2363 2727
rect 2359 2721 2363 2722
rect 2431 2726 2435 2727
rect 2431 2721 2435 2722
rect 2495 2726 2499 2727
rect 2495 2721 2499 2722
rect 2607 2726 2611 2727
rect 2607 2721 2611 2722
rect 2623 2726 2627 2727
rect 2623 2721 2627 2722
rect 2743 2726 2747 2727
rect 2743 2721 2747 2722
rect 2775 2726 2779 2727
rect 2775 2721 2779 2722
rect 2863 2726 2867 2727
rect 2863 2721 2867 2722
rect 2927 2726 2931 2727
rect 2927 2721 2931 2722
rect 2983 2726 2987 2727
rect 2983 2721 2987 2722
rect 3071 2726 3075 2727
rect 3071 2721 3075 2722
rect 3103 2726 3107 2727
rect 3103 2721 3107 2722
rect 3215 2726 3219 2727
rect 3215 2721 3219 2722
rect 3359 2726 3363 2727
rect 3359 2721 3363 2722
rect 3479 2726 3483 2727
rect 3479 2721 3483 2722
rect 3575 2726 3579 2727
rect 3575 2721 3579 2722
rect 110 2708 116 2709
rect 110 2704 111 2708
rect 115 2704 116 2708
rect 110 2703 116 2704
rect 1822 2708 1828 2709
rect 1822 2704 1823 2708
rect 1827 2704 1828 2708
rect 1864 2706 1866 2721
rect 1888 2716 1890 2721
rect 2048 2716 2050 2721
rect 2208 2716 2210 2721
rect 2360 2716 2362 2721
rect 2496 2716 2498 2721
rect 2624 2716 2626 2721
rect 2744 2716 2746 2721
rect 2864 2716 2866 2721
rect 2984 2716 2986 2721
rect 3104 2716 3106 2721
rect 1886 2715 1892 2716
rect 1886 2711 1887 2715
rect 1891 2711 1892 2715
rect 1886 2710 1892 2711
rect 2046 2715 2052 2716
rect 2046 2711 2047 2715
rect 2051 2711 2052 2715
rect 2046 2710 2052 2711
rect 2206 2715 2212 2716
rect 2206 2711 2207 2715
rect 2211 2711 2212 2715
rect 2206 2710 2212 2711
rect 2358 2715 2364 2716
rect 2358 2711 2359 2715
rect 2363 2711 2364 2715
rect 2358 2710 2364 2711
rect 2494 2715 2500 2716
rect 2494 2711 2495 2715
rect 2499 2711 2500 2715
rect 2494 2710 2500 2711
rect 2622 2715 2628 2716
rect 2622 2711 2623 2715
rect 2627 2711 2628 2715
rect 2622 2710 2628 2711
rect 2742 2715 2748 2716
rect 2742 2711 2743 2715
rect 2747 2711 2748 2715
rect 2742 2710 2748 2711
rect 2862 2715 2868 2716
rect 2862 2711 2863 2715
rect 2867 2711 2868 2715
rect 2862 2710 2868 2711
rect 2982 2715 2988 2716
rect 2982 2711 2983 2715
rect 2987 2711 2988 2715
rect 2982 2710 2988 2711
rect 3102 2715 3108 2716
rect 3102 2711 3103 2715
rect 3107 2711 3108 2715
rect 3102 2710 3108 2711
rect 3576 2706 3578 2721
rect 1822 2703 1828 2704
rect 1862 2705 1868 2706
rect 1862 2701 1863 2705
rect 1867 2701 1868 2705
rect 1862 2700 1868 2701
rect 3574 2705 3580 2706
rect 3574 2701 3575 2705
rect 3579 2701 3580 2705
rect 3574 2700 3580 2701
rect 110 2691 116 2692
rect 110 2687 111 2691
rect 115 2687 116 2691
rect 110 2686 116 2687
rect 1822 2691 1828 2692
rect 1822 2687 1823 2691
rect 1827 2687 1828 2691
rect 1822 2686 1828 2687
rect 1862 2688 1868 2689
rect 112 2667 114 2686
rect 134 2681 140 2682
rect 134 2677 135 2681
rect 139 2677 140 2681
rect 134 2676 140 2677
rect 222 2681 228 2682
rect 222 2677 223 2681
rect 227 2677 228 2681
rect 222 2676 228 2677
rect 342 2681 348 2682
rect 342 2677 343 2681
rect 347 2677 348 2681
rect 342 2676 348 2677
rect 470 2681 476 2682
rect 470 2677 471 2681
rect 475 2677 476 2681
rect 470 2676 476 2677
rect 606 2681 612 2682
rect 606 2677 607 2681
rect 611 2677 612 2681
rect 606 2676 612 2677
rect 750 2681 756 2682
rect 750 2677 751 2681
rect 755 2677 756 2681
rect 750 2676 756 2677
rect 894 2681 900 2682
rect 894 2677 895 2681
rect 899 2677 900 2681
rect 894 2676 900 2677
rect 1038 2681 1044 2682
rect 1038 2677 1039 2681
rect 1043 2677 1044 2681
rect 1038 2676 1044 2677
rect 136 2667 138 2676
rect 224 2667 226 2676
rect 344 2667 346 2676
rect 472 2667 474 2676
rect 608 2667 610 2676
rect 752 2667 754 2676
rect 896 2667 898 2676
rect 1040 2667 1042 2676
rect 1824 2667 1826 2686
rect 1862 2684 1863 2688
rect 1867 2684 1868 2688
rect 1862 2683 1868 2684
rect 3574 2688 3580 2689
rect 3574 2684 3575 2688
rect 3579 2684 3580 2688
rect 3574 2683 3580 2684
rect 111 2666 115 2667
rect 111 2661 115 2662
rect 135 2666 139 2667
rect 135 2661 139 2662
rect 223 2666 227 2667
rect 223 2661 227 2662
rect 231 2666 235 2667
rect 231 2661 235 2662
rect 343 2666 347 2667
rect 343 2661 347 2662
rect 351 2666 355 2667
rect 351 2661 355 2662
rect 471 2666 475 2667
rect 471 2661 475 2662
rect 583 2666 587 2667
rect 583 2661 587 2662
rect 607 2666 611 2667
rect 607 2661 611 2662
rect 695 2666 699 2667
rect 695 2661 699 2662
rect 751 2666 755 2667
rect 751 2661 755 2662
rect 799 2666 803 2667
rect 799 2661 803 2662
rect 895 2666 899 2667
rect 895 2661 899 2662
rect 903 2666 907 2667
rect 903 2661 907 2662
rect 999 2666 1003 2667
rect 999 2661 1003 2662
rect 1039 2666 1043 2667
rect 1039 2661 1043 2662
rect 1103 2666 1107 2667
rect 1103 2661 1107 2662
rect 1207 2666 1211 2667
rect 1207 2661 1211 2662
rect 1311 2666 1315 2667
rect 1311 2661 1315 2662
rect 1823 2666 1827 2667
rect 1823 2661 1827 2662
rect 112 2646 114 2661
rect 136 2656 138 2661
rect 232 2656 234 2661
rect 352 2656 354 2661
rect 472 2656 474 2661
rect 584 2656 586 2661
rect 696 2656 698 2661
rect 800 2656 802 2661
rect 904 2656 906 2661
rect 1000 2656 1002 2661
rect 1104 2656 1106 2661
rect 1208 2656 1210 2661
rect 1312 2656 1314 2661
rect 134 2655 140 2656
rect 134 2651 135 2655
rect 139 2651 140 2655
rect 134 2650 140 2651
rect 230 2655 236 2656
rect 230 2651 231 2655
rect 235 2651 236 2655
rect 230 2650 236 2651
rect 350 2655 356 2656
rect 350 2651 351 2655
rect 355 2651 356 2655
rect 350 2650 356 2651
rect 470 2655 476 2656
rect 470 2651 471 2655
rect 475 2651 476 2655
rect 470 2650 476 2651
rect 582 2655 588 2656
rect 582 2651 583 2655
rect 587 2651 588 2655
rect 582 2650 588 2651
rect 694 2655 700 2656
rect 694 2651 695 2655
rect 699 2651 700 2655
rect 694 2650 700 2651
rect 798 2655 804 2656
rect 798 2651 799 2655
rect 803 2651 804 2655
rect 798 2650 804 2651
rect 902 2655 908 2656
rect 902 2651 903 2655
rect 907 2651 908 2655
rect 902 2650 908 2651
rect 998 2655 1004 2656
rect 998 2651 999 2655
rect 1003 2651 1004 2655
rect 998 2650 1004 2651
rect 1102 2655 1108 2656
rect 1102 2651 1103 2655
rect 1107 2651 1108 2655
rect 1102 2650 1108 2651
rect 1206 2655 1212 2656
rect 1206 2651 1207 2655
rect 1211 2651 1212 2655
rect 1206 2650 1212 2651
rect 1310 2655 1316 2656
rect 1310 2651 1311 2655
rect 1315 2651 1316 2655
rect 1310 2650 1316 2651
rect 1824 2646 1826 2661
rect 1864 2651 1866 2683
rect 1894 2675 1900 2676
rect 1894 2671 1895 2675
rect 1899 2671 1900 2675
rect 1894 2670 1900 2671
rect 2054 2675 2060 2676
rect 2054 2671 2055 2675
rect 2059 2671 2060 2675
rect 2054 2670 2060 2671
rect 2214 2675 2220 2676
rect 2214 2671 2215 2675
rect 2219 2671 2220 2675
rect 2214 2670 2220 2671
rect 2366 2675 2372 2676
rect 2366 2671 2367 2675
rect 2371 2671 2372 2675
rect 2366 2670 2372 2671
rect 2502 2675 2508 2676
rect 2502 2671 2503 2675
rect 2507 2671 2508 2675
rect 2502 2670 2508 2671
rect 2630 2675 2636 2676
rect 2630 2671 2631 2675
rect 2635 2671 2636 2675
rect 2630 2670 2636 2671
rect 2750 2675 2756 2676
rect 2750 2671 2751 2675
rect 2755 2671 2756 2675
rect 2750 2670 2756 2671
rect 2870 2675 2876 2676
rect 2870 2671 2871 2675
rect 2875 2671 2876 2675
rect 2870 2670 2876 2671
rect 2990 2675 2996 2676
rect 2990 2671 2991 2675
rect 2995 2671 2996 2675
rect 2990 2670 2996 2671
rect 3110 2675 3116 2676
rect 3110 2671 3111 2675
rect 3115 2671 3116 2675
rect 3110 2670 3116 2671
rect 1896 2651 1898 2670
rect 2056 2651 2058 2670
rect 2216 2651 2218 2670
rect 2368 2651 2370 2670
rect 2504 2651 2506 2670
rect 2632 2651 2634 2670
rect 2752 2651 2754 2670
rect 2872 2651 2874 2670
rect 2992 2651 2994 2670
rect 3112 2651 3114 2670
rect 3576 2651 3578 2683
rect 1863 2650 1867 2651
rect 110 2645 116 2646
rect 110 2641 111 2645
rect 115 2641 116 2645
rect 110 2640 116 2641
rect 1822 2645 1828 2646
rect 1863 2645 1867 2646
rect 1895 2650 1899 2651
rect 1895 2645 1899 2646
rect 1999 2650 2003 2651
rect 1999 2645 2003 2646
rect 2055 2650 2059 2651
rect 2055 2645 2059 2646
rect 2119 2650 2123 2651
rect 2119 2645 2123 2646
rect 2215 2650 2219 2651
rect 2215 2645 2219 2646
rect 2239 2650 2243 2651
rect 2239 2645 2243 2646
rect 2351 2650 2355 2651
rect 2351 2645 2355 2646
rect 2367 2650 2371 2651
rect 2367 2645 2371 2646
rect 2455 2650 2459 2651
rect 2455 2645 2459 2646
rect 2503 2650 2507 2651
rect 2503 2645 2507 2646
rect 2551 2650 2555 2651
rect 2551 2645 2555 2646
rect 2631 2650 2635 2651
rect 2631 2645 2635 2646
rect 2655 2650 2659 2651
rect 2655 2645 2659 2646
rect 2751 2650 2755 2651
rect 2751 2645 2755 2646
rect 2759 2650 2763 2651
rect 2759 2645 2763 2646
rect 2863 2650 2867 2651
rect 2863 2645 2867 2646
rect 2871 2650 2875 2651
rect 2871 2645 2875 2646
rect 2991 2650 2995 2651
rect 2991 2645 2995 2646
rect 3111 2650 3115 2651
rect 3111 2645 3115 2646
rect 3575 2650 3579 2651
rect 3575 2645 3579 2646
rect 1822 2641 1823 2645
rect 1827 2641 1828 2645
rect 1822 2640 1828 2641
rect 110 2628 116 2629
rect 110 2624 111 2628
rect 115 2624 116 2628
rect 110 2623 116 2624
rect 1822 2628 1828 2629
rect 1822 2624 1823 2628
rect 1827 2624 1828 2628
rect 1822 2623 1828 2624
rect 112 2595 114 2623
rect 142 2615 148 2616
rect 142 2611 143 2615
rect 147 2611 148 2615
rect 142 2610 148 2611
rect 238 2615 244 2616
rect 238 2611 239 2615
rect 243 2611 244 2615
rect 238 2610 244 2611
rect 358 2615 364 2616
rect 358 2611 359 2615
rect 363 2611 364 2615
rect 358 2610 364 2611
rect 478 2615 484 2616
rect 478 2611 479 2615
rect 483 2611 484 2615
rect 478 2610 484 2611
rect 590 2615 596 2616
rect 590 2611 591 2615
rect 595 2611 596 2615
rect 590 2610 596 2611
rect 702 2615 708 2616
rect 702 2611 703 2615
rect 707 2611 708 2615
rect 702 2610 708 2611
rect 806 2615 812 2616
rect 806 2611 807 2615
rect 811 2611 812 2615
rect 806 2610 812 2611
rect 910 2615 916 2616
rect 910 2611 911 2615
rect 915 2611 916 2615
rect 910 2610 916 2611
rect 1006 2615 1012 2616
rect 1006 2611 1007 2615
rect 1011 2611 1012 2615
rect 1006 2610 1012 2611
rect 1110 2615 1116 2616
rect 1110 2611 1111 2615
rect 1115 2611 1116 2615
rect 1110 2610 1116 2611
rect 1214 2615 1220 2616
rect 1214 2611 1215 2615
rect 1219 2611 1220 2615
rect 1214 2610 1220 2611
rect 1318 2615 1324 2616
rect 1318 2611 1319 2615
rect 1323 2611 1324 2615
rect 1318 2610 1324 2611
rect 144 2595 146 2610
rect 240 2595 242 2610
rect 360 2595 362 2610
rect 480 2595 482 2610
rect 592 2595 594 2610
rect 704 2595 706 2610
rect 808 2595 810 2610
rect 912 2595 914 2610
rect 1008 2595 1010 2610
rect 1112 2595 1114 2610
rect 1216 2595 1218 2610
rect 1320 2595 1322 2610
rect 1824 2595 1826 2623
rect 1864 2621 1866 2645
rect 1896 2634 1898 2645
rect 2000 2634 2002 2645
rect 2120 2634 2122 2645
rect 2240 2634 2242 2645
rect 2352 2634 2354 2645
rect 2456 2634 2458 2645
rect 2552 2634 2554 2645
rect 2656 2634 2658 2645
rect 2760 2634 2762 2645
rect 2864 2634 2866 2645
rect 1894 2633 1900 2634
rect 1894 2629 1895 2633
rect 1899 2629 1900 2633
rect 1894 2628 1900 2629
rect 1998 2633 2004 2634
rect 1998 2629 1999 2633
rect 2003 2629 2004 2633
rect 1998 2628 2004 2629
rect 2118 2633 2124 2634
rect 2118 2629 2119 2633
rect 2123 2629 2124 2633
rect 2118 2628 2124 2629
rect 2238 2633 2244 2634
rect 2238 2629 2239 2633
rect 2243 2629 2244 2633
rect 2238 2628 2244 2629
rect 2350 2633 2356 2634
rect 2350 2629 2351 2633
rect 2355 2629 2356 2633
rect 2350 2628 2356 2629
rect 2454 2633 2460 2634
rect 2454 2629 2455 2633
rect 2459 2629 2460 2633
rect 2454 2628 2460 2629
rect 2550 2633 2556 2634
rect 2550 2629 2551 2633
rect 2555 2629 2556 2633
rect 2550 2628 2556 2629
rect 2654 2633 2660 2634
rect 2654 2629 2655 2633
rect 2659 2629 2660 2633
rect 2654 2628 2660 2629
rect 2758 2633 2764 2634
rect 2758 2629 2759 2633
rect 2763 2629 2764 2633
rect 2758 2628 2764 2629
rect 2862 2633 2868 2634
rect 2862 2629 2863 2633
rect 2867 2629 2868 2633
rect 2862 2628 2868 2629
rect 3576 2621 3578 2645
rect 1862 2620 1868 2621
rect 1862 2616 1863 2620
rect 1867 2616 1868 2620
rect 1862 2615 1868 2616
rect 3574 2620 3580 2621
rect 3574 2616 3575 2620
rect 3579 2616 3580 2620
rect 3574 2615 3580 2616
rect 1862 2603 1868 2604
rect 1862 2599 1863 2603
rect 1867 2599 1868 2603
rect 1862 2598 1868 2599
rect 3574 2603 3580 2604
rect 3574 2599 3575 2603
rect 3579 2599 3580 2603
rect 3574 2598 3580 2599
rect 111 2594 115 2595
rect 111 2589 115 2590
rect 143 2594 147 2595
rect 143 2589 147 2590
rect 239 2594 243 2595
rect 239 2589 243 2590
rect 271 2594 275 2595
rect 271 2589 275 2590
rect 359 2594 363 2595
rect 359 2589 363 2590
rect 415 2594 419 2595
rect 415 2589 419 2590
rect 479 2594 483 2595
rect 479 2589 483 2590
rect 551 2594 555 2595
rect 551 2589 555 2590
rect 591 2594 595 2595
rect 591 2589 595 2590
rect 679 2594 683 2595
rect 679 2589 683 2590
rect 703 2594 707 2595
rect 703 2589 707 2590
rect 807 2594 811 2595
rect 807 2589 811 2590
rect 911 2594 915 2595
rect 911 2589 915 2590
rect 927 2594 931 2595
rect 927 2589 931 2590
rect 1007 2594 1011 2595
rect 1007 2589 1011 2590
rect 1047 2594 1051 2595
rect 1047 2589 1051 2590
rect 1111 2594 1115 2595
rect 1111 2589 1115 2590
rect 1175 2594 1179 2595
rect 1175 2589 1179 2590
rect 1215 2594 1219 2595
rect 1215 2589 1219 2590
rect 1319 2594 1323 2595
rect 1319 2589 1323 2590
rect 1823 2594 1827 2595
rect 1823 2589 1827 2590
rect 112 2565 114 2589
rect 144 2578 146 2589
rect 272 2578 274 2589
rect 416 2578 418 2589
rect 552 2578 554 2589
rect 680 2578 682 2589
rect 808 2578 810 2589
rect 928 2578 930 2589
rect 1048 2578 1050 2589
rect 1176 2578 1178 2589
rect 142 2577 148 2578
rect 142 2573 143 2577
rect 147 2573 148 2577
rect 142 2572 148 2573
rect 270 2577 276 2578
rect 270 2573 271 2577
rect 275 2573 276 2577
rect 270 2572 276 2573
rect 414 2577 420 2578
rect 414 2573 415 2577
rect 419 2573 420 2577
rect 414 2572 420 2573
rect 550 2577 556 2578
rect 550 2573 551 2577
rect 555 2573 556 2577
rect 550 2572 556 2573
rect 678 2577 684 2578
rect 678 2573 679 2577
rect 683 2573 684 2577
rect 678 2572 684 2573
rect 806 2577 812 2578
rect 806 2573 807 2577
rect 811 2573 812 2577
rect 806 2572 812 2573
rect 926 2577 932 2578
rect 926 2573 927 2577
rect 931 2573 932 2577
rect 926 2572 932 2573
rect 1046 2577 1052 2578
rect 1046 2573 1047 2577
rect 1051 2573 1052 2577
rect 1046 2572 1052 2573
rect 1174 2577 1180 2578
rect 1174 2573 1175 2577
rect 1179 2573 1180 2577
rect 1174 2572 1180 2573
rect 1824 2565 1826 2589
rect 1864 2579 1866 2598
rect 1886 2593 1892 2594
rect 1886 2589 1887 2593
rect 1891 2589 1892 2593
rect 1886 2588 1892 2589
rect 1990 2593 1996 2594
rect 1990 2589 1991 2593
rect 1995 2589 1996 2593
rect 1990 2588 1996 2589
rect 2110 2593 2116 2594
rect 2110 2589 2111 2593
rect 2115 2589 2116 2593
rect 2110 2588 2116 2589
rect 2230 2593 2236 2594
rect 2230 2589 2231 2593
rect 2235 2589 2236 2593
rect 2230 2588 2236 2589
rect 2342 2593 2348 2594
rect 2342 2589 2343 2593
rect 2347 2589 2348 2593
rect 2342 2588 2348 2589
rect 2446 2593 2452 2594
rect 2446 2589 2447 2593
rect 2451 2589 2452 2593
rect 2446 2588 2452 2589
rect 2542 2593 2548 2594
rect 2542 2589 2543 2593
rect 2547 2589 2548 2593
rect 2542 2588 2548 2589
rect 2646 2593 2652 2594
rect 2646 2589 2647 2593
rect 2651 2589 2652 2593
rect 2646 2588 2652 2589
rect 2750 2593 2756 2594
rect 2750 2589 2751 2593
rect 2755 2589 2756 2593
rect 2750 2588 2756 2589
rect 2854 2593 2860 2594
rect 2854 2589 2855 2593
rect 2859 2589 2860 2593
rect 2854 2588 2860 2589
rect 1888 2579 1890 2588
rect 1992 2579 1994 2588
rect 2112 2579 2114 2588
rect 2232 2579 2234 2588
rect 2344 2579 2346 2588
rect 2448 2579 2450 2588
rect 2544 2579 2546 2588
rect 2648 2579 2650 2588
rect 2752 2579 2754 2588
rect 2856 2579 2858 2588
rect 3576 2579 3578 2598
rect 1863 2578 1867 2579
rect 1863 2573 1867 2574
rect 1887 2578 1891 2579
rect 1887 2573 1891 2574
rect 1991 2578 1995 2579
rect 1991 2573 1995 2574
rect 2111 2578 2115 2579
rect 2111 2573 2115 2574
rect 2231 2578 2235 2579
rect 2231 2573 2235 2574
rect 2343 2578 2347 2579
rect 2343 2573 2347 2574
rect 2351 2578 2355 2579
rect 2351 2573 2355 2574
rect 2447 2578 2451 2579
rect 2447 2573 2451 2574
rect 2471 2578 2475 2579
rect 2471 2573 2475 2574
rect 2543 2578 2547 2579
rect 2543 2573 2547 2574
rect 2591 2578 2595 2579
rect 2591 2573 2595 2574
rect 2647 2578 2651 2579
rect 2647 2573 2651 2574
rect 2711 2578 2715 2579
rect 2711 2573 2715 2574
rect 2751 2578 2755 2579
rect 2751 2573 2755 2574
rect 2831 2578 2835 2579
rect 2831 2573 2835 2574
rect 2855 2578 2859 2579
rect 2855 2573 2859 2574
rect 3575 2578 3579 2579
rect 3575 2573 3579 2574
rect 110 2564 116 2565
rect 110 2560 111 2564
rect 115 2560 116 2564
rect 110 2559 116 2560
rect 1822 2564 1828 2565
rect 1822 2560 1823 2564
rect 1827 2560 1828 2564
rect 1822 2559 1828 2560
rect 1864 2558 1866 2573
rect 1888 2568 1890 2573
rect 1992 2568 1994 2573
rect 2112 2568 2114 2573
rect 2232 2568 2234 2573
rect 2352 2568 2354 2573
rect 2472 2568 2474 2573
rect 2592 2568 2594 2573
rect 2712 2568 2714 2573
rect 2832 2568 2834 2573
rect 1886 2567 1892 2568
rect 1886 2563 1887 2567
rect 1891 2563 1892 2567
rect 1886 2562 1892 2563
rect 1990 2567 1996 2568
rect 1990 2563 1991 2567
rect 1995 2563 1996 2567
rect 1990 2562 1996 2563
rect 2110 2567 2116 2568
rect 2110 2563 2111 2567
rect 2115 2563 2116 2567
rect 2110 2562 2116 2563
rect 2230 2567 2236 2568
rect 2230 2563 2231 2567
rect 2235 2563 2236 2567
rect 2230 2562 2236 2563
rect 2350 2567 2356 2568
rect 2350 2563 2351 2567
rect 2355 2563 2356 2567
rect 2350 2562 2356 2563
rect 2470 2567 2476 2568
rect 2470 2563 2471 2567
rect 2475 2563 2476 2567
rect 2470 2562 2476 2563
rect 2590 2567 2596 2568
rect 2590 2563 2591 2567
rect 2595 2563 2596 2567
rect 2590 2562 2596 2563
rect 2710 2567 2716 2568
rect 2710 2563 2711 2567
rect 2715 2563 2716 2567
rect 2710 2562 2716 2563
rect 2830 2567 2836 2568
rect 2830 2563 2831 2567
rect 2835 2563 2836 2567
rect 2830 2562 2836 2563
rect 3576 2558 3578 2573
rect 1862 2557 1868 2558
rect 1862 2553 1863 2557
rect 1867 2553 1868 2557
rect 1862 2552 1868 2553
rect 3574 2557 3580 2558
rect 3574 2553 3575 2557
rect 3579 2553 3580 2557
rect 3574 2552 3580 2553
rect 110 2547 116 2548
rect 110 2543 111 2547
rect 115 2543 116 2547
rect 110 2542 116 2543
rect 1822 2547 1828 2548
rect 1822 2543 1823 2547
rect 1827 2543 1828 2547
rect 1822 2542 1828 2543
rect 112 2527 114 2542
rect 134 2537 140 2538
rect 134 2533 135 2537
rect 139 2533 140 2537
rect 134 2532 140 2533
rect 262 2537 268 2538
rect 262 2533 263 2537
rect 267 2533 268 2537
rect 262 2532 268 2533
rect 406 2537 412 2538
rect 406 2533 407 2537
rect 411 2533 412 2537
rect 406 2532 412 2533
rect 542 2537 548 2538
rect 542 2533 543 2537
rect 547 2533 548 2537
rect 542 2532 548 2533
rect 670 2537 676 2538
rect 670 2533 671 2537
rect 675 2533 676 2537
rect 670 2532 676 2533
rect 798 2537 804 2538
rect 798 2533 799 2537
rect 803 2533 804 2537
rect 798 2532 804 2533
rect 918 2537 924 2538
rect 918 2533 919 2537
rect 923 2533 924 2537
rect 918 2532 924 2533
rect 1038 2537 1044 2538
rect 1038 2533 1039 2537
rect 1043 2533 1044 2537
rect 1038 2532 1044 2533
rect 1166 2537 1172 2538
rect 1166 2533 1167 2537
rect 1171 2533 1172 2537
rect 1166 2532 1172 2533
rect 136 2527 138 2532
rect 264 2527 266 2532
rect 408 2527 410 2532
rect 544 2527 546 2532
rect 672 2527 674 2532
rect 800 2527 802 2532
rect 920 2527 922 2532
rect 1040 2527 1042 2532
rect 1168 2527 1170 2532
rect 1824 2527 1826 2542
rect 1862 2540 1868 2541
rect 1862 2536 1863 2540
rect 1867 2536 1868 2540
rect 1862 2535 1868 2536
rect 3574 2540 3580 2541
rect 3574 2536 3575 2540
rect 3579 2536 3580 2540
rect 3574 2535 3580 2536
rect 111 2526 115 2527
rect 111 2521 115 2522
rect 135 2526 139 2527
rect 135 2521 139 2522
rect 263 2526 267 2527
rect 263 2521 267 2522
rect 279 2526 283 2527
rect 279 2521 283 2522
rect 407 2526 411 2527
rect 407 2521 411 2522
rect 439 2526 443 2527
rect 439 2521 443 2522
rect 543 2526 547 2527
rect 543 2521 547 2522
rect 591 2526 595 2527
rect 591 2521 595 2522
rect 671 2526 675 2527
rect 671 2521 675 2522
rect 735 2526 739 2527
rect 735 2521 739 2522
rect 799 2526 803 2527
rect 799 2521 803 2522
rect 871 2526 875 2527
rect 871 2521 875 2522
rect 919 2526 923 2527
rect 919 2521 923 2522
rect 1007 2526 1011 2527
rect 1007 2521 1011 2522
rect 1039 2526 1043 2527
rect 1039 2521 1043 2522
rect 1143 2526 1147 2527
rect 1143 2521 1147 2522
rect 1167 2526 1171 2527
rect 1167 2521 1171 2522
rect 1279 2526 1283 2527
rect 1279 2521 1283 2522
rect 1823 2526 1827 2527
rect 1823 2521 1827 2522
rect 112 2506 114 2521
rect 136 2516 138 2521
rect 280 2516 282 2521
rect 440 2516 442 2521
rect 592 2516 594 2521
rect 736 2516 738 2521
rect 872 2516 874 2521
rect 1008 2516 1010 2521
rect 1144 2516 1146 2521
rect 1280 2516 1282 2521
rect 134 2515 140 2516
rect 134 2511 135 2515
rect 139 2511 140 2515
rect 134 2510 140 2511
rect 278 2515 284 2516
rect 278 2511 279 2515
rect 283 2511 284 2515
rect 278 2510 284 2511
rect 438 2515 444 2516
rect 438 2511 439 2515
rect 443 2511 444 2515
rect 438 2510 444 2511
rect 590 2515 596 2516
rect 590 2511 591 2515
rect 595 2511 596 2515
rect 590 2510 596 2511
rect 734 2515 740 2516
rect 734 2511 735 2515
rect 739 2511 740 2515
rect 734 2510 740 2511
rect 870 2515 876 2516
rect 870 2511 871 2515
rect 875 2511 876 2515
rect 870 2510 876 2511
rect 1006 2515 1012 2516
rect 1006 2511 1007 2515
rect 1011 2511 1012 2515
rect 1006 2510 1012 2511
rect 1142 2515 1148 2516
rect 1142 2511 1143 2515
rect 1147 2511 1148 2515
rect 1142 2510 1148 2511
rect 1278 2515 1284 2516
rect 1278 2511 1279 2515
rect 1283 2511 1284 2515
rect 1278 2510 1284 2511
rect 1824 2506 1826 2521
rect 1864 2507 1866 2535
rect 1894 2527 1900 2528
rect 1894 2523 1895 2527
rect 1899 2523 1900 2527
rect 1894 2522 1900 2523
rect 1998 2527 2004 2528
rect 1998 2523 1999 2527
rect 2003 2523 2004 2527
rect 1998 2522 2004 2523
rect 2118 2527 2124 2528
rect 2118 2523 2119 2527
rect 2123 2523 2124 2527
rect 2118 2522 2124 2523
rect 2238 2527 2244 2528
rect 2238 2523 2239 2527
rect 2243 2523 2244 2527
rect 2238 2522 2244 2523
rect 2358 2527 2364 2528
rect 2358 2523 2359 2527
rect 2363 2523 2364 2527
rect 2358 2522 2364 2523
rect 2478 2527 2484 2528
rect 2478 2523 2479 2527
rect 2483 2523 2484 2527
rect 2478 2522 2484 2523
rect 2598 2527 2604 2528
rect 2598 2523 2599 2527
rect 2603 2523 2604 2527
rect 2598 2522 2604 2523
rect 2718 2527 2724 2528
rect 2718 2523 2719 2527
rect 2723 2523 2724 2527
rect 2718 2522 2724 2523
rect 2838 2527 2844 2528
rect 2838 2523 2839 2527
rect 2843 2523 2844 2527
rect 2838 2522 2844 2523
rect 1896 2507 1898 2522
rect 2000 2507 2002 2522
rect 2120 2507 2122 2522
rect 2240 2507 2242 2522
rect 2360 2507 2362 2522
rect 2480 2507 2482 2522
rect 2600 2507 2602 2522
rect 2720 2507 2722 2522
rect 2840 2507 2842 2522
rect 3576 2507 3578 2535
rect 1863 2506 1867 2507
rect 110 2505 116 2506
rect 110 2501 111 2505
rect 115 2501 116 2505
rect 110 2500 116 2501
rect 1822 2505 1828 2506
rect 1822 2501 1823 2505
rect 1827 2501 1828 2505
rect 1863 2501 1867 2502
rect 1895 2506 1899 2507
rect 1895 2501 1899 2502
rect 1999 2506 2003 2507
rect 1999 2501 2003 2502
rect 2031 2506 2035 2507
rect 2031 2501 2035 2502
rect 2119 2506 2123 2507
rect 2119 2501 2123 2502
rect 2191 2506 2195 2507
rect 2191 2501 2195 2502
rect 2239 2506 2243 2507
rect 2239 2501 2243 2502
rect 2343 2506 2347 2507
rect 2343 2501 2347 2502
rect 2359 2506 2363 2507
rect 2359 2501 2363 2502
rect 2479 2506 2483 2507
rect 2479 2501 2483 2502
rect 2487 2506 2491 2507
rect 2487 2501 2491 2502
rect 2599 2506 2603 2507
rect 2599 2501 2603 2502
rect 2623 2506 2627 2507
rect 2623 2501 2627 2502
rect 2719 2506 2723 2507
rect 2719 2501 2723 2502
rect 2751 2506 2755 2507
rect 2751 2501 2755 2502
rect 2839 2506 2843 2507
rect 2839 2501 2843 2502
rect 2879 2506 2883 2507
rect 2879 2501 2883 2502
rect 3015 2506 3019 2507
rect 3015 2501 3019 2502
rect 3575 2506 3579 2507
rect 3575 2501 3579 2502
rect 1822 2500 1828 2501
rect 110 2488 116 2489
rect 110 2484 111 2488
rect 115 2484 116 2488
rect 110 2483 116 2484
rect 1822 2488 1828 2489
rect 1822 2484 1823 2488
rect 1827 2484 1828 2488
rect 1822 2483 1828 2484
rect 112 2459 114 2483
rect 142 2475 148 2476
rect 142 2471 143 2475
rect 147 2471 148 2475
rect 142 2470 148 2471
rect 286 2475 292 2476
rect 286 2471 287 2475
rect 291 2471 292 2475
rect 286 2470 292 2471
rect 446 2475 452 2476
rect 446 2471 447 2475
rect 451 2471 452 2475
rect 446 2470 452 2471
rect 598 2475 604 2476
rect 598 2471 599 2475
rect 603 2471 604 2475
rect 598 2470 604 2471
rect 742 2475 748 2476
rect 742 2471 743 2475
rect 747 2471 748 2475
rect 742 2470 748 2471
rect 878 2475 884 2476
rect 878 2471 879 2475
rect 883 2471 884 2475
rect 878 2470 884 2471
rect 1014 2475 1020 2476
rect 1014 2471 1015 2475
rect 1019 2471 1020 2475
rect 1014 2470 1020 2471
rect 1150 2475 1156 2476
rect 1150 2471 1151 2475
rect 1155 2471 1156 2475
rect 1150 2470 1156 2471
rect 1286 2475 1292 2476
rect 1286 2471 1287 2475
rect 1291 2471 1292 2475
rect 1286 2470 1292 2471
rect 144 2459 146 2470
rect 288 2459 290 2470
rect 448 2459 450 2470
rect 600 2459 602 2470
rect 744 2459 746 2470
rect 880 2459 882 2470
rect 1016 2459 1018 2470
rect 1152 2459 1154 2470
rect 1288 2459 1290 2470
rect 1824 2459 1826 2483
rect 1864 2477 1866 2501
rect 1896 2490 1898 2501
rect 2032 2490 2034 2501
rect 2192 2490 2194 2501
rect 2344 2490 2346 2501
rect 2488 2490 2490 2501
rect 2624 2490 2626 2501
rect 2752 2490 2754 2501
rect 2880 2490 2882 2501
rect 3016 2490 3018 2501
rect 1894 2489 1900 2490
rect 1894 2485 1895 2489
rect 1899 2485 1900 2489
rect 1894 2484 1900 2485
rect 2030 2489 2036 2490
rect 2030 2485 2031 2489
rect 2035 2485 2036 2489
rect 2030 2484 2036 2485
rect 2190 2489 2196 2490
rect 2190 2485 2191 2489
rect 2195 2485 2196 2489
rect 2190 2484 2196 2485
rect 2342 2489 2348 2490
rect 2342 2485 2343 2489
rect 2347 2485 2348 2489
rect 2342 2484 2348 2485
rect 2486 2489 2492 2490
rect 2486 2485 2487 2489
rect 2491 2485 2492 2489
rect 2486 2484 2492 2485
rect 2622 2489 2628 2490
rect 2622 2485 2623 2489
rect 2627 2485 2628 2489
rect 2622 2484 2628 2485
rect 2750 2489 2756 2490
rect 2750 2485 2751 2489
rect 2755 2485 2756 2489
rect 2750 2484 2756 2485
rect 2878 2489 2884 2490
rect 2878 2485 2879 2489
rect 2883 2485 2884 2489
rect 2878 2484 2884 2485
rect 3014 2489 3020 2490
rect 3014 2485 3015 2489
rect 3019 2485 3020 2489
rect 3014 2484 3020 2485
rect 3576 2477 3578 2501
rect 1862 2476 1868 2477
rect 1862 2472 1863 2476
rect 1867 2472 1868 2476
rect 1862 2471 1868 2472
rect 3574 2476 3580 2477
rect 3574 2472 3575 2476
rect 3579 2472 3580 2476
rect 3574 2471 3580 2472
rect 1862 2459 1868 2460
rect 111 2458 115 2459
rect 111 2453 115 2454
rect 143 2458 147 2459
rect 143 2453 147 2454
rect 191 2458 195 2459
rect 191 2453 195 2454
rect 287 2458 291 2459
rect 287 2453 291 2454
rect 319 2458 323 2459
rect 319 2453 323 2454
rect 447 2458 451 2459
rect 447 2453 451 2454
rect 455 2458 459 2459
rect 455 2453 459 2454
rect 591 2458 595 2459
rect 591 2453 595 2454
rect 599 2458 603 2459
rect 599 2453 603 2454
rect 727 2458 731 2459
rect 727 2453 731 2454
rect 743 2458 747 2459
rect 743 2453 747 2454
rect 863 2458 867 2459
rect 863 2453 867 2454
rect 879 2458 883 2459
rect 879 2453 883 2454
rect 999 2458 1003 2459
rect 999 2453 1003 2454
rect 1015 2458 1019 2459
rect 1015 2453 1019 2454
rect 1135 2458 1139 2459
rect 1135 2453 1139 2454
rect 1151 2458 1155 2459
rect 1151 2453 1155 2454
rect 1271 2458 1275 2459
rect 1271 2453 1275 2454
rect 1287 2458 1291 2459
rect 1287 2453 1291 2454
rect 1407 2458 1411 2459
rect 1407 2453 1411 2454
rect 1823 2458 1827 2459
rect 1862 2455 1863 2459
rect 1867 2455 1868 2459
rect 1862 2454 1868 2455
rect 3574 2459 3580 2460
rect 3574 2455 3575 2459
rect 3579 2455 3580 2459
rect 3574 2454 3580 2455
rect 1823 2453 1827 2454
rect 112 2429 114 2453
rect 192 2442 194 2453
rect 320 2442 322 2453
rect 456 2442 458 2453
rect 592 2442 594 2453
rect 728 2442 730 2453
rect 864 2442 866 2453
rect 1000 2442 1002 2453
rect 1136 2442 1138 2453
rect 1272 2442 1274 2453
rect 1408 2442 1410 2453
rect 190 2441 196 2442
rect 190 2437 191 2441
rect 195 2437 196 2441
rect 190 2436 196 2437
rect 318 2441 324 2442
rect 318 2437 319 2441
rect 323 2437 324 2441
rect 318 2436 324 2437
rect 454 2441 460 2442
rect 454 2437 455 2441
rect 459 2437 460 2441
rect 454 2436 460 2437
rect 590 2441 596 2442
rect 590 2437 591 2441
rect 595 2437 596 2441
rect 590 2436 596 2437
rect 726 2441 732 2442
rect 726 2437 727 2441
rect 731 2437 732 2441
rect 726 2436 732 2437
rect 862 2441 868 2442
rect 862 2437 863 2441
rect 867 2437 868 2441
rect 862 2436 868 2437
rect 998 2441 1004 2442
rect 998 2437 999 2441
rect 1003 2437 1004 2441
rect 998 2436 1004 2437
rect 1134 2441 1140 2442
rect 1134 2437 1135 2441
rect 1139 2437 1140 2441
rect 1134 2436 1140 2437
rect 1270 2441 1276 2442
rect 1270 2437 1271 2441
rect 1275 2437 1276 2441
rect 1270 2436 1276 2437
rect 1406 2441 1412 2442
rect 1406 2437 1407 2441
rect 1411 2437 1412 2441
rect 1406 2436 1412 2437
rect 1824 2429 1826 2453
rect 1864 2439 1866 2454
rect 1886 2449 1892 2450
rect 1886 2445 1887 2449
rect 1891 2445 1892 2449
rect 1886 2444 1892 2445
rect 2022 2449 2028 2450
rect 2022 2445 2023 2449
rect 2027 2445 2028 2449
rect 2022 2444 2028 2445
rect 2182 2449 2188 2450
rect 2182 2445 2183 2449
rect 2187 2445 2188 2449
rect 2182 2444 2188 2445
rect 2334 2449 2340 2450
rect 2334 2445 2335 2449
rect 2339 2445 2340 2449
rect 2334 2444 2340 2445
rect 2478 2449 2484 2450
rect 2478 2445 2479 2449
rect 2483 2445 2484 2449
rect 2478 2444 2484 2445
rect 2614 2449 2620 2450
rect 2614 2445 2615 2449
rect 2619 2445 2620 2449
rect 2614 2444 2620 2445
rect 2742 2449 2748 2450
rect 2742 2445 2743 2449
rect 2747 2445 2748 2449
rect 2742 2444 2748 2445
rect 2870 2449 2876 2450
rect 2870 2445 2871 2449
rect 2875 2445 2876 2449
rect 2870 2444 2876 2445
rect 3006 2449 3012 2450
rect 3006 2445 3007 2449
rect 3011 2445 3012 2449
rect 3006 2444 3012 2445
rect 1888 2439 1890 2444
rect 2024 2439 2026 2444
rect 2184 2439 2186 2444
rect 2336 2439 2338 2444
rect 2480 2439 2482 2444
rect 2616 2439 2618 2444
rect 2744 2439 2746 2444
rect 2872 2439 2874 2444
rect 3008 2439 3010 2444
rect 3576 2439 3578 2454
rect 1863 2438 1867 2439
rect 1863 2433 1867 2434
rect 1887 2438 1891 2439
rect 1887 2433 1891 2434
rect 2015 2438 2019 2439
rect 2015 2433 2019 2434
rect 2023 2438 2027 2439
rect 2023 2433 2027 2434
rect 2175 2438 2179 2439
rect 2175 2433 2179 2434
rect 2183 2438 2187 2439
rect 2183 2433 2187 2434
rect 2335 2438 2339 2439
rect 2335 2433 2339 2434
rect 2479 2438 2483 2439
rect 2479 2433 2483 2434
rect 2495 2438 2499 2439
rect 2495 2433 2499 2434
rect 2615 2438 2619 2439
rect 2615 2433 2619 2434
rect 2647 2438 2651 2439
rect 2647 2433 2651 2434
rect 2743 2438 2747 2439
rect 2743 2433 2747 2434
rect 2799 2438 2803 2439
rect 2799 2433 2803 2434
rect 2871 2438 2875 2439
rect 2871 2433 2875 2434
rect 2951 2438 2955 2439
rect 2951 2433 2955 2434
rect 3007 2438 3011 2439
rect 3007 2433 3011 2434
rect 3111 2438 3115 2439
rect 3111 2433 3115 2434
rect 3575 2438 3579 2439
rect 3575 2433 3579 2434
rect 110 2428 116 2429
rect 110 2424 111 2428
rect 115 2424 116 2428
rect 110 2423 116 2424
rect 1822 2428 1828 2429
rect 1822 2424 1823 2428
rect 1827 2424 1828 2428
rect 1822 2423 1828 2424
rect 1864 2418 1866 2433
rect 1888 2428 1890 2433
rect 2016 2428 2018 2433
rect 2176 2428 2178 2433
rect 2336 2428 2338 2433
rect 2496 2428 2498 2433
rect 2648 2428 2650 2433
rect 2800 2428 2802 2433
rect 2952 2428 2954 2433
rect 3112 2428 3114 2433
rect 1886 2427 1892 2428
rect 1886 2423 1887 2427
rect 1891 2423 1892 2427
rect 1886 2422 1892 2423
rect 2014 2427 2020 2428
rect 2014 2423 2015 2427
rect 2019 2423 2020 2427
rect 2014 2422 2020 2423
rect 2174 2427 2180 2428
rect 2174 2423 2175 2427
rect 2179 2423 2180 2427
rect 2174 2422 2180 2423
rect 2334 2427 2340 2428
rect 2334 2423 2335 2427
rect 2339 2423 2340 2427
rect 2334 2422 2340 2423
rect 2494 2427 2500 2428
rect 2494 2423 2495 2427
rect 2499 2423 2500 2427
rect 2494 2422 2500 2423
rect 2646 2427 2652 2428
rect 2646 2423 2647 2427
rect 2651 2423 2652 2427
rect 2646 2422 2652 2423
rect 2798 2427 2804 2428
rect 2798 2423 2799 2427
rect 2803 2423 2804 2427
rect 2798 2422 2804 2423
rect 2950 2427 2956 2428
rect 2950 2423 2951 2427
rect 2955 2423 2956 2427
rect 2950 2422 2956 2423
rect 3110 2427 3116 2428
rect 3110 2423 3111 2427
rect 3115 2423 3116 2427
rect 3110 2422 3116 2423
rect 3576 2418 3578 2433
rect 1862 2417 1868 2418
rect 1862 2413 1863 2417
rect 1867 2413 1868 2417
rect 1862 2412 1868 2413
rect 3574 2417 3580 2418
rect 3574 2413 3575 2417
rect 3579 2413 3580 2417
rect 3574 2412 3580 2413
rect 110 2411 116 2412
rect 110 2407 111 2411
rect 115 2407 116 2411
rect 110 2406 116 2407
rect 1822 2411 1828 2412
rect 1822 2407 1823 2411
rect 1827 2407 1828 2411
rect 1822 2406 1828 2407
rect 112 2379 114 2406
rect 182 2401 188 2402
rect 182 2397 183 2401
rect 187 2397 188 2401
rect 182 2396 188 2397
rect 310 2401 316 2402
rect 310 2397 311 2401
rect 315 2397 316 2401
rect 310 2396 316 2397
rect 446 2401 452 2402
rect 446 2397 447 2401
rect 451 2397 452 2401
rect 446 2396 452 2397
rect 582 2401 588 2402
rect 582 2397 583 2401
rect 587 2397 588 2401
rect 582 2396 588 2397
rect 718 2401 724 2402
rect 718 2397 719 2401
rect 723 2397 724 2401
rect 718 2396 724 2397
rect 854 2401 860 2402
rect 854 2397 855 2401
rect 859 2397 860 2401
rect 854 2396 860 2397
rect 990 2401 996 2402
rect 990 2397 991 2401
rect 995 2397 996 2401
rect 990 2396 996 2397
rect 1126 2401 1132 2402
rect 1126 2397 1127 2401
rect 1131 2397 1132 2401
rect 1126 2396 1132 2397
rect 1262 2401 1268 2402
rect 1262 2397 1263 2401
rect 1267 2397 1268 2401
rect 1262 2396 1268 2397
rect 1398 2401 1404 2402
rect 1398 2397 1399 2401
rect 1403 2397 1404 2401
rect 1398 2396 1404 2397
rect 184 2379 186 2396
rect 312 2379 314 2396
rect 448 2379 450 2396
rect 584 2379 586 2396
rect 720 2379 722 2396
rect 856 2379 858 2396
rect 992 2379 994 2396
rect 1128 2379 1130 2396
rect 1264 2379 1266 2396
rect 1400 2379 1402 2396
rect 1824 2379 1826 2406
rect 1862 2400 1868 2401
rect 1862 2396 1863 2400
rect 1867 2396 1868 2400
rect 1862 2395 1868 2396
rect 3574 2400 3580 2401
rect 3574 2396 3575 2400
rect 3579 2396 3580 2400
rect 3574 2395 3580 2396
rect 111 2378 115 2379
rect 111 2373 115 2374
rect 159 2378 163 2379
rect 159 2373 163 2374
rect 183 2378 187 2379
rect 183 2373 187 2374
rect 247 2378 251 2379
rect 247 2373 251 2374
rect 311 2378 315 2379
rect 311 2373 315 2374
rect 335 2378 339 2379
rect 335 2373 339 2374
rect 439 2378 443 2379
rect 439 2373 443 2374
rect 447 2378 451 2379
rect 447 2373 451 2374
rect 559 2378 563 2379
rect 559 2373 563 2374
rect 583 2378 587 2379
rect 583 2373 587 2374
rect 687 2378 691 2379
rect 687 2373 691 2374
rect 719 2378 723 2379
rect 719 2373 723 2374
rect 815 2378 819 2379
rect 815 2373 819 2374
rect 855 2378 859 2379
rect 855 2373 859 2374
rect 951 2378 955 2379
rect 951 2373 955 2374
rect 991 2378 995 2379
rect 991 2373 995 2374
rect 1079 2378 1083 2379
rect 1079 2373 1083 2374
rect 1127 2378 1131 2379
rect 1127 2373 1131 2374
rect 1207 2378 1211 2379
rect 1207 2373 1211 2374
rect 1263 2378 1267 2379
rect 1263 2373 1267 2374
rect 1327 2378 1331 2379
rect 1327 2373 1331 2374
rect 1399 2378 1403 2379
rect 1399 2373 1403 2374
rect 1455 2378 1459 2379
rect 1455 2373 1459 2374
rect 1583 2378 1587 2379
rect 1583 2373 1587 2374
rect 1823 2378 1827 2379
rect 1823 2373 1827 2374
rect 112 2358 114 2373
rect 160 2368 162 2373
rect 248 2368 250 2373
rect 336 2368 338 2373
rect 440 2368 442 2373
rect 560 2368 562 2373
rect 688 2368 690 2373
rect 816 2368 818 2373
rect 952 2368 954 2373
rect 1080 2368 1082 2373
rect 1208 2368 1210 2373
rect 1328 2368 1330 2373
rect 1456 2368 1458 2373
rect 1584 2368 1586 2373
rect 158 2367 164 2368
rect 158 2363 159 2367
rect 163 2363 164 2367
rect 158 2362 164 2363
rect 246 2367 252 2368
rect 246 2363 247 2367
rect 251 2363 252 2367
rect 246 2362 252 2363
rect 334 2367 340 2368
rect 334 2363 335 2367
rect 339 2363 340 2367
rect 334 2362 340 2363
rect 438 2367 444 2368
rect 438 2363 439 2367
rect 443 2363 444 2367
rect 438 2362 444 2363
rect 558 2367 564 2368
rect 558 2363 559 2367
rect 563 2363 564 2367
rect 558 2362 564 2363
rect 686 2367 692 2368
rect 686 2363 687 2367
rect 691 2363 692 2367
rect 686 2362 692 2363
rect 814 2367 820 2368
rect 814 2363 815 2367
rect 819 2363 820 2367
rect 814 2362 820 2363
rect 950 2367 956 2368
rect 950 2363 951 2367
rect 955 2363 956 2367
rect 950 2362 956 2363
rect 1078 2367 1084 2368
rect 1078 2363 1079 2367
rect 1083 2363 1084 2367
rect 1078 2362 1084 2363
rect 1206 2367 1212 2368
rect 1206 2363 1207 2367
rect 1211 2363 1212 2367
rect 1206 2362 1212 2363
rect 1326 2367 1332 2368
rect 1326 2363 1327 2367
rect 1331 2363 1332 2367
rect 1326 2362 1332 2363
rect 1454 2367 1460 2368
rect 1454 2363 1455 2367
rect 1459 2363 1460 2367
rect 1454 2362 1460 2363
rect 1582 2367 1588 2368
rect 1582 2363 1583 2367
rect 1587 2363 1588 2367
rect 1582 2362 1588 2363
rect 1824 2358 1826 2373
rect 1864 2367 1866 2395
rect 1894 2387 1900 2388
rect 1894 2383 1895 2387
rect 1899 2383 1900 2387
rect 1894 2382 1900 2383
rect 2022 2387 2028 2388
rect 2022 2383 2023 2387
rect 2027 2383 2028 2387
rect 2022 2382 2028 2383
rect 2182 2387 2188 2388
rect 2182 2383 2183 2387
rect 2187 2383 2188 2387
rect 2182 2382 2188 2383
rect 2342 2387 2348 2388
rect 2342 2383 2343 2387
rect 2347 2383 2348 2387
rect 2342 2382 2348 2383
rect 2502 2387 2508 2388
rect 2502 2383 2503 2387
rect 2507 2383 2508 2387
rect 2502 2382 2508 2383
rect 2654 2387 2660 2388
rect 2654 2383 2655 2387
rect 2659 2383 2660 2387
rect 2654 2382 2660 2383
rect 2806 2387 2812 2388
rect 2806 2383 2807 2387
rect 2811 2383 2812 2387
rect 2806 2382 2812 2383
rect 2958 2387 2964 2388
rect 2958 2383 2959 2387
rect 2963 2383 2964 2387
rect 2958 2382 2964 2383
rect 3118 2387 3124 2388
rect 3118 2383 3119 2387
rect 3123 2383 3124 2387
rect 3118 2382 3124 2383
rect 1896 2367 1898 2382
rect 2024 2367 2026 2382
rect 2184 2367 2186 2382
rect 2344 2367 2346 2382
rect 2504 2367 2506 2382
rect 2656 2367 2658 2382
rect 2808 2367 2810 2382
rect 2960 2367 2962 2382
rect 3120 2367 3122 2382
rect 3576 2367 3578 2395
rect 1863 2366 1867 2367
rect 1863 2361 1867 2362
rect 1895 2366 1899 2367
rect 1895 2361 1899 2362
rect 1927 2366 1931 2367
rect 1927 2361 1931 2362
rect 2023 2366 2027 2367
rect 2023 2361 2027 2362
rect 2087 2366 2091 2367
rect 2087 2361 2091 2362
rect 2183 2366 2187 2367
rect 2183 2361 2187 2362
rect 2247 2366 2251 2367
rect 2247 2361 2251 2362
rect 2343 2366 2347 2367
rect 2343 2361 2347 2362
rect 2407 2366 2411 2367
rect 2407 2361 2411 2362
rect 2503 2366 2507 2367
rect 2503 2361 2507 2362
rect 2559 2366 2563 2367
rect 2559 2361 2563 2362
rect 2655 2366 2659 2367
rect 2655 2361 2659 2362
rect 2703 2366 2707 2367
rect 2703 2361 2707 2362
rect 2807 2366 2811 2367
rect 2807 2361 2811 2362
rect 2831 2366 2835 2367
rect 2831 2361 2835 2362
rect 2951 2366 2955 2367
rect 2951 2361 2955 2362
rect 2959 2366 2963 2367
rect 2959 2361 2963 2362
rect 3071 2366 3075 2367
rect 3071 2361 3075 2362
rect 3119 2366 3123 2367
rect 3119 2361 3123 2362
rect 3183 2366 3187 2367
rect 3183 2361 3187 2362
rect 3287 2366 3291 2367
rect 3287 2361 3291 2362
rect 3399 2366 3403 2367
rect 3399 2361 3403 2362
rect 3487 2366 3491 2367
rect 3487 2361 3491 2362
rect 3575 2366 3579 2367
rect 3575 2361 3579 2362
rect 110 2357 116 2358
rect 110 2353 111 2357
rect 115 2353 116 2357
rect 110 2352 116 2353
rect 1822 2357 1828 2358
rect 1822 2353 1823 2357
rect 1827 2353 1828 2357
rect 1822 2352 1828 2353
rect 110 2340 116 2341
rect 110 2336 111 2340
rect 115 2336 116 2340
rect 110 2335 116 2336
rect 1822 2340 1828 2341
rect 1822 2336 1823 2340
rect 1827 2336 1828 2340
rect 1864 2337 1866 2361
rect 1928 2350 1930 2361
rect 2088 2350 2090 2361
rect 2248 2350 2250 2361
rect 2408 2350 2410 2361
rect 2560 2350 2562 2361
rect 2704 2350 2706 2361
rect 2832 2350 2834 2361
rect 2952 2350 2954 2361
rect 3072 2350 3074 2361
rect 3184 2350 3186 2361
rect 3288 2350 3290 2361
rect 3400 2350 3402 2361
rect 3488 2350 3490 2361
rect 1926 2349 1932 2350
rect 1926 2345 1927 2349
rect 1931 2345 1932 2349
rect 1926 2344 1932 2345
rect 2086 2349 2092 2350
rect 2086 2345 2087 2349
rect 2091 2345 2092 2349
rect 2086 2344 2092 2345
rect 2246 2349 2252 2350
rect 2246 2345 2247 2349
rect 2251 2345 2252 2349
rect 2246 2344 2252 2345
rect 2406 2349 2412 2350
rect 2406 2345 2407 2349
rect 2411 2345 2412 2349
rect 2406 2344 2412 2345
rect 2558 2349 2564 2350
rect 2558 2345 2559 2349
rect 2563 2345 2564 2349
rect 2558 2344 2564 2345
rect 2702 2349 2708 2350
rect 2702 2345 2703 2349
rect 2707 2345 2708 2349
rect 2702 2344 2708 2345
rect 2830 2349 2836 2350
rect 2830 2345 2831 2349
rect 2835 2345 2836 2349
rect 2830 2344 2836 2345
rect 2950 2349 2956 2350
rect 2950 2345 2951 2349
rect 2955 2345 2956 2349
rect 2950 2344 2956 2345
rect 3070 2349 3076 2350
rect 3070 2345 3071 2349
rect 3075 2345 3076 2349
rect 3070 2344 3076 2345
rect 3182 2349 3188 2350
rect 3182 2345 3183 2349
rect 3187 2345 3188 2349
rect 3182 2344 3188 2345
rect 3286 2349 3292 2350
rect 3286 2345 3287 2349
rect 3291 2345 3292 2349
rect 3286 2344 3292 2345
rect 3398 2349 3404 2350
rect 3398 2345 3399 2349
rect 3403 2345 3404 2349
rect 3398 2344 3404 2345
rect 3486 2349 3492 2350
rect 3486 2345 3487 2349
rect 3491 2345 3492 2349
rect 3486 2344 3492 2345
rect 3576 2337 3578 2361
rect 1822 2335 1828 2336
rect 1862 2336 1868 2337
rect 112 2303 114 2335
rect 166 2327 172 2328
rect 166 2323 167 2327
rect 171 2323 172 2327
rect 166 2322 172 2323
rect 254 2327 260 2328
rect 254 2323 255 2327
rect 259 2323 260 2327
rect 254 2322 260 2323
rect 342 2327 348 2328
rect 342 2323 343 2327
rect 347 2323 348 2327
rect 342 2322 348 2323
rect 446 2327 452 2328
rect 446 2323 447 2327
rect 451 2323 452 2327
rect 446 2322 452 2323
rect 566 2327 572 2328
rect 566 2323 567 2327
rect 571 2323 572 2327
rect 566 2322 572 2323
rect 694 2327 700 2328
rect 694 2323 695 2327
rect 699 2323 700 2327
rect 694 2322 700 2323
rect 822 2327 828 2328
rect 822 2323 823 2327
rect 827 2323 828 2327
rect 822 2322 828 2323
rect 958 2327 964 2328
rect 958 2323 959 2327
rect 963 2323 964 2327
rect 958 2322 964 2323
rect 1086 2327 1092 2328
rect 1086 2323 1087 2327
rect 1091 2323 1092 2327
rect 1086 2322 1092 2323
rect 1214 2327 1220 2328
rect 1214 2323 1215 2327
rect 1219 2323 1220 2327
rect 1214 2322 1220 2323
rect 1334 2327 1340 2328
rect 1334 2323 1335 2327
rect 1339 2323 1340 2327
rect 1334 2322 1340 2323
rect 1462 2327 1468 2328
rect 1462 2323 1463 2327
rect 1467 2323 1468 2327
rect 1462 2322 1468 2323
rect 1590 2327 1596 2328
rect 1590 2323 1591 2327
rect 1595 2323 1596 2327
rect 1590 2322 1596 2323
rect 168 2303 170 2322
rect 256 2303 258 2322
rect 344 2303 346 2322
rect 448 2303 450 2322
rect 568 2303 570 2322
rect 696 2303 698 2322
rect 824 2303 826 2322
rect 960 2303 962 2322
rect 1088 2303 1090 2322
rect 1216 2303 1218 2322
rect 1336 2303 1338 2322
rect 1464 2303 1466 2322
rect 1592 2303 1594 2322
rect 1824 2303 1826 2335
rect 1862 2332 1863 2336
rect 1867 2332 1868 2336
rect 1862 2331 1868 2332
rect 3574 2336 3580 2337
rect 3574 2332 3575 2336
rect 3579 2332 3580 2336
rect 3574 2331 3580 2332
rect 1862 2319 1868 2320
rect 1862 2315 1863 2319
rect 1867 2315 1868 2319
rect 1862 2314 1868 2315
rect 3574 2319 3580 2320
rect 3574 2315 3575 2319
rect 3579 2315 3580 2319
rect 3574 2314 3580 2315
rect 111 2302 115 2303
rect 111 2297 115 2298
rect 167 2302 171 2303
rect 167 2297 171 2298
rect 255 2302 259 2303
rect 255 2297 259 2298
rect 343 2302 347 2303
rect 343 2297 347 2298
rect 447 2302 451 2303
rect 447 2297 451 2298
rect 567 2302 571 2303
rect 567 2297 571 2298
rect 695 2302 699 2303
rect 695 2297 699 2298
rect 823 2302 827 2303
rect 823 2297 827 2298
rect 863 2302 867 2303
rect 863 2297 867 2298
rect 959 2302 963 2303
rect 959 2297 963 2298
rect 1023 2302 1027 2303
rect 1023 2297 1027 2298
rect 1087 2302 1091 2303
rect 1087 2297 1091 2298
rect 1175 2302 1179 2303
rect 1175 2297 1179 2298
rect 1215 2302 1219 2303
rect 1215 2297 1219 2298
rect 1319 2302 1323 2303
rect 1319 2297 1323 2298
rect 1335 2302 1339 2303
rect 1335 2297 1339 2298
rect 1463 2302 1467 2303
rect 1463 2297 1467 2298
rect 1591 2302 1595 2303
rect 1591 2297 1595 2298
rect 1599 2302 1603 2303
rect 1599 2297 1603 2298
rect 1735 2302 1739 2303
rect 1735 2297 1739 2298
rect 1823 2302 1827 2303
rect 1823 2297 1827 2298
rect 112 2273 114 2297
rect 696 2286 698 2297
rect 864 2286 866 2297
rect 1024 2286 1026 2297
rect 1176 2286 1178 2297
rect 1320 2286 1322 2297
rect 1464 2286 1466 2297
rect 1600 2286 1602 2297
rect 1736 2286 1738 2297
rect 694 2285 700 2286
rect 694 2281 695 2285
rect 699 2281 700 2285
rect 694 2280 700 2281
rect 862 2285 868 2286
rect 862 2281 863 2285
rect 867 2281 868 2285
rect 862 2280 868 2281
rect 1022 2285 1028 2286
rect 1022 2281 1023 2285
rect 1027 2281 1028 2285
rect 1022 2280 1028 2281
rect 1174 2285 1180 2286
rect 1174 2281 1175 2285
rect 1179 2281 1180 2285
rect 1174 2280 1180 2281
rect 1318 2285 1324 2286
rect 1318 2281 1319 2285
rect 1323 2281 1324 2285
rect 1318 2280 1324 2281
rect 1462 2285 1468 2286
rect 1462 2281 1463 2285
rect 1467 2281 1468 2285
rect 1462 2280 1468 2281
rect 1598 2285 1604 2286
rect 1598 2281 1599 2285
rect 1603 2281 1604 2285
rect 1598 2280 1604 2281
rect 1734 2285 1740 2286
rect 1734 2281 1735 2285
rect 1739 2281 1740 2285
rect 1734 2280 1740 2281
rect 1824 2273 1826 2297
rect 1864 2295 1866 2314
rect 1918 2309 1924 2310
rect 1918 2305 1919 2309
rect 1923 2305 1924 2309
rect 1918 2304 1924 2305
rect 2078 2309 2084 2310
rect 2078 2305 2079 2309
rect 2083 2305 2084 2309
rect 2078 2304 2084 2305
rect 2238 2309 2244 2310
rect 2238 2305 2239 2309
rect 2243 2305 2244 2309
rect 2238 2304 2244 2305
rect 2398 2309 2404 2310
rect 2398 2305 2399 2309
rect 2403 2305 2404 2309
rect 2398 2304 2404 2305
rect 2550 2309 2556 2310
rect 2550 2305 2551 2309
rect 2555 2305 2556 2309
rect 2550 2304 2556 2305
rect 2694 2309 2700 2310
rect 2694 2305 2695 2309
rect 2699 2305 2700 2309
rect 2694 2304 2700 2305
rect 2822 2309 2828 2310
rect 2822 2305 2823 2309
rect 2827 2305 2828 2309
rect 2822 2304 2828 2305
rect 2942 2309 2948 2310
rect 2942 2305 2943 2309
rect 2947 2305 2948 2309
rect 2942 2304 2948 2305
rect 3062 2309 3068 2310
rect 3062 2305 3063 2309
rect 3067 2305 3068 2309
rect 3062 2304 3068 2305
rect 3174 2309 3180 2310
rect 3174 2305 3175 2309
rect 3179 2305 3180 2309
rect 3174 2304 3180 2305
rect 3278 2309 3284 2310
rect 3278 2305 3279 2309
rect 3283 2305 3284 2309
rect 3278 2304 3284 2305
rect 3390 2309 3396 2310
rect 3390 2305 3391 2309
rect 3395 2305 3396 2309
rect 3390 2304 3396 2305
rect 3478 2309 3484 2310
rect 3478 2305 3479 2309
rect 3483 2305 3484 2309
rect 3478 2304 3484 2305
rect 1920 2295 1922 2304
rect 2080 2295 2082 2304
rect 2240 2295 2242 2304
rect 2400 2295 2402 2304
rect 2552 2295 2554 2304
rect 2696 2295 2698 2304
rect 2824 2295 2826 2304
rect 2944 2295 2946 2304
rect 3064 2295 3066 2304
rect 3176 2295 3178 2304
rect 3280 2295 3282 2304
rect 3392 2295 3394 2304
rect 3480 2295 3482 2304
rect 3576 2295 3578 2314
rect 1863 2294 1867 2295
rect 1863 2289 1867 2290
rect 1919 2294 1923 2295
rect 1919 2289 1923 2290
rect 1975 2294 1979 2295
rect 1975 2289 1979 2290
rect 2079 2294 2083 2295
rect 2079 2289 2083 2290
rect 2143 2294 2147 2295
rect 2143 2289 2147 2290
rect 2239 2294 2243 2295
rect 2239 2289 2243 2290
rect 2311 2294 2315 2295
rect 2311 2289 2315 2290
rect 2399 2294 2403 2295
rect 2399 2289 2403 2290
rect 2479 2294 2483 2295
rect 2479 2289 2483 2290
rect 2551 2294 2555 2295
rect 2551 2289 2555 2290
rect 2639 2294 2643 2295
rect 2639 2289 2643 2290
rect 2695 2294 2699 2295
rect 2695 2289 2699 2290
rect 2783 2294 2787 2295
rect 2783 2289 2787 2290
rect 2823 2294 2827 2295
rect 2823 2289 2827 2290
rect 2919 2294 2923 2295
rect 2919 2289 2923 2290
rect 2943 2294 2947 2295
rect 2943 2289 2947 2290
rect 3039 2294 3043 2295
rect 3039 2289 3043 2290
rect 3063 2294 3067 2295
rect 3063 2289 3067 2290
rect 3159 2294 3163 2295
rect 3159 2289 3163 2290
rect 3175 2294 3179 2295
rect 3175 2289 3179 2290
rect 3271 2294 3275 2295
rect 3271 2289 3275 2290
rect 3279 2294 3283 2295
rect 3279 2289 3283 2290
rect 3383 2294 3387 2295
rect 3383 2289 3387 2290
rect 3391 2294 3395 2295
rect 3391 2289 3395 2290
rect 3479 2294 3483 2295
rect 3479 2289 3483 2290
rect 3575 2294 3579 2295
rect 3575 2289 3579 2290
rect 1864 2274 1866 2289
rect 1976 2284 1978 2289
rect 2144 2284 2146 2289
rect 2312 2284 2314 2289
rect 2480 2284 2482 2289
rect 2640 2284 2642 2289
rect 2784 2284 2786 2289
rect 2920 2284 2922 2289
rect 3040 2284 3042 2289
rect 3160 2284 3162 2289
rect 3272 2284 3274 2289
rect 3384 2284 3386 2289
rect 3480 2284 3482 2289
rect 1974 2283 1980 2284
rect 1974 2279 1975 2283
rect 1979 2279 1980 2283
rect 1974 2278 1980 2279
rect 2142 2283 2148 2284
rect 2142 2279 2143 2283
rect 2147 2279 2148 2283
rect 2142 2278 2148 2279
rect 2310 2283 2316 2284
rect 2310 2279 2311 2283
rect 2315 2279 2316 2283
rect 2310 2278 2316 2279
rect 2478 2283 2484 2284
rect 2478 2279 2479 2283
rect 2483 2279 2484 2283
rect 2478 2278 2484 2279
rect 2638 2283 2644 2284
rect 2638 2279 2639 2283
rect 2643 2279 2644 2283
rect 2638 2278 2644 2279
rect 2782 2283 2788 2284
rect 2782 2279 2783 2283
rect 2787 2279 2788 2283
rect 2782 2278 2788 2279
rect 2918 2283 2924 2284
rect 2918 2279 2919 2283
rect 2923 2279 2924 2283
rect 2918 2278 2924 2279
rect 3038 2283 3044 2284
rect 3038 2279 3039 2283
rect 3043 2279 3044 2283
rect 3038 2278 3044 2279
rect 3158 2283 3164 2284
rect 3158 2279 3159 2283
rect 3163 2279 3164 2283
rect 3158 2278 3164 2279
rect 3270 2283 3276 2284
rect 3270 2279 3271 2283
rect 3275 2279 3276 2283
rect 3270 2278 3276 2279
rect 3382 2283 3388 2284
rect 3382 2279 3383 2283
rect 3387 2279 3388 2283
rect 3382 2278 3388 2279
rect 3478 2283 3484 2284
rect 3478 2279 3479 2283
rect 3483 2279 3484 2283
rect 3478 2278 3484 2279
rect 3576 2274 3578 2289
rect 1862 2273 1868 2274
rect 110 2272 116 2273
rect 110 2268 111 2272
rect 115 2268 116 2272
rect 110 2267 116 2268
rect 1822 2272 1828 2273
rect 1822 2268 1823 2272
rect 1827 2268 1828 2272
rect 1862 2269 1863 2273
rect 1867 2269 1868 2273
rect 1862 2268 1868 2269
rect 3574 2273 3580 2274
rect 3574 2269 3575 2273
rect 3579 2269 3580 2273
rect 3574 2268 3580 2269
rect 1822 2267 1828 2268
rect 1862 2256 1868 2257
rect 110 2255 116 2256
rect 110 2251 111 2255
rect 115 2251 116 2255
rect 110 2250 116 2251
rect 1822 2255 1828 2256
rect 1822 2251 1823 2255
rect 1827 2251 1828 2255
rect 1862 2252 1863 2256
rect 1867 2252 1868 2256
rect 1862 2251 1868 2252
rect 3574 2256 3580 2257
rect 3574 2252 3575 2256
rect 3579 2252 3580 2256
rect 3574 2251 3580 2252
rect 1822 2250 1828 2251
rect 112 2227 114 2250
rect 686 2245 692 2246
rect 686 2241 687 2245
rect 691 2241 692 2245
rect 686 2240 692 2241
rect 854 2245 860 2246
rect 854 2241 855 2245
rect 859 2241 860 2245
rect 854 2240 860 2241
rect 1014 2245 1020 2246
rect 1014 2241 1015 2245
rect 1019 2241 1020 2245
rect 1014 2240 1020 2241
rect 1166 2245 1172 2246
rect 1166 2241 1167 2245
rect 1171 2241 1172 2245
rect 1166 2240 1172 2241
rect 1310 2245 1316 2246
rect 1310 2241 1311 2245
rect 1315 2241 1316 2245
rect 1310 2240 1316 2241
rect 1454 2245 1460 2246
rect 1454 2241 1455 2245
rect 1459 2241 1460 2245
rect 1454 2240 1460 2241
rect 1590 2245 1596 2246
rect 1590 2241 1591 2245
rect 1595 2241 1596 2245
rect 1590 2240 1596 2241
rect 1726 2245 1732 2246
rect 1726 2241 1727 2245
rect 1731 2241 1732 2245
rect 1726 2240 1732 2241
rect 688 2227 690 2240
rect 856 2227 858 2240
rect 1016 2227 1018 2240
rect 1168 2227 1170 2240
rect 1312 2227 1314 2240
rect 1456 2227 1458 2240
rect 1592 2227 1594 2240
rect 1728 2227 1730 2240
rect 1824 2227 1826 2250
rect 1864 2227 1866 2251
rect 1982 2243 1988 2244
rect 1982 2239 1983 2243
rect 1987 2239 1988 2243
rect 1982 2238 1988 2239
rect 2150 2243 2156 2244
rect 2150 2239 2151 2243
rect 2155 2239 2156 2243
rect 2150 2238 2156 2239
rect 2318 2243 2324 2244
rect 2318 2239 2319 2243
rect 2323 2239 2324 2243
rect 2318 2238 2324 2239
rect 2486 2243 2492 2244
rect 2486 2239 2487 2243
rect 2491 2239 2492 2243
rect 2486 2238 2492 2239
rect 2646 2243 2652 2244
rect 2646 2239 2647 2243
rect 2651 2239 2652 2243
rect 2646 2238 2652 2239
rect 2790 2243 2796 2244
rect 2790 2239 2791 2243
rect 2795 2239 2796 2243
rect 2790 2238 2796 2239
rect 2926 2243 2932 2244
rect 2926 2239 2927 2243
rect 2931 2239 2932 2243
rect 2926 2238 2932 2239
rect 3046 2243 3052 2244
rect 3046 2239 3047 2243
rect 3051 2239 3052 2243
rect 3046 2238 3052 2239
rect 3166 2243 3172 2244
rect 3166 2239 3167 2243
rect 3171 2239 3172 2243
rect 3166 2238 3172 2239
rect 3278 2243 3284 2244
rect 3278 2239 3279 2243
rect 3283 2239 3284 2243
rect 3278 2238 3284 2239
rect 3390 2243 3396 2244
rect 3390 2239 3391 2243
rect 3395 2239 3396 2243
rect 3390 2238 3396 2239
rect 3486 2243 3492 2244
rect 3486 2239 3487 2243
rect 3491 2239 3492 2243
rect 3486 2238 3492 2239
rect 1984 2227 1986 2238
rect 2152 2227 2154 2238
rect 2320 2227 2322 2238
rect 2488 2227 2490 2238
rect 2648 2227 2650 2238
rect 2792 2227 2794 2238
rect 2928 2227 2930 2238
rect 3048 2227 3050 2238
rect 3168 2227 3170 2238
rect 3280 2227 3282 2238
rect 3392 2227 3394 2238
rect 3488 2227 3490 2238
rect 3576 2227 3578 2251
rect 111 2226 115 2227
rect 111 2221 115 2222
rect 535 2226 539 2227
rect 535 2221 539 2222
rect 687 2226 691 2227
rect 687 2221 691 2222
rect 719 2226 723 2227
rect 719 2221 723 2222
rect 855 2226 859 2227
rect 855 2221 859 2222
rect 895 2226 899 2227
rect 895 2221 899 2222
rect 1015 2226 1019 2227
rect 1015 2221 1019 2222
rect 1071 2226 1075 2227
rect 1071 2221 1075 2222
rect 1167 2226 1171 2227
rect 1167 2221 1171 2222
rect 1239 2226 1243 2227
rect 1239 2221 1243 2222
rect 1311 2226 1315 2227
rect 1311 2221 1315 2222
rect 1407 2226 1411 2227
rect 1407 2221 1411 2222
rect 1455 2226 1459 2227
rect 1455 2221 1459 2222
rect 1575 2226 1579 2227
rect 1575 2221 1579 2222
rect 1591 2226 1595 2227
rect 1591 2221 1595 2222
rect 1727 2226 1731 2227
rect 1727 2221 1731 2222
rect 1823 2226 1827 2227
rect 1823 2221 1827 2222
rect 1863 2226 1867 2227
rect 1863 2221 1867 2222
rect 1983 2226 1987 2227
rect 1983 2221 1987 2222
rect 2007 2226 2011 2227
rect 2007 2221 2011 2222
rect 2151 2226 2155 2227
rect 2151 2221 2155 2222
rect 2167 2226 2171 2227
rect 2167 2221 2171 2222
rect 2319 2226 2323 2227
rect 2319 2221 2323 2222
rect 2335 2226 2339 2227
rect 2335 2221 2339 2222
rect 2487 2226 2491 2227
rect 2487 2221 2491 2222
rect 2519 2226 2523 2227
rect 2519 2221 2523 2222
rect 2647 2226 2651 2227
rect 2647 2221 2651 2222
rect 2711 2226 2715 2227
rect 2711 2221 2715 2222
rect 2791 2226 2795 2227
rect 2791 2221 2795 2222
rect 2903 2226 2907 2227
rect 2903 2221 2907 2222
rect 2927 2226 2931 2227
rect 2927 2221 2931 2222
rect 3047 2226 3051 2227
rect 3047 2221 3051 2222
rect 3103 2226 3107 2227
rect 3103 2221 3107 2222
rect 3167 2226 3171 2227
rect 3167 2221 3171 2222
rect 3279 2226 3283 2227
rect 3279 2221 3283 2222
rect 3303 2226 3307 2227
rect 3303 2221 3307 2222
rect 3391 2226 3395 2227
rect 3391 2221 3395 2222
rect 3487 2226 3491 2227
rect 3487 2221 3491 2222
rect 3575 2226 3579 2227
rect 3575 2221 3579 2222
rect 112 2206 114 2221
rect 536 2216 538 2221
rect 720 2216 722 2221
rect 896 2216 898 2221
rect 1072 2216 1074 2221
rect 1240 2216 1242 2221
rect 1408 2216 1410 2221
rect 1576 2216 1578 2221
rect 1728 2216 1730 2221
rect 534 2215 540 2216
rect 534 2211 535 2215
rect 539 2211 540 2215
rect 534 2210 540 2211
rect 718 2215 724 2216
rect 718 2211 719 2215
rect 723 2211 724 2215
rect 718 2210 724 2211
rect 894 2215 900 2216
rect 894 2211 895 2215
rect 899 2211 900 2215
rect 894 2210 900 2211
rect 1070 2215 1076 2216
rect 1070 2211 1071 2215
rect 1075 2211 1076 2215
rect 1070 2210 1076 2211
rect 1238 2215 1244 2216
rect 1238 2211 1239 2215
rect 1243 2211 1244 2215
rect 1238 2210 1244 2211
rect 1406 2215 1412 2216
rect 1406 2211 1407 2215
rect 1411 2211 1412 2215
rect 1406 2210 1412 2211
rect 1574 2215 1580 2216
rect 1574 2211 1575 2215
rect 1579 2211 1580 2215
rect 1574 2210 1580 2211
rect 1726 2215 1732 2216
rect 1726 2211 1727 2215
rect 1731 2211 1732 2215
rect 1726 2210 1732 2211
rect 1824 2206 1826 2221
rect 110 2205 116 2206
rect 110 2201 111 2205
rect 115 2201 116 2205
rect 110 2200 116 2201
rect 1822 2205 1828 2206
rect 1822 2201 1823 2205
rect 1827 2201 1828 2205
rect 1822 2200 1828 2201
rect 1864 2197 1866 2221
rect 2008 2210 2010 2221
rect 2168 2210 2170 2221
rect 2336 2210 2338 2221
rect 2520 2210 2522 2221
rect 2712 2210 2714 2221
rect 2904 2210 2906 2221
rect 3104 2210 3106 2221
rect 3304 2210 3306 2221
rect 3488 2210 3490 2221
rect 2006 2209 2012 2210
rect 2006 2205 2007 2209
rect 2011 2205 2012 2209
rect 2006 2204 2012 2205
rect 2166 2209 2172 2210
rect 2166 2205 2167 2209
rect 2171 2205 2172 2209
rect 2166 2204 2172 2205
rect 2334 2209 2340 2210
rect 2334 2205 2335 2209
rect 2339 2205 2340 2209
rect 2334 2204 2340 2205
rect 2518 2209 2524 2210
rect 2518 2205 2519 2209
rect 2523 2205 2524 2209
rect 2518 2204 2524 2205
rect 2710 2209 2716 2210
rect 2710 2205 2711 2209
rect 2715 2205 2716 2209
rect 2710 2204 2716 2205
rect 2902 2209 2908 2210
rect 2902 2205 2903 2209
rect 2907 2205 2908 2209
rect 2902 2204 2908 2205
rect 3102 2209 3108 2210
rect 3102 2205 3103 2209
rect 3107 2205 3108 2209
rect 3102 2204 3108 2205
rect 3302 2209 3308 2210
rect 3302 2205 3303 2209
rect 3307 2205 3308 2209
rect 3302 2204 3308 2205
rect 3486 2209 3492 2210
rect 3486 2205 3487 2209
rect 3491 2205 3492 2209
rect 3486 2204 3492 2205
rect 3576 2197 3578 2221
rect 1862 2196 1868 2197
rect 1862 2192 1863 2196
rect 1867 2192 1868 2196
rect 1862 2191 1868 2192
rect 3574 2196 3580 2197
rect 3574 2192 3575 2196
rect 3579 2192 3580 2196
rect 3574 2191 3580 2192
rect 110 2188 116 2189
rect 110 2184 111 2188
rect 115 2184 116 2188
rect 110 2183 116 2184
rect 1822 2188 1828 2189
rect 1822 2184 1823 2188
rect 1827 2184 1828 2188
rect 1822 2183 1828 2184
rect 112 2159 114 2183
rect 542 2175 548 2176
rect 542 2171 543 2175
rect 547 2171 548 2175
rect 542 2170 548 2171
rect 726 2175 732 2176
rect 726 2171 727 2175
rect 731 2171 732 2175
rect 726 2170 732 2171
rect 902 2175 908 2176
rect 902 2171 903 2175
rect 907 2171 908 2175
rect 902 2170 908 2171
rect 1078 2175 1084 2176
rect 1078 2171 1079 2175
rect 1083 2171 1084 2175
rect 1078 2170 1084 2171
rect 1246 2175 1252 2176
rect 1246 2171 1247 2175
rect 1251 2171 1252 2175
rect 1246 2170 1252 2171
rect 1414 2175 1420 2176
rect 1414 2171 1415 2175
rect 1419 2171 1420 2175
rect 1414 2170 1420 2171
rect 1582 2175 1588 2176
rect 1582 2171 1583 2175
rect 1587 2171 1588 2175
rect 1582 2170 1588 2171
rect 1734 2175 1740 2176
rect 1734 2171 1735 2175
rect 1739 2171 1740 2175
rect 1734 2170 1740 2171
rect 544 2159 546 2170
rect 728 2159 730 2170
rect 904 2159 906 2170
rect 1080 2159 1082 2170
rect 1248 2159 1250 2170
rect 1416 2159 1418 2170
rect 1584 2159 1586 2170
rect 1736 2159 1738 2170
rect 1824 2159 1826 2183
rect 1862 2179 1868 2180
rect 1862 2175 1863 2179
rect 1867 2175 1868 2179
rect 1862 2174 1868 2175
rect 3574 2179 3580 2180
rect 3574 2175 3575 2179
rect 3579 2175 3580 2179
rect 3574 2174 3580 2175
rect 111 2158 115 2159
rect 111 2153 115 2154
rect 495 2158 499 2159
rect 495 2153 499 2154
rect 543 2158 547 2159
rect 543 2153 547 2154
rect 623 2158 627 2159
rect 623 2153 627 2154
rect 727 2158 731 2159
rect 727 2153 731 2154
rect 759 2158 763 2159
rect 759 2153 763 2154
rect 895 2158 899 2159
rect 895 2153 899 2154
rect 903 2158 907 2159
rect 903 2153 907 2154
rect 1039 2158 1043 2159
rect 1039 2153 1043 2154
rect 1079 2158 1083 2159
rect 1079 2153 1083 2154
rect 1183 2158 1187 2159
rect 1183 2153 1187 2154
rect 1247 2158 1251 2159
rect 1247 2153 1251 2154
rect 1327 2158 1331 2159
rect 1327 2153 1331 2154
rect 1415 2158 1419 2159
rect 1415 2153 1419 2154
rect 1471 2158 1475 2159
rect 1471 2153 1475 2154
rect 1583 2158 1587 2159
rect 1583 2153 1587 2154
rect 1623 2158 1627 2159
rect 1623 2153 1627 2154
rect 1735 2158 1739 2159
rect 1735 2153 1739 2154
rect 1823 2158 1827 2159
rect 1823 2153 1827 2154
rect 112 2129 114 2153
rect 496 2142 498 2153
rect 624 2142 626 2153
rect 760 2142 762 2153
rect 896 2142 898 2153
rect 1040 2142 1042 2153
rect 1184 2142 1186 2153
rect 1328 2142 1330 2153
rect 1472 2142 1474 2153
rect 1624 2142 1626 2153
rect 494 2141 500 2142
rect 494 2137 495 2141
rect 499 2137 500 2141
rect 494 2136 500 2137
rect 622 2141 628 2142
rect 622 2137 623 2141
rect 627 2137 628 2141
rect 622 2136 628 2137
rect 758 2141 764 2142
rect 758 2137 759 2141
rect 763 2137 764 2141
rect 758 2136 764 2137
rect 894 2141 900 2142
rect 894 2137 895 2141
rect 899 2137 900 2141
rect 894 2136 900 2137
rect 1038 2141 1044 2142
rect 1038 2137 1039 2141
rect 1043 2137 1044 2141
rect 1038 2136 1044 2137
rect 1182 2141 1188 2142
rect 1182 2137 1183 2141
rect 1187 2137 1188 2141
rect 1182 2136 1188 2137
rect 1326 2141 1332 2142
rect 1326 2137 1327 2141
rect 1331 2137 1332 2141
rect 1326 2136 1332 2137
rect 1470 2141 1476 2142
rect 1470 2137 1471 2141
rect 1475 2137 1476 2141
rect 1470 2136 1476 2137
rect 1622 2141 1628 2142
rect 1622 2137 1623 2141
rect 1627 2137 1628 2141
rect 1622 2136 1628 2137
rect 1824 2129 1826 2153
rect 1864 2151 1866 2174
rect 1998 2169 2004 2170
rect 1998 2165 1999 2169
rect 2003 2165 2004 2169
rect 1998 2164 2004 2165
rect 2158 2169 2164 2170
rect 2158 2165 2159 2169
rect 2163 2165 2164 2169
rect 2158 2164 2164 2165
rect 2326 2169 2332 2170
rect 2326 2165 2327 2169
rect 2331 2165 2332 2169
rect 2326 2164 2332 2165
rect 2510 2169 2516 2170
rect 2510 2165 2511 2169
rect 2515 2165 2516 2169
rect 2510 2164 2516 2165
rect 2702 2169 2708 2170
rect 2702 2165 2703 2169
rect 2707 2165 2708 2169
rect 2702 2164 2708 2165
rect 2894 2169 2900 2170
rect 2894 2165 2895 2169
rect 2899 2165 2900 2169
rect 2894 2164 2900 2165
rect 3094 2169 3100 2170
rect 3094 2165 3095 2169
rect 3099 2165 3100 2169
rect 3094 2164 3100 2165
rect 3294 2169 3300 2170
rect 3294 2165 3295 2169
rect 3299 2165 3300 2169
rect 3294 2164 3300 2165
rect 3478 2169 3484 2170
rect 3478 2165 3479 2169
rect 3483 2165 3484 2169
rect 3478 2164 3484 2165
rect 2000 2151 2002 2164
rect 2160 2151 2162 2164
rect 2328 2151 2330 2164
rect 2512 2151 2514 2164
rect 2704 2151 2706 2164
rect 2896 2151 2898 2164
rect 3096 2151 3098 2164
rect 3296 2151 3298 2164
rect 3480 2151 3482 2164
rect 3576 2151 3578 2174
rect 1863 2150 1867 2151
rect 1863 2145 1867 2146
rect 1999 2150 2003 2151
rect 1999 2145 2003 2146
rect 2023 2150 2027 2151
rect 2023 2145 2027 2146
rect 2159 2150 2163 2151
rect 2159 2145 2163 2146
rect 2167 2150 2171 2151
rect 2167 2145 2171 2146
rect 2319 2150 2323 2151
rect 2319 2145 2323 2146
rect 2327 2150 2331 2151
rect 2327 2145 2331 2146
rect 2471 2150 2475 2151
rect 2471 2145 2475 2146
rect 2511 2150 2515 2151
rect 2511 2145 2515 2146
rect 2615 2150 2619 2151
rect 2615 2145 2619 2146
rect 2703 2150 2707 2151
rect 2703 2145 2707 2146
rect 2759 2150 2763 2151
rect 2759 2145 2763 2146
rect 2895 2150 2899 2151
rect 2895 2145 2899 2146
rect 3023 2150 3027 2151
rect 3023 2145 3027 2146
rect 3095 2150 3099 2151
rect 3095 2145 3099 2146
rect 3143 2150 3147 2151
rect 3143 2145 3147 2146
rect 3263 2150 3267 2151
rect 3263 2145 3267 2146
rect 3295 2150 3299 2151
rect 3295 2145 3299 2146
rect 3383 2150 3387 2151
rect 3383 2145 3387 2146
rect 3479 2150 3483 2151
rect 3479 2145 3483 2146
rect 3575 2150 3579 2151
rect 3575 2145 3579 2146
rect 1864 2130 1866 2145
rect 2024 2140 2026 2145
rect 2168 2140 2170 2145
rect 2320 2140 2322 2145
rect 2472 2140 2474 2145
rect 2616 2140 2618 2145
rect 2760 2140 2762 2145
rect 2896 2140 2898 2145
rect 3024 2140 3026 2145
rect 3144 2140 3146 2145
rect 3264 2140 3266 2145
rect 3384 2140 3386 2145
rect 3480 2140 3482 2145
rect 2022 2139 2028 2140
rect 2022 2135 2023 2139
rect 2027 2135 2028 2139
rect 2022 2134 2028 2135
rect 2166 2139 2172 2140
rect 2166 2135 2167 2139
rect 2171 2135 2172 2139
rect 2166 2134 2172 2135
rect 2318 2139 2324 2140
rect 2318 2135 2319 2139
rect 2323 2135 2324 2139
rect 2318 2134 2324 2135
rect 2470 2139 2476 2140
rect 2470 2135 2471 2139
rect 2475 2135 2476 2139
rect 2470 2134 2476 2135
rect 2614 2139 2620 2140
rect 2614 2135 2615 2139
rect 2619 2135 2620 2139
rect 2614 2134 2620 2135
rect 2758 2139 2764 2140
rect 2758 2135 2759 2139
rect 2763 2135 2764 2139
rect 2758 2134 2764 2135
rect 2894 2139 2900 2140
rect 2894 2135 2895 2139
rect 2899 2135 2900 2139
rect 2894 2134 2900 2135
rect 3022 2139 3028 2140
rect 3022 2135 3023 2139
rect 3027 2135 3028 2139
rect 3022 2134 3028 2135
rect 3142 2139 3148 2140
rect 3142 2135 3143 2139
rect 3147 2135 3148 2139
rect 3142 2134 3148 2135
rect 3262 2139 3268 2140
rect 3262 2135 3263 2139
rect 3267 2135 3268 2139
rect 3262 2134 3268 2135
rect 3382 2139 3388 2140
rect 3382 2135 3383 2139
rect 3387 2135 3388 2139
rect 3382 2134 3388 2135
rect 3478 2139 3484 2140
rect 3478 2135 3479 2139
rect 3483 2135 3484 2139
rect 3478 2134 3484 2135
rect 3576 2130 3578 2145
rect 1862 2129 1868 2130
rect 110 2128 116 2129
rect 110 2124 111 2128
rect 115 2124 116 2128
rect 110 2123 116 2124
rect 1822 2128 1828 2129
rect 1822 2124 1823 2128
rect 1827 2124 1828 2128
rect 1862 2125 1863 2129
rect 1867 2125 1868 2129
rect 1862 2124 1868 2125
rect 3574 2129 3580 2130
rect 3574 2125 3575 2129
rect 3579 2125 3580 2129
rect 3574 2124 3580 2125
rect 1822 2123 1828 2124
rect 1862 2112 1868 2113
rect 110 2111 116 2112
rect 110 2107 111 2111
rect 115 2107 116 2111
rect 110 2106 116 2107
rect 1822 2111 1828 2112
rect 1822 2107 1823 2111
rect 1827 2107 1828 2111
rect 1862 2108 1863 2112
rect 1867 2108 1868 2112
rect 1862 2107 1868 2108
rect 3574 2112 3580 2113
rect 3574 2108 3575 2112
rect 3579 2108 3580 2112
rect 3574 2107 3580 2108
rect 1822 2106 1828 2107
rect 112 2087 114 2106
rect 486 2101 492 2102
rect 486 2097 487 2101
rect 491 2097 492 2101
rect 486 2096 492 2097
rect 614 2101 620 2102
rect 614 2097 615 2101
rect 619 2097 620 2101
rect 614 2096 620 2097
rect 750 2101 756 2102
rect 750 2097 751 2101
rect 755 2097 756 2101
rect 750 2096 756 2097
rect 886 2101 892 2102
rect 886 2097 887 2101
rect 891 2097 892 2101
rect 886 2096 892 2097
rect 1030 2101 1036 2102
rect 1030 2097 1031 2101
rect 1035 2097 1036 2101
rect 1030 2096 1036 2097
rect 1174 2101 1180 2102
rect 1174 2097 1175 2101
rect 1179 2097 1180 2101
rect 1174 2096 1180 2097
rect 1318 2101 1324 2102
rect 1318 2097 1319 2101
rect 1323 2097 1324 2101
rect 1318 2096 1324 2097
rect 1462 2101 1468 2102
rect 1462 2097 1463 2101
rect 1467 2097 1468 2101
rect 1462 2096 1468 2097
rect 1614 2101 1620 2102
rect 1614 2097 1615 2101
rect 1619 2097 1620 2101
rect 1614 2096 1620 2097
rect 488 2087 490 2096
rect 616 2087 618 2096
rect 752 2087 754 2096
rect 888 2087 890 2096
rect 1032 2087 1034 2096
rect 1176 2087 1178 2096
rect 1320 2087 1322 2096
rect 1464 2087 1466 2096
rect 1616 2087 1618 2096
rect 1824 2087 1826 2106
rect 111 2086 115 2087
rect 111 2081 115 2082
rect 319 2086 323 2087
rect 319 2081 323 2082
rect 431 2086 435 2087
rect 431 2081 435 2082
rect 487 2086 491 2087
rect 487 2081 491 2082
rect 551 2086 555 2087
rect 551 2081 555 2082
rect 615 2086 619 2087
rect 615 2081 619 2082
rect 679 2086 683 2087
rect 679 2081 683 2082
rect 751 2086 755 2087
rect 751 2081 755 2082
rect 799 2086 803 2087
rect 799 2081 803 2082
rect 887 2086 891 2087
rect 887 2081 891 2082
rect 919 2086 923 2087
rect 919 2081 923 2082
rect 1031 2086 1035 2087
rect 1031 2081 1035 2082
rect 1039 2086 1043 2087
rect 1039 2081 1043 2082
rect 1159 2086 1163 2087
rect 1159 2081 1163 2082
rect 1175 2086 1179 2087
rect 1175 2081 1179 2082
rect 1279 2086 1283 2087
rect 1279 2081 1283 2082
rect 1319 2086 1323 2087
rect 1319 2081 1323 2082
rect 1407 2086 1411 2087
rect 1407 2081 1411 2082
rect 1463 2086 1467 2087
rect 1463 2081 1467 2082
rect 1615 2086 1619 2087
rect 1615 2081 1619 2082
rect 1823 2086 1827 2087
rect 1823 2081 1827 2082
rect 112 2066 114 2081
rect 320 2076 322 2081
rect 432 2076 434 2081
rect 552 2076 554 2081
rect 680 2076 682 2081
rect 800 2076 802 2081
rect 920 2076 922 2081
rect 1040 2076 1042 2081
rect 1160 2076 1162 2081
rect 1280 2076 1282 2081
rect 1408 2076 1410 2081
rect 318 2075 324 2076
rect 318 2071 319 2075
rect 323 2071 324 2075
rect 318 2070 324 2071
rect 430 2075 436 2076
rect 430 2071 431 2075
rect 435 2071 436 2075
rect 430 2070 436 2071
rect 550 2075 556 2076
rect 550 2071 551 2075
rect 555 2071 556 2075
rect 550 2070 556 2071
rect 678 2075 684 2076
rect 678 2071 679 2075
rect 683 2071 684 2075
rect 678 2070 684 2071
rect 798 2075 804 2076
rect 798 2071 799 2075
rect 803 2071 804 2075
rect 798 2070 804 2071
rect 918 2075 924 2076
rect 918 2071 919 2075
rect 923 2071 924 2075
rect 918 2070 924 2071
rect 1038 2075 1044 2076
rect 1038 2071 1039 2075
rect 1043 2071 1044 2075
rect 1038 2070 1044 2071
rect 1158 2075 1164 2076
rect 1158 2071 1159 2075
rect 1163 2071 1164 2075
rect 1158 2070 1164 2071
rect 1278 2075 1284 2076
rect 1278 2071 1279 2075
rect 1283 2071 1284 2075
rect 1278 2070 1284 2071
rect 1406 2075 1412 2076
rect 1406 2071 1407 2075
rect 1411 2071 1412 2075
rect 1406 2070 1412 2071
rect 1824 2066 1826 2081
rect 1864 2079 1866 2107
rect 2030 2099 2036 2100
rect 2030 2095 2031 2099
rect 2035 2095 2036 2099
rect 2030 2094 2036 2095
rect 2174 2099 2180 2100
rect 2174 2095 2175 2099
rect 2179 2095 2180 2099
rect 2174 2094 2180 2095
rect 2326 2099 2332 2100
rect 2326 2095 2327 2099
rect 2331 2095 2332 2099
rect 2326 2094 2332 2095
rect 2478 2099 2484 2100
rect 2478 2095 2479 2099
rect 2483 2095 2484 2099
rect 2478 2094 2484 2095
rect 2622 2099 2628 2100
rect 2622 2095 2623 2099
rect 2627 2095 2628 2099
rect 2622 2094 2628 2095
rect 2766 2099 2772 2100
rect 2766 2095 2767 2099
rect 2771 2095 2772 2099
rect 2766 2094 2772 2095
rect 2902 2099 2908 2100
rect 2902 2095 2903 2099
rect 2907 2095 2908 2099
rect 2902 2094 2908 2095
rect 3030 2099 3036 2100
rect 3030 2095 3031 2099
rect 3035 2095 3036 2099
rect 3030 2094 3036 2095
rect 3150 2099 3156 2100
rect 3150 2095 3151 2099
rect 3155 2095 3156 2099
rect 3150 2094 3156 2095
rect 3270 2099 3276 2100
rect 3270 2095 3271 2099
rect 3275 2095 3276 2099
rect 3270 2094 3276 2095
rect 3390 2099 3396 2100
rect 3390 2095 3391 2099
rect 3395 2095 3396 2099
rect 3390 2094 3396 2095
rect 3486 2099 3492 2100
rect 3486 2095 3487 2099
rect 3491 2095 3492 2099
rect 3486 2094 3492 2095
rect 2032 2079 2034 2094
rect 2176 2079 2178 2094
rect 2328 2079 2330 2094
rect 2480 2079 2482 2094
rect 2624 2079 2626 2094
rect 2768 2079 2770 2094
rect 2904 2079 2906 2094
rect 3032 2079 3034 2094
rect 3152 2079 3154 2094
rect 3272 2079 3274 2094
rect 3392 2079 3394 2094
rect 3488 2079 3490 2094
rect 3576 2079 3578 2107
rect 1863 2078 1867 2079
rect 1863 2073 1867 2074
rect 1983 2078 1987 2079
rect 1983 2073 1987 2074
rect 2031 2078 2035 2079
rect 2031 2073 2035 2074
rect 2143 2078 2147 2079
rect 2143 2073 2147 2074
rect 2175 2078 2179 2079
rect 2175 2073 2179 2074
rect 2311 2078 2315 2079
rect 2311 2073 2315 2074
rect 2327 2078 2331 2079
rect 2327 2073 2331 2074
rect 2471 2078 2475 2079
rect 2471 2073 2475 2074
rect 2479 2078 2483 2079
rect 2479 2073 2483 2074
rect 2623 2078 2627 2079
rect 2623 2073 2627 2074
rect 2631 2078 2635 2079
rect 2631 2073 2635 2074
rect 2767 2078 2771 2079
rect 2767 2073 2771 2074
rect 2775 2078 2779 2079
rect 2775 2073 2779 2074
rect 2903 2078 2907 2079
rect 2903 2073 2907 2074
rect 2911 2078 2915 2079
rect 2911 2073 2915 2074
rect 3031 2078 3035 2079
rect 3031 2073 3035 2074
rect 3039 2078 3043 2079
rect 3039 2073 3043 2074
rect 3151 2078 3155 2079
rect 3151 2073 3155 2074
rect 3159 2078 3163 2079
rect 3159 2073 3163 2074
rect 3271 2078 3275 2079
rect 3271 2073 3275 2074
rect 3279 2078 3283 2079
rect 3279 2073 3283 2074
rect 3391 2078 3395 2079
rect 3391 2073 3395 2074
rect 3487 2078 3491 2079
rect 3487 2073 3491 2074
rect 3575 2078 3579 2079
rect 3575 2073 3579 2074
rect 110 2065 116 2066
rect 110 2061 111 2065
rect 115 2061 116 2065
rect 110 2060 116 2061
rect 1822 2065 1828 2066
rect 1822 2061 1823 2065
rect 1827 2061 1828 2065
rect 1822 2060 1828 2061
rect 1864 2049 1866 2073
rect 1984 2062 1986 2073
rect 2144 2062 2146 2073
rect 2312 2062 2314 2073
rect 2472 2062 2474 2073
rect 2632 2062 2634 2073
rect 2776 2062 2778 2073
rect 2912 2062 2914 2073
rect 3040 2062 3042 2073
rect 3160 2062 3162 2073
rect 3280 2062 3282 2073
rect 3392 2062 3394 2073
rect 3488 2062 3490 2073
rect 1982 2061 1988 2062
rect 1982 2057 1983 2061
rect 1987 2057 1988 2061
rect 1982 2056 1988 2057
rect 2142 2061 2148 2062
rect 2142 2057 2143 2061
rect 2147 2057 2148 2061
rect 2142 2056 2148 2057
rect 2310 2061 2316 2062
rect 2310 2057 2311 2061
rect 2315 2057 2316 2061
rect 2310 2056 2316 2057
rect 2470 2061 2476 2062
rect 2470 2057 2471 2061
rect 2475 2057 2476 2061
rect 2470 2056 2476 2057
rect 2630 2061 2636 2062
rect 2630 2057 2631 2061
rect 2635 2057 2636 2061
rect 2630 2056 2636 2057
rect 2774 2061 2780 2062
rect 2774 2057 2775 2061
rect 2779 2057 2780 2061
rect 2774 2056 2780 2057
rect 2910 2061 2916 2062
rect 2910 2057 2911 2061
rect 2915 2057 2916 2061
rect 2910 2056 2916 2057
rect 3038 2061 3044 2062
rect 3038 2057 3039 2061
rect 3043 2057 3044 2061
rect 3038 2056 3044 2057
rect 3158 2061 3164 2062
rect 3158 2057 3159 2061
rect 3163 2057 3164 2061
rect 3158 2056 3164 2057
rect 3278 2061 3284 2062
rect 3278 2057 3279 2061
rect 3283 2057 3284 2061
rect 3278 2056 3284 2057
rect 3390 2061 3396 2062
rect 3390 2057 3391 2061
rect 3395 2057 3396 2061
rect 3390 2056 3396 2057
rect 3486 2061 3492 2062
rect 3486 2057 3487 2061
rect 3491 2057 3492 2061
rect 3486 2056 3492 2057
rect 3576 2049 3578 2073
rect 110 2048 116 2049
rect 110 2044 111 2048
rect 115 2044 116 2048
rect 110 2043 116 2044
rect 1822 2048 1828 2049
rect 1822 2044 1823 2048
rect 1827 2044 1828 2048
rect 1822 2043 1828 2044
rect 1862 2048 1868 2049
rect 1862 2044 1863 2048
rect 1867 2044 1868 2048
rect 1862 2043 1868 2044
rect 3574 2048 3580 2049
rect 3574 2044 3575 2048
rect 3579 2044 3580 2048
rect 3574 2043 3580 2044
rect 112 2015 114 2043
rect 326 2035 332 2036
rect 326 2031 327 2035
rect 331 2031 332 2035
rect 326 2030 332 2031
rect 438 2035 444 2036
rect 438 2031 439 2035
rect 443 2031 444 2035
rect 438 2030 444 2031
rect 558 2035 564 2036
rect 558 2031 559 2035
rect 563 2031 564 2035
rect 558 2030 564 2031
rect 686 2035 692 2036
rect 686 2031 687 2035
rect 691 2031 692 2035
rect 686 2030 692 2031
rect 806 2035 812 2036
rect 806 2031 807 2035
rect 811 2031 812 2035
rect 806 2030 812 2031
rect 926 2035 932 2036
rect 926 2031 927 2035
rect 931 2031 932 2035
rect 926 2030 932 2031
rect 1046 2035 1052 2036
rect 1046 2031 1047 2035
rect 1051 2031 1052 2035
rect 1046 2030 1052 2031
rect 1166 2035 1172 2036
rect 1166 2031 1167 2035
rect 1171 2031 1172 2035
rect 1166 2030 1172 2031
rect 1286 2035 1292 2036
rect 1286 2031 1287 2035
rect 1291 2031 1292 2035
rect 1286 2030 1292 2031
rect 1414 2035 1420 2036
rect 1414 2031 1415 2035
rect 1419 2031 1420 2035
rect 1414 2030 1420 2031
rect 328 2015 330 2030
rect 440 2015 442 2030
rect 560 2015 562 2030
rect 688 2015 690 2030
rect 808 2015 810 2030
rect 928 2015 930 2030
rect 1048 2015 1050 2030
rect 1168 2015 1170 2030
rect 1288 2015 1290 2030
rect 1416 2015 1418 2030
rect 1824 2015 1826 2043
rect 1862 2031 1868 2032
rect 1862 2027 1863 2031
rect 1867 2027 1868 2031
rect 1862 2026 1868 2027
rect 3574 2031 3580 2032
rect 3574 2027 3575 2031
rect 3579 2027 3580 2031
rect 3574 2026 3580 2027
rect 111 2014 115 2015
rect 111 2009 115 2010
rect 183 2014 187 2015
rect 183 2009 187 2010
rect 295 2014 299 2015
rect 295 2009 299 2010
rect 327 2014 331 2015
rect 327 2009 331 2010
rect 415 2014 419 2015
rect 415 2009 419 2010
rect 439 2014 443 2015
rect 439 2009 443 2010
rect 535 2014 539 2015
rect 535 2009 539 2010
rect 559 2014 563 2015
rect 559 2009 563 2010
rect 655 2014 659 2015
rect 655 2009 659 2010
rect 687 2014 691 2015
rect 687 2009 691 2010
rect 775 2014 779 2015
rect 775 2009 779 2010
rect 807 2014 811 2015
rect 807 2009 811 2010
rect 895 2014 899 2015
rect 895 2009 899 2010
rect 927 2014 931 2015
rect 927 2009 931 2010
rect 1015 2014 1019 2015
rect 1015 2009 1019 2010
rect 1047 2014 1051 2015
rect 1047 2009 1051 2010
rect 1135 2014 1139 2015
rect 1135 2009 1139 2010
rect 1167 2014 1171 2015
rect 1167 2009 1171 2010
rect 1255 2014 1259 2015
rect 1255 2009 1259 2010
rect 1287 2014 1291 2015
rect 1287 2009 1291 2010
rect 1415 2014 1419 2015
rect 1415 2009 1419 2010
rect 1823 2014 1827 2015
rect 1864 2011 1866 2026
rect 1974 2021 1980 2022
rect 1974 2017 1975 2021
rect 1979 2017 1980 2021
rect 1974 2016 1980 2017
rect 2134 2021 2140 2022
rect 2134 2017 2135 2021
rect 2139 2017 2140 2021
rect 2134 2016 2140 2017
rect 2302 2021 2308 2022
rect 2302 2017 2303 2021
rect 2307 2017 2308 2021
rect 2302 2016 2308 2017
rect 2462 2021 2468 2022
rect 2462 2017 2463 2021
rect 2467 2017 2468 2021
rect 2462 2016 2468 2017
rect 2622 2021 2628 2022
rect 2622 2017 2623 2021
rect 2627 2017 2628 2021
rect 2622 2016 2628 2017
rect 2766 2021 2772 2022
rect 2766 2017 2767 2021
rect 2771 2017 2772 2021
rect 2766 2016 2772 2017
rect 2902 2021 2908 2022
rect 2902 2017 2903 2021
rect 2907 2017 2908 2021
rect 2902 2016 2908 2017
rect 3030 2021 3036 2022
rect 3030 2017 3031 2021
rect 3035 2017 3036 2021
rect 3030 2016 3036 2017
rect 3150 2021 3156 2022
rect 3150 2017 3151 2021
rect 3155 2017 3156 2021
rect 3150 2016 3156 2017
rect 3270 2021 3276 2022
rect 3270 2017 3271 2021
rect 3275 2017 3276 2021
rect 3270 2016 3276 2017
rect 3382 2021 3388 2022
rect 3382 2017 3383 2021
rect 3387 2017 3388 2021
rect 3382 2016 3388 2017
rect 3478 2021 3484 2022
rect 3478 2017 3479 2021
rect 3483 2017 3484 2021
rect 3478 2016 3484 2017
rect 1976 2011 1978 2016
rect 2136 2011 2138 2016
rect 2304 2011 2306 2016
rect 2464 2011 2466 2016
rect 2624 2011 2626 2016
rect 2768 2011 2770 2016
rect 2904 2011 2906 2016
rect 3032 2011 3034 2016
rect 3152 2011 3154 2016
rect 3272 2011 3274 2016
rect 3384 2011 3386 2016
rect 3480 2011 3482 2016
rect 3576 2011 3578 2026
rect 1823 2009 1827 2010
rect 1863 2010 1867 2011
rect 112 1985 114 2009
rect 184 1998 186 2009
rect 296 1998 298 2009
rect 416 1998 418 2009
rect 536 1998 538 2009
rect 656 1998 658 2009
rect 776 1998 778 2009
rect 896 1998 898 2009
rect 1016 1998 1018 2009
rect 1136 1998 1138 2009
rect 1256 1998 1258 2009
rect 182 1997 188 1998
rect 182 1993 183 1997
rect 187 1993 188 1997
rect 182 1992 188 1993
rect 294 1997 300 1998
rect 294 1993 295 1997
rect 299 1993 300 1997
rect 294 1992 300 1993
rect 414 1997 420 1998
rect 414 1993 415 1997
rect 419 1993 420 1997
rect 414 1992 420 1993
rect 534 1997 540 1998
rect 534 1993 535 1997
rect 539 1993 540 1997
rect 534 1992 540 1993
rect 654 1997 660 1998
rect 654 1993 655 1997
rect 659 1993 660 1997
rect 654 1992 660 1993
rect 774 1997 780 1998
rect 774 1993 775 1997
rect 779 1993 780 1997
rect 774 1992 780 1993
rect 894 1997 900 1998
rect 894 1993 895 1997
rect 899 1993 900 1997
rect 894 1992 900 1993
rect 1014 1997 1020 1998
rect 1014 1993 1015 1997
rect 1019 1993 1020 1997
rect 1014 1992 1020 1993
rect 1134 1997 1140 1998
rect 1134 1993 1135 1997
rect 1139 1993 1140 1997
rect 1134 1992 1140 1993
rect 1254 1997 1260 1998
rect 1254 1993 1255 1997
rect 1259 1993 1260 1997
rect 1254 1992 1260 1993
rect 1824 1985 1826 2009
rect 1863 2005 1867 2006
rect 1887 2010 1891 2011
rect 1887 2005 1891 2006
rect 1975 2010 1979 2011
rect 1975 2005 1979 2006
rect 2031 2010 2035 2011
rect 2031 2005 2035 2006
rect 2135 2010 2139 2011
rect 2135 2005 2139 2006
rect 2199 2010 2203 2011
rect 2199 2005 2203 2006
rect 2303 2010 2307 2011
rect 2303 2005 2307 2006
rect 2375 2010 2379 2011
rect 2375 2005 2379 2006
rect 2463 2010 2467 2011
rect 2463 2005 2467 2006
rect 2543 2010 2547 2011
rect 2543 2005 2547 2006
rect 2623 2010 2627 2011
rect 2623 2005 2627 2006
rect 2711 2010 2715 2011
rect 2711 2005 2715 2006
rect 2767 2010 2771 2011
rect 2767 2005 2771 2006
rect 2871 2010 2875 2011
rect 2871 2005 2875 2006
rect 2903 2010 2907 2011
rect 2903 2005 2907 2006
rect 3031 2010 3035 2011
rect 3031 2005 3035 2006
rect 3039 2010 3043 2011
rect 3039 2005 3043 2006
rect 3151 2010 3155 2011
rect 3151 2005 3155 2006
rect 3207 2010 3211 2011
rect 3207 2005 3211 2006
rect 3271 2010 3275 2011
rect 3271 2005 3275 2006
rect 3383 2010 3387 2011
rect 3383 2005 3387 2006
rect 3479 2010 3483 2011
rect 3479 2005 3483 2006
rect 3575 2010 3579 2011
rect 3575 2005 3579 2006
rect 1864 1990 1866 2005
rect 1888 2000 1890 2005
rect 2032 2000 2034 2005
rect 2200 2000 2202 2005
rect 2376 2000 2378 2005
rect 2544 2000 2546 2005
rect 2712 2000 2714 2005
rect 2872 2000 2874 2005
rect 3040 2000 3042 2005
rect 3208 2000 3210 2005
rect 1886 1999 1892 2000
rect 1886 1995 1887 1999
rect 1891 1995 1892 1999
rect 1886 1994 1892 1995
rect 2030 1999 2036 2000
rect 2030 1995 2031 1999
rect 2035 1995 2036 1999
rect 2030 1994 2036 1995
rect 2198 1999 2204 2000
rect 2198 1995 2199 1999
rect 2203 1995 2204 1999
rect 2198 1994 2204 1995
rect 2374 1999 2380 2000
rect 2374 1995 2375 1999
rect 2379 1995 2380 1999
rect 2374 1994 2380 1995
rect 2542 1999 2548 2000
rect 2542 1995 2543 1999
rect 2547 1995 2548 1999
rect 2542 1994 2548 1995
rect 2710 1999 2716 2000
rect 2710 1995 2711 1999
rect 2715 1995 2716 1999
rect 2710 1994 2716 1995
rect 2870 1999 2876 2000
rect 2870 1995 2871 1999
rect 2875 1995 2876 1999
rect 2870 1994 2876 1995
rect 3038 1999 3044 2000
rect 3038 1995 3039 1999
rect 3043 1995 3044 1999
rect 3038 1994 3044 1995
rect 3206 1999 3212 2000
rect 3206 1995 3207 1999
rect 3211 1995 3212 1999
rect 3206 1994 3212 1995
rect 3576 1990 3578 2005
rect 1862 1989 1868 1990
rect 1862 1985 1863 1989
rect 1867 1985 1868 1989
rect 110 1984 116 1985
rect 110 1980 111 1984
rect 115 1980 116 1984
rect 110 1979 116 1980
rect 1822 1984 1828 1985
rect 1862 1984 1868 1985
rect 3574 1989 3580 1990
rect 3574 1985 3575 1989
rect 3579 1985 3580 1989
rect 3574 1984 3580 1985
rect 1822 1980 1823 1984
rect 1827 1980 1828 1984
rect 1822 1979 1828 1980
rect 1862 1972 1868 1973
rect 1862 1968 1863 1972
rect 1867 1968 1868 1972
rect 110 1967 116 1968
rect 110 1963 111 1967
rect 115 1963 116 1967
rect 110 1962 116 1963
rect 1822 1967 1828 1968
rect 1862 1967 1868 1968
rect 3574 1972 3580 1973
rect 3574 1968 3575 1972
rect 3579 1968 3580 1972
rect 3574 1967 3580 1968
rect 1822 1963 1823 1967
rect 1827 1963 1828 1967
rect 1822 1962 1828 1963
rect 112 1943 114 1962
rect 174 1957 180 1958
rect 174 1953 175 1957
rect 179 1953 180 1957
rect 174 1952 180 1953
rect 286 1957 292 1958
rect 286 1953 287 1957
rect 291 1953 292 1957
rect 286 1952 292 1953
rect 406 1957 412 1958
rect 406 1953 407 1957
rect 411 1953 412 1957
rect 406 1952 412 1953
rect 526 1957 532 1958
rect 526 1953 527 1957
rect 531 1953 532 1957
rect 526 1952 532 1953
rect 646 1957 652 1958
rect 646 1953 647 1957
rect 651 1953 652 1957
rect 646 1952 652 1953
rect 766 1957 772 1958
rect 766 1953 767 1957
rect 771 1953 772 1957
rect 766 1952 772 1953
rect 886 1957 892 1958
rect 886 1953 887 1957
rect 891 1953 892 1957
rect 886 1952 892 1953
rect 1006 1957 1012 1958
rect 1006 1953 1007 1957
rect 1011 1953 1012 1957
rect 1006 1952 1012 1953
rect 1126 1957 1132 1958
rect 1126 1953 1127 1957
rect 1131 1953 1132 1957
rect 1126 1952 1132 1953
rect 1246 1957 1252 1958
rect 1246 1953 1247 1957
rect 1251 1953 1252 1957
rect 1246 1952 1252 1953
rect 176 1943 178 1952
rect 288 1943 290 1952
rect 408 1943 410 1952
rect 528 1943 530 1952
rect 648 1943 650 1952
rect 768 1943 770 1952
rect 888 1943 890 1952
rect 1008 1943 1010 1952
rect 1128 1943 1130 1952
rect 1248 1943 1250 1952
rect 1824 1943 1826 1962
rect 111 1942 115 1943
rect 111 1937 115 1938
rect 135 1942 139 1943
rect 135 1937 139 1938
rect 175 1942 179 1943
rect 175 1937 179 1938
rect 223 1942 227 1943
rect 223 1937 227 1938
rect 287 1942 291 1943
rect 287 1937 291 1938
rect 351 1942 355 1943
rect 351 1937 355 1938
rect 407 1942 411 1943
rect 407 1937 411 1938
rect 495 1942 499 1943
rect 495 1937 499 1938
rect 527 1942 531 1943
rect 527 1937 531 1938
rect 647 1942 651 1943
rect 647 1937 651 1938
rect 655 1942 659 1943
rect 655 1937 659 1938
rect 767 1942 771 1943
rect 767 1937 771 1938
rect 839 1942 843 1943
rect 839 1937 843 1938
rect 887 1942 891 1943
rect 887 1937 891 1938
rect 1007 1942 1011 1943
rect 1007 1937 1011 1938
rect 1039 1942 1043 1943
rect 1039 1937 1043 1938
rect 1127 1942 1131 1943
rect 1127 1937 1131 1938
rect 1247 1942 1251 1943
rect 1247 1937 1251 1938
rect 1463 1942 1467 1943
rect 1463 1937 1467 1938
rect 1823 1942 1827 1943
rect 1823 1937 1827 1938
rect 112 1922 114 1937
rect 136 1932 138 1937
rect 224 1932 226 1937
rect 352 1932 354 1937
rect 496 1932 498 1937
rect 656 1932 658 1937
rect 840 1932 842 1937
rect 1040 1932 1042 1937
rect 1248 1932 1250 1937
rect 1464 1932 1466 1937
rect 134 1931 140 1932
rect 134 1927 135 1931
rect 139 1927 140 1931
rect 134 1926 140 1927
rect 222 1931 228 1932
rect 222 1927 223 1931
rect 227 1927 228 1931
rect 222 1926 228 1927
rect 350 1931 356 1932
rect 350 1927 351 1931
rect 355 1927 356 1931
rect 350 1926 356 1927
rect 494 1931 500 1932
rect 494 1927 495 1931
rect 499 1927 500 1931
rect 494 1926 500 1927
rect 654 1931 660 1932
rect 654 1927 655 1931
rect 659 1927 660 1931
rect 654 1926 660 1927
rect 838 1931 844 1932
rect 838 1927 839 1931
rect 843 1927 844 1931
rect 838 1926 844 1927
rect 1038 1931 1044 1932
rect 1038 1927 1039 1931
rect 1043 1927 1044 1931
rect 1038 1926 1044 1927
rect 1246 1931 1252 1932
rect 1246 1927 1247 1931
rect 1251 1927 1252 1931
rect 1246 1926 1252 1927
rect 1462 1931 1468 1932
rect 1462 1927 1463 1931
rect 1467 1927 1468 1931
rect 1462 1926 1468 1927
rect 1824 1922 1826 1937
rect 1864 1935 1866 1967
rect 1894 1959 1900 1960
rect 1894 1955 1895 1959
rect 1899 1955 1900 1959
rect 1894 1954 1900 1955
rect 2038 1959 2044 1960
rect 2038 1955 2039 1959
rect 2043 1955 2044 1959
rect 2038 1954 2044 1955
rect 2206 1959 2212 1960
rect 2206 1955 2207 1959
rect 2211 1955 2212 1959
rect 2206 1954 2212 1955
rect 2382 1959 2388 1960
rect 2382 1955 2383 1959
rect 2387 1955 2388 1959
rect 2382 1954 2388 1955
rect 2550 1959 2556 1960
rect 2550 1955 2551 1959
rect 2555 1955 2556 1959
rect 2550 1954 2556 1955
rect 2718 1959 2724 1960
rect 2718 1955 2719 1959
rect 2723 1955 2724 1959
rect 2718 1954 2724 1955
rect 2878 1959 2884 1960
rect 2878 1955 2879 1959
rect 2883 1955 2884 1959
rect 2878 1954 2884 1955
rect 3046 1959 3052 1960
rect 3046 1955 3047 1959
rect 3051 1955 3052 1959
rect 3046 1954 3052 1955
rect 3214 1959 3220 1960
rect 3214 1955 3215 1959
rect 3219 1955 3220 1959
rect 3214 1954 3220 1955
rect 1896 1935 1898 1954
rect 2040 1935 2042 1954
rect 2208 1935 2210 1954
rect 2384 1935 2386 1954
rect 2552 1935 2554 1954
rect 2720 1935 2722 1954
rect 2880 1935 2882 1954
rect 3048 1935 3050 1954
rect 3216 1935 3218 1954
rect 3576 1935 3578 1967
rect 1863 1934 1867 1935
rect 1863 1929 1867 1930
rect 1895 1934 1899 1935
rect 1895 1929 1899 1930
rect 1991 1934 1995 1935
rect 1991 1929 1995 1930
rect 2039 1934 2043 1935
rect 2039 1929 2043 1930
rect 2119 1934 2123 1935
rect 2119 1929 2123 1930
rect 2207 1934 2211 1935
rect 2207 1929 2211 1930
rect 2255 1934 2259 1935
rect 2255 1929 2259 1930
rect 2383 1934 2387 1935
rect 2383 1929 2387 1930
rect 2511 1934 2515 1935
rect 2511 1929 2515 1930
rect 2551 1934 2555 1935
rect 2551 1929 2555 1930
rect 2631 1934 2635 1935
rect 2631 1929 2635 1930
rect 2719 1934 2723 1935
rect 2719 1929 2723 1930
rect 2751 1934 2755 1935
rect 2751 1929 2755 1930
rect 2879 1934 2883 1935
rect 2879 1929 2883 1930
rect 3007 1934 3011 1935
rect 3007 1929 3011 1930
rect 3047 1934 3051 1935
rect 3047 1929 3051 1930
rect 3215 1934 3219 1935
rect 3215 1929 3219 1930
rect 3575 1934 3579 1935
rect 3575 1929 3579 1930
rect 110 1921 116 1922
rect 110 1917 111 1921
rect 115 1917 116 1921
rect 110 1916 116 1917
rect 1822 1921 1828 1922
rect 1822 1917 1823 1921
rect 1827 1917 1828 1921
rect 1822 1916 1828 1917
rect 1864 1905 1866 1929
rect 1896 1918 1898 1929
rect 1992 1918 1994 1929
rect 2120 1918 2122 1929
rect 2256 1918 2258 1929
rect 2384 1918 2386 1929
rect 2512 1918 2514 1929
rect 2632 1918 2634 1929
rect 2752 1918 2754 1929
rect 2880 1918 2882 1929
rect 3008 1918 3010 1929
rect 1894 1917 1900 1918
rect 1894 1913 1895 1917
rect 1899 1913 1900 1917
rect 1894 1912 1900 1913
rect 1990 1917 1996 1918
rect 1990 1913 1991 1917
rect 1995 1913 1996 1917
rect 1990 1912 1996 1913
rect 2118 1917 2124 1918
rect 2118 1913 2119 1917
rect 2123 1913 2124 1917
rect 2118 1912 2124 1913
rect 2254 1917 2260 1918
rect 2254 1913 2255 1917
rect 2259 1913 2260 1917
rect 2254 1912 2260 1913
rect 2382 1917 2388 1918
rect 2382 1913 2383 1917
rect 2387 1913 2388 1917
rect 2382 1912 2388 1913
rect 2510 1917 2516 1918
rect 2510 1913 2511 1917
rect 2515 1913 2516 1917
rect 2510 1912 2516 1913
rect 2630 1917 2636 1918
rect 2630 1913 2631 1917
rect 2635 1913 2636 1917
rect 2630 1912 2636 1913
rect 2750 1917 2756 1918
rect 2750 1913 2751 1917
rect 2755 1913 2756 1917
rect 2750 1912 2756 1913
rect 2878 1917 2884 1918
rect 2878 1913 2879 1917
rect 2883 1913 2884 1917
rect 2878 1912 2884 1913
rect 3006 1917 3012 1918
rect 3006 1913 3007 1917
rect 3011 1913 3012 1917
rect 3006 1912 3012 1913
rect 3576 1905 3578 1929
rect 110 1904 116 1905
rect 110 1900 111 1904
rect 115 1900 116 1904
rect 110 1899 116 1900
rect 1822 1904 1828 1905
rect 1822 1900 1823 1904
rect 1827 1900 1828 1904
rect 1822 1899 1828 1900
rect 1862 1904 1868 1905
rect 1862 1900 1863 1904
rect 1867 1900 1868 1904
rect 1862 1899 1868 1900
rect 3574 1904 3580 1905
rect 3574 1900 3575 1904
rect 3579 1900 3580 1904
rect 3574 1899 3580 1900
rect 112 1867 114 1899
rect 142 1891 148 1892
rect 142 1887 143 1891
rect 147 1887 148 1891
rect 142 1886 148 1887
rect 230 1891 236 1892
rect 230 1887 231 1891
rect 235 1887 236 1891
rect 230 1886 236 1887
rect 358 1891 364 1892
rect 358 1887 359 1891
rect 363 1887 364 1891
rect 358 1886 364 1887
rect 502 1891 508 1892
rect 502 1887 503 1891
rect 507 1887 508 1891
rect 502 1886 508 1887
rect 662 1891 668 1892
rect 662 1887 663 1891
rect 667 1887 668 1891
rect 662 1886 668 1887
rect 846 1891 852 1892
rect 846 1887 847 1891
rect 851 1887 852 1891
rect 846 1886 852 1887
rect 1046 1891 1052 1892
rect 1046 1887 1047 1891
rect 1051 1887 1052 1891
rect 1046 1886 1052 1887
rect 1254 1891 1260 1892
rect 1254 1887 1255 1891
rect 1259 1887 1260 1891
rect 1254 1886 1260 1887
rect 1470 1891 1476 1892
rect 1470 1887 1471 1891
rect 1475 1887 1476 1891
rect 1470 1886 1476 1887
rect 144 1867 146 1886
rect 232 1867 234 1886
rect 360 1867 362 1886
rect 504 1867 506 1886
rect 664 1867 666 1886
rect 848 1867 850 1886
rect 1048 1867 1050 1886
rect 1256 1867 1258 1886
rect 1472 1867 1474 1886
rect 1824 1867 1826 1899
rect 1862 1887 1868 1888
rect 1862 1883 1863 1887
rect 1867 1883 1868 1887
rect 1862 1882 1868 1883
rect 3574 1887 3580 1888
rect 3574 1883 3575 1887
rect 3579 1883 3580 1887
rect 3574 1882 3580 1883
rect 111 1866 115 1867
rect 111 1861 115 1862
rect 143 1866 147 1867
rect 143 1861 147 1862
rect 231 1866 235 1867
rect 231 1861 235 1862
rect 271 1866 275 1867
rect 271 1861 275 1862
rect 359 1866 363 1867
rect 359 1861 363 1862
rect 415 1866 419 1867
rect 415 1861 419 1862
rect 503 1866 507 1867
rect 503 1861 507 1862
rect 559 1866 563 1867
rect 559 1861 563 1862
rect 663 1866 667 1867
rect 663 1861 667 1862
rect 695 1866 699 1867
rect 695 1861 699 1862
rect 823 1866 827 1867
rect 823 1861 827 1862
rect 847 1866 851 1867
rect 847 1861 851 1862
rect 943 1866 947 1867
rect 943 1861 947 1862
rect 1047 1866 1051 1867
rect 1047 1861 1051 1862
rect 1055 1866 1059 1867
rect 1055 1861 1059 1862
rect 1159 1866 1163 1867
rect 1159 1861 1163 1862
rect 1255 1866 1259 1867
rect 1255 1861 1259 1862
rect 1263 1866 1267 1867
rect 1263 1861 1267 1862
rect 1359 1866 1363 1867
rect 1359 1861 1363 1862
rect 1455 1866 1459 1867
rect 1455 1861 1459 1862
rect 1471 1866 1475 1867
rect 1471 1861 1475 1862
rect 1551 1866 1555 1867
rect 1551 1861 1555 1862
rect 1647 1866 1651 1867
rect 1647 1861 1651 1862
rect 1735 1866 1739 1867
rect 1735 1861 1739 1862
rect 1823 1866 1827 1867
rect 1823 1861 1827 1862
rect 112 1837 114 1861
rect 144 1850 146 1861
rect 272 1850 274 1861
rect 416 1850 418 1861
rect 560 1850 562 1861
rect 696 1850 698 1861
rect 824 1850 826 1861
rect 944 1850 946 1861
rect 1056 1850 1058 1861
rect 1160 1850 1162 1861
rect 1264 1850 1266 1861
rect 1360 1850 1362 1861
rect 1456 1850 1458 1861
rect 1552 1850 1554 1861
rect 1648 1850 1650 1861
rect 1736 1850 1738 1861
rect 142 1849 148 1850
rect 142 1845 143 1849
rect 147 1845 148 1849
rect 142 1844 148 1845
rect 270 1849 276 1850
rect 270 1845 271 1849
rect 275 1845 276 1849
rect 270 1844 276 1845
rect 414 1849 420 1850
rect 414 1845 415 1849
rect 419 1845 420 1849
rect 414 1844 420 1845
rect 558 1849 564 1850
rect 558 1845 559 1849
rect 563 1845 564 1849
rect 558 1844 564 1845
rect 694 1849 700 1850
rect 694 1845 695 1849
rect 699 1845 700 1849
rect 694 1844 700 1845
rect 822 1849 828 1850
rect 822 1845 823 1849
rect 827 1845 828 1849
rect 822 1844 828 1845
rect 942 1849 948 1850
rect 942 1845 943 1849
rect 947 1845 948 1849
rect 942 1844 948 1845
rect 1054 1849 1060 1850
rect 1054 1845 1055 1849
rect 1059 1845 1060 1849
rect 1054 1844 1060 1845
rect 1158 1849 1164 1850
rect 1158 1845 1159 1849
rect 1163 1845 1164 1849
rect 1158 1844 1164 1845
rect 1262 1849 1268 1850
rect 1262 1845 1263 1849
rect 1267 1845 1268 1849
rect 1262 1844 1268 1845
rect 1358 1849 1364 1850
rect 1358 1845 1359 1849
rect 1363 1845 1364 1849
rect 1358 1844 1364 1845
rect 1454 1849 1460 1850
rect 1454 1845 1455 1849
rect 1459 1845 1460 1849
rect 1454 1844 1460 1845
rect 1550 1849 1556 1850
rect 1550 1845 1551 1849
rect 1555 1845 1556 1849
rect 1550 1844 1556 1845
rect 1646 1849 1652 1850
rect 1646 1845 1647 1849
rect 1651 1845 1652 1849
rect 1646 1844 1652 1845
rect 1734 1849 1740 1850
rect 1734 1845 1735 1849
rect 1739 1845 1740 1849
rect 1734 1844 1740 1845
rect 1824 1837 1826 1861
rect 1864 1859 1866 1882
rect 1886 1877 1892 1878
rect 1886 1873 1887 1877
rect 1891 1873 1892 1877
rect 1886 1872 1892 1873
rect 1982 1877 1988 1878
rect 1982 1873 1983 1877
rect 1987 1873 1988 1877
rect 1982 1872 1988 1873
rect 2110 1877 2116 1878
rect 2110 1873 2111 1877
rect 2115 1873 2116 1877
rect 2110 1872 2116 1873
rect 2246 1877 2252 1878
rect 2246 1873 2247 1877
rect 2251 1873 2252 1877
rect 2246 1872 2252 1873
rect 2374 1877 2380 1878
rect 2374 1873 2375 1877
rect 2379 1873 2380 1877
rect 2374 1872 2380 1873
rect 2502 1877 2508 1878
rect 2502 1873 2503 1877
rect 2507 1873 2508 1877
rect 2502 1872 2508 1873
rect 2622 1877 2628 1878
rect 2622 1873 2623 1877
rect 2627 1873 2628 1877
rect 2622 1872 2628 1873
rect 2742 1877 2748 1878
rect 2742 1873 2743 1877
rect 2747 1873 2748 1877
rect 2742 1872 2748 1873
rect 2870 1877 2876 1878
rect 2870 1873 2871 1877
rect 2875 1873 2876 1877
rect 2870 1872 2876 1873
rect 2998 1877 3004 1878
rect 2998 1873 2999 1877
rect 3003 1873 3004 1877
rect 2998 1872 3004 1873
rect 1888 1859 1890 1872
rect 1984 1859 1986 1872
rect 2112 1859 2114 1872
rect 2248 1859 2250 1872
rect 2376 1859 2378 1872
rect 2504 1859 2506 1872
rect 2624 1859 2626 1872
rect 2744 1859 2746 1872
rect 2872 1859 2874 1872
rect 3000 1859 3002 1872
rect 3576 1859 3578 1882
rect 1863 1858 1867 1859
rect 1863 1853 1867 1854
rect 1887 1858 1891 1859
rect 1887 1853 1891 1854
rect 1983 1858 1987 1859
rect 1983 1853 1987 1854
rect 2111 1858 2115 1859
rect 2111 1853 2115 1854
rect 2223 1858 2227 1859
rect 2223 1853 2227 1854
rect 2247 1858 2251 1859
rect 2247 1853 2251 1854
rect 2359 1858 2363 1859
rect 2359 1853 2363 1854
rect 2375 1858 2379 1859
rect 2375 1853 2379 1854
rect 2495 1858 2499 1859
rect 2495 1853 2499 1854
rect 2503 1858 2507 1859
rect 2503 1853 2507 1854
rect 2623 1858 2627 1859
rect 2623 1853 2627 1854
rect 2743 1858 2747 1859
rect 2743 1853 2747 1854
rect 2863 1858 2867 1859
rect 2863 1853 2867 1854
rect 2871 1858 2875 1859
rect 2871 1853 2875 1854
rect 2991 1858 2995 1859
rect 2991 1853 2995 1854
rect 2999 1858 3003 1859
rect 2999 1853 3003 1854
rect 3575 1858 3579 1859
rect 3575 1853 3579 1854
rect 1864 1838 1866 1853
rect 2224 1848 2226 1853
rect 2360 1848 2362 1853
rect 2496 1848 2498 1853
rect 2624 1848 2626 1853
rect 2744 1848 2746 1853
rect 2864 1848 2866 1853
rect 2992 1848 2994 1853
rect 2222 1847 2228 1848
rect 2222 1843 2223 1847
rect 2227 1843 2228 1847
rect 2222 1842 2228 1843
rect 2358 1847 2364 1848
rect 2358 1843 2359 1847
rect 2363 1843 2364 1847
rect 2358 1842 2364 1843
rect 2494 1847 2500 1848
rect 2494 1843 2495 1847
rect 2499 1843 2500 1847
rect 2494 1842 2500 1843
rect 2622 1847 2628 1848
rect 2622 1843 2623 1847
rect 2627 1843 2628 1847
rect 2622 1842 2628 1843
rect 2742 1847 2748 1848
rect 2742 1843 2743 1847
rect 2747 1843 2748 1847
rect 2742 1842 2748 1843
rect 2862 1847 2868 1848
rect 2862 1843 2863 1847
rect 2867 1843 2868 1847
rect 2862 1842 2868 1843
rect 2990 1847 2996 1848
rect 2990 1843 2991 1847
rect 2995 1843 2996 1847
rect 2990 1842 2996 1843
rect 3576 1838 3578 1853
rect 1862 1837 1868 1838
rect 110 1836 116 1837
rect 110 1832 111 1836
rect 115 1832 116 1836
rect 110 1831 116 1832
rect 1822 1836 1828 1837
rect 1822 1832 1823 1836
rect 1827 1832 1828 1836
rect 1862 1833 1863 1837
rect 1867 1833 1868 1837
rect 1862 1832 1868 1833
rect 3574 1837 3580 1838
rect 3574 1833 3575 1837
rect 3579 1833 3580 1837
rect 3574 1832 3580 1833
rect 1822 1831 1828 1832
rect 1862 1820 1868 1821
rect 110 1819 116 1820
rect 110 1815 111 1819
rect 115 1815 116 1819
rect 110 1814 116 1815
rect 1822 1819 1828 1820
rect 1822 1815 1823 1819
rect 1827 1815 1828 1819
rect 1862 1816 1863 1820
rect 1867 1816 1868 1820
rect 1862 1815 1868 1816
rect 3574 1820 3580 1821
rect 3574 1816 3575 1820
rect 3579 1816 3580 1820
rect 3574 1815 3580 1816
rect 1822 1814 1828 1815
rect 112 1787 114 1814
rect 134 1809 140 1810
rect 134 1805 135 1809
rect 139 1805 140 1809
rect 134 1804 140 1805
rect 262 1809 268 1810
rect 262 1805 263 1809
rect 267 1805 268 1809
rect 262 1804 268 1805
rect 406 1809 412 1810
rect 406 1805 407 1809
rect 411 1805 412 1809
rect 406 1804 412 1805
rect 550 1809 556 1810
rect 550 1805 551 1809
rect 555 1805 556 1809
rect 550 1804 556 1805
rect 686 1809 692 1810
rect 686 1805 687 1809
rect 691 1805 692 1809
rect 686 1804 692 1805
rect 814 1809 820 1810
rect 814 1805 815 1809
rect 819 1805 820 1809
rect 814 1804 820 1805
rect 934 1809 940 1810
rect 934 1805 935 1809
rect 939 1805 940 1809
rect 934 1804 940 1805
rect 1046 1809 1052 1810
rect 1046 1805 1047 1809
rect 1051 1805 1052 1809
rect 1046 1804 1052 1805
rect 1150 1809 1156 1810
rect 1150 1805 1151 1809
rect 1155 1805 1156 1809
rect 1150 1804 1156 1805
rect 1254 1809 1260 1810
rect 1254 1805 1255 1809
rect 1259 1805 1260 1809
rect 1254 1804 1260 1805
rect 1350 1809 1356 1810
rect 1350 1805 1351 1809
rect 1355 1805 1356 1809
rect 1350 1804 1356 1805
rect 1446 1809 1452 1810
rect 1446 1805 1447 1809
rect 1451 1805 1452 1809
rect 1446 1804 1452 1805
rect 1542 1809 1548 1810
rect 1542 1805 1543 1809
rect 1547 1805 1548 1809
rect 1542 1804 1548 1805
rect 1638 1809 1644 1810
rect 1638 1805 1639 1809
rect 1643 1805 1644 1809
rect 1638 1804 1644 1805
rect 1726 1809 1732 1810
rect 1726 1805 1727 1809
rect 1731 1805 1732 1809
rect 1726 1804 1732 1805
rect 136 1787 138 1804
rect 264 1787 266 1804
rect 408 1787 410 1804
rect 552 1787 554 1804
rect 688 1787 690 1804
rect 816 1787 818 1804
rect 936 1787 938 1804
rect 1048 1787 1050 1804
rect 1152 1787 1154 1804
rect 1256 1787 1258 1804
rect 1352 1787 1354 1804
rect 1448 1787 1450 1804
rect 1544 1787 1546 1804
rect 1640 1787 1642 1804
rect 1728 1787 1730 1804
rect 1824 1787 1826 1814
rect 1864 1787 1866 1815
rect 2230 1807 2236 1808
rect 2230 1803 2231 1807
rect 2235 1803 2236 1807
rect 2230 1802 2236 1803
rect 2366 1807 2372 1808
rect 2366 1803 2367 1807
rect 2371 1803 2372 1807
rect 2366 1802 2372 1803
rect 2502 1807 2508 1808
rect 2502 1803 2503 1807
rect 2507 1803 2508 1807
rect 2502 1802 2508 1803
rect 2630 1807 2636 1808
rect 2630 1803 2631 1807
rect 2635 1803 2636 1807
rect 2630 1802 2636 1803
rect 2750 1807 2756 1808
rect 2750 1803 2751 1807
rect 2755 1803 2756 1807
rect 2750 1802 2756 1803
rect 2870 1807 2876 1808
rect 2870 1803 2871 1807
rect 2875 1803 2876 1807
rect 2870 1802 2876 1803
rect 2998 1807 3004 1808
rect 2998 1803 2999 1807
rect 3003 1803 3004 1807
rect 2998 1802 3004 1803
rect 2232 1787 2234 1802
rect 2368 1787 2370 1802
rect 2504 1787 2506 1802
rect 2632 1787 2634 1802
rect 2752 1787 2754 1802
rect 2872 1787 2874 1802
rect 3000 1787 3002 1802
rect 3576 1787 3578 1815
rect 111 1786 115 1787
rect 111 1781 115 1782
rect 135 1786 139 1787
rect 135 1781 139 1782
rect 263 1786 267 1787
rect 263 1781 267 1782
rect 303 1786 307 1787
rect 303 1781 307 1782
rect 407 1786 411 1787
rect 407 1781 411 1782
rect 495 1786 499 1787
rect 495 1781 499 1782
rect 551 1786 555 1787
rect 551 1781 555 1782
rect 687 1786 691 1787
rect 687 1781 691 1782
rect 815 1786 819 1787
rect 815 1781 819 1782
rect 871 1786 875 1787
rect 871 1781 875 1782
rect 935 1786 939 1787
rect 935 1781 939 1782
rect 1047 1786 1051 1787
rect 1047 1781 1051 1782
rect 1151 1786 1155 1787
rect 1151 1781 1155 1782
rect 1215 1786 1219 1787
rect 1215 1781 1219 1782
rect 1255 1786 1259 1787
rect 1255 1781 1259 1782
rect 1351 1786 1355 1787
rect 1351 1781 1355 1782
rect 1375 1786 1379 1787
rect 1375 1781 1379 1782
rect 1447 1786 1451 1787
rect 1447 1781 1451 1782
rect 1535 1786 1539 1787
rect 1535 1781 1539 1782
rect 1543 1786 1547 1787
rect 1543 1781 1547 1782
rect 1639 1786 1643 1787
rect 1639 1781 1643 1782
rect 1703 1786 1707 1787
rect 1703 1781 1707 1782
rect 1727 1786 1731 1787
rect 1727 1781 1731 1782
rect 1823 1786 1827 1787
rect 1823 1781 1827 1782
rect 1863 1786 1867 1787
rect 1863 1781 1867 1782
rect 2231 1786 2235 1787
rect 2231 1781 2235 1782
rect 2271 1786 2275 1787
rect 2271 1781 2275 1782
rect 2359 1786 2363 1787
rect 2359 1781 2363 1782
rect 2367 1786 2371 1787
rect 2367 1781 2371 1782
rect 2455 1786 2459 1787
rect 2455 1781 2459 1782
rect 2503 1786 2507 1787
rect 2503 1781 2507 1782
rect 2559 1786 2563 1787
rect 2559 1781 2563 1782
rect 2631 1786 2635 1787
rect 2631 1781 2635 1782
rect 2663 1786 2667 1787
rect 2663 1781 2667 1782
rect 2751 1786 2755 1787
rect 2751 1781 2755 1782
rect 2759 1786 2763 1787
rect 2759 1781 2763 1782
rect 2863 1786 2867 1787
rect 2863 1781 2867 1782
rect 2871 1786 2875 1787
rect 2871 1781 2875 1782
rect 2967 1786 2971 1787
rect 2967 1781 2971 1782
rect 2999 1786 3003 1787
rect 2999 1781 3003 1782
rect 3071 1786 3075 1787
rect 3071 1781 3075 1782
rect 3175 1786 3179 1787
rect 3175 1781 3179 1782
rect 3575 1786 3579 1787
rect 3575 1781 3579 1782
rect 112 1766 114 1781
rect 136 1776 138 1781
rect 304 1776 306 1781
rect 496 1776 498 1781
rect 688 1776 690 1781
rect 872 1776 874 1781
rect 1048 1776 1050 1781
rect 1216 1776 1218 1781
rect 1376 1776 1378 1781
rect 1536 1776 1538 1781
rect 1704 1776 1706 1781
rect 134 1775 140 1776
rect 134 1771 135 1775
rect 139 1771 140 1775
rect 134 1770 140 1771
rect 302 1775 308 1776
rect 302 1771 303 1775
rect 307 1771 308 1775
rect 302 1770 308 1771
rect 494 1775 500 1776
rect 494 1771 495 1775
rect 499 1771 500 1775
rect 494 1770 500 1771
rect 686 1775 692 1776
rect 686 1771 687 1775
rect 691 1771 692 1775
rect 686 1770 692 1771
rect 870 1775 876 1776
rect 870 1771 871 1775
rect 875 1771 876 1775
rect 870 1770 876 1771
rect 1046 1775 1052 1776
rect 1046 1771 1047 1775
rect 1051 1771 1052 1775
rect 1046 1770 1052 1771
rect 1214 1775 1220 1776
rect 1214 1771 1215 1775
rect 1219 1771 1220 1775
rect 1214 1770 1220 1771
rect 1374 1775 1380 1776
rect 1374 1771 1375 1775
rect 1379 1771 1380 1775
rect 1374 1770 1380 1771
rect 1534 1775 1540 1776
rect 1534 1771 1535 1775
rect 1539 1771 1540 1775
rect 1534 1770 1540 1771
rect 1702 1775 1708 1776
rect 1702 1771 1703 1775
rect 1707 1771 1708 1775
rect 1702 1770 1708 1771
rect 1824 1766 1826 1781
rect 110 1765 116 1766
rect 110 1761 111 1765
rect 115 1761 116 1765
rect 110 1760 116 1761
rect 1822 1765 1828 1766
rect 1822 1761 1823 1765
rect 1827 1761 1828 1765
rect 1822 1760 1828 1761
rect 1864 1757 1866 1781
rect 2272 1770 2274 1781
rect 2360 1770 2362 1781
rect 2456 1770 2458 1781
rect 2560 1770 2562 1781
rect 2664 1770 2666 1781
rect 2760 1770 2762 1781
rect 2864 1770 2866 1781
rect 2968 1770 2970 1781
rect 3072 1770 3074 1781
rect 3176 1770 3178 1781
rect 2270 1769 2276 1770
rect 2270 1765 2271 1769
rect 2275 1765 2276 1769
rect 2270 1764 2276 1765
rect 2358 1769 2364 1770
rect 2358 1765 2359 1769
rect 2363 1765 2364 1769
rect 2358 1764 2364 1765
rect 2454 1769 2460 1770
rect 2454 1765 2455 1769
rect 2459 1765 2460 1769
rect 2454 1764 2460 1765
rect 2558 1769 2564 1770
rect 2558 1765 2559 1769
rect 2563 1765 2564 1769
rect 2558 1764 2564 1765
rect 2662 1769 2668 1770
rect 2662 1765 2663 1769
rect 2667 1765 2668 1769
rect 2662 1764 2668 1765
rect 2758 1769 2764 1770
rect 2758 1765 2759 1769
rect 2763 1765 2764 1769
rect 2758 1764 2764 1765
rect 2862 1769 2868 1770
rect 2862 1765 2863 1769
rect 2867 1765 2868 1769
rect 2862 1764 2868 1765
rect 2966 1769 2972 1770
rect 2966 1765 2967 1769
rect 2971 1765 2972 1769
rect 2966 1764 2972 1765
rect 3070 1769 3076 1770
rect 3070 1765 3071 1769
rect 3075 1765 3076 1769
rect 3070 1764 3076 1765
rect 3174 1769 3180 1770
rect 3174 1765 3175 1769
rect 3179 1765 3180 1769
rect 3174 1764 3180 1765
rect 3576 1757 3578 1781
rect 1862 1756 1868 1757
rect 1862 1752 1863 1756
rect 1867 1752 1868 1756
rect 1862 1751 1868 1752
rect 3574 1756 3580 1757
rect 3574 1752 3575 1756
rect 3579 1752 3580 1756
rect 3574 1751 3580 1752
rect 110 1748 116 1749
rect 110 1744 111 1748
rect 115 1744 116 1748
rect 110 1743 116 1744
rect 1822 1748 1828 1749
rect 1822 1744 1823 1748
rect 1827 1744 1828 1748
rect 1822 1743 1828 1744
rect 112 1715 114 1743
rect 142 1735 148 1736
rect 142 1731 143 1735
rect 147 1731 148 1735
rect 142 1730 148 1731
rect 310 1735 316 1736
rect 310 1731 311 1735
rect 315 1731 316 1735
rect 310 1730 316 1731
rect 502 1735 508 1736
rect 502 1731 503 1735
rect 507 1731 508 1735
rect 502 1730 508 1731
rect 694 1735 700 1736
rect 694 1731 695 1735
rect 699 1731 700 1735
rect 694 1730 700 1731
rect 878 1735 884 1736
rect 878 1731 879 1735
rect 883 1731 884 1735
rect 878 1730 884 1731
rect 1054 1735 1060 1736
rect 1054 1731 1055 1735
rect 1059 1731 1060 1735
rect 1054 1730 1060 1731
rect 1222 1735 1228 1736
rect 1222 1731 1223 1735
rect 1227 1731 1228 1735
rect 1222 1730 1228 1731
rect 1382 1735 1388 1736
rect 1382 1731 1383 1735
rect 1387 1731 1388 1735
rect 1382 1730 1388 1731
rect 1542 1735 1548 1736
rect 1542 1731 1543 1735
rect 1547 1731 1548 1735
rect 1542 1730 1548 1731
rect 1710 1735 1716 1736
rect 1710 1731 1711 1735
rect 1715 1731 1716 1735
rect 1710 1730 1716 1731
rect 144 1715 146 1730
rect 312 1715 314 1730
rect 504 1715 506 1730
rect 696 1715 698 1730
rect 880 1715 882 1730
rect 1056 1715 1058 1730
rect 1224 1715 1226 1730
rect 1384 1715 1386 1730
rect 1544 1715 1546 1730
rect 1712 1715 1714 1730
rect 1824 1715 1826 1743
rect 1862 1739 1868 1740
rect 1862 1735 1863 1739
rect 1867 1735 1868 1739
rect 1862 1734 1868 1735
rect 3574 1739 3580 1740
rect 3574 1735 3575 1739
rect 3579 1735 3580 1739
rect 3574 1734 3580 1735
rect 1864 1715 1866 1734
rect 2262 1729 2268 1730
rect 2262 1725 2263 1729
rect 2267 1725 2268 1729
rect 2262 1724 2268 1725
rect 2350 1729 2356 1730
rect 2350 1725 2351 1729
rect 2355 1725 2356 1729
rect 2350 1724 2356 1725
rect 2446 1729 2452 1730
rect 2446 1725 2447 1729
rect 2451 1725 2452 1729
rect 2446 1724 2452 1725
rect 2550 1729 2556 1730
rect 2550 1725 2551 1729
rect 2555 1725 2556 1729
rect 2550 1724 2556 1725
rect 2654 1729 2660 1730
rect 2654 1725 2655 1729
rect 2659 1725 2660 1729
rect 2654 1724 2660 1725
rect 2750 1729 2756 1730
rect 2750 1725 2751 1729
rect 2755 1725 2756 1729
rect 2750 1724 2756 1725
rect 2854 1729 2860 1730
rect 2854 1725 2855 1729
rect 2859 1725 2860 1729
rect 2854 1724 2860 1725
rect 2958 1729 2964 1730
rect 2958 1725 2959 1729
rect 2963 1725 2964 1729
rect 2958 1724 2964 1725
rect 3062 1729 3068 1730
rect 3062 1725 3063 1729
rect 3067 1725 3068 1729
rect 3062 1724 3068 1725
rect 3166 1729 3172 1730
rect 3166 1725 3167 1729
rect 3171 1725 3172 1729
rect 3166 1724 3172 1725
rect 2264 1715 2266 1724
rect 2352 1715 2354 1724
rect 2448 1715 2450 1724
rect 2552 1715 2554 1724
rect 2656 1715 2658 1724
rect 2752 1715 2754 1724
rect 2856 1715 2858 1724
rect 2960 1715 2962 1724
rect 3064 1715 3066 1724
rect 3168 1715 3170 1724
rect 3576 1715 3578 1734
rect 111 1714 115 1715
rect 111 1709 115 1710
rect 143 1714 147 1715
rect 143 1709 147 1710
rect 287 1714 291 1715
rect 287 1709 291 1710
rect 311 1714 315 1715
rect 311 1709 315 1710
rect 471 1714 475 1715
rect 471 1709 475 1710
rect 503 1714 507 1715
rect 503 1709 507 1710
rect 655 1714 659 1715
rect 655 1709 659 1710
rect 695 1714 699 1715
rect 695 1709 699 1710
rect 839 1714 843 1715
rect 839 1709 843 1710
rect 879 1714 883 1715
rect 879 1709 883 1710
rect 1023 1714 1027 1715
rect 1023 1709 1027 1710
rect 1055 1714 1059 1715
rect 1055 1709 1059 1710
rect 1191 1714 1195 1715
rect 1191 1709 1195 1710
rect 1223 1714 1227 1715
rect 1223 1709 1227 1710
rect 1359 1714 1363 1715
rect 1359 1709 1363 1710
rect 1383 1714 1387 1715
rect 1383 1709 1387 1710
rect 1527 1714 1531 1715
rect 1527 1709 1531 1710
rect 1543 1714 1547 1715
rect 1543 1709 1547 1710
rect 1695 1714 1699 1715
rect 1695 1709 1699 1710
rect 1711 1714 1715 1715
rect 1711 1709 1715 1710
rect 1823 1714 1827 1715
rect 1823 1709 1827 1710
rect 1863 1714 1867 1715
rect 1863 1709 1867 1710
rect 2247 1714 2251 1715
rect 2247 1709 2251 1710
rect 2263 1714 2267 1715
rect 2263 1709 2267 1710
rect 2351 1714 2355 1715
rect 2351 1709 2355 1710
rect 2367 1714 2371 1715
rect 2367 1709 2371 1710
rect 2447 1714 2451 1715
rect 2447 1709 2451 1710
rect 2495 1714 2499 1715
rect 2495 1709 2499 1710
rect 2551 1714 2555 1715
rect 2551 1709 2555 1710
rect 2623 1714 2627 1715
rect 2623 1709 2627 1710
rect 2655 1714 2659 1715
rect 2655 1709 2659 1710
rect 2751 1714 2755 1715
rect 2751 1709 2755 1710
rect 2759 1714 2763 1715
rect 2759 1709 2763 1710
rect 2855 1714 2859 1715
rect 2855 1709 2859 1710
rect 2887 1714 2891 1715
rect 2887 1709 2891 1710
rect 2959 1714 2963 1715
rect 2959 1709 2963 1710
rect 3015 1714 3019 1715
rect 3015 1709 3019 1710
rect 3063 1714 3067 1715
rect 3063 1709 3067 1710
rect 3135 1714 3139 1715
rect 3135 1709 3139 1710
rect 3167 1714 3171 1715
rect 3167 1709 3171 1710
rect 3247 1714 3251 1715
rect 3247 1709 3251 1710
rect 3367 1714 3371 1715
rect 3367 1709 3371 1710
rect 3479 1714 3483 1715
rect 3479 1709 3483 1710
rect 3575 1714 3579 1715
rect 3575 1709 3579 1710
rect 112 1685 114 1709
rect 144 1698 146 1709
rect 288 1698 290 1709
rect 472 1698 474 1709
rect 656 1698 658 1709
rect 840 1698 842 1709
rect 1024 1698 1026 1709
rect 1192 1698 1194 1709
rect 1360 1698 1362 1709
rect 1528 1698 1530 1709
rect 1696 1698 1698 1709
rect 142 1697 148 1698
rect 142 1693 143 1697
rect 147 1693 148 1697
rect 142 1692 148 1693
rect 286 1697 292 1698
rect 286 1693 287 1697
rect 291 1693 292 1697
rect 286 1692 292 1693
rect 470 1697 476 1698
rect 470 1693 471 1697
rect 475 1693 476 1697
rect 470 1692 476 1693
rect 654 1697 660 1698
rect 654 1693 655 1697
rect 659 1693 660 1697
rect 654 1692 660 1693
rect 838 1697 844 1698
rect 838 1693 839 1697
rect 843 1693 844 1697
rect 838 1692 844 1693
rect 1022 1697 1028 1698
rect 1022 1693 1023 1697
rect 1027 1693 1028 1697
rect 1022 1692 1028 1693
rect 1190 1697 1196 1698
rect 1190 1693 1191 1697
rect 1195 1693 1196 1697
rect 1190 1692 1196 1693
rect 1358 1697 1364 1698
rect 1358 1693 1359 1697
rect 1363 1693 1364 1697
rect 1358 1692 1364 1693
rect 1526 1697 1532 1698
rect 1526 1693 1527 1697
rect 1531 1693 1532 1697
rect 1526 1692 1532 1693
rect 1694 1697 1700 1698
rect 1694 1693 1695 1697
rect 1699 1693 1700 1697
rect 1694 1692 1700 1693
rect 1824 1685 1826 1709
rect 1864 1694 1866 1709
rect 2248 1704 2250 1709
rect 2368 1704 2370 1709
rect 2496 1704 2498 1709
rect 2624 1704 2626 1709
rect 2760 1704 2762 1709
rect 2888 1704 2890 1709
rect 3016 1704 3018 1709
rect 3136 1704 3138 1709
rect 3248 1704 3250 1709
rect 3368 1704 3370 1709
rect 3480 1704 3482 1709
rect 2246 1703 2252 1704
rect 2246 1699 2247 1703
rect 2251 1699 2252 1703
rect 2246 1698 2252 1699
rect 2366 1703 2372 1704
rect 2366 1699 2367 1703
rect 2371 1699 2372 1703
rect 2366 1698 2372 1699
rect 2494 1703 2500 1704
rect 2494 1699 2495 1703
rect 2499 1699 2500 1703
rect 2494 1698 2500 1699
rect 2622 1703 2628 1704
rect 2622 1699 2623 1703
rect 2627 1699 2628 1703
rect 2622 1698 2628 1699
rect 2758 1703 2764 1704
rect 2758 1699 2759 1703
rect 2763 1699 2764 1703
rect 2758 1698 2764 1699
rect 2886 1703 2892 1704
rect 2886 1699 2887 1703
rect 2891 1699 2892 1703
rect 2886 1698 2892 1699
rect 3014 1703 3020 1704
rect 3014 1699 3015 1703
rect 3019 1699 3020 1703
rect 3014 1698 3020 1699
rect 3134 1703 3140 1704
rect 3134 1699 3135 1703
rect 3139 1699 3140 1703
rect 3134 1698 3140 1699
rect 3246 1703 3252 1704
rect 3246 1699 3247 1703
rect 3251 1699 3252 1703
rect 3246 1698 3252 1699
rect 3366 1703 3372 1704
rect 3366 1699 3367 1703
rect 3371 1699 3372 1703
rect 3366 1698 3372 1699
rect 3478 1703 3484 1704
rect 3478 1699 3479 1703
rect 3483 1699 3484 1703
rect 3478 1698 3484 1699
rect 3576 1694 3578 1709
rect 1862 1693 1868 1694
rect 1862 1689 1863 1693
rect 1867 1689 1868 1693
rect 1862 1688 1868 1689
rect 3574 1693 3580 1694
rect 3574 1689 3575 1693
rect 3579 1689 3580 1693
rect 3574 1688 3580 1689
rect 110 1684 116 1685
rect 110 1680 111 1684
rect 115 1680 116 1684
rect 110 1679 116 1680
rect 1822 1684 1828 1685
rect 1822 1680 1823 1684
rect 1827 1680 1828 1684
rect 1822 1679 1828 1680
rect 1862 1676 1868 1677
rect 1862 1672 1863 1676
rect 1867 1672 1868 1676
rect 1862 1671 1868 1672
rect 3574 1676 3580 1677
rect 3574 1672 3575 1676
rect 3579 1672 3580 1676
rect 3574 1671 3580 1672
rect 110 1667 116 1668
rect 110 1663 111 1667
rect 115 1663 116 1667
rect 110 1662 116 1663
rect 1822 1667 1828 1668
rect 1822 1663 1823 1667
rect 1827 1663 1828 1667
rect 1822 1662 1828 1663
rect 112 1639 114 1662
rect 134 1657 140 1658
rect 134 1653 135 1657
rect 139 1653 140 1657
rect 134 1652 140 1653
rect 278 1657 284 1658
rect 278 1653 279 1657
rect 283 1653 284 1657
rect 278 1652 284 1653
rect 462 1657 468 1658
rect 462 1653 463 1657
rect 467 1653 468 1657
rect 462 1652 468 1653
rect 646 1657 652 1658
rect 646 1653 647 1657
rect 651 1653 652 1657
rect 646 1652 652 1653
rect 830 1657 836 1658
rect 830 1653 831 1657
rect 835 1653 836 1657
rect 830 1652 836 1653
rect 1014 1657 1020 1658
rect 1014 1653 1015 1657
rect 1019 1653 1020 1657
rect 1014 1652 1020 1653
rect 1182 1657 1188 1658
rect 1182 1653 1183 1657
rect 1187 1653 1188 1657
rect 1182 1652 1188 1653
rect 1350 1657 1356 1658
rect 1350 1653 1351 1657
rect 1355 1653 1356 1657
rect 1350 1652 1356 1653
rect 1518 1657 1524 1658
rect 1518 1653 1519 1657
rect 1523 1653 1524 1657
rect 1518 1652 1524 1653
rect 1686 1657 1692 1658
rect 1686 1653 1687 1657
rect 1691 1653 1692 1657
rect 1686 1652 1692 1653
rect 136 1639 138 1652
rect 280 1639 282 1652
rect 464 1639 466 1652
rect 648 1639 650 1652
rect 832 1639 834 1652
rect 1016 1639 1018 1652
rect 1184 1639 1186 1652
rect 1352 1639 1354 1652
rect 1520 1639 1522 1652
rect 1688 1639 1690 1652
rect 1824 1639 1826 1662
rect 1864 1643 1866 1671
rect 2254 1663 2260 1664
rect 2254 1659 2255 1663
rect 2259 1659 2260 1663
rect 2254 1658 2260 1659
rect 2374 1663 2380 1664
rect 2374 1659 2375 1663
rect 2379 1659 2380 1663
rect 2374 1658 2380 1659
rect 2502 1663 2508 1664
rect 2502 1659 2503 1663
rect 2507 1659 2508 1663
rect 2502 1658 2508 1659
rect 2630 1663 2636 1664
rect 2630 1659 2631 1663
rect 2635 1659 2636 1663
rect 2630 1658 2636 1659
rect 2766 1663 2772 1664
rect 2766 1659 2767 1663
rect 2771 1659 2772 1663
rect 2766 1658 2772 1659
rect 2894 1663 2900 1664
rect 2894 1659 2895 1663
rect 2899 1659 2900 1663
rect 2894 1658 2900 1659
rect 3022 1663 3028 1664
rect 3022 1659 3023 1663
rect 3027 1659 3028 1663
rect 3022 1658 3028 1659
rect 3142 1663 3148 1664
rect 3142 1659 3143 1663
rect 3147 1659 3148 1663
rect 3142 1658 3148 1659
rect 3254 1663 3260 1664
rect 3254 1659 3255 1663
rect 3259 1659 3260 1663
rect 3254 1658 3260 1659
rect 3374 1663 3380 1664
rect 3374 1659 3375 1663
rect 3379 1659 3380 1663
rect 3374 1658 3380 1659
rect 3486 1663 3492 1664
rect 3486 1659 3487 1663
rect 3491 1659 3492 1663
rect 3486 1658 3492 1659
rect 2256 1643 2258 1658
rect 2376 1643 2378 1658
rect 2504 1643 2506 1658
rect 2632 1643 2634 1658
rect 2768 1643 2770 1658
rect 2896 1643 2898 1658
rect 3024 1643 3026 1658
rect 3144 1643 3146 1658
rect 3256 1643 3258 1658
rect 3376 1643 3378 1658
rect 3488 1643 3490 1658
rect 3576 1643 3578 1671
rect 1863 1642 1867 1643
rect 111 1638 115 1639
rect 111 1633 115 1634
rect 135 1638 139 1639
rect 135 1633 139 1634
rect 271 1638 275 1639
rect 271 1633 275 1634
rect 279 1638 283 1639
rect 279 1633 283 1634
rect 447 1638 451 1639
rect 447 1633 451 1634
rect 463 1638 467 1639
rect 463 1633 467 1634
rect 631 1638 635 1639
rect 631 1633 635 1634
rect 647 1638 651 1639
rect 647 1633 651 1634
rect 815 1638 819 1639
rect 815 1633 819 1634
rect 831 1638 835 1639
rect 831 1633 835 1634
rect 991 1638 995 1639
rect 991 1633 995 1634
rect 1015 1638 1019 1639
rect 1015 1633 1019 1634
rect 1151 1638 1155 1639
rect 1151 1633 1155 1634
rect 1183 1638 1187 1639
rect 1183 1633 1187 1634
rect 1303 1638 1307 1639
rect 1303 1633 1307 1634
rect 1351 1638 1355 1639
rect 1351 1633 1355 1634
rect 1455 1638 1459 1639
rect 1455 1633 1459 1634
rect 1519 1638 1523 1639
rect 1519 1633 1523 1634
rect 1599 1638 1603 1639
rect 1599 1633 1603 1634
rect 1687 1638 1691 1639
rect 1687 1633 1691 1634
rect 1727 1638 1731 1639
rect 1727 1633 1731 1634
rect 1823 1638 1827 1639
rect 1863 1637 1867 1638
rect 2151 1642 2155 1643
rect 2151 1637 2155 1638
rect 2255 1642 2259 1643
rect 2255 1637 2259 1638
rect 2343 1642 2347 1643
rect 2343 1637 2347 1638
rect 2375 1642 2379 1643
rect 2375 1637 2379 1638
rect 2503 1642 2507 1643
rect 2503 1637 2507 1638
rect 2527 1642 2531 1643
rect 2527 1637 2531 1638
rect 2631 1642 2635 1643
rect 2631 1637 2635 1638
rect 2703 1642 2707 1643
rect 2703 1637 2707 1638
rect 2767 1642 2771 1643
rect 2767 1637 2771 1638
rect 2871 1642 2875 1643
rect 2871 1637 2875 1638
rect 2895 1642 2899 1643
rect 2895 1637 2899 1638
rect 3023 1642 3027 1643
rect 3023 1637 3027 1638
rect 3031 1642 3035 1643
rect 3031 1637 3035 1638
rect 3143 1642 3147 1643
rect 3143 1637 3147 1638
rect 3191 1642 3195 1643
rect 3191 1637 3195 1638
rect 3255 1642 3259 1643
rect 3255 1637 3259 1638
rect 3351 1642 3355 1643
rect 3351 1637 3355 1638
rect 3375 1642 3379 1643
rect 3375 1637 3379 1638
rect 3487 1642 3491 1643
rect 3487 1637 3491 1638
rect 3575 1642 3579 1643
rect 3575 1637 3579 1638
rect 1823 1633 1827 1634
rect 112 1618 114 1633
rect 136 1628 138 1633
rect 272 1628 274 1633
rect 448 1628 450 1633
rect 632 1628 634 1633
rect 816 1628 818 1633
rect 992 1628 994 1633
rect 1152 1628 1154 1633
rect 1304 1628 1306 1633
rect 1456 1628 1458 1633
rect 1600 1628 1602 1633
rect 1728 1628 1730 1633
rect 134 1627 140 1628
rect 134 1623 135 1627
rect 139 1623 140 1627
rect 134 1622 140 1623
rect 270 1627 276 1628
rect 270 1623 271 1627
rect 275 1623 276 1627
rect 270 1622 276 1623
rect 446 1627 452 1628
rect 446 1623 447 1627
rect 451 1623 452 1627
rect 446 1622 452 1623
rect 630 1627 636 1628
rect 630 1623 631 1627
rect 635 1623 636 1627
rect 630 1622 636 1623
rect 814 1627 820 1628
rect 814 1623 815 1627
rect 819 1623 820 1627
rect 814 1622 820 1623
rect 990 1627 996 1628
rect 990 1623 991 1627
rect 995 1623 996 1627
rect 990 1622 996 1623
rect 1150 1627 1156 1628
rect 1150 1623 1151 1627
rect 1155 1623 1156 1627
rect 1150 1622 1156 1623
rect 1302 1627 1308 1628
rect 1302 1623 1303 1627
rect 1307 1623 1308 1627
rect 1302 1622 1308 1623
rect 1454 1627 1460 1628
rect 1454 1623 1455 1627
rect 1459 1623 1460 1627
rect 1454 1622 1460 1623
rect 1598 1627 1604 1628
rect 1598 1623 1599 1627
rect 1603 1623 1604 1627
rect 1598 1622 1604 1623
rect 1726 1627 1732 1628
rect 1726 1623 1727 1627
rect 1731 1623 1732 1627
rect 1726 1622 1732 1623
rect 1824 1618 1826 1633
rect 110 1617 116 1618
rect 110 1613 111 1617
rect 115 1613 116 1617
rect 110 1612 116 1613
rect 1822 1617 1828 1618
rect 1822 1613 1823 1617
rect 1827 1613 1828 1617
rect 1864 1613 1866 1637
rect 2152 1626 2154 1637
rect 2344 1626 2346 1637
rect 2528 1626 2530 1637
rect 2704 1626 2706 1637
rect 2872 1626 2874 1637
rect 3032 1626 3034 1637
rect 3192 1626 3194 1637
rect 3352 1626 3354 1637
rect 3488 1626 3490 1637
rect 2150 1625 2156 1626
rect 2150 1621 2151 1625
rect 2155 1621 2156 1625
rect 2150 1620 2156 1621
rect 2342 1625 2348 1626
rect 2342 1621 2343 1625
rect 2347 1621 2348 1625
rect 2342 1620 2348 1621
rect 2526 1625 2532 1626
rect 2526 1621 2527 1625
rect 2531 1621 2532 1625
rect 2526 1620 2532 1621
rect 2702 1625 2708 1626
rect 2702 1621 2703 1625
rect 2707 1621 2708 1625
rect 2702 1620 2708 1621
rect 2870 1625 2876 1626
rect 2870 1621 2871 1625
rect 2875 1621 2876 1625
rect 2870 1620 2876 1621
rect 3030 1625 3036 1626
rect 3030 1621 3031 1625
rect 3035 1621 3036 1625
rect 3030 1620 3036 1621
rect 3190 1625 3196 1626
rect 3190 1621 3191 1625
rect 3195 1621 3196 1625
rect 3190 1620 3196 1621
rect 3350 1625 3356 1626
rect 3350 1621 3351 1625
rect 3355 1621 3356 1625
rect 3350 1620 3356 1621
rect 3486 1625 3492 1626
rect 3486 1621 3487 1625
rect 3491 1621 3492 1625
rect 3486 1620 3492 1621
rect 3576 1613 3578 1637
rect 1822 1612 1828 1613
rect 1862 1612 1868 1613
rect 1862 1608 1863 1612
rect 1867 1608 1868 1612
rect 1862 1607 1868 1608
rect 3574 1612 3580 1613
rect 3574 1608 3575 1612
rect 3579 1608 3580 1612
rect 3574 1607 3580 1608
rect 110 1600 116 1601
rect 110 1596 111 1600
rect 115 1596 116 1600
rect 110 1595 116 1596
rect 1822 1600 1828 1601
rect 1822 1596 1823 1600
rect 1827 1596 1828 1600
rect 1822 1595 1828 1596
rect 1862 1595 1868 1596
rect 112 1571 114 1595
rect 142 1587 148 1588
rect 142 1583 143 1587
rect 147 1583 148 1587
rect 142 1582 148 1583
rect 278 1587 284 1588
rect 278 1583 279 1587
rect 283 1583 284 1587
rect 278 1582 284 1583
rect 454 1587 460 1588
rect 454 1583 455 1587
rect 459 1583 460 1587
rect 454 1582 460 1583
rect 638 1587 644 1588
rect 638 1583 639 1587
rect 643 1583 644 1587
rect 638 1582 644 1583
rect 822 1587 828 1588
rect 822 1583 823 1587
rect 827 1583 828 1587
rect 822 1582 828 1583
rect 998 1587 1004 1588
rect 998 1583 999 1587
rect 1003 1583 1004 1587
rect 998 1582 1004 1583
rect 1158 1587 1164 1588
rect 1158 1583 1159 1587
rect 1163 1583 1164 1587
rect 1158 1582 1164 1583
rect 1310 1587 1316 1588
rect 1310 1583 1311 1587
rect 1315 1583 1316 1587
rect 1310 1582 1316 1583
rect 1462 1587 1468 1588
rect 1462 1583 1463 1587
rect 1467 1583 1468 1587
rect 1462 1582 1468 1583
rect 1606 1587 1612 1588
rect 1606 1583 1607 1587
rect 1611 1583 1612 1587
rect 1606 1582 1612 1583
rect 1734 1587 1740 1588
rect 1734 1583 1735 1587
rect 1739 1583 1740 1587
rect 1734 1582 1740 1583
rect 144 1571 146 1582
rect 280 1571 282 1582
rect 456 1571 458 1582
rect 640 1571 642 1582
rect 824 1571 826 1582
rect 1000 1571 1002 1582
rect 1160 1571 1162 1582
rect 1312 1571 1314 1582
rect 1464 1571 1466 1582
rect 1608 1571 1610 1582
rect 1736 1571 1738 1582
rect 1824 1571 1826 1595
rect 1862 1591 1863 1595
rect 1867 1591 1868 1595
rect 1862 1590 1868 1591
rect 3574 1595 3580 1596
rect 3574 1591 3575 1595
rect 3579 1591 3580 1595
rect 3574 1590 3580 1591
rect 1864 1575 1866 1590
rect 2142 1585 2148 1586
rect 2142 1581 2143 1585
rect 2147 1581 2148 1585
rect 2142 1580 2148 1581
rect 2334 1585 2340 1586
rect 2334 1581 2335 1585
rect 2339 1581 2340 1585
rect 2334 1580 2340 1581
rect 2518 1585 2524 1586
rect 2518 1581 2519 1585
rect 2523 1581 2524 1585
rect 2518 1580 2524 1581
rect 2694 1585 2700 1586
rect 2694 1581 2695 1585
rect 2699 1581 2700 1585
rect 2694 1580 2700 1581
rect 2862 1585 2868 1586
rect 2862 1581 2863 1585
rect 2867 1581 2868 1585
rect 2862 1580 2868 1581
rect 3022 1585 3028 1586
rect 3022 1581 3023 1585
rect 3027 1581 3028 1585
rect 3022 1580 3028 1581
rect 3182 1585 3188 1586
rect 3182 1581 3183 1585
rect 3187 1581 3188 1585
rect 3182 1580 3188 1581
rect 3342 1585 3348 1586
rect 3342 1581 3343 1585
rect 3347 1581 3348 1585
rect 3342 1580 3348 1581
rect 3478 1585 3484 1586
rect 3478 1581 3479 1585
rect 3483 1581 3484 1585
rect 3478 1580 3484 1581
rect 2144 1575 2146 1580
rect 2336 1575 2338 1580
rect 2520 1575 2522 1580
rect 2696 1575 2698 1580
rect 2864 1575 2866 1580
rect 3024 1575 3026 1580
rect 3184 1575 3186 1580
rect 3344 1575 3346 1580
rect 3480 1575 3482 1580
rect 3576 1575 3578 1590
rect 1863 1574 1867 1575
rect 111 1570 115 1571
rect 111 1565 115 1566
rect 143 1570 147 1571
rect 143 1565 147 1566
rect 271 1570 275 1571
rect 271 1565 275 1566
rect 279 1570 283 1571
rect 279 1565 283 1566
rect 431 1570 435 1571
rect 431 1565 435 1566
rect 455 1570 459 1571
rect 455 1565 459 1566
rect 599 1570 603 1571
rect 599 1565 603 1566
rect 639 1570 643 1571
rect 639 1565 643 1566
rect 767 1570 771 1571
rect 767 1565 771 1566
rect 823 1570 827 1571
rect 823 1565 827 1566
rect 935 1570 939 1571
rect 935 1565 939 1566
rect 999 1570 1003 1571
rect 999 1565 1003 1566
rect 1103 1570 1107 1571
rect 1103 1565 1107 1566
rect 1159 1570 1163 1571
rect 1159 1565 1163 1566
rect 1263 1570 1267 1571
rect 1263 1565 1267 1566
rect 1311 1570 1315 1571
rect 1311 1565 1315 1566
rect 1423 1570 1427 1571
rect 1423 1565 1427 1566
rect 1463 1570 1467 1571
rect 1463 1565 1467 1566
rect 1591 1570 1595 1571
rect 1591 1565 1595 1566
rect 1607 1570 1611 1571
rect 1607 1565 1611 1566
rect 1735 1570 1739 1571
rect 1735 1565 1739 1566
rect 1823 1570 1827 1571
rect 1863 1569 1867 1570
rect 2087 1574 2091 1575
rect 2087 1569 2091 1570
rect 2143 1574 2147 1575
rect 2143 1569 2147 1570
rect 2279 1574 2283 1575
rect 2279 1569 2283 1570
rect 2335 1574 2339 1575
rect 2335 1569 2339 1570
rect 2455 1574 2459 1575
rect 2455 1569 2459 1570
rect 2519 1574 2523 1575
rect 2519 1569 2523 1570
rect 2623 1574 2627 1575
rect 2623 1569 2627 1570
rect 2695 1574 2699 1575
rect 2695 1569 2699 1570
rect 2791 1574 2795 1575
rect 2791 1569 2795 1570
rect 2863 1574 2867 1575
rect 2863 1569 2867 1570
rect 2951 1574 2955 1575
rect 2951 1569 2955 1570
rect 3023 1574 3027 1575
rect 3023 1569 3027 1570
rect 3111 1574 3115 1575
rect 3111 1569 3115 1570
rect 3183 1574 3187 1575
rect 3183 1569 3187 1570
rect 3271 1574 3275 1575
rect 3271 1569 3275 1570
rect 3343 1574 3347 1575
rect 3343 1569 3347 1570
rect 3431 1574 3435 1575
rect 3431 1569 3435 1570
rect 3479 1574 3483 1575
rect 3479 1569 3483 1570
rect 3575 1574 3579 1575
rect 3575 1569 3579 1570
rect 1823 1565 1827 1566
rect 112 1541 114 1565
rect 144 1554 146 1565
rect 272 1554 274 1565
rect 432 1554 434 1565
rect 600 1554 602 1565
rect 768 1554 770 1565
rect 936 1554 938 1565
rect 1104 1554 1106 1565
rect 1264 1554 1266 1565
rect 1424 1554 1426 1565
rect 1592 1554 1594 1565
rect 1736 1554 1738 1565
rect 142 1553 148 1554
rect 142 1549 143 1553
rect 147 1549 148 1553
rect 142 1548 148 1549
rect 270 1553 276 1554
rect 270 1549 271 1553
rect 275 1549 276 1553
rect 270 1548 276 1549
rect 430 1553 436 1554
rect 430 1549 431 1553
rect 435 1549 436 1553
rect 430 1548 436 1549
rect 598 1553 604 1554
rect 598 1549 599 1553
rect 603 1549 604 1553
rect 598 1548 604 1549
rect 766 1553 772 1554
rect 766 1549 767 1553
rect 771 1549 772 1553
rect 766 1548 772 1549
rect 934 1553 940 1554
rect 934 1549 935 1553
rect 939 1549 940 1553
rect 934 1548 940 1549
rect 1102 1553 1108 1554
rect 1102 1549 1103 1553
rect 1107 1549 1108 1553
rect 1102 1548 1108 1549
rect 1262 1553 1268 1554
rect 1262 1549 1263 1553
rect 1267 1549 1268 1553
rect 1262 1548 1268 1549
rect 1422 1553 1428 1554
rect 1422 1549 1423 1553
rect 1427 1549 1428 1553
rect 1422 1548 1428 1549
rect 1590 1553 1596 1554
rect 1590 1549 1591 1553
rect 1595 1549 1596 1553
rect 1590 1548 1596 1549
rect 1734 1553 1740 1554
rect 1734 1549 1735 1553
rect 1739 1549 1740 1553
rect 1734 1548 1740 1549
rect 1824 1541 1826 1565
rect 1864 1554 1866 1569
rect 2088 1564 2090 1569
rect 2280 1564 2282 1569
rect 2456 1564 2458 1569
rect 2624 1564 2626 1569
rect 2792 1564 2794 1569
rect 2952 1564 2954 1569
rect 3112 1564 3114 1569
rect 3272 1564 3274 1569
rect 3432 1564 3434 1569
rect 2086 1563 2092 1564
rect 2086 1559 2087 1563
rect 2091 1559 2092 1563
rect 2086 1558 2092 1559
rect 2278 1563 2284 1564
rect 2278 1559 2279 1563
rect 2283 1559 2284 1563
rect 2278 1558 2284 1559
rect 2454 1563 2460 1564
rect 2454 1559 2455 1563
rect 2459 1559 2460 1563
rect 2454 1558 2460 1559
rect 2622 1563 2628 1564
rect 2622 1559 2623 1563
rect 2627 1559 2628 1563
rect 2622 1558 2628 1559
rect 2790 1563 2796 1564
rect 2790 1559 2791 1563
rect 2795 1559 2796 1563
rect 2790 1558 2796 1559
rect 2950 1563 2956 1564
rect 2950 1559 2951 1563
rect 2955 1559 2956 1563
rect 2950 1558 2956 1559
rect 3110 1563 3116 1564
rect 3110 1559 3111 1563
rect 3115 1559 3116 1563
rect 3110 1558 3116 1559
rect 3270 1563 3276 1564
rect 3270 1559 3271 1563
rect 3275 1559 3276 1563
rect 3270 1558 3276 1559
rect 3430 1563 3436 1564
rect 3430 1559 3431 1563
rect 3435 1559 3436 1563
rect 3430 1558 3436 1559
rect 3576 1554 3578 1569
rect 1862 1553 1868 1554
rect 1862 1549 1863 1553
rect 1867 1549 1868 1553
rect 1862 1548 1868 1549
rect 3574 1553 3580 1554
rect 3574 1549 3575 1553
rect 3579 1549 3580 1553
rect 3574 1548 3580 1549
rect 110 1540 116 1541
rect 110 1536 111 1540
rect 115 1536 116 1540
rect 110 1535 116 1536
rect 1822 1540 1828 1541
rect 1822 1536 1823 1540
rect 1827 1536 1828 1540
rect 1822 1535 1828 1536
rect 1862 1536 1868 1537
rect 1862 1532 1863 1536
rect 1867 1532 1868 1536
rect 1862 1531 1868 1532
rect 3574 1536 3580 1537
rect 3574 1532 3575 1536
rect 3579 1532 3580 1536
rect 3574 1531 3580 1532
rect 110 1523 116 1524
rect 110 1519 111 1523
rect 115 1519 116 1523
rect 110 1518 116 1519
rect 1822 1523 1828 1524
rect 1822 1519 1823 1523
rect 1827 1519 1828 1523
rect 1822 1518 1828 1519
rect 112 1499 114 1518
rect 134 1513 140 1514
rect 134 1509 135 1513
rect 139 1509 140 1513
rect 134 1508 140 1509
rect 262 1513 268 1514
rect 262 1509 263 1513
rect 267 1509 268 1513
rect 262 1508 268 1509
rect 422 1513 428 1514
rect 422 1509 423 1513
rect 427 1509 428 1513
rect 422 1508 428 1509
rect 590 1513 596 1514
rect 590 1509 591 1513
rect 595 1509 596 1513
rect 590 1508 596 1509
rect 758 1513 764 1514
rect 758 1509 759 1513
rect 763 1509 764 1513
rect 758 1508 764 1509
rect 926 1513 932 1514
rect 926 1509 927 1513
rect 931 1509 932 1513
rect 926 1508 932 1509
rect 1094 1513 1100 1514
rect 1094 1509 1095 1513
rect 1099 1509 1100 1513
rect 1094 1508 1100 1509
rect 1254 1513 1260 1514
rect 1254 1509 1255 1513
rect 1259 1509 1260 1513
rect 1254 1508 1260 1509
rect 1414 1513 1420 1514
rect 1414 1509 1415 1513
rect 1419 1509 1420 1513
rect 1414 1508 1420 1509
rect 1582 1513 1588 1514
rect 1582 1509 1583 1513
rect 1587 1509 1588 1513
rect 1582 1508 1588 1509
rect 1726 1513 1732 1514
rect 1726 1509 1727 1513
rect 1731 1509 1732 1513
rect 1726 1508 1732 1509
rect 136 1499 138 1508
rect 264 1499 266 1508
rect 424 1499 426 1508
rect 592 1499 594 1508
rect 760 1499 762 1508
rect 928 1499 930 1508
rect 1096 1499 1098 1508
rect 1256 1499 1258 1508
rect 1416 1499 1418 1508
rect 1584 1499 1586 1508
rect 1728 1499 1730 1508
rect 1824 1499 1826 1518
rect 1864 1499 1866 1531
rect 2094 1523 2100 1524
rect 2094 1519 2095 1523
rect 2099 1519 2100 1523
rect 2094 1518 2100 1519
rect 2286 1523 2292 1524
rect 2286 1519 2287 1523
rect 2291 1519 2292 1523
rect 2286 1518 2292 1519
rect 2462 1523 2468 1524
rect 2462 1519 2463 1523
rect 2467 1519 2468 1523
rect 2462 1518 2468 1519
rect 2630 1523 2636 1524
rect 2630 1519 2631 1523
rect 2635 1519 2636 1523
rect 2630 1518 2636 1519
rect 2798 1523 2804 1524
rect 2798 1519 2799 1523
rect 2803 1519 2804 1523
rect 2798 1518 2804 1519
rect 2958 1523 2964 1524
rect 2958 1519 2959 1523
rect 2963 1519 2964 1523
rect 2958 1518 2964 1519
rect 3118 1523 3124 1524
rect 3118 1519 3119 1523
rect 3123 1519 3124 1523
rect 3118 1518 3124 1519
rect 3278 1523 3284 1524
rect 3278 1519 3279 1523
rect 3283 1519 3284 1523
rect 3278 1518 3284 1519
rect 3438 1523 3444 1524
rect 3438 1519 3439 1523
rect 3443 1519 3444 1523
rect 3438 1518 3444 1519
rect 2096 1499 2098 1518
rect 2288 1499 2290 1518
rect 2464 1499 2466 1518
rect 2632 1499 2634 1518
rect 2800 1499 2802 1518
rect 2960 1499 2962 1518
rect 3120 1499 3122 1518
rect 3280 1499 3282 1518
rect 3440 1499 3442 1518
rect 3576 1499 3578 1531
rect 111 1498 115 1499
rect 111 1493 115 1494
rect 135 1498 139 1499
rect 135 1493 139 1494
rect 183 1498 187 1499
rect 183 1493 187 1494
rect 263 1498 267 1499
rect 263 1493 267 1494
rect 327 1498 331 1499
rect 327 1493 331 1494
rect 423 1498 427 1499
rect 423 1493 427 1494
rect 471 1498 475 1499
rect 471 1493 475 1494
rect 591 1498 595 1499
rect 591 1493 595 1494
rect 607 1498 611 1499
rect 607 1493 611 1494
rect 743 1498 747 1499
rect 743 1493 747 1494
rect 759 1498 763 1499
rect 759 1493 763 1494
rect 871 1498 875 1499
rect 871 1493 875 1494
rect 927 1498 931 1499
rect 927 1493 931 1494
rect 991 1498 995 1499
rect 991 1493 995 1494
rect 1095 1498 1099 1499
rect 1095 1493 1099 1494
rect 1119 1498 1123 1499
rect 1119 1493 1123 1494
rect 1247 1498 1251 1499
rect 1247 1493 1251 1494
rect 1255 1498 1259 1499
rect 1255 1493 1259 1494
rect 1375 1498 1379 1499
rect 1375 1493 1379 1494
rect 1415 1498 1419 1499
rect 1415 1493 1419 1494
rect 1583 1498 1587 1499
rect 1583 1493 1587 1494
rect 1727 1498 1731 1499
rect 1727 1493 1731 1494
rect 1823 1498 1827 1499
rect 1823 1493 1827 1494
rect 1863 1498 1867 1499
rect 1863 1493 1867 1494
rect 1895 1498 1899 1499
rect 1895 1493 1899 1494
rect 1991 1498 1995 1499
rect 1991 1493 1995 1494
rect 2095 1498 2099 1499
rect 2095 1493 2099 1494
rect 2119 1498 2123 1499
rect 2119 1493 2123 1494
rect 2247 1498 2251 1499
rect 2247 1493 2251 1494
rect 2287 1498 2291 1499
rect 2287 1493 2291 1494
rect 2383 1498 2387 1499
rect 2383 1493 2387 1494
rect 2463 1498 2467 1499
rect 2463 1493 2467 1494
rect 2535 1498 2539 1499
rect 2535 1493 2539 1494
rect 2631 1498 2635 1499
rect 2631 1493 2635 1494
rect 2703 1498 2707 1499
rect 2703 1493 2707 1494
rect 2799 1498 2803 1499
rect 2799 1493 2803 1494
rect 2887 1498 2891 1499
rect 2887 1493 2891 1494
rect 2959 1498 2963 1499
rect 2959 1493 2963 1494
rect 3087 1498 3091 1499
rect 3087 1493 3091 1494
rect 3119 1498 3123 1499
rect 3119 1493 3123 1494
rect 3279 1498 3283 1499
rect 3279 1493 3283 1494
rect 3295 1498 3299 1499
rect 3295 1493 3299 1494
rect 3439 1498 3443 1499
rect 3439 1493 3443 1494
rect 3487 1498 3491 1499
rect 3487 1493 3491 1494
rect 3575 1498 3579 1499
rect 3575 1493 3579 1494
rect 112 1478 114 1493
rect 184 1488 186 1493
rect 328 1488 330 1493
rect 472 1488 474 1493
rect 608 1488 610 1493
rect 744 1488 746 1493
rect 872 1488 874 1493
rect 992 1488 994 1493
rect 1120 1488 1122 1493
rect 1248 1488 1250 1493
rect 1376 1488 1378 1493
rect 182 1487 188 1488
rect 182 1483 183 1487
rect 187 1483 188 1487
rect 182 1482 188 1483
rect 326 1487 332 1488
rect 326 1483 327 1487
rect 331 1483 332 1487
rect 326 1482 332 1483
rect 470 1487 476 1488
rect 470 1483 471 1487
rect 475 1483 476 1487
rect 470 1482 476 1483
rect 606 1487 612 1488
rect 606 1483 607 1487
rect 611 1483 612 1487
rect 606 1482 612 1483
rect 742 1487 748 1488
rect 742 1483 743 1487
rect 747 1483 748 1487
rect 742 1482 748 1483
rect 870 1487 876 1488
rect 870 1483 871 1487
rect 875 1483 876 1487
rect 870 1482 876 1483
rect 990 1487 996 1488
rect 990 1483 991 1487
rect 995 1483 996 1487
rect 990 1482 996 1483
rect 1118 1487 1124 1488
rect 1118 1483 1119 1487
rect 1123 1483 1124 1487
rect 1118 1482 1124 1483
rect 1246 1487 1252 1488
rect 1246 1483 1247 1487
rect 1251 1483 1252 1487
rect 1246 1482 1252 1483
rect 1374 1487 1380 1488
rect 1374 1483 1375 1487
rect 1379 1483 1380 1487
rect 1374 1482 1380 1483
rect 1824 1478 1826 1493
rect 110 1477 116 1478
rect 110 1473 111 1477
rect 115 1473 116 1477
rect 110 1472 116 1473
rect 1822 1477 1828 1478
rect 1822 1473 1823 1477
rect 1827 1473 1828 1477
rect 1822 1472 1828 1473
rect 1864 1469 1866 1493
rect 1896 1482 1898 1493
rect 1992 1482 1994 1493
rect 2120 1482 2122 1493
rect 2248 1482 2250 1493
rect 2384 1482 2386 1493
rect 2536 1482 2538 1493
rect 2704 1482 2706 1493
rect 2888 1482 2890 1493
rect 3088 1482 3090 1493
rect 3296 1482 3298 1493
rect 3488 1482 3490 1493
rect 1894 1481 1900 1482
rect 1894 1477 1895 1481
rect 1899 1477 1900 1481
rect 1894 1476 1900 1477
rect 1990 1481 1996 1482
rect 1990 1477 1991 1481
rect 1995 1477 1996 1481
rect 1990 1476 1996 1477
rect 2118 1481 2124 1482
rect 2118 1477 2119 1481
rect 2123 1477 2124 1481
rect 2118 1476 2124 1477
rect 2246 1481 2252 1482
rect 2246 1477 2247 1481
rect 2251 1477 2252 1481
rect 2246 1476 2252 1477
rect 2382 1481 2388 1482
rect 2382 1477 2383 1481
rect 2387 1477 2388 1481
rect 2382 1476 2388 1477
rect 2534 1481 2540 1482
rect 2534 1477 2535 1481
rect 2539 1477 2540 1481
rect 2534 1476 2540 1477
rect 2702 1481 2708 1482
rect 2702 1477 2703 1481
rect 2707 1477 2708 1481
rect 2702 1476 2708 1477
rect 2886 1481 2892 1482
rect 2886 1477 2887 1481
rect 2891 1477 2892 1481
rect 2886 1476 2892 1477
rect 3086 1481 3092 1482
rect 3086 1477 3087 1481
rect 3091 1477 3092 1481
rect 3086 1476 3092 1477
rect 3294 1481 3300 1482
rect 3294 1477 3295 1481
rect 3299 1477 3300 1481
rect 3294 1476 3300 1477
rect 3486 1481 3492 1482
rect 3486 1477 3487 1481
rect 3491 1477 3492 1481
rect 3486 1476 3492 1477
rect 3576 1469 3578 1493
rect 1862 1468 1868 1469
rect 1862 1464 1863 1468
rect 1867 1464 1868 1468
rect 1862 1463 1868 1464
rect 3574 1468 3580 1469
rect 3574 1464 3575 1468
rect 3579 1464 3580 1468
rect 3574 1463 3580 1464
rect 110 1460 116 1461
rect 110 1456 111 1460
rect 115 1456 116 1460
rect 110 1455 116 1456
rect 1822 1460 1828 1461
rect 1822 1456 1823 1460
rect 1827 1456 1828 1460
rect 1822 1455 1828 1456
rect 112 1423 114 1455
rect 190 1447 196 1448
rect 190 1443 191 1447
rect 195 1443 196 1447
rect 190 1442 196 1443
rect 334 1447 340 1448
rect 334 1443 335 1447
rect 339 1443 340 1447
rect 334 1442 340 1443
rect 478 1447 484 1448
rect 478 1443 479 1447
rect 483 1443 484 1447
rect 478 1442 484 1443
rect 614 1447 620 1448
rect 614 1443 615 1447
rect 619 1443 620 1447
rect 614 1442 620 1443
rect 750 1447 756 1448
rect 750 1443 751 1447
rect 755 1443 756 1447
rect 750 1442 756 1443
rect 878 1447 884 1448
rect 878 1443 879 1447
rect 883 1443 884 1447
rect 878 1442 884 1443
rect 998 1447 1004 1448
rect 998 1443 999 1447
rect 1003 1443 1004 1447
rect 998 1442 1004 1443
rect 1126 1447 1132 1448
rect 1126 1443 1127 1447
rect 1131 1443 1132 1447
rect 1126 1442 1132 1443
rect 1254 1447 1260 1448
rect 1254 1443 1255 1447
rect 1259 1443 1260 1447
rect 1254 1442 1260 1443
rect 1382 1447 1388 1448
rect 1382 1443 1383 1447
rect 1387 1443 1388 1447
rect 1382 1442 1388 1443
rect 192 1423 194 1442
rect 336 1423 338 1442
rect 480 1423 482 1442
rect 616 1423 618 1442
rect 752 1423 754 1442
rect 880 1423 882 1442
rect 1000 1423 1002 1442
rect 1128 1423 1130 1442
rect 1256 1423 1258 1442
rect 1384 1423 1386 1442
rect 1824 1423 1826 1455
rect 1862 1451 1868 1452
rect 1862 1447 1863 1451
rect 1867 1447 1868 1451
rect 1862 1446 1868 1447
rect 3574 1451 3580 1452
rect 3574 1447 3575 1451
rect 3579 1447 3580 1451
rect 3574 1446 3580 1447
rect 1864 1427 1866 1446
rect 1886 1441 1892 1442
rect 1886 1437 1887 1441
rect 1891 1437 1892 1441
rect 1886 1436 1892 1437
rect 1982 1441 1988 1442
rect 1982 1437 1983 1441
rect 1987 1437 1988 1441
rect 1982 1436 1988 1437
rect 2110 1441 2116 1442
rect 2110 1437 2111 1441
rect 2115 1437 2116 1441
rect 2110 1436 2116 1437
rect 2238 1441 2244 1442
rect 2238 1437 2239 1441
rect 2243 1437 2244 1441
rect 2238 1436 2244 1437
rect 2374 1441 2380 1442
rect 2374 1437 2375 1441
rect 2379 1437 2380 1441
rect 2374 1436 2380 1437
rect 2526 1441 2532 1442
rect 2526 1437 2527 1441
rect 2531 1437 2532 1441
rect 2526 1436 2532 1437
rect 2694 1441 2700 1442
rect 2694 1437 2695 1441
rect 2699 1437 2700 1441
rect 2694 1436 2700 1437
rect 2878 1441 2884 1442
rect 2878 1437 2879 1441
rect 2883 1437 2884 1441
rect 2878 1436 2884 1437
rect 3078 1441 3084 1442
rect 3078 1437 3079 1441
rect 3083 1437 3084 1441
rect 3078 1436 3084 1437
rect 3286 1441 3292 1442
rect 3286 1437 3287 1441
rect 3291 1437 3292 1441
rect 3286 1436 3292 1437
rect 3478 1441 3484 1442
rect 3478 1437 3479 1441
rect 3483 1437 3484 1441
rect 3478 1436 3484 1437
rect 1888 1427 1890 1436
rect 1984 1427 1986 1436
rect 2112 1427 2114 1436
rect 2240 1427 2242 1436
rect 2376 1427 2378 1436
rect 2528 1427 2530 1436
rect 2696 1427 2698 1436
rect 2880 1427 2882 1436
rect 3080 1427 3082 1436
rect 3288 1427 3290 1436
rect 3480 1427 3482 1436
rect 3576 1427 3578 1446
rect 1863 1426 1867 1427
rect 111 1422 115 1423
rect 111 1417 115 1418
rect 191 1422 195 1423
rect 191 1417 195 1418
rect 199 1422 203 1423
rect 199 1417 203 1418
rect 335 1422 339 1423
rect 335 1417 339 1418
rect 463 1422 467 1423
rect 463 1417 467 1418
rect 479 1422 483 1423
rect 479 1417 483 1418
rect 583 1422 587 1423
rect 583 1417 587 1418
rect 615 1422 619 1423
rect 615 1417 619 1418
rect 703 1422 707 1423
rect 703 1417 707 1418
rect 751 1422 755 1423
rect 751 1417 755 1418
rect 815 1422 819 1423
rect 815 1417 819 1418
rect 879 1422 883 1423
rect 879 1417 883 1418
rect 919 1422 923 1423
rect 919 1417 923 1418
rect 999 1422 1003 1423
rect 999 1417 1003 1418
rect 1015 1422 1019 1423
rect 1015 1417 1019 1418
rect 1119 1422 1123 1423
rect 1119 1417 1123 1418
rect 1127 1422 1131 1423
rect 1127 1417 1131 1418
rect 1223 1422 1227 1423
rect 1223 1417 1227 1418
rect 1255 1422 1259 1423
rect 1255 1417 1259 1418
rect 1327 1422 1331 1423
rect 1327 1417 1331 1418
rect 1383 1422 1387 1423
rect 1383 1417 1387 1418
rect 1823 1422 1827 1423
rect 1863 1421 1867 1422
rect 1887 1426 1891 1427
rect 1887 1421 1891 1422
rect 1975 1426 1979 1427
rect 1975 1421 1979 1422
rect 1983 1426 1987 1427
rect 1983 1421 1987 1422
rect 2071 1426 2075 1427
rect 2071 1421 2075 1422
rect 2111 1426 2115 1427
rect 2111 1421 2115 1422
rect 2183 1426 2187 1427
rect 2183 1421 2187 1422
rect 2239 1426 2243 1427
rect 2239 1421 2243 1422
rect 2303 1426 2307 1427
rect 2303 1421 2307 1422
rect 2375 1426 2379 1427
rect 2375 1421 2379 1422
rect 2439 1426 2443 1427
rect 2439 1421 2443 1422
rect 2527 1426 2531 1427
rect 2527 1421 2531 1422
rect 2607 1426 2611 1427
rect 2607 1421 2611 1422
rect 2695 1426 2699 1427
rect 2695 1421 2699 1422
rect 2807 1426 2811 1427
rect 2807 1421 2811 1422
rect 2879 1426 2883 1427
rect 2879 1421 2883 1422
rect 3031 1426 3035 1427
rect 3031 1421 3035 1422
rect 3079 1426 3083 1427
rect 3079 1421 3083 1422
rect 3263 1426 3267 1427
rect 3263 1421 3267 1422
rect 3287 1426 3291 1427
rect 3287 1421 3291 1422
rect 3479 1426 3483 1427
rect 3479 1421 3483 1422
rect 3575 1426 3579 1427
rect 3575 1421 3579 1422
rect 1823 1417 1827 1418
rect 112 1393 114 1417
rect 200 1406 202 1417
rect 336 1406 338 1417
rect 464 1406 466 1417
rect 584 1406 586 1417
rect 704 1406 706 1417
rect 816 1406 818 1417
rect 920 1406 922 1417
rect 1016 1406 1018 1417
rect 1120 1406 1122 1417
rect 1224 1406 1226 1417
rect 1328 1406 1330 1417
rect 198 1405 204 1406
rect 198 1401 199 1405
rect 203 1401 204 1405
rect 198 1400 204 1401
rect 334 1405 340 1406
rect 334 1401 335 1405
rect 339 1401 340 1405
rect 334 1400 340 1401
rect 462 1405 468 1406
rect 462 1401 463 1405
rect 467 1401 468 1405
rect 462 1400 468 1401
rect 582 1405 588 1406
rect 582 1401 583 1405
rect 587 1401 588 1405
rect 582 1400 588 1401
rect 702 1405 708 1406
rect 702 1401 703 1405
rect 707 1401 708 1405
rect 702 1400 708 1401
rect 814 1405 820 1406
rect 814 1401 815 1405
rect 819 1401 820 1405
rect 814 1400 820 1401
rect 918 1405 924 1406
rect 918 1401 919 1405
rect 923 1401 924 1405
rect 918 1400 924 1401
rect 1014 1405 1020 1406
rect 1014 1401 1015 1405
rect 1019 1401 1020 1405
rect 1014 1400 1020 1401
rect 1118 1405 1124 1406
rect 1118 1401 1119 1405
rect 1123 1401 1124 1405
rect 1118 1400 1124 1401
rect 1222 1405 1228 1406
rect 1222 1401 1223 1405
rect 1227 1401 1228 1405
rect 1222 1400 1228 1401
rect 1326 1405 1332 1406
rect 1326 1401 1327 1405
rect 1331 1401 1332 1405
rect 1326 1400 1332 1401
rect 1824 1393 1826 1417
rect 1864 1406 1866 1421
rect 1888 1416 1890 1421
rect 1976 1416 1978 1421
rect 2072 1416 2074 1421
rect 2184 1416 2186 1421
rect 2304 1416 2306 1421
rect 2440 1416 2442 1421
rect 2608 1416 2610 1421
rect 2808 1416 2810 1421
rect 3032 1416 3034 1421
rect 3264 1416 3266 1421
rect 3480 1416 3482 1421
rect 1886 1415 1892 1416
rect 1886 1411 1887 1415
rect 1891 1411 1892 1415
rect 1886 1410 1892 1411
rect 1974 1415 1980 1416
rect 1974 1411 1975 1415
rect 1979 1411 1980 1415
rect 1974 1410 1980 1411
rect 2070 1415 2076 1416
rect 2070 1411 2071 1415
rect 2075 1411 2076 1415
rect 2070 1410 2076 1411
rect 2182 1415 2188 1416
rect 2182 1411 2183 1415
rect 2187 1411 2188 1415
rect 2182 1410 2188 1411
rect 2302 1415 2308 1416
rect 2302 1411 2303 1415
rect 2307 1411 2308 1415
rect 2302 1410 2308 1411
rect 2438 1415 2444 1416
rect 2438 1411 2439 1415
rect 2443 1411 2444 1415
rect 2438 1410 2444 1411
rect 2606 1415 2612 1416
rect 2606 1411 2607 1415
rect 2611 1411 2612 1415
rect 2606 1410 2612 1411
rect 2806 1415 2812 1416
rect 2806 1411 2807 1415
rect 2811 1411 2812 1415
rect 2806 1410 2812 1411
rect 3030 1415 3036 1416
rect 3030 1411 3031 1415
rect 3035 1411 3036 1415
rect 3030 1410 3036 1411
rect 3262 1415 3268 1416
rect 3262 1411 3263 1415
rect 3267 1411 3268 1415
rect 3262 1410 3268 1411
rect 3478 1415 3484 1416
rect 3478 1411 3479 1415
rect 3483 1411 3484 1415
rect 3478 1410 3484 1411
rect 3576 1406 3578 1421
rect 1862 1405 1868 1406
rect 1862 1401 1863 1405
rect 1867 1401 1868 1405
rect 1862 1400 1868 1401
rect 3574 1405 3580 1406
rect 3574 1401 3575 1405
rect 3579 1401 3580 1405
rect 3574 1400 3580 1401
rect 110 1392 116 1393
rect 110 1388 111 1392
rect 115 1388 116 1392
rect 110 1387 116 1388
rect 1822 1392 1828 1393
rect 1822 1388 1823 1392
rect 1827 1388 1828 1392
rect 1822 1387 1828 1388
rect 1862 1388 1868 1389
rect 1862 1384 1863 1388
rect 1867 1384 1868 1388
rect 1862 1383 1868 1384
rect 3574 1388 3580 1389
rect 3574 1384 3575 1388
rect 3579 1384 3580 1388
rect 3574 1383 3580 1384
rect 110 1375 116 1376
rect 110 1371 111 1375
rect 115 1371 116 1375
rect 110 1370 116 1371
rect 1822 1375 1828 1376
rect 1822 1371 1823 1375
rect 1827 1371 1828 1375
rect 1822 1370 1828 1371
rect 112 1351 114 1370
rect 190 1365 196 1366
rect 190 1361 191 1365
rect 195 1361 196 1365
rect 190 1360 196 1361
rect 326 1365 332 1366
rect 326 1361 327 1365
rect 331 1361 332 1365
rect 326 1360 332 1361
rect 454 1365 460 1366
rect 454 1361 455 1365
rect 459 1361 460 1365
rect 454 1360 460 1361
rect 574 1365 580 1366
rect 574 1361 575 1365
rect 579 1361 580 1365
rect 574 1360 580 1361
rect 694 1365 700 1366
rect 694 1361 695 1365
rect 699 1361 700 1365
rect 694 1360 700 1361
rect 806 1365 812 1366
rect 806 1361 807 1365
rect 811 1361 812 1365
rect 806 1360 812 1361
rect 910 1365 916 1366
rect 910 1361 911 1365
rect 915 1361 916 1365
rect 910 1360 916 1361
rect 1006 1365 1012 1366
rect 1006 1361 1007 1365
rect 1011 1361 1012 1365
rect 1006 1360 1012 1361
rect 1110 1365 1116 1366
rect 1110 1361 1111 1365
rect 1115 1361 1116 1365
rect 1110 1360 1116 1361
rect 1214 1365 1220 1366
rect 1214 1361 1215 1365
rect 1219 1361 1220 1365
rect 1214 1360 1220 1361
rect 1318 1365 1324 1366
rect 1318 1361 1319 1365
rect 1323 1361 1324 1365
rect 1318 1360 1324 1361
rect 192 1351 194 1360
rect 328 1351 330 1360
rect 456 1351 458 1360
rect 576 1351 578 1360
rect 696 1351 698 1360
rect 808 1351 810 1360
rect 912 1351 914 1360
rect 1008 1351 1010 1360
rect 1112 1351 1114 1360
rect 1216 1351 1218 1360
rect 1320 1351 1322 1360
rect 1824 1351 1826 1370
rect 1864 1355 1866 1383
rect 1894 1375 1900 1376
rect 1894 1371 1895 1375
rect 1899 1371 1900 1375
rect 1894 1370 1900 1371
rect 1982 1375 1988 1376
rect 1982 1371 1983 1375
rect 1987 1371 1988 1375
rect 1982 1370 1988 1371
rect 2078 1375 2084 1376
rect 2078 1371 2079 1375
rect 2083 1371 2084 1375
rect 2078 1370 2084 1371
rect 2190 1375 2196 1376
rect 2190 1371 2191 1375
rect 2195 1371 2196 1375
rect 2190 1370 2196 1371
rect 2310 1375 2316 1376
rect 2310 1371 2311 1375
rect 2315 1371 2316 1375
rect 2310 1370 2316 1371
rect 2446 1375 2452 1376
rect 2446 1371 2447 1375
rect 2451 1371 2452 1375
rect 2446 1370 2452 1371
rect 2614 1375 2620 1376
rect 2614 1371 2615 1375
rect 2619 1371 2620 1375
rect 2614 1370 2620 1371
rect 2814 1375 2820 1376
rect 2814 1371 2815 1375
rect 2819 1371 2820 1375
rect 2814 1370 2820 1371
rect 3038 1375 3044 1376
rect 3038 1371 3039 1375
rect 3043 1371 3044 1375
rect 3038 1370 3044 1371
rect 3270 1375 3276 1376
rect 3270 1371 3271 1375
rect 3275 1371 3276 1375
rect 3270 1370 3276 1371
rect 3486 1375 3492 1376
rect 3486 1371 3487 1375
rect 3491 1371 3492 1375
rect 3486 1370 3492 1371
rect 1896 1355 1898 1370
rect 1984 1355 1986 1370
rect 2080 1355 2082 1370
rect 2192 1355 2194 1370
rect 2312 1355 2314 1370
rect 2448 1355 2450 1370
rect 2616 1355 2618 1370
rect 2816 1355 2818 1370
rect 3040 1355 3042 1370
rect 3272 1355 3274 1370
rect 3488 1355 3490 1370
rect 3576 1355 3578 1383
rect 1863 1354 1867 1355
rect 111 1350 115 1351
rect 111 1345 115 1346
rect 191 1350 195 1351
rect 191 1345 195 1346
rect 231 1350 235 1351
rect 231 1345 235 1346
rect 327 1350 331 1351
rect 327 1345 331 1346
rect 383 1350 387 1351
rect 383 1345 387 1346
rect 455 1350 459 1351
rect 455 1345 459 1346
rect 543 1350 547 1351
rect 543 1345 547 1346
rect 575 1350 579 1351
rect 575 1345 579 1346
rect 695 1350 699 1351
rect 695 1345 699 1346
rect 703 1350 707 1351
rect 703 1345 707 1346
rect 807 1350 811 1351
rect 807 1345 811 1346
rect 871 1350 875 1351
rect 871 1345 875 1346
rect 911 1350 915 1351
rect 911 1345 915 1346
rect 1007 1350 1011 1351
rect 1007 1345 1011 1346
rect 1039 1350 1043 1351
rect 1039 1345 1043 1346
rect 1111 1350 1115 1351
rect 1111 1345 1115 1346
rect 1207 1350 1211 1351
rect 1207 1345 1211 1346
rect 1215 1350 1219 1351
rect 1215 1345 1219 1346
rect 1319 1350 1323 1351
rect 1319 1345 1323 1346
rect 1375 1350 1379 1351
rect 1375 1345 1379 1346
rect 1823 1350 1827 1351
rect 1863 1349 1867 1350
rect 1895 1354 1899 1355
rect 1895 1349 1899 1350
rect 1983 1354 1987 1355
rect 1983 1349 1987 1350
rect 2079 1354 2083 1355
rect 2079 1349 2083 1350
rect 2103 1354 2107 1355
rect 2103 1349 2107 1350
rect 2191 1354 2195 1355
rect 2191 1349 2195 1350
rect 2223 1354 2227 1355
rect 2223 1349 2227 1350
rect 2311 1354 2315 1355
rect 2311 1349 2315 1350
rect 2359 1354 2363 1355
rect 2359 1349 2363 1350
rect 2447 1354 2451 1355
rect 2447 1349 2451 1350
rect 2511 1354 2515 1355
rect 2511 1349 2515 1350
rect 2615 1354 2619 1355
rect 2615 1349 2619 1350
rect 2687 1354 2691 1355
rect 2687 1349 2691 1350
rect 2815 1354 2819 1355
rect 2815 1349 2819 1350
rect 2871 1354 2875 1355
rect 2871 1349 2875 1350
rect 3039 1354 3043 1355
rect 3039 1349 3043 1350
rect 3071 1354 3075 1355
rect 3071 1349 3075 1350
rect 3271 1354 3275 1355
rect 3271 1349 3275 1350
rect 3279 1354 3283 1355
rect 3279 1349 3283 1350
rect 3487 1354 3491 1355
rect 3487 1349 3491 1350
rect 3575 1354 3579 1355
rect 3575 1349 3579 1350
rect 1823 1345 1827 1346
rect 112 1330 114 1345
rect 232 1340 234 1345
rect 384 1340 386 1345
rect 544 1340 546 1345
rect 704 1340 706 1345
rect 872 1340 874 1345
rect 1040 1340 1042 1345
rect 1208 1340 1210 1345
rect 1376 1340 1378 1345
rect 230 1339 236 1340
rect 230 1335 231 1339
rect 235 1335 236 1339
rect 230 1334 236 1335
rect 382 1339 388 1340
rect 382 1335 383 1339
rect 387 1335 388 1339
rect 382 1334 388 1335
rect 542 1339 548 1340
rect 542 1335 543 1339
rect 547 1335 548 1339
rect 542 1334 548 1335
rect 702 1339 708 1340
rect 702 1335 703 1339
rect 707 1335 708 1339
rect 702 1334 708 1335
rect 870 1339 876 1340
rect 870 1335 871 1339
rect 875 1335 876 1339
rect 870 1334 876 1335
rect 1038 1339 1044 1340
rect 1038 1335 1039 1339
rect 1043 1335 1044 1339
rect 1038 1334 1044 1335
rect 1206 1339 1212 1340
rect 1206 1335 1207 1339
rect 1211 1335 1212 1339
rect 1206 1334 1212 1335
rect 1374 1339 1380 1340
rect 1374 1335 1375 1339
rect 1379 1335 1380 1339
rect 1374 1334 1380 1335
rect 1824 1330 1826 1345
rect 110 1329 116 1330
rect 110 1325 111 1329
rect 115 1325 116 1329
rect 110 1324 116 1325
rect 1822 1329 1828 1330
rect 1822 1325 1823 1329
rect 1827 1325 1828 1329
rect 1864 1325 1866 1349
rect 1896 1338 1898 1349
rect 1984 1338 1986 1349
rect 2104 1338 2106 1349
rect 2224 1338 2226 1349
rect 2360 1338 2362 1349
rect 2512 1338 2514 1349
rect 2688 1338 2690 1349
rect 2872 1338 2874 1349
rect 3072 1338 3074 1349
rect 3280 1338 3282 1349
rect 3488 1338 3490 1349
rect 1894 1337 1900 1338
rect 1894 1333 1895 1337
rect 1899 1333 1900 1337
rect 1894 1332 1900 1333
rect 1982 1337 1988 1338
rect 1982 1333 1983 1337
rect 1987 1333 1988 1337
rect 1982 1332 1988 1333
rect 2102 1337 2108 1338
rect 2102 1333 2103 1337
rect 2107 1333 2108 1337
rect 2102 1332 2108 1333
rect 2222 1337 2228 1338
rect 2222 1333 2223 1337
rect 2227 1333 2228 1337
rect 2222 1332 2228 1333
rect 2358 1337 2364 1338
rect 2358 1333 2359 1337
rect 2363 1333 2364 1337
rect 2358 1332 2364 1333
rect 2510 1337 2516 1338
rect 2510 1333 2511 1337
rect 2515 1333 2516 1337
rect 2510 1332 2516 1333
rect 2686 1337 2692 1338
rect 2686 1333 2687 1337
rect 2691 1333 2692 1337
rect 2686 1332 2692 1333
rect 2870 1337 2876 1338
rect 2870 1333 2871 1337
rect 2875 1333 2876 1337
rect 2870 1332 2876 1333
rect 3070 1337 3076 1338
rect 3070 1333 3071 1337
rect 3075 1333 3076 1337
rect 3070 1332 3076 1333
rect 3278 1337 3284 1338
rect 3278 1333 3279 1337
rect 3283 1333 3284 1337
rect 3278 1332 3284 1333
rect 3486 1337 3492 1338
rect 3486 1333 3487 1337
rect 3491 1333 3492 1337
rect 3486 1332 3492 1333
rect 3576 1325 3578 1349
rect 1822 1324 1828 1325
rect 1862 1324 1868 1325
rect 1862 1320 1863 1324
rect 1867 1320 1868 1324
rect 1862 1319 1868 1320
rect 3574 1324 3580 1325
rect 3574 1320 3575 1324
rect 3579 1320 3580 1324
rect 3574 1319 3580 1320
rect 110 1312 116 1313
rect 110 1308 111 1312
rect 115 1308 116 1312
rect 110 1307 116 1308
rect 1822 1312 1828 1313
rect 1822 1308 1823 1312
rect 1827 1308 1828 1312
rect 1822 1307 1828 1308
rect 1862 1307 1868 1308
rect 112 1283 114 1307
rect 238 1299 244 1300
rect 238 1295 239 1299
rect 243 1295 244 1299
rect 238 1294 244 1295
rect 390 1299 396 1300
rect 390 1295 391 1299
rect 395 1295 396 1299
rect 390 1294 396 1295
rect 550 1299 556 1300
rect 550 1295 551 1299
rect 555 1295 556 1299
rect 550 1294 556 1295
rect 710 1299 716 1300
rect 710 1295 711 1299
rect 715 1295 716 1299
rect 710 1294 716 1295
rect 878 1299 884 1300
rect 878 1295 879 1299
rect 883 1295 884 1299
rect 878 1294 884 1295
rect 1046 1299 1052 1300
rect 1046 1295 1047 1299
rect 1051 1295 1052 1299
rect 1046 1294 1052 1295
rect 1214 1299 1220 1300
rect 1214 1295 1215 1299
rect 1219 1295 1220 1299
rect 1214 1294 1220 1295
rect 1382 1299 1388 1300
rect 1382 1295 1383 1299
rect 1387 1295 1388 1299
rect 1382 1294 1388 1295
rect 240 1283 242 1294
rect 392 1283 394 1294
rect 552 1283 554 1294
rect 712 1283 714 1294
rect 880 1283 882 1294
rect 1048 1283 1050 1294
rect 1216 1283 1218 1294
rect 1384 1283 1386 1294
rect 1824 1283 1826 1307
rect 1862 1303 1863 1307
rect 1867 1303 1868 1307
rect 1862 1302 1868 1303
rect 3574 1307 3580 1308
rect 3574 1303 3575 1307
rect 3579 1303 3580 1307
rect 3574 1302 3580 1303
rect 111 1282 115 1283
rect 111 1277 115 1278
rect 215 1282 219 1283
rect 215 1277 219 1278
rect 239 1282 243 1283
rect 239 1277 243 1278
rect 359 1282 363 1283
rect 359 1277 363 1278
rect 391 1282 395 1283
rect 391 1277 395 1278
rect 519 1282 523 1283
rect 519 1277 523 1278
rect 551 1282 555 1283
rect 551 1277 555 1278
rect 679 1282 683 1283
rect 679 1277 683 1278
rect 711 1282 715 1283
rect 711 1277 715 1278
rect 839 1282 843 1283
rect 839 1277 843 1278
rect 879 1282 883 1283
rect 879 1277 883 1278
rect 999 1282 1003 1283
rect 999 1277 1003 1278
rect 1047 1282 1051 1283
rect 1047 1277 1051 1278
rect 1151 1282 1155 1283
rect 1151 1277 1155 1278
rect 1215 1282 1219 1283
rect 1215 1277 1219 1278
rect 1295 1282 1299 1283
rect 1295 1277 1299 1278
rect 1383 1282 1387 1283
rect 1383 1277 1387 1278
rect 1439 1282 1443 1283
rect 1439 1277 1443 1278
rect 1591 1282 1595 1283
rect 1591 1277 1595 1278
rect 1823 1282 1827 1283
rect 1823 1277 1827 1278
rect 112 1253 114 1277
rect 216 1266 218 1277
rect 360 1266 362 1277
rect 520 1266 522 1277
rect 680 1266 682 1277
rect 840 1266 842 1277
rect 1000 1266 1002 1277
rect 1152 1266 1154 1277
rect 1296 1266 1298 1277
rect 1440 1266 1442 1277
rect 1592 1266 1594 1277
rect 214 1265 220 1266
rect 214 1261 215 1265
rect 219 1261 220 1265
rect 214 1260 220 1261
rect 358 1265 364 1266
rect 358 1261 359 1265
rect 363 1261 364 1265
rect 358 1260 364 1261
rect 518 1265 524 1266
rect 518 1261 519 1265
rect 523 1261 524 1265
rect 518 1260 524 1261
rect 678 1265 684 1266
rect 678 1261 679 1265
rect 683 1261 684 1265
rect 678 1260 684 1261
rect 838 1265 844 1266
rect 838 1261 839 1265
rect 843 1261 844 1265
rect 838 1260 844 1261
rect 998 1265 1004 1266
rect 998 1261 999 1265
rect 1003 1261 1004 1265
rect 998 1260 1004 1261
rect 1150 1265 1156 1266
rect 1150 1261 1151 1265
rect 1155 1261 1156 1265
rect 1150 1260 1156 1261
rect 1294 1265 1300 1266
rect 1294 1261 1295 1265
rect 1299 1261 1300 1265
rect 1294 1260 1300 1261
rect 1438 1265 1444 1266
rect 1438 1261 1439 1265
rect 1443 1261 1444 1265
rect 1438 1260 1444 1261
rect 1590 1265 1596 1266
rect 1590 1261 1591 1265
rect 1595 1261 1596 1265
rect 1590 1260 1596 1261
rect 1824 1253 1826 1277
rect 1864 1275 1866 1302
rect 1886 1297 1892 1298
rect 1886 1293 1887 1297
rect 1891 1293 1892 1297
rect 1886 1292 1892 1293
rect 1974 1297 1980 1298
rect 1974 1293 1975 1297
rect 1979 1293 1980 1297
rect 1974 1292 1980 1293
rect 2094 1297 2100 1298
rect 2094 1293 2095 1297
rect 2099 1293 2100 1297
rect 2094 1292 2100 1293
rect 2214 1297 2220 1298
rect 2214 1293 2215 1297
rect 2219 1293 2220 1297
rect 2214 1292 2220 1293
rect 2350 1297 2356 1298
rect 2350 1293 2351 1297
rect 2355 1293 2356 1297
rect 2350 1292 2356 1293
rect 2502 1297 2508 1298
rect 2502 1293 2503 1297
rect 2507 1293 2508 1297
rect 2502 1292 2508 1293
rect 2678 1297 2684 1298
rect 2678 1293 2679 1297
rect 2683 1293 2684 1297
rect 2678 1292 2684 1293
rect 2862 1297 2868 1298
rect 2862 1293 2863 1297
rect 2867 1293 2868 1297
rect 2862 1292 2868 1293
rect 3062 1297 3068 1298
rect 3062 1293 3063 1297
rect 3067 1293 3068 1297
rect 3062 1292 3068 1293
rect 3270 1297 3276 1298
rect 3270 1293 3271 1297
rect 3275 1293 3276 1297
rect 3270 1292 3276 1293
rect 3478 1297 3484 1298
rect 3478 1293 3479 1297
rect 3483 1293 3484 1297
rect 3478 1292 3484 1293
rect 1888 1275 1890 1292
rect 1976 1275 1978 1292
rect 2096 1275 2098 1292
rect 2216 1275 2218 1292
rect 2352 1275 2354 1292
rect 2504 1275 2506 1292
rect 2680 1275 2682 1292
rect 2864 1275 2866 1292
rect 3064 1275 3066 1292
rect 3272 1275 3274 1292
rect 3480 1275 3482 1292
rect 3576 1275 3578 1302
rect 1863 1274 1867 1275
rect 1863 1269 1867 1270
rect 1887 1274 1891 1275
rect 1887 1269 1891 1270
rect 1975 1274 1979 1275
rect 1975 1269 1979 1270
rect 2055 1274 2059 1275
rect 2055 1269 2059 1270
rect 2095 1274 2099 1275
rect 2095 1269 2099 1270
rect 2143 1274 2147 1275
rect 2143 1269 2147 1270
rect 2215 1274 2219 1275
rect 2215 1269 2219 1270
rect 2239 1274 2243 1275
rect 2239 1269 2243 1270
rect 2335 1274 2339 1275
rect 2335 1269 2339 1270
rect 2351 1274 2355 1275
rect 2351 1269 2355 1270
rect 2431 1274 2435 1275
rect 2431 1269 2435 1270
rect 2503 1274 2507 1275
rect 2503 1269 2507 1270
rect 2551 1274 2555 1275
rect 2551 1269 2555 1270
rect 2679 1274 2683 1275
rect 2679 1269 2683 1270
rect 2687 1274 2691 1275
rect 2687 1269 2691 1270
rect 2855 1274 2859 1275
rect 2855 1269 2859 1270
rect 2863 1274 2867 1275
rect 2863 1269 2867 1270
rect 3039 1274 3043 1275
rect 3039 1269 3043 1270
rect 3063 1274 3067 1275
rect 3063 1269 3067 1270
rect 3231 1274 3235 1275
rect 3231 1269 3235 1270
rect 3271 1274 3275 1275
rect 3271 1269 3275 1270
rect 3431 1274 3435 1275
rect 3431 1269 3435 1270
rect 3479 1274 3483 1275
rect 3479 1269 3483 1270
rect 3575 1274 3579 1275
rect 3575 1269 3579 1270
rect 1864 1254 1866 1269
rect 2056 1264 2058 1269
rect 2144 1264 2146 1269
rect 2240 1264 2242 1269
rect 2336 1264 2338 1269
rect 2432 1264 2434 1269
rect 2552 1264 2554 1269
rect 2688 1264 2690 1269
rect 2856 1264 2858 1269
rect 3040 1264 3042 1269
rect 3232 1264 3234 1269
rect 3432 1264 3434 1269
rect 2054 1263 2060 1264
rect 2054 1259 2055 1263
rect 2059 1259 2060 1263
rect 2054 1258 2060 1259
rect 2142 1263 2148 1264
rect 2142 1259 2143 1263
rect 2147 1259 2148 1263
rect 2142 1258 2148 1259
rect 2238 1263 2244 1264
rect 2238 1259 2239 1263
rect 2243 1259 2244 1263
rect 2238 1258 2244 1259
rect 2334 1263 2340 1264
rect 2334 1259 2335 1263
rect 2339 1259 2340 1263
rect 2334 1258 2340 1259
rect 2430 1263 2436 1264
rect 2430 1259 2431 1263
rect 2435 1259 2436 1263
rect 2430 1258 2436 1259
rect 2550 1263 2556 1264
rect 2550 1259 2551 1263
rect 2555 1259 2556 1263
rect 2550 1258 2556 1259
rect 2686 1263 2692 1264
rect 2686 1259 2687 1263
rect 2691 1259 2692 1263
rect 2686 1258 2692 1259
rect 2854 1263 2860 1264
rect 2854 1259 2855 1263
rect 2859 1259 2860 1263
rect 2854 1258 2860 1259
rect 3038 1263 3044 1264
rect 3038 1259 3039 1263
rect 3043 1259 3044 1263
rect 3038 1258 3044 1259
rect 3230 1263 3236 1264
rect 3230 1259 3231 1263
rect 3235 1259 3236 1263
rect 3230 1258 3236 1259
rect 3430 1263 3436 1264
rect 3430 1259 3431 1263
rect 3435 1259 3436 1263
rect 3430 1258 3436 1259
rect 3576 1254 3578 1269
rect 1862 1253 1868 1254
rect 110 1252 116 1253
rect 110 1248 111 1252
rect 115 1248 116 1252
rect 110 1247 116 1248
rect 1822 1252 1828 1253
rect 1822 1248 1823 1252
rect 1827 1248 1828 1252
rect 1862 1249 1863 1253
rect 1867 1249 1868 1253
rect 1862 1248 1868 1249
rect 3574 1253 3580 1254
rect 3574 1249 3575 1253
rect 3579 1249 3580 1253
rect 3574 1248 3580 1249
rect 1822 1247 1828 1248
rect 1862 1236 1868 1237
rect 110 1235 116 1236
rect 110 1231 111 1235
rect 115 1231 116 1235
rect 110 1230 116 1231
rect 1822 1235 1828 1236
rect 1822 1231 1823 1235
rect 1827 1231 1828 1235
rect 1862 1232 1863 1236
rect 1867 1232 1868 1236
rect 1862 1231 1868 1232
rect 3574 1236 3580 1237
rect 3574 1232 3575 1236
rect 3579 1232 3580 1236
rect 3574 1231 3580 1232
rect 1822 1230 1828 1231
rect 112 1207 114 1230
rect 206 1225 212 1226
rect 206 1221 207 1225
rect 211 1221 212 1225
rect 206 1220 212 1221
rect 350 1225 356 1226
rect 350 1221 351 1225
rect 355 1221 356 1225
rect 350 1220 356 1221
rect 510 1225 516 1226
rect 510 1221 511 1225
rect 515 1221 516 1225
rect 510 1220 516 1221
rect 670 1225 676 1226
rect 670 1221 671 1225
rect 675 1221 676 1225
rect 670 1220 676 1221
rect 830 1225 836 1226
rect 830 1221 831 1225
rect 835 1221 836 1225
rect 830 1220 836 1221
rect 990 1225 996 1226
rect 990 1221 991 1225
rect 995 1221 996 1225
rect 990 1220 996 1221
rect 1142 1225 1148 1226
rect 1142 1221 1143 1225
rect 1147 1221 1148 1225
rect 1142 1220 1148 1221
rect 1286 1225 1292 1226
rect 1286 1221 1287 1225
rect 1291 1221 1292 1225
rect 1286 1220 1292 1221
rect 1430 1225 1436 1226
rect 1430 1221 1431 1225
rect 1435 1221 1436 1225
rect 1430 1220 1436 1221
rect 1582 1225 1588 1226
rect 1582 1221 1583 1225
rect 1587 1221 1588 1225
rect 1582 1220 1588 1221
rect 208 1207 210 1220
rect 352 1207 354 1220
rect 512 1207 514 1220
rect 672 1207 674 1220
rect 832 1207 834 1220
rect 992 1207 994 1220
rect 1144 1207 1146 1220
rect 1288 1207 1290 1220
rect 1432 1207 1434 1220
rect 1584 1207 1586 1220
rect 1824 1207 1826 1230
rect 111 1206 115 1207
rect 111 1201 115 1202
rect 135 1206 139 1207
rect 135 1201 139 1202
rect 207 1206 211 1207
rect 207 1201 211 1202
rect 271 1206 275 1207
rect 271 1201 275 1202
rect 351 1206 355 1207
rect 351 1201 355 1202
rect 423 1206 427 1207
rect 423 1201 427 1202
rect 511 1206 515 1207
rect 511 1201 515 1202
rect 575 1206 579 1207
rect 575 1201 579 1202
rect 671 1206 675 1207
rect 671 1201 675 1202
rect 727 1206 731 1207
rect 727 1201 731 1202
rect 831 1206 835 1207
rect 831 1201 835 1202
rect 887 1206 891 1207
rect 887 1201 891 1202
rect 991 1206 995 1207
rect 991 1201 995 1202
rect 1055 1206 1059 1207
rect 1055 1201 1059 1202
rect 1143 1206 1147 1207
rect 1143 1201 1147 1202
rect 1231 1206 1235 1207
rect 1231 1201 1235 1202
rect 1287 1206 1291 1207
rect 1287 1201 1291 1202
rect 1415 1206 1419 1207
rect 1415 1201 1419 1202
rect 1431 1206 1435 1207
rect 1431 1201 1435 1202
rect 1583 1206 1587 1207
rect 1583 1201 1587 1202
rect 1599 1206 1603 1207
rect 1599 1201 1603 1202
rect 1823 1206 1827 1207
rect 1864 1203 1866 1231
rect 2062 1223 2068 1224
rect 2062 1219 2063 1223
rect 2067 1219 2068 1223
rect 2062 1218 2068 1219
rect 2150 1223 2156 1224
rect 2150 1219 2151 1223
rect 2155 1219 2156 1223
rect 2150 1218 2156 1219
rect 2246 1223 2252 1224
rect 2246 1219 2247 1223
rect 2251 1219 2252 1223
rect 2246 1218 2252 1219
rect 2342 1223 2348 1224
rect 2342 1219 2343 1223
rect 2347 1219 2348 1223
rect 2342 1218 2348 1219
rect 2438 1223 2444 1224
rect 2438 1219 2439 1223
rect 2443 1219 2444 1223
rect 2438 1218 2444 1219
rect 2558 1223 2564 1224
rect 2558 1219 2559 1223
rect 2563 1219 2564 1223
rect 2558 1218 2564 1219
rect 2694 1223 2700 1224
rect 2694 1219 2695 1223
rect 2699 1219 2700 1223
rect 2694 1218 2700 1219
rect 2862 1223 2868 1224
rect 2862 1219 2863 1223
rect 2867 1219 2868 1223
rect 2862 1218 2868 1219
rect 3046 1223 3052 1224
rect 3046 1219 3047 1223
rect 3051 1219 3052 1223
rect 3046 1218 3052 1219
rect 3238 1223 3244 1224
rect 3238 1219 3239 1223
rect 3243 1219 3244 1223
rect 3238 1218 3244 1219
rect 3438 1223 3444 1224
rect 3438 1219 3439 1223
rect 3443 1219 3444 1223
rect 3438 1218 3444 1219
rect 2064 1203 2066 1218
rect 2152 1203 2154 1218
rect 2248 1203 2250 1218
rect 2344 1203 2346 1218
rect 2440 1203 2442 1218
rect 2560 1203 2562 1218
rect 2696 1203 2698 1218
rect 2864 1203 2866 1218
rect 3048 1203 3050 1218
rect 3240 1203 3242 1218
rect 3440 1203 3442 1218
rect 3576 1203 3578 1231
rect 1823 1201 1827 1202
rect 1863 1202 1867 1203
rect 112 1186 114 1201
rect 136 1196 138 1201
rect 272 1196 274 1201
rect 424 1196 426 1201
rect 576 1196 578 1201
rect 728 1196 730 1201
rect 888 1196 890 1201
rect 1056 1196 1058 1201
rect 1232 1196 1234 1201
rect 1416 1196 1418 1201
rect 1600 1196 1602 1201
rect 134 1195 140 1196
rect 134 1191 135 1195
rect 139 1191 140 1195
rect 134 1190 140 1191
rect 270 1195 276 1196
rect 270 1191 271 1195
rect 275 1191 276 1195
rect 270 1190 276 1191
rect 422 1195 428 1196
rect 422 1191 423 1195
rect 427 1191 428 1195
rect 422 1190 428 1191
rect 574 1195 580 1196
rect 574 1191 575 1195
rect 579 1191 580 1195
rect 574 1190 580 1191
rect 726 1195 732 1196
rect 726 1191 727 1195
rect 731 1191 732 1195
rect 726 1190 732 1191
rect 886 1195 892 1196
rect 886 1191 887 1195
rect 891 1191 892 1195
rect 886 1190 892 1191
rect 1054 1195 1060 1196
rect 1054 1191 1055 1195
rect 1059 1191 1060 1195
rect 1054 1190 1060 1191
rect 1230 1195 1236 1196
rect 1230 1191 1231 1195
rect 1235 1191 1236 1195
rect 1230 1190 1236 1191
rect 1414 1195 1420 1196
rect 1414 1191 1415 1195
rect 1419 1191 1420 1195
rect 1414 1190 1420 1191
rect 1598 1195 1604 1196
rect 1598 1191 1599 1195
rect 1603 1191 1604 1195
rect 1598 1190 1604 1191
rect 1824 1186 1826 1201
rect 1863 1197 1867 1198
rect 2039 1202 2043 1203
rect 2039 1197 2043 1198
rect 2063 1202 2067 1203
rect 2063 1197 2067 1198
rect 2151 1202 2155 1203
rect 2151 1197 2155 1198
rect 2247 1202 2251 1203
rect 2247 1197 2251 1198
rect 2279 1202 2283 1203
rect 2279 1197 2283 1198
rect 2343 1202 2347 1203
rect 2343 1197 2347 1198
rect 2415 1202 2419 1203
rect 2415 1197 2419 1198
rect 2439 1202 2443 1203
rect 2439 1197 2443 1198
rect 2559 1202 2563 1203
rect 2559 1197 2563 1198
rect 2695 1202 2699 1203
rect 2695 1197 2699 1198
rect 2711 1202 2715 1203
rect 2711 1197 2715 1198
rect 2863 1202 2867 1203
rect 2863 1197 2867 1198
rect 3015 1202 3019 1203
rect 3015 1197 3019 1198
rect 3047 1202 3051 1203
rect 3047 1197 3051 1198
rect 3167 1202 3171 1203
rect 3167 1197 3171 1198
rect 3239 1202 3243 1203
rect 3239 1197 3243 1198
rect 3327 1202 3331 1203
rect 3327 1197 3331 1198
rect 3439 1202 3443 1203
rect 3439 1197 3443 1198
rect 3487 1202 3491 1203
rect 3487 1197 3491 1198
rect 3575 1202 3579 1203
rect 3575 1197 3579 1198
rect 110 1185 116 1186
rect 110 1181 111 1185
rect 115 1181 116 1185
rect 110 1180 116 1181
rect 1822 1185 1828 1186
rect 1822 1181 1823 1185
rect 1827 1181 1828 1185
rect 1822 1180 1828 1181
rect 1864 1173 1866 1197
rect 2040 1186 2042 1197
rect 2152 1186 2154 1197
rect 2280 1186 2282 1197
rect 2416 1186 2418 1197
rect 2560 1186 2562 1197
rect 2712 1186 2714 1197
rect 2864 1186 2866 1197
rect 3016 1186 3018 1197
rect 3168 1186 3170 1197
rect 3328 1186 3330 1197
rect 3488 1186 3490 1197
rect 2038 1185 2044 1186
rect 2038 1181 2039 1185
rect 2043 1181 2044 1185
rect 2038 1180 2044 1181
rect 2150 1185 2156 1186
rect 2150 1181 2151 1185
rect 2155 1181 2156 1185
rect 2150 1180 2156 1181
rect 2278 1185 2284 1186
rect 2278 1181 2279 1185
rect 2283 1181 2284 1185
rect 2278 1180 2284 1181
rect 2414 1185 2420 1186
rect 2414 1181 2415 1185
rect 2419 1181 2420 1185
rect 2414 1180 2420 1181
rect 2558 1185 2564 1186
rect 2558 1181 2559 1185
rect 2563 1181 2564 1185
rect 2558 1180 2564 1181
rect 2710 1185 2716 1186
rect 2710 1181 2711 1185
rect 2715 1181 2716 1185
rect 2710 1180 2716 1181
rect 2862 1185 2868 1186
rect 2862 1181 2863 1185
rect 2867 1181 2868 1185
rect 2862 1180 2868 1181
rect 3014 1185 3020 1186
rect 3014 1181 3015 1185
rect 3019 1181 3020 1185
rect 3014 1180 3020 1181
rect 3166 1185 3172 1186
rect 3166 1181 3167 1185
rect 3171 1181 3172 1185
rect 3166 1180 3172 1181
rect 3326 1185 3332 1186
rect 3326 1181 3327 1185
rect 3331 1181 3332 1185
rect 3326 1180 3332 1181
rect 3486 1185 3492 1186
rect 3486 1181 3487 1185
rect 3491 1181 3492 1185
rect 3486 1180 3492 1181
rect 3576 1173 3578 1197
rect 1862 1172 1868 1173
rect 110 1168 116 1169
rect 110 1164 111 1168
rect 115 1164 116 1168
rect 110 1163 116 1164
rect 1822 1168 1828 1169
rect 1822 1164 1823 1168
rect 1827 1164 1828 1168
rect 1862 1168 1863 1172
rect 1867 1168 1868 1172
rect 1862 1167 1868 1168
rect 3574 1172 3580 1173
rect 3574 1168 3575 1172
rect 3579 1168 3580 1172
rect 3574 1167 3580 1168
rect 1822 1163 1828 1164
rect 112 1139 114 1163
rect 142 1155 148 1156
rect 142 1151 143 1155
rect 147 1151 148 1155
rect 142 1150 148 1151
rect 278 1155 284 1156
rect 278 1151 279 1155
rect 283 1151 284 1155
rect 278 1150 284 1151
rect 430 1155 436 1156
rect 430 1151 431 1155
rect 435 1151 436 1155
rect 430 1150 436 1151
rect 582 1155 588 1156
rect 582 1151 583 1155
rect 587 1151 588 1155
rect 582 1150 588 1151
rect 734 1155 740 1156
rect 734 1151 735 1155
rect 739 1151 740 1155
rect 734 1150 740 1151
rect 894 1155 900 1156
rect 894 1151 895 1155
rect 899 1151 900 1155
rect 894 1150 900 1151
rect 1062 1155 1068 1156
rect 1062 1151 1063 1155
rect 1067 1151 1068 1155
rect 1062 1150 1068 1151
rect 1238 1155 1244 1156
rect 1238 1151 1239 1155
rect 1243 1151 1244 1155
rect 1238 1150 1244 1151
rect 1422 1155 1428 1156
rect 1422 1151 1423 1155
rect 1427 1151 1428 1155
rect 1422 1150 1428 1151
rect 1606 1155 1612 1156
rect 1606 1151 1607 1155
rect 1611 1151 1612 1155
rect 1606 1150 1612 1151
rect 144 1139 146 1150
rect 280 1139 282 1150
rect 432 1139 434 1150
rect 584 1139 586 1150
rect 736 1139 738 1150
rect 896 1139 898 1150
rect 1064 1139 1066 1150
rect 1240 1139 1242 1150
rect 1424 1139 1426 1150
rect 1608 1139 1610 1150
rect 1824 1139 1826 1163
rect 1862 1155 1868 1156
rect 1862 1151 1863 1155
rect 1867 1151 1868 1155
rect 1862 1150 1868 1151
rect 3574 1155 3580 1156
rect 3574 1151 3575 1155
rect 3579 1151 3580 1155
rect 3574 1150 3580 1151
rect 111 1138 115 1139
rect 111 1133 115 1134
rect 143 1138 147 1139
rect 143 1133 147 1134
rect 279 1138 283 1139
rect 279 1133 283 1134
rect 295 1138 299 1139
rect 295 1133 299 1134
rect 431 1138 435 1139
rect 431 1133 435 1134
rect 479 1138 483 1139
rect 479 1133 483 1134
rect 583 1138 587 1139
rect 583 1133 587 1134
rect 663 1138 667 1139
rect 663 1133 667 1134
rect 735 1138 739 1139
rect 735 1133 739 1134
rect 847 1138 851 1139
rect 847 1133 851 1134
rect 895 1138 899 1139
rect 895 1133 899 1134
rect 1031 1138 1035 1139
rect 1031 1133 1035 1134
rect 1063 1138 1067 1139
rect 1063 1133 1067 1134
rect 1207 1138 1211 1139
rect 1207 1133 1211 1134
rect 1239 1138 1243 1139
rect 1239 1133 1243 1134
rect 1391 1138 1395 1139
rect 1391 1133 1395 1134
rect 1423 1138 1427 1139
rect 1423 1133 1427 1134
rect 1575 1138 1579 1139
rect 1575 1133 1579 1134
rect 1607 1138 1611 1139
rect 1607 1133 1611 1134
rect 1735 1138 1739 1139
rect 1735 1133 1739 1134
rect 1823 1138 1827 1139
rect 1823 1133 1827 1134
rect 112 1109 114 1133
rect 144 1122 146 1133
rect 296 1122 298 1133
rect 480 1122 482 1133
rect 664 1122 666 1133
rect 848 1122 850 1133
rect 1032 1122 1034 1133
rect 1208 1122 1210 1133
rect 1392 1122 1394 1133
rect 1576 1122 1578 1133
rect 1736 1122 1738 1133
rect 142 1121 148 1122
rect 142 1117 143 1121
rect 147 1117 148 1121
rect 142 1116 148 1117
rect 294 1121 300 1122
rect 294 1117 295 1121
rect 299 1117 300 1121
rect 294 1116 300 1117
rect 478 1121 484 1122
rect 478 1117 479 1121
rect 483 1117 484 1121
rect 478 1116 484 1117
rect 662 1121 668 1122
rect 662 1117 663 1121
rect 667 1117 668 1121
rect 662 1116 668 1117
rect 846 1121 852 1122
rect 846 1117 847 1121
rect 851 1117 852 1121
rect 846 1116 852 1117
rect 1030 1121 1036 1122
rect 1030 1117 1031 1121
rect 1035 1117 1036 1121
rect 1030 1116 1036 1117
rect 1206 1121 1212 1122
rect 1206 1117 1207 1121
rect 1211 1117 1212 1121
rect 1206 1116 1212 1117
rect 1390 1121 1396 1122
rect 1390 1117 1391 1121
rect 1395 1117 1396 1121
rect 1390 1116 1396 1117
rect 1574 1121 1580 1122
rect 1574 1117 1575 1121
rect 1579 1117 1580 1121
rect 1574 1116 1580 1117
rect 1734 1121 1740 1122
rect 1734 1117 1735 1121
rect 1739 1117 1740 1121
rect 1734 1116 1740 1117
rect 1824 1109 1826 1133
rect 1864 1123 1866 1150
rect 2030 1145 2036 1146
rect 2030 1141 2031 1145
rect 2035 1141 2036 1145
rect 2030 1140 2036 1141
rect 2142 1145 2148 1146
rect 2142 1141 2143 1145
rect 2147 1141 2148 1145
rect 2142 1140 2148 1141
rect 2270 1145 2276 1146
rect 2270 1141 2271 1145
rect 2275 1141 2276 1145
rect 2270 1140 2276 1141
rect 2406 1145 2412 1146
rect 2406 1141 2407 1145
rect 2411 1141 2412 1145
rect 2406 1140 2412 1141
rect 2550 1145 2556 1146
rect 2550 1141 2551 1145
rect 2555 1141 2556 1145
rect 2550 1140 2556 1141
rect 2702 1145 2708 1146
rect 2702 1141 2703 1145
rect 2707 1141 2708 1145
rect 2702 1140 2708 1141
rect 2854 1145 2860 1146
rect 2854 1141 2855 1145
rect 2859 1141 2860 1145
rect 2854 1140 2860 1141
rect 3006 1145 3012 1146
rect 3006 1141 3007 1145
rect 3011 1141 3012 1145
rect 3006 1140 3012 1141
rect 3158 1145 3164 1146
rect 3158 1141 3159 1145
rect 3163 1141 3164 1145
rect 3158 1140 3164 1141
rect 3318 1145 3324 1146
rect 3318 1141 3319 1145
rect 3323 1141 3324 1145
rect 3318 1140 3324 1141
rect 3478 1145 3484 1146
rect 3478 1141 3479 1145
rect 3483 1141 3484 1145
rect 3478 1140 3484 1141
rect 2032 1123 2034 1140
rect 2144 1123 2146 1140
rect 2272 1123 2274 1140
rect 2408 1123 2410 1140
rect 2552 1123 2554 1140
rect 2704 1123 2706 1140
rect 2856 1123 2858 1140
rect 3008 1123 3010 1140
rect 3160 1123 3162 1140
rect 3320 1123 3322 1140
rect 3480 1123 3482 1140
rect 3576 1123 3578 1150
rect 1863 1122 1867 1123
rect 1863 1117 1867 1118
rect 1943 1122 1947 1123
rect 1943 1117 1947 1118
rect 2031 1122 2035 1123
rect 2031 1117 2035 1118
rect 2087 1122 2091 1123
rect 2087 1117 2091 1118
rect 2143 1122 2147 1123
rect 2143 1117 2147 1118
rect 2231 1122 2235 1123
rect 2231 1117 2235 1118
rect 2271 1122 2275 1123
rect 2271 1117 2275 1118
rect 2383 1122 2387 1123
rect 2383 1117 2387 1118
rect 2407 1122 2411 1123
rect 2407 1117 2411 1118
rect 2535 1122 2539 1123
rect 2535 1117 2539 1118
rect 2551 1122 2555 1123
rect 2551 1117 2555 1118
rect 2687 1122 2691 1123
rect 2687 1117 2691 1118
rect 2703 1122 2707 1123
rect 2703 1117 2707 1118
rect 2839 1122 2843 1123
rect 2839 1117 2843 1118
rect 2855 1122 2859 1123
rect 2855 1117 2859 1118
rect 2991 1122 2995 1123
rect 2991 1117 2995 1118
rect 3007 1122 3011 1123
rect 3007 1117 3011 1118
rect 3151 1122 3155 1123
rect 3151 1117 3155 1118
rect 3159 1122 3163 1123
rect 3159 1117 3163 1118
rect 3319 1122 3323 1123
rect 3319 1117 3323 1118
rect 3479 1122 3483 1123
rect 3479 1117 3483 1118
rect 3575 1122 3579 1123
rect 3575 1117 3579 1118
rect 110 1108 116 1109
rect 110 1104 111 1108
rect 115 1104 116 1108
rect 110 1103 116 1104
rect 1822 1108 1828 1109
rect 1822 1104 1823 1108
rect 1827 1104 1828 1108
rect 1822 1103 1828 1104
rect 1864 1102 1866 1117
rect 1944 1112 1946 1117
rect 2088 1112 2090 1117
rect 2232 1112 2234 1117
rect 2384 1112 2386 1117
rect 2536 1112 2538 1117
rect 2688 1112 2690 1117
rect 2840 1112 2842 1117
rect 2992 1112 2994 1117
rect 3152 1112 3154 1117
rect 3320 1112 3322 1117
rect 3480 1112 3482 1117
rect 1942 1111 1948 1112
rect 1942 1107 1943 1111
rect 1947 1107 1948 1111
rect 1942 1106 1948 1107
rect 2086 1111 2092 1112
rect 2086 1107 2087 1111
rect 2091 1107 2092 1111
rect 2086 1106 2092 1107
rect 2230 1111 2236 1112
rect 2230 1107 2231 1111
rect 2235 1107 2236 1111
rect 2230 1106 2236 1107
rect 2382 1111 2388 1112
rect 2382 1107 2383 1111
rect 2387 1107 2388 1111
rect 2382 1106 2388 1107
rect 2534 1111 2540 1112
rect 2534 1107 2535 1111
rect 2539 1107 2540 1111
rect 2534 1106 2540 1107
rect 2686 1111 2692 1112
rect 2686 1107 2687 1111
rect 2691 1107 2692 1111
rect 2686 1106 2692 1107
rect 2838 1111 2844 1112
rect 2838 1107 2839 1111
rect 2843 1107 2844 1111
rect 2838 1106 2844 1107
rect 2990 1111 2996 1112
rect 2990 1107 2991 1111
rect 2995 1107 2996 1111
rect 2990 1106 2996 1107
rect 3150 1111 3156 1112
rect 3150 1107 3151 1111
rect 3155 1107 3156 1111
rect 3150 1106 3156 1107
rect 3318 1111 3324 1112
rect 3318 1107 3319 1111
rect 3323 1107 3324 1111
rect 3318 1106 3324 1107
rect 3478 1111 3484 1112
rect 3478 1107 3479 1111
rect 3483 1107 3484 1111
rect 3478 1106 3484 1107
rect 3576 1102 3578 1117
rect 1862 1101 1868 1102
rect 1862 1097 1863 1101
rect 1867 1097 1868 1101
rect 1862 1096 1868 1097
rect 3574 1101 3580 1102
rect 3574 1097 3575 1101
rect 3579 1097 3580 1101
rect 3574 1096 3580 1097
rect 110 1091 116 1092
rect 110 1087 111 1091
rect 115 1087 116 1091
rect 110 1086 116 1087
rect 1822 1091 1828 1092
rect 1822 1087 1823 1091
rect 1827 1087 1828 1091
rect 1822 1086 1828 1087
rect 112 1071 114 1086
rect 134 1081 140 1082
rect 134 1077 135 1081
rect 139 1077 140 1081
rect 134 1076 140 1077
rect 286 1081 292 1082
rect 286 1077 287 1081
rect 291 1077 292 1081
rect 286 1076 292 1077
rect 470 1081 476 1082
rect 470 1077 471 1081
rect 475 1077 476 1081
rect 470 1076 476 1077
rect 654 1081 660 1082
rect 654 1077 655 1081
rect 659 1077 660 1081
rect 654 1076 660 1077
rect 838 1081 844 1082
rect 838 1077 839 1081
rect 843 1077 844 1081
rect 838 1076 844 1077
rect 1022 1081 1028 1082
rect 1022 1077 1023 1081
rect 1027 1077 1028 1081
rect 1022 1076 1028 1077
rect 1198 1081 1204 1082
rect 1198 1077 1199 1081
rect 1203 1077 1204 1081
rect 1198 1076 1204 1077
rect 1382 1081 1388 1082
rect 1382 1077 1383 1081
rect 1387 1077 1388 1081
rect 1382 1076 1388 1077
rect 1566 1081 1572 1082
rect 1566 1077 1567 1081
rect 1571 1077 1572 1081
rect 1566 1076 1572 1077
rect 1726 1081 1732 1082
rect 1726 1077 1727 1081
rect 1731 1077 1732 1081
rect 1726 1076 1732 1077
rect 136 1071 138 1076
rect 288 1071 290 1076
rect 472 1071 474 1076
rect 656 1071 658 1076
rect 840 1071 842 1076
rect 1024 1071 1026 1076
rect 1200 1071 1202 1076
rect 1384 1071 1386 1076
rect 1568 1071 1570 1076
rect 1728 1071 1730 1076
rect 1824 1071 1826 1086
rect 1862 1084 1868 1085
rect 1862 1080 1863 1084
rect 1867 1080 1868 1084
rect 1862 1079 1868 1080
rect 3574 1084 3580 1085
rect 3574 1080 3575 1084
rect 3579 1080 3580 1084
rect 3574 1079 3580 1080
rect 111 1070 115 1071
rect 111 1065 115 1066
rect 135 1070 139 1071
rect 135 1065 139 1066
rect 271 1070 275 1071
rect 271 1065 275 1066
rect 287 1070 291 1071
rect 287 1065 291 1066
rect 431 1070 435 1071
rect 431 1065 435 1066
rect 471 1070 475 1071
rect 471 1065 475 1066
rect 583 1070 587 1071
rect 583 1065 587 1066
rect 655 1070 659 1071
rect 655 1065 659 1066
rect 735 1070 739 1071
rect 735 1065 739 1066
rect 839 1070 843 1071
rect 839 1065 843 1066
rect 887 1070 891 1071
rect 887 1065 891 1066
rect 1023 1070 1027 1071
rect 1023 1065 1027 1066
rect 1047 1070 1051 1071
rect 1047 1065 1051 1066
rect 1199 1070 1203 1071
rect 1199 1065 1203 1066
rect 1215 1070 1219 1071
rect 1215 1065 1219 1066
rect 1383 1070 1387 1071
rect 1383 1065 1387 1066
rect 1559 1070 1563 1071
rect 1559 1065 1563 1066
rect 1567 1070 1571 1071
rect 1567 1065 1571 1066
rect 1727 1070 1731 1071
rect 1727 1065 1731 1066
rect 1823 1070 1827 1071
rect 1823 1065 1827 1066
rect 112 1050 114 1065
rect 136 1060 138 1065
rect 272 1060 274 1065
rect 432 1060 434 1065
rect 584 1060 586 1065
rect 736 1060 738 1065
rect 888 1060 890 1065
rect 1048 1060 1050 1065
rect 1216 1060 1218 1065
rect 1384 1060 1386 1065
rect 1560 1060 1562 1065
rect 1728 1060 1730 1065
rect 134 1059 140 1060
rect 134 1055 135 1059
rect 139 1055 140 1059
rect 134 1054 140 1055
rect 270 1059 276 1060
rect 270 1055 271 1059
rect 275 1055 276 1059
rect 270 1054 276 1055
rect 430 1059 436 1060
rect 430 1055 431 1059
rect 435 1055 436 1059
rect 430 1054 436 1055
rect 582 1059 588 1060
rect 582 1055 583 1059
rect 587 1055 588 1059
rect 582 1054 588 1055
rect 734 1059 740 1060
rect 734 1055 735 1059
rect 739 1055 740 1059
rect 734 1054 740 1055
rect 886 1059 892 1060
rect 886 1055 887 1059
rect 891 1055 892 1059
rect 886 1054 892 1055
rect 1046 1059 1052 1060
rect 1046 1055 1047 1059
rect 1051 1055 1052 1059
rect 1046 1054 1052 1055
rect 1214 1059 1220 1060
rect 1214 1055 1215 1059
rect 1219 1055 1220 1059
rect 1214 1054 1220 1055
rect 1382 1059 1388 1060
rect 1382 1055 1383 1059
rect 1387 1055 1388 1059
rect 1382 1054 1388 1055
rect 1558 1059 1564 1060
rect 1558 1055 1559 1059
rect 1563 1055 1564 1059
rect 1558 1054 1564 1055
rect 1726 1059 1732 1060
rect 1726 1055 1727 1059
rect 1731 1055 1732 1059
rect 1726 1054 1732 1055
rect 1824 1050 1826 1065
rect 110 1049 116 1050
rect 110 1045 111 1049
rect 115 1045 116 1049
rect 110 1044 116 1045
rect 1822 1049 1828 1050
rect 1822 1045 1823 1049
rect 1827 1045 1828 1049
rect 1822 1044 1828 1045
rect 1864 1043 1866 1079
rect 1950 1071 1956 1072
rect 1950 1067 1951 1071
rect 1955 1067 1956 1071
rect 1950 1066 1956 1067
rect 2094 1071 2100 1072
rect 2094 1067 2095 1071
rect 2099 1067 2100 1071
rect 2094 1066 2100 1067
rect 2238 1071 2244 1072
rect 2238 1067 2239 1071
rect 2243 1067 2244 1071
rect 2238 1066 2244 1067
rect 2390 1071 2396 1072
rect 2390 1067 2391 1071
rect 2395 1067 2396 1071
rect 2390 1066 2396 1067
rect 2542 1071 2548 1072
rect 2542 1067 2543 1071
rect 2547 1067 2548 1071
rect 2542 1066 2548 1067
rect 2694 1071 2700 1072
rect 2694 1067 2695 1071
rect 2699 1067 2700 1071
rect 2694 1066 2700 1067
rect 2846 1071 2852 1072
rect 2846 1067 2847 1071
rect 2851 1067 2852 1071
rect 2846 1066 2852 1067
rect 2998 1071 3004 1072
rect 2998 1067 2999 1071
rect 3003 1067 3004 1071
rect 2998 1066 3004 1067
rect 3158 1071 3164 1072
rect 3158 1067 3159 1071
rect 3163 1067 3164 1071
rect 3158 1066 3164 1067
rect 3326 1071 3332 1072
rect 3326 1067 3327 1071
rect 3331 1067 3332 1071
rect 3326 1066 3332 1067
rect 3486 1071 3492 1072
rect 3486 1067 3487 1071
rect 3491 1067 3492 1071
rect 3486 1066 3492 1067
rect 1952 1043 1954 1066
rect 2096 1043 2098 1066
rect 2240 1043 2242 1066
rect 2392 1043 2394 1066
rect 2544 1043 2546 1066
rect 2696 1043 2698 1066
rect 2848 1043 2850 1066
rect 3000 1043 3002 1066
rect 3160 1043 3162 1066
rect 3328 1043 3330 1066
rect 3488 1043 3490 1066
rect 3576 1043 3578 1079
rect 1863 1042 1867 1043
rect 1863 1037 1867 1038
rect 1919 1042 1923 1043
rect 1919 1037 1923 1038
rect 1951 1042 1955 1043
rect 1951 1037 1955 1038
rect 2095 1042 2099 1043
rect 2095 1037 2099 1038
rect 2127 1042 2131 1043
rect 2127 1037 2131 1038
rect 2239 1042 2243 1043
rect 2239 1037 2243 1038
rect 2327 1042 2331 1043
rect 2327 1037 2331 1038
rect 2391 1042 2395 1043
rect 2391 1037 2395 1038
rect 2519 1042 2523 1043
rect 2519 1037 2523 1038
rect 2543 1042 2547 1043
rect 2543 1037 2547 1038
rect 2695 1042 2699 1043
rect 2695 1037 2699 1038
rect 2847 1042 2851 1043
rect 2847 1037 2851 1038
rect 2863 1042 2867 1043
rect 2863 1037 2867 1038
rect 2999 1042 3003 1043
rect 2999 1037 3003 1038
rect 3023 1042 3027 1043
rect 3023 1037 3027 1038
rect 3159 1042 3163 1043
rect 3159 1037 3163 1038
rect 3183 1042 3187 1043
rect 3183 1037 3187 1038
rect 3327 1042 3331 1043
rect 3327 1037 3331 1038
rect 3343 1042 3347 1043
rect 3343 1037 3347 1038
rect 3487 1042 3491 1043
rect 3487 1037 3491 1038
rect 3575 1042 3579 1043
rect 3575 1037 3579 1038
rect 110 1032 116 1033
rect 110 1028 111 1032
rect 115 1028 116 1032
rect 110 1027 116 1028
rect 1822 1032 1828 1033
rect 1822 1028 1823 1032
rect 1827 1028 1828 1032
rect 1822 1027 1828 1028
rect 112 999 114 1027
rect 142 1019 148 1020
rect 142 1015 143 1019
rect 147 1015 148 1019
rect 142 1014 148 1015
rect 278 1019 284 1020
rect 278 1015 279 1019
rect 283 1015 284 1019
rect 278 1014 284 1015
rect 438 1019 444 1020
rect 438 1015 439 1019
rect 443 1015 444 1019
rect 438 1014 444 1015
rect 590 1019 596 1020
rect 590 1015 591 1019
rect 595 1015 596 1019
rect 590 1014 596 1015
rect 742 1019 748 1020
rect 742 1015 743 1019
rect 747 1015 748 1019
rect 742 1014 748 1015
rect 894 1019 900 1020
rect 894 1015 895 1019
rect 899 1015 900 1019
rect 894 1014 900 1015
rect 1054 1019 1060 1020
rect 1054 1015 1055 1019
rect 1059 1015 1060 1019
rect 1054 1014 1060 1015
rect 1222 1019 1228 1020
rect 1222 1015 1223 1019
rect 1227 1015 1228 1019
rect 1222 1014 1228 1015
rect 1390 1019 1396 1020
rect 1390 1015 1391 1019
rect 1395 1015 1396 1019
rect 1390 1014 1396 1015
rect 1566 1019 1572 1020
rect 1566 1015 1567 1019
rect 1571 1015 1572 1019
rect 1566 1014 1572 1015
rect 1734 1019 1740 1020
rect 1734 1015 1735 1019
rect 1739 1015 1740 1019
rect 1734 1014 1740 1015
rect 144 999 146 1014
rect 280 999 282 1014
rect 440 999 442 1014
rect 592 999 594 1014
rect 744 999 746 1014
rect 896 999 898 1014
rect 1056 999 1058 1014
rect 1224 999 1226 1014
rect 1392 999 1394 1014
rect 1568 999 1570 1014
rect 1736 999 1738 1014
rect 1824 999 1826 1027
rect 1864 1013 1866 1037
rect 1920 1026 1922 1037
rect 2128 1026 2130 1037
rect 2328 1026 2330 1037
rect 2520 1026 2522 1037
rect 2696 1026 2698 1037
rect 2864 1026 2866 1037
rect 3024 1026 3026 1037
rect 3184 1026 3186 1037
rect 3344 1026 3346 1037
rect 3488 1026 3490 1037
rect 1918 1025 1924 1026
rect 1918 1021 1919 1025
rect 1923 1021 1924 1025
rect 1918 1020 1924 1021
rect 2126 1025 2132 1026
rect 2126 1021 2127 1025
rect 2131 1021 2132 1025
rect 2126 1020 2132 1021
rect 2326 1025 2332 1026
rect 2326 1021 2327 1025
rect 2331 1021 2332 1025
rect 2326 1020 2332 1021
rect 2518 1025 2524 1026
rect 2518 1021 2519 1025
rect 2523 1021 2524 1025
rect 2518 1020 2524 1021
rect 2694 1025 2700 1026
rect 2694 1021 2695 1025
rect 2699 1021 2700 1025
rect 2694 1020 2700 1021
rect 2862 1025 2868 1026
rect 2862 1021 2863 1025
rect 2867 1021 2868 1025
rect 2862 1020 2868 1021
rect 3022 1025 3028 1026
rect 3022 1021 3023 1025
rect 3027 1021 3028 1025
rect 3022 1020 3028 1021
rect 3182 1025 3188 1026
rect 3182 1021 3183 1025
rect 3187 1021 3188 1025
rect 3182 1020 3188 1021
rect 3342 1025 3348 1026
rect 3342 1021 3343 1025
rect 3347 1021 3348 1025
rect 3342 1020 3348 1021
rect 3486 1025 3492 1026
rect 3486 1021 3487 1025
rect 3491 1021 3492 1025
rect 3486 1020 3492 1021
rect 3576 1013 3578 1037
rect 1862 1012 1868 1013
rect 1862 1008 1863 1012
rect 1867 1008 1868 1012
rect 1862 1007 1868 1008
rect 3574 1012 3580 1013
rect 3574 1008 3575 1012
rect 3579 1008 3580 1012
rect 3574 1007 3580 1008
rect 111 998 115 999
rect 111 993 115 994
rect 143 998 147 999
rect 143 993 147 994
rect 279 998 283 999
rect 279 993 283 994
rect 287 998 291 999
rect 287 993 291 994
rect 439 998 443 999
rect 439 993 443 994
rect 463 998 467 999
rect 463 993 467 994
rect 591 998 595 999
rect 591 993 595 994
rect 647 998 651 999
rect 647 993 651 994
rect 743 998 747 999
rect 743 993 747 994
rect 823 998 827 999
rect 823 993 827 994
rect 895 998 899 999
rect 895 993 899 994
rect 999 998 1003 999
rect 999 993 1003 994
rect 1055 998 1059 999
rect 1055 993 1059 994
rect 1167 998 1171 999
rect 1167 993 1171 994
rect 1223 998 1227 999
rect 1223 993 1227 994
rect 1327 998 1331 999
rect 1327 993 1331 994
rect 1391 998 1395 999
rect 1391 993 1395 994
rect 1487 998 1491 999
rect 1487 993 1491 994
rect 1567 998 1571 999
rect 1567 993 1571 994
rect 1655 998 1659 999
rect 1655 993 1659 994
rect 1735 998 1739 999
rect 1735 993 1739 994
rect 1823 998 1827 999
rect 1823 993 1827 994
rect 1862 995 1868 996
rect 112 969 114 993
rect 144 982 146 993
rect 288 982 290 993
rect 464 982 466 993
rect 648 982 650 993
rect 824 982 826 993
rect 1000 982 1002 993
rect 1168 982 1170 993
rect 1328 982 1330 993
rect 1488 982 1490 993
rect 1656 982 1658 993
rect 142 981 148 982
rect 142 977 143 981
rect 147 977 148 981
rect 142 976 148 977
rect 286 981 292 982
rect 286 977 287 981
rect 291 977 292 981
rect 286 976 292 977
rect 462 981 468 982
rect 462 977 463 981
rect 467 977 468 981
rect 462 976 468 977
rect 646 981 652 982
rect 646 977 647 981
rect 651 977 652 981
rect 646 976 652 977
rect 822 981 828 982
rect 822 977 823 981
rect 827 977 828 981
rect 822 976 828 977
rect 998 981 1004 982
rect 998 977 999 981
rect 1003 977 1004 981
rect 998 976 1004 977
rect 1166 981 1172 982
rect 1166 977 1167 981
rect 1171 977 1172 981
rect 1166 976 1172 977
rect 1326 981 1332 982
rect 1326 977 1327 981
rect 1331 977 1332 981
rect 1326 976 1332 977
rect 1486 981 1492 982
rect 1486 977 1487 981
rect 1491 977 1492 981
rect 1486 976 1492 977
rect 1654 981 1660 982
rect 1654 977 1655 981
rect 1659 977 1660 981
rect 1654 976 1660 977
rect 1824 969 1826 993
rect 1862 991 1863 995
rect 1867 991 1868 995
rect 1862 990 1868 991
rect 3574 995 3580 996
rect 3574 991 3575 995
rect 3579 991 3580 995
rect 3574 990 3580 991
rect 1864 971 1866 990
rect 1910 985 1916 986
rect 1910 981 1911 985
rect 1915 981 1916 985
rect 1910 980 1916 981
rect 2118 985 2124 986
rect 2118 981 2119 985
rect 2123 981 2124 985
rect 2118 980 2124 981
rect 2318 985 2324 986
rect 2318 981 2319 985
rect 2323 981 2324 985
rect 2318 980 2324 981
rect 2510 985 2516 986
rect 2510 981 2511 985
rect 2515 981 2516 985
rect 2510 980 2516 981
rect 2686 985 2692 986
rect 2686 981 2687 985
rect 2691 981 2692 985
rect 2686 980 2692 981
rect 2854 985 2860 986
rect 2854 981 2855 985
rect 2859 981 2860 985
rect 2854 980 2860 981
rect 3014 985 3020 986
rect 3014 981 3015 985
rect 3019 981 3020 985
rect 3014 980 3020 981
rect 3174 985 3180 986
rect 3174 981 3175 985
rect 3179 981 3180 985
rect 3174 980 3180 981
rect 3334 985 3340 986
rect 3334 981 3335 985
rect 3339 981 3340 985
rect 3334 980 3340 981
rect 3478 985 3484 986
rect 3478 981 3479 985
rect 3483 981 3484 985
rect 3478 980 3484 981
rect 1912 971 1914 980
rect 2120 971 2122 980
rect 2320 971 2322 980
rect 2512 971 2514 980
rect 2688 971 2690 980
rect 2856 971 2858 980
rect 3016 971 3018 980
rect 3176 971 3178 980
rect 3336 971 3338 980
rect 3480 971 3482 980
rect 3576 971 3578 990
rect 1863 970 1867 971
rect 110 968 116 969
rect 110 964 111 968
rect 115 964 116 968
rect 110 963 116 964
rect 1822 968 1828 969
rect 1822 964 1823 968
rect 1827 964 1828 968
rect 1863 965 1867 966
rect 1887 970 1891 971
rect 1887 965 1891 966
rect 1911 970 1915 971
rect 1911 965 1915 966
rect 2071 970 2075 971
rect 2071 965 2075 966
rect 2119 970 2123 971
rect 2119 965 2123 966
rect 2263 970 2267 971
rect 2263 965 2267 966
rect 2319 970 2323 971
rect 2319 965 2323 966
rect 2455 970 2459 971
rect 2455 965 2459 966
rect 2511 970 2515 971
rect 2511 965 2515 966
rect 2631 970 2635 971
rect 2631 965 2635 966
rect 2687 970 2691 971
rect 2687 965 2691 966
rect 2799 970 2803 971
rect 2799 965 2803 966
rect 2855 970 2859 971
rect 2855 965 2859 966
rect 2951 970 2955 971
rect 2951 965 2955 966
rect 3015 970 3019 971
rect 3015 965 3019 966
rect 3095 970 3099 971
rect 3095 965 3099 966
rect 3175 970 3179 971
rect 3175 965 3179 966
rect 3231 970 3235 971
rect 3231 965 3235 966
rect 3335 970 3339 971
rect 3335 965 3339 966
rect 3367 970 3371 971
rect 3367 965 3371 966
rect 3479 970 3483 971
rect 3479 965 3483 966
rect 3575 970 3579 971
rect 3575 965 3579 966
rect 1822 963 1828 964
rect 110 951 116 952
rect 110 947 111 951
rect 115 947 116 951
rect 110 946 116 947
rect 1822 951 1828 952
rect 1822 947 1823 951
rect 1827 947 1828 951
rect 1864 950 1866 965
rect 1888 960 1890 965
rect 2072 960 2074 965
rect 2264 960 2266 965
rect 2456 960 2458 965
rect 2632 960 2634 965
rect 2800 960 2802 965
rect 2952 960 2954 965
rect 3096 960 3098 965
rect 3232 960 3234 965
rect 3368 960 3370 965
rect 3480 960 3482 965
rect 1886 959 1892 960
rect 1886 955 1887 959
rect 1891 955 1892 959
rect 1886 954 1892 955
rect 2070 959 2076 960
rect 2070 955 2071 959
rect 2075 955 2076 959
rect 2070 954 2076 955
rect 2262 959 2268 960
rect 2262 955 2263 959
rect 2267 955 2268 959
rect 2262 954 2268 955
rect 2454 959 2460 960
rect 2454 955 2455 959
rect 2459 955 2460 959
rect 2454 954 2460 955
rect 2630 959 2636 960
rect 2630 955 2631 959
rect 2635 955 2636 959
rect 2630 954 2636 955
rect 2798 959 2804 960
rect 2798 955 2799 959
rect 2803 955 2804 959
rect 2798 954 2804 955
rect 2950 959 2956 960
rect 2950 955 2951 959
rect 2955 955 2956 959
rect 2950 954 2956 955
rect 3094 959 3100 960
rect 3094 955 3095 959
rect 3099 955 3100 959
rect 3094 954 3100 955
rect 3230 959 3236 960
rect 3230 955 3231 959
rect 3235 955 3236 959
rect 3230 954 3236 955
rect 3366 959 3372 960
rect 3366 955 3367 959
rect 3371 955 3372 959
rect 3366 954 3372 955
rect 3478 959 3484 960
rect 3478 955 3479 959
rect 3483 955 3484 959
rect 3478 954 3484 955
rect 3576 950 3578 965
rect 1822 946 1828 947
rect 1862 949 1868 950
rect 112 923 114 946
rect 134 941 140 942
rect 134 937 135 941
rect 139 937 140 941
rect 134 936 140 937
rect 278 941 284 942
rect 278 937 279 941
rect 283 937 284 941
rect 278 936 284 937
rect 454 941 460 942
rect 454 937 455 941
rect 459 937 460 941
rect 454 936 460 937
rect 638 941 644 942
rect 638 937 639 941
rect 643 937 644 941
rect 638 936 644 937
rect 814 941 820 942
rect 814 937 815 941
rect 819 937 820 941
rect 814 936 820 937
rect 990 941 996 942
rect 990 937 991 941
rect 995 937 996 941
rect 990 936 996 937
rect 1158 941 1164 942
rect 1158 937 1159 941
rect 1163 937 1164 941
rect 1158 936 1164 937
rect 1318 941 1324 942
rect 1318 937 1319 941
rect 1323 937 1324 941
rect 1318 936 1324 937
rect 1478 941 1484 942
rect 1478 937 1479 941
rect 1483 937 1484 941
rect 1478 936 1484 937
rect 1646 941 1652 942
rect 1646 937 1647 941
rect 1651 937 1652 941
rect 1646 936 1652 937
rect 136 923 138 936
rect 280 923 282 936
rect 456 923 458 936
rect 640 923 642 936
rect 816 923 818 936
rect 992 923 994 936
rect 1160 923 1162 936
rect 1320 923 1322 936
rect 1480 923 1482 936
rect 1648 923 1650 936
rect 1824 923 1826 946
rect 1862 945 1863 949
rect 1867 945 1868 949
rect 1862 944 1868 945
rect 3574 949 3580 950
rect 3574 945 3575 949
rect 3579 945 3580 949
rect 3574 944 3580 945
rect 1862 932 1868 933
rect 1862 928 1863 932
rect 1867 928 1868 932
rect 1862 927 1868 928
rect 3574 932 3580 933
rect 3574 928 3575 932
rect 3579 928 3580 932
rect 3574 927 3580 928
rect 111 922 115 923
rect 111 917 115 918
rect 135 922 139 923
rect 135 917 139 918
rect 271 922 275 923
rect 271 917 275 918
rect 279 922 283 923
rect 279 917 283 918
rect 439 922 443 923
rect 439 917 443 918
rect 455 922 459 923
rect 455 917 459 918
rect 607 922 611 923
rect 607 917 611 918
rect 639 922 643 923
rect 639 917 643 918
rect 775 922 779 923
rect 775 917 779 918
rect 815 922 819 923
rect 815 917 819 918
rect 935 922 939 923
rect 935 917 939 918
rect 991 922 995 923
rect 991 917 995 918
rect 1095 922 1099 923
rect 1095 917 1099 918
rect 1159 922 1163 923
rect 1159 917 1163 918
rect 1247 922 1251 923
rect 1247 917 1251 918
rect 1319 922 1323 923
rect 1319 917 1323 918
rect 1399 922 1403 923
rect 1399 917 1403 918
rect 1479 922 1483 923
rect 1479 917 1483 918
rect 1551 922 1555 923
rect 1551 917 1555 918
rect 1647 922 1651 923
rect 1647 917 1651 918
rect 1823 922 1827 923
rect 1823 917 1827 918
rect 112 902 114 917
rect 136 912 138 917
rect 272 912 274 917
rect 440 912 442 917
rect 608 912 610 917
rect 776 912 778 917
rect 936 912 938 917
rect 1096 912 1098 917
rect 1248 912 1250 917
rect 1400 912 1402 917
rect 1552 912 1554 917
rect 134 911 140 912
rect 134 907 135 911
rect 139 907 140 911
rect 134 906 140 907
rect 270 911 276 912
rect 270 907 271 911
rect 275 907 276 911
rect 270 906 276 907
rect 438 911 444 912
rect 438 907 439 911
rect 443 907 444 911
rect 438 906 444 907
rect 606 911 612 912
rect 606 907 607 911
rect 611 907 612 911
rect 606 906 612 907
rect 774 911 780 912
rect 774 907 775 911
rect 779 907 780 911
rect 774 906 780 907
rect 934 911 940 912
rect 934 907 935 911
rect 939 907 940 911
rect 934 906 940 907
rect 1094 911 1100 912
rect 1094 907 1095 911
rect 1099 907 1100 911
rect 1094 906 1100 907
rect 1246 911 1252 912
rect 1246 907 1247 911
rect 1251 907 1252 911
rect 1246 906 1252 907
rect 1398 911 1404 912
rect 1398 907 1399 911
rect 1403 907 1404 911
rect 1398 906 1404 907
rect 1550 911 1556 912
rect 1550 907 1551 911
rect 1555 907 1556 911
rect 1550 906 1556 907
rect 1824 902 1826 917
rect 110 901 116 902
rect 110 897 111 901
rect 115 897 116 901
rect 110 896 116 897
rect 1822 901 1828 902
rect 1822 897 1823 901
rect 1827 897 1828 901
rect 1822 896 1828 897
rect 1864 895 1866 927
rect 1894 919 1900 920
rect 1894 915 1895 919
rect 1899 915 1900 919
rect 1894 914 1900 915
rect 2078 919 2084 920
rect 2078 915 2079 919
rect 2083 915 2084 919
rect 2078 914 2084 915
rect 2270 919 2276 920
rect 2270 915 2271 919
rect 2275 915 2276 919
rect 2270 914 2276 915
rect 2462 919 2468 920
rect 2462 915 2463 919
rect 2467 915 2468 919
rect 2462 914 2468 915
rect 2638 919 2644 920
rect 2638 915 2639 919
rect 2643 915 2644 919
rect 2638 914 2644 915
rect 2806 919 2812 920
rect 2806 915 2807 919
rect 2811 915 2812 919
rect 2806 914 2812 915
rect 2958 919 2964 920
rect 2958 915 2959 919
rect 2963 915 2964 919
rect 2958 914 2964 915
rect 3102 919 3108 920
rect 3102 915 3103 919
rect 3107 915 3108 919
rect 3102 914 3108 915
rect 3238 919 3244 920
rect 3238 915 3239 919
rect 3243 915 3244 919
rect 3238 914 3244 915
rect 3374 919 3380 920
rect 3374 915 3375 919
rect 3379 915 3380 919
rect 3374 914 3380 915
rect 3486 919 3492 920
rect 3486 915 3487 919
rect 3491 915 3492 919
rect 3486 914 3492 915
rect 1896 895 1898 914
rect 2080 895 2082 914
rect 2272 895 2274 914
rect 2464 895 2466 914
rect 2640 895 2642 914
rect 2808 895 2810 914
rect 2960 895 2962 914
rect 3104 895 3106 914
rect 3240 895 3242 914
rect 3376 895 3378 914
rect 3488 895 3490 914
rect 3576 895 3578 927
rect 1863 894 1867 895
rect 1863 889 1867 890
rect 1895 894 1899 895
rect 1895 889 1899 890
rect 2023 894 2027 895
rect 2023 889 2027 890
rect 2079 894 2083 895
rect 2079 889 2083 890
rect 2183 894 2187 895
rect 2183 889 2187 890
rect 2271 894 2275 895
rect 2271 889 2275 890
rect 2351 894 2355 895
rect 2351 889 2355 890
rect 2463 894 2467 895
rect 2463 889 2467 890
rect 2519 894 2523 895
rect 2519 889 2523 890
rect 2639 894 2643 895
rect 2639 889 2643 890
rect 2687 894 2691 895
rect 2687 889 2691 890
rect 2807 894 2811 895
rect 2807 889 2811 890
rect 2839 894 2843 895
rect 2839 889 2843 890
rect 2959 894 2963 895
rect 2959 889 2963 890
rect 2983 894 2987 895
rect 2983 889 2987 890
rect 3103 894 3107 895
rect 3103 889 3107 890
rect 3119 894 3123 895
rect 3119 889 3123 890
rect 3239 894 3243 895
rect 3239 889 3243 890
rect 3247 894 3251 895
rect 3247 889 3251 890
rect 3375 894 3379 895
rect 3375 889 3379 890
rect 3487 894 3491 895
rect 3487 889 3491 890
rect 3575 894 3579 895
rect 3575 889 3579 890
rect 110 884 116 885
rect 110 880 111 884
rect 115 880 116 884
rect 110 879 116 880
rect 1822 884 1828 885
rect 1822 880 1823 884
rect 1827 880 1828 884
rect 1822 879 1828 880
rect 112 855 114 879
rect 142 871 148 872
rect 142 867 143 871
rect 147 867 148 871
rect 142 866 148 867
rect 278 871 284 872
rect 278 867 279 871
rect 283 867 284 871
rect 278 866 284 867
rect 446 871 452 872
rect 446 867 447 871
rect 451 867 452 871
rect 446 866 452 867
rect 614 871 620 872
rect 614 867 615 871
rect 619 867 620 871
rect 614 866 620 867
rect 782 871 788 872
rect 782 867 783 871
rect 787 867 788 871
rect 782 866 788 867
rect 942 871 948 872
rect 942 867 943 871
rect 947 867 948 871
rect 942 866 948 867
rect 1102 871 1108 872
rect 1102 867 1103 871
rect 1107 867 1108 871
rect 1102 866 1108 867
rect 1254 871 1260 872
rect 1254 867 1255 871
rect 1259 867 1260 871
rect 1254 866 1260 867
rect 1406 871 1412 872
rect 1406 867 1407 871
rect 1411 867 1412 871
rect 1406 866 1412 867
rect 1558 871 1564 872
rect 1558 867 1559 871
rect 1563 867 1564 871
rect 1558 866 1564 867
rect 144 855 146 866
rect 280 855 282 866
rect 448 855 450 866
rect 616 855 618 866
rect 784 855 786 866
rect 944 855 946 866
rect 1104 855 1106 866
rect 1256 855 1258 866
rect 1408 855 1410 866
rect 1560 855 1562 866
rect 1824 855 1826 879
rect 1864 865 1866 889
rect 1896 878 1898 889
rect 2024 878 2026 889
rect 2184 878 2186 889
rect 2352 878 2354 889
rect 2520 878 2522 889
rect 2688 878 2690 889
rect 2840 878 2842 889
rect 2984 878 2986 889
rect 3120 878 3122 889
rect 3248 878 3250 889
rect 3376 878 3378 889
rect 3488 878 3490 889
rect 1894 877 1900 878
rect 1894 873 1895 877
rect 1899 873 1900 877
rect 1894 872 1900 873
rect 2022 877 2028 878
rect 2022 873 2023 877
rect 2027 873 2028 877
rect 2022 872 2028 873
rect 2182 877 2188 878
rect 2182 873 2183 877
rect 2187 873 2188 877
rect 2182 872 2188 873
rect 2350 877 2356 878
rect 2350 873 2351 877
rect 2355 873 2356 877
rect 2350 872 2356 873
rect 2518 877 2524 878
rect 2518 873 2519 877
rect 2523 873 2524 877
rect 2518 872 2524 873
rect 2686 877 2692 878
rect 2686 873 2687 877
rect 2691 873 2692 877
rect 2686 872 2692 873
rect 2838 877 2844 878
rect 2838 873 2839 877
rect 2843 873 2844 877
rect 2838 872 2844 873
rect 2982 877 2988 878
rect 2982 873 2983 877
rect 2987 873 2988 877
rect 2982 872 2988 873
rect 3118 877 3124 878
rect 3118 873 3119 877
rect 3123 873 3124 877
rect 3118 872 3124 873
rect 3246 877 3252 878
rect 3246 873 3247 877
rect 3251 873 3252 877
rect 3246 872 3252 873
rect 3374 877 3380 878
rect 3374 873 3375 877
rect 3379 873 3380 877
rect 3374 872 3380 873
rect 3486 877 3492 878
rect 3486 873 3487 877
rect 3491 873 3492 877
rect 3486 872 3492 873
rect 3576 865 3578 889
rect 1862 864 1868 865
rect 1862 860 1863 864
rect 1867 860 1868 864
rect 1862 859 1868 860
rect 3574 864 3580 865
rect 3574 860 3575 864
rect 3579 860 3580 864
rect 3574 859 3580 860
rect 111 854 115 855
rect 111 849 115 850
rect 143 854 147 855
rect 143 849 147 850
rect 279 854 283 855
rect 279 849 283 850
rect 287 854 291 855
rect 287 849 291 850
rect 447 854 451 855
rect 447 849 451 850
rect 463 854 467 855
rect 463 849 467 850
rect 615 854 619 855
rect 615 849 619 850
rect 639 854 643 855
rect 639 849 643 850
rect 783 854 787 855
rect 783 849 787 850
rect 807 854 811 855
rect 807 849 811 850
rect 943 854 947 855
rect 943 849 947 850
rect 983 854 987 855
rect 983 849 987 850
rect 1103 854 1107 855
rect 1103 849 1107 850
rect 1159 854 1163 855
rect 1159 849 1163 850
rect 1255 854 1259 855
rect 1255 849 1259 850
rect 1335 854 1339 855
rect 1335 849 1339 850
rect 1407 854 1411 855
rect 1407 849 1411 850
rect 1511 854 1515 855
rect 1511 849 1515 850
rect 1559 854 1563 855
rect 1559 849 1563 850
rect 1823 854 1827 855
rect 1823 849 1827 850
rect 112 825 114 849
rect 144 838 146 849
rect 288 838 290 849
rect 464 838 466 849
rect 640 838 642 849
rect 808 838 810 849
rect 984 838 986 849
rect 1160 838 1162 849
rect 1336 838 1338 849
rect 1512 838 1514 849
rect 142 837 148 838
rect 142 833 143 837
rect 147 833 148 837
rect 142 832 148 833
rect 286 837 292 838
rect 286 833 287 837
rect 291 833 292 837
rect 286 832 292 833
rect 462 837 468 838
rect 462 833 463 837
rect 467 833 468 837
rect 462 832 468 833
rect 638 837 644 838
rect 638 833 639 837
rect 643 833 644 837
rect 638 832 644 833
rect 806 837 812 838
rect 806 833 807 837
rect 811 833 812 837
rect 806 832 812 833
rect 982 837 988 838
rect 982 833 983 837
rect 987 833 988 837
rect 982 832 988 833
rect 1158 837 1164 838
rect 1158 833 1159 837
rect 1163 833 1164 837
rect 1158 832 1164 833
rect 1334 837 1340 838
rect 1334 833 1335 837
rect 1339 833 1340 837
rect 1334 832 1340 833
rect 1510 837 1516 838
rect 1510 833 1511 837
rect 1515 833 1516 837
rect 1510 832 1516 833
rect 1824 825 1826 849
rect 1862 847 1868 848
rect 1862 843 1863 847
rect 1867 843 1868 847
rect 1862 842 1868 843
rect 3574 847 3580 848
rect 3574 843 3575 847
rect 3579 843 3580 847
rect 3574 842 3580 843
rect 110 824 116 825
rect 110 820 111 824
rect 115 820 116 824
rect 110 819 116 820
rect 1822 824 1828 825
rect 1822 820 1823 824
rect 1827 820 1828 824
rect 1822 819 1828 820
rect 1864 819 1866 842
rect 1886 837 1892 838
rect 1886 833 1887 837
rect 1891 833 1892 837
rect 1886 832 1892 833
rect 2014 837 2020 838
rect 2014 833 2015 837
rect 2019 833 2020 837
rect 2014 832 2020 833
rect 2174 837 2180 838
rect 2174 833 2175 837
rect 2179 833 2180 837
rect 2174 832 2180 833
rect 2342 837 2348 838
rect 2342 833 2343 837
rect 2347 833 2348 837
rect 2342 832 2348 833
rect 2510 837 2516 838
rect 2510 833 2511 837
rect 2515 833 2516 837
rect 2510 832 2516 833
rect 2678 837 2684 838
rect 2678 833 2679 837
rect 2683 833 2684 837
rect 2678 832 2684 833
rect 2830 837 2836 838
rect 2830 833 2831 837
rect 2835 833 2836 837
rect 2830 832 2836 833
rect 2974 837 2980 838
rect 2974 833 2975 837
rect 2979 833 2980 837
rect 2974 832 2980 833
rect 3110 837 3116 838
rect 3110 833 3111 837
rect 3115 833 3116 837
rect 3110 832 3116 833
rect 3238 837 3244 838
rect 3238 833 3239 837
rect 3243 833 3244 837
rect 3238 832 3244 833
rect 3366 837 3372 838
rect 3366 833 3367 837
rect 3371 833 3372 837
rect 3366 832 3372 833
rect 3478 837 3484 838
rect 3478 833 3479 837
rect 3483 833 3484 837
rect 3478 832 3484 833
rect 1888 819 1890 832
rect 2016 819 2018 832
rect 2176 819 2178 832
rect 2344 819 2346 832
rect 2512 819 2514 832
rect 2680 819 2682 832
rect 2832 819 2834 832
rect 2976 819 2978 832
rect 3112 819 3114 832
rect 3240 819 3242 832
rect 3368 819 3370 832
rect 3480 819 3482 832
rect 3576 819 3578 842
rect 1863 818 1867 819
rect 1863 813 1867 814
rect 1887 818 1891 819
rect 1887 813 1891 814
rect 2015 818 2019 819
rect 2015 813 2019 814
rect 2071 818 2075 819
rect 2071 813 2075 814
rect 2175 818 2179 819
rect 2175 813 2179 814
rect 2263 818 2267 819
rect 2263 813 2267 814
rect 2343 818 2347 819
rect 2343 813 2347 814
rect 2447 818 2451 819
rect 2447 813 2451 814
rect 2511 818 2515 819
rect 2511 813 2515 814
rect 2623 818 2627 819
rect 2623 813 2627 814
rect 2679 818 2683 819
rect 2679 813 2683 814
rect 2791 818 2795 819
rect 2791 813 2795 814
rect 2831 818 2835 819
rect 2831 813 2835 814
rect 2943 818 2947 819
rect 2943 813 2947 814
rect 2975 818 2979 819
rect 2975 813 2979 814
rect 3087 818 3091 819
rect 3087 813 3091 814
rect 3111 818 3115 819
rect 3111 813 3115 814
rect 3223 818 3227 819
rect 3223 813 3227 814
rect 3239 818 3243 819
rect 3239 813 3243 814
rect 3359 818 3363 819
rect 3359 813 3363 814
rect 3367 818 3371 819
rect 3367 813 3371 814
rect 3479 818 3483 819
rect 3479 813 3483 814
rect 3575 818 3579 819
rect 3575 813 3579 814
rect 110 807 116 808
rect 110 803 111 807
rect 115 803 116 807
rect 110 802 116 803
rect 1822 807 1828 808
rect 1822 803 1823 807
rect 1827 803 1828 807
rect 1822 802 1828 803
rect 112 783 114 802
rect 134 797 140 798
rect 134 793 135 797
rect 139 793 140 797
rect 134 792 140 793
rect 278 797 284 798
rect 278 793 279 797
rect 283 793 284 797
rect 278 792 284 793
rect 454 797 460 798
rect 454 793 455 797
rect 459 793 460 797
rect 454 792 460 793
rect 630 797 636 798
rect 630 793 631 797
rect 635 793 636 797
rect 630 792 636 793
rect 798 797 804 798
rect 798 793 799 797
rect 803 793 804 797
rect 798 792 804 793
rect 974 797 980 798
rect 974 793 975 797
rect 979 793 980 797
rect 974 792 980 793
rect 1150 797 1156 798
rect 1150 793 1151 797
rect 1155 793 1156 797
rect 1150 792 1156 793
rect 1326 797 1332 798
rect 1326 793 1327 797
rect 1331 793 1332 797
rect 1326 792 1332 793
rect 1502 797 1508 798
rect 1502 793 1503 797
rect 1507 793 1508 797
rect 1502 792 1508 793
rect 136 783 138 792
rect 280 783 282 792
rect 456 783 458 792
rect 632 783 634 792
rect 800 783 802 792
rect 976 783 978 792
rect 1152 783 1154 792
rect 1328 783 1330 792
rect 1504 783 1506 792
rect 1824 783 1826 802
rect 1864 798 1866 813
rect 1888 808 1890 813
rect 2072 808 2074 813
rect 2264 808 2266 813
rect 2448 808 2450 813
rect 2624 808 2626 813
rect 2792 808 2794 813
rect 2944 808 2946 813
rect 3088 808 3090 813
rect 3224 808 3226 813
rect 3360 808 3362 813
rect 3480 808 3482 813
rect 1886 807 1892 808
rect 1886 803 1887 807
rect 1891 803 1892 807
rect 1886 802 1892 803
rect 2070 807 2076 808
rect 2070 803 2071 807
rect 2075 803 2076 807
rect 2070 802 2076 803
rect 2262 807 2268 808
rect 2262 803 2263 807
rect 2267 803 2268 807
rect 2262 802 2268 803
rect 2446 807 2452 808
rect 2446 803 2447 807
rect 2451 803 2452 807
rect 2446 802 2452 803
rect 2622 807 2628 808
rect 2622 803 2623 807
rect 2627 803 2628 807
rect 2622 802 2628 803
rect 2790 807 2796 808
rect 2790 803 2791 807
rect 2795 803 2796 807
rect 2790 802 2796 803
rect 2942 807 2948 808
rect 2942 803 2943 807
rect 2947 803 2948 807
rect 2942 802 2948 803
rect 3086 807 3092 808
rect 3086 803 3087 807
rect 3091 803 3092 807
rect 3086 802 3092 803
rect 3222 807 3228 808
rect 3222 803 3223 807
rect 3227 803 3228 807
rect 3222 802 3228 803
rect 3358 807 3364 808
rect 3358 803 3359 807
rect 3363 803 3364 807
rect 3358 802 3364 803
rect 3478 807 3484 808
rect 3478 803 3479 807
rect 3483 803 3484 807
rect 3478 802 3484 803
rect 3576 798 3578 813
rect 1862 797 1868 798
rect 1862 793 1863 797
rect 1867 793 1868 797
rect 1862 792 1868 793
rect 3574 797 3580 798
rect 3574 793 3575 797
rect 3579 793 3580 797
rect 3574 792 3580 793
rect 111 782 115 783
rect 111 777 115 778
rect 135 782 139 783
rect 135 777 139 778
rect 271 782 275 783
rect 271 777 275 778
rect 279 782 283 783
rect 279 777 283 778
rect 439 782 443 783
rect 439 777 443 778
rect 455 782 459 783
rect 455 777 459 778
rect 607 782 611 783
rect 607 777 611 778
rect 631 782 635 783
rect 631 777 635 778
rect 775 782 779 783
rect 775 777 779 778
rect 799 782 803 783
rect 799 777 803 778
rect 935 782 939 783
rect 935 777 939 778
rect 975 782 979 783
rect 975 777 979 778
rect 1087 782 1091 783
rect 1087 777 1091 778
rect 1151 782 1155 783
rect 1151 777 1155 778
rect 1239 782 1243 783
rect 1239 777 1243 778
rect 1327 782 1331 783
rect 1327 777 1331 778
rect 1391 782 1395 783
rect 1391 777 1395 778
rect 1503 782 1507 783
rect 1503 777 1507 778
rect 1551 782 1555 783
rect 1551 777 1555 778
rect 1823 782 1827 783
rect 1823 777 1827 778
rect 1862 780 1868 781
rect 112 762 114 777
rect 136 772 138 777
rect 272 772 274 777
rect 440 772 442 777
rect 608 772 610 777
rect 776 772 778 777
rect 936 772 938 777
rect 1088 772 1090 777
rect 1240 772 1242 777
rect 1392 772 1394 777
rect 1552 772 1554 777
rect 134 771 140 772
rect 134 767 135 771
rect 139 767 140 771
rect 134 766 140 767
rect 270 771 276 772
rect 270 767 271 771
rect 275 767 276 771
rect 270 766 276 767
rect 438 771 444 772
rect 438 767 439 771
rect 443 767 444 771
rect 438 766 444 767
rect 606 771 612 772
rect 606 767 607 771
rect 611 767 612 771
rect 606 766 612 767
rect 774 771 780 772
rect 774 767 775 771
rect 779 767 780 771
rect 774 766 780 767
rect 934 771 940 772
rect 934 767 935 771
rect 939 767 940 771
rect 934 766 940 767
rect 1086 771 1092 772
rect 1086 767 1087 771
rect 1091 767 1092 771
rect 1086 766 1092 767
rect 1238 771 1244 772
rect 1238 767 1239 771
rect 1243 767 1244 771
rect 1238 766 1244 767
rect 1390 771 1396 772
rect 1390 767 1391 771
rect 1395 767 1396 771
rect 1390 766 1396 767
rect 1550 771 1556 772
rect 1550 767 1551 771
rect 1555 767 1556 771
rect 1550 766 1556 767
rect 1824 762 1826 777
rect 1862 776 1863 780
rect 1867 776 1868 780
rect 1862 775 1868 776
rect 3574 780 3580 781
rect 3574 776 3575 780
rect 3579 776 3580 780
rect 3574 775 3580 776
rect 110 761 116 762
rect 110 757 111 761
rect 115 757 116 761
rect 110 756 116 757
rect 1822 761 1828 762
rect 1822 757 1823 761
rect 1827 757 1828 761
rect 1822 756 1828 757
rect 1864 751 1866 775
rect 1894 767 1900 768
rect 1894 763 1895 767
rect 1899 763 1900 767
rect 1894 762 1900 763
rect 2078 767 2084 768
rect 2078 763 2079 767
rect 2083 763 2084 767
rect 2078 762 2084 763
rect 2270 767 2276 768
rect 2270 763 2271 767
rect 2275 763 2276 767
rect 2270 762 2276 763
rect 2454 767 2460 768
rect 2454 763 2455 767
rect 2459 763 2460 767
rect 2454 762 2460 763
rect 2630 767 2636 768
rect 2630 763 2631 767
rect 2635 763 2636 767
rect 2630 762 2636 763
rect 2798 767 2804 768
rect 2798 763 2799 767
rect 2803 763 2804 767
rect 2798 762 2804 763
rect 2950 767 2956 768
rect 2950 763 2951 767
rect 2955 763 2956 767
rect 2950 762 2956 763
rect 3094 767 3100 768
rect 3094 763 3095 767
rect 3099 763 3100 767
rect 3094 762 3100 763
rect 3230 767 3236 768
rect 3230 763 3231 767
rect 3235 763 3236 767
rect 3230 762 3236 763
rect 3366 767 3372 768
rect 3366 763 3367 767
rect 3371 763 3372 767
rect 3366 762 3372 763
rect 3486 767 3492 768
rect 3486 763 3487 767
rect 3491 763 3492 767
rect 3486 762 3492 763
rect 1896 751 1898 762
rect 2080 751 2082 762
rect 2272 751 2274 762
rect 2456 751 2458 762
rect 2632 751 2634 762
rect 2800 751 2802 762
rect 2952 751 2954 762
rect 3096 751 3098 762
rect 3232 751 3234 762
rect 3368 751 3370 762
rect 3488 751 3490 762
rect 3576 751 3578 775
rect 1863 750 1867 751
rect 1863 745 1867 746
rect 1895 750 1899 751
rect 1895 745 1899 746
rect 2071 750 2075 751
rect 2071 745 2075 746
rect 2079 750 2083 751
rect 2079 745 2083 746
rect 2263 750 2267 751
rect 2263 745 2267 746
rect 2271 750 2275 751
rect 2271 745 2275 746
rect 2447 750 2451 751
rect 2447 745 2451 746
rect 2455 750 2459 751
rect 2455 745 2459 746
rect 2623 750 2627 751
rect 2623 745 2627 746
rect 2631 750 2635 751
rect 2631 745 2635 746
rect 2799 750 2803 751
rect 2799 745 2803 746
rect 2951 750 2955 751
rect 2951 745 2955 746
rect 2975 750 2979 751
rect 2975 745 2979 746
rect 3095 750 3099 751
rect 3095 745 3099 746
rect 3151 750 3155 751
rect 3151 745 3155 746
rect 3231 750 3235 751
rect 3231 745 3235 746
rect 3327 750 3331 751
rect 3327 745 3331 746
rect 3367 750 3371 751
rect 3367 745 3371 746
rect 3487 750 3491 751
rect 3487 745 3491 746
rect 3575 750 3579 751
rect 3575 745 3579 746
rect 110 744 116 745
rect 110 740 111 744
rect 115 740 116 744
rect 110 739 116 740
rect 1822 744 1828 745
rect 1822 740 1823 744
rect 1827 740 1828 744
rect 1822 739 1828 740
rect 112 711 114 739
rect 142 731 148 732
rect 142 727 143 731
rect 147 727 148 731
rect 142 726 148 727
rect 278 731 284 732
rect 278 727 279 731
rect 283 727 284 731
rect 278 726 284 727
rect 446 731 452 732
rect 446 727 447 731
rect 451 727 452 731
rect 446 726 452 727
rect 614 731 620 732
rect 614 727 615 731
rect 619 727 620 731
rect 614 726 620 727
rect 782 731 788 732
rect 782 727 783 731
rect 787 727 788 731
rect 782 726 788 727
rect 942 731 948 732
rect 942 727 943 731
rect 947 727 948 731
rect 942 726 948 727
rect 1094 731 1100 732
rect 1094 727 1095 731
rect 1099 727 1100 731
rect 1094 726 1100 727
rect 1246 731 1252 732
rect 1246 727 1247 731
rect 1251 727 1252 731
rect 1246 726 1252 727
rect 1398 731 1404 732
rect 1398 727 1399 731
rect 1403 727 1404 731
rect 1398 726 1404 727
rect 1558 731 1564 732
rect 1558 727 1559 731
rect 1563 727 1564 731
rect 1558 726 1564 727
rect 144 711 146 726
rect 280 711 282 726
rect 448 711 450 726
rect 616 711 618 726
rect 784 711 786 726
rect 944 711 946 726
rect 1096 711 1098 726
rect 1248 711 1250 726
rect 1400 711 1402 726
rect 1560 711 1562 726
rect 1824 711 1826 739
rect 1864 721 1866 745
rect 1896 734 1898 745
rect 2072 734 2074 745
rect 2264 734 2266 745
rect 2448 734 2450 745
rect 2624 734 2626 745
rect 2800 734 2802 745
rect 2976 734 2978 745
rect 3152 734 3154 745
rect 3328 734 3330 745
rect 3488 734 3490 745
rect 1894 733 1900 734
rect 1894 729 1895 733
rect 1899 729 1900 733
rect 1894 728 1900 729
rect 2070 733 2076 734
rect 2070 729 2071 733
rect 2075 729 2076 733
rect 2070 728 2076 729
rect 2262 733 2268 734
rect 2262 729 2263 733
rect 2267 729 2268 733
rect 2262 728 2268 729
rect 2446 733 2452 734
rect 2446 729 2447 733
rect 2451 729 2452 733
rect 2446 728 2452 729
rect 2622 733 2628 734
rect 2622 729 2623 733
rect 2627 729 2628 733
rect 2622 728 2628 729
rect 2798 733 2804 734
rect 2798 729 2799 733
rect 2803 729 2804 733
rect 2798 728 2804 729
rect 2974 733 2980 734
rect 2974 729 2975 733
rect 2979 729 2980 733
rect 2974 728 2980 729
rect 3150 733 3156 734
rect 3150 729 3151 733
rect 3155 729 3156 733
rect 3150 728 3156 729
rect 3326 733 3332 734
rect 3326 729 3327 733
rect 3331 729 3332 733
rect 3326 728 3332 729
rect 3486 733 3492 734
rect 3486 729 3487 733
rect 3491 729 3492 733
rect 3486 728 3492 729
rect 3576 721 3578 745
rect 1862 720 1868 721
rect 1862 716 1863 720
rect 1867 716 1868 720
rect 1862 715 1868 716
rect 3574 720 3580 721
rect 3574 716 3575 720
rect 3579 716 3580 720
rect 3574 715 3580 716
rect 111 710 115 711
rect 111 705 115 706
rect 143 710 147 711
rect 143 705 147 706
rect 279 710 283 711
rect 279 705 283 706
rect 287 710 291 711
rect 287 705 291 706
rect 447 710 451 711
rect 447 705 451 706
rect 455 710 459 711
rect 455 705 459 706
rect 615 710 619 711
rect 615 705 619 706
rect 623 710 627 711
rect 623 705 627 706
rect 783 710 787 711
rect 783 705 787 706
rect 791 710 795 711
rect 791 705 795 706
rect 943 710 947 711
rect 943 705 947 706
rect 959 710 963 711
rect 959 705 963 706
rect 1095 710 1099 711
rect 1095 705 1099 706
rect 1119 710 1123 711
rect 1119 705 1123 706
rect 1247 710 1251 711
rect 1247 705 1251 706
rect 1279 710 1283 711
rect 1279 705 1283 706
rect 1399 710 1403 711
rect 1399 705 1403 706
rect 1439 710 1443 711
rect 1439 705 1443 706
rect 1559 710 1563 711
rect 1559 705 1563 706
rect 1599 710 1603 711
rect 1599 705 1603 706
rect 1823 710 1827 711
rect 1823 705 1827 706
rect 112 681 114 705
rect 144 694 146 705
rect 288 694 290 705
rect 456 694 458 705
rect 624 694 626 705
rect 792 694 794 705
rect 960 694 962 705
rect 1120 694 1122 705
rect 1280 694 1282 705
rect 1440 694 1442 705
rect 1600 694 1602 705
rect 142 693 148 694
rect 142 689 143 693
rect 147 689 148 693
rect 142 688 148 689
rect 286 693 292 694
rect 286 689 287 693
rect 291 689 292 693
rect 286 688 292 689
rect 454 693 460 694
rect 454 689 455 693
rect 459 689 460 693
rect 454 688 460 689
rect 622 693 628 694
rect 622 689 623 693
rect 627 689 628 693
rect 622 688 628 689
rect 790 693 796 694
rect 790 689 791 693
rect 795 689 796 693
rect 790 688 796 689
rect 958 693 964 694
rect 958 689 959 693
rect 963 689 964 693
rect 958 688 964 689
rect 1118 693 1124 694
rect 1118 689 1119 693
rect 1123 689 1124 693
rect 1118 688 1124 689
rect 1278 693 1284 694
rect 1278 689 1279 693
rect 1283 689 1284 693
rect 1278 688 1284 689
rect 1438 693 1444 694
rect 1438 689 1439 693
rect 1443 689 1444 693
rect 1438 688 1444 689
rect 1598 693 1604 694
rect 1598 689 1599 693
rect 1603 689 1604 693
rect 1598 688 1604 689
rect 1824 681 1826 705
rect 1862 703 1868 704
rect 1862 699 1863 703
rect 1867 699 1868 703
rect 1862 698 1868 699
rect 3574 703 3580 704
rect 3574 699 3575 703
rect 3579 699 3580 703
rect 3574 698 3580 699
rect 110 680 116 681
rect 110 676 111 680
rect 115 676 116 680
rect 110 675 116 676
rect 1822 680 1828 681
rect 1822 676 1823 680
rect 1827 676 1828 680
rect 1864 679 1866 698
rect 1886 693 1892 694
rect 1886 689 1887 693
rect 1891 689 1892 693
rect 1886 688 1892 689
rect 2062 693 2068 694
rect 2062 689 2063 693
rect 2067 689 2068 693
rect 2062 688 2068 689
rect 2254 693 2260 694
rect 2254 689 2255 693
rect 2259 689 2260 693
rect 2254 688 2260 689
rect 2438 693 2444 694
rect 2438 689 2439 693
rect 2443 689 2444 693
rect 2438 688 2444 689
rect 2614 693 2620 694
rect 2614 689 2615 693
rect 2619 689 2620 693
rect 2614 688 2620 689
rect 2790 693 2796 694
rect 2790 689 2791 693
rect 2795 689 2796 693
rect 2790 688 2796 689
rect 2966 693 2972 694
rect 2966 689 2967 693
rect 2971 689 2972 693
rect 2966 688 2972 689
rect 3142 693 3148 694
rect 3142 689 3143 693
rect 3147 689 3148 693
rect 3142 688 3148 689
rect 3318 693 3324 694
rect 3318 689 3319 693
rect 3323 689 3324 693
rect 3318 688 3324 689
rect 3478 693 3484 694
rect 3478 689 3479 693
rect 3483 689 3484 693
rect 3478 688 3484 689
rect 1888 679 1890 688
rect 2064 679 2066 688
rect 2256 679 2258 688
rect 2440 679 2442 688
rect 2616 679 2618 688
rect 2792 679 2794 688
rect 2968 679 2970 688
rect 3144 679 3146 688
rect 3320 679 3322 688
rect 3480 679 3482 688
rect 3576 679 3578 698
rect 1822 675 1828 676
rect 1863 678 1867 679
rect 1863 673 1867 674
rect 1887 678 1891 679
rect 1887 673 1891 674
rect 1975 678 1979 679
rect 1975 673 1979 674
rect 2063 678 2067 679
rect 2063 673 2067 674
rect 2095 678 2099 679
rect 2095 673 2099 674
rect 2223 678 2227 679
rect 2223 673 2227 674
rect 2255 678 2259 679
rect 2255 673 2259 674
rect 2351 678 2355 679
rect 2351 673 2355 674
rect 2439 678 2443 679
rect 2439 673 2443 674
rect 2479 678 2483 679
rect 2479 673 2483 674
rect 2615 678 2619 679
rect 2615 673 2619 674
rect 2767 678 2771 679
rect 2767 673 2771 674
rect 2791 678 2795 679
rect 2791 673 2795 674
rect 2935 678 2939 679
rect 2935 673 2939 674
rect 2967 678 2971 679
rect 2967 673 2971 674
rect 3119 678 3123 679
rect 3119 673 3123 674
rect 3143 678 3147 679
rect 3143 673 3147 674
rect 3311 678 3315 679
rect 3311 673 3315 674
rect 3319 678 3323 679
rect 3319 673 3323 674
rect 3479 678 3483 679
rect 3479 673 3483 674
rect 3575 678 3579 679
rect 3575 673 3579 674
rect 110 663 116 664
rect 110 659 111 663
rect 115 659 116 663
rect 110 658 116 659
rect 1822 663 1828 664
rect 1822 659 1823 663
rect 1827 659 1828 663
rect 1822 658 1828 659
rect 1864 658 1866 673
rect 1888 668 1890 673
rect 1976 668 1978 673
rect 2096 668 2098 673
rect 2224 668 2226 673
rect 2352 668 2354 673
rect 2480 668 2482 673
rect 2616 668 2618 673
rect 2768 668 2770 673
rect 2936 668 2938 673
rect 3120 668 3122 673
rect 3312 668 3314 673
rect 3480 668 3482 673
rect 1886 667 1892 668
rect 1886 663 1887 667
rect 1891 663 1892 667
rect 1886 662 1892 663
rect 1974 667 1980 668
rect 1974 663 1975 667
rect 1979 663 1980 667
rect 1974 662 1980 663
rect 2094 667 2100 668
rect 2094 663 2095 667
rect 2099 663 2100 667
rect 2094 662 2100 663
rect 2222 667 2228 668
rect 2222 663 2223 667
rect 2227 663 2228 667
rect 2222 662 2228 663
rect 2350 667 2356 668
rect 2350 663 2351 667
rect 2355 663 2356 667
rect 2350 662 2356 663
rect 2478 667 2484 668
rect 2478 663 2479 667
rect 2483 663 2484 667
rect 2478 662 2484 663
rect 2614 667 2620 668
rect 2614 663 2615 667
rect 2619 663 2620 667
rect 2614 662 2620 663
rect 2766 667 2772 668
rect 2766 663 2767 667
rect 2771 663 2772 667
rect 2766 662 2772 663
rect 2934 667 2940 668
rect 2934 663 2935 667
rect 2939 663 2940 667
rect 2934 662 2940 663
rect 3118 667 3124 668
rect 3118 663 3119 667
rect 3123 663 3124 667
rect 3118 662 3124 663
rect 3310 667 3316 668
rect 3310 663 3311 667
rect 3315 663 3316 667
rect 3310 662 3316 663
rect 3478 667 3484 668
rect 3478 663 3479 667
rect 3483 663 3484 667
rect 3478 662 3484 663
rect 3576 658 3578 673
rect 112 635 114 658
rect 134 653 140 654
rect 134 649 135 653
rect 139 649 140 653
rect 134 648 140 649
rect 278 653 284 654
rect 278 649 279 653
rect 283 649 284 653
rect 278 648 284 649
rect 446 653 452 654
rect 446 649 447 653
rect 451 649 452 653
rect 446 648 452 649
rect 614 653 620 654
rect 614 649 615 653
rect 619 649 620 653
rect 614 648 620 649
rect 782 653 788 654
rect 782 649 783 653
rect 787 649 788 653
rect 782 648 788 649
rect 950 653 956 654
rect 950 649 951 653
rect 955 649 956 653
rect 950 648 956 649
rect 1110 653 1116 654
rect 1110 649 1111 653
rect 1115 649 1116 653
rect 1110 648 1116 649
rect 1270 653 1276 654
rect 1270 649 1271 653
rect 1275 649 1276 653
rect 1270 648 1276 649
rect 1430 653 1436 654
rect 1430 649 1431 653
rect 1435 649 1436 653
rect 1430 648 1436 649
rect 1590 653 1596 654
rect 1590 649 1591 653
rect 1595 649 1596 653
rect 1590 648 1596 649
rect 136 635 138 648
rect 280 635 282 648
rect 448 635 450 648
rect 616 635 618 648
rect 784 635 786 648
rect 952 635 954 648
rect 1112 635 1114 648
rect 1272 635 1274 648
rect 1432 635 1434 648
rect 1592 635 1594 648
rect 1824 635 1826 658
rect 1862 657 1868 658
rect 1862 653 1863 657
rect 1867 653 1868 657
rect 1862 652 1868 653
rect 3574 657 3580 658
rect 3574 653 3575 657
rect 3579 653 3580 657
rect 3574 652 3580 653
rect 1862 640 1868 641
rect 1862 636 1863 640
rect 1867 636 1868 640
rect 1862 635 1868 636
rect 3574 640 3580 641
rect 3574 636 3575 640
rect 3579 636 3580 640
rect 3574 635 3580 636
rect 111 634 115 635
rect 111 629 115 630
rect 135 634 139 635
rect 135 629 139 630
rect 279 634 283 635
rect 279 629 283 630
rect 287 634 291 635
rect 287 629 291 630
rect 447 634 451 635
rect 447 629 451 630
rect 455 634 459 635
rect 455 629 459 630
rect 615 634 619 635
rect 615 629 619 630
rect 631 634 635 635
rect 631 629 635 630
rect 783 634 787 635
rect 783 629 787 630
rect 799 634 803 635
rect 799 629 803 630
rect 951 634 955 635
rect 951 629 955 630
rect 967 634 971 635
rect 967 629 971 630
rect 1111 634 1115 635
rect 1111 629 1115 630
rect 1119 634 1123 635
rect 1119 629 1123 630
rect 1271 634 1275 635
rect 1271 629 1275 630
rect 1415 634 1419 635
rect 1415 629 1419 630
rect 1431 634 1435 635
rect 1431 629 1435 630
rect 1559 634 1563 635
rect 1559 629 1563 630
rect 1591 634 1595 635
rect 1591 629 1595 630
rect 1711 634 1715 635
rect 1711 629 1715 630
rect 1823 634 1827 635
rect 1823 629 1827 630
rect 112 614 114 629
rect 136 624 138 629
rect 288 624 290 629
rect 456 624 458 629
rect 632 624 634 629
rect 800 624 802 629
rect 968 624 970 629
rect 1120 624 1122 629
rect 1272 624 1274 629
rect 1416 624 1418 629
rect 1560 624 1562 629
rect 1712 624 1714 629
rect 134 623 140 624
rect 134 619 135 623
rect 139 619 140 623
rect 134 618 140 619
rect 286 623 292 624
rect 286 619 287 623
rect 291 619 292 623
rect 286 618 292 619
rect 454 623 460 624
rect 454 619 455 623
rect 459 619 460 623
rect 454 618 460 619
rect 630 623 636 624
rect 630 619 631 623
rect 635 619 636 623
rect 630 618 636 619
rect 798 623 804 624
rect 798 619 799 623
rect 803 619 804 623
rect 798 618 804 619
rect 966 623 972 624
rect 966 619 967 623
rect 971 619 972 623
rect 966 618 972 619
rect 1118 623 1124 624
rect 1118 619 1119 623
rect 1123 619 1124 623
rect 1118 618 1124 619
rect 1270 623 1276 624
rect 1270 619 1271 623
rect 1275 619 1276 623
rect 1270 618 1276 619
rect 1414 623 1420 624
rect 1414 619 1415 623
rect 1419 619 1420 623
rect 1414 618 1420 619
rect 1558 623 1564 624
rect 1558 619 1559 623
rect 1563 619 1564 623
rect 1558 618 1564 619
rect 1710 623 1716 624
rect 1710 619 1711 623
rect 1715 619 1716 623
rect 1710 618 1716 619
rect 1824 614 1826 629
rect 110 613 116 614
rect 110 609 111 613
rect 115 609 116 613
rect 110 608 116 609
rect 1822 613 1828 614
rect 1822 609 1823 613
rect 1827 609 1828 613
rect 1822 608 1828 609
rect 1864 607 1866 635
rect 1894 627 1900 628
rect 1894 623 1895 627
rect 1899 623 1900 627
rect 1894 622 1900 623
rect 1982 627 1988 628
rect 1982 623 1983 627
rect 1987 623 1988 627
rect 1982 622 1988 623
rect 2102 627 2108 628
rect 2102 623 2103 627
rect 2107 623 2108 627
rect 2102 622 2108 623
rect 2230 627 2236 628
rect 2230 623 2231 627
rect 2235 623 2236 627
rect 2230 622 2236 623
rect 2358 627 2364 628
rect 2358 623 2359 627
rect 2363 623 2364 627
rect 2358 622 2364 623
rect 2486 627 2492 628
rect 2486 623 2487 627
rect 2491 623 2492 627
rect 2486 622 2492 623
rect 2622 627 2628 628
rect 2622 623 2623 627
rect 2627 623 2628 627
rect 2622 622 2628 623
rect 2774 627 2780 628
rect 2774 623 2775 627
rect 2779 623 2780 627
rect 2774 622 2780 623
rect 2942 627 2948 628
rect 2942 623 2943 627
rect 2947 623 2948 627
rect 2942 622 2948 623
rect 3126 627 3132 628
rect 3126 623 3127 627
rect 3131 623 3132 627
rect 3126 622 3132 623
rect 3318 627 3324 628
rect 3318 623 3319 627
rect 3323 623 3324 627
rect 3318 622 3324 623
rect 3486 627 3492 628
rect 3486 623 3487 627
rect 3491 623 3492 627
rect 3486 622 3492 623
rect 1896 607 1898 622
rect 1984 607 1986 622
rect 2104 607 2106 622
rect 2232 607 2234 622
rect 2360 607 2362 622
rect 2488 607 2490 622
rect 2624 607 2626 622
rect 2776 607 2778 622
rect 2944 607 2946 622
rect 3128 607 3130 622
rect 3320 607 3322 622
rect 3488 607 3490 622
rect 3576 607 3578 635
rect 1863 606 1867 607
rect 1863 601 1867 602
rect 1895 606 1899 607
rect 1895 601 1899 602
rect 1983 606 1987 607
rect 1983 601 1987 602
rect 2047 606 2051 607
rect 2047 601 2051 602
rect 2103 606 2107 607
rect 2103 601 2107 602
rect 2215 606 2219 607
rect 2215 601 2219 602
rect 2231 606 2235 607
rect 2231 601 2235 602
rect 2359 606 2363 607
rect 2359 601 2363 602
rect 2391 606 2395 607
rect 2391 601 2395 602
rect 2487 606 2491 607
rect 2487 601 2491 602
rect 2583 606 2587 607
rect 2583 601 2587 602
rect 2623 606 2627 607
rect 2623 601 2627 602
rect 2775 606 2779 607
rect 2775 601 2779 602
rect 2799 606 2803 607
rect 2799 601 2803 602
rect 2943 606 2947 607
rect 2943 601 2947 602
rect 3023 606 3027 607
rect 3023 601 3027 602
rect 3127 606 3131 607
rect 3127 601 3131 602
rect 3255 606 3259 607
rect 3255 601 3259 602
rect 3319 606 3323 607
rect 3319 601 3323 602
rect 3487 606 3491 607
rect 3487 601 3491 602
rect 3575 606 3579 607
rect 3575 601 3579 602
rect 110 596 116 597
rect 110 592 111 596
rect 115 592 116 596
rect 110 591 116 592
rect 1822 596 1828 597
rect 1822 592 1823 596
rect 1827 592 1828 596
rect 1822 591 1828 592
rect 112 563 114 591
rect 142 583 148 584
rect 142 579 143 583
rect 147 579 148 583
rect 142 578 148 579
rect 294 583 300 584
rect 294 579 295 583
rect 299 579 300 583
rect 294 578 300 579
rect 462 583 468 584
rect 462 579 463 583
rect 467 579 468 583
rect 462 578 468 579
rect 638 583 644 584
rect 638 579 639 583
rect 643 579 644 583
rect 638 578 644 579
rect 806 583 812 584
rect 806 579 807 583
rect 811 579 812 583
rect 806 578 812 579
rect 974 583 980 584
rect 974 579 975 583
rect 979 579 980 583
rect 974 578 980 579
rect 1126 583 1132 584
rect 1126 579 1127 583
rect 1131 579 1132 583
rect 1126 578 1132 579
rect 1278 583 1284 584
rect 1278 579 1279 583
rect 1283 579 1284 583
rect 1278 578 1284 579
rect 1422 583 1428 584
rect 1422 579 1423 583
rect 1427 579 1428 583
rect 1422 578 1428 579
rect 1566 583 1572 584
rect 1566 579 1567 583
rect 1571 579 1572 583
rect 1566 578 1572 579
rect 1718 583 1724 584
rect 1718 579 1719 583
rect 1723 579 1724 583
rect 1718 578 1724 579
rect 144 563 146 578
rect 296 563 298 578
rect 464 563 466 578
rect 640 563 642 578
rect 808 563 810 578
rect 976 563 978 578
rect 1128 563 1130 578
rect 1280 563 1282 578
rect 1424 563 1426 578
rect 1568 563 1570 578
rect 1720 563 1722 578
rect 1824 563 1826 591
rect 1864 577 1866 601
rect 1896 590 1898 601
rect 2048 590 2050 601
rect 2216 590 2218 601
rect 2392 590 2394 601
rect 2584 590 2586 601
rect 2800 590 2802 601
rect 3024 590 3026 601
rect 3256 590 3258 601
rect 3488 590 3490 601
rect 1894 589 1900 590
rect 1894 585 1895 589
rect 1899 585 1900 589
rect 1894 584 1900 585
rect 2046 589 2052 590
rect 2046 585 2047 589
rect 2051 585 2052 589
rect 2046 584 2052 585
rect 2214 589 2220 590
rect 2214 585 2215 589
rect 2219 585 2220 589
rect 2214 584 2220 585
rect 2390 589 2396 590
rect 2390 585 2391 589
rect 2395 585 2396 589
rect 2390 584 2396 585
rect 2582 589 2588 590
rect 2582 585 2583 589
rect 2587 585 2588 589
rect 2582 584 2588 585
rect 2798 589 2804 590
rect 2798 585 2799 589
rect 2803 585 2804 589
rect 2798 584 2804 585
rect 3022 589 3028 590
rect 3022 585 3023 589
rect 3027 585 3028 589
rect 3022 584 3028 585
rect 3254 589 3260 590
rect 3254 585 3255 589
rect 3259 585 3260 589
rect 3254 584 3260 585
rect 3486 589 3492 590
rect 3486 585 3487 589
rect 3491 585 3492 589
rect 3486 584 3492 585
rect 3576 577 3578 601
rect 1862 576 1868 577
rect 1862 572 1863 576
rect 1867 572 1868 576
rect 1862 571 1868 572
rect 3574 576 3580 577
rect 3574 572 3575 576
rect 3579 572 3580 576
rect 3574 571 3580 572
rect 111 562 115 563
rect 111 557 115 558
rect 143 562 147 563
rect 143 557 147 558
rect 151 562 155 563
rect 151 557 155 558
rect 295 562 299 563
rect 295 557 299 558
rect 311 562 315 563
rect 311 557 315 558
rect 463 562 467 563
rect 463 557 467 558
rect 471 562 475 563
rect 471 557 475 558
rect 631 562 635 563
rect 631 557 635 558
rect 639 562 643 563
rect 639 557 643 558
rect 783 562 787 563
rect 783 557 787 558
rect 807 562 811 563
rect 807 557 811 558
rect 927 562 931 563
rect 927 557 931 558
rect 975 562 979 563
rect 975 557 979 558
rect 1063 562 1067 563
rect 1063 557 1067 558
rect 1127 562 1131 563
rect 1127 557 1131 558
rect 1191 562 1195 563
rect 1191 557 1195 558
rect 1279 562 1283 563
rect 1279 557 1283 558
rect 1311 562 1315 563
rect 1311 557 1315 558
rect 1423 562 1427 563
rect 1423 557 1427 558
rect 1535 562 1539 563
rect 1535 557 1539 558
rect 1567 562 1571 563
rect 1567 557 1571 558
rect 1647 562 1651 563
rect 1647 557 1651 558
rect 1719 562 1723 563
rect 1719 557 1723 558
rect 1735 562 1739 563
rect 1735 557 1739 558
rect 1823 562 1827 563
rect 1823 557 1827 558
rect 1862 559 1868 560
rect 112 533 114 557
rect 152 546 154 557
rect 312 546 314 557
rect 472 546 474 557
rect 632 546 634 557
rect 784 546 786 557
rect 928 546 930 557
rect 1064 546 1066 557
rect 1192 546 1194 557
rect 1312 546 1314 557
rect 1424 546 1426 557
rect 1536 546 1538 557
rect 1648 546 1650 557
rect 1736 546 1738 557
rect 150 545 156 546
rect 150 541 151 545
rect 155 541 156 545
rect 150 540 156 541
rect 310 545 316 546
rect 310 541 311 545
rect 315 541 316 545
rect 310 540 316 541
rect 470 545 476 546
rect 470 541 471 545
rect 475 541 476 545
rect 470 540 476 541
rect 630 545 636 546
rect 630 541 631 545
rect 635 541 636 545
rect 630 540 636 541
rect 782 545 788 546
rect 782 541 783 545
rect 787 541 788 545
rect 782 540 788 541
rect 926 545 932 546
rect 926 541 927 545
rect 931 541 932 545
rect 926 540 932 541
rect 1062 545 1068 546
rect 1062 541 1063 545
rect 1067 541 1068 545
rect 1062 540 1068 541
rect 1190 545 1196 546
rect 1190 541 1191 545
rect 1195 541 1196 545
rect 1190 540 1196 541
rect 1310 545 1316 546
rect 1310 541 1311 545
rect 1315 541 1316 545
rect 1310 540 1316 541
rect 1422 545 1428 546
rect 1422 541 1423 545
rect 1427 541 1428 545
rect 1422 540 1428 541
rect 1534 545 1540 546
rect 1534 541 1535 545
rect 1539 541 1540 545
rect 1534 540 1540 541
rect 1646 545 1652 546
rect 1646 541 1647 545
rect 1651 541 1652 545
rect 1646 540 1652 541
rect 1734 545 1740 546
rect 1734 541 1735 545
rect 1739 541 1740 545
rect 1734 540 1740 541
rect 1824 533 1826 557
rect 1862 555 1863 559
rect 1867 555 1868 559
rect 1862 554 1868 555
rect 3574 559 3580 560
rect 3574 555 3575 559
rect 3579 555 3580 559
rect 3574 554 3580 555
rect 110 532 116 533
rect 110 528 111 532
rect 115 528 116 532
rect 110 527 116 528
rect 1822 532 1828 533
rect 1822 528 1823 532
rect 1827 528 1828 532
rect 1864 531 1866 554
rect 1886 549 1892 550
rect 1886 545 1887 549
rect 1891 545 1892 549
rect 1886 544 1892 545
rect 2038 549 2044 550
rect 2038 545 2039 549
rect 2043 545 2044 549
rect 2038 544 2044 545
rect 2206 549 2212 550
rect 2206 545 2207 549
rect 2211 545 2212 549
rect 2206 544 2212 545
rect 2382 549 2388 550
rect 2382 545 2383 549
rect 2387 545 2388 549
rect 2382 544 2388 545
rect 2574 549 2580 550
rect 2574 545 2575 549
rect 2579 545 2580 549
rect 2574 544 2580 545
rect 2790 549 2796 550
rect 2790 545 2791 549
rect 2795 545 2796 549
rect 2790 544 2796 545
rect 3014 549 3020 550
rect 3014 545 3015 549
rect 3019 545 3020 549
rect 3014 544 3020 545
rect 3246 549 3252 550
rect 3246 545 3247 549
rect 3251 545 3252 549
rect 3246 544 3252 545
rect 3478 549 3484 550
rect 3478 545 3479 549
rect 3483 545 3484 549
rect 3478 544 3484 545
rect 1888 531 1890 544
rect 2040 531 2042 544
rect 2208 531 2210 544
rect 2384 531 2386 544
rect 2576 531 2578 544
rect 2792 531 2794 544
rect 3016 531 3018 544
rect 3248 531 3250 544
rect 3480 531 3482 544
rect 3576 531 3578 554
rect 1822 527 1828 528
rect 1863 530 1867 531
rect 1863 525 1867 526
rect 1887 530 1891 531
rect 1887 525 1891 526
rect 2039 530 2043 531
rect 2039 525 2043 526
rect 2191 530 2195 531
rect 2191 525 2195 526
rect 2207 530 2211 531
rect 2207 525 2211 526
rect 2279 530 2283 531
rect 2279 525 2283 526
rect 2375 530 2379 531
rect 2375 525 2379 526
rect 2383 530 2387 531
rect 2383 525 2387 526
rect 2487 530 2491 531
rect 2487 525 2491 526
rect 2575 530 2579 531
rect 2575 525 2579 526
rect 2631 530 2635 531
rect 2631 525 2635 526
rect 2791 530 2795 531
rect 2791 525 2795 526
rect 2807 530 2811 531
rect 2807 525 2811 526
rect 3007 530 3011 531
rect 3007 525 3011 526
rect 3015 530 3019 531
rect 3015 525 3019 526
rect 3215 530 3219 531
rect 3215 525 3219 526
rect 3247 530 3251 531
rect 3247 525 3251 526
rect 3431 530 3435 531
rect 3431 525 3435 526
rect 3479 530 3483 531
rect 3479 525 3483 526
rect 3575 530 3579 531
rect 3575 525 3579 526
rect 110 515 116 516
rect 110 511 111 515
rect 115 511 116 515
rect 110 510 116 511
rect 1822 515 1828 516
rect 1822 511 1823 515
rect 1827 511 1828 515
rect 1822 510 1828 511
rect 1864 510 1866 525
rect 2192 520 2194 525
rect 2280 520 2282 525
rect 2376 520 2378 525
rect 2488 520 2490 525
rect 2632 520 2634 525
rect 2808 520 2810 525
rect 3008 520 3010 525
rect 3216 520 3218 525
rect 3432 520 3434 525
rect 2190 519 2196 520
rect 2190 515 2191 519
rect 2195 515 2196 519
rect 2190 514 2196 515
rect 2278 519 2284 520
rect 2278 515 2279 519
rect 2283 515 2284 519
rect 2278 514 2284 515
rect 2374 519 2380 520
rect 2374 515 2375 519
rect 2379 515 2380 519
rect 2374 514 2380 515
rect 2486 519 2492 520
rect 2486 515 2487 519
rect 2491 515 2492 519
rect 2486 514 2492 515
rect 2630 519 2636 520
rect 2630 515 2631 519
rect 2635 515 2636 519
rect 2630 514 2636 515
rect 2806 519 2812 520
rect 2806 515 2807 519
rect 2811 515 2812 519
rect 2806 514 2812 515
rect 3006 519 3012 520
rect 3006 515 3007 519
rect 3011 515 3012 519
rect 3006 514 3012 515
rect 3214 519 3220 520
rect 3214 515 3215 519
rect 3219 515 3220 519
rect 3214 514 3220 515
rect 3430 519 3436 520
rect 3430 515 3431 519
rect 3435 515 3436 519
rect 3430 514 3436 515
rect 3576 510 3578 525
rect 112 487 114 510
rect 142 505 148 506
rect 142 501 143 505
rect 147 501 148 505
rect 142 500 148 501
rect 302 505 308 506
rect 302 501 303 505
rect 307 501 308 505
rect 302 500 308 501
rect 462 505 468 506
rect 462 501 463 505
rect 467 501 468 505
rect 462 500 468 501
rect 622 505 628 506
rect 622 501 623 505
rect 627 501 628 505
rect 622 500 628 501
rect 774 505 780 506
rect 774 501 775 505
rect 779 501 780 505
rect 774 500 780 501
rect 918 505 924 506
rect 918 501 919 505
rect 923 501 924 505
rect 918 500 924 501
rect 1054 505 1060 506
rect 1054 501 1055 505
rect 1059 501 1060 505
rect 1054 500 1060 501
rect 1182 505 1188 506
rect 1182 501 1183 505
rect 1187 501 1188 505
rect 1182 500 1188 501
rect 1302 505 1308 506
rect 1302 501 1303 505
rect 1307 501 1308 505
rect 1302 500 1308 501
rect 1414 505 1420 506
rect 1414 501 1415 505
rect 1419 501 1420 505
rect 1414 500 1420 501
rect 1526 505 1532 506
rect 1526 501 1527 505
rect 1531 501 1532 505
rect 1526 500 1532 501
rect 1638 505 1644 506
rect 1638 501 1639 505
rect 1643 501 1644 505
rect 1638 500 1644 501
rect 1726 505 1732 506
rect 1726 501 1727 505
rect 1731 501 1732 505
rect 1726 500 1732 501
rect 144 487 146 500
rect 304 487 306 500
rect 464 487 466 500
rect 624 487 626 500
rect 776 487 778 500
rect 920 487 922 500
rect 1056 487 1058 500
rect 1184 487 1186 500
rect 1304 487 1306 500
rect 1416 487 1418 500
rect 1528 487 1530 500
rect 1640 487 1642 500
rect 1728 487 1730 500
rect 1824 487 1826 510
rect 1862 509 1868 510
rect 1862 505 1863 509
rect 1867 505 1868 509
rect 1862 504 1868 505
rect 3574 509 3580 510
rect 3574 505 3575 509
rect 3579 505 3580 509
rect 3574 504 3580 505
rect 1862 492 1868 493
rect 1862 488 1863 492
rect 1867 488 1868 492
rect 1862 487 1868 488
rect 3574 492 3580 493
rect 3574 488 3575 492
rect 3579 488 3580 492
rect 3574 487 3580 488
rect 111 486 115 487
rect 111 481 115 482
rect 143 486 147 487
rect 143 481 147 482
rect 159 486 163 487
rect 159 481 163 482
rect 303 486 307 487
rect 303 481 307 482
rect 311 486 315 487
rect 311 481 315 482
rect 463 486 467 487
rect 463 481 467 482
rect 615 486 619 487
rect 615 481 619 482
rect 623 486 627 487
rect 623 481 627 482
rect 759 486 763 487
rect 759 481 763 482
rect 775 486 779 487
rect 775 481 779 482
rect 887 486 891 487
rect 887 481 891 482
rect 919 486 923 487
rect 919 481 923 482
rect 1007 486 1011 487
rect 1007 481 1011 482
rect 1055 486 1059 487
rect 1055 481 1059 482
rect 1127 486 1131 487
rect 1127 481 1131 482
rect 1183 486 1187 487
rect 1183 481 1187 482
rect 1239 486 1243 487
rect 1239 481 1243 482
rect 1303 486 1307 487
rect 1303 481 1307 482
rect 1343 486 1347 487
rect 1343 481 1347 482
rect 1415 486 1419 487
rect 1415 481 1419 482
rect 1439 486 1443 487
rect 1439 481 1443 482
rect 1527 486 1531 487
rect 1527 481 1531 482
rect 1543 486 1547 487
rect 1543 481 1547 482
rect 1639 486 1643 487
rect 1639 481 1643 482
rect 1727 486 1731 487
rect 1727 481 1731 482
rect 1823 486 1827 487
rect 1823 481 1827 482
rect 112 466 114 481
rect 160 476 162 481
rect 312 476 314 481
rect 464 476 466 481
rect 616 476 618 481
rect 760 476 762 481
rect 888 476 890 481
rect 1008 476 1010 481
rect 1128 476 1130 481
rect 1240 476 1242 481
rect 1344 476 1346 481
rect 1440 476 1442 481
rect 1544 476 1546 481
rect 1640 476 1642 481
rect 1728 476 1730 481
rect 158 475 164 476
rect 158 471 159 475
rect 163 471 164 475
rect 158 470 164 471
rect 310 475 316 476
rect 310 471 311 475
rect 315 471 316 475
rect 310 470 316 471
rect 462 475 468 476
rect 462 471 463 475
rect 467 471 468 475
rect 462 470 468 471
rect 614 475 620 476
rect 614 471 615 475
rect 619 471 620 475
rect 614 470 620 471
rect 758 475 764 476
rect 758 471 759 475
rect 763 471 764 475
rect 758 470 764 471
rect 886 475 892 476
rect 886 471 887 475
rect 891 471 892 475
rect 886 470 892 471
rect 1006 475 1012 476
rect 1006 471 1007 475
rect 1011 471 1012 475
rect 1006 470 1012 471
rect 1126 475 1132 476
rect 1126 471 1127 475
rect 1131 471 1132 475
rect 1126 470 1132 471
rect 1238 475 1244 476
rect 1238 471 1239 475
rect 1243 471 1244 475
rect 1238 470 1244 471
rect 1342 475 1348 476
rect 1342 471 1343 475
rect 1347 471 1348 475
rect 1342 470 1348 471
rect 1438 475 1444 476
rect 1438 471 1439 475
rect 1443 471 1444 475
rect 1438 470 1444 471
rect 1542 475 1548 476
rect 1542 471 1543 475
rect 1547 471 1548 475
rect 1542 470 1548 471
rect 1638 475 1644 476
rect 1638 471 1639 475
rect 1643 471 1644 475
rect 1638 470 1644 471
rect 1726 475 1732 476
rect 1726 471 1727 475
rect 1731 471 1732 475
rect 1726 470 1732 471
rect 1824 466 1826 481
rect 110 465 116 466
rect 110 461 111 465
rect 115 461 116 465
rect 110 460 116 461
rect 1822 465 1828 466
rect 1822 461 1823 465
rect 1827 461 1828 465
rect 1822 460 1828 461
rect 1864 455 1866 487
rect 2198 479 2204 480
rect 2198 475 2199 479
rect 2203 475 2204 479
rect 2198 474 2204 475
rect 2286 479 2292 480
rect 2286 475 2287 479
rect 2291 475 2292 479
rect 2286 474 2292 475
rect 2382 479 2388 480
rect 2382 475 2383 479
rect 2387 475 2388 479
rect 2382 474 2388 475
rect 2494 479 2500 480
rect 2494 475 2495 479
rect 2499 475 2500 479
rect 2494 474 2500 475
rect 2638 479 2644 480
rect 2638 475 2639 479
rect 2643 475 2644 479
rect 2638 474 2644 475
rect 2814 479 2820 480
rect 2814 475 2815 479
rect 2819 475 2820 479
rect 2814 474 2820 475
rect 3014 479 3020 480
rect 3014 475 3015 479
rect 3019 475 3020 479
rect 3014 474 3020 475
rect 3222 479 3228 480
rect 3222 475 3223 479
rect 3227 475 3228 479
rect 3222 474 3228 475
rect 3438 479 3444 480
rect 3438 475 3439 479
rect 3443 475 3444 479
rect 3438 474 3444 475
rect 2200 455 2202 474
rect 2288 455 2290 474
rect 2384 455 2386 474
rect 2496 455 2498 474
rect 2640 455 2642 474
rect 2816 455 2818 474
rect 3016 455 3018 474
rect 3224 455 3226 474
rect 3440 455 3442 474
rect 3576 455 3578 487
rect 1863 454 1867 455
rect 1863 449 1867 450
rect 1895 454 1899 455
rect 1895 449 1899 450
rect 2039 454 2043 455
rect 2039 449 2043 450
rect 2199 454 2203 455
rect 2199 449 2203 450
rect 2207 454 2211 455
rect 2207 449 2211 450
rect 2287 454 2291 455
rect 2287 449 2291 450
rect 2383 454 2387 455
rect 2383 449 2387 450
rect 2495 454 2499 455
rect 2495 449 2499 450
rect 2575 454 2579 455
rect 2575 449 2579 450
rect 2639 454 2643 455
rect 2639 449 2643 450
rect 2783 454 2787 455
rect 2783 449 2787 450
rect 2815 454 2819 455
rect 2815 449 2819 450
rect 3007 454 3011 455
rect 3007 449 3011 450
rect 3015 454 3019 455
rect 3015 449 3019 450
rect 3223 454 3227 455
rect 3223 449 3227 450
rect 3239 454 3243 455
rect 3239 449 3243 450
rect 3439 454 3443 455
rect 3439 449 3443 450
rect 3471 454 3475 455
rect 3471 449 3475 450
rect 3575 454 3579 455
rect 3575 449 3579 450
rect 110 448 116 449
rect 110 444 111 448
rect 115 444 116 448
rect 110 443 116 444
rect 1822 448 1828 449
rect 1822 444 1823 448
rect 1827 444 1828 448
rect 1822 443 1828 444
rect 112 419 114 443
rect 166 435 172 436
rect 166 431 167 435
rect 171 431 172 435
rect 166 430 172 431
rect 318 435 324 436
rect 318 431 319 435
rect 323 431 324 435
rect 318 430 324 431
rect 470 435 476 436
rect 470 431 471 435
rect 475 431 476 435
rect 470 430 476 431
rect 622 435 628 436
rect 622 431 623 435
rect 627 431 628 435
rect 622 430 628 431
rect 766 435 772 436
rect 766 431 767 435
rect 771 431 772 435
rect 766 430 772 431
rect 894 435 900 436
rect 894 431 895 435
rect 899 431 900 435
rect 894 430 900 431
rect 1014 435 1020 436
rect 1014 431 1015 435
rect 1019 431 1020 435
rect 1014 430 1020 431
rect 1134 435 1140 436
rect 1134 431 1135 435
rect 1139 431 1140 435
rect 1134 430 1140 431
rect 1246 435 1252 436
rect 1246 431 1247 435
rect 1251 431 1252 435
rect 1246 430 1252 431
rect 1350 435 1356 436
rect 1350 431 1351 435
rect 1355 431 1356 435
rect 1350 430 1356 431
rect 1446 435 1452 436
rect 1446 431 1447 435
rect 1451 431 1452 435
rect 1446 430 1452 431
rect 1550 435 1556 436
rect 1550 431 1551 435
rect 1555 431 1556 435
rect 1550 430 1556 431
rect 1646 435 1652 436
rect 1646 431 1647 435
rect 1651 431 1652 435
rect 1646 430 1652 431
rect 1734 435 1740 436
rect 1734 431 1735 435
rect 1739 431 1740 435
rect 1734 430 1740 431
rect 168 419 170 430
rect 320 419 322 430
rect 472 419 474 430
rect 624 419 626 430
rect 768 419 770 430
rect 896 419 898 430
rect 1016 419 1018 430
rect 1136 419 1138 430
rect 1248 419 1250 430
rect 1352 419 1354 430
rect 1448 419 1450 430
rect 1552 419 1554 430
rect 1648 419 1650 430
rect 1736 419 1738 430
rect 1824 419 1826 443
rect 1864 425 1866 449
rect 1896 438 1898 449
rect 2040 438 2042 449
rect 2208 438 2210 449
rect 2384 438 2386 449
rect 2576 438 2578 449
rect 2784 438 2786 449
rect 3008 438 3010 449
rect 3240 438 3242 449
rect 3472 438 3474 449
rect 1894 437 1900 438
rect 1894 433 1895 437
rect 1899 433 1900 437
rect 1894 432 1900 433
rect 2038 437 2044 438
rect 2038 433 2039 437
rect 2043 433 2044 437
rect 2038 432 2044 433
rect 2206 437 2212 438
rect 2206 433 2207 437
rect 2211 433 2212 437
rect 2206 432 2212 433
rect 2382 437 2388 438
rect 2382 433 2383 437
rect 2387 433 2388 437
rect 2382 432 2388 433
rect 2574 437 2580 438
rect 2574 433 2575 437
rect 2579 433 2580 437
rect 2574 432 2580 433
rect 2782 437 2788 438
rect 2782 433 2783 437
rect 2787 433 2788 437
rect 2782 432 2788 433
rect 3006 437 3012 438
rect 3006 433 3007 437
rect 3011 433 3012 437
rect 3006 432 3012 433
rect 3238 437 3244 438
rect 3238 433 3239 437
rect 3243 433 3244 437
rect 3238 432 3244 433
rect 3470 437 3476 438
rect 3470 433 3471 437
rect 3475 433 3476 437
rect 3470 432 3476 433
rect 3576 425 3578 449
rect 1862 424 1868 425
rect 1862 420 1863 424
rect 1867 420 1868 424
rect 1862 419 1868 420
rect 3574 424 3580 425
rect 3574 420 3575 424
rect 3579 420 3580 424
rect 3574 419 3580 420
rect 111 418 115 419
rect 111 413 115 414
rect 151 418 155 419
rect 151 413 155 414
rect 167 418 171 419
rect 167 413 171 414
rect 271 418 275 419
rect 271 413 275 414
rect 319 418 323 419
rect 319 413 323 414
rect 407 418 411 419
rect 407 413 411 414
rect 471 418 475 419
rect 471 413 475 414
rect 551 418 555 419
rect 551 413 555 414
rect 623 418 627 419
rect 623 413 627 414
rect 711 418 715 419
rect 711 413 715 414
rect 767 418 771 419
rect 767 413 771 414
rect 887 418 891 419
rect 887 413 891 414
rect 895 418 899 419
rect 895 413 899 414
rect 1015 418 1019 419
rect 1015 413 1019 414
rect 1063 418 1067 419
rect 1063 413 1067 414
rect 1135 418 1139 419
rect 1135 413 1139 414
rect 1247 418 1251 419
rect 1247 413 1251 414
rect 1351 418 1355 419
rect 1351 413 1355 414
rect 1439 418 1443 419
rect 1439 413 1443 414
rect 1447 418 1451 419
rect 1447 413 1451 414
rect 1551 418 1555 419
rect 1551 413 1555 414
rect 1639 418 1643 419
rect 1639 413 1643 414
rect 1647 418 1651 419
rect 1647 413 1651 414
rect 1735 418 1739 419
rect 1735 413 1739 414
rect 1823 418 1827 419
rect 1823 413 1827 414
rect 112 389 114 413
rect 152 402 154 413
rect 272 402 274 413
rect 408 402 410 413
rect 552 402 554 413
rect 712 402 714 413
rect 888 402 890 413
rect 1064 402 1066 413
rect 1248 402 1250 413
rect 1440 402 1442 413
rect 1640 402 1642 413
rect 150 401 156 402
rect 150 397 151 401
rect 155 397 156 401
rect 150 396 156 397
rect 270 401 276 402
rect 270 397 271 401
rect 275 397 276 401
rect 270 396 276 397
rect 406 401 412 402
rect 406 397 407 401
rect 411 397 412 401
rect 406 396 412 397
rect 550 401 556 402
rect 550 397 551 401
rect 555 397 556 401
rect 550 396 556 397
rect 710 401 716 402
rect 710 397 711 401
rect 715 397 716 401
rect 710 396 716 397
rect 886 401 892 402
rect 886 397 887 401
rect 891 397 892 401
rect 886 396 892 397
rect 1062 401 1068 402
rect 1062 397 1063 401
rect 1067 397 1068 401
rect 1062 396 1068 397
rect 1246 401 1252 402
rect 1246 397 1247 401
rect 1251 397 1252 401
rect 1246 396 1252 397
rect 1438 401 1444 402
rect 1438 397 1439 401
rect 1443 397 1444 401
rect 1438 396 1444 397
rect 1638 401 1644 402
rect 1638 397 1639 401
rect 1643 397 1644 401
rect 1638 396 1644 397
rect 1824 389 1826 413
rect 1862 407 1868 408
rect 1862 403 1863 407
rect 1867 403 1868 407
rect 1862 402 1868 403
rect 3574 407 3580 408
rect 3574 403 3575 407
rect 3579 403 3580 407
rect 3574 402 3580 403
rect 110 388 116 389
rect 110 384 111 388
rect 115 384 116 388
rect 110 383 116 384
rect 1822 388 1828 389
rect 1822 384 1823 388
rect 1827 384 1828 388
rect 1864 387 1866 402
rect 1886 397 1892 398
rect 1886 393 1887 397
rect 1891 393 1892 397
rect 1886 392 1892 393
rect 2030 397 2036 398
rect 2030 393 2031 397
rect 2035 393 2036 397
rect 2030 392 2036 393
rect 2198 397 2204 398
rect 2198 393 2199 397
rect 2203 393 2204 397
rect 2198 392 2204 393
rect 2374 397 2380 398
rect 2374 393 2375 397
rect 2379 393 2380 397
rect 2374 392 2380 393
rect 2566 397 2572 398
rect 2566 393 2567 397
rect 2571 393 2572 397
rect 2566 392 2572 393
rect 2774 397 2780 398
rect 2774 393 2775 397
rect 2779 393 2780 397
rect 2774 392 2780 393
rect 2998 397 3004 398
rect 2998 393 2999 397
rect 3003 393 3004 397
rect 2998 392 3004 393
rect 3230 397 3236 398
rect 3230 393 3231 397
rect 3235 393 3236 397
rect 3230 392 3236 393
rect 3462 397 3468 398
rect 3462 393 3463 397
rect 3467 393 3468 397
rect 3462 392 3468 393
rect 1888 387 1890 392
rect 2032 387 2034 392
rect 2200 387 2202 392
rect 2376 387 2378 392
rect 2568 387 2570 392
rect 2776 387 2778 392
rect 3000 387 3002 392
rect 3232 387 3234 392
rect 3464 387 3466 392
rect 3576 387 3578 402
rect 1822 383 1828 384
rect 1863 386 1867 387
rect 1863 381 1867 382
rect 1887 386 1891 387
rect 1887 381 1891 382
rect 1975 386 1979 387
rect 1975 381 1979 382
rect 2031 386 2035 387
rect 2031 381 2035 382
rect 2063 386 2067 387
rect 2063 381 2067 382
rect 2151 386 2155 387
rect 2151 381 2155 382
rect 2199 386 2203 387
rect 2199 381 2203 382
rect 2263 386 2267 387
rect 2263 381 2267 382
rect 2375 386 2379 387
rect 2375 381 2379 382
rect 2383 386 2387 387
rect 2383 381 2387 382
rect 2519 386 2523 387
rect 2519 381 2523 382
rect 2567 386 2571 387
rect 2567 381 2571 382
rect 2671 386 2675 387
rect 2671 381 2675 382
rect 2775 386 2779 387
rect 2775 381 2779 382
rect 2847 386 2851 387
rect 2847 381 2851 382
rect 2999 386 3003 387
rect 2999 381 3003 382
rect 3031 386 3035 387
rect 3031 381 3035 382
rect 3231 386 3235 387
rect 3231 381 3235 382
rect 3431 386 3435 387
rect 3431 381 3435 382
rect 3463 386 3467 387
rect 3463 381 3467 382
rect 3575 386 3579 387
rect 3575 381 3579 382
rect 110 371 116 372
rect 110 367 111 371
rect 115 367 116 371
rect 110 366 116 367
rect 1822 371 1828 372
rect 1822 367 1823 371
rect 1827 367 1828 371
rect 1822 366 1828 367
rect 1864 366 1866 381
rect 1888 376 1890 381
rect 1976 376 1978 381
rect 2064 376 2066 381
rect 2152 376 2154 381
rect 2264 376 2266 381
rect 2384 376 2386 381
rect 2520 376 2522 381
rect 2672 376 2674 381
rect 2848 376 2850 381
rect 3032 376 3034 381
rect 3232 376 3234 381
rect 3432 376 3434 381
rect 1886 375 1892 376
rect 1886 371 1887 375
rect 1891 371 1892 375
rect 1886 370 1892 371
rect 1974 375 1980 376
rect 1974 371 1975 375
rect 1979 371 1980 375
rect 1974 370 1980 371
rect 2062 375 2068 376
rect 2062 371 2063 375
rect 2067 371 2068 375
rect 2062 370 2068 371
rect 2150 375 2156 376
rect 2150 371 2151 375
rect 2155 371 2156 375
rect 2150 370 2156 371
rect 2262 375 2268 376
rect 2262 371 2263 375
rect 2267 371 2268 375
rect 2262 370 2268 371
rect 2382 375 2388 376
rect 2382 371 2383 375
rect 2387 371 2388 375
rect 2382 370 2388 371
rect 2518 375 2524 376
rect 2518 371 2519 375
rect 2523 371 2524 375
rect 2518 370 2524 371
rect 2670 375 2676 376
rect 2670 371 2671 375
rect 2675 371 2676 375
rect 2670 370 2676 371
rect 2846 375 2852 376
rect 2846 371 2847 375
rect 2851 371 2852 375
rect 2846 370 2852 371
rect 3030 375 3036 376
rect 3030 371 3031 375
rect 3035 371 3036 375
rect 3030 370 3036 371
rect 3230 375 3236 376
rect 3230 371 3231 375
rect 3235 371 3236 375
rect 3230 370 3236 371
rect 3430 375 3436 376
rect 3430 371 3431 375
rect 3435 371 3436 375
rect 3430 370 3436 371
rect 3576 366 3578 381
rect 112 335 114 366
rect 142 361 148 362
rect 142 357 143 361
rect 147 357 148 361
rect 142 356 148 357
rect 262 361 268 362
rect 262 357 263 361
rect 267 357 268 361
rect 262 356 268 357
rect 398 361 404 362
rect 398 357 399 361
rect 403 357 404 361
rect 398 356 404 357
rect 542 361 548 362
rect 542 357 543 361
rect 547 357 548 361
rect 542 356 548 357
rect 702 361 708 362
rect 702 357 703 361
rect 707 357 708 361
rect 702 356 708 357
rect 878 361 884 362
rect 878 357 879 361
rect 883 357 884 361
rect 878 356 884 357
rect 1054 361 1060 362
rect 1054 357 1055 361
rect 1059 357 1060 361
rect 1054 356 1060 357
rect 1238 361 1244 362
rect 1238 357 1239 361
rect 1243 357 1244 361
rect 1238 356 1244 357
rect 1430 361 1436 362
rect 1430 357 1431 361
rect 1435 357 1436 361
rect 1430 356 1436 357
rect 1630 361 1636 362
rect 1630 357 1631 361
rect 1635 357 1636 361
rect 1630 356 1636 357
rect 144 335 146 356
rect 264 335 266 356
rect 400 335 402 356
rect 544 335 546 356
rect 704 335 706 356
rect 880 335 882 356
rect 1056 335 1058 356
rect 1240 335 1242 356
rect 1432 335 1434 356
rect 1632 335 1634 356
rect 1824 335 1826 366
rect 1862 365 1868 366
rect 1862 361 1863 365
rect 1867 361 1868 365
rect 1862 360 1868 361
rect 3574 365 3580 366
rect 3574 361 3575 365
rect 3579 361 3580 365
rect 3574 360 3580 361
rect 1862 348 1868 349
rect 1862 344 1863 348
rect 1867 344 1868 348
rect 1862 343 1868 344
rect 3574 348 3580 349
rect 3574 344 3575 348
rect 3579 344 3580 348
rect 3574 343 3580 344
rect 111 334 115 335
rect 111 329 115 330
rect 135 334 139 335
rect 135 329 139 330
rect 143 334 147 335
rect 143 329 147 330
rect 223 334 227 335
rect 223 329 227 330
rect 263 334 267 335
rect 263 329 267 330
rect 311 334 315 335
rect 311 329 315 330
rect 399 334 403 335
rect 399 329 403 330
rect 487 334 491 335
rect 487 329 491 330
rect 543 334 547 335
rect 543 329 547 330
rect 575 334 579 335
rect 575 329 579 330
rect 663 334 667 335
rect 663 329 667 330
rect 703 334 707 335
rect 703 329 707 330
rect 751 334 755 335
rect 751 329 755 330
rect 839 334 843 335
rect 839 329 843 330
rect 879 334 883 335
rect 879 329 883 330
rect 927 334 931 335
rect 927 329 931 330
rect 1015 334 1019 335
rect 1015 329 1019 330
rect 1055 334 1059 335
rect 1055 329 1059 330
rect 1103 334 1107 335
rect 1103 329 1107 330
rect 1191 334 1195 335
rect 1191 329 1195 330
rect 1239 334 1243 335
rect 1239 329 1243 330
rect 1287 334 1291 335
rect 1287 329 1291 330
rect 1383 334 1387 335
rect 1383 329 1387 330
rect 1431 334 1435 335
rect 1431 329 1435 330
rect 1479 334 1483 335
rect 1479 329 1483 330
rect 1575 334 1579 335
rect 1575 329 1579 330
rect 1631 334 1635 335
rect 1631 329 1635 330
rect 1671 334 1675 335
rect 1671 329 1675 330
rect 1823 334 1827 335
rect 1823 329 1827 330
rect 112 314 114 329
rect 136 324 138 329
rect 224 324 226 329
rect 312 324 314 329
rect 400 324 402 329
rect 488 324 490 329
rect 576 324 578 329
rect 664 324 666 329
rect 752 324 754 329
rect 840 324 842 329
rect 928 324 930 329
rect 1016 324 1018 329
rect 1104 324 1106 329
rect 1192 324 1194 329
rect 1288 324 1290 329
rect 1384 324 1386 329
rect 1480 324 1482 329
rect 1576 324 1578 329
rect 1672 324 1674 329
rect 134 323 140 324
rect 134 319 135 323
rect 139 319 140 323
rect 134 318 140 319
rect 222 323 228 324
rect 222 319 223 323
rect 227 319 228 323
rect 222 318 228 319
rect 310 323 316 324
rect 310 319 311 323
rect 315 319 316 323
rect 310 318 316 319
rect 398 323 404 324
rect 398 319 399 323
rect 403 319 404 323
rect 398 318 404 319
rect 486 323 492 324
rect 486 319 487 323
rect 491 319 492 323
rect 486 318 492 319
rect 574 323 580 324
rect 574 319 575 323
rect 579 319 580 323
rect 574 318 580 319
rect 662 323 668 324
rect 662 319 663 323
rect 667 319 668 323
rect 662 318 668 319
rect 750 323 756 324
rect 750 319 751 323
rect 755 319 756 323
rect 750 318 756 319
rect 838 323 844 324
rect 838 319 839 323
rect 843 319 844 323
rect 838 318 844 319
rect 926 323 932 324
rect 926 319 927 323
rect 931 319 932 323
rect 926 318 932 319
rect 1014 323 1020 324
rect 1014 319 1015 323
rect 1019 319 1020 323
rect 1014 318 1020 319
rect 1102 323 1108 324
rect 1102 319 1103 323
rect 1107 319 1108 323
rect 1102 318 1108 319
rect 1190 323 1196 324
rect 1190 319 1191 323
rect 1195 319 1196 323
rect 1190 318 1196 319
rect 1286 323 1292 324
rect 1286 319 1287 323
rect 1291 319 1292 323
rect 1286 318 1292 319
rect 1382 323 1388 324
rect 1382 319 1383 323
rect 1387 319 1388 323
rect 1382 318 1388 319
rect 1478 323 1484 324
rect 1478 319 1479 323
rect 1483 319 1484 323
rect 1478 318 1484 319
rect 1574 323 1580 324
rect 1574 319 1575 323
rect 1579 319 1580 323
rect 1574 318 1580 319
rect 1670 323 1676 324
rect 1670 319 1671 323
rect 1675 319 1676 323
rect 1670 318 1676 319
rect 1824 314 1826 329
rect 1864 319 1866 343
rect 1894 335 1900 336
rect 1894 331 1895 335
rect 1899 331 1900 335
rect 1894 330 1900 331
rect 1982 335 1988 336
rect 1982 331 1983 335
rect 1987 331 1988 335
rect 1982 330 1988 331
rect 2070 335 2076 336
rect 2070 331 2071 335
rect 2075 331 2076 335
rect 2070 330 2076 331
rect 2158 335 2164 336
rect 2158 331 2159 335
rect 2163 331 2164 335
rect 2158 330 2164 331
rect 2270 335 2276 336
rect 2270 331 2271 335
rect 2275 331 2276 335
rect 2270 330 2276 331
rect 2390 335 2396 336
rect 2390 331 2391 335
rect 2395 331 2396 335
rect 2390 330 2396 331
rect 2526 335 2532 336
rect 2526 331 2527 335
rect 2531 331 2532 335
rect 2526 330 2532 331
rect 2678 335 2684 336
rect 2678 331 2679 335
rect 2683 331 2684 335
rect 2678 330 2684 331
rect 2854 335 2860 336
rect 2854 331 2855 335
rect 2859 331 2860 335
rect 2854 330 2860 331
rect 3038 335 3044 336
rect 3038 331 3039 335
rect 3043 331 3044 335
rect 3038 330 3044 331
rect 3238 335 3244 336
rect 3238 331 3239 335
rect 3243 331 3244 335
rect 3238 330 3244 331
rect 3438 335 3444 336
rect 3438 331 3439 335
rect 3443 331 3444 335
rect 3438 330 3444 331
rect 1896 319 1898 330
rect 1984 319 1986 330
rect 2072 319 2074 330
rect 2160 319 2162 330
rect 2272 319 2274 330
rect 2392 319 2394 330
rect 2528 319 2530 330
rect 2680 319 2682 330
rect 2856 319 2858 330
rect 3040 319 3042 330
rect 3240 319 3242 330
rect 3440 319 3442 330
rect 3576 319 3578 343
rect 1863 318 1867 319
rect 110 313 116 314
rect 110 309 111 313
rect 115 309 116 313
rect 110 308 116 309
rect 1822 313 1828 314
rect 1863 313 1867 314
rect 1895 318 1899 319
rect 1895 313 1899 314
rect 1983 318 1987 319
rect 1983 313 1987 314
rect 2071 318 2075 319
rect 2071 313 2075 314
rect 2159 318 2163 319
rect 2159 313 2163 314
rect 2247 318 2251 319
rect 2247 313 2251 314
rect 2271 318 2275 319
rect 2271 313 2275 314
rect 2359 318 2363 319
rect 2359 313 2363 314
rect 2391 318 2395 319
rect 2391 313 2395 314
rect 2471 318 2475 319
rect 2471 313 2475 314
rect 2527 318 2531 319
rect 2527 313 2531 314
rect 2583 318 2587 319
rect 2583 313 2587 314
rect 2679 318 2683 319
rect 2679 313 2683 314
rect 2695 318 2699 319
rect 2695 313 2699 314
rect 2807 318 2811 319
rect 2807 313 2811 314
rect 2855 318 2859 319
rect 2855 313 2859 314
rect 2919 318 2923 319
rect 2919 313 2923 314
rect 3039 318 3043 319
rect 3039 313 3043 314
rect 3159 318 3163 319
rect 3159 313 3163 314
rect 3239 318 3243 319
rect 3239 313 3243 314
rect 3439 318 3443 319
rect 3439 313 3443 314
rect 3575 318 3579 319
rect 3575 313 3579 314
rect 1822 309 1823 313
rect 1827 309 1828 313
rect 1822 308 1828 309
rect 110 296 116 297
rect 110 292 111 296
rect 115 292 116 296
rect 110 291 116 292
rect 1822 296 1828 297
rect 1822 292 1823 296
rect 1827 292 1828 296
rect 1822 291 1828 292
rect 112 263 114 291
rect 142 283 148 284
rect 142 279 143 283
rect 147 279 148 283
rect 142 278 148 279
rect 230 283 236 284
rect 230 279 231 283
rect 235 279 236 283
rect 230 278 236 279
rect 318 283 324 284
rect 318 279 319 283
rect 323 279 324 283
rect 318 278 324 279
rect 406 283 412 284
rect 406 279 407 283
rect 411 279 412 283
rect 406 278 412 279
rect 494 283 500 284
rect 494 279 495 283
rect 499 279 500 283
rect 494 278 500 279
rect 582 283 588 284
rect 582 279 583 283
rect 587 279 588 283
rect 582 278 588 279
rect 670 283 676 284
rect 670 279 671 283
rect 675 279 676 283
rect 670 278 676 279
rect 758 283 764 284
rect 758 279 759 283
rect 763 279 764 283
rect 758 278 764 279
rect 846 283 852 284
rect 846 279 847 283
rect 851 279 852 283
rect 846 278 852 279
rect 934 283 940 284
rect 934 279 935 283
rect 939 279 940 283
rect 934 278 940 279
rect 1022 283 1028 284
rect 1022 279 1023 283
rect 1027 279 1028 283
rect 1022 278 1028 279
rect 1110 283 1116 284
rect 1110 279 1111 283
rect 1115 279 1116 283
rect 1110 278 1116 279
rect 1198 283 1204 284
rect 1198 279 1199 283
rect 1203 279 1204 283
rect 1198 278 1204 279
rect 1294 283 1300 284
rect 1294 279 1295 283
rect 1299 279 1300 283
rect 1294 278 1300 279
rect 1390 283 1396 284
rect 1390 279 1391 283
rect 1395 279 1396 283
rect 1390 278 1396 279
rect 1486 283 1492 284
rect 1486 279 1487 283
rect 1491 279 1492 283
rect 1486 278 1492 279
rect 1582 283 1588 284
rect 1582 279 1583 283
rect 1587 279 1588 283
rect 1582 278 1588 279
rect 1678 283 1684 284
rect 1678 279 1679 283
rect 1683 279 1684 283
rect 1678 278 1684 279
rect 144 263 146 278
rect 232 263 234 278
rect 320 263 322 278
rect 408 263 410 278
rect 496 263 498 278
rect 584 263 586 278
rect 672 263 674 278
rect 760 263 762 278
rect 848 263 850 278
rect 936 263 938 278
rect 1024 263 1026 278
rect 1112 263 1114 278
rect 1200 263 1202 278
rect 1296 263 1298 278
rect 1392 263 1394 278
rect 1488 263 1490 278
rect 1584 263 1586 278
rect 1680 263 1682 278
rect 1824 263 1826 291
rect 1864 289 1866 313
rect 1896 302 1898 313
rect 1984 302 1986 313
rect 2072 302 2074 313
rect 2160 302 2162 313
rect 2248 302 2250 313
rect 2360 302 2362 313
rect 2472 302 2474 313
rect 2584 302 2586 313
rect 2696 302 2698 313
rect 2808 302 2810 313
rect 2920 302 2922 313
rect 3040 302 3042 313
rect 3160 302 3162 313
rect 1894 301 1900 302
rect 1894 297 1895 301
rect 1899 297 1900 301
rect 1894 296 1900 297
rect 1982 301 1988 302
rect 1982 297 1983 301
rect 1987 297 1988 301
rect 1982 296 1988 297
rect 2070 301 2076 302
rect 2070 297 2071 301
rect 2075 297 2076 301
rect 2070 296 2076 297
rect 2158 301 2164 302
rect 2158 297 2159 301
rect 2163 297 2164 301
rect 2158 296 2164 297
rect 2246 301 2252 302
rect 2246 297 2247 301
rect 2251 297 2252 301
rect 2246 296 2252 297
rect 2358 301 2364 302
rect 2358 297 2359 301
rect 2363 297 2364 301
rect 2358 296 2364 297
rect 2470 301 2476 302
rect 2470 297 2471 301
rect 2475 297 2476 301
rect 2470 296 2476 297
rect 2582 301 2588 302
rect 2582 297 2583 301
rect 2587 297 2588 301
rect 2582 296 2588 297
rect 2694 301 2700 302
rect 2694 297 2695 301
rect 2699 297 2700 301
rect 2694 296 2700 297
rect 2806 301 2812 302
rect 2806 297 2807 301
rect 2811 297 2812 301
rect 2806 296 2812 297
rect 2918 301 2924 302
rect 2918 297 2919 301
rect 2923 297 2924 301
rect 2918 296 2924 297
rect 3038 301 3044 302
rect 3038 297 3039 301
rect 3043 297 3044 301
rect 3038 296 3044 297
rect 3158 301 3164 302
rect 3158 297 3159 301
rect 3163 297 3164 301
rect 3158 296 3164 297
rect 3576 289 3578 313
rect 1862 288 1868 289
rect 1862 284 1863 288
rect 1867 284 1868 288
rect 1862 283 1868 284
rect 3574 288 3580 289
rect 3574 284 3575 288
rect 3579 284 3580 288
rect 3574 283 3580 284
rect 1862 271 1868 272
rect 1862 267 1863 271
rect 1867 267 1868 271
rect 1862 266 1868 267
rect 3574 271 3580 272
rect 3574 267 3575 271
rect 3579 267 3580 271
rect 3574 266 3580 267
rect 111 262 115 263
rect 111 257 115 258
rect 143 262 147 263
rect 143 257 147 258
rect 231 262 235 263
rect 231 257 235 258
rect 319 262 323 263
rect 319 257 323 258
rect 407 262 411 263
rect 407 257 411 258
rect 495 262 499 263
rect 495 257 499 258
rect 583 262 587 263
rect 583 257 587 258
rect 671 262 675 263
rect 671 257 675 258
rect 759 262 763 263
rect 759 257 763 258
rect 847 262 851 263
rect 847 257 851 258
rect 935 262 939 263
rect 935 257 939 258
rect 1023 262 1027 263
rect 1023 257 1027 258
rect 1111 262 1115 263
rect 1111 257 1115 258
rect 1199 262 1203 263
rect 1199 257 1203 258
rect 1287 262 1291 263
rect 1287 257 1291 258
rect 1295 262 1299 263
rect 1295 257 1299 258
rect 1375 262 1379 263
rect 1375 257 1379 258
rect 1391 262 1395 263
rect 1391 257 1395 258
rect 1463 262 1467 263
rect 1463 257 1467 258
rect 1487 262 1491 263
rect 1487 257 1491 258
rect 1551 262 1555 263
rect 1551 257 1555 258
rect 1583 262 1587 263
rect 1583 257 1587 258
rect 1639 262 1643 263
rect 1639 257 1643 258
rect 1679 262 1683 263
rect 1679 257 1683 258
rect 1727 262 1731 263
rect 1727 257 1731 258
rect 1823 262 1827 263
rect 1823 257 1827 258
rect 112 233 114 257
rect 144 246 146 257
rect 232 246 234 257
rect 320 246 322 257
rect 408 246 410 257
rect 496 246 498 257
rect 584 246 586 257
rect 672 246 674 257
rect 760 246 762 257
rect 848 246 850 257
rect 936 246 938 257
rect 1024 246 1026 257
rect 1112 246 1114 257
rect 1200 246 1202 257
rect 1288 246 1290 257
rect 1376 246 1378 257
rect 1464 246 1466 257
rect 1552 246 1554 257
rect 1640 246 1642 257
rect 1728 246 1730 257
rect 142 245 148 246
rect 142 241 143 245
rect 147 241 148 245
rect 142 240 148 241
rect 230 245 236 246
rect 230 241 231 245
rect 235 241 236 245
rect 230 240 236 241
rect 318 245 324 246
rect 318 241 319 245
rect 323 241 324 245
rect 318 240 324 241
rect 406 245 412 246
rect 406 241 407 245
rect 411 241 412 245
rect 406 240 412 241
rect 494 245 500 246
rect 494 241 495 245
rect 499 241 500 245
rect 494 240 500 241
rect 582 245 588 246
rect 582 241 583 245
rect 587 241 588 245
rect 582 240 588 241
rect 670 245 676 246
rect 670 241 671 245
rect 675 241 676 245
rect 670 240 676 241
rect 758 245 764 246
rect 758 241 759 245
rect 763 241 764 245
rect 758 240 764 241
rect 846 245 852 246
rect 846 241 847 245
rect 851 241 852 245
rect 846 240 852 241
rect 934 245 940 246
rect 934 241 935 245
rect 939 241 940 245
rect 934 240 940 241
rect 1022 245 1028 246
rect 1022 241 1023 245
rect 1027 241 1028 245
rect 1022 240 1028 241
rect 1110 245 1116 246
rect 1110 241 1111 245
rect 1115 241 1116 245
rect 1110 240 1116 241
rect 1198 245 1204 246
rect 1198 241 1199 245
rect 1203 241 1204 245
rect 1198 240 1204 241
rect 1286 245 1292 246
rect 1286 241 1287 245
rect 1291 241 1292 245
rect 1286 240 1292 241
rect 1374 245 1380 246
rect 1374 241 1375 245
rect 1379 241 1380 245
rect 1374 240 1380 241
rect 1462 245 1468 246
rect 1462 241 1463 245
rect 1467 241 1468 245
rect 1462 240 1468 241
rect 1550 245 1556 246
rect 1550 241 1551 245
rect 1555 241 1556 245
rect 1550 240 1556 241
rect 1638 245 1644 246
rect 1638 241 1639 245
rect 1643 241 1644 245
rect 1638 240 1644 241
rect 1726 245 1732 246
rect 1726 241 1727 245
rect 1731 241 1732 245
rect 1726 240 1732 241
rect 1824 233 1826 257
rect 1864 251 1866 266
rect 1886 261 1892 262
rect 1886 257 1887 261
rect 1891 257 1892 261
rect 1886 256 1892 257
rect 1974 261 1980 262
rect 1974 257 1975 261
rect 1979 257 1980 261
rect 1974 256 1980 257
rect 2062 261 2068 262
rect 2062 257 2063 261
rect 2067 257 2068 261
rect 2062 256 2068 257
rect 2150 261 2156 262
rect 2150 257 2151 261
rect 2155 257 2156 261
rect 2150 256 2156 257
rect 2238 261 2244 262
rect 2238 257 2239 261
rect 2243 257 2244 261
rect 2238 256 2244 257
rect 2350 261 2356 262
rect 2350 257 2351 261
rect 2355 257 2356 261
rect 2350 256 2356 257
rect 2462 261 2468 262
rect 2462 257 2463 261
rect 2467 257 2468 261
rect 2462 256 2468 257
rect 2574 261 2580 262
rect 2574 257 2575 261
rect 2579 257 2580 261
rect 2574 256 2580 257
rect 2686 261 2692 262
rect 2686 257 2687 261
rect 2691 257 2692 261
rect 2686 256 2692 257
rect 2798 261 2804 262
rect 2798 257 2799 261
rect 2803 257 2804 261
rect 2798 256 2804 257
rect 2910 261 2916 262
rect 2910 257 2911 261
rect 2915 257 2916 261
rect 2910 256 2916 257
rect 3030 261 3036 262
rect 3030 257 3031 261
rect 3035 257 3036 261
rect 3030 256 3036 257
rect 3150 261 3156 262
rect 3150 257 3151 261
rect 3155 257 3156 261
rect 3150 256 3156 257
rect 1888 251 1890 256
rect 1976 251 1978 256
rect 2064 251 2066 256
rect 2152 251 2154 256
rect 2240 251 2242 256
rect 2352 251 2354 256
rect 2464 251 2466 256
rect 2576 251 2578 256
rect 2688 251 2690 256
rect 2800 251 2802 256
rect 2912 251 2914 256
rect 3032 251 3034 256
rect 3152 251 3154 256
rect 3576 251 3578 266
rect 1863 250 1867 251
rect 1863 245 1867 246
rect 1887 250 1891 251
rect 1887 245 1891 246
rect 1975 250 1979 251
rect 1975 245 1979 246
rect 2063 250 2067 251
rect 2063 245 2067 246
rect 2151 250 2155 251
rect 2151 245 2155 246
rect 2239 250 2243 251
rect 2239 245 2243 246
rect 2263 250 2267 251
rect 2263 245 2267 246
rect 2351 250 2355 251
rect 2351 245 2355 246
rect 2399 250 2403 251
rect 2399 245 2403 246
rect 2463 250 2467 251
rect 2463 245 2467 246
rect 2535 250 2539 251
rect 2535 245 2539 246
rect 2575 250 2579 251
rect 2575 245 2579 246
rect 2679 250 2683 251
rect 2679 245 2683 246
rect 2687 250 2691 251
rect 2687 245 2691 246
rect 2799 250 2803 251
rect 2799 245 2803 246
rect 2815 250 2819 251
rect 2815 245 2819 246
rect 2911 250 2915 251
rect 2911 245 2915 246
rect 2951 250 2955 251
rect 2951 245 2955 246
rect 3031 250 3035 251
rect 3031 245 3035 246
rect 3087 250 3091 251
rect 3087 245 3091 246
rect 3151 250 3155 251
rect 3151 245 3155 246
rect 3223 250 3227 251
rect 3223 245 3227 246
rect 3359 250 3363 251
rect 3359 245 3363 246
rect 3479 250 3483 251
rect 3479 245 3483 246
rect 3575 250 3579 251
rect 3575 245 3579 246
rect 110 232 116 233
rect 110 228 111 232
rect 115 228 116 232
rect 110 227 116 228
rect 1822 232 1828 233
rect 1822 228 1823 232
rect 1827 228 1828 232
rect 1864 230 1866 245
rect 1888 240 1890 245
rect 1976 240 1978 245
rect 2064 240 2066 245
rect 2152 240 2154 245
rect 2264 240 2266 245
rect 2400 240 2402 245
rect 2536 240 2538 245
rect 2680 240 2682 245
rect 2816 240 2818 245
rect 2952 240 2954 245
rect 3088 240 3090 245
rect 3224 240 3226 245
rect 3360 240 3362 245
rect 3480 240 3482 245
rect 1886 239 1892 240
rect 1886 235 1887 239
rect 1891 235 1892 239
rect 1886 234 1892 235
rect 1974 239 1980 240
rect 1974 235 1975 239
rect 1979 235 1980 239
rect 1974 234 1980 235
rect 2062 239 2068 240
rect 2062 235 2063 239
rect 2067 235 2068 239
rect 2062 234 2068 235
rect 2150 239 2156 240
rect 2150 235 2151 239
rect 2155 235 2156 239
rect 2150 234 2156 235
rect 2262 239 2268 240
rect 2262 235 2263 239
rect 2267 235 2268 239
rect 2262 234 2268 235
rect 2398 239 2404 240
rect 2398 235 2399 239
rect 2403 235 2404 239
rect 2398 234 2404 235
rect 2534 239 2540 240
rect 2534 235 2535 239
rect 2539 235 2540 239
rect 2534 234 2540 235
rect 2678 239 2684 240
rect 2678 235 2679 239
rect 2683 235 2684 239
rect 2678 234 2684 235
rect 2814 239 2820 240
rect 2814 235 2815 239
rect 2819 235 2820 239
rect 2814 234 2820 235
rect 2950 239 2956 240
rect 2950 235 2951 239
rect 2955 235 2956 239
rect 2950 234 2956 235
rect 3086 239 3092 240
rect 3086 235 3087 239
rect 3091 235 3092 239
rect 3086 234 3092 235
rect 3222 239 3228 240
rect 3222 235 3223 239
rect 3227 235 3228 239
rect 3222 234 3228 235
rect 3358 239 3364 240
rect 3358 235 3359 239
rect 3363 235 3364 239
rect 3358 234 3364 235
rect 3478 239 3484 240
rect 3478 235 3479 239
rect 3483 235 3484 239
rect 3478 234 3484 235
rect 3576 230 3578 245
rect 1822 227 1828 228
rect 1862 229 1868 230
rect 1862 225 1863 229
rect 1867 225 1868 229
rect 1862 224 1868 225
rect 3574 229 3580 230
rect 3574 225 3575 229
rect 3579 225 3580 229
rect 3574 224 3580 225
rect 110 215 116 216
rect 110 211 111 215
rect 115 211 116 215
rect 110 210 116 211
rect 1822 215 1828 216
rect 1822 211 1823 215
rect 1827 211 1828 215
rect 1822 210 1828 211
rect 1862 212 1868 213
rect 112 195 114 210
rect 134 205 140 206
rect 134 201 135 205
rect 139 201 140 205
rect 134 200 140 201
rect 222 205 228 206
rect 222 201 223 205
rect 227 201 228 205
rect 222 200 228 201
rect 310 205 316 206
rect 310 201 311 205
rect 315 201 316 205
rect 310 200 316 201
rect 398 205 404 206
rect 398 201 399 205
rect 403 201 404 205
rect 398 200 404 201
rect 486 205 492 206
rect 486 201 487 205
rect 491 201 492 205
rect 486 200 492 201
rect 574 205 580 206
rect 574 201 575 205
rect 579 201 580 205
rect 574 200 580 201
rect 662 205 668 206
rect 662 201 663 205
rect 667 201 668 205
rect 662 200 668 201
rect 750 205 756 206
rect 750 201 751 205
rect 755 201 756 205
rect 750 200 756 201
rect 838 205 844 206
rect 838 201 839 205
rect 843 201 844 205
rect 838 200 844 201
rect 926 205 932 206
rect 926 201 927 205
rect 931 201 932 205
rect 926 200 932 201
rect 1014 205 1020 206
rect 1014 201 1015 205
rect 1019 201 1020 205
rect 1014 200 1020 201
rect 1102 205 1108 206
rect 1102 201 1103 205
rect 1107 201 1108 205
rect 1102 200 1108 201
rect 1190 205 1196 206
rect 1190 201 1191 205
rect 1195 201 1196 205
rect 1190 200 1196 201
rect 1278 205 1284 206
rect 1278 201 1279 205
rect 1283 201 1284 205
rect 1278 200 1284 201
rect 1366 205 1372 206
rect 1366 201 1367 205
rect 1371 201 1372 205
rect 1366 200 1372 201
rect 1454 205 1460 206
rect 1454 201 1455 205
rect 1459 201 1460 205
rect 1454 200 1460 201
rect 1542 205 1548 206
rect 1542 201 1543 205
rect 1547 201 1548 205
rect 1542 200 1548 201
rect 1630 205 1636 206
rect 1630 201 1631 205
rect 1635 201 1636 205
rect 1630 200 1636 201
rect 1718 205 1724 206
rect 1718 201 1719 205
rect 1723 201 1724 205
rect 1718 200 1724 201
rect 136 195 138 200
rect 224 195 226 200
rect 312 195 314 200
rect 400 195 402 200
rect 488 195 490 200
rect 576 195 578 200
rect 664 195 666 200
rect 752 195 754 200
rect 840 195 842 200
rect 928 195 930 200
rect 1016 195 1018 200
rect 1104 195 1106 200
rect 1192 195 1194 200
rect 1280 195 1282 200
rect 1368 195 1370 200
rect 1456 195 1458 200
rect 1544 195 1546 200
rect 1632 195 1634 200
rect 1720 195 1722 200
rect 1824 195 1826 210
rect 1862 208 1863 212
rect 1867 208 1868 212
rect 1862 207 1868 208
rect 3574 212 3580 213
rect 3574 208 3575 212
rect 3579 208 3580 212
rect 3574 207 3580 208
rect 111 194 115 195
rect 111 189 115 190
rect 135 194 139 195
rect 135 189 139 190
rect 223 194 227 195
rect 223 189 227 190
rect 311 194 315 195
rect 311 189 315 190
rect 399 194 403 195
rect 399 189 403 190
rect 487 194 491 195
rect 487 189 491 190
rect 575 194 579 195
rect 575 189 579 190
rect 663 194 667 195
rect 663 189 667 190
rect 751 194 755 195
rect 751 189 755 190
rect 839 194 843 195
rect 839 189 843 190
rect 927 194 931 195
rect 927 189 931 190
rect 1015 194 1019 195
rect 1015 189 1019 190
rect 1103 194 1107 195
rect 1103 189 1107 190
rect 1191 194 1195 195
rect 1191 189 1195 190
rect 1279 194 1283 195
rect 1279 189 1283 190
rect 1367 194 1371 195
rect 1367 189 1371 190
rect 1455 194 1459 195
rect 1455 189 1459 190
rect 1543 194 1547 195
rect 1543 189 1547 190
rect 1631 194 1635 195
rect 1631 189 1635 190
rect 1719 194 1723 195
rect 1719 189 1723 190
rect 1823 194 1827 195
rect 1823 189 1827 190
rect 1864 151 1866 207
rect 1894 199 1900 200
rect 1894 195 1895 199
rect 1899 195 1900 199
rect 1894 194 1900 195
rect 1982 199 1988 200
rect 1982 195 1983 199
rect 1987 195 1988 199
rect 1982 194 1988 195
rect 2070 199 2076 200
rect 2070 195 2071 199
rect 2075 195 2076 199
rect 2070 194 2076 195
rect 2158 199 2164 200
rect 2158 195 2159 199
rect 2163 195 2164 199
rect 2158 194 2164 195
rect 2270 199 2276 200
rect 2270 195 2271 199
rect 2275 195 2276 199
rect 2270 194 2276 195
rect 2406 199 2412 200
rect 2406 195 2407 199
rect 2411 195 2412 199
rect 2406 194 2412 195
rect 2542 199 2548 200
rect 2542 195 2543 199
rect 2547 195 2548 199
rect 2542 194 2548 195
rect 2686 199 2692 200
rect 2686 195 2687 199
rect 2691 195 2692 199
rect 2686 194 2692 195
rect 2822 199 2828 200
rect 2822 195 2823 199
rect 2827 195 2828 199
rect 2822 194 2828 195
rect 2958 199 2964 200
rect 2958 195 2959 199
rect 2963 195 2964 199
rect 2958 194 2964 195
rect 3094 199 3100 200
rect 3094 195 3095 199
rect 3099 195 3100 199
rect 3094 194 3100 195
rect 3230 199 3236 200
rect 3230 195 3231 199
rect 3235 195 3236 199
rect 3230 194 3236 195
rect 3366 199 3372 200
rect 3366 195 3367 199
rect 3371 195 3372 199
rect 3366 194 3372 195
rect 3486 199 3492 200
rect 3486 195 3487 199
rect 3491 195 3492 199
rect 3486 194 3492 195
rect 1896 151 1898 194
rect 1984 151 1986 194
rect 2072 151 2074 194
rect 2160 151 2162 194
rect 2272 151 2274 194
rect 2408 151 2410 194
rect 2544 151 2546 194
rect 2688 151 2690 194
rect 2824 151 2826 194
rect 2960 151 2962 194
rect 3096 151 3098 194
rect 3232 151 3234 194
rect 3368 151 3370 194
rect 3488 151 3490 194
rect 3576 151 3578 207
rect 1863 150 1867 151
rect 1863 145 1867 146
rect 1895 150 1899 151
rect 1895 145 1899 146
rect 1983 150 1987 151
rect 1983 145 1987 146
rect 2071 150 2075 151
rect 2071 145 2075 146
rect 2159 150 2163 151
rect 2159 145 2163 146
rect 2271 150 2275 151
rect 2271 145 2275 146
rect 2407 150 2411 151
rect 2407 145 2411 146
rect 2543 150 2547 151
rect 2543 145 2547 146
rect 2687 150 2691 151
rect 2687 145 2691 146
rect 2783 150 2787 151
rect 2783 145 2787 146
rect 2823 150 2827 151
rect 2823 145 2827 146
rect 2871 150 2875 151
rect 2871 145 2875 146
rect 2959 150 2963 151
rect 2959 145 2963 146
rect 3047 150 3051 151
rect 3047 145 3051 146
rect 3095 150 3099 151
rect 3095 145 3099 146
rect 3135 150 3139 151
rect 3135 145 3139 146
rect 3223 150 3227 151
rect 3223 145 3227 146
rect 3231 150 3235 151
rect 3231 145 3235 146
rect 3311 150 3315 151
rect 3311 145 3315 146
rect 3367 150 3371 151
rect 3367 145 3371 146
rect 3399 150 3403 151
rect 3399 145 3403 146
rect 3487 150 3491 151
rect 3487 145 3491 146
rect 3575 150 3579 151
rect 3575 145 3579 146
rect 1864 121 1866 145
rect 2784 134 2786 145
rect 2872 134 2874 145
rect 2960 134 2962 145
rect 3048 134 3050 145
rect 3136 134 3138 145
rect 3224 134 3226 145
rect 3312 134 3314 145
rect 3400 134 3402 145
rect 3488 134 3490 145
rect 2782 133 2788 134
rect 2782 129 2783 133
rect 2787 129 2788 133
rect 2782 128 2788 129
rect 2870 133 2876 134
rect 2870 129 2871 133
rect 2875 129 2876 133
rect 2870 128 2876 129
rect 2958 133 2964 134
rect 2958 129 2959 133
rect 2963 129 2964 133
rect 2958 128 2964 129
rect 3046 133 3052 134
rect 3046 129 3047 133
rect 3051 129 3052 133
rect 3046 128 3052 129
rect 3134 133 3140 134
rect 3134 129 3135 133
rect 3139 129 3140 133
rect 3134 128 3140 129
rect 3222 133 3228 134
rect 3222 129 3223 133
rect 3227 129 3228 133
rect 3222 128 3228 129
rect 3310 133 3316 134
rect 3310 129 3311 133
rect 3315 129 3316 133
rect 3310 128 3316 129
rect 3398 133 3404 134
rect 3398 129 3399 133
rect 3403 129 3404 133
rect 3398 128 3404 129
rect 3486 133 3492 134
rect 3486 129 3487 133
rect 3491 129 3492 133
rect 3486 128 3492 129
rect 3576 121 3578 145
rect 1862 120 1868 121
rect 1862 116 1863 120
rect 1867 116 1868 120
rect 1862 115 1868 116
rect 3574 120 3580 121
rect 3574 116 3575 120
rect 3579 116 3580 120
rect 3574 115 3580 116
rect 1862 103 1868 104
rect 1862 99 1863 103
rect 1867 99 1868 103
rect 1862 98 1868 99
rect 3574 103 3580 104
rect 3574 99 3575 103
rect 3579 99 3580 103
rect 3574 98 3580 99
rect 1864 83 1866 98
rect 2774 93 2780 94
rect 2774 89 2775 93
rect 2779 89 2780 93
rect 2774 88 2780 89
rect 2862 93 2868 94
rect 2862 89 2863 93
rect 2867 89 2868 93
rect 2862 88 2868 89
rect 2950 93 2956 94
rect 2950 89 2951 93
rect 2955 89 2956 93
rect 2950 88 2956 89
rect 3038 93 3044 94
rect 3038 89 3039 93
rect 3043 89 3044 93
rect 3038 88 3044 89
rect 3126 93 3132 94
rect 3126 89 3127 93
rect 3131 89 3132 93
rect 3126 88 3132 89
rect 3214 93 3220 94
rect 3214 89 3215 93
rect 3219 89 3220 93
rect 3214 88 3220 89
rect 3302 93 3308 94
rect 3302 89 3303 93
rect 3307 89 3308 93
rect 3302 88 3308 89
rect 3390 93 3396 94
rect 3390 89 3391 93
rect 3395 89 3396 93
rect 3390 88 3396 89
rect 3478 93 3484 94
rect 3478 89 3479 93
rect 3483 89 3484 93
rect 3478 88 3484 89
rect 2776 83 2778 88
rect 2864 83 2866 88
rect 2952 83 2954 88
rect 3040 83 3042 88
rect 3128 83 3130 88
rect 3216 83 3218 88
rect 3304 83 3306 88
rect 3392 83 3394 88
rect 3480 83 3482 88
rect 3576 83 3578 98
rect 1863 82 1867 83
rect 1863 77 1867 78
rect 2775 82 2779 83
rect 2775 77 2779 78
rect 2863 82 2867 83
rect 2863 77 2867 78
rect 2951 82 2955 83
rect 2951 77 2955 78
rect 3039 82 3043 83
rect 3039 77 3043 78
rect 3127 82 3131 83
rect 3127 77 3131 78
rect 3215 82 3219 83
rect 3215 77 3219 78
rect 3303 82 3307 83
rect 3303 77 3307 78
rect 3391 82 3395 83
rect 3391 77 3395 78
rect 3479 82 3483 83
rect 3479 77 3483 78
rect 3575 82 3579 83
rect 3575 77 3579 78
<< m4c >>
rect 111 3666 115 3670
rect 135 3666 139 3670
rect 223 3666 227 3670
rect 1823 3666 1827 3670
rect 111 3598 115 3602
rect 143 3598 147 3602
rect 231 3598 235 3602
rect 319 3598 323 3602
rect 407 3598 411 3602
rect 495 3598 499 3602
rect 1823 3598 1827 3602
rect 1863 3590 1867 3594
rect 1887 3590 1891 3594
rect 1975 3590 1979 3594
rect 2063 3590 2067 3594
rect 2151 3590 2155 3594
rect 2239 3590 2243 3594
rect 2327 3590 2331 3594
rect 2431 3590 2435 3594
rect 2535 3590 2539 3594
rect 2631 3590 2635 3594
rect 2727 3590 2731 3594
rect 2823 3590 2827 3594
rect 2919 3590 2923 3594
rect 3015 3590 3019 3594
rect 3119 3590 3123 3594
rect 3223 3590 3227 3594
rect 3575 3590 3579 3594
rect 111 3530 115 3534
rect 135 3530 139 3534
rect 223 3530 227 3534
rect 247 3530 251 3534
rect 311 3530 315 3534
rect 375 3530 379 3534
rect 399 3530 403 3534
rect 487 3530 491 3534
rect 503 3530 507 3534
rect 623 3530 627 3534
rect 743 3530 747 3534
rect 863 3530 867 3534
rect 975 3530 979 3534
rect 1079 3530 1083 3534
rect 1175 3530 1179 3534
rect 1271 3530 1275 3534
rect 1367 3530 1371 3534
rect 1471 3530 1475 3534
rect 1575 3530 1579 3534
rect 1823 3530 1827 3534
rect 1863 3522 1867 3526
rect 1895 3522 1899 3526
rect 1983 3522 1987 3526
rect 2071 3522 2075 3526
rect 2103 3522 2107 3526
rect 2159 3522 2163 3526
rect 2231 3522 2235 3526
rect 2247 3522 2251 3526
rect 2335 3522 2339 3526
rect 2367 3522 2371 3526
rect 2439 3522 2443 3526
rect 2511 3522 2515 3526
rect 2543 3522 2547 3526
rect 2639 3522 2643 3526
rect 2655 3522 2659 3526
rect 2735 3522 2739 3526
rect 2791 3522 2795 3526
rect 2831 3522 2835 3526
rect 2927 3522 2931 3526
rect 2935 3522 2939 3526
rect 3023 3522 3027 3526
rect 3079 3522 3083 3526
rect 3127 3522 3131 3526
rect 3223 3522 3227 3526
rect 3231 3522 3235 3526
rect 3575 3522 3579 3526
rect 111 3462 115 3466
rect 175 3462 179 3466
rect 255 3462 259 3466
rect 303 3462 307 3466
rect 383 3462 387 3466
rect 447 3462 451 3466
rect 511 3462 515 3466
rect 591 3462 595 3466
rect 631 3462 635 3466
rect 743 3462 747 3466
rect 751 3462 755 3466
rect 871 3462 875 3466
rect 895 3462 899 3466
rect 983 3462 987 3466
rect 1039 3462 1043 3466
rect 1087 3462 1091 3466
rect 1183 3462 1187 3466
rect 1279 3462 1283 3466
rect 1327 3462 1331 3466
rect 1375 3462 1379 3466
rect 1479 3462 1483 3466
rect 1583 3462 1587 3466
rect 1823 3462 1827 3466
rect 1863 3446 1867 3450
rect 1887 3446 1891 3450
rect 1975 3446 1979 3450
rect 2023 3446 2027 3450
rect 2095 3446 2099 3450
rect 2191 3446 2195 3450
rect 2223 3446 2227 3450
rect 2359 3446 2363 3450
rect 2367 3446 2371 3450
rect 2503 3446 2507 3450
rect 2543 3446 2547 3450
rect 2647 3446 2651 3450
rect 2711 3446 2715 3450
rect 2783 3446 2787 3450
rect 2871 3446 2875 3450
rect 2927 3446 2931 3450
rect 3031 3446 3035 3450
rect 3071 3446 3075 3450
rect 3191 3446 3195 3450
rect 3215 3446 3219 3450
rect 3359 3446 3363 3450
rect 3575 3446 3579 3450
rect 111 3394 115 3398
rect 135 3394 139 3398
rect 167 3394 171 3398
rect 263 3394 267 3398
rect 295 3394 299 3398
rect 407 3394 411 3398
rect 439 3394 443 3398
rect 567 3394 571 3398
rect 583 3394 587 3398
rect 727 3394 731 3398
rect 735 3394 739 3398
rect 887 3394 891 3398
rect 1031 3394 1035 3398
rect 1047 3394 1051 3398
rect 1175 3394 1179 3398
rect 1207 3394 1211 3398
rect 1319 3394 1323 3398
rect 1367 3394 1371 3398
rect 1471 3394 1475 3398
rect 1527 3394 1531 3398
rect 1823 3394 1827 3398
rect 1863 3370 1867 3374
rect 1895 3370 1899 3374
rect 2031 3370 2035 3374
rect 2199 3370 2203 3374
rect 2375 3370 2379 3374
rect 2551 3370 2555 3374
rect 2719 3370 2723 3374
rect 2879 3370 2883 3374
rect 3039 3370 3043 3374
rect 3191 3370 3195 3374
rect 3199 3370 3203 3374
rect 3343 3370 3347 3374
rect 3367 3370 3371 3374
rect 3487 3370 3491 3374
rect 3575 3370 3579 3374
rect 111 3322 115 3326
rect 143 3322 147 3326
rect 207 3322 211 3326
rect 271 3322 275 3326
rect 335 3322 339 3326
rect 415 3322 419 3326
rect 479 3322 483 3326
rect 575 3322 579 3326
rect 639 3322 643 3326
rect 735 3322 739 3326
rect 807 3322 811 3326
rect 895 3322 899 3326
rect 983 3322 987 3326
rect 1055 3322 1059 3326
rect 1167 3322 1171 3326
rect 1215 3322 1219 3326
rect 1351 3322 1355 3326
rect 1375 3322 1379 3326
rect 1535 3322 1539 3326
rect 1543 3322 1547 3326
rect 1823 3322 1827 3326
rect 1863 3302 1867 3306
rect 1887 3302 1891 3306
rect 2007 3302 2011 3306
rect 2023 3302 2027 3306
rect 2151 3302 2155 3306
rect 2191 3302 2195 3306
rect 2303 3302 2307 3306
rect 2367 3302 2371 3306
rect 2463 3302 2467 3306
rect 2543 3302 2547 3306
rect 2631 3302 2635 3306
rect 2711 3302 2715 3306
rect 2799 3302 2803 3306
rect 2871 3302 2875 3306
rect 2967 3302 2971 3306
rect 3031 3302 3035 3306
rect 3135 3302 3139 3306
rect 3183 3302 3187 3306
rect 3311 3302 3315 3306
rect 3335 3302 3339 3306
rect 3479 3302 3483 3306
rect 3575 3302 3579 3306
rect 111 3250 115 3254
rect 199 3250 203 3254
rect 327 3250 331 3254
rect 367 3250 371 3254
rect 471 3250 475 3254
rect 503 3250 507 3254
rect 631 3250 635 3254
rect 639 3250 643 3254
rect 783 3250 787 3254
rect 799 3250 803 3254
rect 935 3250 939 3254
rect 975 3250 979 3254
rect 1095 3250 1099 3254
rect 1159 3250 1163 3254
rect 1255 3250 1259 3254
rect 1343 3250 1347 3254
rect 1415 3250 1419 3254
rect 1535 3250 1539 3254
rect 1575 3250 1579 3254
rect 1823 3250 1827 3254
rect 1863 3226 1867 3230
rect 1895 3226 1899 3230
rect 2015 3226 2019 3230
rect 2023 3226 2027 3230
rect 2159 3226 2163 3230
rect 2175 3226 2179 3230
rect 2311 3226 2315 3230
rect 2327 3226 2331 3230
rect 2463 3226 2467 3230
rect 2471 3226 2475 3230
rect 2599 3226 2603 3230
rect 2639 3226 2643 3230
rect 2735 3226 2739 3230
rect 2807 3226 2811 3230
rect 2871 3226 2875 3230
rect 2975 3226 2979 3230
rect 3015 3226 3019 3230
rect 3143 3226 3147 3230
rect 3167 3226 3171 3230
rect 3319 3226 3323 3230
rect 3327 3226 3331 3230
rect 3487 3226 3491 3230
rect 3575 3226 3579 3230
rect 111 3174 115 3178
rect 375 3174 379 3178
rect 447 3174 451 3178
rect 511 3174 515 3178
rect 559 3174 563 3178
rect 647 3174 651 3178
rect 687 3174 691 3178
rect 791 3174 795 3178
rect 823 3174 827 3178
rect 943 3174 947 3178
rect 975 3174 979 3178
rect 1103 3174 1107 3178
rect 1135 3174 1139 3178
rect 1263 3174 1267 3178
rect 1295 3174 1299 3178
rect 1423 3174 1427 3178
rect 1463 3174 1467 3178
rect 1583 3174 1587 3178
rect 1639 3174 1643 3178
rect 1823 3174 1827 3178
rect 1863 3154 1867 3158
rect 1887 3154 1891 3158
rect 2015 3154 2019 3158
rect 2047 3154 2051 3158
rect 2167 3154 2171 3158
rect 2199 3154 2203 3158
rect 2319 3154 2323 3158
rect 2351 3154 2355 3158
rect 2455 3154 2459 3158
rect 2511 3154 2515 3158
rect 2591 3154 2595 3158
rect 2679 3154 2683 3158
rect 2727 3154 2731 3158
rect 2863 3154 2867 3158
rect 2871 3154 2875 3158
rect 3007 3154 3011 3158
rect 3071 3154 3075 3158
rect 3159 3154 3163 3158
rect 3287 3154 3291 3158
rect 3319 3154 3323 3158
rect 3479 3154 3483 3158
rect 3575 3154 3579 3158
rect 111 3098 115 3102
rect 439 3098 443 3102
rect 551 3098 555 3102
rect 663 3098 667 3102
rect 679 3098 683 3102
rect 783 3098 787 3102
rect 815 3098 819 3102
rect 903 3098 907 3102
rect 967 3098 971 3102
rect 1031 3098 1035 3102
rect 1127 3098 1131 3102
rect 1159 3098 1163 3102
rect 1287 3098 1291 3102
rect 1423 3098 1427 3102
rect 1455 3098 1459 3102
rect 1559 3098 1563 3102
rect 1631 3098 1635 3102
rect 1695 3098 1699 3102
rect 1823 3098 1827 3102
rect 1863 3078 1867 3082
rect 1895 3078 1899 3082
rect 1919 3078 1923 3082
rect 2055 3078 2059 3082
rect 2087 3078 2091 3082
rect 2207 3078 2211 3082
rect 2279 3078 2283 3082
rect 2359 3078 2363 3082
rect 2487 3078 2491 3082
rect 2519 3078 2523 3082
rect 2687 3078 2691 3082
rect 2719 3078 2723 3082
rect 2879 3078 2883 3082
rect 2975 3078 2979 3082
rect 3079 3078 3083 3082
rect 3239 3078 3243 3082
rect 3295 3078 3299 3082
rect 3487 3078 3491 3082
rect 3575 3078 3579 3082
rect 111 3026 115 3030
rect 559 3026 563 3030
rect 575 3026 579 3030
rect 671 3026 675 3030
rect 703 3026 707 3030
rect 791 3026 795 3030
rect 831 3026 835 3030
rect 911 3026 915 3030
rect 967 3026 971 3030
rect 1039 3026 1043 3030
rect 1103 3026 1107 3030
rect 1167 3026 1171 3030
rect 1239 3026 1243 3030
rect 1295 3026 1299 3030
rect 1367 3026 1371 3030
rect 1431 3026 1435 3030
rect 1495 3026 1499 3030
rect 1567 3026 1571 3030
rect 1623 3026 1627 3030
rect 1703 3026 1707 3030
rect 1735 3026 1739 3030
rect 1823 3026 1827 3030
rect 1863 3006 1867 3010
rect 1911 3006 1915 3010
rect 2023 3006 2027 3010
rect 2079 3006 2083 3010
rect 2159 3006 2163 3010
rect 2271 3006 2275 3010
rect 2287 3006 2291 3010
rect 2415 3006 2419 3010
rect 2479 3006 2483 3010
rect 2535 3006 2539 3010
rect 2663 3006 2667 3010
rect 2711 3006 2715 3010
rect 2807 3006 2811 3010
rect 2967 3006 2971 3010
rect 3143 3006 3147 3010
rect 3231 3006 3235 3010
rect 3319 3006 3323 3010
rect 3479 3006 3483 3010
rect 3575 3006 3579 3010
rect 111 2958 115 2962
rect 495 2958 499 2962
rect 567 2958 571 2962
rect 639 2958 643 2962
rect 695 2958 699 2962
rect 783 2958 787 2962
rect 823 2958 827 2962
rect 919 2958 923 2962
rect 959 2958 963 2962
rect 1055 2958 1059 2962
rect 1095 2958 1099 2962
rect 1183 2958 1187 2962
rect 1231 2958 1235 2962
rect 1303 2958 1307 2962
rect 1359 2958 1363 2962
rect 1415 2958 1419 2962
rect 1487 2958 1491 2962
rect 1527 2958 1531 2962
rect 1615 2958 1619 2962
rect 1639 2958 1643 2962
rect 1727 2958 1731 2962
rect 1823 2958 1827 2962
rect 1863 2930 1867 2934
rect 1895 2930 1899 2934
rect 2031 2930 2035 2934
rect 2167 2930 2171 2934
rect 2175 2930 2179 2934
rect 2295 2930 2299 2934
rect 2423 2930 2427 2934
rect 2495 2930 2499 2934
rect 2543 2930 2547 2934
rect 2671 2930 2675 2934
rect 2815 2930 2819 2934
rect 2823 2930 2827 2934
rect 2975 2930 2979 2934
rect 3151 2930 3155 2934
rect 3167 2930 3171 2934
rect 3327 2930 3331 2934
rect 3487 2930 3491 2934
rect 3575 2930 3579 2934
rect 111 2886 115 2890
rect 327 2886 331 2890
rect 455 2886 459 2890
rect 503 2886 507 2890
rect 591 2886 595 2890
rect 647 2886 651 2890
rect 727 2886 731 2890
rect 791 2886 795 2890
rect 871 2886 875 2890
rect 927 2886 931 2890
rect 1007 2886 1011 2890
rect 1063 2886 1067 2890
rect 1143 2886 1147 2890
rect 1191 2886 1195 2890
rect 1279 2886 1283 2890
rect 1311 2886 1315 2890
rect 1415 2886 1419 2890
rect 1423 2886 1427 2890
rect 1535 2886 1539 2890
rect 1551 2886 1555 2890
rect 1647 2886 1651 2890
rect 1735 2886 1739 2890
rect 1823 2886 1827 2890
rect 1863 2862 1867 2866
rect 1887 2862 1891 2866
rect 2023 2862 2027 2866
rect 2167 2862 2171 2866
rect 2191 2862 2195 2866
rect 2359 2862 2363 2866
rect 2487 2862 2491 2866
rect 2519 2862 2523 2866
rect 2671 2862 2675 2866
rect 2807 2862 2811 2866
rect 2815 2862 2819 2866
rect 2935 2862 2939 2866
rect 3055 2862 3059 2866
rect 3159 2862 3163 2866
rect 3167 2862 3171 2866
rect 3279 2862 3283 2866
rect 3391 2862 3395 2866
rect 3479 2862 3483 2866
rect 3575 2862 3579 2866
rect 111 2810 115 2814
rect 167 2810 171 2814
rect 295 2810 299 2814
rect 319 2810 323 2814
rect 423 2810 427 2814
rect 447 2810 451 2814
rect 559 2810 563 2814
rect 583 2810 587 2814
rect 695 2810 699 2814
rect 719 2810 723 2814
rect 823 2810 827 2814
rect 863 2810 867 2814
rect 951 2810 955 2814
rect 999 2810 1003 2814
rect 1079 2810 1083 2814
rect 1135 2810 1139 2814
rect 1207 2810 1211 2814
rect 1271 2810 1275 2814
rect 1343 2810 1347 2814
rect 1407 2810 1411 2814
rect 1543 2810 1547 2814
rect 1823 2810 1827 2814
rect 1863 2794 1867 2798
rect 1895 2794 1899 2798
rect 2031 2794 2035 2798
rect 2063 2794 2067 2798
rect 2199 2794 2203 2798
rect 2255 2794 2259 2798
rect 2367 2794 2371 2798
rect 2439 2794 2443 2798
rect 2527 2794 2531 2798
rect 2615 2794 2619 2798
rect 2679 2794 2683 2798
rect 2783 2794 2787 2798
rect 2815 2794 2819 2798
rect 2935 2794 2939 2798
rect 2943 2794 2947 2798
rect 3063 2794 3067 2798
rect 3079 2794 3083 2798
rect 3175 2794 3179 2798
rect 3223 2794 3227 2798
rect 3287 2794 3291 2798
rect 3367 2794 3371 2798
rect 3399 2794 3403 2798
rect 3487 2794 3491 2798
rect 3575 2794 3579 2798
rect 111 2734 115 2738
rect 143 2734 147 2738
rect 175 2734 179 2738
rect 231 2734 235 2738
rect 303 2734 307 2738
rect 351 2734 355 2738
rect 431 2734 435 2738
rect 479 2734 483 2738
rect 567 2734 571 2738
rect 615 2734 619 2738
rect 703 2734 707 2738
rect 759 2734 763 2738
rect 831 2734 835 2738
rect 903 2734 907 2738
rect 959 2734 963 2738
rect 1047 2734 1051 2738
rect 1087 2734 1091 2738
rect 1215 2734 1219 2738
rect 1351 2734 1355 2738
rect 1823 2734 1827 2738
rect 1863 2722 1867 2726
rect 1887 2722 1891 2726
rect 2047 2722 2051 2726
rect 2055 2722 2059 2726
rect 2207 2722 2211 2726
rect 2247 2722 2251 2726
rect 2359 2722 2363 2726
rect 2431 2722 2435 2726
rect 2495 2722 2499 2726
rect 2607 2722 2611 2726
rect 2623 2722 2627 2726
rect 2743 2722 2747 2726
rect 2775 2722 2779 2726
rect 2863 2722 2867 2726
rect 2927 2722 2931 2726
rect 2983 2722 2987 2726
rect 3071 2722 3075 2726
rect 3103 2722 3107 2726
rect 3215 2722 3219 2726
rect 3359 2722 3363 2726
rect 3479 2722 3483 2726
rect 3575 2722 3579 2726
rect 111 2662 115 2666
rect 135 2662 139 2666
rect 223 2662 227 2666
rect 231 2662 235 2666
rect 343 2662 347 2666
rect 351 2662 355 2666
rect 471 2662 475 2666
rect 583 2662 587 2666
rect 607 2662 611 2666
rect 695 2662 699 2666
rect 751 2662 755 2666
rect 799 2662 803 2666
rect 895 2662 899 2666
rect 903 2662 907 2666
rect 999 2662 1003 2666
rect 1039 2662 1043 2666
rect 1103 2662 1107 2666
rect 1207 2662 1211 2666
rect 1311 2662 1315 2666
rect 1823 2662 1827 2666
rect 1863 2646 1867 2650
rect 1895 2646 1899 2650
rect 1999 2646 2003 2650
rect 2055 2646 2059 2650
rect 2119 2646 2123 2650
rect 2215 2646 2219 2650
rect 2239 2646 2243 2650
rect 2351 2646 2355 2650
rect 2367 2646 2371 2650
rect 2455 2646 2459 2650
rect 2503 2646 2507 2650
rect 2551 2646 2555 2650
rect 2631 2646 2635 2650
rect 2655 2646 2659 2650
rect 2751 2646 2755 2650
rect 2759 2646 2763 2650
rect 2863 2646 2867 2650
rect 2871 2646 2875 2650
rect 2991 2646 2995 2650
rect 3111 2646 3115 2650
rect 3575 2646 3579 2650
rect 111 2590 115 2594
rect 143 2590 147 2594
rect 239 2590 243 2594
rect 271 2590 275 2594
rect 359 2590 363 2594
rect 415 2590 419 2594
rect 479 2590 483 2594
rect 551 2590 555 2594
rect 591 2590 595 2594
rect 679 2590 683 2594
rect 703 2590 707 2594
rect 807 2590 811 2594
rect 911 2590 915 2594
rect 927 2590 931 2594
rect 1007 2590 1011 2594
rect 1047 2590 1051 2594
rect 1111 2590 1115 2594
rect 1175 2590 1179 2594
rect 1215 2590 1219 2594
rect 1319 2590 1323 2594
rect 1823 2590 1827 2594
rect 1863 2574 1867 2578
rect 1887 2574 1891 2578
rect 1991 2574 1995 2578
rect 2111 2574 2115 2578
rect 2231 2574 2235 2578
rect 2343 2574 2347 2578
rect 2351 2574 2355 2578
rect 2447 2574 2451 2578
rect 2471 2574 2475 2578
rect 2543 2574 2547 2578
rect 2591 2574 2595 2578
rect 2647 2574 2651 2578
rect 2711 2574 2715 2578
rect 2751 2574 2755 2578
rect 2831 2574 2835 2578
rect 2855 2574 2859 2578
rect 3575 2574 3579 2578
rect 111 2522 115 2526
rect 135 2522 139 2526
rect 263 2522 267 2526
rect 279 2522 283 2526
rect 407 2522 411 2526
rect 439 2522 443 2526
rect 543 2522 547 2526
rect 591 2522 595 2526
rect 671 2522 675 2526
rect 735 2522 739 2526
rect 799 2522 803 2526
rect 871 2522 875 2526
rect 919 2522 923 2526
rect 1007 2522 1011 2526
rect 1039 2522 1043 2526
rect 1143 2522 1147 2526
rect 1167 2522 1171 2526
rect 1279 2522 1283 2526
rect 1823 2522 1827 2526
rect 1863 2502 1867 2506
rect 1895 2502 1899 2506
rect 1999 2502 2003 2506
rect 2031 2502 2035 2506
rect 2119 2502 2123 2506
rect 2191 2502 2195 2506
rect 2239 2502 2243 2506
rect 2343 2502 2347 2506
rect 2359 2502 2363 2506
rect 2479 2502 2483 2506
rect 2487 2502 2491 2506
rect 2599 2502 2603 2506
rect 2623 2502 2627 2506
rect 2719 2502 2723 2506
rect 2751 2502 2755 2506
rect 2839 2502 2843 2506
rect 2879 2502 2883 2506
rect 3015 2502 3019 2506
rect 3575 2502 3579 2506
rect 111 2454 115 2458
rect 143 2454 147 2458
rect 191 2454 195 2458
rect 287 2454 291 2458
rect 319 2454 323 2458
rect 447 2454 451 2458
rect 455 2454 459 2458
rect 591 2454 595 2458
rect 599 2454 603 2458
rect 727 2454 731 2458
rect 743 2454 747 2458
rect 863 2454 867 2458
rect 879 2454 883 2458
rect 999 2454 1003 2458
rect 1015 2454 1019 2458
rect 1135 2454 1139 2458
rect 1151 2454 1155 2458
rect 1271 2454 1275 2458
rect 1287 2454 1291 2458
rect 1407 2454 1411 2458
rect 1823 2454 1827 2458
rect 1863 2434 1867 2438
rect 1887 2434 1891 2438
rect 2015 2434 2019 2438
rect 2023 2434 2027 2438
rect 2175 2434 2179 2438
rect 2183 2434 2187 2438
rect 2335 2434 2339 2438
rect 2479 2434 2483 2438
rect 2495 2434 2499 2438
rect 2615 2434 2619 2438
rect 2647 2434 2651 2438
rect 2743 2434 2747 2438
rect 2799 2434 2803 2438
rect 2871 2434 2875 2438
rect 2951 2434 2955 2438
rect 3007 2434 3011 2438
rect 3111 2434 3115 2438
rect 3575 2434 3579 2438
rect 111 2374 115 2378
rect 159 2374 163 2378
rect 183 2374 187 2378
rect 247 2374 251 2378
rect 311 2374 315 2378
rect 335 2374 339 2378
rect 439 2374 443 2378
rect 447 2374 451 2378
rect 559 2374 563 2378
rect 583 2374 587 2378
rect 687 2374 691 2378
rect 719 2374 723 2378
rect 815 2374 819 2378
rect 855 2374 859 2378
rect 951 2374 955 2378
rect 991 2374 995 2378
rect 1079 2374 1083 2378
rect 1127 2374 1131 2378
rect 1207 2374 1211 2378
rect 1263 2374 1267 2378
rect 1327 2374 1331 2378
rect 1399 2374 1403 2378
rect 1455 2374 1459 2378
rect 1583 2374 1587 2378
rect 1823 2374 1827 2378
rect 1863 2362 1867 2366
rect 1895 2362 1899 2366
rect 1927 2362 1931 2366
rect 2023 2362 2027 2366
rect 2087 2362 2091 2366
rect 2183 2362 2187 2366
rect 2247 2362 2251 2366
rect 2343 2362 2347 2366
rect 2407 2362 2411 2366
rect 2503 2362 2507 2366
rect 2559 2362 2563 2366
rect 2655 2362 2659 2366
rect 2703 2362 2707 2366
rect 2807 2362 2811 2366
rect 2831 2362 2835 2366
rect 2951 2362 2955 2366
rect 2959 2362 2963 2366
rect 3071 2362 3075 2366
rect 3119 2362 3123 2366
rect 3183 2362 3187 2366
rect 3287 2362 3291 2366
rect 3399 2362 3403 2366
rect 3487 2362 3491 2366
rect 3575 2362 3579 2366
rect 111 2298 115 2302
rect 167 2298 171 2302
rect 255 2298 259 2302
rect 343 2298 347 2302
rect 447 2298 451 2302
rect 567 2298 571 2302
rect 695 2298 699 2302
rect 823 2298 827 2302
rect 863 2298 867 2302
rect 959 2298 963 2302
rect 1023 2298 1027 2302
rect 1087 2298 1091 2302
rect 1175 2298 1179 2302
rect 1215 2298 1219 2302
rect 1319 2298 1323 2302
rect 1335 2298 1339 2302
rect 1463 2298 1467 2302
rect 1591 2298 1595 2302
rect 1599 2298 1603 2302
rect 1735 2298 1739 2302
rect 1823 2298 1827 2302
rect 1863 2290 1867 2294
rect 1919 2290 1923 2294
rect 1975 2290 1979 2294
rect 2079 2290 2083 2294
rect 2143 2290 2147 2294
rect 2239 2290 2243 2294
rect 2311 2290 2315 2294
rect 2399 2290 2403 2294
rect 2479 2290 2483 2294
rect 2551 2290 2555 2294
rect 2639 2290 2643 2294
rect 2695 2290 2699 2294
rect 2783 2290 2787 2294
rect 2823 2290 2827 2294
rect 2919 2290 2923 2294
rect 2943 2290 2947 2294
rect 3039 2290 3043 2294
rect 3063 2290 3067 2294
rect 3159 2290 3163 2294
rect 3175 2290 3179 2294
rect 3271 2290 3275 2294
rect 3279 2290 3283 2294
rect 3383 2290 3387 2294
rect 3391 2290 3395 2294
rect 3479 2290 3483 2294
rect 3575 2290 3579 2294
rect 111 2222 115 2226
rect 535 2222 539 2226
rect 687 2222 691 2226
rect 719 2222 723 2226
rect 855 2222 859 2226
rect 895 2222 899 2226
rect 1015 2222 1019 2226
rect 1071 2222 1075 2226
rect 1167 2222 1171 2226
rect 1239 2222 1243 2226
rect 1311 2222 1315 2226
rect 1407 2222 1411 2226
rect 1455 2222 1459 2226
rect 1575 2222 1579 2226
rect 1591 2222 1595 2226
rect 1727 2222 1731 2226
rect 1823 2222 1827 2226
rect 1863 2222 1867 2226
rect 1983 2222 1987 2226
rect 2007 2222 2011 2226
rect 2151 2222 2155 2226
rect 2167 2222 2171 2226
rect 2319 2222 2323 2226
rect 2335 2222 2339 2226
rect 2487 2222 2491 2226
rect 2519 2222 2523 2226
rect 2647 2222 2651 2226
rect 2711 2222 2715 2226
rect 2791 2222 2795 2226
rect 2903 2222 2907 2226
rect 2927 2222 2931 2226
rect 3047 2222 3051 2226
rect 3103 2222 3107 2226
rect 3167 2222 3171 2226
rect 3279 2222 3283 2226
rect 3303 2222 3307 2226
rect 3391 2222 3395 2226
rect 3487 2222 3491 2226
rect 3575 2222 3579 2226
rect 111 2154 115 2158
rect 495 2154 499 2158
rect 543 2154 547 2158
rect 623 2154 627 2158
rect 727 2154 731 2158
rect 759 2154 763 2158
rect 895 2154 899 2158
rect 903 2154 907 2158
rect 1039 2154 1043 2158
rect 1079 2154 1083 2158
rect 1183 2154 1187 2158
rect 1247 2154 1251 2158
rect 1327 2154 1331 2158
rect 1415 2154 1419 2158
rect 1471 2154 1475 2158
rect 1583 2154 1587 2158
rect 1623 2154 1627 2158
rect 1735 2154 1739 2158
rect 1823 2154 1827 2158
rect 1863 2146 1867 2150
rect 1999 2146 2003 2150
rect 2023 2146 2027 2150
rect 2159 2146 2163 2150
rect 2167 2146 2171 2150
rect 2319 2146 2323 2150
rect 2327 2146 2331 2150
rect 2471 2146 2475 2150
rect 2511 2146 2515 2150
rect 2615 2146 2619 2150
rect 2703 2146 2707 2150
rect 2759 2146 2763 2150
rect 2895 2146 2899 2150
rect 3023 2146 3027 2150
rect 3095 2146 3099 2150
rect 3143 2146 3147 2150
rect 3263 2146 3267 2150
rect 3295 2146 3299 2150
rect 3383 2146 3387 2150
rect 3479 2146 3483 2150
rect 3575 2146 3579 2150
rect 111 2082 115 2086
rect 319 2082 323 2086
rect 431 2082 435 2086
rect 487 2082 491 2086
rect 551 2082 555 2086
rect 615 2082 619 2086
rect 679 2082 683 2086
rect 751 2082 755 2086
rect 799 2082 803 2086
rect 887 2082 891 2086
rect 919 2082 923 2086
rect 1031 2082 1035 2086
rect 1039 2082 1043 2086
rect 1159 2082 1163 2086
rect 1175 2082 1179 2086
rect 1279 2082 1283 2086
rect 1319 2082 1323 2086
rect 1407 2082 1411 2086
rect 1463 2082 1467 2086
rect 1615 2082 1619 2086
rect 1823 2082 1827 2086
rect 1863 2074 1867 2078
rect 1983 2074 1987 2078
rect 2031 2074 2035 2078
rect 2143 2074 2147 2078
rect 2175 2074 2179 2078
rect 2311 2074 2315 2078
rect 2327 2074 2331 2078
rect 2471 2074 2475 2078
rect 2479 2074 2483 2078
rect 2623 2074 2627 2078
rect 2631 2074 2635 2078
rect 2767 2074 2771 2078
rect 2775 2074 2779 2078
rect 2903 2074 2907 2078
rect 2911 2074 2915 2078
rect 3031 2074 3035 2078
rect 3039 2074 3043 2078
rect 3151 2074 3155 2078
rect 3159 2074 3163 2078
rect 3271 2074 3275 2078
rect 3279 2074 3283 2078
rect 3391 2074 3395 2078
rect 3487 2074 3491 2078
rect 3575 2074 3579 2078
rect 111 2010 115 2014
rect 183 2010 187 2014
rect 295 2010 299 2014
rect 327 2010 331 2014
rect 415 2010 419 2014
rect 439 2010 443 2014
rect 535 2010 539 2014
rect 559 2010 563 2014
rect 655 2010 659 2014
rect 687 2010 691 2014
rect 775 2010 779 2014
rect 807 2010 811 2014
rect 895 2010 899 2014
rect 927 2010 931 2014
rect 1015 2010 1019 2014
rect 1047 2010 1051 2014
rect 1135 2010 1139 2014
rect 1167 2010 1171 2014
rect 1255 2010 1259 2014
rect 1287 2010 1291 2014
rect 1415 2010 1419 2014
rect 1823 2010 1827 2014
rect 1863 2006 1867 2010
rect 1887 2006 1891 2010
rect 1975 2006 1979 2010
rect 2031 2006 2035 2010
rect 2135 2006 2139 2010
rect 2199 2006 2203 2010
rect 2303 2006 2307 2010
rect 2375 2006 2379 2010
rect 2463 2006 2467 2010
rect 2543 2006 2547 2010
rect 2623 2006 2627 2010
rect 2711 2006 2715 2010
rect 2767 2006 2771 2010
rect 2871 2006 2875 2010
rect 2903 2006 2907 2010
rect 3031 2006 3035 2010
rect 3039 2006 3043 2010
rect 3151 2006 3155 2010
rect 3207 2006 3211 2010
rect 3271 2006 3275 2010
rect 3383 2006 3387 2010
rect 3479 2006 3483 2010
rect 3575 2006 3579 2010
rect 111 1938 115 1942
rect 135 1938 139 1942
rect 175 1938 179 1942
rect 223 1938 227 1942
rect 287 1938 291 1942
rect 351 1938 355 1942
rect 407 1938 411 1942
rect 495 1938 499 1942
rect 527 1938 531 1942
rect 647 1938 651 1942
rect 655 1938 659 1942
rect 767 1938 771 1942
rect 839 1938 843 1942
rect 887 1938 891 1942
rect 1007 1938 1011 1942
rect 1039 1938 1043 1942
rect 1127 1938 1131 1942
rect 1247 1938 1251 1942
rect 1463 1938 1467 1942
rect 1823 1938 1827 1942
rect 1863 1930 1867 1934
rect 1895 1930 1899 1934
rect 1991 1930 1995 1934
rect 2039 1930 2043 1934
rect 2119 1930 2123 1934
rect 2207 1930 2211 1934
rect 2255 1930 2259 1934
rect 2383 1930 2387 1934
rect 2511 1930 2515 1934
rect 2551 1930 2555 1934
rect 2631 1930 2635 1934
rect 2719 1930 2723 1934
rect 2751 1930 2755 1934
rect 2879 1930 2883 1934
rect 3007 1930 3011 1934
rect 3047 1930 3051 1934
rect 3215 1930 3219 1934
rect 3575 1930 3579 1934
rect 111 1862 115 1866
rect 143 1862 147 1866
rect 231 1862 235 1866
rect 271 1862 275 1866
rect 359 1862 363 1866
rect 415 1862 419 1866
rect 503 1862 507 1866
rect 559 1862 563 1866
rect 663 1862 667 1866
rect 695 1862 699 1866
rect 823 1862 827 1866
rect 847 1862 851 1866
rect 943 1862 947 1866
rect 1047 1862 1051 1866
rect 1055 1862 1059 1866
rect 1159 1862 1163 1866
rect 1255 1862 1259 1866
rect 1263 1862 1267 1866
rect 1359 1862 1363 1866
rect 1455 1862 1459 1866
rect 1471 1862 1475 1866
rect 1551 1862 1555 1866
rect 1647 1862 1651 1866
rect 1735 1862 1739 1866
rect 1823 1862 1827 1866
rect 1863 1854 1867 1858
rect 1887 1854 1891 1858
rect 1983 1854 1987 1858
rect 2111 1854 2115 1858
rect 2223 1854 2227 1858
rect 2247 1854 2251 1858
rect 2359 1854 2363 1858
rect 2375 1854 2379 1858
rect 2495 1854 2499 1858
rect 2503 1854 2507 1858
rect 2623 1854 2627 1858
rect 2743 1854 2747 1858
rect 2863 1854 2867 1858
rect 2871 1854 2875 1858
rect 2991 1854 2995 1858
rect 2999 1854 3003 1858
rect 3575 1854 3579 1858
rect 111 1782 115 1786
rect 135 1782 139 1786
rect 263 1782 267 1786
rect 303 1782 307 1786
rect 407 1782 411 1786
rect 495 1782 499 1786
rect 551 1782 555 1786
rect 687 1782 691 1786
rect 815 1782 819 1786
rect 871 1782 875 1786
rect 935 1782 939 1786
rect 1047 1782 1051 1786
rect 1151 1782 1155 1786
rect 1215 1782 1219 1786
rect 1255 1782 1259 1786
rect 1351 1782 1355 1786
rect 1375 1782 1379 1786
rect 1447 1782 1451 1786
rect 1535 1782 1539 1786
rect 1543 1782 1547 1786
rect 1639 1782 1643 1786
rect 1703 1782 1707 1786
rect 1727 1782 1731 1786
rect 1823 1782 1827 1786
rect 1863 1782 1867 1786
rect 2231 1782 2235 1786
rect 2271 1782 2275 1786
rect 2359 1782 2363 1786
rect 2367 1782 2371 1786
rect 2455 1782 2459 1786
rect 2503 1782 2507 1786
rect 2559 1782 2563 1786
rect 2631 1782 2635 1786
rect 2663 1782 2667 1786
rect 2751 1782 2755 1786
rect 2759 1782 2763 1786
rect 2863 1782 2867 1786
rect 2871 1782 2875 1786
rect 2967 1782 2971 1786
rect 2999 1782 3003 1786
rect 3071 1782 3075 1786
rect 3175 1782 3179 1786
rect 3575 1782 3579 1786
rect 111 1710 115 1714
rect 143 1710 147 1714
rect 287 1710 291 1714
rect 311 1710 315 1714
rect 471 1710 475 1714
rect 503 1710 507 1714
rect 655 1710 659 1714
rect 695 1710 699 1714
rect 839 1710 843 1714
rect 879 1710 883 1714
rect 1023 1710 1027 1714
rect 1055 1710 1059 1714
rect 1191 1710 1195 1714
rect 1223 1710 1227 1714
rect 1359 1710 1363 1714
rect 1383 1710 1387 1714
rect 1527 1710 1531 1714
rect 1543 1710 1547 1714
rect 1695 1710 1699 1714
rect 1711 1710 1715 1714
rect 1823 1710 1827 1714
rect 1863 1710 1867 1714
rect 2247 1710 2251 1714
rect 2263 1710 2267 1714
rect 2351 1710 2355 1714
rect 2367 1710 2371 1714
rect 2447 1710 2451 1714
rect 2495 1710 2499 1714
rect 2551 1710 2555 1714
rect 2623 1710 2627 1714
rect 2655 1710 2659 1714
rect 2751 1710 2755 1714
rect 2759 1710 2763 1714
rect 2855 1710 2859 1714
rect 2887 1710 2891 1714
rect 2959 1710 2963 1714
rect 3015 1710 3019 1714
rect 3063 1710 3067 1714
rect 3135 1710 3139 1714
rect 3167 1710 3171 1714
rect 3247 1710 3251 1714
rect 3367 1710 3371 1714
rect 3479 1710 3483 1714
rect 3575 1710 3579 1714
rect 111 1634 115 1638
rect 135 1634 139 1638
rect 271 1634 275 1638
rect 279 1634 283 1638
rect 447 1634 451 1638
rect 463 1634 467 1638
rect 631 1634 635 1638
rect 647 1634 651 1638
rect 815 1634 819 1638
rect 831 1634 835 1638
rect 991 1634 995 1638
rect 1015 1634 1019 1638
rect 1151 1634 1155 1638
rect 1183 1634 1187 1638
rect 1303 1634 1307 1638
rect 1351 1634 1355 1638
rect 1455 1634 1459 1638
rect 1519 1634 1523 1638
rect 1599 1634 1603 1638
rect 1687 1634 1691 1638
rect 1727 1634 1731 1638
rect 1823 1634 1827 1638
rect 1863 1638 1867 1642
rect 2151 1638 2155 1642
rect 2255 1638 2259 1642
rect 2343 1638 2347 1642
rect 2375 1638 2379 1642
rect 2503 1638 2507 1642
rect 2527 1638 2531 1642
rect 2631 1638 2635 1642
rect 2703 1638 2707 1642
rect 2767 1638 2771 1642
rect 2871 1638 2875 1642
rect 2895 1638 2899 1642
rect 3023 1638 3027 1642
rect 3031 1638 3035 1642
rect 3143 1638 3147 1642
rect 3191 1638 3195 1642
rect 3255 1638 3259 1642
rect 3351 1638 3355 1642
rect 3375 1638 3379 1642
rect 3487 1638 3491 1642
rect 3575 1638 3579 1642
rect 111 1566 115 1570
rect 143 1566 147 1570
rect 271 1566 275 1570
rect 279 1566 283 1570
rect 431 1566 435 1570
rect 455 1566 459 1570
rect 599 1566 603 1570
rect 639 1566 643 1570
rect 767 1566 771 1570
rect 823 1566 827 1570
rect 935 1566 939 1570
rect 999 1566 1003 1570
rect 1103 1566 1107 1570
rect 1159 1566 1163 1570
rect 1263 1566 1267 1570
rect 1311 1566 1315 1570
rect 1423 1566 1427 1570
rect 1463 1566 1467 1570
rect 1591 1566 1595 1570
rect 1607 1566 1611 1570
rect 1735 1566 1739 1570
rect 1823 1566 1827 1570
rect 1863 1570 1867 1574
rect 2087 1570 2091 1574
rect 2143 1570 2147 1574
rect 2279 1570 2283 1574
rect 2335 1570 2339 1574
rect 2455 1570 2459 1574
rect 2519 1570 2523 1574
rect 2623 1570 2627 1574
rect 2695 1570 2699 1574
rect 2791 1570 2795 1574
rect 2863 1570 2867 1574
rect 2951 1570 2955 1574
rect 3023 1570 3027 1574
rect 3111 1570 3115 1574
rect 3183 1570 3187 1574
rect 3271 1570 3275 1574
rect 3343 1570 3347 1574
rect 3431 1570 3435 1574
rect 3479 1570 3483 1574
rect 3575 1570 3579 1574
rect 111 1494 115 1498
rect 135 1494 139 1498
rect 183 1494 187 1498
rect 263 1494 267 1498
rect 327 1494 331 1498
rect 423 1494 427 1498
rect 471 1494 475 1498
rect 591 1494 595 1498
rect 607 1494 611 1498
rect 743 1494 747 1498
rect 759 1494 763 1498
rect 871 1494 875 1498
rect 927 1494 931 1498
rect 991 1494 995 1498
rect 1095 1494 1099 1498
rect 1119 1494 1123 1498
rect 1247 1494 1251 1498
rect 1255 1494 1259 1498
rect 1375 1494 1379 1498
rect 1415 1494 1419 1498
rect 1583 1494 1587 1498
rect 1727 1494 1731 1498
rect 1823 1494 1827 1498
rect 1863 1494 1867 1498
rect 1895 1494 1899 1498
rect 1991 1494 1995 1498
rect 2095 1494 2099 1498
rect 2119 1494 2123 1498
rect 2247 1494 2251 1498
rect 2287 1494 2291 1498
rect 2383 1494 2387 1498
rect 2463 1494 2467 1498
rect 2535 1494 2539 1498
rect 2631 1494 2635 1498
rect 2703 1494 2707 1498
rect 2799 1494 2803 1498
rect 2887 1494 2891 1498
rect 2959 1494 2963 1498
rect 3087 1494 3091 1498
rect 3119 1494 3123 1498
rect 3279 1494 3283 1498
rect 3295 1494 3299 1498
rect 3439 1494 3443 1498
rect 3487 1494 3491 1498
rect 3575 1494 3579 1498
rect 111 1418 115 1422
rect 191 1418 195 1422
rect 199 1418 203 1422
rect 335 1418 339 1422
rect 463 1418 467 1422
rect 479 1418 483 1422
rect 583 1418 587 1422
rect 615 1418 619 1422
rect 703 1418 707 1422
rect 751 1418 755 1422
rect 815 1418 819 1422
rect 879 1418 883 1422
rect 919 1418 923 1422
rect 999 1418 1003 1422
rect 1015 1418 1019 1422
rect 1119 1418 1123 1422
rect 1127 1418 1131 1422
rect 1223 1418 1227 1422
rect 1255 1418 1259 1422
rect 1327 1418 1331 1422
rect 1383 1418 1387 1422
rect 1823 1418 1827 1422
rect 1863 1422 1867 1426
rect 1887 1422 1891 1426
rect 1975 1422 1979 1426
rect 1983 1422 1987 1426
rect 2071 1422 2075 1426
rect 2111 1422 2115 1426
rect 2183 1422 2187 1426
rect 2239 1422 2243 1426
rect 2303 1422 2307 1426
rect 2375 1422 2379 1426
rect 2439 1422 2443 1426
rect 2527 1422 2531 1426
rect 2607 1422 2611 1426
rect 2695 1422 2699 1426
rect 2807 1422 2811 1426
rect 2879 1422 2883 1426
rect 3031 1422 3035 1426
rect 3079 1422 3083 1426
rect 3263 1422 3267 1426
rect 3287 1422 3291 1426
rect 3479 1422 3483 1426
rect 3575 1422 3579 1426
rect 111 1346 115 1350
rect 191 1346 195 1350
rect 231 1346 235 1350
rect 327 1346 331 1350
rect 383 1346 387 1350
rect 455 1346 459 1350
rect 543 1346 547 1350
rect 575 1346 579 1350
rect 695 1346 699 1350
rect 703 1346 707 1350
rect 807 1346 811 1350
rect 871 1346 875 1350
rect 911 1346 915 1350
rect 1007 1346 1011 1350
rect 1039 1346 1043 1350
rect 1111 1346 1115 1350
rect 1207 1346 1211 1350
rect 1215 1346 1219 1350
rect 1319 1346 1323 1350
rect 1375 1346 1379 1350
rect 1823 1346 1827 1350
rect 1863 1350 1867 1354
rect 1895 1350 1899 1354
rect 1983 1350 1987 1354
rect 2079 1350 2083 1354
rect 2103 1350 2107 1354
rect 2191 1350 2195 1354
rect 2223 1350 2227 1354
rect 2311 1350 2315 1354
rect 2359 1350 2363 1354
rect 2447 1350 2451 1354
rect 2511 1350 2515 1354
rect 2615 1350 2619 1354
rect 2687 1350 2691 1354
rect 2815 1350 2819 1354
rect 2871 1350 2875 1354
rect 3039 1350 3043 1354
rect 3071 1350 3075 1354
rect 3271 1350 3275 1354
rect 3279 1350 3283 1354
rect 3487 1350 3491 1354
rect 3575 1350 3579 1354
rect 111 1278 115 1282
rect 215 1278 219 1282
rect 239 1278 243 1282
rect 359 1278 363 1282
rect 391 1278 395 1282
rect 519 1278 523 1282
rect 551 1278 555 1282
rect 679 1278 683 1282
rect 711 1278 715 1282
rect 839 1278 843 1282
rect 879 1278 883 1282
rect 999 1278 1003 1282
rect 1047 1278 1051 1282
rect 1151 1278 1155 1282
rect 1215 1278 1219 1282
rect 1295 1278 1299 1282
rect 1383 1278 1387 1282
rect 1439 1278 1443 1282
rect 1591 1278 1595 1282
rect 1823 1278 1827 1282
rect 1863 1270 1867 1274
rect 1887 1270 1891 1274
rect 1975 1270 1979 1274
rect 2055 1270 2059 1274
rect 2095 1270 2099 1274
rect 2143 1270 2147 1274
rect 2215 1270 2219 1274
rect 2239 1270 2243 1274
rect 2335 1270 2339 1274
rect 2351 1270 2355 1274
rect 2431 1270 2435 1274
rect 2503 1270 2507 1274
rect 2551 1270 2555 1274
rect 2679 1270 2683 1274
rect 2687 1270 2691 1274
rect 2855 1270 2859 1274
rect 2863 1270 2867 1274
rect 3039 1270 3043 1274
rect 3063 1270 3067 1274
rect 3231 1270 3235 1274
rect 3271 1270 3275 1274
rect 3431 1270 3435 1274
rect 3479 1270 3483 1274
rect 3575 1270 3579 1274
rect 111 1202 115 1206
rect 135 1202 139 1206
rect 207 1202 211 1206
rect 271 1202 275 1206
rect 351 1202 355 1206
rect 423 1202 427 1206
rect 511 1202 515 1206
rect 575 1202 579 1206
rect 671 1202 675 1206
rect 727 1202 731 1206
rect 831 1202 835 1206
rect 887 1202 891 1206
rect 991 1202 995 1206
rect 1055 1202 1059 1206
rect 1143 1202 1147 1206
rect 1231 1202 1235 1206
rect 1287 1202 1291 1206
rect 1415 1202 1419 1206
rect 1431 1202 1435 1206
rect 1583 1202 1587 1206
rect 1599 1202 1603 1206
rect 1823 1202 1827 1206
rect 1863 1198 1867 1202
rect 2039 1198 2043 1202
rect 2063 1198 2067 1202
rect 2151 1198 2155 1202
rect 2247 1198 2251 1202
rect 2279 1198 2283 1202
rect 2343 1198 2347 1202
rect 2415 1198 2419 1202
rect 2439 1198 2443 1202
rect 2559 1198 2563 1202
rect 2695 1198 2699 1202
rect 2711 1198 2715 1202
rect 2863 1198 2867 1202
rect 3015 1198 3019 1202
rect 3047 1198 3051 1202
rect 3167 1198 3171 1202
rect 3239 1198 3243 1202
rect 3327 1198 3331 1202
rect 3439 1198 3443 1202
rect 3487 1198 3491 1202
rect 3575 1198 3579 1202
rect 111 1134 115 1138
rect 143 1134 147 1138
rect 279 1134 283 1138
rect 295 1134 299 1138
rect 431 1134 435 1138
rect 479 1134 483 1138
rect 583 1134 587 1138
rect 663 1134 667 1138
rect 735 1134 739 1138
rect 847 1134 851 1138
rect 895 1134 899 1138
rect 1031 1134 1035 1138
rect 1063 1134 1067 1138
rect 1207 1134 1211 1138
rect 1239 1134 1243 1138
rect 1391 1134 1395 1138
rect 1423 1134 1427 1138
rect 1575 1134 1579 1138
rect 1607 1134 1611 1138
rect 1735 1134 1739 1138
rect 1823 1134 1827 1138
rect 1863 1118 1867 1122
rect 1943 1118 1947 1122
rect 2031 1118 2035 1122
rect 2087 1118 2091 1122
rect 2143 1118 2147 1122
rect 2231 1118 2235 1122
rect 2271 1118 2275 1122
rect 2383 1118 2387 1122
rect 2407 1118 2411 1122
rect 2535 1118 2539 1122
rect 2551 1118 2555 1122
rect 2687 1118 2691 1122
rect 2703 1118 2707 1122
rect 2839 1118 2843 1122
rect 2855 1118 2859 1122
rect 2991 1118 2995 1122
rect 3007 1118 3011 1122
rect 3151 1118 3155 1122
rect 3159 1118 3163 1122
rect 3319 1118 3323 1122
rect 3479 1118 3483 1122
rect 3575 1118 3579 1122
rect 111 1066 115 1070
rect 135 1066 139 1070
rect 271 1066 275 1070
rect 287 1066 291 1070
rect 431 1066 435 1070
rect 471 1066 475 1070
rect 583 1066 587 1070
rect 655 1066 659 1070
rect 735 1066 739 1070
rect 839 1066 843 1070
rect 887 1066 891 1070
rect 1023 1066 1027 1070
rect 1047 1066 1051 1070
rect 1199 1066 1203 1070
rect 1215 1066 1219 1070
rect 1383 1066 1387 1070
rect 1559 1066 1563 1070
rect 1567 1066 1571 1070
rect 1727 1066 1731 1070
rect 1823 1066 1827 1070
rect 1863 1038 1867 1042
rect 1919 1038 1923 1042
rect 1951 1038 1955 1042
rect 2095 1038 2099 1042
rect 2127 1038 2131 1042
rect 2239 1038 2243 1042
rect 2327 1038 2331 1042
rect 2391 1038 2395 1042
rect 2519 1038 2523 1042
rect 2543 1038 2547 1042
rect 2695 1038 2699 1042
rect 2847 1038 2851 1042
rect 2863 1038 2867 1042
rect 2999 1038 3003 1042
rect 3023 1038 3027 1042
rect 3159 1038 3163 1042
rect 3183 1038 3187 1042
rect 3327 1038 3331 1042
rect 3343 1038 3347 1042
rect 3487 1038 3491 1042
rect 3575 1038 3579 1042
rect 111 994 115 998
rect 143 994 147 998
rect 279 994 283 998
rect 287 994 291 998
rect 439 994 443 998
rect 463 994 467 998
rect 591 994 595 998
rect 647 994 651 998
rect 743 994 747 998
rect 823 994 827 998
rect 895 994 899 998
rect 999 994 1003 998
rect 1055 994 1059 998
rect 1167 994 1171 998
rect 1223 994 1227 998
rect 1327 994 1331 998
rect 1391 994 1395 998
rect 1487 994 1491 998
rect 1567 994 1571 998
rect 1655 994 1659 998
rect 1735 994 1739 998
rect 1823 994 1827 998
rect 1863 966 1867 970
rect 1887 966 1891 970
rect 1911 966 1915 970
rect 2071 966 2075 970
rect 2119 966 2123 970
rect 2263 966 2267 970
rect 2319 966 2323 970
rect 2455 966 2459 970
rect 2511 966 2515 970
rect 2631 966 2635 970
rect 2687 966 2691 970
rect 2799 966 2803 970
rect 2855 966 2859 970
rect 2951 966 2955 970
rect 3015 966 3019 970
rect 3095 966 3099 970
rect 3175 966 3179 970
rect 3231 966 3235 970
rect 3335 966 3339 970
rect 3367 966 3371 970
rect 3479 966 3483 970
rect 3575 966 3579 970
rect 111 918 115 922
rect 135 918 139 922
rect 271 918 275 922
rect 279 918 283 922
rect 439 918 443 922
rect 455 918 459 922
rect 607 918 611 922
rect 639 918 643 922
rect 775 918 779 922
rect 815 918 819 922
rect 935 918 939 922
rect 991 918 995 922
rect 1095 918 1099 922
rect 1159 918 1163 922
rect 1247 918 1251 922
rect 1319 918 1323 922
rect 1399 918 1403 922
rect 1479 918 1483 922
rect 1551 918 1555 922
rect 1647 918 1651 922
rect 1823 918 1827 922
rect 1863 890 1867 894
rect 1895 890 1899 894
rect 2023 890 2027 894
rect 2079 890 2083 894
rect 2183 890 2187 894
rect 2271 890 2275 894
rect 2351 890 2355 894
rect 2463 890 2467 894
rect 2519 890 2523 894
rect 2639 890 2643 894
rect 2687 890 2691 894
rect 2807 890 2811 894
rect 2839 890 2843 894
rect 2959 890 2963 894
rect 2983 890 2987 894
rect 3103 890 3107 894
rect 3119 890 3123 894
rect 3239 890 3243 894
rect 3247 890 3251 894
rect 3375 890 3379 894
rect 3487 890 3491 894
rect 3575 890 3579 894
rect 111 850 115 854
rect 143 850 147 854
rect 279 850 283 854
rect 287 850 291 854
rect 447 850 451 854
rect 463 850 467 854
rect 615 850 619 854
rect 639 850 643 854
rect 783 850 787 854
rect 807 850 811 854
rect 943 850 947 854
rect 983 850 987 854
rect 1103 850 1107 854
rect 1159 850 1163 854
rect 1255 850 1259 854
rect 1335 850 1339 854
rect 1407 850 1411 854
rect 1511 850 1515 854
rect 1559 850 1563 854
rect 1823 850 1827 854
rect 1863 814 1867 818
rect 1887 814 1891 818
rect 2015 814 2019 818
rect 2071 814 2075 818
rect 2175 814 2179 818
rect 2263 814 2267 818
rect 2343 814 2347 818
rect 2447 814 2451 818
rect 2511 814 2515 818
rect 2623 814 2627 818
rect 2679 814 2683 818
rect 2791 814 2795 818
rect 2831 814 2835 818
rect 2943 814 2947 818
rect 2975 814 2979 818
rect 3087 814 3091 818
rect 3111 814 3115 818
rect 3223 814 3227 818
rect 3239 814 3243 818
rect 3359 814 3363 818
rect 3367 814 3371 818
rect 3479 814 3483 818
rect 3575 814 3579 818
rect 111 778 115 782
rect 135 778 139 782
rect 271 778 275 782
rect 279 778 283 782
rect 439 778 443 782
rect 455 778 459 782
rect 607 778 611 782
rect 631 778 635 782
rect 775 778 779 782
rect 799 778 803 782
rect 935 778 939 782
rect 975 778 979 782
rect 1087 778 1091 782
rect 1151 778 1155 782
rect 1239 778 1243 782
rect 1327 778 1331 782
rect 1391 778 1395 782
rect 1503 778 1507 782
rect 1551 778 1555 782
rect 1823 778 1827 782
rect 1863 746 1867 750
rect 1895 746 1899 750
rect 2071 746 2075 750
rect 2079 746 2083 750
rect 2263 746 2267 750
rect 2271 746 2275 750
rect 2447 746 2451 750
rect 2455 746 2459 750
rect 2623 746 2627 750
rect 2631 746 2635 750
rect 2799 746 2803 750
rect 2951 746 2955 750
rect 2975 746 2979 750
rect 3095 746 3099 750
rect 3151 746 3155 750
rect 3231 746 3235 750
rect 3327 746 3331 750
rect 3367 746 3371 750
rect 3487 746 3491 750
rect 3575 746 3579 750
rect 111 706 115 710
rect 143 706 147 710
rect 279 706 283 710
rect 287 706 291 710
rect 447 706 451 710
rect 455 706 459 710
rect 615 706 619 710
rect 623 706 627 710
rect 783 706 787 710
rect 791 706 795 710
rect 943 706 947 710
rect 959 706 963 710
rect 1095 706 1099 710
rect 1119 706 1123 710
rect 1247 706 1251 710
rect 1279 706 1283 710
rect 1399 706 1403 710
rect 1439 706 1443 710
rect 1559 706 1563 710
rect 1599 706 1603 710
rect 1823 706 1827 710
rect 1863 674 1867 678
rect 1887 674 1891 678
rect 1975 674 1979 678
rect 2063 674 2067 678
rect 2095 674 2099 678
rect 2223 674 2227 678
rect 2255 674 2259 678
rect 2351 674 2355 678
rect 2439 674 2443 678
rect 2479 674 2483 678
rect 2615 674 2619 678
rect 2767 674 2771 678
rect 2791 674 2795 678
rect 2935 674 2939 678
rect 2967 674 2971 678
rect 3119 674 3123 678
rect 3143 674 3147 678
rect 3311 674 3315 678
rect 3319 674 3323 678
rect 3479 674 3483 678
rect 3575 674 3579 678
rect 111 630 115 634
rect 135 630 139 634
rect 279 630 283 634
rect 287 630 291 634
rect 447 630 451 634
rect 455 630 459 634
rect 615 630 619 634
rect 631 630 635 634
rect 783 630 787 634
rect 799 630 803 634
rect 951 630 955 634
rect 967 630 971 634
rect 1111 630 1115 634
rect 1119 630 1123 634
rect 1271 630 1275 634
rect 1415 630 1419 634
rect 1431 630 1435 634
rect 1559 630 1563 634
rect 1591 630 1595 634
rect 1711 630 1715 634
rect 1823 630 1827 634
rect 1863 602 1867 606
rect 1895 602 1899 606
rect 1983 602 1987 606
rect 2047 602 2051 606
rect 2103 602 2107 606
rect 2215 602 2219 606
rect 2231 602 2235 606
rect 2359 602 2363 606
rect 2391 602 2395 606
rect 2487 602 2491 606
rect 2583 602 2587 606
rect 2623 602 2627 606
rect 2775 602 2779 606
rect 2799 602 2803 606
rect 2943 602 2947 606
rect 3023 602 3027 606
rect 3127 602 3131 606
rect 3255 602 3259 606
rect 3319 602 3323 606
rect 3487 602 3491 606
rect 3575 602 3579 606
rect 111 558 115 562
rect 143 558 147 562
rect 151 558 155 562
rect 295 558 299 562
rect 311 558 315 562
rect 463 558 467 562
rect 471 558 475 562
rect 631 558 635 562
rect 639 558 643 562
rect 783 558 787 562
rect 807 558 811 562
rect 927 558 931 562
rect 975 558 979 562
rect 1063 558 1067 562
rect 1127 558 1131 562
rect 1191 558 1195 562
rect 1279 558 1283 562
rect 1311 558 1315 562
rect 1423 558 1427 562
rect 1535 558 1539 562
rect 1567 558 1571 562
rect 1647 558 1651 562
rect 1719 558 1723 562
rect 1735 558 1739 562
rect 1823 558 1827 562
rect 1863 526 1867 530
rect 1887 526 1891 530
rect 2039 526 2043 530
rect 2191 526 2195 530
rect 2207 526 2211 530
rect 2279 526 2283 530
rect 2375 526 2379 530
rect 2383 526 2387 530
rect 2487 526 2491 530
rect 2575 526 2579 530
rect 2631 526 2635 530
rect 2791 526 2795 530
rect 2807 526 2811 530
rect 3007 526 3011 530
rect 3015 526 3019 530
rect 3215 526 3219 530
rect 3247 526 3251 530
rect 3431 526 3435 530
rect 3479 526 3483 530
rect 3575 526 3579 530
rect 111 482 115 486
rect 143 482 147 486
rect 159 482 163 486
rect 303 482 307 486
rect 311 482 315 486
rect 463 482 467 486
rect 615 482 619 486
rect 623 482 627 486
rect 759 482 763 486
rect 775 482 779 486
rect 887 482 891 486
rect 919 482 923 486
rect 1007 482 1011 486
rect 1055 482 1059 486
rect 1127 482 1131 486
rect 1183 482 1187 486
rect 1239 482 1243 486
rect 1303 482 1307 486
rect 1343 482 1347 486
rect 1415 482 1419 486
rect 1439 482 1443 486
rect 1527 482 1531 486
rect 1543 482 1547 486
rect 1639 482 1643 486
rect 1727 482 1731 486
rect 1823 482 1827 486
rect 1863 450 1867 454
rect 1895 450 1899 454
rect 2039 450 2043 454
rect 2199 450 2203 454
rect 2207 450 2211 454
rect 2287 450 2291 454
rect 2383 450 2387 454
rect 2495 450 2499 454
rect 2575 450 2579 454
rect 2639 450 2643 454
rect 2783 450 2787 454
rect 2815 450 2819 454
rect 3007 450 3011 454
rect 3015 450 3019 454
rect 3223 450 3227 454
rect 3239 450 3243 454
rect 3439 450 3443 454
rect 3471 450 3475 454
rect 3575 450 3579 454
rect 111 414 115 418
rect 151 414 155 418
rect 167 414 171 418
rect 271 414 275 418
rect 319 414 323 418
rect 407 414 411 418
rect 471 414 475 418
rect 551 414 555 418
rect 623 414 627 418
rect 711 414 715 418
rect 767 414 771 418
rect 887 414 891 418
rect 895 414 899 418
rect 1015 414 1019 418
rect 1063 414 1067 418
rect 1135 414 1139 418
rect 1247 414 1251 418
rect 1351 414 1355 418
rect 1439 414 1443 418
rect 1447 414 1451 418
rect 1551 414 1555 418
rect 1639 414 1643 418
rect 1647 414 1651 418
rect 1735 414 1739 418
rect 1823 414 1827 418
rect 1863 382 1867 386
rect 1887 382 1891 386
rect 1975 382 1979 386
rect 2031 382 2035 386
rect 2063 382 2067 386
rect 2151 382 2155 386
rect 2199 382 2203 386
rect 2263 382 2267 386
rect 2375 382 2379 386
rect 2383 382 2387 386
rect 2519 382 2523 386
rect 2567 382 2571 386
rect 2671 382 2675 386
rect 2775 382 2779 386
rect 2847 382 2851 386
rect 2999 382 3003 386
rect 3031 382 3035 386
rect 3231 382 3235 386
rect 3431 382 3435 386
rect 3463 382 3467 386
rect 3575 382 3579 386
rect 111 330 115 334
rect 135 330 139 334
rect 143 330 147 334
rect 223 330 227 334
rect 263 330 267 334
rect 311 330 315 334
rect 399 330 403 334
rect 487 330 491 334
rect 543 330 547 334
rect 575 330 579 334
rect 663 330 667 334
rect 703 330 707 334
rect 751 330 755 334
rect 839 330 843 334
rect 879 330 883 334
rect 927 330 931 334
rect 1015 330 1019 334
rect 1055 330 1059 334
rect 1103 330 1107 334
rect 1191 330 1195 334
rect 1239 330 1243 334
rect 1287 330 1291 334
rect 1383 330 1387 334
rect 1431 330 1435 334
rect 1479 330 1483 334
rect 1575 330 1579 334
rect 1631 330 1635 334
rect 1671 330 1675 334
rect 1823 330 1827 334
rect 1863 314 1867 318
rect 1895 314 1899 318
rect 1983 314 1987 318
rect 2071 314 2075 318
rect 2159 314 2163 318
rect 2247 314 2251 318
rect 2271 314 2275 318
rect 2359 314 2363 318
rect 2391 314 2395 318
rect 2471 314 2475 318
rect 2527 314 2531 318
rect 2583 314 2587 318
rect 2679 314 2683 318
rect 2695 314 2699 318
rect 2807 314 2811 318
rect 2855 314 2859 318
rect 2919 314 2923 318
rect 3039 314 3043 318
rect 3159 314 3163 318
rect 3239 314 3243 318
rect 3439 314 3443 318
rect 3575 314 3579 318
rect 111 258 115 262
rect 143 258 147 262
rect 231 258 235 262
rect 319 258 323 262
rect 407 258 411 262
rect 495 258 499 262
rect 583 258 587 262
rect 671 258 675 262
rect 759 258 763 262
rect 847 258 851 262
rect 935 258 939 262
rect 1023 258 1027 262
rect 1111 258 1115 262
rect 1199 258 1203 262
rect 1287 258 1291 262
rect 1295 258 1299 262
rect 1375 258 1379 262
rect 1391 258 1395 262
rect 1463 258 1467 262
rect 1487 258 1491 262
rect 1551 258 1555 262
rect 1583 258 1587 262
rect 1639 258 1643 262
rect 1679 258 1683 262
rect 1727 258 1731 262
rect 1823 258 1827 262
rect 1863 246 1867 250
rect 1887 246 1891 250
rect 1975 246 1979 250
rect 2063 246 2067 250
rect 2151 246 2155 250
rect 2239 246 2243 250
rect 2263 246 2267 250
rect 2351 246 2355 250
rect 2399 246 2403 250
rect 2463 246 2467 250
rect 2535 246 2539 250
rect 2575 246 2579 250
rect 2679 246 2683 250
rect 2687 246 2691 250
rect 2799 246 2803 250
rect 2815 246 2819 250
rect 2911 246 2915 250
rect 2951 246 2955 250
rect 3031 246 3035 250
rect 3087 246 3091 250
rect 3151 246 3155 250
rect 3223 246 3227 250
rect 3359 246 3363 250
rect 3479 246 3483 250
rect 3575 246 3579 250
rect 111 190 115 194
rect 135 190 139 194
rect 223 190 227 194
rect 311 190 315 194
rect 399 190 403 194
rect 487 190 491 194
rect 575 190 579 194
rect 663 190 667 194
rect 751 190 755 194
rect 839 190 843 194
rect 927 190 931 194
rect 1015 190 1019 194
rect 1103 190 1107 194
rect 1191 190 1195 194
rect 1279 190 1283 194
rect 1367 190 1371 194
rect 1455 190 1459 194
rect 1543 190 1547 194
rect 1631 190 1635 194
rect 1719 190 1723 194
rect 1823 190 1827 194
rect 1863 146 1867 150
rect 1895 146 1899 150
rect 1983 146 1987 150
rect 2071 146 2075 150
rect 2159 146 2163 150
rect 2271 146 2275 150
rect 2407 146 2411 150
rect 2543 146 2547 150
rect 2687 146 2691 150
rect 2783 146 2787 150
rect 2823 146 2827 150
rect 2871 146 2875 150
rect 2959 146 2963 150
rect 3047 146 3051 150
rect 3095 146 3099 150
rect 3135 146 3139 150
rect 3223 146 3227 150
rect 3231 146 3235 150
rect 3311 146 3315 150
rect 3367 146 3371 150
rect 3399 146 3403 150
rect 3487 146 3491 150
rect 3575 146 3579 150
rect 1863 78 1867 82
rect 2775 78 2779 82
rect 2863 78 2867 82
rect 2951 78 2955 82
rect 3039 78 3043 82
rect 3127 78 3131 82
rect 3215 78 3219 82
rect 3303 78 3307 82
rect 3391 78 3395 82
rect 3479 78 3483 82
rect 3575 78 3579 82
<< m4 >>
rect 84 3665 85 3671
rect 91 3670 1835 3671
rect 91 3666 111 3670
rect 115 3666 135 3670
rect 139 3666 223 3670
rect 227 3666 1823 3670
rect 1827 3666 1835 3670
rect 91 3665 1835 3666
rect 1841 3665 1842 3671
rect 1834 3607 1835 3613
rect 1841 3607 1866 3613
rect 96 3597 97 3603
rect 103 3602 1847 3603
rect 103 3598 111 3602
rect 115 3598 143 3602
rect 147 3598 231 3602
rect 235 3598 319 3602
rect 323 3598 407 3602
rect 411 3598 495 3602
rect 499 3598 1823 3602
rect 1827 3598 1847 3602
rect 103 3597 1847 3598
rect 1853 3597 1854 3603
rect 1860 3595 1866 3607
rect 1860 3594 3599 3595
rect 1860 3590 1863 3594
rect 1867 3590 1887 3594
rect 1891 3590 1975 3594
rect 1979 3590 2063 3594
rect 2067 3590 2151 3594
rect 2155 3590 2239 3594
rect 2243 3590 2327 3594
rect 2331 3590 2431 3594
rect 2435 3590 2535 3594
rect 2539 3590 2631 3594
rect 2635 3590 2727 3594
rect 2731 3590 2823 3594
rect 2827 3590 2919 3594
rect 2923 3590 3015 3594
rect 3019 3590 3119 3594
rect 3123 3590 3223 3594
rect 3227 3590 3575 3594
rect 3579 3590 3599 3594
rect 1860 3589 3599 3590
rect 3605 3589 3606 3595
rect 84 3529 85 3535
rect 91 3534 1835 3535
rect 91 3530 111 3534
rect 115 3530 135 3534
rect 139 3530 223 3534
rect 227 3530 247 3534
rect 251 3530 311 3534
rect 315 3530 375 3534
rect 379 3530 399 3534
rect 403 3530 487 3534
rect 491 3530 503 3534
rect 507 3530 623 3534
rect 627 3530 743 3534
rect 747 3530 863 3534
rect 867 3530 975 3534
rect 979 3530 1079 3534
rect 1083 3530 1175 3534
rect 1179 3530 1271 3534
rect 1275 3530 1367 3534
rect 1371 3530 1471 3534
rect 1475 3530 1575 3534
rect 1579 3530 1823 3534
rect 1827 3530 1835 3534
rect 91 3529 1835 3530
rect 1841 3529 1842 3535
rect 1846 3521 1847 3527
rect 1853 3526 3611 3527
rect 1853 3522 1863 3526
rect 1867 3522 1895 3526
rect 1899 3522 1983 3526
rect 1987 3522 2071 3526
rect 2075 3522 2103 3526
rect 2107 3522 2159 3526
rect 2163 3522 2231 3526
rect 2235 3522 2247 3526
rect 2251 3522 2335 3526
rect 2339 3522 2367 3526
rect 2371 3522 2439 3526
rect 2443 3522 2511 3526
rect 2515 3522 2543 3526
rect 2547 3522 2639 3526
rect 2643 3522 2655 3526
rect 2659 3522 2735 3526
rect 2739 3522 2791 3526
rect 2795 3522 2831 3526
rect 2835 3522 2927 3526
rect 2931 3522 2935 3526
rect 2939 3522 3023 3526
rect 3027 3522 3079 3526
rect 3083 3522 3127 3526
rect 3131 3522 3223 3526
rect 3227 3522 3231 3526
rect 3235 3522 3575 3526
rect 3579 3522 3611 3526
rect 1853 3521 3611 3522
rect 3617 3521 3618 3527
rect 96 3461 97 3467
rect 103 3466 1847 3467
rect 103 3462 111 3466
rect 115 3462 175 3466
rect 179 3462 255 3466
rect 259 3462 303 3466
rect 307 3462 383 3466
rect 387 3462 447 3466
rect 451 3462 511 3466
rect 515 3462 591 3466
rect 595 3462 631 3466
rect 635 3462 743 3466
rect 747 3462 751 3466
rect 755 3462 871 3466
rect 875 3462 895 3466
rect 899 3462 983 3466
rect 987 3462 1039 3466
rect 1043 3462 1087 3466
rect 1091 3462 1183 3466
rect 1187 3462 1279 3466
rect 1283 3462 1327 3466
rect 1331 3462 1375 3466
rect 1379 3462 1479 3466
rect 1483 3462 1583 3466
rect 1587 3462 1823 3466
rect 1827 3462 1847 3466
rect 103 3461 1847 3462
rect 1853 3461 1854 3467
rect 1834 3445 1835 3451
rect 1841 3450 3599 3451
rect 1841 3446 1863 3450
rect 1867 3446 1887 3450
rect 1891 3446 1975 3450
rect 1979 3446 2023 3450
rect 2027 3446 2095 3450
rect 2099 3446 2191 3450
rect 2195 3446 2223 3450
rect 2227 3446 2359 3450
rect 2363 3446 2367 3450
rect 2371 3446 2503 3450
rect 2507 3446 2543 3450
rect 2547 3446 2647 3450
rect 2651 3446 2711 3450
rect 2715 3446 2783 3450
rect 2787 3446 2871 3450
rect 2875 3446 2927 3450
rect 2931 3446 3031 3450
rect 3035 3446 3071 3450
rect 3075 3446 3191 3450
rect 3195 3446 3215 3450
rect 3219 3446 3359 3450
rect 3363 3446 3575 3450
rect 3579 3446 3599 3450
rect 1841 3445 3599 3446
rect 3605 3445 3606 3451
rect 84 3393 85 3399
rect 91 3398 1835 3399
rect 91 3394 111 3398
rect 115 3394 135 3398
rect 139 3394 167 3398
rect 171 3394 263 3398
rect 267 3394 295 3398
rect 299 3394 407 3398
rect 411 3394 439 3398
rect 443 3394 567 3398
rect 571 3394 583 3398
rect 587 3394 727 3398
rect 731 3394 735 3398
rect 739 3394 887 3398
rect 891 3394 1031 3398
rect 1035 3394 1047 3398
rect 1051 3394 1175 3398
rect 1179 3394 1207 3398
rect 1211 3394 1319 3398
rect 1323 3394 1367 3398
rect 1371 3394 1471 3398
rect 1475 3394 1527 3398
rect 1531 3394 1823 3398
rect 1827 3394 1835 3398
rect 91 3393 1835 3394
rect 1841 3393 1842 3399
rect 1846 3369 1847 3375
rect 1853 3374 3611 3375
rect 1853 3370 1863 3374
rect 1867 3370 1895 3374
rect 1899 3370 2031 3374
rect 2035 3370 2199 3374
rect 2203 3370 2375 3374
rect 2379 3370 2551 3374
rect 2555 3370 2719 3374
rect 2723 3370 2879 3374
rect 2883 3370 3039 3374
rect 3043 3370 3191 3374
rect 3195 3370 3199 3374
rect 3203 3370 3343 3374
rect 3347 3370 3367 3374
rect 3371 3370 3487 3374
rect 3491 3370 3575 3374
rect 3579 3370 3611 3374
rect 1853 3369 3611 3370
rect 3617 3369 3618 3375
rect 96 3321 97 3327
rect 103 3326 1847 3327
rect 103 3322 111 3326
rect 115 3322 143 3326
rect 147 3322 207 3326
rect 211 3322 271 3326
rect 275 3322 335 3326
rect 339 3322 415 3326
rect 419 3322 479 3326
rect 483 3322 575 3326
rect 579 3322 639 3326
rect 643 3322 735 3326
rect 739 3322 807 3326
rect 811 3322 895 3326
rect 899 3322 983 3326
rect 987 3322 1055 3326
rect 1059 3322 1167 3326
rect 1171 3322 1215 3326
rect 1219 3322 1351 3326
rect 1355 3322 1375 3326
rect 1379 3322 1535 3326
rect 1539 3322 1543 3326
rect 1547 3322 1823 3326
rect 1827 3322 1847 3326
rect 103 3321 1847 3322
rect 1853 3321 1854 3327
rect 1834 3301 1835 3307
rect 1841 3306 3599 3307
rect 1841 3302 1863 3306
rect 1867 3302 1887 3306
rect 1891 3302 2007 3306
rect 2011 3302 2023 3306
rect 2027 3302 2151 3306
rect 2155 3302 2191 3306
rect 2195 3302 2303 3306
rect 2307 3302 2367 3306
rect 2371 3302 2463 3306
rect 2467 3302 2543 3306
rect 2547 3302 2631 3306
rect 2635 3302 2711 3306
rect 2715 3302 2799 3306
rect 2803 3302 2871 3306
rect 2875 3302 2967 3306
rect 2971 3302 3031 3306
rect 3035 3302 3135 3306
rect 3139 3302 3183 3306
rect 3187 3302 3311 3306
rect 3315 3302 3335 3306
rect 3339 3302 3479 3306
rect 3483 3302 3575 3306
rect 3579 3302 3599 3306
rect 1841 3301 3599 3302
rect 3605 3301 3606 3307
rect 84 3249 85 3255
rect 91 3254 1835 3255
rect 91 3250 111 3254
rect 115 3250 199 3254
rect 203 3250 327 3254
rect 331 3250 367 3254
rect 371 3250 471 3254
rect 475 3250 503 3254
rect 507 3250 631 3254
rect 635 3250 639 3254
rect 643 3250 783 3254
rect 787 3250 799 3254
rect 803 3250 935 3254
rect 939 3250 975 3254
rect 979 3250 1095 3254
rect 1099 3250 1159 3254
rect 1163 3250 1255 3254
rect 1259 3250 1343 3254
rect 1347 3250 1415 3254
rect 1419 3250 1535 3254
rect 1539 3250 1575 3254
rect 1579 3250 1823 3254
rect 1827 3250 1835 3254
rect 91 3249 1835 3250
rect 1841 3249 1842 3255
rect 1846 3225 1847 3231
rect 1853 3230 3611 3231
rect 1853 3226 1863 3230
rect 1867 3226 1895 3230
rect 1899 3226 2015 3230
rect 2019 3226 2023 3230
rect 2027 3226 2159 3230
rect 2163 3226 2175 3230
rect 2179 3226 2311 3230
rect 2315 3226 2327 3230
rect 2331 3226 2463 3230
rect 2467 3226 2471 3230
rect 2475 3226 2599 3230
rect 2603 3226 2639 3230
rect 2643 3226 2735 3230
rect 2739 3226 2807 3230
rect 2811 3226 2871 3230
rect 2875 3226 2975 3230
rect 2979 3226 3015 3230
rect 3019 3226 3143 3230
rect 3147 3226 3167 3230
rect 3171 3226 3319 3230
rect 3323 3226 3327 3230
rect 3331 3226 3487 3230
rect 3491 3226 3575 3230
rect 3579 3226 3611 3230
rect 1853 3225 3611 3226
rect 3617 3225 3618 3231
rect 96 3173 97 3179
rect 103 3178 1847 3179
rect 103 3174 111 3178
rect 115 3174 375 3178
rect 379 3174 447 3178
rect 451 3174 511 3178
rect 515 3174 559 3178
rect 563 3174 647 3178
rect 651 3174 687 3178
rect 691 3174 791 3178
rect 795 3174 823 3178
rect 827 3174 943 3178
rect 947 3174 975 3178
rect 979 3174 1103 3178
rect 1107 3174 1135 3178
rect 1139 3174 1263 3178
rect 1267 3174 1295 3178
rect 1299 3174 1423 3178
rect 1427 3174 1463 3178
rect 1467 3174 1583 3178
rect 1587 3174 1639 3178
rect 1643 3174 1823 3178
rect 1827 3174 1847 3178
rect 103 3173 1847 3174
rect 1853 3173 1854 3179
rect 1834 3153 1835 3159
rect 1841 3158 3599 3159
rect 1841 3154 1863 3158
rect 1867 3154 1887 3158
rect 1891 3154 2015 3158
rect 2019 3154 2047 3158
rect 2051 3154 2167 3158
rect 2171 3154 2199 3158
rect 2203 3154 2319 3158
rect 2323 3154 2351 3158
rect 2355 3154 2455 3158
rect 2459 3154 2511 3158
rect 2515 3154 2591 3158
rect 2595 3154 2679 3158
rect 2683 3154 2727 3158
rect 2731 3154 2863 3158
rect 2867 3154 2871 3158
rect 2875 3154 3007 3158
rect 3011 3154 3071 3158
rect 3075 3154 3159 3158
rect 3163 3154 3287 3158
rect 3291 3154 3319 3158
rect 3323 3154 3479 3158
rect 3483 3154 3575 3158
rect 3579 3154 3599 3158
rect 1841 3153 3599 3154
rect 3605 3153 3606 3159
rect 84 3097 85 3103
rect 91 3102 1835 3103
rect 91 3098 111 3102
rect 115 3098 439 3102
rect 443 3098 551 3102
rect 555 3098 663 3102
rect 667 3098 679 3102
rect 683 3098 783 3102
rect 787 3098 815 3102
rect 819 3098 903 3102
rect 907 3098 967 3102
rect 971 3098 1031 3102
rect 1035 3098 1127 3102
rect 1131 3098 1159 3102
rect 1163 3098 1287 3102
rect 1291 3098 1423 3102
rect 1427 3098 1455 3102
rect 1459 3098 1559 3102
rect 1563 3098 1631 3102
rect 1635 3098 1695 3102
rect 1699 3098 1823 3102
rect 1827 3098 1835 3102
rect 91 3097 1835 3098
rect 1841 3097 1842 3103
rect 1846 3077 1847 3083
rect 1853 3082 3611 3083
rect 1853 3078 1863 3082
rect 1867 3078 1895 3082
rect 1899 3078 1919 3082
rect 1923 3078 2055 3082
rect 2059 3078 2087 3082
rect 2091 3078 2207 3082
rect 2211 3078 2279 3082
rect 2283 3078 2359 3082
rect 2363 3078 2487 3082
rect 2491 3078 2519 3082
rect 2523 3078 2687 3082
rect 2691 3078 2719 3082
rect 2723 3078 2879 3082
rect 2883 3078 2975 3082
rect 2979 3078 3079 3082
rect 3083 3078 3239 3082
rect 3243 3078 3295 3082
rect 3299 3078 3487 3082
rect 3491 3078 3575 3082
rect 3579 3078 3611 3082
rect 1853 3077 3611 3078
rect 3617 3077 3618 3083
rect 96 3025 97 3031
rect 103 3030 1847 3031
rect 103 3026 111 3030
rect 115 3026 559 3030
rect 563 3026 575 3030
rect 579 3026 671 3030
rect 675 3026 703 3030
rect 707 3026 791 3030
rect 795 3026 831 3030
rect 835 3026 911 3030
rect 915 3026 967 3030
rect 971 3026 1039 3030
rect 1043 3026 1103 3030
rect 1107 3026 1167 3030
rect 1171 3026 1239 3030
rect 1243 3026 1295 3030
rect 1299 3026 1367 3030
rect 1371 3026 1431 3030
rect 1435 3026 1495 3030
rect 1499 3026 1567 3030
rect 1571 3026 1623 3030
rect 1627 3026 1703 3030
rect 1707 3026 1735 3030
rect 1739 3026 1823 3030
rect 1827 3026 1847 3030
rect 103 3025 1847 3026
rect 1853 3025 1854 3031
rect 1834 3005 1835 3011
rect 1841 3010 3599 3011
rect 1841 3006 1863 3010
rect 1867 3006 1911 3010
rect 1915 3006 2023 3010
rect 2027 3006 2079 3010
rect 2083 3006 2159 3010
rect 2163 3006 2271 3010
rect 2275 3006 2287 3010
rect 2291 3006 2415 3010
rect 2419 3006 2479 3010
rect 2483 3006 2535 3010
rect 2539 3006 2663 3010
rect 2667 3006 2711 3010
rect 2715 3006 2807 3010
rect 2811 3006 2967 3010
rect 2971 3006 3143 3010
rect 3147 3006 3231 3010
rect 3235 3006 3319 3010
rect 3323 3006 3479 3010
rect 3483 3006 3575 3010
rect 3579 3006 3599 3010
rect 1841 3005 3599 3006
rect 3605 3005 3606 3011
rect 84 2957 85 2963
rect 91 2962 1835 2963
rect 91 2958 111 2962
rect 115 2958 495 2962
rect 499 2958 567 2962
rect 571 2958 639 2962
rect 643 2958 695 2962
rect 699 2958 783 2962
rect 787 2958 823 2962
rect 827 2958 919 2962
rect 923 2958 959 2962
rect 963 2958 1055 2962
rect 1059 2958 1095 2962
rect 1099 2958 1183 2962
rect 1187 2958 1231 2962
rect 1235 2958 1303 2962
rect 1307 2958 1359 2962
rect 1363 2958 1415 2962
rect 1419 2958 1487 2962
rect 1491 2958 1527 2962
rect 1531 2958 1615 2962
rect 1619 2958 1639 2962
rect 1643 2958 1727 2962
rect 1731 2958 1823 2962
rect 1827 2958 1835 2962
rect 91 2957 1835 2958
rect 1841 2957 1842 2963
rect 1846 2929 1847 2935
rect 1853 2934 3611 2935
rect 1853 2930 1863 2934
rect 1867 2930 1895 2934
rect 1899 2930 2031 2934
rect 2035 2930 2167 2934
rect 2171 2930 2175 2934
rect 2179 2930 2295 2934
rect 2299 2930 2423 2934
rect 2427 2930 2495 2934
rect 2499 2930 2543 2934
rect 2547 2930 2671 2934
rect 2675 2930 2815 2934
rect 2819 2930 2823 2934
rect 2827 2930 2975 2934
rect 2979 2930 3151 2934
rect 3155 2930 3167 2934
rect 3171 2930 3327 2934
rect 3331 2930 3487 2934
rect 3491 2930 3575 2934
rect 3579 2930 3611 2934
rect 1853 2929 3611 2930
rect 3617 2929 3618 2935
rect 96 2885 97 2891
rect 103 2890 1847 2891
rect 103 2886 111 2890
rect 115 2886 327 2890
rect 331 2886 455 2890
rect 459 2886 503 2890
rect 507 2886 591 2890
rect 595 2886 647 2890
rect 651 2886 727 2890
rect 731 2886 791 2890
rect 795 2886 871 2890
rect 875 2886 927 2890
rect 931 2886 1007 2890
rect 1011 2886 1063 2890
rect 1067 2886 1143 2890
rect 1147 2886 1191 2890
rect 1195 2886 1279 2890
rect 1283 2886 1311 2890
rect 1315 2886 1415 2890
rect 1419 2886 1423 2890
rect 1427 2886 1535 2890
rect 1539 2886 1551 2890
rect 1555 2886 1647 2890
rect 1651 2886 1735 2890
rect 1739 2886 1823 2890
rect 1827 2886 1847 2890
rect 103 2885 1847 2886
rect 1853 2885 1854 2891
rect 1834 2861 1835 2867
rect 1841 2866 3599 2867
rect 1841 2862 1863 2866
rect 1867 2862 1887 2866
rect 1891 2862 2023 2866
rect 2027 2862 2167 2866
rect 2171 2862 2191 2866
rect 2195 2862 2359 2866
rect 2363 2862 2487 2866
rect 2491 2862 2519 2866
rect 2523 2862 2671 2866
rect 2675 2862 2807 2866
rect 2811 2862 2815 2866
rect 2819 2862 2935 2866
rect 2939 2862 3055 2866
rect 3059 2862 3159 2866
rect 3163 2862 3167 2866
rect 3171 2862 3279 2866
rect 3283 2862 3391 2866
rect 3395 2862 3479 2866
rect 3483 2862 3575 2866
rect 3579 2862 3599 2866
rect 1841 2861 3599 2862
rect 3605 2861 3606 2867
rect 84 2809 85 2815
rect 91 2814 1835 2815
rect 91 2810 111 2814
rect 115 2810 167 2814
rect 171 2810 295 2814
rect 299 2810 319 2814
rect 323 2810 423 2814
rect 427 2810 447 2814
rect 451 2810 559 2814
rect 563 2810 583 2814
rect 587 2810 695 2814
rect 699 2810 719 2814
rect 723 2810 823 2814
rect 827 2810 863 2814
rect 867 2810 951 2814
rect 955 2810 999 2814
rect 1003 2810 1079 2814
rect 1083 2810 1135 2814
rect 1139 2810 1207 2814
rect 1211 2810 1271 2814
rect 1275 2810 1343 2814
rect 1347 2810 1407 2814
rect 1411 2810 1543 2814
rect 1547 2810 1823 2814
rect 1827 2810 1835 2814
rect 91 2809 1835 2810
rect 1841 2809 1842 2815
rect 1846 2793 1847 2799
rect 1853 2798 3611 2799
rect 1853 2794 1863 2798
rect 1867 2794 1895 2798
rect 1899 2794 2031 2798
rect 2035 2794 2063 2798
rect 2067 2794 2199 2798
rect 2203 2794 2255 2798
rect 2259 2794 2367 2798
rect 2371 2794 2439 2798
rect 2443 2794 2527 2798
rect 2531 2794 2615 2798
rect 2619 2794 2679 2798
rect 2683 2794 2783 2798
rect 2787 2794 2815 2798
rect 2819 2794 2935 2798
rect 2939 2794 2943 2798
rect 2947 2794 3063 2798
rect 3067 2794 3079 2798
rect 3083 2794 3175 2798
rect 3179 2794 3223 2798
rect 3227 2794 3287 2798
rect 3291 2794 3367 2798
rect 3371 2794 3399 2798
rect 3403 2794 3487 2798
rect 3491 2794 3575 2798
rect 3579 2794 3611 2798
rect 1853 2793 3611 2794
rect 3617 2793 3618 2799
rect 96 2733 97 2739
rect 103 2738 1847 2739
rect 103 2734 111 2738
rect 115 2734 143 2738
rect 147 2734 175 2738
rect 179 2734 231 2738
rect 235 2734 303 2738
rect 307 2734 351 2738
rect 355 2734 431 2738
rect 435 2734 479 2738
rect 483 2734 567 2738
rect 571 2734 615 2738
rect 619 2734 703 2738
rect 707 2734 759 2738
rect 763 2734 831 2738
rect 835 2734 903 2738
rect 907 2734 959 2738
rect 963 2734 1047 2738
rect 1051 2734 1087 2738
rect 1091 2734 1215 2738
rect 1219 2734 1351 2738
rect 1355 2734 1823 2738
rect 1827 2734 1847 2738
rect 103 2733 1847 2734
rect 1853 2733 1854 2739
rect 1834 2721 1835 2727
rect 1841 2726 3599 2727
rect 1841 2722 1863 2726
rect 1867 2722 1887 2726
rect 1891 2722 2047 2726
rect 2051 2722 2055 2726
rect 2059 2722 2207 2726
rect 2211 2722 2247 2726
rect 2251 2722 2359 2726
rect 2363 2722 2431 2726
rect 2435 2722 2495 2726
rect 2499 2722 2607 2726
rect 2611 2722 2623 2726
rect 2627 2722 2743 2726
rect 2747 2722 2775 2726
rect 2779 2722 2863 2726
rect 2867 2722 2927 2726
rect 2931 2722 2983 2726
rect 2987 2722 3071 2726
rect 3075 2722 3103 2726
rect 3107 2722 3215 2726
rect 3219 2722 3359 2726
rect 3363 2722 3479 2726
rect 3483 2722 3575 2726
rect 3579 2722 3599 2726
rect 1841 2721 3599 2722
rect 3605 2721 3606 2727
rect 84 2661 85 2667
rect 91 2666 1835 2667
rect 91 2662 111 2666
rect 115 2662 135 2666
rect 139 2662 223 2666
rect 227 2662 231 2666
rect 235 2662 343 2666
rect 347 2662 351 2666
rect 355 2662 471 2666
rect 475 2662 583 2666
rect 587 2662 607 2666
rect 611 2662 695 2666
rect 699 2662 751 2666
rect 755 2662 799 2666
rect 803 2662 895 2666
rect 899 2662 903 2666
rect 907 2662 999 2666
rect 1003 2662 1039 2666
rect 1043 2662 1103 2666
rect 1107 2662 1207 2666
rect 1211 2662 1311 2666
rect 1315 2662 1823 2666
rect 1827 2662 1835 2666
rect 91 2661 1835 2662
rect 1841 2661 1842 2667
rect 1846 2645 1847 2651
rect 1853 2650 3611 2651
rect 1853 2646 1863 2650
rect 1867 2646 1895 2650
rect 1899 2646 1999 2650
rect 2003 2646 2055 2650
rect 2059 2646 2119 2650
rect 2123 2646 2215 2650
rect 2219 2646 2239 2650
rect 2243 2646 2351 2650
rect 2355 2646 2367 2650
rect 2371 2646 2455 2650
rect 2459 2646 2503 2650
rect 2507 2646 2551 2650
rect 2555 2646 2631 2650
rect 2635 2646 2655 2650
rect 2659 2646 2751 2650
rect 2755 2646 2759 2650
rect 2763 2646 2863 2650
rect 2867 2646 2871 2650
rect 2875 2646 2991 2650
rect 2995 2646 3111 2650
rect 3115 2646 3575 2650
rect 3579 2646 3611 2650
rect 1853 2645 3611 2646
rect 3617 2645 3618 2651
rect 96 2589 97 2595
rect 103 2594 1847 2595
rect 103 2590 111 2594
rect 115 2590 143 2594
rect 147 2590 239 2594
rect 243 2590 271 2594
rect 275 2590 359 2594
rect 363 2590 415 2594
rect 419 2590 479 2594
rect 483 2590 551 2594
rect 555 2590 591 2594
rect 595 2590 679 2594
rect 683 2590 703 2594
rect 707 2590 807 2594
rect 811 2590 911 2594
rect 915 2590 927 2594
rect 931 2590 1007 2594
rect 1011 2590 1047 2594
rect 1051 2590 1111 2594
rect 1115 2590 1175 2594
rect 1179 2590 1215 2594
rect 1219 2590 1319 2594
rect 1323 2590 1823 2594
rect 1827 2590 1847 2594
rect 103 2589 1847 2590
rect 1853 2589 1854 2595
rect 1834 2573 1835 2579
rect 1841 2578 3599 2579
rect 1841 2574 1863 2578
rect 1867 2574 1887 2578
rect 1891 2574 1991 2578
rect 1995 2574 2111 2578
rect 2115 2574 2231 2578
rect 2235 2574 2343 2578
rect 2347 2574 2351 2578
rect 2355 2574 2447 2578
rect 2451 2574 2471 2578
rect 2475 2574 2543 2578
rect 2547 2574 2591 2578
rect 2595 2574 2647 2578
rect 2651 2574 2711 2578
rect 2715 2574 2751 2578
rect 2755 2574 2831 2578
rect 2835 2574 2855 2578
rect 2859 2574 3575 2578
rect 3579 2574 3599 2578
rect 1841 2573 3599 2574
rect 3605 2573 3606 2579
rect 84 2521 85 2527
rect 91 2526 1835 2527
rect 91 2522 111 2526
rect 115 2522 135 2526
rect 139 2522 263 2526
rect 267 2522 279 2526
rect 283 2522 407 2526
rect 411 2522 439 2526
rect 443 2522 543 2526
rect 547 2522 591 2526
rect 595 2522 671 2526
rect 675 2522 735 2526
rect 739 2522 799 2526
rect 803 2522 871 2526
rect 875 2522 919 2526
rect 923 2522 1007 2526
rect 1011 2522 1039 2526
rect 1043 2522 1143 2526
rect 1147 2522 1167 2526
rect 1171 2522 1279 2526
rect 1283 2522 1823 2526
rect 1827 2522 1835 2526
rect 91 2521 1835 2522
rect 1841 2521 1842 2527
rect 1846 2501 1847 2507
rect 1853 2506 3611 2507
rect 1853 2502 1863 2506
rect 1867 2502 1895 2506
rect 1899 2502 1999 2506
rect 2003 2502 2031 2506
rect 2035 2502 2119 2506
rect 2123 2502 2191 2506
rect 2195 2502 2239 2506
rect 2243 2502 2343 2506
rect 2347 2502 2359 2506
rect 2363 2502 2479 2506
rect 2483 2502 2487 2506
rect 2491 2502 2599 2506
rect 2603 2502 2623 2506
rect 2627 2502 2719 2506
rect 2723 2502 2751 2506
rect 2755 2502 2839 2506
rect 2843 2502 2879 2506
rect 2883 2502 3015 2506
rect 3019 2502 3575 2506
rect 3579 2502 3611 2506
rect 1853 2501 3611 2502
rect 3617 2501 3618 2507
rect 96 2453 97 2459
rect 103 2458 1847 2459
rect 103 2454 111 2458
rect 115 2454 143 2458
rect 147 2454 191 2458
rect 195 2454 287 2458
rect 291 2454 319 2458
rect 323 2454 447 2458
rect 451 2454 455 2458
rect 459 2454 591 2458
rect 595 2454 599 2458
rect 603 2454 727 2458
rect 731 2454 743 2458
rect 747 2454 863 2458
rect 867 2454 879 2458
rect 883 2454 999 2458
rect 1003 2454 1015 2458
rect 1019 2454 1135 2458
rect 1139 2454 1151 2458
rect 1155 2454 1271 2458
rect 1275 2454 1287 2458
rect 1291 2454 1407 2458
rect 1411 2454 1823 2458
rect 1827 2454 1847 2458
rect 103 2453 1847 2454
rect 1853 2453 1854 2459
rect 1834 2433 1835 2439
rect 1841 2438 3599 2439
rect 1841 2434 1863 2438
rect 1867 2434 1887 2438
rect 1891 2434 2015 2438
rect 2019 2434 2023 2438
rect 2027 2434 2175 2438
rect 2179 2434 2183 2438
rect 2187 2434 2335 2438
rect 2339 2434 2479 2438
rect 2483 2434 2495 2438
rect 2499 2434 2615 2438
rect 2619 2434 2647 2438
rect 2651 2434 2743 2438
rect 2747 2434 2799 2438
rect 2803 2434 2871 2438
rect 2875 2434 2951 2438
rect 2955 2434 3007 2438
rect 3011 2434 3111 2438
rect 3115 2434 3575 2438
rect 3579 2434 3599 2438
rect 1841 2433 3599 2434
rect 3605 2433 3606 2439
rect 84 2373 85 2379
rect 91 2378 1835 2379
rect 91 2374 111 2378
rect 115 2374 159 2378
rect 163 2374 183 2378
rect 187 2374 247 2378
rect 251 2374 311 2378
rect 315 2374 335 2378
rect 339 2374 439 2378
rect 443 2374 447 2378
rect 451 2374 559 2378
rect 563 2374 583 2378
rect 587 2374 687 2378
rect 691 2374 719 2378
rect 723 2374 815 2378
rect 819 2374 855 2378
rect 859 2374 951 2378
rect 955 2374 991 2378
rect 995 2374 1079 2378
rect 1083 2374 1127 2378
rect 1131 2374 1207 2378
rect 1211 2374 1263 2378
rect 1267 2374 1327 2378
rect 1331 2374 1399 2378
rect 1403 2374 1455 2378
rect 1459 2374 1583 2378
rect 1587 2374 1823 2378
rect 1827 2374 1835 2378
rect 91 2373 1835 2374
rect 1841 2373 1842 2379
rect 1846 2361 1847 2367
rect 1853 2366 3611 2367
rect 1853 2362 1863 2366
rect 1867 2362 1895 2366
rect 1899 2362 1927 2366
rect 1931 2362 2023 2366
rect 2027 2362 2087 2366
rect 2091 2362 2183 2366
rect 2187 2362 2247 2366
rect 2251 2362 2343 2366
rect 2347 2362 2407 2366
rect 2411 2362 2503 2366
rect 2507 2362 2559 2366
rect 2563 2362 2655 2366
rect 2659 2362 2703 2366
rect 2707 2362 2807 2366
rect 2811 2362 2831 2366
rect 2835 2362 2951 2366
rect 2955 2362 2959 2366
rect 2963 2362 3071 2366
rect 3075 2362 3119 2366
rect 3123 2362 3183 2366
rect 3187 2362 3287 2366
rect 3291 2362 3399 2366
rect 3403 2362 3487 2366
rect 3491 2362 3575 2366
rect 3579 2362 3611 2366
rect 1853 2361 3611 2362
rect 3617 2361 3618 2367
rect 1834 2307 1835 2313
rect 1841 2307 1866 2313
rect 96 2297 97 2303
rect 103 2302 1847 2303
rect 103 2298 111 2302
rect 115 2298 167 2302
rect 171 2298 255 2302
rect 259 2298 343 2302
rect 347 2298 447 2302
rect 451 2298 567 2302
rect 571 2298 695 2302
rect 699 2298 823 2302
rect 827 2298 863 2302
rect 867 2298 959 2302
rect 963 2298 1023 2302
rect 1027 2298 1087 2302
rect 1091 2298 1175 2302
rect 1179 2298 1215 2302
rect 1219 2298 1319 2302
rect 1323 2298 1335 2302
rect 1339 2298 1463 2302
rect 1467 2298 1591 2302
rect 1595 2298 1599 2302
rect 1603 2298 1735 2302
rect 1739 2298 1823 2302
rect 1827 2298 1847 2302
rect 103 2297 1847 2298
rect 1853 2297 1854 2303
rect 1860 2295 1866 2307
rect 1860 2294 3599 2295
rect 1860 2290 1863 2294
rect 1867 2290 1919 2294
rect 1923 2290 1975 2294
rect 1979 2290 2079 2294
rect 2083 2290 2143 2294
rect 2147 2290 2239 2294
rect 2243 2290 2311 2294
rect 2315 2290 2399 2294
rect 2403 2290 2479 2294
rect 2483 2290 2551 2294
rect 2555 2290 2639 2294
rect 2643 2290 2695 2294
rect 2699 2290 2783 2294
rect 2787 2290 2823 2294
rect 2827 2290 2919 2294
rect 2923 2290 2943 2294
rect 2947 2290 3039 2294
rect 3043 2290 3063 2294
rect 3067 2290 3159 2294
rect 3163 2290 3175 2294
rect 3179 2290 3271 2294
rect 3275 2290 3279 2294
rect 3283 2290 3383 2294
rect 3387 2290 3391 2294
rect 3395 2290 3479 2294
rect 3483 2290 3575 2294
rect 3579 2290 3599 2294
rect 1860 2289 3599 2290
rect 3605 2289 3606 2295
rect 84 2221 85 2227
rect 91 2226 1835 2227
rect 91 2222 111 2226
rect 115 2222 535 2226
rect 539 2222 687 2226
rect 691 2222 719 2226
rect 723 2222 855 2226
rect 859 2222 895 2226
rect 899 2222 1015 2226
rect 1019 2222 1071 2226
rect 1075 2222 1167 2226
rect 1171 2222 1239 2226
rect 1243 2222 1311 2226
rect 1315 2222 1407 2226
rect 1411 2222 1455 2226
rect 1459 2222 1575 2226
rect 1579 2222 1591 2226
rect 1595 2222 1727 2226
rect 1731 2222 1823 2226
rect 1827 2222 1835 2226
rect 91 2221 1835 2222
rect 1841 2221 1842 2227
rect 1846 2221 1847 2227
rect 1853 2226 3611 2227
rect 1853 2222 1863 2226
rect 1867 2222 1983 2226
rect 1987 2222 2007 2226
rect 2011 2222 2151 2226
rect 2155 2222 2167 2226
rect 2171 2222 2319 2226
rect 2323 2222 2335 2226
rect 2339 2222 2487 2226
rect 2491 2222 2519 2226
rect 2523 2222 2647 2226
rect 2651 2222 2711 2226
rect 2715 2222 2791 2226
rect 2795 2222 2903 2226
rect 2907 2222 2927 2226
rect 2931 2222 3047 2226
rect 3051 2222 3103 2226
rect 3107 2222 3167 2226
rect 3171 2222 3279 2226
rect 3283 2222 3303 2226
rect 3307 2222 3391 2226
rect 3395 2222 3487 2226
rect 3491 2222 3575 2226
rect 3579 2222 3611 2226
rect 1853 2221 3611 2222
rect 3617 2221 3618 2227
rect 1834 2163 1835 2169
rect 1841 2163 1866 2169
rect 96 2153 97 2159
rect 103 2158 1847 2159
rect 103 2154 111 2158
rect 115 2154 495 2158
rect 499 2154 543 2158
rect 547 2154 623 2158
rect 627 2154 727 2158
rect 731 2154 759 2158
rect 763 2154 895 2158
rect 899 2154 903 2158
rect 907 2154 1039 2158
rect 1043 2154 1079 2158
rect 1083 2154 1183 2158
rect 1187 2154 1247 2158
rect 1251 2154 1327 2158
rect 1331 2154 1415 2158
rect 1419 2154 1471 2158
rect 1475 2154 1583 2158
rect 1587 2154 1623 2158
rect 1627 2154 1735 2158
rect 1739 2154 1823 2158
rect 1827 2154 1847 2158
rect 103 2153 1847 2154
rect 1853 2153 1854 2159
rect 1860 2151 1866 2163
rect 1860 2150 3599 2151
rect 1860 2146 1863 2150
rect 1867 2146 1999 2150
rect 2003 2146 2023 2150
rect 2027 2146 2159 2150
rect 2163 2146 2167 2150
rect 2171 2146 2319 2150
rect 2323 2146 2327 2150
rect 2331 2146 2471 2150
rect 2475 2146 2511 2150
rect 2515 2146 2615 2150
rect 2619 2146 2703 2150
rect 2707 2146 2759 2150
rect 2763 2146 2895 2150
rect 2899 2146 3023 2150
rect 3027 2146 3095 2150
rect 3099 2146 3143 2150
rect 3147 2146 3263 2150
rect 3267 2146 3295 2150
rect 3299 2146 3383 2150
rect 3387 2146 3479 2150
rect 3483 2146 3575 2150
rect 3579 2146 3599 2150
rect 1860 2145 3599 2146
rect 3605 2145 3606 2151
rect 84 2081 85 2087
rect 91 2086 1835 2087
rect 91 2082 111 2086
rect 115 2082 319 2086
rect 323 2082 431 2086
rect 435 2082 487 2086
rect 491 2082 551 2086
rect 555 2082 615 2086
rect 619 2082 679 2086
rect 683 2082 751 2086
rect 755 2082 799 2086
rect 803 2082 887 2086
rect 891 2082 919 2086
rect 923 2082 1031 2086
rect 1035 2082 1039 2086
rect 1043 2082 1159 2086
rect 1163 2082 1175 2086
rect 1179 2082 1279 2086
rect 1283 2082 1319 2086
rect 1323 2082 1407 2086
rect 1411 2082 1463 2086
rect 1467 2082 1615 2086
rect 1619 2082 1823 2086
rect 1827 2082 1835 2086
rect 91 2081 1835 2082
rect 1841 2081 1842 2087
rect 1846 2073 1847 2079
rect 1853 2078 3611 2079
rect 1853 2074 1863 2078
rect 1867 2074 1983 2078
rect 1987 2074 2031 2078
rect 2035 2074 2143 2078
rect 2147 2074 2175 2078
rect 2179 2074 2311 2078
rect 2315 2074 2327 2078
rect 2331 2074 2471 2078
rect 2475 2074 2479 2078
rect 2483 2074 2623 2078
rect 2627 2074 2631 2078
rect 2635 2074 2767 2078
rect 2771 2074 2775 2078
rect 2779 2074 2903 2078
rect 2907 2074 2911 2078
rect 2915 2074 3031 2078
rect 3035 2074 3039 2078
rect 3043 2074 3151 2078
rect 3155 2074 3159 2078
rect 3163 2074 3271 2078
rect 3275 2074 3279 2078
rect 3283 2074 3391 2078
rect 3395 2074 3487 2078
rect 3491 2074 3575 2078
rect 3579 2074 3611 2078
rect 1853 2073 3611 2074
rect 3617 2073 3618 2079
rect 1834 2019 1835 2025
rect 1841 2019 1866 2025
rect 96 2009 97 2015
rect 103 2014 1847 2015
rect 103 2010 111 2014
rect 115 2010 183 2014
rect 187 2010 295 2014
rect 299 2010 327 2014
rect 331 2010 415 2014
rect 419 2010 439 2014
rect 443 2010 535 2014
rect 539 2010 559 2014
rect 563 2010 655 2014
rect 659 2010 687 2014
rect 691 2010 775 2014
rect 779 2010 807 2014
rect 811 2010 895 2014
rect 899 2010 927 2014
rect 931 2010 1015 2014
rect 1019 2010 1047 2014
rect 1051 2010 1135 2014
rect 1139 2010 1167 2014
rect 1171 2010 1255 2014
rect 1259 2010 1287 2014
rect 1291 2010 1415 2014
rect 1419 2010 1823 2014
rect 1827 2010 1847 2014
rect 103 2009 1847 2010
rect 1853 2009 1854 2015
rect 1860 2011 1866 2019
rect 1860 2010 3599 2011
rect 1860 2006 1863 2010
rect 1867 2006 1887 2010
rect 1891 2006 1975 2010
rect 1979 2006 2031 2010
rect 2035 2006 2135 2010
rect 2139 2006 2199 2010
rect 2203 2006 2303 2010
rect 2307 2006 2375 2010
rect 2379 2006 2463 2010
rect 2467 2006 2543 2010
rect 2547 2006 2623 2010
rect 2627 2006 2711 2010
rect 2715 2006 2767 2010
rect 2771 2006 2871 2010
rect 2875 2006 2903 2010
rect 2907 2006 3031 2010
rect 3035 2006 3039 2010
rect 3043 2006 3151 2010
rect 3155 2006 3207 2010
rect 3211 2006 3271 2010
rect 3275 2006 3383 2010
rect 3387 2006 3479 2010
rect 3483 2006 3575 2010
rect 3579 2006 3599 2010
rect 1860 2005 3599 2006
rect 3605 2005 3606 2011
rect 84 1937 85 1943
rect 91 1942 1835 1943
rect 91 1938 111 1942
rect 115 1938 135 1942
rect 139 1938 175 1942
rect 179 1938 223 1942
rect 227 1938 287 1942
rect 291 1938 351 1942
rect 355 1938 407 1942
rect 411 1938 495 1942
rect 499 1938 527 1942
rect 531 1938 647 1942
rect 651 1938 655 1942
rect 659 1938 767 1942
rect 771 1938 839 1942
rect 843 1938 887 1942
rect 891 1938 1007 1942
rect 1011 1938 1039 1942
rect 1043 1938 1127 1942
rect 1131 1938 1247 1942
rect 1251 1938 1463 1942
rect 1467 1938 1823 1942
rect 1827 1938 1835 1942
rect 91 1937 1835 1938
rect 1841 1937 1842 1943
rect 1846 1929 1847 1935
rect 1853 1934 3611 1935
rect 1853 1930 1863 1934
rect 1867 1930 1895 1934
rect 1899 1930 1991 1934
rect 1995 1930 2039 1934
rect 2043 1930 2119 1934
rect 2123 1930 2207 1934
rect 2211 1930 2255 1934
rect 2259 1930 2383 1934
rect 2387 1930 2511 1934
rect 2515 1930 2551 1934
rect 2555 1930 2631 1934
rect 2635 1930 2719 1934
rect 2723 1930 2751 1934
rect 2755 1930 2879 1934
rect 2883 1930 3007 1934
rect 3011 1930 3047 1934
rect 3051 1930 3215 1934
rect 3219 1930 3575 1934
rect 3579 1930 3611 1934
rect 1853 1929 3611 1930
rect 3617 1929 3618 1935
rect 1834 1871 1835 1877
rect 1841 1871 1866 1877
rect 96 1861 97 1867
rect 103 1866 1847 1867
rect 103 1862 111 1866
rect 115 1862 143 1866
rect 147 1862 231 1866
rect 235 1862 271 1866
rect 275 1862 359 1866
rect 363 1862 415 1866
rect 419 1862 503 1866
rect 507 1862 559 1866
rect 563 1862 663 1866
rect 667 1862 695 1866
rect 699 1862 823 1866
rect 827 1862 847 1866
rect 851 1862 943 1866
rect 947 1862 1047 1866
rect 1051 1862 1055 1866
rect 1059 1862 1159 1866
rect 1163 1862 1255 1866
rect 1259 1862 1263 1866
rect 1267 1862 1359 1866
rect 1363 1862 1455 1866
rect 1459 1862 1471 1866
rect 1475 1862 1551 1866
rect 1555 1862 1647 1866
rect 1651 1862 1735 1866
rect 1739 1862 1823 1866
rect 1827 1862 1847 1866
rect 103 1861 1847 1862
rect 1853 1861 1854 1867
rect 1860 1859 1866 1871
rect 1860 1858 3599 1859
rect 1860 1854 1863 1858
rect 1867 1854 1887 1858
rect 1891 1854 1983 1858
rect 1987 1854 2111 1858
rect 2115 1854 2223 1858
rect 2227 1854 2247 1858
rect 2251 1854 2359 1858
rect 2363 1854 2375 1858
rect 2379 1854 2495 1858
rect 2499 1854 2503 1858
rect 2507 1854 2623 1858
rect 2627 1854 2743 1858
rect 2747 1854 2863 1858
rect 2867 1854 2871 1858
rect 2875 1854 2991 1858
rect 2995 1854 2999 1858
rect 3003 1854 3575 1858
rect 3579 1854 3599 1858
rect 1860 1853 3599 1854
rect 3605 1853 3606 1859
rect 84 1781 85 1787
rect 91 1786 1835 1787
rect 91 1782 111 1786
rect 115 1782 135 1786
rect 139 1782 263 1786
rect 267 1782 303 1786
rect 307 1782 407 1786
rect 411 1782 495 1786
rect 499 1782 551 1786
rect 555 1782 687 1786
rect 691 1782 815 1786
rect 819 1782 871 1786
rect 875 1782 935 1786
rect 939 1782 1047 1786
rect 1051 1782 1151 1786
rect 1155 1782 1215 1786
rect 1219 1782 1255 1786
rect 1259 1782 1351 1786
rect 1355 1782 1375 1786
rect 1379 1782 1447 1786
rect 1451 1782 1535 1786
rect 1539 1782 1543 1786
rect 1547 1782 1639 1786
rect 1643 1782 1703 1786
rect 1707 1782 1727 1786
rect 1731 1782 1823 1786
rect 1827 1782 1835 1786
rect 91 1781 1835 1782
rect 1841 1781 1842 1787
rect 1846 1781 1847 1787
rect 1853 1786 3611 1787
rect 1853 1782 1863 1786
rect 1867 1782 2231 1786
rect 2235 1782 2271 1786
rect 2275 1782 2359 1786
rect 2363 1782 2367 1786
rect 2371 1782 2455 1786
rect 2459 1782 2503 1786
rect 2507 1782 2559 1786
rect 2563 1782 2631 1786
rect 2635 1782 2663 1786
rect 2667 1782 2751 1786
rect 2755 1782 2759 1786
rect 2763 1782 2863 1786
rect 2867 1782 2871 1786
rect 2875 1782 2967 1786
rect 2971 1782 2999 1786
rect 3003 1782 3071 1786
rect 3075 1782 3175 1786
rect 3179 1782 3575 1786
rect 3579 1782 3611 1786
rect 1853 1781 3611 1782
rect 3617 1781 3618 1787
rect 1834 1719 1835 1725
rect 1841 1719 1866 1725
rect 1860 1715 1866 1719
rect 96 1709 97 1715
rect 103 1714 1847 1715
rect 103 1710 111 1714
rect 115 1710 143 1714
rect 147 1710 287 1714
rect 291 1710 311 1714
rect 315 1710 471 1714
rect 475 1710 503 1714
rect 507 1710 655 1714
rect 659 1710 695 1714
rect 699 1710 839 1714
rect 843 1710 879 1714
rect 883 1710 1023 1714
rect 1027 1710 1055 1714
rect 1059 1710 1191 1714
rect 1195 1710 1223 1714
rect 1227 1710 1359 1714
rect 1363 1710 1383 1714
rect 1387 1710 1527 1714
rect 1531 1710 1543 1714
rect 1547 1710 1695 1714
rect 1699 1710 1711 1714
rect 1715 1710 1823 1714
rect 1827 1710 1847 1714
rect 103 1709 1847 1710
rect 1853 1709 1854 1715
rect 1860 1714 3599 1715
rect 1860 1710 1863 1714
rect 1867 1710 2247 1714
rect 2251 1710 2263 1714
rect 2267 1710 2351 1714
rect 2355 1710 2367 1714
rect 2371 1710 2447 1714
rect 2451 1710 2495 1714
rect 2499 1710 2551 1714
rect 2555 1710 2623 1714
rect 2627 1710 2655 1714
rect 2659 1710 2751 1714
rect 2755 1710 2759 1714
rect 2763 1710 2855 1714
rect 2859 1710 2887 1714
rect 2891 1710 2959 1714
rect 2963 1710 3015 1714
rect 3019 1710 3063 1714
rect 3067 1710 3135 1714
rect 3139 1710 3167 1714
rect 3171 1710 3247 1714
rect 3251 1710 3367 1714
rect 3371 1710 3479 1714
rect 3483 1710 3575 1714
rect 3579 1710 3599 1714
rect 1860 1709 3599 1710
rect 3605 1709 3606 1715
rect 84 1633 85 1639
rect 91 1638 1835 1639
rect 91 1634 111 1638
rect 115 1634 135 1638
rect 139 1634 271 1638
rect 275 1634 279 1638
rect 283 1634 447 1638
rect 451 1634 463 1638
rect 467 1634 631 1638
rect 635 1634 647 1638
rect 651 1634 815 1638
rect 819 1634 831 1638
rect 835 1634 991 1638
rect 995 1634 1015 1638
rect 1019 1634 1151 1638
rect 1155 1634 1183 1638
rect 1187 1634 1303 1638
rect 1307 1634 1351 1638
rect 1355 1634 1455 1638
rect 1459 1634 1519 1638
rect 1523 1634 1599 1638
rect 1603 1634 1687 1638
rect 1691 1634 1727 1638
rect 1731 1634 1823 1638
rect 1827 1634 1835 1638
rect 91 1633 1835 1634
rect 1841 1633 1842 1639
rect 1846 1637 1847 1643
rect 1853 1642 3611 1643
rect 1853 1638 1863 1642
rect 1867 1638 2151 1642
rect 2155 1638 2255 1642
rect 2259 1638 2343 1642
rect 2347 1638 2375 1642
rect 2379 1638 2503 1642
rect 2507 1638 2527 1642
rect 2531 1638 2631 1642
rect 2635 1638 2703 1642
rect 2707 1638 2767 1642
rect 2771 1638 2871 1642
rect 2875 1638 2895 1642
rect 2899 1638 3023 1642
rect 3027 1638 3031 1642
rect 3035 1638 3143 1642
rect 3147 1638 3191 1642
rect 3195 1638 3255 1642
rect 3259 1638 3351 1642
rect 3355 1638 3375 1642
rect 3379 1638 3487 1642
rect 3491 1638 3575 1642
rect 3579 1638 3611 1642
rect 1853 1637 3611 1638
rect 3617 1637 3618 1643
rect 1834 1575 1835 1581
rect 1841 1575 1866 1581
rect 1860 1574 3599 1575
rect 96 1565 97 1571
rect 103 1570 1847 1571
rect 103 1566 111 1570
rect 115 1566 143 1570
rect 147 1566 271 1570
rect 275 1566 279 1570
rect 283 1566 431 1570
rect 435 1566 455 1570
rect 459 1566 599 1570
rect 603 1566 639 1570
rect 643 1566 767 1570
rect 771 1566 823 1570
rect 827 1566 935 1570
rect 939 1566 999 1570
rect 1003 1566 1103 1570
rect 1107 1566 1159 1570
rect 1163 1566 1263 1570
rect 1267 1566 1311 1570
rect 1315 1566 1423 1570
rect 1427 1566 1463 1570
rect 1467 1566 1591 1570
rect 1595 1566 1607 1570
rect 1611 1566 1735 1570
rect 1739 1566 1823 1570
rect 1827 1566 1847 1570
rect 103 1565 1847 1566
rect 1853 1565 1854 1571
rect 1860 1570 1863 1574
rect 1867 1570 2087 1574
rect 2091 1570 2143 1574
rect 2147 1570 2279 1574
rect 2283 1570 2335 1574
rect 2339 1570 2455 1574
rect 2459 1570 2519 1574
rect 2523 1570 2623 1574
rect 2627 1570 2695 1574
rect 2699 1570 2791 1574
rect 2795 1570 2863 1574
rect 2867 1570 2951 1574
rect 2955 1570 3023 1574
rect 3027 1570 3111 1574
rect 3115 1570 3183 1574
rect 3187 1570 3271 1574
rect 3275 1570 3343 1574
rect 3347 1570 3431 1574
rect 3435 1570 3479 1574
rect 3483 1570 3575 1574
rect 3579 1570 3599 1574
rect 1860 1569 3599 1570
rect 3605 1569 3606 1575
rect 84 1493 85 1499
rect 91 1498 1835 1499
rect 91 1494 111 1498
rect 115 1494 135 1498
rect 139 1494 183 1498
rect 187 1494 263 1498
rect 267 1494 327 1498
rect 331 1494 423 1498
rect 427 1494 471 1498
rect 475 1494 591 1498
rect 595 1494 607 1498
rect 611 1494 743 1498
rect 747 1494 759 1498
rect 763 1494 871 1498
rect 875 1494 927 1498
rect 931 1494 991 1498
rect 995 1494 1095 1498
rect 1099 1494 1119 1498
rect 1123 1494 1247 1498
rect 1251 1494 1255 1498
rect 1259 1494 1375 1498
rect 1379 1494 1415 1498
rect 1419 1494 1583 1498
rect 1587 1494 1727 1498
rect 1731 1494 1823 1498
rect 1827 1494 1835 1498
rect 91 1493 1835 1494
rect 1841 1493 1842 1499
rect 1846 1493 1847 1499
rect 1853 1498 3611 1499
rect 1853 1494 1863 1498
rect 1867 1494 1895 1498
rect 1899 1494 1991 1498
rect 1995 1494 2095 1498
rect 2099 1494 2119 1498
rect 2123 1494 2247 1498
rect 2251 1494 2287 1498
rect 2291 1494 2383 1498
rect 2387 1494 2463 1498
rect 2467 1494 2535 1498
rect 2539 1494 2631 1498
rect 2635 1494 2703 1498
rect 2707 1494 2799 1498
rect 2803 1494 2887 1498
rect 2891 1494 2959 1498
rect 2963 1494 3087 1498
rect 3091 1494 3119 1498
rect 3123 1494 3279 1498
rect 3283 1494 3295 1498
rect 3299 1494 3439 1498
rect 3443 1494 3487 1498
rect 3491 1494 3575 1498
rect 3579 1494 3611 1498
rect 1853 1493 3611 1494
rect 3617 1493 3618 1499
rect 1834 1427 1835 1433
rect 1841 1427 1866 1433
rect 1860 1426 3599 1427
rect 96 1417 97 1423
rect 103 1422 1847 1423
rect 103 1418 111 1422
rect 115 1418 191 1422
rect 195 1418 199 1422
rect 203 1418 335 1422
rect 339 1418 463 1422
rect 467 1418 479 1422
rect 483 1418 583 1422
rect 587 1418 615 1422
rect 619 1418 703 1422
rect 707 1418 751 1422
rect 755 1418 815 1422
rect 819 1418 879 1422
rect 883 1418 919 1422
rect 923 1418 999 1422
rect 1003 1418 1015 1422
rect 1019 1418 1119 1422
rect 1123 1418 1127 1422
rect 1131 1418 1223 1422
rect 1227 1418 1255 1422
rect 1259 1418 1327 1422
rect 1331 1418 1383 1422
rect 1387 1418 1823 1422
rect 1827 1418 1847 1422
rect 103 1417 1847 1418
rect 1853 1417 1854 1423
rect 1860 1422 1863 1426
rect 1867 1422 1887 1426
rect 1891 1422 1975 1426
rect 1979 1422 1983 1426
rect 1987 1422 2071 1426
rect 2075 1422 2111 1426
rect 2115 1422 2183 1426
rect 2187 1422 2239 1426
rect 2243 1422 2303 1426
rect 2307 1422 2375 1426
rect 2379 1422 2439 1426
rect 2443 1422 2527 1426
rect 2531 1422 2607 1426
rect 2611 1422 2695 1426
rect 2699 1422 2807 1426
rect 2811 1422 2879 1426
rect 2883 1422 3031 1426
rect 3035 1422 3079 1426
rect 3083 1422 3263 1426
rect 3267 1422 3287 1426
rect 3291 1422 3479 1426
rect 3483 1422 3575 1426
rect 3579 1422 3599 1426
rect 1860 1421 3599 1422
rect 3605 1421 3606 1427
rect 84 1345 85 1351
rect 91 1350 1835 1351
rect 91 1346 111 1350
rect 115 1346 191 1350
rect 195 1346 231 1350
rect 235 1346 327 1350
rect 331 1346 383 1350
rect 387 1346 455 1350
rect 459 1346 543 1350
rect 547 1346 575 1350
rect 579 1346 695 1350
rect 699 1346 703 1350
rect 707 1346 807 1350
rect 811 1346 871 1350
rect 875 1346 911 1350
rect 915 1346 1007 1350
rect 1011 1346 1039 1350
rect 1043 1346 1111 1350
rect 1115 1346 1207 1350
rect 1211 1346 1215 1350
rect 1219 1346 1319 1350
rect 1323 1346 1375 1350
rect 1379 1346 1823 1350
rect 1827 1346 1835 1350
rect 91 1345 1835 1346
rect 1841 1345 1842 1351
rect 1846 1349 1847 1355
rect 1853 1354 3611 1355
rect 1853 1350 1863 1354
rect 1867 1350 1895 1354
rect 1899 1350 1983 1354
rect 1987 1350 2079 1354
rect 2083 1350 2103 1354
rect 2107 1350 2191 1354
rect 2195 1350 2223 1354
rect 2227 1350 2311 1354
rect 2315 1350 2359 1354
rect 2363 1350 2447 1354
rect 2451 1350 2511 1354
rect 2515 1350 2615 1354
rect 2619 1350 2687 1354
rect 2691 1350 2815 1354
rect 2819 1350 2871 1354
rect 2875 1350 3039 1354
rect 3043 1350 3071 1354
rect 3075 1350 3271 1354
rect 3275 1350 3279 1354
rect 3283 1350 3487 1354
rect 3491 1350 3575 1354
rect 3579 1350 3611 1354
rect 1853 1349 3611 1350
rect 3617 1349 3618 1355
rect 1834 1287 1835 1293
rect 1841 1287 1866 1293
rect 96 1277 97 1283
rect 103 1282 1847 1283
rect 103 1278 111 1282
rect 115 1278 215 1282
rect 219 1278 239 1282
rect 243 1278 359 1282
rect 363 1278 391 1282
rect 395 1278 519 1282
rect 523 1278 551 1282
rect 555 1278 679 1282
rect 683 1278 711 1282
rect 715 1278 839 1282
rect 843 1278 879 1282
rect 883 1278 999 1282
rect 1003 1278 1047 1282
rect 1051 1278 1151 1282
rect 1155 1278 1215 1282
rect 1219 1278 1295 1282
rect 1299 1278 1383 1282
rect 1387 1278 1439 1282
rect 1443 1278 1591 1282
rect 1595 1278 1823 1282
rect 1827 1278 1847 1282
rect 103 1277 1847 1278
rect 1853 1277 1854 1283
rect 1860 1275 1866 1287
rect 1860 1274 3599 1275
rect 1860 1270 1863 1274
rect 1867 1270 1887 1274
rect 1891 1270 1975 1274
rect 1979 1270 2055 1274
rect 2059 1270 2095 1274
rect 2099 1270 2143 1274
rect 2147 1270 2215 1274
rect 2219 1270 2239 1274
rect 2243 1270 2335 1274
rect 2339 1270 2351 1274
rect 2355 1270 2431 1274
rect 2435 1270 2503 1274
rect 2507 1270 2551 1274
rect 2555 1270 2679 1274
rect 2683 1270 2687 1274
rect 2691 1270 2855 1274
rect 2859 1270 2863 1274
rect 2867 1270 3039 1274
rect 3043 1270 3063 1274
rect 3067 1270 3231 1274
rect 3235 1270 3271 1274
rect 3275 1270 3431 1274
rect 3435 1270 3479 1274
rect 3483 1270 3575 1274
rect 3579 1270 3599 1274
rect 1860 1269 3599 1270
rect 3605 1269 3606 1275
rect 84 1201 85 1207
rect 91 1206 1835 1207
rect 91 1202 111 1206
rect 115 1202 135 1206
rect 139 1202 207 1206
rect 211 1202 271 1206
rect 275 1202 351 1206
rect 355 1202 423 1206
rect 427 1202 511 1206
rect 515 1202 575 1206
rect 579 1202 671 1206
rect 675 1202 727 1206
rect 731 1202 831 1206
rect 835 1202 887 1206
rect 891 1202 991 1206
rect 995 1202 1055 1206
rect 1059 1202 1143 1206
rect 1147 1202 1231 1206
rect 1235 1202 1287 1206
rect 1291 1202 1415 1206
rect 1419 1202 1431 1206
rect 1435 1202 1583 1206
rect 1587 1202 1599 1206
rect 1603 1202 1823 1206
rect 1827 1202 1835 1206
rect 91 1201 1835 1202
rect 1841 1201 1842 1207
rect 1846 1197 1847 1203
rect 1853 1202 3611 1203
rect 1853 1198 1863 1202
rect 1867 1198 2039 1202
rect 2043 1198 2063 1202
rect 2067 1198 2151 1202
rect 2155 1198 2247 1202
rect 2251 1198 2279 1202
rect 2283 1198 2343 1202
rect 2347 1198 2415 1202
rect 2419 1198 2439 1202
rect 2443 1198 2559 1202
rect 2563 1198 2695 1202
rect 2699 1198 2711 1202
rect 2715 1198 2863 1202
rect 2867 1198 3015 1202
rect 3019 1198 3047 1202
rect 3051 1198 3167 1202
rect 3171 1198 3239 1202
rect 3243 1198 3327 1202
rect 3331 1198 3439 1202
rect 3443 1198 3487 1202
rect 3491 1198 3575 1202
rect 3579 1198 3611 1202
rect 1853 1197 3611 1198
rect 3617 1197 3618 1203
rect 96 1133 97 1139
rect 103 1138 1847 1139
rect 103 1134 111 1138
rect 115 1134 143 1138
rect 147 1134 279 1138
rect 283 1134 295 1138
rect 299 1134 431 1138
rect 435 1134 479 1138
rect 483 1134 583 1138
rect 587 1134 663 1138
rect 667 1134 735 1138
rect 739 1134 847 1138
rect 851 1134 895 1138
rect 899 1134 1031 1138
rect 1035 1134 1063 1138
rect 1067 1134 1207 1138
rect 1211 1134 1239 1138
rect 1243 1134 1391 1138
rect 1395 1134 1423 1138
rect 1427 1134 1575 1138
rect 1579 1134 1607 1138
rect 1611 1134 1735 1138
rect 1739 1134 1823 1138
rect 1827 1134 1847 1138
rect 103 1133 1847 1134
rect 1853 1133 1854 1139
rect 1834 1117 1835 1123
rect 1841 1122 3599 1123
rect 1841 1118 1863 1122
rect 1867 1118 1943 1122
rect 1947 1118 2031 1122
rect 2035 1118 2087 1122
rect 2091 1118 2143 1122
rect 2147 1118 2231 1122
rect 2235 1118 2271 1122
rect 2275 1118 2383 1122
rect 2387 1118 2407 1122
rect 2411 1118 2535 1122
rect 2539 1118 2551 1122
rect 2555 1118 2687 1122
rect 2691 1118 2703 1122
rect 2707 1118 2839 1122
rect 2843 1118 2855 1122
rect 2859 1118 2991 1122
rect 2995 1118 3007 1122
rect 3011 1118 3151 1122
rect 3155 1118 3159 1122
rect 3163 1118 3319 1122
rect 3323 1118 3479 1122
rect 3483 1118 3575 1122
rect 3579 1118 3599 1122
rect 1841 1117 3599 1118
rect 3605 1117 3606 1123
rect 84 1065 85 1071
rect 91 1070 1835 1071
rect 91 1066 111 1070
rect 115 1066 135 1070
rect 139 1066 271 1070
rect 275 1066 287 1070
rect 291 1066 431 1070
rect 435 1066 471 1070
rect 475 1066 583 1070
rect 587 1066 655 1070
rect 659 1066 735 1070
rect 739 1066 839 1070
rect 843 1066 887 1070
rect 891 1066 1023 1070
rect 1027 1066 1047 1070
rect 1051 1066 1199 1070
rect 1203 1066 1215 1070
rect 1219 1066 1383 1070
rect 1387 1066 1559 1070
rect 1563 1066 1567 1070
rect 1571 1066 1727 1070
rect 1731 1066 1823 1070
rect 1827 1066 1835 1070
rect 91 1065 1835 1066
rect 1841 1065 1842 1071
rect 1846 1037 1847 1043
rect 1853 1042 3611 1043
rect 1853 1038 1863 1042
rect 1867 1038 1919 1042
rect 1923 1038 1951 1042
rect 1955 1038 2095 1042
rect 2099 1038 2127 1042
rect 2131 1038 2239 1042
rect 2243 1038 2327 1042
rect 2331 1038 2391 1042
rect 2395 1038 2519 1042
rect 2523 1038 2543 1042
rect 2547 1038 2695 1042
rect 2699 1038 2847 1042
rect 2851 1038 2863 1042
rect 2867 1038 2999 1042
rect 3003 1038 3023 1042
rect 3027 1038 3159 1042
rect 3163 1038 3183 1042
rect 3187 1038 3327 1042
rect 3331 1038 3343 1042
rect 3347 1038 3487 1042
rect 3491 1038 3575 1042
rect 3579 1038 3611 1042
rect 1853 1037 3611 1038
rect 3617 1037 3618 1043
rect 96 993 97 999
rect 103 998 1847 999
rect 103 994 111 998
rect 115 994 143 998
rect 147 994 279 998
rect 283 994 287 998
rect 291 994 439 998
rect 443 994 463 998
rect 467 994 591 998
rect 595 994 647 998
rect 651 994 743 998
rect 747 994 823 998
rect 827 994 895 998
rect 899 994 999 998
rect 1003 994 1055 998
rect 1059 994 1167 998
rect 1171 994 1223 998
rect 1227 994 1327 998
rect 1331 994 1391 998
rect 1395 994 1487 998
rect 1491 994 1567 998
rect 1571 994 1655 998
rect 1659 994 1735 998
rect 1739 994 1823 998
rect 1827 994 1847 998
rect 103 993 1847 994
rect 1853 993 1854 999
rect 1834 965 1835 971
rect 1841 970 3599 971
rect 1841 966 1863 970
rect 1867 966 1887 970
rect 1891 966 1911 970
rect 1915 966 2071 970
rect 2075 966 2119 970
rect 2123 966 2263 970
rect 2267 966 2319 970
rect 2323 966 2455 970
rect 2459 966 2511 970
rect 2515 966 2631 970
rect 2635 966 2687 970
rect 2691 966 2799 970
rect 2803 966 2855 970
rect 2859 966 2951 970
rect 2955 966 3015 970
rect 3019 966 3095 970
rect 3099 966 3175 970
rect 3179 966 3231 970
rect 3235 966 3335 970
rect 3339 966 3367 970
rect 3371 966 3479 970
rect 3483 966 3575 970
rect 3579 966 3599 970
rect 1841 965 3599 966
rect 3605 965 3606 971
rect 84 917 85 923
rect 91 922 1835 923
rect 91 918 111 922
rect 115 918 135 922
rect 139 918 271 922
rect 275 918 279 922
rect 283 918 439 922
rect 443 918 455 922
rect 459 918 607 922
rect 611 918 639 922
rect 643 918 775 922
rect 779 918 815 922
rect 819 918 935 922
rect 939 918 991 922
rect 995 918 1095 922
rect 1099 918 1159 922
rect 1163 918 1247 922
rect 1251 918 1319 922
rect 1323 918 1399 922
rect 1403 918 1479 922
rect 1483 918 1551 922
rect 1555 918 1647 922
rect 1651 918 1823 922
rect 1827 918 1835 922
rect 91 917 1835 918
rect 1841 917 1842 923
rect 1846 889 1847 895
rect 1853 894 3611 895
rect 1853 890 1863 894
rect 1867 890 1895 894
rect 1899 890 2023 894
rect 2027 890 2079 894
rect 2083 890 2183 894
rect 2187 890 2271 894
rect 2275 890 2351 894
rect 2355 890 2463 894
rect 2467 890 2519 894
rect 2523 890 2639 894
rect 2643 890 2687 894
rect 2691 890 2807 894
rect 2811 890 2839 894
rect 2843 890 2959 894
rect 2963 890 2983 894
rect 2987 890 3103 894
rect 3107 890 3119 894
rect 3123 890 3239 894
rect 3243 890 3247 894
rect 3251 890 3375 894
rect 3379 890 3487 894
rect 3491 890 3575 894
rect 3579 890 3611 894
rect 1853 889 3611 890
rect 3617 889 3618 895
rect 96 849 97 855
rect 103 854 1847 855
rect 103 850 111 854
rect 115 850 143 854
rect 147 850 279 854
rect 283 850 287 854
rect 291 850 447 854
rect 451 850 463 854
rect 467 850 615 854
rect 619 850 639 854
rect 643 850 783 854
rect 787 850 807 854
rect 811 850 943 854
rect 947 850 983 854
rect 987 850 1103 854
rect 1107 850 1159 854
rect 1163 850 1255 854
rect 1259 850 1335 854
rect 1339 850 1407 854
rect 1411 850 1511 854
rect 1515 850 1559 854
rect 1563 850 1823 854
rect 1827 850 1847 854
rect 103 849 1847 850
rect 1853 849 1854 855
rect 1834 813 1835 819
rect 1841 818 3599 819
rect 1841 814 1863 818
rect 1867 814 1887 818
rect 1891 814 2015 818
rect 2019 814 2071 818
rect 2075 814 2175 818
rect 2179 814 2263 818
rect 2267 814 2343 818
rect 2347 814 2447 818
rect 2451 814 2511 818
rect 2515 814 2623 818
rect 2627 814 2679 818
rect 2683 814 2791 818
rect 2795 814 2831 818
rect 2835 814 2943 818
rect 2947 814 2975 818
rect 2979 814 3087 818
rect 3091 814 3111 818
rect 3115 814 3223 818
rect 3227 814 3239 818
rect 3243 814 3359 818
rect 3363 814 3367 818
rect 3371 814 3479 818
rect 3483 814 3575 818
rect 3579 814 3599 818
rect 1841 813 3599 814
rect 3605 813 3606 819
rect 84 777 85 783
rect 91 782 1835 783
rect 91 778 111 782
rect 115 778 135 782
rect 139 778 271 782
rect 275 778 279 782
rect 283 778 439 782
rect 443 778 455 782
rect 459 778 607 782
rect 611 778 631 782
rect 635 778 775 782
rect 779 778 799 782
rect 803 778 935 782
rect 939 778 975 782
rect 979 778 1087 782
rect 1091 778 1151 782
rect 1155 778 1239 782
rect 1243 778 1327 782
rect 1331 778 1391 782
rect 1395 778 1503 782
rect 1507 778 1551 782
rect 1555 778 1823 782
rect 1827 778 1835 782
rect 91 777 1835 778
rect 1841 777 1842 783
rect 1846 745 1847 751
rect 1853 750 3611 751
rect 1853 746 1863 750
rect 1867 746 1895 750
rect 1899 746 2071 750
rect 2075 746 2079 750
rect 2083 746 2263 750
rect 2267 746 2271 750
rect 2275 746 2447 750
rect 2451 746 2455 750
rect 2459 746 2623 750
rect 2627 746 2631 750
rect 2635 746 2799 750
rect 2803 746 2951 750
rect 2955 746 2975 750
rect 2979 746 3095 750
rect 3099 746 3151 750
rect 3155 746 3231 750
rect 3235 746 3327 750
rect 3331 746 3367 750
rect 3371 746 3487 750
rect 3491 746 3575 750
rect 3579 746 3611 750
rect 1853 745 3611 746
rect 3617 745 3618 751
rect 96 705 97 711
rect 103 710 1847 711
rect 103 706 111 710
rect 115 706 143 710
rect 147 706 279 710
rect 283 706 287 710
rect 291 706 447 710
rect 451 706 455 710
rect 459 706 615 710
rect 619 706 623 710
rect 627 706 783 710
rect 787 706 791 710
rect 795 706 943 710
rect 947 706 959 710
rect 963 706 1095 710
rect 1099 706 1119 710
rect 1123 706 1247 710
rect 1251 706 1279 710
rect 1283 706 1399 710
rect 1403 706 1439 710
rect 1443 706 1559 710
rect 1563 706 1599 710
rect 1603 706 1823 710
rect 1827 706 1847 710
rect 103 705 1847 706
rect 1853 705 1854 711
rect 1834 673 1835 679
rect 1841 678 3599 679
rect 1841 674 1863 678
rect 1867 674 1887 678
rect 1891 674 1975 678
rect 1979 674 2063 678
rect 2067 674 2095 678
rect 2099 674 2223 678
rect 2227 674 2255 678
rect 2259 674 2351 678
rect 2355 674 2439 678
rect 2443 674 2479 678
rect 2483 674 2615 678
rect 2619 674 2767 678
rect 2771 674 2791 678
rect 2795 674 2935 678
rect 2939 674 2967 678
rect 2971 674 3119 678
rect 3123 674 3143 678
rect 3147 674 3311 678
rect 3315 674 3319 678
rect 3323 674 3479 678
rect 3483 674 3575 678
rect 3579 674 3599 678
rect 1841 673 3599 674
rect 3605 673 3606 679
rect 84 629 85 635
rect 91 634 1835 635
rect 91 630 111 634
rect 115 630 135 634
rect 139 630 279 634
rect 283 630 287 634
rect 291 630 447 634
rect 451 630 455 634
rect 459 630 615 634
rect 619 630 631 634
rect 635 630 783 634
rect 787 630 799 634
rect 803 630 951 634
rect 955 630 967 634
rect 971 630 1111 634
rect 1115 630 1119 634
rect 1123 630 1271 634
rect 1275 630 1415 634
rect 1419 630 1431 634
rect 1435 630 1559 634
rect 1563 630 1591 634
rect 1595 630 1711 634
rect 1715 630 1823 634
rect 1827 630 1835 634
rect 91 629 1835 630
rect 1841 629 1842 635
rect 1846 601 1847 607
rect 1853 606 3611 607
rect 1853 602 1863 606
rect 1867 602 1895 606
rect 1899 602 1983 606
rect 1987 602 2047 606
rect 2051 602 2103 606
rect 2107 602 2215 606
rect 2219 602 2231 606
rect 2235 602 2359 606
rect 2363 602 2391 606
rect 2395 602 2487 606
rect 2491 602 2583 606
rect 2587 602 2623 606
rect 2627 602 2775 606
rect 2779 602 2799 606
rect 2803 602 2943 606
rect 2947 602 3023 606
rect 3027 602 3127 606
rect 3131 602 3255 606
rect 3259 602 3319 606
rect 3323 602 3487 606
rect 3491 602 3575 606
rect 3579 602 3611 606
rect 1853 601 3611 602
rect 3617 601 3618 607
rect 96 557 97 563
rect 103 562 1847 563
rect 103 558 111 562
rect 115 558 143 562
rect 147 558 151 562
rect 155 558 295 562
rect 299 558 311 562
rect 315 558 463 562
rect 467 558 471 562
rect 475 558 631 562
rect 635 558 639 562
rect 643 558 783 562
rect 787 558 807 562
rect 811 558 927 562
rect 931 558 975 562
rect 979 558 1063 562
rect 1067 558 1127 562
rect 1131 558 1191 562
rect 1195 558 1279 562
rect 1283 558 1311 562
rect 1315 558 1423 562
rect 1427 558 1535 562
rect 1539 558 1567 562
rect 1571 558 1647 562
rect 1651 558 1719 562
rect 1723 558 1735 562
rect 1739 558 1823 562
rect 1827 558 1847 562
rect 103 557 1847 558
rect 1853 557 1854 563
rect 1834 525 1835 531
rect 1841 530 3599 531
rect 1841 526 1863 530
rect 1867 526 1887 530
rect 1891 526 2039 530
rect 2043 526 2191 530
rect 2195 526 2207 530
rect 2211 526 2279 530
rect 2283 526 2375 530
rect 2379 526 2383 530
rect 2387 526 2487 530
rect 2491 526 2575 530
rect 2579 526 2631 530
rect 2635 526 2791 530
rect 2795 526 2807 530
rect 2811 526 3007 530
rect 3011 526 3015 530
rect 3019 526 3215 530
rect 3219 526 3247 530
rect 3251 526 3431 530
rect 3435 526 3479 530
rect 3483 526 3575 530
rect 3579 526 3599 530
rect 1841 525 3599 526
rect 3605 525 3606 531
rect 84 481 85 487
rect 91 486 1835 487
rect 91 482 111 486
rect 115 482 143 486
rect 147 482 159 486
rect 163 482 303 486
rect 307 482 311 486
rect 315 482 463 486
rect 467 482 615 486
rect 619 482 623 486
rect 627 482 759 486
rect 763 482 775 486
rect 779 482 887 486
rect 891 482 919 486
rect 923 482 1007 486
rect 1011 482 1055 486
rect 1059 482 1127 486
rect 1131 482 1183 486
rect 1187 482 1239 486
rect 1243 482 1303 486
rect 1307 482 1343 486
rect 1347 482 1415 486
rect 1419 482 1439 486
rect 1443 482 1527 486
rect 1531 482 1543 486
rect 1547 482 1639 486
rect 1643 482 1727 486
rect 1731 482 1823 486
rect 1827 482 1835 486
rect 91 481 1835 482
rect 1841 481 1842 487
rect 1846 449 1847 455
rect 1853 454 3611 455
rect 1853 450 1863 454
rect 1867 450 1895 454
rect 1899 450 2039 454
rect 2043 450 2199 454
rect 2203 450 2207 454
rect 2211 450 2287 454
rect 2291 450 2383 454
rect 2387 450 2495 454
rect 2499 450 2575 454
rect 2579 450 2639 454
rect 2643 450 2783 454
rect 2787 450 2815 454
rect 2819 450 3007 454
rect 3011 450 3015 454
rect 3019 450 3223 454
rect 3227 450 3239 454
rect 3243 450 3439 454
rect 3443 450 3471 454
rect 3475 450 3575 454
rect 3579 450 3611 454
rect 1853 449 3611 450
rect 3617 449 3618 455
rect 96 413 97 419
rect 103 418 1847 419
rect 103 414 111 418
rect 115 414 151 418
rect 155 414 167 418
rect 171 414 271 418
rect 275 414 319 418
rect 323 414 407 418
rect 411 414 471 418
rect 475 414 551 418
rect 555 414 623 418
rect 627 414 711 418
rect 715 414 767 418
rect 771 414 887 418
rect 891 414 895 418
rect 899 414 1015 418
rect 1019 414 1063 418
rect 1067 414 1135 418
rect 1139 414 1247 418
rect 1251 414 1351 418
rect 1355 414 1439 418
rect 1443 414 1447 418
rect 1451 414 1551 418
rect 1555 414 1639 418
rect 1643 414 1647 418
rect 1651 414 1735 418
rect 1739 414 1823 418
rect 1827 414 1847 418
rect 103 413 1847 414
rect 1853 413 1854 419
rect 1834 381 1835 387
rect 1841 386 3599 387
rect 1841 382 1863 386
rect 1867 382 1887 386
rect 1891 382 1975 386
rect 1979 382 2031 386
rect 2035 382 2063 386
rect 2067 382 2151 386
rect 2155 382 2199 386
rect 2203 382 2263 386
rect 2267 382 2375 386
rect 2379 382 2383 386
rect 2387 382 2519 386
rect 2523 382 2567 386
rect 2571 382 2671 386
rect 2675 382 2775 386
rect 2779 382 2847 386
rect 2851 382 2999 386
rect 3003 382 3031 386
rect 3035 382 3231 386
rect 3235 382 3431 386
rect 3435 382 3463 386
rect 3467 382 3575 386
rect 3579 382 3599 386
rect 1841 381 3599 382
rect 3605 381 3606 387
rect 84 329 85 335
rect 91 334 1835 335
rect 91 330 111 334
rect 115 330 135 334
rect 139 330 143 334
rect 147 330 223 334
rect 227 330 263 334
rect 267 330 311 334
rect 315 330 399 334
rect 403 330 487 334
rect 491 330 543 334
rect 547 330 575 334
rect 579 330 663 334
rect 667 330 703 334
rect 707 330 751 334
rect 755 330 839 334
rect 843 330 879 334
rect 883 330 927 334
rect 931 330 1015 334
rect 1019 330 1055 334
rect 1059 330 1103 334
rect 1107 330 1191 334
rect 1195 330 1239 334
rect 1243 330 1287 334
rect 1291 330 1383 334
rect 1387 330 1431 334
rect 1435 330 1479 334
rect 1483 330 1575 334
rect 1579 330 1631 334
rect 1635 330 1671 334
rect 1675 330 1823 334
rect 1827 330 1835 334
rect 91 329 1835 330
rect 1841 329 1842 335
rect 1846 313 1847 319
rect 1853 318 3611 319
rect 1853 314 1863 318
rect 1867 314 1895 318
rect 1899 314 1983 318
rect 1987 314 2071 318
rect 2075 314 2159 318
rect 2163 314 2247 318
rect 2251 314 2271 318
rect 2275 314 2359 318
rect 2363 314 2391 318
rect 2395 314 2471 318
rect 2475 314 2527 318
rect 2531 314 2583 318
rect 2587 314 2679 318
rect 2683 314 2695 318
rect 2699 314 2807 318
rect 2811 314 2855 318
rect 2859 314 2919 318
rect 2923 314 3039 318
rect 3043 314 3159 318
rect 3163 314 3239 318
rect 3243 314 3439 318
rect 3443 314 3575 318
rect 3579 314 3611 318
rect 1853 313 3611 314
rect 3617 313 3618 319
rect 96 257 97 263
rect 103 262 1847 263
rect 103 258 111 262
rect 115 258 143 262
rect 147 258 231 262
rect 235 258 319 262
rect 323 258 407 262
rect 411 258 495 262
rect 499 258 583 262
rect 587 258 671 262
rect 675 258 759 262
rect 763 258 847 262
rect 851 258 935 262
rect 939 258 1023 262
rect 1027 258 1111 262
rect 1115 258 1199 262
rect 1203 258 1287 262
rect 1291 258 1295 262
rect 1299 258 1375 262
rect 1379 258 1391 262
rect 1395 258 1463 262
rect 1467 258 1487 262
rect 1491 258 1551 262
rect 1555 258 1583 262
rect 1587 258 1639 262
rect 1643 258 1679 262
rect 1683 258 1727 262
rect 1731 258 1823 262
rect 1827 258 1847 262
rect 103 257 1847 258
rect 1853 257 1854 263
rect 1834 245 1835 251
rect 1841 250 3599 251
rect 1841 246 1863 250
rect 1867 246 1887 250
rect 1891 246 1975 250
rect 1979 246 2063 250
rect 2067 246 2151 250
rect 2155 246 2239 250
rect 2243 246 2263 250
rect 2267 246 2351 250
rect 2355 246 2399 250
rect 2403 246 2463 250
rect 2467 246 2535 250
rect 2539 246 2575 250
rect 2579 246 2679 250
rect 2683 246 2687 250
rect 2691 246 2799 250
rect 2803 246 2815 250
rect 2819 246 2911 250
rect 2915 246 2951 250
rect 2955 246 3031 250
rect 3035 246 3087 250
rect 3091 246 3151 250
rect 3155 246 3223 250
rect 3227 246 3359 250
rect 3363 246 3479 250
rect 3483 246 3575 250
rect 3579 246 3599 250
rect 1841 245 3599 246
rect 3605 245 3606 251
rect 84 189 85 195
rect 91 194 1835 195
rect 91 190 111 194
rect 115 190 135 194
rect 139 190 223 194
rect 227 190 311 194
rect 315 190 399 194
rect 403 190 487 194
rect 491 190 575 194
rect 579 190 663 194
rect 667 190 751 194
rect 755 190 839 194
rect 843 190 927 194
rect 931 190 1015 194
rect 1019 190 1103 194
rect 1107 190 1191 194
rect 1195 190 1279 194
rect 1283 190 1367 194
rect 1371 190 1455 194
rect 1459 190 1543 194
rect 1547 190 1631 194
rect 1635 190 1719 194
rect 1723 190 1823 194
rect 1827 190 1835 194
rect 91 189 1835 190
rect 1841 189 1842 195
rect 1846 145 1847 151
rect 1853 150 3611 151
rect 1853 146 1863 150
rect 1867 146 1895 150
rect 1899 146 1983 150
rect 1987 146 2071 150
rect 2075 146 2159 150
rect 2163 146 2271 150
rect 2275 146 2407 150
rect 2411 146 2543 150
rect 2547 146 2687 150
rect 2691 146 2783 150
rect 2787 146 2823 150
rect 2827 146 2871 150
rect 2875 146 2959 150
rect 2963 146 3047 150
rect 3051 146 3095 150
rect 3099 146 3135 150
rect 3139 146 3223 150
rect 3227 146 3231 150
rect 3235 146 3311 150
rect 3315 146 3367 150
rect 3371 146 3399 150
rect 3403 146 3487 150
rect 3491 146 3575 150
rect 3579 146 3611 150
rect 1853 145 3611 146
rect 3617 145 3618 151
rect 1834 77 1835 83
rect 1841 82 3599 83
rect 1841 78 1863 82
rect 1867 78 2775 82
rect 2779 78 2863 82
rect 2867 78 2951 82
rect 2955 78 3039 82
rect 3043 78 3127 82
rect 3131 78 3215 82
rect 3219 78 3303 82
rect 3307 78 3391 82
rect 3395 78 3479 82
rect 3483 78 3575 82
rect 3579 78 3599 82
rect 1841 77 3599 78
rect 3605 77 3606 83
<< m5c >>
rect 85 3665 91 3671
rect 1835 3665 1841 3671
rect 1835 3607 1841 3613
rect 97 3597 103 3603
rect 1847 3597 1853 3603
rect 3599 3589 3605 3595
rect 85 3529 91 3535
rect 1835 3529 1841 3535
rect 1847 3521 1853 3527
rect 3611 3521 3617 3527
rect 97 3461 103 3467
rect 1847 3461 1853 3467
rect 1835 3445 1841 3451
rect 3599 3445 3605 3451
rect 85 3393 91 3399
rect 1835 3393 1841 3399
rect 1847 3369 1853 3375
rect 3611 3369 3617 3375
rect 97 3321 103 3327
rect 1847 3321 1853 3327
rect 1835 3301 1841 3307
rect 3599 3301 3605 3307
rect 85 3249 91 3255
rect 1835 3249 1841 3255
rect 1847 3225 1853 3231
rect 3611 3225 3617 3231
rect 97 3173 103 3179
rect 1847 3173 1853 3179
rect 1835 3153 1841 3159
rect 3599 3153 3605 3159
rect 85 3097 91 3103
rect 1835 3097 1841 3103
rect 1847 3077 1853 3083
rect 3611 3077 3617 3083
rect 97 3025 103 3031
rect 1847 3025 1853 3031
rect 1835 3005 1841 3011
rect 3599 3005 3605 3011
rect 85 2957 91 2963
rect 1835 2957 1841 2963
rect 1847 2929 1853 2935
rect 3611 2929 3617 2935
rect 97 2885 103 2891
rect 1847 2885 1853 2891
rect 1835 2861 1841 2867
rect 3599 2861 3605 2867
rect 85 2809 91 2815
rect 1835 2809 1841 2815
rect 1847 2793 1853 2799
rect 3611 2793 3617 2799
rect 97 2733 103 2739
rect 1847 2733 1853 2739
rect 1835 2721 1841 2727
rect 3599 2721 3605 2727
rect 85 2661 91 2667
rect 1835 2661 1841 2667
rect 1847 2645 1853 2651
rect 3611 2645 3617 2651
rect 97 2589 103 2595
rect 1847 2589 1853 2595
rect 1835 2573 1841 2579
rect 3599 2573 3605 2579
rect 85 2521 91 2527
rect 1835 2521 1841 2527
rect 1847 2501 1853 2507
rect 3611 2501 3617 2507
rect 97 2453 103 2459
rect 1847 2453 1853 2459
rect 1835 2433 1841 2439
rect 3599 2433 3605 2439
rect 85 2373 91 2379
rect 1835 2373 1841 2379
rect 1847 2361 1853 2367
rect 3611 2361 3617 2367
rect 1835 2307 1841 2313
rect 97 2297 103 2303
rect 1847 2297 1853 2303
rect 3599 2289 3605 2295
rect 85 2221 91 2227
rect 1835 2221 1841 2227
rect 1847 2221 1853 2227
rect 3611 2221 3617 2227
rect 1835 2163 1841 2169
rect 97 2153 103 2159
rect 1847 2153 1853 2159
rect 3599 2145 3605 2151
rect 85 2081 91 2087
rect 1835 2081 1841 2087
rect 1847 2073 1853 2079
rect 3611 2073 3617 2079
rect 1835 2019 1841 2025
rect 97 2009 103 2015
rect 1847 2009 1853 2015
rect 3599 2005 3605 2011
rect 85 1937 91 1943
rect 1835 1937 1841 1943
rect 1847 1929 1853 1935
rect 3611 1929 3617 1935
rect 1835 1871 1841 1877
rect 97 1861 103 1867
rect 1847 1861 1853 1867
rect 3599 1853 3605 1859
rect 85 1781 91 1787
rect 1835 1781 1841 1787
rect 1847 1781 1853 1787
rect 3611 1781 3617 1787
rect 1835 1719 1841 1725
rect 97 1709 103 1715
rect 1847 1709 1853 1715
rect 3599 1709 3605 1715
rect 85 1633 91 1639
rect 1835 1633 1841 1639
rect 1847 1637 1853 1643
rect 3611 1637 3617 1643
rect 1835 1575 1841 1581
rect 97 1565 103 1571
rect 1847 1565 1853 1571
rect 3599 1569 3605 1575
rect 85 1493 91 1499
rect 1835 1493 1841 1499
rect 1847 1493 1853 1499
rect 3611 1493 3617 1499
rect 1835 1427 1841 1433
rect 97 1417 103 1423
rect 1847 1417 1853 1423
rect 3599 1421 3605 1427
rect 85 1345 91 1351
rect 1835 1345 1841 1351
rect 1847 1349 1853 1355
rect 3611 1349 3617 1355
rect 1835 1287 1841 1293
rect 97 1277 103 1283
rect 1847 1277 1853 1283
rect 3599 1269 3605 1275
rect 85 1201 91 1207
rect 1835 1201 1841 1207
rect 1847 1197 1853 1203
rect 3611 1197 3617 1203
rect 97 1133 103 1139
rect 1847 1133 1853 1139
rect 1835 1117 1841 1123
rect 3599 1117 3605 1123
rect 85 1065 91 1071
rect 1835 1065 1841 1071
rect 1847 1037 1853 1043
rect 3611 1037 3617 1043
rect 97 993 103 999
rect 1847 993 1853 999
rect 1835 965 1841 971
rect 3599 965 3605 971
rect 85 917 91 923
rect 1835 917 1841 923
rect 1847 889 1853 895
rect 3611 889 3617 895
rect 97 849 103 855
rect 1847 849 1853 855
rect 1835 813 1841 819
rect 3599 813 3605 819
rect 85 777 91 783
rect 1835 777 1841 783
rect 1847 745 1853 751
rect 3611 745 3617 751
rect 97 705 103 711
rect 1847 705 1853 711
rect 1835 673 1841 679
rect 3599 673 3605 679
rect 85 629 91 635
rect 1835 629 1841 635
rect 1847 601 1853 607
rect 3611 601 3617 607
rect 97 557 103 563
rect 1847 557 1853 563
rect 1835 525 1841 531
rect 3599 525 3605 531
rect 85 481 91 487
rect 1835 481 1841 487
rect 1847 449 1853 455
rect 3611 449 3617 455
rect 97 413 103 419
rect 1847 413 1853 419
rect 1835 381 1841 387
rect 3599 381 3605 387
rect 85 329 91 335
rect 1835 329 1841 335
rect 1847 313 1853 319
rect 3611 313 3617 319
rect 97 257 103 263
rect 1847 257 1853 263
rect 1835 245 1841 251
rect 3599 245 3605 251
rect 85 189 91 195
rect 1835 189 1841 195
rect 1847 145 1853 151
rect 3611 145 3617 151
rect 1835 77 1841 83
rect 3599 77 3605 83
<< m5 >>
rect 84 3671 92 3672
rect 84 3665 85 3671
rect 91 3665 92 3671
rect 84 3535 92 3665
rect 84 3529 85 3535
rect 91 3529 92 3535
rect 84 3399 92 3529
rect 84 3393 85 3399
rect 91 3393 92 3399
rect 84 3255 92 3393
rect 84 3249 85 3255
rect 91 3249 92 3255
rect 84 3103 92 3249
rect 84 3097 85 3103
rect 91 3097 92 3103
rect 84 2963 92 3097
rect 84 2957 85 2963
rect 91 2957 92 2963
rect 84 2815 92 2957
rect 84 2809 85 2815
rect 91 2809 92 2815
rect 84 2667 92 2809
rect 84 2661 85 2667
rect 91 2661 92 2667
rect 84 2527 92 2661
rect 84 2521 85 2527
rect 91 2521 92 2527
rect 84 2379 92 2521
rect 84 2373 85 2379
rect 91 2373 92 2379
rect 84 2227 92 2373
rect 84 2221 85 2227
rect 91 2221 92 2227
rect 84 2087 92 2221
rect 84 2081 85 2087
rect 91 2081 92 2087
rect 84 1943 92 2081
rect 84 1937 85 1943
rect 91 1937 92 1943
rect 84 1787 92 1937
rect 84 1781 85 1787
rect 91 1781 92 1787
rect 84 1639 92 1781
rect 84 1633 85 1639
rect 91 1633 92 1639
rect 84 1499 92 1633
rect 84 1493 85 1499
rect 91 1493 92 1499
rect 84 1351 92 1493
rect 84 1345 85 1351
rect 91 1345 92 1351
rect 84 1207 92 1345
rect 84 1201 85 1207
rect 91 1201 92 1207
rect 84 1071 92 1201
rect 84 1065 85 1071
rect 91 1065 92 1071
rect 84 923 92 1065
rect 84 917 85 923
rect 91 917 92 923
rect 84 783 92 917
rect 84 777 85 783
rect 91 777 92 783
rect 84 635 92 777
rect 84 629 85 635
rect 91 629 92 635
rect 84 487 92 629
rect 84 481 85 487
rect 91 481 92 487
rect 84 335 92 481
rect 84 329 85 335
rect 91 329 92 335
rect 84 195 92 329
rect 84 189 85 195
rect 91 189 92 195
rect 84 72 92 189
rect 96 3603 104 3672
rect 96 3597 97 3603
rect 103 3597 104 3603
rect 96 3467 104 3597
rect 96 3461 97 3467
rect 103 3461 104 3467
rect 96 3327 104 3461
rect 96 3321 97 3327
rect 103 3321 104 3327
rect 96 3179 104 3321
rect 96 3173 97 3179
rect 103 3173 104 3179
rect 96 3031 104 3173
rect 96 3025 97 3031
rect 103 3025 104 3031
rect 96 2891 104 3025
rect 96 2885 97 2891
rect 103 2885 104 2891
rect 96 2739 104 2885
rect 96 2733 97 2739
rect 103 2733 104 2739
rect 96 2595 104 2733
rect 96 2589 97 2595
rect 103 2589 104 2595
rect 96 2459 104 2589
rect 96 2453 97 2459
rect 103 2453 104 2459
rect 96 2303 104 2453
rect 96 2297 97 2303
rect 103 2297 104 2303
rect 96 2159 104 2297
rect 96 2153 97 2159
rect 103 2153 104 2159
rect 96 2015 104 2153
rect 96 2009 97 2015
rect 103 2009 104 2015
rect 96 1867 104 2009
rect 96 1861 97 1867
rect 103 1861 104 1867
rect 96 1715 104 1861
rect 96 1709 97 1715
rect 103 1709 104 1715
rect 96 1571 104 1709
rect 96 1565 97 1571
rect 103 1565 104 1571
rect 96 1423 104 1565
rect 96 1417 97 1423
rect 103 1417 104 1423
rect 96 1283 104 1417
rect 96 1277 97 1283
rect 103 1277 104 1283
rect 96 1139 104 1277
rect 96 1133 97 1139
rect 103 1133 104 1139
rect 96 999 104 1133
rect 96 993 97 999
rect 103 993 104 999
rect 96 855 104 993
rect 96 849 97 855
rect 103 849 104 855
rect 96 711 104 849
rect 96 705 97 711
rect 103 705 104 711
rect 96 563 104 705
rect 96 557 97 563
rect 103 557 104 563
rect 96 419 104 557
rect 96 413 97 419
rect 103 413 104 419
rect 96 263 104 413
rect 96 257 97 263
rect 103 257 104 263
rect 96 72 104 257
rect 1834 3671 1842 3672
rect 1834 3665 1835 3671
rect 1841 3665 1842 3671
rect 1834 3613 1842 3665
rect 1834 3607 1835 3613
rect 1841 3607 1842 3613
rect 1834 3535 1842 3607
rect 1834 3529 1835 3535
rect 1841 3529 1842 3535
rect 1834 3451 1842 3529
rect 1834 3445 1835 3451
rect 1841 3445 1842 3451
rect 1834 3399 1842 3445
rect 1834 3393 1835 3399
rect 1841 3393 1842 3399
rect 1834 3307 1842 3393
rect 1834 3301 1835 3307
rect 1841 3301 1842 3307
rect 1834 3255 1842 3301
rect 1834 3249 1835 3255
rect 1841 3249 1842 3255
rect 1834 3159 1842 3249
rect 1834 3153 1835 3159
rect 1841 3153 1842 3159
rect 1834 3103 1842 3153
rect 1834 3097 1835 3103
rect 1841 3097 1842 3103
rect 1834 3011 1842 3097
rect 1834 3005 1835 3011
rect 1841 3005 1842 3011
rect 1834 2963 1842 3005
rect 1834 2957 1835 2963
rect 1841 2957 1842 2963
rect 1834 2867 1842 2957
rect 1834 2861 1835 2867
rect 1841 2861 1842 2867
rect 1834 2815 1842 2861
rect 1834 2809 1835 2815
rect 1841 2809 1842 2815
rect 1834 2727 1842 2809
rect 1834 2721 1835 2727
rect 1841 2721 1842 2727
rect 1834 2667 1842 2721
rect 1834 2661 1835 2667
rect 1841 2661 1842 2667
rect 1834 2579 1842 2661
rect 1834 2573 1835 2579
rect 1841 2573 1842 2579
rect 1834 2527 1842 2573
rect 1834 2521 1835 2527
rect 1841 2521 1842 2527
rect 1834 2439 1842 2521
rect 1834 2433 1835 2439
rect 1841 2433 1842 2439
rect 1834 2379 1842 2433
rect 1834 2373 1835 2379
rect 1841 2373 1842 2379
rect 1834 2313 1842 2373
rect 1834 2307 1835 2313
rect 1841 2307 1842 2313
rect 1834 2227 1842 2307
rect 1834 2221 1835 2227
rect 1841 2221 1842 2227
rect 1834 2169 1842 2221
rect 1834 2163 1835 2169
rect 1841 2163 1842 2169
rect 1834 2087 1842 2163
rect 1834 2081 1835 2087
rect 1841 2081 1842 2087
rect 1834 2025 1842 2081
rect 1834 2019 1835 2025
rect 1841 2019 1842 2025
rect 1834 1943 1842 2019
rect 1834 1937 1835 1943
rect 1841 1937 1842 1943
rect 1834 1877 1842 1937
rect 1834 1871 1835 1877
rect 1841 1871 1842 1877
rect 1834 1787 1842 1871
rect 1834 1781 1835 1787
rect 1841 1781 1842 1787
rect 1834 1725 1842 1781
rect 1834 1719 1835 1725
rect 1841 1719 1842 1725
rect 1834 1639 1842 1719
rect 1834 1633 1835 1639
rect 1841 1633 1842 1639
rect 1834 1581 1842 1633
rect 1834 1575 1835 1581
rect 1841 1575 1842 1581
rect 1834 1499 1842 1575
rect 1834 1493 1835 1499
rect 1841 1493 1842 1499
rect 1834 1433 1842 1493
rect 1834 1427 1835 1433
rect 1841 1427 1842 1433
rect 1834 1351 1842 1427
rect 1834 1345 1835 1351
rect 1841 1345 1842 1351
rect 1834 1293 1842 1345
rect 1834 1287 1835 1293
rect 1841 1287 1842 1293
rect 1834 1207 1842 1287
rect 1834 1201 1835 1207
rect 1841 1201 1842 1207
rect 1834 1123 1842 1201
rect 1834 1117 1835 1123
rect 1841 1117 1842 1123
rect 1834 1071 1842 1117
rect 1834 1065 1835 1071
rect 1841 1065 1842 1071
rect 1834 971 1842 1065
rect 1834 965 1835 971
rect 1841 965 1842 971
rect 1834 923 1842 965
rect 1834 917 1835 923
rect 1841 917 1842 923
rect 1834 819 1842 917
rect 1834 813 1835 819
rect 1841 813 1842 819
rect 1834 783 1842 813
rect 1834 777 1835 783
rect 1841 777 1842 783
rect 1834 679 1842 777
rect 1834 673 1835 679
rect 1841 673 1842 679
rect 1834 635 1842 673
rect 1834 629 1835 635
rect 1841 629 1842 635
rect 1834 531 1842 629
rect 1834 525 1835 531
rect 1841 525 1842 531
rect 1834 487 1842 525
rect 1834 481 1835 487
rect 1841 481 1842 487
rect 1834 387 1842 481
rect 1834 381 1835 387
rect 1841 381 1842 387
rect 1834 335 1842 381
rect 1834 329 1835 335
rect 1841 329 1842 335
rect 1834 251 1842 329
rect 1834 245 1835 251
rect 1841 245 1842 251
rect 1834 195 1842 245
rect 1834 189 1835 195
rect 1841 189 1842 195
rect 1834 83 1842 189
rect 1834 77 1835 83
rect 1841 77 1842 83
rect 1834 72 1842 77
rect 1846 3603 1854 3672
rect 1846 3597 1847 3603
rect 1853 3597 1854 3603
rect 1846 3527 1854 3597
rect 1846 3521 1847 3527
rect 1853 3521 1854 3527
rect 1846 3467 1854 3521
rect 1846 3461 1847 3467
rect 1853 3461 1854 3467
rect 1846 3375 1854 3461
rect 1846 3369 1847 3375
rect 1853 3369 1854 3375
rect 1846 3327 1854 3369
rect 1846 3321 1847 3327
rect 1853 3321 1854 3327
rect 1846 3231 1854 3321
rect 1846 3225 1847 3231
rect 1853 3225 1854 3231
rect 1846 3179 1854 3225
rect 1846 3173 1847 3179
rect 1853 3173 1854 3179
rect 1846 3083 1854 3173
rect 1846 3077 1847 3083
rect 1853 3077 1854 3083
rect 1846 3031 1854 3077
rect 1846 3025 1847 3031
rect 1853 3025 1854 3031
rect 1846 2935 1854 3025
rect 1846 2929 1847 2935
rect 1853 2929 1854 2935
rect 1846 2891 1854 2929
rect 1846 2885 1847 2891
rect 1853 2885 1854 2891
rect 1846 2799 1854 2885
rect 1846 2793 1847 2799
rect 1853 2793 1854 2799
rect 1846 2739 1854 2793
rect 1846 2733 1847 2739
rect 1853 2733 1854 2739
rect 1846 2651 1854 2733
rect 1846 2645 1847 2651
rect 1853 2645 1854 2651
rect 1846 2595 1854 2645
rect 1846 2589 1847 2595
rect 1853 2589 1854 2595
rect 1846 2507 1854 2589
rect 1846 2501 1847 2507
rect 1853 2501 1854 2507
rect 1846 2459 1854 2501
rect 1846 2453 1847 2459
rect 1853 2453 1854 2459
rect 1846 2367 1854 2453
rect 1846 2361 1847 2367
rect 1853 2361 1854 2367
rect 1846 2303 1854 2361
rect 1846 2297 1847 2303
rect 1853 2297 1854 2303
rect 1846 2227 1854 2297
rect 1846 2221 1847 2227
rect 1853 2221 1854 2227
rect 1846 2159 1854 2221
rect 1846 2153 1847 2159
rect 1853 2153 1854 2159
rect 1846 2079 1854 2153
rect 1846 2073 1847 2079
rect 1853 2073 1854 2079
rect 1846 2015 1854 2073
rect 1846 2009 1847 2015
rect 1853 2009 1854 2015
rect 1846 1935 1854 2009
rect 1846 1929 1847 1935
rect 1853 1929 1854 1935
rect 1846 1867 1854 1929
rect 1846 1861 1847 1867
rect 1853 1861 1854 1867
rect 1846 1787 1854 1861
rect 1846 1781 1847 1787
rect 1853 1781 1854 1787
rect 1846 1715 1854 1781
rect 1846 1709 1847 1715
rect 1853 1709 1854 1715
rect 1846 1643 1854 1709
rect 1846 1637 1847 1643
rect 1853 1637 1854 1643
rect 1846 1571 1854 1637
rect 1846 1565 1847 1571
rect 1853 1565 1854 1571
rect 1846 1499 1854 1565
rect 1846 1493 1847 1499
rect 1853 1493 1854 1499
rect 1846 1423 1854 1493
rect 1846 1417 1847 1423
rect 1853 1417 1854 1423
rect 1846 1355 1854 1417
rect 1846 1349 1847 1355
rect 1853 1349 1854 1355
rect 1846 1283 1854 1349
rect 1846 1277 1847 1283
rect 1853 1277 1854 1283
rect 1846 1203 1854 1277
rect 1846 1197 1847 1203
rect 1853 1197 1854 1203
rect 1846 1139 1854 1197
rect 1846 1133 1847 1139
rect 1853 1133 1854 1139
rect 1846 1043 1854 1133
rect 1846 1037 1847 1043
rect 1853 1037 1854 1043
rect 1846 999 1854 1037
rect 1846 993 1847 999
rect 1853 993 1854 999
rect 1846 895 1854 993
rect 1846 889 1847 895
rect 1853 889 1854 895
rect 1846 855 1854 889
rect 1846 849 1847 855
rect 1853 849 1854 855
rect 1846 751 1854 849
rect 1846 745 1847 751
rect 1853 745 1854 751
rect 1846 711 1854 745
rect 1846 705 1847 711
rect 1853 705 1854 711
rect 1846 607 1854 705
rect 1846 601 1847 607
rect 1853 601 1854 607
rect 1846 563 1854 601
rect 1846 557 1847 563
rect 1853 557 1854 563
rect 1846 455 1854 557
rect 1846 449 1847 455
rect 1853 449 1854 455
rect 1846 419 1854 449
rect 1846 413 1847 419
rect 1853 413 1854 419
rect 1846 319 1854 413
rect 1846 313 1847 319
rect 1853 313 1854 319
rect 1846 263 1854 313
rect 1846 257 1847 263
rect 1853 257 1854 263
rect 1846 151 1854 257
rect 1846 145 1847 151
rect 1853 145 1854 151
rect 1846 72 1854 145
rect 3598 3595 3606 3672
rect 3598 3589 3599 3595
rect 3605 3589 3606 3595
rect 3598 3451 3606 3589
rect 3598 3445 3599 3451
rect 3605 3445 3606 3451
rect 3598 3307 3606 3445
rect 3598 3301 3599 3307
rect 3605 3301 3606 3307
rect 3598 3159 3606 3301
rect 3598 3153 3599 3159
rect 3605 3153 3606 3159
rect 3598 3011 3606 3153
rect 3598 3005 3599 3011
rect 3605 3005 3606 3011
rect 3598 2867 3606 3005
rect 3598 2861 3599 2867
rect 3605 2861 3606 2867
rect 3598 2727 3606 2861
rect 3598 2721 3599 2727
rect 3605 2721 3606 2727
rect 3598 2579 3606 2721
rect 3598 2573 3599 2579
rect 3605 2573 3606 2579
rect 3598 2439 3606 2573
rect 3598 2433 3599 2439
rect 3605 2433 3606 2439
rect 3598 2295 3606 2433
rect 3598 2289 3599 2295
rect 3605 2289 3606 2295
rect 3598 2151 3606 2289
rect 3598 2145 3599 2151
rect 3605 2145 3606 2151
rect 3598 2011 3606 2145
rect 3598 2005 3599 2011
rect 3605 2005 3606 2011
rect 3598 1859 3606 2005
rect 3598 1853 3599 1859
rect 3605 1853 3606 1859
rect 3598 1715 3606 1853
rect 3598 1709 3599 1715
rect 3605 1709 3606 1715
rect 3598 1575 3606 1709
rect 3598 1569 3599 1575
rect 3605 1569 3606 1575
rect 3598 1427 3606 1569
rect 3598 1421 3599 1427
rect 3605 1421 3606 1427
rect 3598 1275 3606 1421
rect 3598 1269 3599 1275
rect 3605 1269 3606 1275
rect 3598 1123 3606 1269
rect 3598 1117 3599 1123
rect 3605 1117 3606 1123
rect 3598 971 3606 1117
rect 3598 965 3599 971
rect 3605 965 3606 971
rect 3598 819 3606 965
rect 3598 813 3599 819
rect 3605 813 3606 819
rect 3598 679 3606 813
rect 3598 673 3599 679
rect 3605 673 3606 679
rect 3598 531 3606 673
rect 3598 525 3599 531
rect 3605 525 3606 531
rect 3598 387 3606 525
rect 3598 381 3599 387
rect 3605 381 3606 387
rect 3598 251 3606 381
rect 3598 245 3599 251
rect 3605 245 3606 251
rect 3598 83 3606 245
rect 3598 77 3599 83
rect 3605 77 3606 83
rect 3598 72 3606 77
rect 3610 3527 3618 3672
rect 3610 3521 3611 3527
rect 3617 3521 3618 3527
rect 3610 3375 3618 3521
rect 3610 3369 3611 3375
rect 3617 3369 3618 3375
rect 3610 3231 3618 3369
rect 3610 3225 3611 3231
rect 3617 3225 3618 3231
rect 3610 3083 3618 3225
rect 3610 3077 3611 3083
rect 3617 3077 3618 3083
rect 3610 2935 3618 3077
rect 3610 2929 3611 2935
rect 3617 2929 3618 2935
rect 3610 2799 3618 2929
rect 3610 2793 3611 2799
rect 3617 2793 3618 2799
rect 3610 2651 3618 2793
rect 3610 2645 3611 2651
rect 3617 2645 3618 2651
rect 3610 2507 3618 2645
rect 3610 2501 3611 2507
rect 3617 2501 3618 2507
rect 3610 2367 3618 2501
rect 3610 2361 3611 2367
rect 3617 2361 3618 2367
rect 3610 2227 3618 2361
rect 3610 2221 3611 2227
rect 3617 2221 3618 2227
rect 3610 2079 3618 2221
rect 3610 2073 3611 2079
rect 3617 2073 3618 2079
rect 3610 1935 3618 2073
rect 3610 1929 3611 1935
rect 3617 1929 3618 1935
rect 3610 1787 3618 1929
rect 3610 1781 3611 1787
rect 3617 1781 3618 1787
rect 3610 1643 3618 1781
rect 3610 1637 3611 1643
rect 3617 1637 3618 1643
rect 3610 1499 3618 1637
rect 3610 1493 3611 1499
rect 3617 1493 3618 1499
rect 3610 1355 3618 1493
rect 3610 1349 3611 1355
rect 3617 1349 3618 1355
rect 3610 1203 3618 1349
rect 3610 1197 3611 1203
rect 3617 1197 3618 1203
rect 3610 1043 3618 1197
rect 3610 1037 3611 1043
rect 3617 1037 3618 1043
rect 3610 895 3618 1037
rect 3610 889 3611 895
rect 3617 889 3618 895
rect 3610 751 3618 889
rect 3610 745 3611 751
rect 3617 745 3618 751
rect 3610 607 3618 745
rect 3610 601 3611 607
rect 3617 601 3618 607
rect 3610 455 3618 601
rect 3610 449 3611 455
rect 3617 449 3618 455
rect 3610 319 3618 449
rect 3610 313 3611 319
rect 3617 313 3618 319
rect 3610 151 3618 313
rect 3610 145 3611 151
rect 3617 145 3618 151
rect 3610 72 3618 145
use circuitwell  npwells
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use circuitppnp  ppnps
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use welltap_svt  __well_tap__191
timestamp 1731220586
transform 1 0 3568 0 -1 3576
box 7 3 12 24
use welltap_svt  __well_tap__190
timestamp 1731220586
transform 1 0 1856 0 -1 3576
box 7 3 12 24
use welltap_svt  __well_tap__189
timestamp 1731220586
transform 1 0 3568 0 1 3472
box 7 3 12 24
use welltap_svt  __well_tap__188
timestamp 1731220586
transform 1 0 1856 0 1 3472
box 7 3 12 24
use welltap_svt  __well_tap__187
timestamp 1731220586
transform 1 0 3568 0 -1 3432
box 7 3 12 24
use welltap_svt  __well_tap__186
timestamp 1731220586
transform 1 0 1856 0 -1 3432
box 7 3 12 24
use welltap_svt  __well_tap__185
timestamp 1731220586
transform 1 0 3568 0 1 3320
box 7 3 12 24
use welltap_svt  __well_tap__184
timestamp 1731220586
transform 1 0 1856 0 1 3320
box 7 3 12 24
use welltap_svt  __well_tap__183
timestamp 1731220586
transform 1 0 3568 0 -1 3288
box 7 3 12 24
use welltap_svt  __well_tap__182
timestamp 1731220586
transform 1 0 1856 0 -1 3288
box 7 3 12 24
use welltap_svt  __well_tap__181
timestamp 1731220586
transform 1 0 3568 0 1 3176
box 7 3 12 24
use welltap_svt  __well_tap__180
timestamp 1731220586
transform 1 0 1856 0 1 3176
box 7 3 12 24
use welltap_svt  __well_tap__179
timestamp 1731220586
transform 1 0 3568 0 -1 3140
box 7 3 12 24
use welltap_svt  __well_tap__178
timestamp 1731220586
transform 1 0 1856 0 -1 3140
box 7 3 12 24
use welltap_svt  __well_tap__177
timestamp 1731220586
transform 1 0 3568 0 1 3028
box 7 3 12 24
use welltap_svt  __well_tap__176
timestamp 1731220586
transform 1 0 1856 0 1 3028
box 7 3 12 24
use welltap_svt  __well_tap__175
timestamp 1731220586
transform 1 0 3568 0 -1 2992
box 7 3 12 24
use welltap_svt  __well_tap__174
timestamp 1731220586
transform 1 0 1856 0 -1 2992
box 7 3 12 24
use welltap_svt  __well_tap__173
timestamp 1731220586
transform 1 0 3568 0 1 2880
box 7 3 12 24
use welltap_svt  __well_tap__172
timestamp 1731220586
transform 1 0 1856 0 1 2880
box 7 3 12 24
use welltap_svt  __well_tap__171
timestamp 1731220586
transform 1 0 3568 0 -1 2848
box 7 3 12 24
use welltap_svt  __well_tap__170
timestamp 1731220586
transform 1 0 1856 0 -1 2848
box 7 3 12 24
use welltap_svt  __well_tap__169
timestamp 1731220586
transform 1 0 3568 0 1 2744
box 7 3 12 24
use welltap_svt  __well_tap__168
timestamp 1731220586
transform 1 0 1856 0 1 2744
box 7 3 12 24
use welltap_svt  __well_tap__167
timestamp 1731220586
transform 1 0 3568 0 -1 2708
box 7 3 12 24
use welltap_svt  __well_tap__166
timestamp 1731220586
transform 1 0 1856 0 -1 2708
box 7 3 12 24
use welltap_svt  __well_tap__165
timestamp 1731220586
transform 1 0 3568 0 1 2596
box 7 3 12 24
use welltap_svt  __well_tap__164
timestamp 1731220586
transform 1 0 1856 0 1 2596
box 7 3 12 24
use welltap_svt  __well_tap__163
timestamp 1731220586
transform 1 0 3568 0 -1 2560
box 7 3 12 24
use welltap_svt  __well_tap__162
timestamp 1731220586
transform 1 0 1856 0 -1 2560
box 7 3 12 24
use welltap_svt  __well_tap__161
timestamp 1731220586
transform 1 0 3568 0 1 2452
box 7 3 12 24
use welltap_svt  __well_tap__160
timestamp 1731220586
transform 1 0 1856 0 1 2452
box 7 3 12 24
use welltap_svt  __well_tap__159
timestamp 1731220586
transform 1 0 3568 0 -1 2420
box 7 3 12 24
use welltap_svt  __well_tap__158
timestamp 1731220586
transform 1 0 1856 0 -1 2420
box 7 3 12 24
use welltap_svt  __well_tap__157
timestamp 1731220586
transform 1 0 3568 0 1 2312
box 7 3 12 24
use welltap_svt  __well_tap__156
timestamp 1731220586
transform 1 0 1856 0 1 2312
box 7 3 12 24
use welltap_svt  __well_tap__155
timestamp 1731220586
transform 1 0 3568 0 -1 2276
box 7 3 12 24
use welltap_svt  __well_tap__154
timestamp 1731220586
transform 1 0 1856 0 -1 2276
box 7 3 12 24
use welltap_svt  __well_tap__153
timestamp 1731220586
transform 1 0 3568 0 1 2172
box 7 3 12 24
use welltap_svt  __well_tap__152
timestamp 1731220586
transform 1 0 1856 0 1 2172
box 7 3 12 24
use welltap_svt  __well_tap__151
timestamp 1731220586
transform 1 0 3568 0 -1 2132
box 7 3 12 24
use welltap_svt  __well_tap__150
timestamp 1731220586
transform 1 0 1856 0 -1 2132
box 7 3 12 24
use welltap_svt  __well_tap__149
timestamp 1731220586
transform 1 0 3568 0 1 2024
box 7 3 12 24
use welltap_svt  __well_tap__148
timestamp 1731220586
transform 1 0 1856 0 1 2024
box 7 3 12 24
use welltap_svt  __well_tap__147
timestamp 1731220586
transform 1 0 3568 0 -1 1992
box 7 3 12 24
use welltap_svt  __well_tap__146
timestamp 1731220586
transform 1 0 1856 0 -1 1992
box 7 3 12 24
use welltap_svt  __well_tap__145
timestamp 1731220586
transform 1 0 3568 0 1 1880
box 7 3 12 24
use welltap_svt  __well_tap__144
timestamp 1731220586
transform 1 0 1856 0 1 1880
box 7 3 12 24
use welltap_svt  __well_tap__143
timestamp 1731220586
transform 1 0 3568 0 -1 1840
box 7 3 12 24
use welltap_svt  __well_tap__142
timestamp 1731220586
transform 1 0 1856 0 -1 1840
box 7 3 12 24
use welltap_svt  __well_tap__141
timestamp 1731220586
transform 1 0 3568 0 1 1732
box 7 3 12 24
use welltap_svt  __well_tap__140
timestamp 1731220586
transform 1 0 1856 0 1 1732
box 7 3 12 24
use welltap_svt  __well_tap__139
timestamp 1731220586
transform 1 0 3568 0 -1 1696
box 7 3 12 24
use welltap_svt  __well_tap__138
timestamp 1731220586
transform 1 0 1856 0 -1 1696
box 7 3 12 24
use welltap_svt  __well_tap__137
timestamp 1731220586
transform 1 0 3568 0 1 1588
box 7 3 12 24
use welltap_svt  __well_tap__136
timestamp 1731220586
transform 1 0 1856 0 1 1588
box 7 3 12 24
use welltap_svt  __well_tap__135
timestamp 1731220586
transform 1 0 3568 0 -1 1556
box 7 3 12 24
use welltap_svt  __well_tap__134
timestamp 1731220586
transform 1 0 1856 0 -1 1556
box 7 3 12 24
use welltap_svt  __well_tap__133
timestamp 1731220586
transform 1 0 3568 0 1 1444
box 7 3 12 24
use welltap_svt  __well_tap__132
timestamp 1731220586
transform 1 0 1856 0 1 1444
box 7 3 12 24
use welltap_svt  __well_tap__131
timestamp 1731220586
transform 1 0 3568 0 -1 1408
box 7 3 12 24
use welltap_svt  __well_tap__130
timestamp 1731220586
transform 1 0 1856 0 -1 1408
box 7 3 12 24
use welltap_svt  __well_tap__129
timestamp 1731220586
transform 1 0 3568 0 1 1300
box 7 3 12 24
use welltap_svt  __well_tap__128
timestamp 1731220586
transform 1 0 1856 0 1 1300
box 7 3 12 24
use welltap_svt  __well_tap__127
timestamp 1731220586
transform 1 0 3568 0 -1 1256
box 7 3 12 24
use welltap_svt  __well_tap__126
timestamp 1731220586
transform 1 0 1856 0 -1 1256
box 7 3 12 24
use welltap_svt  __well_tap__125
timestamp 1731220586
transform 1 0 3568 0 1 1148
box 7 3 12 24
use welltap_svt  __well_tap__124
timestamp 1731220586
transform 1 0 1856 0 1 1148
box 7 3 12 24
use welltap_svt  __well_tap__123
timestamp 1731220586
transform 1 0 3568 0 -1 1104
box 7 3 12 24
use welltap_svt  __well_tap__122
timestamp 1731220586
transform 1 0 1856 0 -1 1104
box 7 3 12 24
use welltap_svt  __well_tap__121
timestamp 1731220586
transform 1 0 3568 0 1 988
box 7 3 12 24
use welltap_svt  __well_tap__120
timestamp 1731220586
transform 1 0 1856 0 1 988
box 7 3 12 24
use welltap_svt  __well_tap__119
timestamp 1731220586
transform 1 0 3568 0 -1 952
box 7 3 12 24
use welltap_svt  __well_tap__118
timestamp 1731220586
transform 1 0 1856 0 -1 952
box 7 3 12 24
use welltap_svt  __well_tap__117
timestamp 1731220586
transform 1 0 3568 0 1 840
box 7 3 12 24
use welltap_svt  __well_tap__116
timestamp 1731220586
transform 1 0 1856 0 1 840
box 7 3 12 24
use welltap_svt  __well_tap__115
timestamp 1731220586
transform 1 0 3568 0 -1 800
box 7 3 12 24
use welltap_svt  __well_tap__114
timestamp 1731220586
transform 1 0 1856 0 -1 800
box 7 3 12 24
use welltap_svt  __well_tap__113
timestamp 1731220586
transform 1 0 3568 0 1 696
box 7 3 12 24
use welltap_svt  __well_tap__112
timestamp 1731220586
transform 1 0 1856 0 1 696
box 7 3 12 24
use welltap_svt  __well_tap__111
timestamp 1731220586
transform 1 0 3568 0 -1 660
box 7 3 12 24
use welltap_svt  __well_tap__110
timestamp 1731220586
transform 1 0 1856 0 -1 660
box 7 3 12 24
use welltap_svt  __well_tap__109
timestamp 1731220586
transform 1 0 3568 0 1 552
box 7 3 12 24
use welltap_svt  __well_tap__108
timestamp 1731220586
transform 1 0 1856 0 1 552
box 7 3 12 24
use welltap_svt  __well_tap__107
timestamp 1731220586
transform 1 0 3568 0 -1 512
box 7 3 12 24
use welltap_svt  __well_tap__106
timestamp 1731220586
transform 1 0 1856 0 -1 512
box 7 3 12 24
use welltap_svt  __well_tap__105
timestamp 1731220586
transform 1 0 3568 0 1 400
box 7 3 12 24
use welltap_svt  __well_tap__104
timestamp 1731220586
transform 1 0 1856 0 1 400
box 7 3 12 24
use welltap_svt  __well_tap__103
timestamp 1731220586
transform 1 0 3568 0 -1 368
box 7 3 12 24
use welltap_svt  __well_tap__102
timestamp 1731220586
transform 1 0 1856 0 -1 368
box 7 3 12 24
use welltap_svt  __well_tap__101
timestamp 1731220586
transform 1 0 3568 0 1 264
box 7 3 12 24
use welltap_svt  __well_tap__100
timestamp 1731220586
transform 1 0 1856 0 1 264
box 7 3 12 24
use welltap_svt  __well_tap__99
timestamp 1731220586
transform 1 0 3568 0 -1 232
box 7 3 12 24
use welltap_svt  __well_tap__98
timestamp 1731220586
transform 1 0 1856 0 -1 232
box 7 3 12 24
use welltap_svt  __well_tap__97
timestamp 1731220586
transform 1 0 3568 0 1 96
box 7 3 12 24
use welltap_svt  __well_tap__96
timestamp 1731220586
transform 1 0 1856 0 1 96
box 7 3 12 24
use welltap_svt  __well_tap__95
timestamp 1731220586
transform 1 0 1816 0 -1 3652
box 7 3 12 24
use welltap_svt  __well_tap__94
timestamp 1731220586
transform 1 0 104 0 -1 3652
box 7 3 12 24
use welltap_svt  __well_tap__93
timestamp 1731220586
transform 1 0 1816 0 1 3548
box 7 3 12 24
use welltap_svt  __well_tap__92
timestamp 1731220586
transform 1 0 104 0 1 3548
box 7 3 12 24
use welltap_svt  __well_tap__91
timestamp 1731220586
transform 1 0 1816 0 -1 3516
box 7 3 12 24
use welltap_svt  __well_tap__90
timestamp 1731220586
transform 1 0 104 0 -1 3516
box 7 3 12 24
use welltap_svt  __well_tap__89
timestamp 1731220586
transform 1 0 1816 0 1 3412
box 7 3 12 24
use welltap_svt  __well_tap__88
timestamp 1731220586
transform 1 0 104 0 1 3412
box 7 3 12 24
use welltap_svt  __well_tap__87
timestamp 1731220586
transform 1 0 1816 0 -1 3380
box 7 3 12 24
use welltap_svt  __well_tap__86
timestamp 1731220586
transform 1 0 104 0 -1 3380
box 7 3 12 24
use welltap_svt  __well_tap__85
timestamp 1731220586
transform 1 0 1816 0 1 3272
box 7 3 12 24
use welltap_svt  __well_tap__84
timestamp 1731220586
transform 1 0 104 0 1 3272
box 7 3 12 24
use welltap_svt  __well_tap__83
timestamp 1731220586
transform 1 0 1816 0 -1 3236
box 7 3 12 24
use welltap_svt  __well_tap__82
timestamp 1731220586
transform 1 0 104 0 -1 3236
box 7 3 12 24
use welltap_svt  __well_tap__81
timestamp 1731220586
transform 1 0 1816 0 1 3124
box 7 3 12 24
use welltap_svt  __well_tap__80
timestamp 1731220586
transform 1 0 104 0 1 3124
box 7 3 12 24
use welltap_svt  __well_tap__79
timestamp 1731220586
transform 1 0 1816 0 -1 3084
box 7 3 12 24
use welltap_svt  __well_tap__78
timestamp 1731220586
transform 1 0 104 0 -1 3084
box 7 3 12 24
use welltap_svt  __well_tap__77
timestamp 1731220586
transform 1 0 1816 0 1 2976
box 7 3 12 24
use welltap_svt  __well_tap__76
timestamp 1731220586
transform 1 0 104 0 1 2976
box 7 3 12 24
use welltap_svt  __well_tap__75
timestamp 1731220586
transform 1 0 1816 0 -1 2944
box 7 3 12 24
use welltap_svt  __well_tap__74
timestamp 1731220586
transform 1 0 104 0 -1 2944
box 7 3 12 24
use welltap_svt  __well_tap__73
timestamp 1731220586
transform 1 0 1816 0 1 2836
box 7 3 12 24
use welltap_svt  __well_tap__72
timestamp 1731220586
transform 1 0 104 0 1 2836
box 7 3 12 24
use welltap_svt  __well_tap__71
timestamp 1731220586
transform 1 0 1816 0 -1 2796
box 7 3 12 24
use welltap_svt  __well_tap__70
timestamp 1731220586
transform 1 0 104 0 -1 2796
box 7 3 12 24
use welltap_svt  __well_tap__69
timestamp 1731220586
transform 1 0 1816 0 1 2684
box 7 3 12 24
use welltap_svt  __well_tap__68
timestamp 1731220586
transform 1 0 104 0 1 2684
box 7 3 12 24
use welltap_svt  __well_tap__67
timestamp 1731220586
transform 1 0 1816 0 -1 2648
box 7 3 12 24
use welltap_svt  __well_tap__66
timestamp 1731220586
transform 1 0 104 0 -1 2648
box 7 3 12 24
use welltap_svt  __well_tap__65
timestamp 1731220586
transform 1 0 1816 0 1 2540
box 7 3 12 24
use welltap_svt  __well_tap__64
timestamp 1731220586
transform 1 0 104 0 1 2540
box 7 3 12 24
use welltap_svt  __well_tap__63
timestamp 1731220586
transform 1 0 1816 0 -1 2508
box 7 3 12 24
use welltap_svt  __well_tap__62
timestamp 1731220586
transform 1 0 104 0 -1 2508
box 7 3 12 24
use welltap_svt  __well_tap__61
timestamp 1731220586
transform 1 0 1816 0 1 2404
box 7 3 12 24
use welltap_svt  __well_tap__60
timestamp 1731220586
transform 1 0 104 0 1 2404
box 7 3 12 24
use welltap_svt  __well_tap__59
timestamp 1731220586
transform 1 0 1816 0 -1 2360
box 7 3 12 24
use welltap_svt  __well_tap__58
timestamp 1731220586
transform 1 0 104 0 -1 2360
box 7 3 12 24
use welltap_svt  __well_tap__57
timestamp 1731220586
transform 1 0 1816 0 1 2248
box 7 3 12 24
use welltap_svt  __well_tap__56
timestamp 1731220586
transform 1 0 104 0 1 2248
box 7 3 12 24
use welltap_svt  __well_tap__55
timestamp 1731220586
transform 1 0 1816 0 -1 2208
box 7 3 12 24
use welltap_svt  __well_tap__54
timestamp 1731220586
transform 1 0 104 0 -1 2208
box 7 3 12 24
use welltap_svt  __well_tap__53
timestamp 1731220586
transform 1 0 1816 0 1 2104
box 7 3 12 24
use welltap_svt  __well_tap__52
timestamp 1731220586
transform 1 0 104 0 1 2104
box 7 3 12 24
use welltap_svt  __well_tap__51
timestamp 1731220586
transform 1 0 1816 0 -1 2068
box 7 3 12 24
use welltap_svt  __well_tap__50
timestamp 1731220586
transform 1 0 104 0 -1 2068
box 7 3 12 24
use welltap_svt  __well_tap__49
timestamp 1731220586
transform 1 0 1816 0 1 1960
box 7 3 12 24
use welltap_svt  __well_tap__48
timestamp 1731220586
transform 1 0 104 0 1 1960
box 7 3 12 24
use welltap_svt  __well_tap__47
timestamp 1731220586
transform 1 0 1816 0 -1 1924
box 7 3 12 24
use welltap_svt  __well_tap__46
timestamp 1731220586
transform 1 0 104 0 -1 1924
box 7 3 12 24
use welltap_svt  __well_tap__45
timestamp 1731220586
transform 1 0 1816 0 1 1812
box 7 3 12 24
use welltap_svt  __well_tap__44
timestamp 1731220586
transform 1 0 104 0 1 1812
box 7 3 12 24
use welltap_svt  __well_tap__43
timestamp 1731220586
transform 1 0 1816 0 -1 1768
box 7 3 12 24
use welltap_svt  __well_tap__42
timestamp 1731220586
transform 1 0 104 0 -1 1768
box 7 3 12 24
use welltap_svt  __well_tap__41
timestamp 1731220586
transform 1 0 1816 0 1 1660
box 7 3 12 24
use welltap_svt  __well_tap__40
timestamp 1731220586
transform 1 0 104 0 1 1660
box 7 3 12 24
use welltap_svt  __well_tap__39
timestamp 1731220586
transform 1 0 1816 0 -1 1620
box 7 3 12 24
use welltap_svt  __well_tap__38
timestamp 1731220586
transform 1 0 104 0 -1 1620
box 7 3 12 24
use welltap_svt  __well_tap__37
timestamp 1731220586
transform 1 0 1816 0 1 1516
box 7 3 12 24
use welltap_svt  __well_tap__36
timestamp 1731220586
transform 1 0 104 0 1 1516
box 7 3 12 24
use welltap_svt  __well_tap__35
timestamp 1731220586
transform 1 0 1816 0 -1 1480
box 7 3 12 24
use welltap_svt  __well_tap__34
timestamp 1731220586
transform 1 0 104 0 -1 1480
box 7 3 12 24
use welltap_svt  __well_tap__33
timestamp 1731220586
transform 1 0 1816 0 1 1368
box 7 3 12 24
use welltap_svt  __well_tap__32
timestamp 1731220586
transform 1 0 104 0 1 1368
box 7 3 12 24
use welltap_svt  __well_tap__31
timestamp 1731220586
transform 1 0 1816 0 -1 1332
box 7 3 12 24
use welltap_svt  __well_tap__30
timestamp 1731220586
transform 1 0 104 0 -1 1332
box 7 3 12 24
use welltap_svt  __well_tap__29
timestamp 1731220586
transform 1 0 1816 0 1 1228
box 7 3 12 24
use welltap_svt  __well_tap__28
timestamp 1731220586
transform 1 0 104 0 1 1228
box 7 3 12 24
use welltap_svt  __well_tap__27
timestamp 1731220586
transform 1 0 1816 0 -1 1188
box 7 3 12 24
use welltap_svt  __well_tap__26
timestamp 1731220586
transform 1 0 104 0 -1 1188
box 7 3 12 24
use welltap_svt  __well_tap__25
timestamp 1731220586
transform 1 0 1816 0 1 1084
box 7 3 12 24
use welltap_svt  __well_tap__24
timestamp 1731220586
transform 1 0 104 0 1 1084
box 7 3 12 24
use welltap_svt  __well_tap__23
timestamp 1731220586
transform 1 0 1816 0 -1 1052
box 7 3 12 24
use welltap_svt  __well_tap__22
timestamp 1731220586
transform 1 0 104 0 -1 1052
box 7 3 12 24
use welltap_svt  __well_tap__21
timestamp 1731220586
transform 1 0 1816 0 1 944
box 7 3 12 24
use welltap_svt  __well_tap__20
timestamp 1731220586
transform 1 0 104 0 1 944
box 7 3 12 24
use welltap_svt  __well_tap__19
timestamp 1731220586
transform 1 0 1816 0 -1 904
box 7 3 12 24
use welltap_svt  __well_tap__18
timestamp 1731220586
transform 1 0 104 0 -1 904
box 7 3 12 24
use welltap_svt  __well_tap__17
timestamp 1731220586
transform 1 0 1816 0 1 800
box 7 3 12 24
use welltap_svt  __well_tap__16
timestamp 1731220586
transform 1 0 104 0 1 800
box 7 3 12 24
use welltap_svt  __well_tap__15
timestamp 1731220586
transform 1 0 1816 0 -1 764
box 7 3 12 24
use welltap_svt  __well_tap__14
timestamp 1731220586
transform 1 0 104 0 -1 764
box 7 3 12 24
use welltap_svt  __well_tap__13
timestamp 1731220586
transform 1 0 1816 0 1 656
box 7 3 12 24
use welltap_svt  __well_tap__12
timestamp 1731220586
transform 1 0 104 0 1 656
box 7 3 12 24
use welltap_svt  __well_tap__11
timestamp 1731220586
transform 1 0 1816 0 -1 616
box 7 3 12 24
use welltap_svt  __well_tap__10
timestamp 1731220586
transform 1 0 104 0 -1 616
box 7 3 12 24
use welltap_svt  __well_tap__9
timestamp 1731220586
transform 1 0 1816 0 1 508
box 7 3 12 24
use welltap_svt  __well_tap__8
timestamp 1731220586
transform 1 0 104 0 1 508
box 7 3 12 24
use welltap_svt  __well_tap__7
timestamp 1731220586
transform 1 0 1816 0 -1 468
box 7 3 12 24
use welltap_svt  __well_tap__6
timestamp 1731220586
transform 1 0 104 0 -1 468
box 7 3 12 24
use welltap_svt  __well_tap__5
timestamp 1731220586
transform 1 0 1816 0 1 364
box 7 3 12 24
use welltap_svt  __well_tap__4
timestamp 1731220586
transform 1 0 104 0 1 364
box 7 3 12 24
use welltap_svt  __well_tap__3
timestamp 1731220586
transform 1 0 1816 0 -1 316
box 7 3 12 24
use welltap_svt  __well_tap__2
timestamp 1731220586
transform 1 0 104 0 -1 316
box 7 3 12 24
use welltap_svt  __well_tap__1
timestamp 1731220586
transform 1 0 1816 0 1 208
box 7 3 12 24
use welltap_svt  __well_tap__0
timestamp 1731220586
transform 1 0 104 0 1 208
box 7 3 12 24
use _0_0std_0_0cells_0_0MUX2X1  tst_5999_6
timestamp 1731220586
transform 1 0 3384 0 1 80
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5998_6
timestamp 1731220586
transform 1 0 3472 0 1 80
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5997_6
timestamp 1731220586
transform 1 0 3472 0 -1 248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5996_6
timestamp 1731220586
transform 1 0 3456 0 1 384
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5995_6
timestamp 1731220586
transform 1 0 3424 0 -1 528
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5994_6
timestamp 1731220586
transform 1 0 3424 0 -1 384
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5993_6
timestamp 1731220586
transform 1 0 3352 0 -1 248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5992_6
timestamp 1731220586
transform 1 0 3296 0 1 80
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5991_6
timestamp 1731220586
transform 1 0 3208 0 1 80
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5990_6
timestamp 1731220586
transform 1 0 3120 0 1 80
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5989_6
timestamp 1731220586
transform 1 0 3032 0 1 80
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5988_6
timestamp 1731220586
transform 1 0 2944 0 1 80
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5987_6
timestamp 1731220586
transform 1 0 2856 0 1 80
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5986_6
timestamp 1731220586
transform 1 0 2768 0 1 80
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5985_6
timestamp 1731220586
transform 1 0 3216 0 -1 248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5984_6
timestamp 1731220586
transform 1 0 3080 0 -1 248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5983_6
timestamp 1731220586
transform 1 0 2944 0 -1 248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5982_6
timestamp 1731220586
transform 1 0 2808 0 -1 248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5981_6
timestamp 1731220586
transform 1 0 3144 0 1 248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5980_6
timestamp 1731220586
transform 1 0 3024 0 1 248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5979_6
timestamp 1731220586
transform 1 0 2904 0 1 248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5978_6
timestamp 1731220586
transform 1 0 2792 0 1 248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5977_6
timestamp 1731220586
transform 1 0 2680 0 1 248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5976_6
timestamp 1731220586
transform 1 0 3224 0 -1 384
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5975_6
timestamp 1731220586
transform 1 0 3024 0 -1 384
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5974_6
timestamp 1731220586
transform 1 0 2840 0 -1 384
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5973_6
timestamp 1731220586
transform 1 0 2664 0 -1 384
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5972_6
timestamp 1731220586
transform 1 0 3224 0 1 384
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5971_6
timestamp 1731220586
transform 1 0 2992 0 1 384
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5970_6
timestamp 1731220586
transform 1 0 2768 0 1 384
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5969_6
timestamp 1731220586
transform 1 0 2560 0 1 384
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5968_6
timestamp 1731220586
transform 1 0 2368 0 1 384
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5967_6
timestamp 1731220586
transform 1 0 3208 0 -1 528
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5966_6
timestamp 1731220586
transform 1 0 3000 0 -1 528
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5965_6
timestamp 1731220586
transform 1 0 2800 0 -1 528
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5964_6
timestamp 1731220586
transform 1 0 2624 0 -1 528
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5963_6
timestamp 1731220586
transform 1 0 2480 0 -1 528
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5962_6
timestamp 1731220586
transform 1 0 2376 0 1 536
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5961_6
timestamp 1731220586
transform 1 0 2568 0 1 536
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5960_6
timestamp 1731220586
transform 1 0 3240 0 1 536
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5959_6
timestamp 1731220586
transform 1 0 3008 0 1 536
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5958_6
timestamp 1731220586
transform 1 0 2784 0 1 536
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5957_6
timestamp 1731220586
transform 1 0 2760 0 -1 676
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5956_6
timestamp 1731220586
transform 1 0 2608 0 -1 676
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5955_6
timestamp 1731220586
transform 1 0 3304 0 -1 676
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5954_6
timestamp 1731220586
transform 1 0 3112 0 -1 676
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5953_6
timestamp 1731220586
transform 1 0 2928 0 -1 676
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5952_6
timestamp 1731220586
transform 1 0 2784 0 1 680
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5951_6
timestamp 1731220586
transform 1 0 2608 0 1 680
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5950_6
timestamp 1731220586
transform 1 0 2960 0 1 680
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5949_6
timestamp 1731220586
transform 1 0 3312 0 1 680
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5948_6
timestamp 1731220586
transform 1 0 3136 0 1 680
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5947_6
timestamp 1731220586
transform 1 0 3080 0 -1 816
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5946_6
timestamp 1731220586
transform 1 0 2936 0 -1 816
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5945_6
timestamp 1731220586
transform 1 0 2784 0 -1 816
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5944_6
timestamp 1731220586
transform 1 0 2824 0 1 824
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5943_6
timestamp 1731220586
transform 1 0 2968 0 1 824
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5942_6
timestamp 1731220586
transform 1 0 3104 0 1 824
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5941_6
timestamp 1731220586
transform 1 0 3232 0 1 824
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5940_6
timestamp 1731220586
transform 1 0 3360 0 1 824
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5939_6
timestamp 1731220586
transform 1 0 3352 0 -1 816
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5938_6
timestamp 1731220586
transform 1 0 3216 0 -1 816
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5937_6
timestamp 1731220586
transform 1 0 3472 0 -1 816
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5936_6
timestamp 1731220586
transform 1 0 3472 0 1 536
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5935_6
timestamp 1731220586
transform 1 0 3472 0 -1 676
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5934_6
timestamp 1731220586
transform 1 0 3472 0 1 680
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5933_6
timestamp 1731220586
transform 1 0 3472 0 1 824
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5932_6
timestamp 1731220586
transform 1 0 3472 0 -1 968
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5931_6
timestamp 1731220586
transform 1 0 3472 0 1 972
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5930_6
timestamp 1731220586
transform 1 0 3472 0 -1 1120
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5929_6
timestamp 1731220586
transform 1 0 3472 0 1 1132
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5928_6
timestamp 1731220586
transform 1 0 3424 0 -1 1272
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5927_6
timestamp 1731220586
transform 1 0 3472 0 1 1284
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5926_6
timestamp 1731220586
transform 1 0 3472 0 -1 1424
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5925_6
timestamp 1731220586
transform 1 0 3472 0 1 1428
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5924_6
timestamp 1731220586
transform 1 0 3472 0 1 1572
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5923_6
timestamp 1731220586
transform 1 0 3472 0 -1 1712
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5922_6
timestamp 1731220586
transform 1 0 3424 0 -1 1572
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5921_6
timestamp 1731220586
transform 1 0 3264 0 1 1284
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5920_6
timestamp 1731220586
transform 1 0 3152 0 1 1132
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5919_6
timestamp 1731220586
transform 1 0 3312 0 1 1132
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5918_6
timestamp 1731220586
transform 1 0 3312 0 -1 1120
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5917_6
timestamp 1731220586
transform 1 0 3328 0 1 972
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5916_6
timestamp 1731220586
transform 1 0 3360 0 -1 968
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5915_6
timestamp 1731220586
transform 1 0 3224 0 -1 968
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5914_6
timestamp 1731220586
transform 1 0 3088 0 -1 968
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5913_6
timestamp 1731220586
transform 1 0 2944 0 -1 968
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5912_6
timestamp 1731220586
transform 1 0 2792 0 -1 968
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5911_6
timestamp 1731220586
transform 1 0 3168 0 1 972
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5910_6
timestamp 1731220586
transform 1 0 3008 0 1 972
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5909_6
timestamp 1731220586
transform 1 0 2848 0 1 972
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5908_6
timestamp 1731220586
transform 1 0 2680 0 1 972
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5907_6
timestamp 1731220586
transform 1 0 3144 0 -1 1120
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5906_6
timestamp 1731220586
transform 1 0 2984 0 -1 1120
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5905_6
timestamp 1731220586
transform 1 0 2832 0 -1 1120
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5904_6
timestamp 1731220586
transform 1 0 2680 0 -1 1120
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5903_6
timestamp 1731220586
transform 1 0 2696 0 1 1132
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5902_6
timestamp 1731220586
transform 1 0 2848 0 1 1132
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5901_6
timestamp 1731220586
transform 1 0 3000 0 1 1132
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5900_6
timestamp 1731220586
transform 1 0 3224 0 -1 1272
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5899_6
timestamp 1731220586
transform 1 0 3032 0 -1 1272
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5898_6
timestamp 1731220586
transform 1 0 2848 0 -1 1272
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5897_6
timestamp 1731220586
transform 1 0 2680 0 -1 1272
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5896_6
timestamp 1731220586
transform 1 0 2544 0 -1 1272
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5895_6
timestamp 1731220586
transform 1 0 3056 0 1 1284
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5894_6
timestamp 1731220586
transform 1 0 2856 0 1 1284
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5893_6
timestamp 1731220586
transform 1 0 2672 0 1 1284
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5892_6
timestamp 1731220586
transform 1 0 2496 0 1 1284
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5891_6
timestamp 1731220586
transform 1 0 2344 0 1 1284
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5890_6
timestamp 1731220586
transform 1 0 2432 0 -1 1424
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5889_6
timestamp 1731220586
transform 1 0 2600 0 -1 1424
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5888_6
timestamp 1731220586
transform 1 0 3256 0 -1 1424
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5887_6
timestamp 1731220586
transform 1 0 3024 0 -1 1424
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5886_6
timestamp 1731220586
transform 1 0 2800 0 -1 1424
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5885_6
timestamp 1731220586
transform 1 0 2688 0 1 1428
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5884_6
timestamp 1731220586
transform 1 0 2520 0 1 1428
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5883_6
timestamp 1731220586
transform 1 0 2872 0 1 1428
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5882_6
timestamp 1731220586
transform 1 0 3280 0 1 1428
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5881_6
timestamp 1731220586
transform 1 0 3072 0 1 1428
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5880_6
timestamp 1731220586
transform 1 0 2944 0 -1 1572
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5879_6
timestamp 1731220586
transform 1 0 2784 0 -1 1572
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5878_6
timestamp 1731220586
transform 1 0 2616 0 -1 1572
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5877_6
timestamp 1731220586
transform 1 0 3264 0 -1 1572
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5876_6
timestamp 1731220586
transform 1 0 3104 0 -1 1572
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5875_6
timestamp 1731220586
transform 1 0 3016 0 1 1572
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5874_6
timestamp 1731220586
transform 1 0 2856 0 1 1572
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5873_6
timestamp 1731220586
transform 1 0 3176 0 1 1572
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5872_6
timestamp 1731220586
transform 1 0 3336 0 1 1572
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5871_6
timestamp 1731220586
transform 1 0 3360 0 -1 1712
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5870_6
timestamp 1731220586
transform 1 0 3240 0 -1 1712
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5869_6
timestamp 1731220586
transform 1 0 3128 0 -1 1712
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5868_6
timestamp 1731220586
transform 1 0 3008 0 -1 1712
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5867_6
timestamp 1731220586
transform 1 0 2880 0 -1 1712
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5866_6
timestamp 1731220586
transform 1 0 3160 0 1 1716
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5865_6
timestamp 1731220586
transform 1 0 3056 0 1 1716
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5864_6
timestamp 1731220586
transform 1 0 2952 0 1 1716
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5863_6
timestamp 1731220586
transform 1 0 2848 0 1 1716
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5862_6
timestamp 1731220586
transform 1 0 2744 0 1 1716
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5861_6
timestamp 1731220586
transform 1 0 2984 0 -1 1856
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5860_6
timestamp 1731220586
transform 1 0 2856 0 -1 1856
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5859_6
timestamp 1731220586
transform 1 0 2736 0 -1 1856
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5858_6
timestamp 1731220586
transform 1 0 2616 0 -1 1856
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5857_6
timestamp 1731220586
transform 1 0 2488 0 -1 1856
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5856_6
timestamp 1731220586
transform 1 0 2496 0 1 1864
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5855_6
timestamp 1731220586
transform 1 0 2616 0 1 1864
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5854_6
timestamp 1731220586
transform 1 0 2736 0 1 1864
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5853_6
timestamp 1731220586
transform 1 0 2864 0 1 1864
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5852_6
timestamp 1731220586
transform 1 0 2992 0 1 1864
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5851_6
timestamp 1731220586
transform 1 0 2864 0 -1 2008
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5850_6
timestamp 1731220586
transform 1 0 2704 0 -1 2008
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5849_6
timestamp 1731220586
transform 1 0 3200 0 -1 2008
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5848_6
timestamp 1731220586
transform 1 0 3032 0 -1 2008
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5847_6
timestamp 1731220586
transform 1 0 2896 0 1 2008
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5846_6
timestamp 1731220586
transform 1 0 2760 0 1 2008
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5845_6
timestamp 1731220586
transform 1 0 2888 0 -1 2148
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5844_6
timestamp 1731220586
transform 1 0 3016 0 -1 2148
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5843_6
timestamp 1731220586
transform 1 0 3136 0 -1 2148
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5842_6
timestamp 1731220586
transform 1 0 3256 0 -1 2148
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5841_6
timestamp 1731220586
transform 1 0 3144 0 1 2008
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5840_6
timestamp 1731220586
transform 1 0 3024 0 1 2008
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5839_6
timestamp 1731220586
transform 1 0 3264 0 1 2008
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5838_6
timestamp 1731220586
transform 1 0 3376 0 1 2008
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5837_6
timestamp 1731220586
transform 1 0 3472 0 1 2008
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5836_6
timestamp 1731220586
transform 1 0 3376 0 -1 2148
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5835_6
timestamp 1731220586
transform 1 0 3472 0 -1 2148
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5834_6
timestamp 1731220586
transform 1 0 3472 0 1 2156
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5833_6
timestamp 1731220586
transform 1 0 3472 0 -1 2292
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5832_6
timestamp 1731220586
transform 1 0 3472 0 1 2296
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5831_6
timestamp 1731220586
transform 1 0 3384 0 1 2296
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5830_6
timestamp 1731220586
transform 1 0 3272 0 1 2296
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5829_6
timestamp 1731220586
transform 1 0 3264 0 -1 2292
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5828_6
timestamp 1731220586
transform 1 0 3376 0 -1 2292
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5827_6
timestamp 1731220586
transform 1 0 3288 0 1 2156
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5826_6
timestamp 1731220586
transform 1 0 3088 0 1 2156
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5825_6
timestamp 1731220586
transform 1 0 3152 0 -1 2292
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5824_6
timestamp 1731220586
transform 1 0 3032 0 -1 2292
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5823_6
timestamp 1731220586
transform 1 0 2912 0 -1 2292
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5822_6
timestamp 1731220586
transform 1 0 2776 0 -1 2292
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5821_6
timestamp 1731220586
transform 1 0 3168 0 1 2296
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5820_6
timestamp 1731220586
transform 1 0 3056 0 1 2296
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5819_6
timestamp 1731220586
transform 1 0 2936 0 1 2296
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5818_6
timestamp 1731220586
transform 1 0 2816 0 1 2296
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5817_6
timestamp 1731220586
transform 1 0 2688 0 1 2296
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5816_6
timestamp 1731220586
transform 1 0 3104 0 -1 2436
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5815_6
timestamp 1731220586
transform 1 0 2944 0 -1 2436
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5814_6
timestamp 1731220586
transform 1 0 2792 0 -1 2436
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5813_6
timestamp 1731220586
transform 1 0 2640 0 -1 2436
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5812_6
timestamp 1731220586
transform 1 0 3000 0 1 2436
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5811_6
timestamp 1731220586
transform 1 0 2864 0 1 2436
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5810_6
timestamp 1731220586
transform 1 0 2736 0 1 2436
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5809_6
timestamp 1731220586
transform 1 0 2608 0 1 2436
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5808_6
timestamp 1731220586
transform 1 0 2472 0 1 2436
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5807_6
timestamp 1731220586
transform 1 0 2824 0 -1 2576
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5806_6
timestamp 1731220586
transform 1 0 2704 0 -1 2576
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5805_6
timestamp 1731220586
transform 1 0 2584 0 -1 2576
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5804_6
timestamp 1731220586
transform 1 0 2464 0 -1 2576
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5803_6
timestamp 1731220586
transform 1 0 2440 0 1 2580
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5802_6
timestamp 1731220586
transform 1 0 2536 0 1 2580
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5801_6
timestamp 1731220586
transform 1 0 2848 0 1 2580
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5800_6
timestamp 1731220586
transform 1 0 2744 0 1 2580
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5799_6
timestamp 1731220586
transform 1 0 2640 0 1 2580
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5798_6
timestamp 1731220586
transform 1 0 2616 0 -1 2724
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5797_6
timestamp 1731220586
transform 1 0 2736 0 -1 2724
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5796_6
timestamp 1731220586
transform 1 0 2856 0 -1 2724
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5795_6
timestamp 1731220586
transform 1 0 3096 0 -1 2724
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5794_6
timestamp 1731220586
transform 1 0 2976 0 -1 2724
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5793_6
timestamp 1731220586
transform 1 0 2920 0 1 2728
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5792_6
timestamp 1731220586
transform 1 0 2768 0 1 2728
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5791_6
timestamp 1731220586
transform 1 0 3208 0 1 2728
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5790_6
timestamp 1731220586
transform 1 0 3064 0 1 2728
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5789_6
timestamp 1731220586
transform 1 0 2928 0 -1 2864
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5788_6
timestamp 1731220586
transform 1 0 2800 0 -1 2864
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5787_6
timestamp 1731220586
transform 1 0 2664 0 -1 2864
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5786_6
timestamp 1731220586
transform 1 0 3048 0 -1 2864
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5785_6
timestamp 1731220586
transform 1 0 3152 0 1 2864
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5784_6
timestamp 1731220586
transform 1 0 3160 0 -1 2864
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5783_6
timestamp 1731220586
transform 1 0 3272 0 -1 2864
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5782_6
timestamp 1731220586
transform 1 0 3384 0 -1 2864
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5781_6
timestamp 1731220586
transform 1 0 3352 0 1 2728
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5780_6
timestamp 1731220586
transform 1 0 3472 0 1 2728
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5779_6
timestamp 1731220586
transform 1 0 3472 0 -1 2864
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5778_6
timestamp 1731220586
transform 1 0 3472 0 1 2864
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5777_6
timestamp 1731220586
transform 1 0 3472 0 -1 3008
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5776_6
timestamp 1731220586
transform 1 0 3472 0 1 3012
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5775_6
timestamp 1731220586
transform 1 0 3472 0 -1 3156
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5774_6
timestamp 1731220586
transform 1 0 3472 0 1 3160
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5773_6
timestamp 1731220586
transform 1 0 3472 0 -1 3304
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5772_6
timestamp 1731220586
transform 1 0 3304 0 -1 3304
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5771_6
timestamp 1731220586
transform 1 0 3472 0 1 3304
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5770_6
timestamp 1731220586
transform 1 0 3328 0 1 3304
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5769_6
timestamp 1731220586
transform 1 0 3176 0 1 3304
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5768_6
timestamp 1731220586
transform 1 0 3024 0 1 3304
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5767_6
timestamp 1731220586
transform 1 0 3352 0 -1 3448
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5766_6
timestamp 1731220586
transform 1 0 3184 0 -1 3448
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5765_6
timestamp 1731220586
transform 1 0 3024 0 -1 3448
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5764_6
timestamp 1731220586
transform 1 0 2864 0 -1 3448
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5763_6
timestamp 1731220586
transform 1 0 2920 0 1 3456
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5762_6
timestamp 1731220586
transform 1 0 3064 0 1 3456
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5761_6
timestamp 1731220586
transform 1 0 3208 0 1 3456
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5760_6
timestamp 1731220586
transform 1 0 3216 0 -1 3592
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5759_6
timestamp 1731220586
transform 1 0 3112 0 -1 3592
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5758_6
timestamp 1731220586
transform 1 0 3008 0 -1 3592
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5757_6
timestamp 1731220586
transform 1 0 2912 0 -1 3592
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5756_6
timestamp 1731220586
transform 1 0 2816 0 -1 3592
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5755_6
timestamp 1731220586
transform 1 0 2720 0 -1 3592
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5754_6
timestamp 1731220586
transform 1 0 2624 0 -1 3592
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5753_6
timestamp 1731220586
transform 1 0 2640 0 1 3456
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5752_6
timestamp 1731220586
transform 1 0 2776 0 1 3456
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5751_6
timestamp 1731220586
transform 1 0 2704 0 -1 3448
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5750_6
timestamp 1731220586
transform 1 0 2704 0 1 3304
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5749_6
timestamp 1731220586
transform 1 0 2864 0 1 3304
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5748_6
timestamp 1731220586
transform 1 0 2792 0 -1 3304
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5747_6
timestamp 1731220586
transform 1 0 2960 0 -1 3304
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5746_6
timestamp 1731220586
transform 1 0 3128 0 -1 3304
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5745_6
timestamp 1731220586
transform 1 0 3312 0 1 3160
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5744_6
timestamp 1731220586
transform 1 0 3152 0 1 3160
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5743_6
timestamp 1731220586
transform 1 0 3000 0 1 3160
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5742_6
timestamp 1731220586
transform 1 0 2856 0 1 3160
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5741_6
timestamp 1731220586
transform 1 0 2720 0 1 3160
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5740_6
timestamp 1731220586
transform 1 0 2864 0 -1 3156
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5739_6
timestamp 1731220586
transform 1 0 3064 0 -1 3156
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5738_6
timestamp 1731220586
transform 1 0 3280 0 -1 3156
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5737_6
timestamp 1731220586
transform 1 0 3224 0 1 3012
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5736_6
timestamp 1731220586
transform 1 0 3312 0 -1 3008
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5735_6
timestamp 1731220586
transform 1 0 3136 0 -1 3008
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5734_6
timestamp 1731220586
transform 1 0 2960 0 -1 3008
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5733_6
timestamp 1731220586
transform 1 0 2800 0 -1 3008
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5732_6
timestamp 1731220586
transform 1 0 2656 0 -1 3008
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5731_6
timestamp 1731220586
transform 1 0 2528 0 -1 3008
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5730_6
timestamp 1731220586
transform 1 0 2408 0 -1 3008
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5729_6
timestamp 1731220586
transform 1 0 2472 0 1 3012
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5728_6
timestamp 1731220586
transform 1 0 2960 0 1 3012
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5727_6
timestamp 1731220586
transform 1 0 2704 0 1 3012
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5726_6
timestamp 1731220586
transform 1 0 2672 0 -1 3156
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5725_6
timestamp 1731220586
transform 1 0 2504 0 -1 3156
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5724_6
timestamp 1731220586
transform 1 0 2344 0 -1 3156
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5723_6
timestamp 1731220586
transform 1 0 2192 0 -1 3156
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5722_6
timestamp 1731220586
transform 1 0 2584 0 1 3160
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5721_6
timestamp 1731220586
transform 1 0 2448 0 1 3160
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5720_6
timestamp 1731220586
transform 1 0 2312 0 1 3160
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5719_6
timestamp 1731220586
transform 1 0 2160 0 1 3160
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5718_6
timestamp 1731220586
transform 1 0 2624 0 -1 3304
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5717_6
timestamp 1731220586
transform 1 0 2456 0 -1 3304
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5716_6
timestamp 1731220586
transform 1 0 2296 0 -1 3304
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5715_6
timestamp 1731220586
transform 1 0 2144 0 -1 3304
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5714_6
timestamp 1731220586
transform 1 0 2536 0 1 3304
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5713_6
timestamp 1731220586
transform 1 0 2360 0 1 3304
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5712_6
timestamp 1731220586
transform 1 0 2184 0 1 3304
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5711_6
timestamp 1731220586
transform 1 0 2016 0 1 3304
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5710_6
timestamp 1731220586
transform 1 0 2184 0 -1 3448
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5709_6
timestamp 1731220586
transform 1 0 2360 0 -1 3448
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5708_6
timestamp 1731220586
transform 1 0 2536 0 -1 3448
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5707_6
timestamp 1731220586
transform 1 0 2496 0 1 3456
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5706_6
timestamp 1731220586
transform 1 0 2352 0 1 3456
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5705_6
timestamp 1731220586
transform 1 0 2216 0 1 3456
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5704_6
timestamp 1731220586
transform 1 0 2088 0 1 3456
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5703_6
timestamp 1731220586
transform 1 0 2528 0 -1 3592
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5702_6
timestamp 1731220586
transform 1 0 2424 0 -1 3592
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5701_6
timestamp 1731220586
transform 1 0 2320 0 -1 3592
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5700_6
timestamp 1731220586
transform 1 0 2232 0 -1 3592
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5699_6
timestamp 1731220586
transform 1 0 2144 0 -1 3592
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5698_6
timestamp 1731220586
transform 1 0 2056 0 -1 3592
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5697_6
timestamp 1731220586
transform 1 0 1968 0 -1 3592
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5696_6
timestamp 1731220586
transform 1 0 1880 0 -1 3592
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5695_6
timestamp 1731220586
transform 1 0 1880 0 1 3456
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5694_6
timestamp 1731220586
transform 1 0 1968 0 1 3456
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5693_6
timestamp 1731220586
transform 1 0 2016 0 -1 3448
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5692_6
timestamp 1731220586
transform 1 0 1880 0 -1 3448
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5691_6
timestamp 1731220586
transform 1 0 1880 0 1 3304
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5690_6
timestamp 1731220586
transform 1 0 1880 0 -1 3304
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5689_6
timestamp 1731220586
transform 1 0 2000 0 -1 3304
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5688_6
timestamp 1731220586
transform 1 0 1880 0 1 3160
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5687_6
timestamp 1731220586
transform 1 0 2008 0 1 3160
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5686_6
timestamp 1731220586
transform 1 0 2040 0 -1 3156
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5685_6
timestamp 1731220586
transform 1 0 1880 0 -1 3156
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5684_6
timestamp 1731220586
transform 1 0 1904 0 1 3012
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5683_6
timestamp 1731220586
transform 1 0 2072 0 1 3012
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5682_6
timestamp 1731220586
transform 1 0 2264 0 1 3012
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5681_6
timestamp 1731220586
transform 1 0 2280 0 -1 3008
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5680_6
timestamp 1731220586
transform 1 0 2152 0 -1 3008
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5679_6
timestamp 1731220586
transform 1 0 2016 0 -1 3008
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5678_6
timestamp 1731220586
transform 1 0 2160 0 1 2864
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5677_6
timestamp 1731220586
transform 1 0 2480 0 1 2864
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5676_6
timestamp 1731220586
transform 1 0 2808 0 1 2864
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5675_6
timestamp 1731220586
transform 1 0 2512 0 -1 2864
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5674_6
timestamp 1731220586
transform 1 0 2352 0 -1 2864
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5673_6
timestamp 1731220586
transform 1 0 2184 0 -1 2864
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5672_6
timestamp 1731220586
transform 1 0 2240 0 1 2728
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5671_6
timestamp 1731220586
transform 1 0 2424 0 1 2728
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5670_6
timestamp 1731220586
transform 1 0 2600 0 1 2728
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5669_6
timestamp 1731220586
transform 1 0 2488 0 -1 2724
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5668_6
timestamp 1731220586
transform 1 0 2352 0 -1 2724
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5667_6
timestamp 1731220586
transform 1 0 2200 0 -1 2724
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5666_6
timestamp 1731220586
transform 1 0 2336 0 1 2580
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5665_6
timestamp 1731220586
transform 1 0 2224 0 1 2580
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5664_6
timestamp 1731220586
transform 1 0 2104 0 1 2580
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5663_6
timestamp 1731220586
transform 1 0 2104 0 -1 2576
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5662_6
timestamp 1731220586
transform 1 0 2224 0 -1 2576
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5661_6
timestamp 1731220586
transform 1 0 2344 0 -1 2576
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5660_6
timestamp 1731220586
transform 1 0 2328 0 1 2436
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5659_6
timestamp 1731220586
transform 1 0 2176 0 1 2436
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5658_6
timestamp 1731220586
transform 1 0 2168 0 -1 2436
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5657_6
timestamp 1731220586
transform 1 0 2328 0 -1 2436
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5656_6
timestamp 1731220586
transform 1 0 2488 0 -1 2436
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5655_6
timestamp 1731220586
transform 1 0 2392 0 1 2296
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5654_6
timestamp 1731220586
transform 1 0 2232 0 1 2296
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5653_6
timestamp 1731220586
transform 1 0 2544 0 1 2296
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5652_6
timestamp 1731220586
transform 1 0 2632 0 -1 2292
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5651_6
timestamp 1731220586
transform 1 0 2472 0 -1 2292
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5650_6
timestamp 1731220586
transform 1 0 2304 0 -1 2292
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5649_6
timestamp 1731220586
transform 1 0 2504 0 1 2156
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5648_6
timestamp 1731220586
transform 1 0 2696 0 1 2156
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5647_6
timestamp 1731220586
transform 1 0 2888 0 1 2156
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5646_6
timestamp 1731220586
transform 1 0 2752 0 -1 2148
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5645_6
timestamp 1731220586
transform 1 0 2608 0 -1 2148
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5644_6
timestamp 1731220586
transform 1 0 2464 0 -1 2148
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5643_6
timestamp 1731220586
transform 1 0 2312 0 -1 2148
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5642_6
timestamp 1731220586
transform 1 0 2296 0 1 2008
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5641_6
timestamp 1731220586
transform 1 0 2456 0 1 2008
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5640_6
timestamp 1731220586
transform 1 0 2616 0 1 2008
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5639_6
timestamp 1731220586
transform 1 0 2536 0 -1 2008
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5638_6
timestamp 1731220586
transform 1 0 2368 0 -1 2008
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5637_6
timestamp 1731220586
transform 1 0 2240 0 1 1864
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5636_6
timestamp 1731220586
transform 1 0 2368 0 1 1864
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5635_6
timestamp 1731220586
transform 1 0 2352 0 -1 1856
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5634_6
timestamp 1731220586
transform 1 0 2216 0 -1 1856
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5633_6
timestamp 1731220586
transform 1 0 2256 0 1 1716
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5632_6
timestamp 1731220586
transform 1 0 2344 0 1 1716
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5631_6
timestamp 1731220586
transform 1 0 2440 0 1 1716
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5630_6
timestamp 1731220586
transform 1 0 2544 0 1 1716
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5629_6
timestamp 1731220586
transform 1 0 2648 0 1 1716
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5628_6
timestamp 1731220586
transform 1 0 2752 0 -1 1712
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5627_6
timestamp 1731220586
transform 1 0 2616 0 -1 1712
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5626_6
timestamp 1731220586
transform 1 0 2488 0 -1 1712
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5625_6
timestamp 1731220586
transform 1 0 2360 0 -1 1712
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5624_6
timestamp 1731220586
transform 1 0 2240 0 -1 1712
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5623_6
timestamp 1731220586
transform 1 0 2688 0 1 1572
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5622_6
timestamp 1731220586
transform 1 0 2512 0 1 1572
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5621_6
timestamp 1731220586
transform 1 0 2328 0 1 1572
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5620_6
timestamp 1731220586
transform 1 0 2136 0 1 1572
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5619_6
timestamp 1731220586
transform 1 0 2080 0 -1 1572
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5618_6
timestamp 1731220586
transform 1 0 2448 0 -1 1572
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5617_6
timestamp 1731220586
transform 1 0 2272 0 -1 1572
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5616_6
timestamp 1731220586
transform 1 0 2104 0 1 1428
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5615_6
timestamp 1731220586
transform 1 0 2232 0 1 1428
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5614_6
timestamp 1731220586
transform 1 0 2368 0 1 1428
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5613_6
timestamp 1731220586
transform 1 0 2296 0 -1 1424
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5612_6
timestamp 1731220586
transform 1 0 2176 0 -1 1424
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5611_6
timestamp 1731220586
transform 1 0 2208 0 1 1284
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5610_6
timestamp 1731220586
transform 1 0 2088 0 1 1284
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5609_6
timestamp 1731220586
transform 1 0 1968 0 1 1284
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5608_6
timestamp 1731220586
transform 1 0 1880 0 1 1284
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5607_6
timestamp 1731220586
transform 1 0 1880 0 -1 1424
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5606_6
timestamp 1731220586
transform 1 0 1968 0 -1 1424
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5605_6
timestamp 1731220586
transform 1 0 2064 0 -1 1424
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5604_6
timestamp 1731220586
transform 1 0 1976 0 1 1428
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5603_6
timestamp 1731220586
transform 1 0 1880 0 1 1428
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5602_6
timestamp 1731220586
transform 1 0 1720 0 1 1500
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5601_6
timestamp 1731220586
transform 1 0 1576 0 1 1500
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5600_6
timestamp 1731220586
transform 1 0 1448 0 -1 1636
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5599_6
timestamp 1731220586
transform 1 0 1592 0 -1 1636
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5598_6
timestamp 1731220586
transform 1 0 1720 0 -1 1636
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5597_6
timestamp 1731220586
transform 1 0 1680 0 1 1644
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5596_6
timestamp 1731220586
transform 1 0 1696 0 -1 1784
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5595_6
timestamp 1731220586
transform 1 0 1368 0 -1 1784
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5594_6
timestamp 1731220586
transform 1 0 1344 0 1 1796
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5593_6
timestamp 1731220586
transform 1 0 1248 0 1 1796
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5592_6
timestamp 1731220586
transform 1 0 1440 0 1 1796
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5591_6
timestamp 1731220586
transform 1 0 1456 0 -1 1940
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5590_6
timestamp 1731220586
transform 1 0 1144 0 1 1796
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5589_6
timestamp 1731220586
transform 1 0 1040 0 1 1796
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5588_6
timestamp 1731220586
transform 1 0 1208 0 -1 1784
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5587_6
timestamp 1731220586
transform 1 0 1040 0 -1 1784
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5586_6
timestamp 1731220586
transform 1 0 1008 0 1 1644
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5585_6
timestamp 1731220586
transform 1 0 984 0 -1 1636
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5584_6
timestamp 1731220586
transform 1 0 1088 0 1 1500
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5583_6
timestamp 1731220586
transform 1 0 920 0 1 1500
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5582_6
timestamp 1731220586
transform 1 0 864 0 -1 1496
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5581_6
timestamp 1731220586
transform 1 0 984 0 -1 1496
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5580_6
timestamp 1731220586
transform 1 0 1112 0 -1 1496
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5579_6
timestamp 1731220586
transform 1 0 1104 0 1 1352
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5578_6
timestamp 1731220586
transform 1 0 1000 0 1 1352
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5577_6
timestamp 1731220586
transform 1 0 904 0 1 1352
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5576_6
timestamp 1731220586
transform 1 0 800 0 1 1352
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5575_6
timestamp 1731220586
transform 1 0 696 0 -1 1348
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5574_6
timestamp 1731220586
transform 1 0 568 0 1 1352
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5573_6
timestamp 1731220586
transform 1 0 448 0 1 1352
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5572_6
timestamp 1731220586
transform 1 0 688 0 1 1352
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5571_6
timestamp 1731220586
transform 1 0 736 0 -1 1496
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5570_6
timestamp 1731220586
transform 1 0 600 0 -1 1496
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5569_6
timestamp 1731220586
transform 1 0 464 0 -1 1496
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5568_6
timestamp 1731220586
transform 1 0 320 0 -1 1496
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5567_6
timestamp 1731220586
transform 1 0 416 0 1 1500
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5566_6
timestamp 1731220586
transform 1 0 584 0 1 1500
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5565_6
timestamp 1731220586
transform 1 0 752 0 1 1500
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5564_6
timestamp 1731220586
transform 1 0 808 0 -1 1636
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5563_6
timestamp 1731220586
transform 1 0 624 0 -1 1636
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5562_6
timestamp 1731220586
transform 1 0 440 0 -1 1636
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5561_6
timestamp 1731220586
transform 1 0 264 0 -1 1636
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5560_6
timestamp 1731220586
transform 1 0 272 0 1 1644
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5559_6
timestamp 1731220586
transform 1 0 456 0 1 1644
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5558_6
timestamp 1731220586
transform 1 0 640 0 1 1644
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5557_6
timestamp 1731220586
transform 1 0 824 0 1 1644
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5556_6
timestamp 1731220586
transform 1 0 864 0 -1 1784
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5555_6
timestamp 1731220586
transform 1 0 680 0 -1 1784
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5554_6
timestamp 1731220586
transform 1 0 488 0 -1 1784
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5553_6
timestamp 1731220586
transform 1 0 544 0 1 1796
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5552_6
timestamp 1731220586
transform 1 0 680 0 1 1796
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5551_6
timestamp 1731220586
transform 1 0 808 0 1 1796
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5550_6
timestamp 1731220586
transform 1 0 928 0 1 1796
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5549_6
timestamp 1731220586
transform 1 0 1240 0 -1 1940
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5548_6
timestamp 1731220586
transform 1 0 1032 0 -1 1940
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5547_6
timestamp 1731220586
transform 1 0 832 0 -1 1940
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5546_6
timestamp 1731220586
transform 1 0 760 0 1 1944
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5545_6
timestamp 1731220586
transform 1 0 880 0 1 1944
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5544_6
timestamp 1731220586
transform 1 0 1000 0 1 1944
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5543_6
timestamp 1731220586
transform 1 0 1240 0 1 1944
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5542_6
timestamp 1731220586
transform 1 0 1120 0 1 1944
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5541_6
timestamp 1731220586
transform 1 0 1032 0 -1 2084
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5540_6
timestamp 1731220586
transform 1 0 912 0 -1 2084
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5539_6
timestamp 1731220586
transform 1 0 1152 0 -1 2084
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5538_6
timestamp 1731220586
transform 1 0 1272 0 -1 2084
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5537_6
timestamp 1731220586
transform 1 0 1400 0 -1 2084
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5536_6
timestamp 1731220586
transform 1 0 1312 0 1 2088
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5535_6
timestamp 1731220586
transform 1 0 1168 0 1 2088
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5534_6
timestamp 1731220586
transform 1 0 1456 0 1 2088
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5533_6
timestamp 1731220586
transform 1 0 1608 0 1 2088
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5532_6
timestamp 1731220586
transform 1 0 1720 0 -1 2224
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5531_6
timestamp 1731220586
transform 1 0 1568 0 -1 2224
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5530_6
timestamp 1731220586
transform 1 0 1400 0 -1 2224
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5529_6
timestamp 1731220586
transform 1 0 1232 0 -1 2224
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5528_6
timestamp 1731220586
transform 1 0 1720 0 1 2232
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5527_6
timestamp 1731220586
transform 1 0 1584 0 1 2232
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5526_6
timestamp 1731220586
transform 1 0 1448 0 1 2232
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5525_6
timestamp 1731220586
transform 1 0 1304 0 1 2232
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5524_6
timestamp 1731220586
transform 1 0 1160 0 1 2232
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5523_6
timestamp 1731220586
transform 1 0 1576 0 -1 2376
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5522_6
timestamp 1731220586
transform 1 0 1448 0 -1 2376
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5521_6
timestamp 1731220586
transform 1 0 1320 0 -1 2376
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5520_6
timestamp 1731220586
transform 1 0 1200 0 -1 2376
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5519_6
timestamp 1731220586
transform 1 0 1072 0 -1 2376
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5518_6
timestamp 1731220586
transform 1 0 1392 0 1 2388
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5517_6
timestamp 1731220586
transform 1 0 1256 0 1 2388
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5516_6
timestamp 1731220586
transform 1 0 1120 0 1 2388
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5515_6
timestamp 1731220586
transform 1 0 984 0 1 2388
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5514_6
timestamp 1731220586
transform 1 0 1272 0 -1 2524
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5513_6
timestamp 1731220586
transform 1 0 1136 0 -1 2524
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5512_6
timestamp 1731220586
transform 1 0 1000 0 -1 2524
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5511_6
timestamp 1731220586
transform 1 0 864 0 -1 2524
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5510_6
timestamp 1731220586
transform 1 0 912 0 1 2524
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5509_6
timestamp 1731220586
transform 1 0 1032 0 1 2524
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5508_6
timestamp 1731220586
transform 1 0 1160 0 1 2524
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5507_6
timestamp 1731220586
transform 1 0 1304 0 -1 2664
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5506_6
timestamp 1731220586
transform 1 0 1200 0 -1 2664
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5505_6
timestamp 1731220586
transform 1 0 1096 0 -1 2664
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5504_6
timestamp 1731220586
transform 1 0 992 0 -1 2664
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5503_6
timestamp 1731220586
transform 1 0 896 0 -1 2664
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5502_6
timestamp 1731220586
transform 1 0 792 0 -1 2664
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5501_6
timestamp 1731220586
transform 1 0 688 0 -1 2664
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5500_6
timestamp 1731220586
transform 1 0 792 0 1 2524
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5499_6
timestamp 1731220586
transform 1 0 728 0 -1 2524
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5498_6
timestamp 1731220586
transform 1 0 848 0 1 2388
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5497_6
timestamp 1731220586
transform 1 0 944 0 -1 2376
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5496_6
timestamp 1731220586
transform 1 0 848 0 1 2232
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5495_6
timestamp 1731220586
transform 1 0 680 0 1 2232
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5494_6
timestamp 1731220586
transform 1 0 1008 0 1 2232
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5493_6
timestamp 1731220586
transform 1 0 1064 0 -1 2224
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5492_6
timestamp 1731220586
transform 1 0 888 0 -1 2224
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5491_6
timestamp 1731220586
transform 1 0 712 0 -1 2224
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5490_6
timestamp 1731220586
transform 1 0 528 0 -1 2224
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5489_6
timestamp 1731220586
transform 1 0 1024 0 1 2088
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5488_6
timestamp 1731220586
transform 1 0 880 0 1 2088
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5487_6
timestamp 1731220586
transform 1 0 744 0 1 2088
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5486_6
timestamp 1731220586
transform 1 0 608 0 1 2088
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5485_6
timestamp 1731220586
transform 1 0 480 0 1 2088
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5484_6
timestamp 1731220586
transform 1 0 792 0 -1 2084
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5483_6
timestamp 1731220586
transform 1 0 672 0 -1 2084
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5482_6
timestamp 1731220586
transform 1 0 544 0 -1 2084
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5481_6
timestamp 1731220586
transform 1 0 424 0 -1 2084
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5480_6
timestamp 1731220586
transform 1 0 312 0 -1 2084
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5479_6
timestamp 1731220586
transform 1 0 640 0 1 1944
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5478_6
timestamp 1731220586
transform 1 0 520 0 1 1944
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5477_6
timestamp 1731220586
transform 1 0 400 0 1 1944
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5476_6
timestamp 1731220586
transform 1 0 280 0 1 1944
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5475_6
timestamp 1731220586
transform 1 0 168 0 1 1944
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5474_6
timestamp 1731220586
transform 1 0 648 0 -1 1940
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5473_6
timestamp 1731220586
transform 1 0 488 0 -1 1940
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5472_6
timestamp 1731220586
transform 1 0 344 0 -1 1940
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5471_6
timestamp 1731220586
transform 1 0 216 0 -1 1940
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5470_6
timestamp 1731220586
transform 1 0 128 0 -1 1940
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5469_6
timestamp 1731220586
transform 1 0 128 0 1 1796
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5468_6
timestamp 1731220586
transform 1 0 256 0 1 1796
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5467_6
timestamp 1731220586
transform 1 0 400 0 1 1796
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5466_6
timestamp 1731220586
transform 1 0 296 0 -1 1784
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5465_6
timestamp 1731220586
transform 1 0 128 0 -1 1784
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5464_6
timestamp 1731220586
transform 1 0 128 0 1 1644
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5463_6
timestamp 1731220586
transform 1 0 128 0 -1 1636
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5462_6
timestamp 1731220586
transform 1 0 128 0 1 1500
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5461_6
timestamp 1731220586
transform 1 0 256 0 1 1500
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5460_6
timestamp 1731220586
transform 1 0 176 0 -1 1496
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5459_6
timestamp 1731220586
transform 1 0 184 0 1 1352
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5458_6
timestamp 1731220586
transform 1 0 320 0 1 1352
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5457_6
timestamp 1731220586
transform 1 0 224 0 -1 1348
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5456_6
timestamp 1731220586
transform 1 0 376 0 -1 1348
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5455_6
timestamp 1731220586
transform 1 0 536 0 -1 1348
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5454_6
timestamp 1731220586
transform 1 0 864 0 -1 1348
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5453_6
timestamp 1731220586
transform 1 0 824 0 1 1212
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5452_6
timestamp 1731220586
transform 1 0 664 0 1 1212
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5451_6
timestamp 1731220586
transform 1 0 504 0 1 1212
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5450_6
timestamp 1731220586
transform 1 0 344 0 1 1212
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5449_6
timestamp 1731220586
transform 1 0 200 0 1 1212
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5448_6
timestamp 1731220586
transform 1 0 128 0 -1 1204
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5447_6
timestamp 1731220586
transform 1 0 264 0 -1 1204
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5446_6
timestamp 1731220586
transform 1 0 416 0 -1 1204
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5445_6
timestamp 1731220586
transform 1 0 280 0 1 1068
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5444_6
timestamp 1731220586
transform 1 0 128 0 1 1068
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5443_6
timestamp 1731220586
transform 1 0 128 0 -1 1068
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5442_6
timestamp 1731220586
transform 1 0 272 0 1 928
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5441_6
timestamp 1731220586
transform 1 0 128 0 1 928
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5440_6
timestamp 1731220586
transform 1 0 128 0 -1 920
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5439_6
timestamp 1731220586
transform 1 0 264 0 -1 920
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5438_6
timestamp 1731220586
transform 1 0 128 0 1 784
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5437_6
timestamp 1731220586
transform 1 0 128 0 -1 780
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5436_6
timestamp 1731220586
transform 1 0 264 0 -1 780
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5435_6
timestamp 1731220586
transform 1 0 272 0 1 640
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5434_6
timestamp 1731220586
transform 1 0 128 0 1 640
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5433_6
timestamp 1731220586
transform 1 0 128 0 -1 632
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5432_6
timestamp 1731220586
transform 1 0 280 0 -1 632
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5431_6
timestamp 1731220586
transform 1 0 296 0 1 492
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5430_6
timestamp 1731220586
transform 1 0 136 0 1 492
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5429_6
timestamp 1731220586
transform 1 0 152 0 -1 484
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5428_6
timestamp 1731220586
transform 1 0 304 0 -1 484
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5427_6
timestamp 1731220586
transform 1 0 256 0 1 348
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5426_6
timestamp 1731220586
transform 1 0 136 0 1 348
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5425_6
timestamp 1731220586
transform 1 0 392 0 1 348
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5424_6
timestamp 1731220586
transform 1 0 392 0 -1 332
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5423_6
timestamp 1731220586
transform 1 0 304 0 -1 332
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5422_6
timestamp 1731220586
transform 1 0 216 0 -1 332
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5421_6
timestamp 1731220586
transform 1 0 128 0 -1 332
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5420_6
timestamp 1731220586
transform 1 0 128 0 1 192
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5419_6
timestamp 1731220586
transform 1 0 216 0 1 192
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5418_6
timestamp 1731220586
transform 1 0 304 0 1 192
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5417_6
timestamp 1731220586
transform 1 0 392 0 1 192
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5416_6
timestamp 1731220586
transform 1 0 480 0 1 192
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5415_6
timestamp 1731220586
transform 1 0 568 0 1 192
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5414_6
timestamp 1731220586
transform 1 0 656 0 1 192
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5413_6
timestamp 1731220586
transform 1 0 920 0 1 192
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5412_6
timestamp 1731220586
transform 1 0 832 0 1 192
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5411_6
timestamp 1731220586
transform 1 0 744 0 1 192
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5410_6
timestamp 1731220586
transform 1 0 656 0 -1 332
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5409_6
timestamp 1731220586
transform 1 0 568 0 -1 332
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5408_6
timestamp 1731220586
transform 1 0 480 0 -1 332
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5407_6
timestamp 1731220586
transform 1 0 744 0 -1 332
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5406_6
timestamp 1731220586
transform 1 0 832 0 -1 332
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5405_6
timestamp 1731220586
transform 1 0 872 0 1 348
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5404_6
timestamp 1731220586
transform 1 0 696 0 1 348
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5403_6
timestamp 1731220586
transform 1 0 536 0 1 348
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5402_6
timestamp 1731220586
transform 1 0 456 0 -1 484
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5401_6
timestamp 1731220586
transform 1 0 608 0 -1 484
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5400_6
timestamp 1731220586
transform 1 0 752 0 -1 484
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5399_6
timestamp 1731220586
transform 1 0 768 0 1 492
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5398_6
timestamp 1731220586
transform 1 0 616 0 1 492
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5397_6
timestamp 1731220586
transform 1 0 456 0 1 492
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5396_6
timestamp 1731220586
transform 1 0 448 0 -1 632
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5395_6
timestamp 1731220586
transform 1 0 624 0 -1 632
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5394_6
timestamp 1731220586
transform 1 0 792 0 -1 632
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5393_6
timestamp 1731220586
transform 1 0 776 0 1 640
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5392_6
timestamp 1731220586
transform 1 0 608 0 1 640
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5391_6
timestamp 1731220586
transform 1 0 440 0 1 640
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5390_6
timestamp 1731220586
transform 1 0 432 0 -1 780
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5389_6
timestamp 1731220586
transform 1 0 600 0 -1 780
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5388_6
timestamp 1731220586
transform 1 0 768 0 -1 780
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5387_6
timestamp 1731220586
transform 1 0 792 0 1 784
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5386_6
timestamp 1731220586
transform 1 0 624 0 1 784
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5385_6
timestamp 1731220586
transform 1 0 448 0 1 784
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5384_6
timestamp 1731220586
transform 1 0 272 0 1 784
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5383_6
timestamp 1731220586
transform 1 0 432 0 -1 920
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5382_6
timestamp 1731220586
transform 1 0 768 0 -1 920
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5381_6
timestamp 1731220586
transform 1 0 600 0 -1 920
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5380_6
timestamp 1731220586
transform 1 0 448 0 1 928
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5379_6
timestamp 1731220586
transform 1 0 632 0 1 928
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5378_6
timestamp 1731220586
transform 1 0 808 0 1 928
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5377_6
timestamp 1731220586
transform 1 0 728 0 -1 1068
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5376_6
timestamp 1731220586
transform 1 0 576 0 -1 1068
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5375_6
timestamp 1731220586
transform 1 0 424 0 -1 1068
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5374_6
timestamp 1731220586
transform 1 0 264 0 -1 1068
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5373_6
timestamp 1731220586
transform 1 0 464 0 1 1068
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5372_6
timestamp 1731220586
transform 1 0 832 0 1 1068
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5371_6
timestamp 1731220586
transform 1 0 648 0 1 1068
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5370_6
timestamp 1731220586
transform 1 0 568 0 -1 1204
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5369_6
timestamp 1731220586
transform 1 0 720 0 -1 1204
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5368_6
timestamp 1731220586
transform 1 0 880 0 -1 1204
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5367_6
timestamp 1731220586
transform 1 0 1048 0 -1 1204
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5366_6
timestamp 1731220586
transform 1 0 1224 0 -1 1204
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5365_6
timestamp 1731220586
transform 1 0 1192 0 1 1068
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5364_6
timestamp 1731220586
transform 1 0 1016 0 1 1068
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5363_6
timestamp 1731220586
transform 1 0 880 0 -1 1068
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5362_6
timestamp 1731220586
transform 1 0 1040 0 -1 1068
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5361_6
timestamp 1731220586
transform 1 0 1376 0 -1 1068
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5360_6
timestamp 1731220586
transform 1 0 1208 0 -1 1068
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5359_6
timestamp 1731220586
transform 1 0 1152 0 1 928
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5358_6
timestamp 1731220586
transform 1 0 984 0 1 928
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5357_6
timestamp 1731220586
transform 1 0 928 0 -1 920
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5356_6
timestamp 1731220586
transform 1 0 1088 0 -1 920
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5355_6
timestamp 1731220586
transform 1 0 968 0 1 784
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5354_6
timestamp 1731220586
transform 1 0 1144 0 1 784
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5353_6
timestamp 1731220586
transform 1 0 1080 0 -1 780
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5352_6
timestamp 1731220586
transform 1 0 928 0 -1 780
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5351_6
timestamp 1731220586
transform 1 0 944 0 1 640
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5350_6
timestamp 1731220586
transform 1 0 1104 0 1 640
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5349_6
timestamp 1731220586
transform 1 0 1112 0 -1 632
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5348_6
timestamp 1731220586
transform 1 0 960 0 -1 632
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5347_6
timestamp 1731220586
transform 1 0 912 0 1 492
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5346_6
timestamp 1731220586
transform 1 0 1048 0 1 492
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5345_6
timestamp 1731220586
transform 1 0 1000 0 -1 484
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5344_6
timestamp 1731220586
transform 1 0 880 0 -1 484
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5343_6
timestamp 1731220586
transform 1 0 1232 0 1 348
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5342_6
timestamp 1731220586
transform 1 0 1048 0 1 348
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5341_6
timestamp 1731220586
transform 1 0 1008 0 -1 332
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5340_6
timestamp 1731220586
transform 1 0 920 0 -1 332
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5339_6
timestamp 1731220586
transform 1 0 1096 0 -1 332
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5338_6
timestamp 1731220586
transform 1 0 1184 0 -1 332
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5337_6
timestamp 1731220586
transform 1 0 1184 0 1 192
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5336_6
timestamp 1731220586
transform 1 0 1096 0 1 192
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5335_6
timestamp 1731220586
transform 1 0 1008 0 1 192
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5334_6
timestamp 1731220586
transform 1 0 1272 0 1 192
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5333_6
timestamp 1731220586
transform 1 0 1360 0 1 192
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5332_6
timestamp 1731220586
transform 1 0 1448 0 1 192
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5331_6
timestamp 1731220586
transform 1 0 1712 0 1 192
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5330_6
timestamp 1731220586
transform 1 0 1624 0 1 192
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5329_6
timestamp 1731220586
transform 1 0 1536 0 1 192
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5328_6
timestamp 1731220586
transform 1 0 1472 0 -1 332
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5327_6
timestamp 1731220586
transform 1 0 1376 0 -1 332
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5326_6
timestamp 1731220586
transform 1 0 1280 0 -1 332
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5325_6
timestamp 1731220586
transform 1 0 1568 0 -1 332
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5324_6
timestamp 1731220586
transform 1 0 1664 0 -1 332
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5323_6
timestamp 1731220586
transform 1 0 1624 0 1 348
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5322_6
timestamp 1731220586
transform 1 0 1424 0 1 348
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5321_6
timestamp 1731220586
transform 1 0 1336 0 -1 484
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5320_6
timestamp 1731220586
transform 1 0 1232 0 -1 484
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5319_6
timestamp 1731220586
transform 1 0 1120 0 -1 484
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5318_6
timestamp 1731220586
transform 1 0 1520 0 1 492
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5317_6
timestamp 1731220586
transform 1 0 1632 0 1 492
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5316_6
timestamp 1731220586
transform 1 0 1720 0 1 492
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5315_6
timestamp 1731220586
transform 1 0 1880 0 1 536
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5314_6
timestamp 1731220586
transform 1 0 1880 0 -1 676
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5313_6
timestamp 1731220586
transform 1 0 1968 0 -1 676
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5312_6
timestamp 1731220586
transform 1 0 2088 0 -1 676
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5311_6
timestamp 1731220586
transform 1 0 2056 0 1 680
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5310_6
timestamp 1731220586
transform 1 0 1880 0 1 680
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5309_6
timestamp 1731220586
transform 1 0 2064 0 -1 816
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5308_6
timestamp 1731220586
transform 1 0 1880 0 -1 816
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5307_6
timestamp 1731220586
transform 1 0 1880 0 1 824
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5306_6
timestamp 1731220586
transform 1 0 2008 0 1 824
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5305_6
timestamp 1731220586
transform 1 0 2168 0 1 824
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5304_6
timestamp 1731220586
transform 1 0 2064 0 -1 968
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5303_6
timestamp 1731220586
transform 1 0 1880 0 -1 968
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5302_6
timestamp 1731220586
transform 1 0 1904 0 1 972
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5301_6
timestamp 1731220586
transform 1 0 2112 0 1 972
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5300_6
timestamp 1731220586
transform 1 0 2224 0 -1 1120
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5299_6
timestamp 1731220586
transform 1 0 2080 0 -1 1120
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5298_6
timestamp 1731220586
transform 1 0 1936 0 -1 1120
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5297_6
timestamp 1731220586
transform 1 0 2024 0 1 1132
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5296_6
timestamp 1731220586
transform 1 0 2264 0 1 1132
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5295_6
timestamp 1731220586
transform 1 0 2136 0 1 1132
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5294_6
timestamp 1731220586
transform 1 0 2048 0 -1 1272
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5293_6
timestamp 1731220586
transform 1 0 2136 0 -1 1272
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5292_6
timestamp 1731220586
transform 1 0 2232 0 -1 1272
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5291_6
timestamp 1731220586
transform 1 0 2328 0 -1 1272
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5290_6
timestamp 1731220586
transform 1 0 2424 0 -1 1272
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5289_6
timestamp 1731220586
transform 1 0 2400 0 1 1132
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5288_6
timestamp 1731220586
transform 1 0 2544 0 1 1132
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5287_6
timestamp 1731220586
transform 1 0 2528 0 -1 1120
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5286_6
timestamp 1731220586
transform 1 0 2376 0 -1 1120
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5285_6
timestamp 1731220586
transform 1 0 2312 0 1 972
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5284_6
timestamp 1731220586
transform 1 0 2504 0 1 972
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5283_6
timestamp 1731220586
transform 1 0 2624 0 -1 968
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5282_6
timestamp 1731220586
transform 1 0 2448 0 -1 968
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5281_6
timestamp 1731220586
transform 1 0 2256 0 -1 968
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5280_6
timestamp 1731220586
transform 1 0 2336 0 1 824
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5279_6
timestamp 1731220586
transform 1 0 2504 0 1 824
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5278_6
timestamp 1731220586
transform 1 0 2672 0 1 824
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5277_6
timestamp 1731220586
transform 1 0 2616 0 -1 816
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5276_6
timestamp 1731220586
transform 1 0 2440 0 -1 816
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5275_6
timestamp 1731220586
transform 1 0 2256 0 -1 816
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5274_6
timestamp 1731220586
transform 1 0 2248 0 1 680
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5273_6
timestamp 1731220586
transform 1 0 2432 0 1 680
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5272_6
timestamp 1731220586
transform 1 0 2472 0 -1 676
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5271_6
timestamp 1731220586
transform 1 0 2344 0 -1 676
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5270_6
timestamp 1731220586
transform 1 0 2216 0 -1 676
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5269_6
timestamp 1731220586
transform 1 0 2200 0 1 536
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5268_6
timestamp 1731220586
transform 1 0 2032 0 1 536
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5267_6
timestamp 1731220586
transform 1 0 2368 0 -1 528
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5266_6
timestamp 1731220586
transform 1 0 2272 0 -1 528
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5265_6
timestamp 1731220586
transform 1 0 2184 0 -1 528
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5264_6
timestamp 1731220586
transform 1 0 2024 0 1 384
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5263_6
timestamp 1731220586
transform 1 0 2192 0 1 384
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5262_6
timestamp 1731220586
transform 1 0 2256 0 -1 384
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5261_6
timestamp 1731220586
transform 1 0 2376 0 -1 384
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5260_6
timestamp 1731220586
transform 1 0 2512 0 -1 384
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5259_6
timestamp 1731220586
transform 1 0 2456 0 1 248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5258_6
timestamp 1731220586
transform 1 0 2344 0 1 248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5257_6
timestamp 1731220586
transform 1 0 2568 0 1 248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5256_6
timestamp 1731220586
transform 1 0 2672 0 -1 248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5255_6
timestamp 1731220586
transform 1 0 2528 0 -1 248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5254_6
timestamp 1731220586
transform 1 0 2392 0 -1 248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5253_6
timestamp 1731220586
transform 1 0 2256 0 -1 248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5252_6
timestamp 1731220586
transform 1 0 2144 0 -1 248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5251_6
timestamp 1731220586
transform 1 0 2056 0 -1 248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5250_6
timestamp 1731220586
transform 1 0 1968 0 -1 248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5249_6
timestamp 1731220586
transform 1 0 1880 0 -1 248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5248_6
timestamp 1731220586
transform 1 0 2232 0 1 248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5247_6
timestamp 1731220586
transform 1 0 2144 0 1 248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5246_6
timestamp 1731220586
transform 1 0 2056 0 1 248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5245_6
timestamp 1731220586
transform 1 0 1968 0 1 248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5244_6
timestamp 1731220586
transform 1 0 1880 0 1 248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5243_6
timestamp 1731220586
transform 1 0 2144 0 -1 384
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5242_6
timestamp 1731220586
transform 1 0 2056 0 -1 384
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5241_6
timestamp 1731220586
transform 1 0 1968 0 -1 384
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5240_6
timestamp 1731220586
transform 1 0 1880 0 -1 384
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5239_6
timestamp 1731220586
transform 1 0 1880 0 1 384
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5238_6
timestamp 1731220586
transform 1 0 1720 0 -1 484
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5237_6
timestamp 1731220586
transform 1 0 1632 0 -1 484
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5236_6
timestamp 1731220586
transform 1 0 1536 0 -1 484
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5235_6
timestamp 1731220586
transform 1 0 1432 0 -1 484
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5234_6
timestamp 1731220586
transform 1 0 1408 0 1 492
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5233_6
timestamp 1731220586
transform 1 0 1296 0 1 492
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5232_6
timestamp 1731220586
transform 1 0 1176 0 1 492
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5231_6
timestamp 1731220586
transform 1 0 1704 0 -1 632
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5230_6
timestamp 1731220586
transform 1 0 1552 0 -1 632
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5229_6
timestamp 1731220586
transform 1 0 1408 0 -1 632
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5228_6
timestamp 1731220586
transform 1 0 1264 0 -1 632
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5227_6
timestamp 1731220586
transform 1 0 1264 0 1 640
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5226_6
timestamp 1731220586
transform 1 0 1424 0 1 640
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5225_6
timestamp 1731220586
transform 1 0 1584 0 1 640
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5224_6
timestamp 1731220586
transform 1 0 1544 0 -1 780
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5223_6
timestamp 1731220586
transform 1 0 1384 0 -1 780
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5222_6
timestamp 1731220586
transform 1 0 1232 0 -1 780
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5221_6
timestamp 1731220586
transform 1 0 1320 0 1 784
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5220_6
timestamp 1731220586
transform 1 0 1496 0 1 784
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5219_6
timestamp 1731220586
transform 1 0 1392 0 -1 920
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5218_6
timestamp 1731220586
transform 1 0 1240 0 -1 920
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5217_6
timestamp 1731220586
transform 1 0 1544 0 -1 920
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5216_6
timestamp 1731220586
transform 1 0 1472 0 1 928
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5215_6
timestamp 1731220586
transform 1 0 1312 0 1 928
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5214_6
timestamp 1731220586
transform 1 0 1640 0 1 928
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5213_6
timestamp 1731220586
transform 1 0 1552 0 -1 1068
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5212_6
timestamp 1731220586
transform 1 0 1720 0 -1 1068
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5211_6
timestamp 1731220586
transform 1 0 1720 0 1 1068
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5210_6
timestamp 1731220586
transform 1 0 1560 0 1 1068
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5209_6
timestamp 1731220586
transform 1 0 1376 0 1 1068
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5208_6
timestamp 1731220586
transform 1 0 1408 0 -1 1204
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5207_6
timestamp 1731220586
transform 1 0 1592 0 -1 1204
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5206_6
timestamp 1731220586
transform 1 0 1576 0 1 1212
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5205_6
timestamp 1731220586
transform 1 0 1424 0 1 1212
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5204_6
timestamp 1731220586
transform 1 0 1280 0 1 1212
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5203_6
timestamp 1731220586
transform 1 0 1136 0 1 1212
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5202_6
timestamp 1731220586
transform 1 0 984 0 1 1212
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5201_6
timestamp 1731220586
transform 1 0 1032 0 -1 1348
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5200_6
timestamp 1731220586
transform 1 0 1200 0 -1 1348
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5199_6
timestamp 1731220586
transform 1 0 1368 0 -1 1348
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5198_6
timestamp 1731220586
transform 1 0 1312 0 1 1352
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5197_6
timestamp 1731220586
transform 1 0 1208 0 1 1352
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5196_6
timestamp 1731220586
transform 1 0 1240 0 -1 1496
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5195_6
timestamp 1731220586
transform 1 0 1368 0 -1 1496
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5194_6
timestamp 1731220586
transform 1 0 1408 0 1 1500
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5193_6
timestamp 1731220586
transform 1 0 1248 0 1 1500
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5192_6
timestamp 1731220586
transform 1 0 1296 0 -1 1636
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5191_6
timestamp 1731220586
transform 1 0 1144 0 -1 1636
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5190_6
timestamp 1731220586
transform 1 0 1176 0 1 1644
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5189_6
timestamp 1731220586
transform 1 0 1344 0 1 1644
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5188_6
timestamp 1731220586
transform 1 0 1512 0 1 1644
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5187_6
timestamp 1731220586
transform 1 0 1528 0 -1 1784
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5186_6
timestamp 1731220586
transform 1 0 1536 0 1 1796
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5185_6
timestamp 1731220586
transform 1 0 1632 0 1 1796
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5184_6
timestamp 1731220586
transform 1 0 1720 0 1 1796
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5183_6
timestamp 1731220586
transform 1 0 1880 0 1 1864
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5182_6
timestamp 1731220586
transform 1 0 2104 0 1 1864
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5181_6
timestamp 1731220586
transform 1 0 1976 0 1 1864
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5180_6
timestamp 1731220586
transform 1 0 1880 0 -1 2008
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5179_6
timestamp 1731220586
transform 1 0 2024 0 -1 2008
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5178_6
timestamp 1731220586
transform 1 0 2192 0 -1 2008
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5177_6
timestamp 1731220586
transform 1 0 2128 0 1 2008
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5176_6
timestamp 1731220586
transform 1 0 1968 0 1 2008
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5175_6
timestamp 1731220586
transform 1 0 2016 0 -1 2148
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5174_6
timestamp 1731220586
transform 1 0 2160 0 -1 2148
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5173_6
timestamp 1731220586
transform 1 0 2320 0 1 2156
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5172_6
timestamp 1731220586
transform 1 0 2152 0 1 2156
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5171_6
timestamp 1731220586
transform 1 0 1992 0 1 2156
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5170_6
timestamp 1731220586
transform 1 0 1968 0 -1 2292
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5169_6
timestamp 1731220586
transform 1 0 2136 0 -1 2292
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5168_6
timestamp 1731220586
transform 1 0 2072 0 1 2296
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5167_6
timestamp 1731220586
transform 1 0 1912 0 1 2296
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5166_6
timestamp 1731220586
transform 1 0 1880 0 -1 2436
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5165_6
timestamp 1731220586
transform 1 0 2008 0 -1 2436
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5164_6
timestamp 1731220586
transform 1 0 2016 0 1 2436
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5163_6
timestamp 1731220586
transform 1 0 1880 0 1 2436
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5162_6
timestamp 1731220586
transform 1 0 1880 0 -1 2576
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5161_6
timestamp 1731220586
transform 1 0 1984 0 -1 2576
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5160_6
timestamp 1731220586
transform 1 0 1984 0 1 2580
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5159_6
timestamp 1731220586
transform 1 0 1880 0 1 2580
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5158_6
timestamp 1731220586
transform 1 0 1880 0 -1 2724
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5157_6
timestamp 1731220586
transform 1 0 2040 0 -1 2724
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5156_6
timestamp 1731220586
transform 1 0 1880 0 1 2728
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5155_6
timestamp 1731220586
transform 1 0 2048 0 1 2728
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5154_6
timestamp 1731220586
transform 1 0 2016 0 -1 2864
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5153_6
timestamp 1731220586
transform 1 0 1880 0 -1 2864
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5152_6
timestamp 1731220586
transform 1 0 1880 0 1 2864
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5151_6
timestamp 1731220586
transform 1 0 1720 0 -1 2960
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5150_6
timestamp 1731220586
transform 1 0 1632 0 -1 2960
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5149_6
timestamp 1731220586
transform 1 0 1720 0 1 2960
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5148_6
timestamp 1731220586
transform 1 0 1688 0 -1 3100
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5147_6
timestamp 1731220586
transform 1 0 1552 0 -1 3100
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5146_6
timestamp 1731220586
transform 1 0 1448 0 1 3108
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5145_6
timestamp 1731220586
transform 1 0 1624 0 1 3108
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5144_6
timestamp 1731220586
transform 1 0 1568 0 -1 3252
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5143_6
timestamp 1731220586
transform 1 0 1408 0 -1 3252
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5142_6
timestamp 1731220586
transform 1 0 1336 0 1 3256
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5141_6
timestamp 1731220586
transform 1 0 1528 0 1 3256
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5140_6
timestamp 1731220586
transform 1 0 1520 0 -1 3396
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5139_6
timestamp 1731220586
transform 1 0 1360 0 -1 3396
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5138_6
timestamp 1731220586
transform 1 0 1200 0 -1 3396
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5137_6
timestamp 1731220586
transform 1 0 1168 0 1 3396
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5136_6
timestamp 1731220586
transform 1 0 1312 0 1 3396
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5135_6
timestamp 1731220586
transform 1 0 1464 0 1 3396
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5134_6
timestamp 1731220586
transform 1 0 1568 0 -1 3532
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5133_6
timestamp 1731220586
transform 1 0 1464 0 -1 3532
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5132_6
timestamp 1731220586
transform 1 0 1360 0 -1 3532
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5131_6
timestamp 1731220586
transform 1 0 1264 0 -1 3532
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5130_6
timestamp 1731220586
transform 1 0 1168 0 -1 3532
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5129_6
timestamp 1731220586
transform 1 0 1072 0 -1 3532
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5128_6
timestamp 1731220586
transform 1 0 968 0 -1 3532
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5127_6
timestamp 1731220586
transform 1 0 856 0 -1 3532
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5126_6
timestamp 1731220586
transform 1 0 736 0 -1 3532
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5125_6
timestamp 1731220586
transform 1 0 880 0 1 3396
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5124_6
timestamp 1731220586
transform 1 0 1024 0 1 3396
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5123_6
timestamp 1731220586
transform 1 0 1040 0 -1 3396
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5122_6
timestamp 1731220586
transform 1 0 880 0 -1 3396
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5121_6
timestamp 1731220586
transform 1 0 968 0 1 3256
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5120_6
timestamp 1731220586
transform 1 0 1152 0 1 3256
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5119_6
timestamp 1731220586
transform 1 0 1088 0 -1 3252
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5118_6
timestamp 1731220586
transform 1 0 928 0 -1 3252
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5117_6
timestamp 1731220586
transform 1 0 1248 0 -1 3252
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5116_6
timestamp 1731220586
transform 1 0 1120 0 1 3108
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5115_6
timestamp 1731220586
transform 1 0 1280 0 1 3108
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5114_6
timestamp 1731220586
transform 1 0 1416 0 -1 3100
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5113_6
timestamp 1731220586
transform 1 0 1280 0 -1 3100
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5112_6
timestamp 1731220586
transform 1 0 1152 0 -1 3100
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5111_6
timestamp 1731220586
transform 1 0 1224 0 1 2960
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5110_6
timestamp 1731220586
transform 1 0 1352 0 1 2960
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5109_6
timestamp 1731220586
transform 1 0 1480 0 1 2960
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5108_6
timestamp 1731220586
transform 1 0 1608 0 1 2960
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5107_6
timestamp 1731220586
transform 1 0 1520 0 -1 2960
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5106_6
timestamp 1731220586
transform 1 0 1408 0 -1 2960
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5105_6
timestamp 1731220586
transform 1 0 1296 0 -1 2960
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5104_6
timestamp 1731220586
transform 1 0 1176 0 -1 2960
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5103_6
timestamp 1731220586
transform 1 0 1048 0 -1 2960
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5102_6
timestamp 1731220586
transform 1 0 1536 0 1 2820
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5101_6
timestamp 1731220586
transform 1 0 1400 0 1 2820
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5100_6
timestamp 1731220586
transform 1 0 1264 0 1 2820
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_599_6
timestamp 1731220586
transform 1 0 1128 0 1 2820
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_598_6
timestamp 1731220586
transform 1 0 992 0 1 2820
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_597_6
timestamp 1731220586
transform 1 0 1336 0 -1 2812
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_596_6
timestamp 1731220586
transform 1 0 1200 0 -1 2812
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_595_6
timestamp 1731220586
transform 1 0 1072 0 -1 2812
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_594_6
timestamp 1731220586
transform 1 0 944 0 -1 2812
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_593_6
timestamp 1731220586
transform 1 0 816 0 -1 2812
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_592_6
timestamp 1731220586
transform 1 0 1032 0 1 2668
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_591_6
timestamp 1731220586
transform 1 0 888 0 1 2668
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_590_6
timestamp 1731220586
transform 1 0 744 0 1 2668
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_589_6
timestamp 1731220586
transform 1 0 576 0 -1 2664
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_588_6
timestamp 1731220586
transform 1 0 536 0 1 2524
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_587_6
timestamp 1731220586
transform 1 0 664 0 1 2524
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_586_6
timestamp 1731220586
transform 1 0 584 0 -1 2524
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_585_6
timestamp 1731220586
transform 1 0 576 0 1 2388
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_584_6
timestamp 1731220586
transform 1 0 712 0 1 2388
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_583_6
timestamp 1731220586
transform 1 0 808 0 -1 2376
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_582_6
timestamp 1731220586
transform 1 0 680 0 -1 2376
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_581_6
timestamp 1731220586
transform 1 0 552 0 -1 2376
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_580_6
timestamp 1731220586
transform 1 0 432 0 -1 2376
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_579_6
timestamp 1731220586
transform 1 0 328 0 -1 2376
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_578_6
timestamp 1731220586
transform 1 0 240 0 -1 2376
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_577_6
timestamp 1731220586
transform 1 0 152 0 -1 2376
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_576_6
timestamp 1731220586
transform 1 0 176 0 1 2388
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_575_6
timestamp 1731220586
transform 1 0 304 0 1 2388
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_574_6
timestamp 1731220586
transform 1 0 440 0 1 2388
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_573_6
timestamp 1731220586
transform 1 0 432 0 -1 2524
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_572_6
timestamp 1731220586
transform 1 0 272 0 -1 2524
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_571_6
timestamp 1731220586
transform 1 0 128 0 -1 2524
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_570_6
timestamp 1731220586
transform 1 0 128 0 1 2524
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_569_6
timestamp 1731220586
transform 1 0 256 0 1 2524
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_568_6
timestamp 1731220586
transform 1 0 400 0 1 2524
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_567_6
timestamp 1731220586
transform 1 0 464 0 -1 2664
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_566_6
timestamp 1731220586
transform 1 0 344 0 -1 2664
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_565_6
timestamp 1731220586
transform 1 0 224 0 -1 2664
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_564_6
timestamp 1731220586
transform 1 0 128 0 -1 2664
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_563_6
timestamp 1731220586
transform 1 0 128 0 1 2668
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_562_6
timestamp 1731220586
transform 1 0 216 0 1 2668
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_561_6
timestamp 1731220586
transform 1 0 600 0 1 2668
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_560_6
timestamp 1731220586
transform 1 0 464 0 1 2668
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_559_6
timestamp 1731220586
transform 1 0 336 0 1 2668
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_558_6
timestamp 1731220586
transform 1 0 288 0 -1 2812
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_557_6
timestamp 1731220586
transform 1 0 160 0 -1 2812
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_556_6
timestamp 1731220586
transform 1 0 688 0 -1 2812
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_555_6
timestamp 1731220586
transform 1 0 552 0 -1 2812
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_554_6
timestamp 1731220586
transform 1 0 416 0 -1 2812
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_553_6
timestamp 1731220586
transform 1 0 312 0 1 2820
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_552_6
timestamp 1731220586
transform 1 0 440 0 1 2820
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_551_6
timestamp 1731220586
transform 1 0 576 0 1 2820
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_550_6
timestamp 1731220586
transform 1 0 712 0 1 2820
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_549_6
timestamp 1731220586
transform 1 0 856 0 1 2820
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_548_6
timestamp 1731220586
transform 1 0 912 0 -1 2960
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_547_6
timestamp 1731220586
transform 1 0 776 0 -1 2960
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_546_6
timestamp 1731220586
transform 1 0 632 0 -1 2960
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_545_6
timestamp 1731220586
transform 1 0 488 0 -1 2960
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_544_6
timestamp 1731220586
transform 1 0 560 0 1 2960
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_543_6
timestamp 1731220586
transform 1 0 688 0 1 2960
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_542_6
timestamp 1731220586
transform 1 0 816 0 1 2960
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_541_6
timestamp 1731220586
transform 1 0 952 0 1 2960
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_540_6
timestamp 1731220586
transform 1 0 1088 0 1 2960
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_539_6
timestamp 1731220586
transform 1 0 1024 0 -1 3100
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_538_6
timestamp 1731220586
transform 1 0 896 0 -1 3100
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_537_6
timestamp 1731220586
transform 1 0 776 0 -1 3100
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_536_6
timestamp 1731220586
transform 1 0 656 0 -1 3100
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_535_6
timestamp 1731220586
transform 1 0 544 0 -1 3100
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_534_6
timestamp 1731220586
transform 1 0 960 0 1 3108
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_533_6
timestamp 1731220586
transform 1 0 808 0 1 3108
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_532_6
timestamp 1731220586
transform 1 0 672 0 1 3108
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_531_6
timestamp 1731220586
transform 1 0 544 0 1 3108
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_530_6
timestamp 1731220586
transform 1 0 432 0 1 3108
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_529_6
timestamp 1731220586
transform 1 0 776 0 -1 3252
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_528_6
timestamp 1731220586
transform 1 0 632 0 -1 3252
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_527_6
timestamp 1731220586
transform 1 0 496 0 -1 3252
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_526_6
timestamp 1731220586
transform 1 0 360 0 -1 3252
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_525_6
timestamp 1731220586
transform 1 0 792 0 1 3256
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_524_6
timestamp 1731220586
transform 1 0 624 0 1 3256
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_523_6
timestamp 1731220586
transform 1 0 464 0 1 3256
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_522_6
timestamp 1731220586
transform 1 0 320 0 1 3256
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_521_6
timestamp 1731220586
transform 1 0 192 0 1 3256
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_520_6
timestamp 1731220586
transform 1 0 720 0 -1 3396
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_519_6
timestamp 1731220586
transform 1 0 560 0 -1 3396
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_518_6
timestamp 1731220586
transform 1 0 400 0 -1 3396
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_517_6
timestamp 1731220586
transform 1 0 256 0 -1 3396
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_516_6
timestamp 1731220586
transform 1 0 128 0 -1 3396
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_515_6
timestamp 1731220586
transform 1 0 160 0 1 3396
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_514_6
timestamp 1731220586
transform 1 0 288 0 1 3396
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_513_6
timestamp 1731220586
transform 1 0 432 0 1 3396
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_512_6
timestamp 1731220586
transform 1 0 576 0 1 3396
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_511_6
timestamp 1731220586
transform 1 0 728 0 1 3396
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_510_6
timestamp 1731220586
transform 1 0 616 0 -1 3532
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_59_6
timestamp 1731220586
transform 1 0 496 0 -1 3532
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_58_6
timestamp 1731220586
transform 1 0 368 0 -1 3532
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_57_6
timestamp 1731220586
transform 1 0 240 0 -1 3532
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_56_6
timestamp 1731220586
transform 1 0 480 0 1 3532
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_55_6
timestamp 1731220586
transform 1 0 392 0 1 3532
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_54_6
timestamp 1731220586
transform 1 0 304 0 1 3532
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_53_6
timestamp 1731220586
transform 1 0 216 0 1 3532
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_52_6
timestamp 1731220586
transform 1 0 128 0 1 3532
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_51_6
timestamp 1731220586
transform 1 0 216 0 -1 3668
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_50_6
timestamp 1731220586
transform 1 0 128 0 -1 3668
box 8 4 80 64
<< end >>
