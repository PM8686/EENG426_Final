magic
tech TSMC180
timestamp 1734143631
<< ndiffusion >>
rect 18 31 24 32
rect 18 29 20 31
rect 22 29 24 31
rect 18 22 24 29
rect 26 22 32 32
rect 34 27 40 32
rect 42 31 48 32
rect 42 29 45 31
rect 47 29 48 31
rect 42 27 48 29
rect 34 25 38 27
rect 34 23 35 25
rect 37 23 38 25
rect 34 22 38 23
<< ndcontact >>
rect 20 29 22 31
rect 45 29 47 31
rect 35 23 37 25
<< ntransistor >>
rect 24 22 26 32
rect 32 22 34 32
rect 40 27 42 32
<< pdiffusion >>
rect 18 55 24 56
rect 18 53 19 55
rect 21 53 24 55
rect 18 48 24 53
rect 26 51 32 56
rect 26 49 27 51
rect 29 49 32 51
rect 26 48 32 49
rect 34 55 40 56
rect 34 53 35 55
rect 37 53 40 55
rect 34 48 40 53
rect 42 51 48 56
rect 42 49 45 51
rect 47 49 48 51
rect 42 48 48 49
<< pdcontact >>
rect 19 53 21 55
rect 27 49 29 51
rect 35 53 37 55
rect 45 49 47 51
<< ptransistor >>
rect 24 48 26 56
rect 32 48 34 56
rect 40 48 42 56
<< polysilicon >>
rect 30 63 34 64
rect 30 61 31 63
rect 33 61 34 63
rect 30 60 34 61
rect 24 56 26 59
rect 32 56 34 60
rect 40 56 42 59
rect 24 32 26 48
rect 32 32 34 48
rect 40 41 42 48
rect 40 40 55 41
rect 40 39 52 40
rect 40 32 42 39
rect 51 38 52 39
rect 54 38 55 40
rect 51 37 55 38
rect 40 24 42 27
rect 24 20 26 22
rect 18 19 26 20
rect 32 19 34 22
rect 18 17 19 19
rect 21 18 26 19
rect 21 17 22 18
rect 18 16 22 17
<< polycontact >>
rect 31 61 33 63
rect 52 38 54 40
rect 19 17 21 19
<< m1 >>
rect 18 67 33 70
rect 30 64 33 67
rect 45 67 57 70
rect 30 63 34 64
rect 30 61 31 63
rect 33 61 34 63
rect 30 60 34 61
rect 18 56 23 57
rect 18 53 19 56
rect 22 53 23 56
rect 18 52 23 53
rect 33 56 38 57
rect 33 53 34 56
rect 37 53 38 56
rect 33 52 38 53
rect 45 52 48 67
rect 26 51 30 52
rect 26 49 27 51
rect 29 49 30 51
rect 26 48 30 49
rect 44 51 48 52
rect 44 49 45 51
rect 47 49 48 51
rect 44 48 48 49
rect 26 42 29 48
rect 18 41 23 42
rect 18 38 19 41
rect 22 38 23 41
rect 18 37 23 38
rect 26 41 31 42
rect 26 38 27 41
rect 30 38 31 41
rect 26 37 31 38
rect 20 32 23 37
rect 45 32 48 48
rect 51 41 56 42
rect 51 38 52 41
rect 55 38 56 41
rect 51 37 56 38
rect 19 31 23 32
rect 19 29 20 31
rect 22 29 23 31
rect 19 28 23 29
rect 44 31 48 32
rect 44 29 45 31
rect 47 29 48 31
rect 44 28 48 29
rect 33 25 38 26
rect 33 22 34 25
rect 37 22 38 25
rect 33 21 38 22
rect 18 19 22 20
rect 18 17 19 19
rect 21 17 22 19
rect 18 16 22 17
rect 18 11 21 16
<< m2c >>
rect 19 55 22 56
rect 19 53 21 55
rect 21 53 22 55
rect 34 55 37 56
rect 34 53 35 55
rect 35 53 37 55
rect 19 38 22 41
rect 27 38 30 41
rect 52 40 55 41
rect 52 38 54 40
rect 54 38 55 40
rect 34 23 35 25
rect 35 23 37 25
rect 34 22 37 23
<< m2 >>
rect 7 56 38 57
rect 7 53 19 56
rect 22 53 34 56
rect 37 53 38 56
rect 7 52 38 53
rect 18 41 56 42
rect 18 38 19 41
rect 22 38 27 41
rect 30 38 52 41
rect 55 38 56 41
rect 18 37 56 38
rect 33 25 38 26
rect 33 22 34 25
rect 37 22 38 25
rect 33 10 38 22
<< labels >>
rlabel m1 s 33 61 34 63 6 A
port 1 nsew signal input
rlabel m1 s 31 61 33 63 6 A
port 1 nsew signal input
rlabel m1 s 30 60 34 61 6 A
port 1 nsew signal input
rlabel m1 s 30 61 31 63 6 A
port 1 nsew signal input
rlabel m1 s 30 63 34 64 6 A
port 1 nsew signal input
rlabel m1 s 30 64 33 67 6 A
port 1 nsew signal input
rlabel m1 s 18 67 33 70 6 A
port 1 nsew signal input
rlabel m1 s 21 17 22 19 6 B
port 2 nsew signal input
rlabel m1 s 19 17 21 19 6 B
port 2 nsew signal input
rlabel m1 s 18 11 21 16 6 B
port 2 nsew signal input
rlabel m1 s 18 16 22 17 6 B
port 2 nsew signal input
rlabel m1 s 18 17 19 19 6 B
port 2 nsew signal input
rlabel m1 s 18 19 22 20 6 B
port 2 nsew signal input
rlabel m1 s 47 49 48 51 6 Y
port 3 nsew signal output
rlabel m1 s 47 29 48 31 6 Y
port 3 nsew signal output
rlabel m1 s 45 49 47 51 6 Y
port 3 nsew signal output
rlabel m1 s 45 29 47 31 6 Y
port 3 nsew signal output
rlabel m1 s 45 32 48 48 6 Y
port 3 nsew signal output
rlabel m1 s 44 49 45 51 6 Y
port 3 nsew signal output
rlabel m1 s 44 51 48 52 6 Y
port 3 nsew signal output
rlabel m1 s 45 52 48 67 6 Y
port 3 nsew signal output
rlabel m1 s 45 67 57 70 6 Y
port 3 nsew signal output
rlabel m1 s 44 29 45 31 6 Y
port 3 nsew signal output
rlabel m1 s 44 31 48 32 6 Y
port 3 nsew signal output
rlabel m1 s 44 28 48 29 6 Y
port 3 nsew signal output
rlabel m1 s 44 48 48 49 6 Y
port 3 nsew signal output
rlabel m2 s 37 53 38 56 6 Vdd
port 4 nsew power input
rlabel m2 s 35 53 37 55 6 Vdd
port 4 nsew power input
rlabel m2 s 34 53 35 55 6 Vdd
port 4 nsew power input
rlabel m2 s 34 55 37 56 6 Vdd
port 4 nsew power input
rlabel m2 s 22 53 34 56 6 Vdd
port 4 nsew power input
rlabel m2 s 21 53 22 55 6 Vdd
port 4 nsew power input
rlabel m2 s 19 53 21 55 6 Vdd
port 4 nsew power input
rlabel m2 s 19 55 22 56 6 Vdd
port 4 nsew power input
rlabel m2 s 7 52 38 53 6 Vdd
port 4 nsew power input
rlabel m2 s 7 53 19 56 6 Vdd
port 4 nsew power input
rlabel m2 s 7 56 38 57 6 Vdd
port 4 nsew power input
rlabel m2c s 35 53 37 55 6 Vdd
port 4 nsew power input
rlabel m2c s 34 53 35 55 6 Vdd
port 4 nsew power input
rlabel m2c s 34 55 37 56 6 Vdd
port 4 nsew power input
rlabel m2c s 21 53 22 55 6 Vdd
port 4 nsew power input
rlabel m2c s 19 53 21 55 6 Vdd
port 4 nsew power input
rlabel m2c s 19 55 22 56 6 Vdd
port 4 nsew power input
rlabel m1 s 37 53 38 56 6 Vdd
port 4 nsew power input
rlabel m1 s 35 53 37 55 6 Vdd
port 4 nsew power input
rlabel m1 s 34 53 35 55 6 Vdd
port 4 nsew power input
rlabel m1 s 34 55 37 56 6 Vdd
port 4 nsew power input
rlabel m1 s 33 52 38 53 6 Vdd
port 4 nsew power input
rlabel m1 s 33 53 34 56 6 Vdd
port 4 nsew power input
rlabel m1 s 33 56 38 57 6 Vdd
port 4 nsew power input
rlabel m1 s 22 53 23 56 6 Vdd
port 4 nsew power input
rlabel m1 s 21 53 22 55 6 Vdd
port 4 nsew power input
rlabel m1 s 19 53 21 55 6 Vdd
port 4 nsew power input
rlabel m1 s 19 55 22 56 6 Vdd
port 4 nsew power input
rlabel m1 s 18 52 23 53 6 Vdd
port 4 nsew power input
rlabel m1 s 18 53 19 56 6 Vdd
port 4 nsew power input
rlabel m1 s 18 56 23 57 6 Vdd
port 4 nsew power input
rlabel m2 s 37 22 38 25 6 GND
port 5 nsew ground input
rlabel m2 s 35 23 37 25 6 GND
port 5 nsew ground input
rlabel m2 s 34 22 37 23 6 GND
port 5 nsew ground input
rlabel m2 s 34 23 35 25 6 GND
port 5 nsew ground input
rlabel m2 s 33 10 38 22 6 GND
port 5 nsew ground input
rlabel m2 s 33 22 34 25 6 GND
port 5 nsew ground input
rlabel m2 s 33 25 38 26 6 GND
port 5 nsew ground input
rlabel m2c s 35 23 37 25 6 GND
port 5 nsew ground input
rlabel m2c s 34 22 37 23 6 GND
port 5 nsew ground input
rlabel m2c s 34 23 35 25 6 GND
port 5 nsew ground input
rlabel m1 s 37 22 38 25 6 GND
port 5 nsew ground input
rlabel m1 s 35 23 37 25 6 GND
port 5 nsew ground input
rlabel m1 s 34 22 37 23 6 GND
port 5 nsew ground input
rlabel m1 s 34 23 35 25 6 GND
port 5 nsew ground input
rlabel m1 s 33 21 38 22 6 GND
port 5 nsew ground input
rlabel m1 s 33 22 34 25 6 GND
port 5 nsew ground input
rlabel m1 s 33 25 38 26 6 GND
port 5 nsew ground input
rlabel space 0 0 60 80 1 prboundary
rlabel polysilicon 41 25 41 25 3 _Y
rlabel ndiffusion 38 24 38 24 3 GND
rlabel ndiffusion 43 28 43 28 3 Y
rlabel ndiffusion 43 30 43 30 3 Y
rlabel ndiffusion 43 32 43 32 3 Y
rlabel pdiffusion 43 49 43 49 3 Y
rlabel pdiffusion 43 50 43 50 3 Y
rlabel pdiffusion 43 52 43 52 3 Y
rlabel polysilicon 41 57 41 57 3 _Y
rlabel ntransistor 41 28 41 28 3 _Y
rlabel polysilicon 41 33 41 33 3 _Y
rlabel polysilicon 41 40 41 40 3 _Y
rlabel polysilicon 41 41 41 41 3 _Y
rlabel polysilicon 41 42 41 42 3 _Y
rlabel ptransistor 41 49 41 49 3 _Y
rlabel ndiffusion 35 26 35 26 3 GND
rlabel ndiffusion 35 28 35 28 3 GND
rlabel pdiffusion 35 49 35 49 3 Vdd
rlabel polysilicon 33 57 33 57 3 A
rlabel ntransistor 33 23 33 23 3 A
rlabel polysilicon 33 33 33 33 3 A
rlabel ptransistor 33 49 33 49 3 A
rlabel polysilicon 22 19 22 19 3 B
rlabel polysilicon 33 20 33 20 3 A
rlabel polysilicon 25 21 25 21 3 B
rlabel ntransistor 25 23 25 23 3 B
rlabel polysilicon 25 33 25 33 3 B
rlabel ptransistor 25 49 25 49 3 B
rlabel polysilicon 25 57 25 57 3 B
rlabel ndiffusion 19 23 19 23 3 _Y
rlabel ndiffusion 19 30 19 30 3 _Y
rlabel ndiffusion 19 32 19 32 3 _Y
rlabel pdiffusion 19 49 19 49 3 Vdd
rlabel pdiffusion 19 56 19 56 3 Vdd
rlabel m1 52 38 52 38 3 _Y
rlabel m1 52 39 52 39 3 _Y
rlabel m1 52 42 52 42 3 _Y
rlabel m1 48 50 48 50 3 Y
port 3 e default output
rlabel m1 48 30 48 30 3 Y
port 3 e default output
rlabel pdcontact 46 50 46 50 3 Y
port 3 e default output
rlabel ndcontact 46 30 46 30 3 Y
port 3 e default output
rlabel m1 46 33 46 33 3 Y
port 3 e default output
rlabel m1 45 50 45 50 3 Y
port 3 e default output
rlabel m1 45 52 45 52 3 Y
port 3 e default output
rlabel m1 46 53 46 53 3 Y
port 3 e default output
rlabel m1 46 68 46 68 3 Y
port 3 e
rlabel m1 45 30 45 30 3 Y
port 3 e
rlabel m1 45 32 45 32 3 Y
port 3 e
rlabel m1 34 53 34 53 3 Vdd
rlabel m1 34 54 34 54 3 Vdd
rlabel m1 34 57 34 57 3 Vdd
rlabel m1 34 62 34 62 3 A
port 1 e default input
rlabel polycontact 32 62 32 62 3 A
port 1 e default input
rlabel m1 45 29 45 29 3 Y
port 3 e
rlabel m1 27 39 27 39 3 _Y
rlabel m1 45 49 45 49 3 Y
port 3 e
rlabel m1 30 50 30 50 3 _Y
rlabel m1 31 61 31 61 3 A
port 1 e default input
rlabel m1 31 62 31 62 3 A
port 1 e default input
rlabel m1 31 64 31 64 3 A
port 1 e default input
rlabel m1 31 65 31 65 3 A
port 1 e default input
rlabel m1 23 30 23 30 3 _Y
rlabel pdcontact 28 50 28 50 3 _Y
rlabel m1 22 18 22 18 3 B
port 2 e default input
rlabel m1 34 22 34 22 3 GND
rlabel ndcontact 21 30 21 30 3 _Y
rlabel m1 21 33 21 33 3 _Y
rlabel m1 27 38 27 38 3 _Y
rlabel m1 27 42 27 42 3 _Y
rlabel m1 27 43 27 43 3 _Y
rlabel m1 27 49 27 49 3 _Y
rlabel m1 27 50 27 50 3 _Y
rlabel m1 27 52 27 52 3 _Y
rlabel polycontact 20 18 20 18 3 B
port 2 e default input
rlabel m1 20 29 20 29 3 _Y
rlabel m1 20 30 20 30 3 _Y
rlabel m1 20 32 20 32 3 _Y
rlabel m1 19 12 19 12 3 B
port 2 e
rlabel m1 19 17 19 17 3 B
port 2 e
rlabel m1 19 18 19 18 3 B
port 2 e
rlabel m1 19 20 19 20 3 B
port 2 e
rlabel m1 19 53 19 53 3 Vdd
rlabel m1 19 54 19 54 3 Vdd
rlabel m1 19 57 19 57 3 Vdd
rlabel m1 19 68 19 68 3 A
port 1 e
rlabel m2 56 39 56 39 3 _Y
rlabel m2 55 39 55 39 3 _Y
rlabel m2c 53 39 53 39 3 _Y
rlabel m2 53 41 53 41 3 _Y
rlabel m2 38 54 38 54 3 Vdd
rlabel m2 38 23 38 23 3 GND
rlabel m2c 36 24 36 24 3 GND
rlabel m2 31 39 31 39 3 _Y
rlabel m2c 36 54 36 54 3 Vdd
rlabel m2c 35 23 35 23 3 GND
rlabel m2c 35 24 35 24 3 GND
rlabel m2c 28 39 28 39 3 _Y
rlabel m2c 35 54 35 54 3 Vdd
rlabel m2 35 56 35 56 3 Vdd
rlabel m2 34 11 34 11 3 GND
rlabel m2 34 23 34 23 3 GND
rlabel m2 34 26 34 26 3 GND
rlabel m2 23 39 23 39 3 _Y
rlabel m2 23 54 23 54 3 Vdd
rlabel m2c 20 39 20 39 3 _Y
rlabel m2 22 54 22 54 3 Vdd
rlabel m2 19 38 19 38 3 _Y
rlabel m2 19 39 19 39 3 _Y
rlabel m2 19 42 19 42 3 _Y
rlabel m2c 20 54 20 54 3 Vdd
rlabel m2 20 56 20 56 3 Vdd
rlabel m2 8 53 8 53 3 Vdd
rlabel m2 8 54 8 54 3 Vdd
rlabel m2 8 57 8 57 3 Vdd
<< properties >>
string FIXED_BBOX 0 0 60 80
string LEFclass CORE
string LEFsite CoreSite
string LEFsymmetry X Y
string LEFview TRUE
<< end >>
