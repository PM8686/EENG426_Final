magic
tech TSMC180
timestamp 1734143631
<< m1 >>
rect 6 17 9 20
rect 6 10 9 13
<< labels >>
rlabel m1 s 6 17 9 20 6 Vdd
port 1 nsew power input
rlabel m1 s 6 10 9 13 6 GND
port 2 nsew ground input
<< properties >>
string FIXED_BBOX 0 0 18 30
string LEFclass CORE WELLTAP
string LEFsite CoreSite
string LEFsymmetry X Y
string LEFview TRUE
<< end >>
