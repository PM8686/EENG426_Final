magic
tech sky130l
timestamp 1731032673
<< ndiffusion >>
rect 8 15 13 16
rect 8 12 9 15
rect 12 12 13 15
rect 8 6 13 12
rect 15 6 20 16
rect 22 14 27 16
rect 22 11 23 14
rect 26 11 27 14
rect 22 10 27 11
rect 29 15 34 16
rect 29 12 30 15
rect 33 12 34 15
rect 29 10 34 12
rect 22 6 26 10
<< ndc >>
rect 9 12 12 15
rect 23 11 26 14
rect 30 12 33 15
<< ntransistor >>
rect 13 6 15 16
rect 20 6 22 16
rect 27 10 29 16
<< pdiffusion >>
rect 8 30 13 31
rect 8 27 9 30
rect 12 27 13 30
rect 8 23 13 27
rect 15 27 20 31
rect 15 24 16 27
rect 19 24 20 27
rect 15 23 20 24
rect 22 30 27 31
rect 22 27 23 30
rect 26 27 27 30
rect 22 23 27 27
rect 29 30 34 31
rect 29 27 30 30
rect 33 27 34 30
rect 29 23 34 27
<< pdc >>
rect 9 27 12 30
rect 16 24 19 27
rect 23 27 26 30
rect 30 27 33 30
<< ptransistor >>
rect 13 23 15 31
rect 20 23 22 31
rect 27 23 29 31
<< polysilicon >>
rect 16 40 22 41
rect 16 37 17 40
rect 20 37 22 40
rect 16 36 22 37
rect 13 31 15 33
rect 20 31 22 36
rect 27 31 29 33
rect 13 16 15 23
rect 20 16 22 23
rect 27 20 29 23
rect 27 19 41 20
rect 27 18 37 19
rect 27 16 29 18
rect 36 16 37 18
rect 40 16 41 19
rect 36 15 41 16
rect 27 8 29 10
rect 13 4 15 6
rect 20 4 22 6
rect 8 3 15 4
rect 8 0 9 3
rect 12 0 15 3
rect 8 -1 15 0
<< pc >>
rect 17 37 20 40
rect 37 16 40 19
rect 9 0 12 3
<< m1 >>
rect 8 40 12 44
rect 9 37 17 40
rect 20 37 21 40
rect 40 35 44 36
rect 30 32 44 35
rect 9 30 12 31
rect 23 30 26 31
rect 9 26 12 27
rect 16 27 19 28
rect 23 26 26 27
rect 30 30 33 32
rect 9 19 12 20
rect 9 15 12 16
rect 16 19 19 24
rect 16 15 19 16
rect 30 15 33 27
rect 37 19 40 20
rect 37 15 40 16
rect 9 11 12 12
rect 23 14 26 15
rect 30 11 33 12
rect 23 8 26 11
rect 23 5 24 8
rect 27 5 28 8
rect 23 4 28 5
rect 1 0 9 3
rect 12 0 13 3
rect 0 -4 4 0
<< m2c >>
rect 9 27 12 30
rect 23 27 26 30
rect 9 16 12 19
rect 16 16 19 19
rect 37 16 40 19
rect 24 5 27 8
<< m2 >>
rect 8 30 27 31
rect 8 27 9 30
rect 12 27 23 30
rect 26 27 27 30
rect 8 26 27 27
rect 8 19 41 20
rect 8 16 9 19
rect 12 16 16 19
rect 19 16 37 19
rect 40 16 41 19
rect 8 15 41 16
rect 23 8 28 9
rect 23 5 24 8
rect 27 5 28 8
rect 23 4 28 5
<< labels >>
rlabel ndiffusion 30 11 30 11 3 Y
rlabel polysilicon 28 17 28 17 3 _Y
rlabel polysilicon 28 22 28 22 3 _Y
rlabel pdiffusion 30 24 30 24 3 Y
rlabel ndiffusion 23 7 23 7 3 GND
rlabel pdiffusion 23 24 23 24 3 Vdd
rlabel polysilicon 21 17 21 17 3 A
rlabel polysilicon 21 22 21 22 3 A
rlabel pdiffusion 16 24 16 24 3 _Y
rlabel polysilicon 14 17 14 17 3 B
rlabel polysilicon 14 22 14 22 3 B
rlabel ndiffusion 9 7 9 7 3 _Y
rlabel pdiffusion 9 24 9 24 3 Vdd
rlabel m1 33 33 33 33 3 Y
rlabel m2 25 5 25 5 3 GND
rlabel m2 9 30 9 30 3 Vdd
rlabel m1 9 41 9 41 3 A
rlabel m1 1 -3 1 -3 3 B
<< end >>
