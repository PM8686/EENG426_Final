magic
tech sky130l
timestamp 1729042338
<< ndiffusion >>
rect 8 10 13 12
rect 8 7 9 10
rect 12 7 13 10
rect 8 6 13 7
rect 15 11 20 12
rect 15 8 16 11
rect 19 8 20 11
rect 15 6 20 8
<< ndc >>
rect 9 7 12 10
rect 16 8 19 11
<< ntransistor >>
rect 13 6 15 12
<< pdiffusion >>
rect 8 26 13 27
rect 8 23 9 26
rect 12 23 13 26
rect 8 19 13 23
rect 15 23 20 27
rect 15 20 16 23
rect 19 20 20 23
rect 15 19 20 20
<< pdc >>
rect 9 23 12 26
rect 16 20 19 23
<< ptransistor >>
rect 13 19 15 27
<< polysilicon >>
rect 13 34 20 35
rect 13 31 16 34
rect 19 31 20 34
rect 13 30 20 31
rect 13 27 15 30
rect 13 12 15 19
rect 13 4 15 6
<< pc >>
rect 16 31 19 34
<< m1 >>
rect 16 34 20 35
rect 8 31 12 32
rect 8 28 9 31
rect 19 31 20 34
rect 16 28 20 31
rect 8 26 12 28
rect 8 23 9 26
rect 8 22 12 23
rect 16 23 20 24
rect 19 20 20 23
rect 16 11 20 20
rect 8 10 12 11
rect 8 7 9 10
rect 8 4 12 7
rect 19 8 20 11
rect 16 4 20 8
<< m2c >>
rect 9 28 12 31
rect 9 7 12 10
<< m2 >>
rect 8 31 13 32
rect 8 28 9 31
rect 12 28 13 31
rect 8 27 13 28
rect 8 10 13 11
rect 8 7 9 10
rect 12 7 13 10
rect 8 6 13 7
<< labels >>
rlabel ndiffusion 16 7 16 7 3 Y
rlabel pdiffusion 16 20 16 20 3 Y
rlabel polysilicon 14 13 14 13 3 A
rlabel polysilicon 14 18 14 18 3 A
rlabel pdiffusion 9 20 9 20 3 Vdd
rlabel m1 17 5 17 5 3 Y
rlabel m1 9 5 9 5 3 GND
rlabel m1 17 29 17 29 3 A
rlabel m2 9 29 9 29 3 Vdd
rlabel m2 9 7 9 7 3 GND
<< end >>
