magic
tech sky130l
timestamp 1731001260
<< m1 >>
rect 144 875 148 911
rect 232 891 236 911
rect 352 735 356 763
rect 840 455 844 479
<< m2c >>
rect 111 1197 115 1201
rect 1111 1197 1115 1201
rect 111 1179 115 1183
rect 1111 1179 1115 1183
rect 111 1129 115 1133
rect 1111 1129 1115 1133
rect 111 1111 115 1115
rect 1111 1111 1115 1115
rect 111 1069 115 1073
rect 1111 1069 1115 1073
rect 111 1051 115 1055
rect 1111 1051 1115 1055
rect 111 1001 115 1005
rect 1111 1001 1115 1005
rect 111 983 115 987
rect 1111 983 1115 987
rect 111 925 115 929
rect 1111 925 1115 929
rect 144 911 148 915
rect 111 907 115 911
rect 232 911 236 915
rect 1111 907 1115 911
rect 232 887 236 891
rect 144 871 148 875
rect 111 849 115 853
rect 1111 849 1115 853
rect 111 831 115 835
rect 1111 831 1115 835
rect 111 777 115 781
rect 1111 777 1115 781
rect 352 763 356 767
rect 111 759 115 763
rect 1111 759 1115 763
rect 352 731 356 735
rect 111 705 115 709
rect 1111 705 1115 709
rect 111 687 115 691
rect 1111 687 1115 691
rect 111 645 115 649
rect 1111 645 1115 649
rect 111 627 115 631
rect 1111 627 1115 631
rect 111 565 115 569
rect 1111 565 1115 569
rect 111 547 115 551
rect 1111 547 1115 551
rect 111 493 115 497
rect 1111 493 1115 497
rect 840 479 844 483
rect 111 475 115 479
rect 1111 475 1115 479
rect 840 451 844 455
rect 111 421 115 425
rect 1111 421 1115 425
rect 111 403 115 407
rect 1111 403 1115 407
rect 111 361 115 365
rect 1111 361 1115 365
rect 111 343 115 347
rect 1111 343 1115 347
rect 111 293 115 297
rect 1111 293 1115 297
rect 111 275 115 279
rect 1111 275 1115 279
rect 111 225 115 229
rect 1111 225 1115 229
rect 111 207 115 211
rect 1111 207 1115 211
rect 111 141 115 145
rect 1111 141 1115 145
rect 111 123 115 127
rect 1111 123 1115 127
<< m2 >>
rect 134 1216 140 1217
rect 134 1212 135 1216
rect 139 1212 140 1216
rect 134 1211 140 1212
rect 222 1216 228 1217
rect 222 1212 223 1216
rect 227 1212 228 1216
rect 222 1211 228 1212
rect 310 1216 316 1217
rect 310 1212 311 1216
rect 315 1212 316 1216
rect 310 1211 316 1212
rect 110 1201 116 1202
rect 110 1197 111 1201
rect 115 1197 116 1201
rect 110 1196 116 1197
rect 1110 1201 1116 1202
rect 1110 1197 1111 1201
rect 1115 1197 1116 1201
rect 1110 1196 1116 1197
rect 202 1187 208 1188
rect 110 1183 116 1184
rect 110 1179 111 1183
rect 115 1179 116 1183
rect 110 1178 116 1179
rect 142 1171 148 1172
rect 142 1167 143 1171
rect 147 1167 148 1171
rect 142 1166 148 1167
rect 162 1163 168 1164
rect 162 1159 163 1163
rect 167 1159 168 1163
rect 196 1162 198 1185
rect 202 1183 203 1187
rect 207 1186 208 1187
rect 290 1187 296 1188
rect 207 1184 249 1186
rect 207 1183 208 1184
rect 202 1182 208 1183
rect 290 1183 291 1187
rect 295 1186 296 1187
rect 295 1184 337 1186
rect 295 1183 296 1184
rect 290 1182 296 1183
rect 1110 1183 1116 1184
rect 1110 1179 1111 1183
rect 1115 1179 1116 1183
rect 1110 1178 1116 1179
rect 230 1171 236 1172
rect 230 1167 231 1171
rect 235 1167 236 1171
rect 230 1166 236 1167
rect 318 1171 324 1172
rect 318 1167 319 1171
rect 323 1167 324 1171
rect 318 1166 324 1167
rect 162 1158 168 1159
rect 192 1160 198 1162
rect 250 1163 256 1164
rect 192 1155 194 1160
rect 250 1159 251 1163
rect 255 1159 256 1163
rect 250 1158 256 1159
rect 410 1163 416 1164
rect 410 1159 411 1163
rect 415 1162 416 1163
rect 415 1160 458 1162
rect 415 1159 416 1160
rect 410 1158 416 1159
rect 270 1155 276 1156
rect 270 1151 271 1155
rect 275 1154 276 1155
rect 358 1155 364 1156
rect 456 1155 458 1160
rect 275 1152 281 1154
rect 275 1151 276 1152
rect 270 1150 276 1151
rect 358 1151 359 1155
rect 363 1154 364 1155
rect 363 1152 369 1154
rect 363 1151 364 1152
rect 358 1150 364 1151
rect 174 1145 180 1146
rect 174 1141 175 1145
rect 179 1141 180 1145
rect 174 1140 180 1141
rect 262 1145 268 1146
rect 262 1141 263 1145
rect 267 1141 268 1145
rect 262 1140 268 1141
rect 350 1145 356 1146
rect 350 1141 351 1145
rect 355 1141 356 1145
rect 350 1140 356 1141
rect 438 1145 444 1146
rect 438 1141 439 1145
rect 443 1141 444 1145
rect 438 1140 444 1141
rect 110 1133 116 1134
rect 110 1129 111 1133
rect 115 1129 116 1133
rect 1110 1133 1116 1134
rect 410 1131 416 1132
rect 410 1130 411 1131
rect 110 1128 116 1129
rect 405 1128 411 1130
rect 258 1127 264 1128
rect 258 1126 259 1127
rect 229 1124 259 1126
rect 258 1123 259 1124
rect 263 1123 264 1127
rect 346 1127 352 1128
rect 346 1126 347 1127
rect 317 1124 347 1126
rect 258 1122 264 1123
rect 346 1123 347 1124
rect 351 1123 352 1127
rect 410 1127 411 1128
rect 415 1127 416 1131
rect 1110 1129 1111 1133
rect 1115 1129 1116 1133
rect 1110 1128 1116 1129
rect 410 1126 416 1127
rect 346 1122 352 1123
rect 110 1115 116 1116
rect 110 1111 111 1115
rect 115 1111 116 1115
rect 110 1110 116 1111
rect 422 1115 428 1116
rect 422 1111 423 1115
rect 427 1114 428 1115
rect 1110 1115 1116 1116
rect 427 1112 449 1114
rect 427 1111 428 1112
rect 422 1110 428 1111
rect 1110 1111 1111 1115
rect 1115 1111 1116 1115
rect 1110 1110 1116 1111
rect 166 1100 172 1101
rect 166 1096 167 1100
rect 171 1096 172 1100
rect 166 1095 172 1096
rect 254 1100 260 1101
rect 254 1096 255 1100
rect 259 1096 260 1100
rect 254 1095 260 1096
rect 342 1100 348 1101
rect 342 1096 343 1100
rect 347 1096 348 1100
rect 342 1095 348 1096
rect 430 1100 436 1101
rect 430 1096 431 1100
rect 435 1096 436 1100
rect 430 1095 436 1096
rect 954 1091 960 1092
rect 398 1088 404 1089
rect 398 1084 399 1088
rect 403 1084 404 1088
rect 398 1083 404 1084
rect 486 1088 492 1089
rect 486 1084 487 1088
rect 491 1084 492 1088
rect 486 1083 492 1084
rect 574 1088 580 1089
rect 574 1084 575 1088
rect 579 1084 580 1088
rect 574 1083 580 1084
rect 662 1088 668 1089
rect 662 1084 663 1088
rect 667 1084 668 1088
rect 662 1083 668 1084
rect 750 1088 756 1089
rect 750 1084 751 1088
rect 755 1084 756 1088
rect 750 1083 756 1084
rect 838 1088 844 1089
rect 838 1084 839 1088
rect 843 1084 844 1088
rect 838 1083 844 1084
rect 926 1088 932 1089
rect 926 1084 927 1088
rect 931 1084 932 1088
rect 954 1087 955 1091
rect 959 1090 960 1091
rect 959 1088 998 1090
rect 959 1087 960 1088
rect 954 1086 960 1087
rect 926 1083 932 1084
rect 996 1074 998 1088
rect 1014 1088 1020 1089
rect 1014 1084 1015 1088
rect 1019 1084 1020 1088
rect 1014 1083 1020 1084
rect 110 1073 116 1074
rect 110 1069 111 1073
rect 115 1069 116 1073
rect 996 1072 1033 1074
rect 1110 1073 1116 1074
rect 110 1068 116 1069
rect 1110 1069 1111 1073
rect 1115 1069 1116 1073
rect 1110 1068 1116 1069
rect 494 1063 500 1064
rect 494 1059 495 1063
rect 499 1059 500 1063
rect 494 1058 500 1059
rect 582 1063 588 1064
rect 582 1059 583 1063
rect 587 1059 588 1063
rect 582 1058 588 1059
rect 670 1063 676 1064
rect 670 1059 671 1063
rect 675 1059 676 1063
rect 758 1063 764 1064
rect 670 1058 676 1059
rect 742 1059 748 1060
rect 742 1058 743 1059
rect 461 1056 498 1058
rect 549 1056 586 1058
rect 637 1056 674 1058
rect 725 1056 743 1058
rect 110 1055 116 1056
rect 110 1051 111 1055
rect 115 1051 116 1055
rect 742 1055 743 1056
rect 747 1055 748 1059
rect 758 1059 759 1063
rect 763 1059 764 1063
rect 934 1063 940 1064
rect 934 1062 935 1063
rect 758 1058 764 1059
rect 919 1060 935 1062
rect 919 1058 921 1060
rect 934 1059 935 1060
rect 939 1059 940 1063
rect 934 1058 940 1059
rect 1022 1063 1028 1064
rect 1022 1059 1023 1063
rect 1027 1059 1028 1063
rect 1022 1058 1028 1059
rect 760 1056 777 1058
rect 901 1056 921 1058
rect 989 1056 1026 1058
rect 742 1054 748 1055
rect 1110 1055 1116 1056
rect 110 1050 116 1051
rect 1110 1051 1111 1055
rect 1115 1051 1116 1055
rect 1110 1050 1116 1051
rect 406 1043 412 1044
rect 406 1039 407 1043
rect 411 1039 412 1043
rect 406 1038 412 1039
rect 494 1043 500 1044
rect 494 1039 495 1043
rect 499 1039 500 1043
rect 494 1038 500 1039
rect 582 1043 588 1044
rect 582 1039 583 1043
rect 587 1039 588 1043
rect 582 1038 588 1039
rect 670 1043 676 1044
rect 670 1039 671 1043
rect 675 1039 676 1043
rect 670 1038 676 1039
rect 758 1043 764 1044
rect 758 1039 759 1043
rect 763 1039 764 1043
rect 758 1038 764 1039
rect 846 1043 852 1044
rect 846 1039 847 1043
rect 851 1039 852 1043
rect 846 1038 852 1039
rect 934 1043 940 1044
rect 934 1039 935 1043
rect 939 1039 940 1043
rect 934 1038 940 1039
rect 1022 1043 1028 1044
rect 1022 1039 1023 1043
rect 1027 1039 1028 1043
rect 1022 1038 1028 1039
rect 422 1035 428 1036
rect 422 1031 423 1035
rect 427 1031 428 1035
rect 422 1030 428 1031
rect 502 1035 508 1036
rect 502 1031 503 1035
rect 507 1034 508 1035
rect 590 1035 596 1036
rect 507 1032 513 1034
rect 507 1031 508 1032
rect 502 1030 508 1031
rect 590 1031 591 1035
rect 595 1034 596 1035
rect 678 1035 684 1036
rect 595 1032 601 1034
rect 595 1031 596 1032
rect 590 1030 596 1031
rect 678 1031 679 1035
rect 683 1034 684 1035
rect 774 1035 780 1036
rect 683 1032 689 1034
rect 683 1031 684 1032
rect 678 1030 684 1031
rect 774 1031 775 1035
rect 779 1031 780 1035
rect 774 1030 780 1031
rect 854 1035 860 1036
rect 854 1031 855 1035
rect 859 1034 860 1035
rect 942 1035 948 1036
rect 859 1032 865 1034
rect 859 1031 860 1032
rect 854 1030 860 1031
rect 942 1031 943 1035
rect 947 1034 948 1035
rect 1030 1035 1036 1036
rect 947 1032 953 1034
rect 947 1031 948 1032
rect 942 1030 948 1031
rect 1030 1031 1031 1035
rect 1035 1034 1036 1035
rect 1035 1032 1041 1034
rect 1035 1031 1036 1032
rect 1030 1030 1036 1031
rect 502 1027 508 1028
rect 414 1023 420 1024
rect 502 1023 503 1027
rect 507 1026 508 1027
rect 590 1027 596 1028
rect 507 1024 513 1026
rect 507 1023 508 1024
rect 414 1019 415 1023
rect 419 1022 420 1023
rect 424 1022 426 1023
rect 502 1022 508 1023
rect 590 1023 591 1027
rect 595 1026 596 1027
rect 766 1027 772 1028
rect 595 1024 601 1026
rect 595 1023 596 1024
rect 590 1022 596 1023
rect 678 1023 684 1024
rect 766 1023 767 1027
rect 771 1026 772 1027
rect 1030 1027 1036 1028
rect 771 1024 777 1026
rect 862 1025 868 1026
rect 771 1023 772 1024
rect 419 1020 426 1022
rect 419 1019 420 1020
rect 414 1018 420 1019
rect 678 1019 679 1023
rect 683 1022 684 1023
rect 688 1022 690 1023
rect 766 1022 772 1023
rect 683 1020 690 1022
rect 862 1021 863 1025
rect 867 1021 868 1025
rect 862 1020 868 1021
rect 954 1025 960 1026
rect 954 1021 955 1025
rect 959 1021 960 1025
rect 1030 1023 1031 1027
rect 1035 1026 1036 1027
rect 1035 1024 1041 1026
rect 1035 1023 1036 1024
rect 1030 1022 1036 1023
rect 954 1020 960 1021
rect 683 1019 684 1020
rect 678 1018 684 1019
rect 406 1017 412 1018
rect 406 1013 407 1017
rect 411 1013 412 1017
rect 406 1012 412 1013
rect 494 1017 500 1018
rect 494 1013 495 1017
rect 499 1013 500 1017
rect 494 1012 500 1013
rect 582 1017 588 1018
rect 582 1013 583 1017
rect 587 1013 588 1017
rect 582 1012 588 1013
rect 670 1017 676 1018
rect 670 1013 671 1017
rect 675 1013 676 1017
rect 670 1012 676 1013
rect 758 1017 764 1018
rect 758 1013 759 1017
rect 763 1013 764 1017
rect 758 1012 764 1013
rect 846 1017 852 1018
rect 846 1013 847 1017
rect 851 1013 852 1017
rect 846 1012 852 1013
rect 934 1017 940 1018
rect 934 1013 935 1017
rect 939 1013 940 1017
rect 934 1012 940 1013
rect 1022 1017 1028 1018
rect 1022 1013 1023 1017
rect 1027 1013 1028 1017
rect 1022 1012 1028 1013
rect 110 1005 116 1006
rect 110 1001 111 1005
rect 115 1001 116 1005
rect 110 1000 116 1001
rect 1110 1005 1116 1006
rect 1110 1001 1111 1005
rect 1115 1001 1116 1005
rect 1110 1000 1116 1001
rect 490 999 496 1000
rect 490 998 491 999
rect 461 996 491 998
rect 490 995 491 996
rect 495 995 496 999
rect 578 999 584 1000
rect 578 998 579 999
rect 549 996 579 998
rect 490 994 496 995
rect 578 995 579 996
rect 583 995 584 999
rect 578 994 584 995
rect 650 999 656 1000
rect 650 995 651 999
rect 655 998 656 999
rect 738 999 744 1000
rect 655 996 689 998
rect 655 995 656 996
rect 650 994 656 995
rect 738 995 739 999
rect 743 998 744 999
rect 846 999 852 1000
rect 743 996 777 998
rect 743 995 744 996
rect 738 994 744 995
rect 846 995 847 999
rect 851 998 852 999
rect 1018 999 1024 1000
rect 1018 998 1019 999
rect 851 996 865 998
rect 989 996 1019 998
rect 851 995 852 996
rect 846 994 852 995
rect 1018 995 1019 996
rect 1023 995 1024 999
rect 1018 994 1024 995
rect 110 987 116 988
rect 110 983 111 987
rect 115 983 116 987
rect 670 987 676 988
rect 670 986 671 987
rect 633 984 671 986
rect 110 982 116 983
rect 670 983 671 984
rect 675 983 676 987
rect 670 982 676 983
rect 1022 987 1028 988
rect 1022 983 1023 987
rect 1027 986 1028 987
rect 1110 987 1116 988
rect 1027 984 1033 986
rect 1027 983 1028 984
rect 1022 982 1028 983
rect 1110 983 1111 987
rect 1115 983 1116 987
rect 1110 982 1116 983
rect 398 972 404 973
rect 398 968 399 972
rect 403 968 404 972
rect 398 967 404 968
rect 486 972 492 973
rect 486 968 487 972
rect 491 968 492 972
rect 486 967 492 968
rect 574 972 580 973
rect 574 968 575 972
rect 579 968 580 972
rect 574 967 580 968
rect 662 972 668 973
rect 662 968 663 972
rect 667 968 668 972
rect 662 967 668 968
rect 750 972 756 973
rect 750 968 751 972
rect 755 968 756 972
rect 750 967 756 968
rect 838 972 844 973
rect 838 968 839 972
rect 843 968 844 972
rect 838 967 844 968
rect 926 972 932 973
rect 926 968 927 972
rect 931 968 932 972
rect 926 967 932 968
rect 1014 972 1020 973
rect 1014 968 1015 972
rect 1019 968 1020 972
rect 1014 967 1020 968
rect 150 944 156 945
rect 150 940 151 944
rect 155 940 156 944
rect 150 939 156 940
rect 270 944 276 945
rect 270 940 271 944
rect 275 940 276 944
rect 270 939 276 940
rect 406 944 412 945
rect 406 940 407 944
rect 411 940 412 944
rect 406 939 412 940
rect 550 944 556 945
rect 550 940 551 944
rect 555 940 556 944
rect 550 939 556 940
rect 710 944 716 945
rect 710 940 711 944
rect 715 940 716 944
rect 710 939 716 940
rect 870 944 876 945
rect 870 940 871 944
rect 875 940 876 944
rect 870 939 876 940
rect 1014 944 1020 945
rect 1014 940 1015 944
rect 1019 940 1020 944
rect 1014 939 1020 940
rect 862 931 868 932
rect 110 929 116 930
rect 110 925 111 929
rect 115 925 116 929
rect 862 927 863 931
rect 867 930 868 931
rect 867 928 889 930
rect 1110 929 1116 930
rect 867 927 868 928
rect 862 926 868 927
rect 110 924 116 925
rect 1110 925 1111 929
rect 1115 925 1116 929
rect 1110 924 1116 925
rect 143 915 149 916
rect 110 911 116 912
rect 110 907 111 911
rect 115 907 116 911
rect 143 911 144 915
rect 148 914 149 915
rect 231 915 237 916
rect 148 912 177 914
rect 148 911 149 912
rect 143 910 149 911
rect 231 911 232 915
rect 236 914 237 915
rect 370 915 376 916
rect 236 912 297 914
rect 236 911 237 912
rect 231 910 237 911
rect 370 911 371 915
rect 375 914 376 915
rect 502 915 508 916
rect 375 912 433 914
rect 375 911 376 912
rect 370 910 376 911
rect 502 911 503 915
rect 507 914 508 915
rect 654 915 660 916
rect 507 912 577 914
rect 507 911 508 912
rect 502 910 508 911
rect 654 911 655 915
rect 659 914 660 915
rect 1082 915 1088 916
rect 1082 914 1083 915
rect 659 912 737 914
rect 1077 912 1083 914
rect 659 911 660 912
rect 654 910 660 911
rect 1082 911 1083 912
rect 1087 911 1088 915
rect 1082 910 1088 911
rect 1110 911 1116 912
rect 110 906 116 907
rect 1110 907 1111 911
rect 1115 907 1116 911
rect 1110 906 1116 907
rect 158 899 164 900
rect 158 895 159 899
rect 163 895 164 899
rect 158 894 164 895
rect 278 899 284 900
rect 278 895 279 899
rect 283 895 284 899
rect 278 894 284 895
rect 414 899 420 900
rect 414 895 415 899
rect 419 895 420 899
rect 414 894 420 895
rect 558 899 564 900
rect 558 895 559 899
rect 563 895 564 899
rect 558 894 564 895
rect 718 899 724 900
rect 718 895 719 899
rect 723 895 724 899
rect 718 894 724 895
rect 878 899 884 900
rect 878 895 879 899
rect 883 895 884 899
rect 878 894 884 895
rect 1022 899 1028 900
rect 1022 895 1023 899
rect 1027 895 1028 899
rect 1022 894 1028 895
rect 231 891 237 892
rect 231 890 232 891
rect 212 888 232 890
rect 176 882 178 885
rect 212 882 214 888
rect 231 887 232 888
rect 236 887 237 891
rect 231 886 237 887
rect 1030 891 1036 892
rect 1030 887 1031 891
rect 1035 890 1036 891
rect 1035 888 1041 890
rect 1035 887 1036 888
rect 1030 886 1036 887
rect 176 880 214 882
rect 218 883 224 884
rect 218 879 219 883
rect 223 882 224 883
rect 296 882 298 885
rect 370 883 376 884
rect 370 882 371 883
rect 223 880 290 882
rect 296 880 371 882
rect 223 879 224 880
rect 218 878 224 879
rect 143 875 149 876
rect 288 875 290 880
rect 370 879 371 880
rect 375 879 376 883
rect 432 882 434 885
rect 502 883 508 884
rect 502 882 503 883
rect 432 880 503 882
rect 370 878 376 879
rect 502 879 503 880
rect 507 879 508 883
rect 576 882 578 885
rect 654 883 660 884
rect 654 882 655 883
rect 576 880 655 882
rect 502 878 508 879
rect 654 879 655 880
rect 659 879 660 883
rect 654 878 660 879
rect 670 883 676 884
rect 670 879 671 883
rect 675 882 676 883
rect 736 882 738 885
rect 675 880 738 882
rect 754 883 760 884
rect 675 879 676 880
rect 670 878 676 879
rect 754 879 755 883
rect 759 882 760 883
rect 896 882 898 885
rect 930 883 936 884
rect 930 882 931 883
rect 759 880 858 882
rect 896 880 931 882
rect 759 879 760 880
rect 754 878 760 879
rect 446 875 452 876
rect 143 871 144 875
rect 148 874 149 875
rect 148 872 161 874
rect 148 871 149 872
rect 143 870 149 871
rect 446 871 447 875
rect 451 874 452 875
rect 638 875 644 876
rect 856 875 858 880
rect 930 879 931 880
rect 935 879 936 883
rect 1082 883 1088 884
rect 1082 882 1083 883
rect 930 878 936 879
rect 1040 880 1083 882
rect 1040 875 1042 880
rect 1082 879 1083 880
rect 1087 879 1088 883
rect 1082 878 1088 879
rect 451 872 457 874
rect 451 871 452 872
rect 446 870 452 871
rect 638 871 639 875
rect 643 874 644 875
rect 643 872 649 874
rect 643 871 644 872
rect 638 870 644 871
rect 142 865 148 866
rect 142 861 143 865
rect 147 861 148 865
rect 142 860 148 861
rect 270 865 276 866
rect 270 861 271 865
rect 275 861 276 865
rect 270 860 276 861
rect 438 865 444 866
rect 438 861 439 865
rect 443 861 444 865
rect 438 860 444 861
rect 630 865 636 866
rect 630 861 631 865
rect 635 861 636 865
rect 630 860 636 861
rect 838 865 844 866
rect 838 861 839 865
rect 843 861 844 865
rect 838 860 844 861
rect 1022 865 1028 866
rect 1022 861 1023 865
rect 1027 861 1028 865
rect 1022 860 1028 861
rect 110 853 116 854
rect 110 849 111 853
rect 115 849 116 853
rect 1110 853 1116 854
rect 218 851 224 852
rect 218 850 219 851
rect 110 848 116 849
rect 197 848 219 850
rect 218 847 219 848
rect 223 847 224 851
rect 754 851 760 852
rect 754 850 755 851
rect 685 848 755 850
rect 218 846 224 847
rect 434 847 440 848
rect 434 846 435 847
rect 325 844 435 846
rect 434 843 435 844
rect 439 843 440 847
rect 626 847 632 848
rect 626 846 627 847
rect 493 844 627 846
rect 434 842 440 843
rect 626 843 627 844
rect 631 843 632 847
rect 754 847 755 848
rect 759 847 760 851
rect 1110 849 1111 853
rect 1115 849 1116 853
rect 1110 848 1116 849
rect 754 846 760 847
rect 626 842 632 843
rect 110 835 116 836
rect 110 831 111 835
rect 115 831 116 835
rect 110 830 116 831
rect 738 835 744 836
rect 738 831 739 835
rect 743 834 744 835
rect 1022 835 1028 836
rect 743 832 849 834
rect 743 831 744 832
rect 738 830 744 831
rect 1022 831 1023 835
rect 1027 834 1028 835
rect 1110 835 1116 836
rect 1027 832 1033 834
rect 1027 831 1028 832
rect 1022 830 1028 831
rect 1110 831 1111 835
rect 1115 831 1116 835
rect 1110 830 1116 831
rect 134 820 140 821
rect 134 816 135 820
rect 139 816 140 820
rect 134 815 140 816
rect 262 820 268 821
rect 262 816 263 820
rect 267 816 268 820
rect 262 815 268 816
rect 430 820 436 821
rect 430 816 431 820
rect 435 816 436 820
rect 430 815 436 816
rect 622 820 628 821
rect 622 816 623 820
rect 627 816 628 820
rect 622 815 628 816
rect 830 820 836 821
rect 830 816 831 820
rect 835 816 836 820
rect 830 815 836 816
rect 1014 820 1020 821
rect 1014 816 1015 820
rect 1019 816 1020 820
rect 1014 815 1020 816
rect 134 796 140 797
rect 134 792 135 796
rect 139 792 140 796
rect 134 791 140 792
rect 238 796 244 797
rect 238 792 239 796
rect 243 792 244 796
rect 238 791 244 792
rect 374 796 380 797
rect 374 792 375 796
rect 379 792 380 796
rect 374 791 380 792
rect 526 796 532 797
rect 526 792 527 796
rect 531 792 532 796
rect 526 791 532 792
rect 694 796 700 797
rect 694 792 695 796
rect 699 792 700 796
rect 694 791 700 792
rect 862 796 868 797
rect 862 792 863 796
rect 867 792 868 796
rect 862 791 868 792
rect 1014 796 1020 797
rect 1014 792 1015 796
rect 1019 792 1020 796
rect 1014 791 1020 792
rect 930 783 936 784
rect 930 782 931 783
rect 110 781 116 782
rect 110 777 111 781
rect 115 777 116 781
rect 921 780 931 782
rect 930 779 931 780
rect 935 779 936 783
rect 930 778 936 779
rect 1110 781 1116 782
rect 110 776 116 777
rect 1110 777 1111 781
rect 1115 777 1116 781
rect 1110 776 1116 777
rect 1022 771 1028 772
rect 210 767 216 768
rect 210 766 211 767
rect 197 764 211 766
rect 110 763 116 764
rect 110 759 111 763
rect 115 759 116 763
rect 210 763 211 764
rect 215 763 216 767
rect 351 767 357 768
rect 351 766 352 767
rect 301 764 352 766
rect 210 762 216 763
rect 351 763 352 764
rect 356 763 357 767
rect 482 767 488 768
rect 482 766 483 767
rect 437 764 483 766
rect 351 762 357 763
rect 482 763 483 764
rect 487 763 488 767
rect 674 767 680 768
rect 674 766 675 767
rect 589 764 675 766
rect 482 762 488 763
rect 674 763 675 764
rect 679 763 680 767
rect 674 762 680 763
rect 682 767 688 768
rect 682 763 683 767
rect 687 766 688 767
rect 1022 767 1023 771
rect 1027 767 1028 771
rect 1022 766 1028 767
rect 687 764 721 766
rect 1024 764 1041 766
rect 687 763 688 764
rect 682 762 688 763
rect 1110 763 1116 764
rect 110 758 116 759
rect 1110 759 1111 763
rect 1115 759 1116 763
rect 1110 758 1116 759
rect 142 751 148 752
rect 142 747 143 751
rect 147 747 148 751
rect 142 746 148 747
rect 246 751 252 752
rect 246 747 247 751
rect 251 747 252 751
rect 246 746 252 747
rect 382 751 388 752
rect 382 747 383 751
rect 387 747 388 751
rect 382 746 388 747
rect 534 751 540 752
rect 534 747 535 751
rect 539 747 540 751
rect 534 746 540 747
rect 702 751 708 752
rect 702 747 703 751
rect 707 747 708 751
rect 702 746 708 747
rect 870 751 876 752
rect 870 747 871 751
rect 875 747 876 751
rect 870 746 876 747
rect 1022 751 1028 752
rect 1022 747 1023 751
rect 1027 747 1028 751
rect 1022 746 1028 747
rect 162 743 168 744
rect 162 739 163 743
rect 167 739 168 743
rect 886 743 892 744
rect 162 738 168 739
rect 248 740 265 742
rect 210 735 216 736
rect 210 731 211 735
rect 215 734 216 735
rect 248 734 250 740
rect 430 739 436 740
rect 215 732 250 734
rect 351 735 357 736
rect 215 731 216 732
rect 210 730 216 731
rect 290 731 296 732
rect 290 727 291 731
rect 295 727 296 731
rect 351 731 352 735
rect 356 734 357 735
rect 400 734 402 737
rect 430 735 431 739
rect 435 738 436 739
rect 582 739 588 740
rect 435 736 466 738
rect 435 735 436 736
rect 430 734 436 735
rect 356 732 402 734
rect 356 731 357 732
rect 464 731 466 736
rect 482 735 488 736
rect 482 731 483 735
rect 487 734 488 735
rect 552 734 554 737
rect 582 735 583 739
rect 587 738 588 739
rect 750 739 756 740
rect 587 736 658 738
rect 587 735 588 736
rect 582 734 588 735
rect 487 732 554 734
rect 487 731 488 732
rect 656 731 658 736
rect 674 735 680 736
rect 674 731 675 735
rect 679 734 680 735
rect 720 734 722 737
rect 750 735 751 739
rect 755 738 756 739
rect 886 739 887 743
rect 891 739 892 743
rect 886 738 892 739
rect 1038 743 1044 744
rect 1038 739 1039 743
rect 1043 739 1044 743
rect 1038 738 1044 739
rect 755 736 850 738
rect 755 735 756 736
rect 750 734 756 735
rect 679 732 722 734
rect 679 731 680 732
rect 848 731 850 736
rect 1030 731 1036 732
rect 351 730 357 731
rect 482 730 488 731
rect 674 730 680 731
rect 290 726 296 727
rect 1030 727 1031 731
rect 1035 730 1036 731
rect 1035 728 1041 730
rect 1035 727 1036 728
rect 1030 726 1036 727
rect 270 721 276 722
rect 270 717 271 721
rect 275 717 276 721
rect 270 716 276 717
rect 446 721 452 722
rect 446 717 447 721
rect 451 717 452 721
rect 446 716 452 717
rect 638 721 644 722
rect 638 717 639 721
rect 643 717 644 721
rect 638 716 644 717
rect 830 721 836 722
rect 830 717 831 721
rect 835 717 836 721
rect 830 716 836 717
rect 1022 721 1028 722
rect 1022 717 1023 721
rect 1027 717 1028 721
rect 1022 716 1028 717
rect 110 709 116 710
rect 110 705 111 709
rect 115 705 116 709
rect 1110 709 1116 710
rect 430 707 436 708
rect 430 706 431 707
rect 110 704 116 705
rect 325 704 431 706
rect 430 703 431 704
rect 435 703 436 707
rect 582 707 588 708
rect 582 706 583 707
rect 501 704 583 706
rect 430 702 436 703
rect 582 703 583 704
rect 587 703 588 707
rect 750 707 756 708
rect 750 706 751 707
rect 693 704 751 706
rect 582 702 588 703
rect 750 703 751 704
rect 755 703 756 707
rect 1110 705 1111 709
rect 1115 705 1116 709
rect 1110 704 1116 705
rect 750 702 756 703
rect 110 691 116 692
rect 110 687 111 691
rect 115 687 116 691
rect 110 686 116 687
rect 738 691 744 692
rect 738 687 739 691
rect 743 690 744 691
rect 1022 691 1028 692
rect 743 688 841 690
rect 743 687 744 688
rect 738 686 744 687
rect 1022 687 1023 691
rect 1027 690 1028 691
rect 1110 691 1116 692
rect 1027 688 1033 690
rect 1027 687 1028 688
rect 1022 686 1028 687
rect 1110 687 1111 691
rect 1115 687 1116 691
rect 1110 686 1116 687
rect 262 676 268 677
rect 262 672 263 676
rect 267 672 268 676
rect 262 671 268 672
rect 438 676 444 677
rect 438 672 439 676
rect 443 672 444 676
rect 438 671 444 672
rect 630 676 636 677
rect 630 672 631 676
rect 635 672 636 676
rect 630 671 636 672
rect 822 676 828 677
rect 822 672 823 676
rect 827 672 828 676
rect 822 671 828 672
rect 1014 676 1020 677
rect 1014 672 1015 676
rect 1019 672 1020 676
rect 1014 671 1020 672
rect 366 664 372 665
rect 366 660 367 664
rect 371 660 372 664
rect 366 659 372 660
rect 462 664 468 665
rect 462 660 463 664
rect 467 660 468 664
rect 462 659 468 660
rect 558 664 564 665
rect 558 660 559 664
rect 563 660 564 664
rect 558 659 564 660
rect 662 664 668 665
rect 662 660 663 664
rect 667 660 668 664
rect 662 659 668 660
rect 774 664 780 665
rect 774 660 775 664
rect 779 660 780 664
rect 774 659 780 660
rect 894 664 900 665
rect 894 660 895 664
rect 899 660 900 664
rect 894 659 900 660
rect 886 651 892 652
rect 110 649 116 650
rect 110 645 111 649
rect 115 645 116 649
rect 886 647 887 651
rect 891 650 892 651
rect 891 648 913 650
rect 1110 649 1116 650
rect 891 647 892 648
rect 886 646 892 647
rect 110 644 116 645
rect 1110 645 1111 649
rect 1115 645 1116 649
rect 1110 644 1116 645
rect 438 635 444 636
rect 438 634 439 635
rect 429 632 439 634
rect 110 631 116 632
rect 110 627 111 631
rect 115 627 116 631
rect 438 631 439 632
rect 443 631 444 635
rect 534 635 540 636
rect 534 634 535 635
rect 525 632 535 634
rect 438 630 444 631
rect 534 631 535 632
rect 539 631 540 635
rect 638 635 644 636
rect 638 634 639 635
rect 621 632 639 634
rect 534 630 540 631
rect 638 631 639 632
rect 643 631 644 635
rect 746 635 752 636
rect 746 634 747 635
rect 725 632 747 634
rect 638 630 644 631
rect 746 631 747 632
rect 751 631 752 635
rect 746 630 752 631
rect 754 635 760 636
rect 754 631 755 635
rect 759 634 760 635
rect 759 632 801 634
rect 759 631 760 632
rect 754 630 760 631
rect 1110 631 1116 632
rect 110 626 116 627
rect 1110 627 1111 631
rect 1115 627 1116 631
rect 1110 626 1116 627
rect 374 619 380 620
rect 374 615 375 619
rect 379 615 380 619
rect 374 614 380 615
rect 470 619 476 620
rect 470 615 471 619
rect 475 615 476 619
rect 470 614 476 615
rect 566 619 572 620
rect 566 615 567 619
rect 571 615 572 619
rect 566 614 572 615
rect 670 619 676 620
rect 670 615 671 619
rect 675 615 676 619
rect 670 614 676 615
rect 782 619 788 620
rect 782 615 783 619
rect 787 615 788 619
rect 782 614 788 615
rect 902 619 908 620
rect 902 615 903 619
rect 907 615 908 619
rect 902 614 908 615
rect 394 611 400 612
rect 394 607 395 611
rect 399 607 400 611
rect 394 606 400 607
rect 922 611 928 612
rect 922 607 923 611
rect 927 607 928 611
rect 922 606 928 607
rect 438 603 444 604
rect 438 599 439 603
rect 443 602 444 603
rect 488 602 490 605
rect 443 600 490 602
rect 534 603 540 604
rect 443 599 444 600
rect 438 598 444 599
rect 534 599 535 603
rect 539 602 540 603
rect 584 602 586 605
rect 539 600 586 602
rect 638 603 644 604
rect 539 599 540 600
rect 534 598 540 599
rect 638 599 639 603
rect 643 602 644 603
rect 688 602 690 605
rect 643 600 690 602
rect 746 603 752 604
rect 643 599 644 600
rect 638 598 644 599
rect 746 599 747 603
rect 751 602 752 603
rect 800 602 802 605
rect 751 600 802 602
rect 751 599 752 600
rect 746 598 752 599
rect 514 591 520 592
rect 514 587 515 591
rect 519 587 520 591
rect 514 586 520 587
rect 590 591 596 592
rect 590 587 591 591
rect 595 590 596 591
rect 678 591 684 592
rect 595 588 601 590
rect 595 587 596 588
rect 590 586 596 587
rect 678 587 679 591
rect 683 590 684 591
rect 766 591 772 592
rect 683 588 689 590
rect 683 587 684 588
rect 678 586 684 587
rect 766 587 767 591
rect 771 590 772 591
rect 854 591 860 592
rect 771 588 777 590
rect 771 587 772 588
rect 766 586 772 587
rect 854 587 855 591
rect 859 590 860 591
rect 950 591 956 592
rect 859 588 865 590
rect 859 587 860 588
rect 854 586 860 587
rect 950 587 951 591
rect 955 587 956 591
rect 950 586 956 587
rect 1030 591 1036 592
rect 1030 587 1031 591
rect 1035 590 1036 591
rect 1035 588 1041 590
rect 1035 587 1036 588
rect 1030 586 1036 587
rect 494 581 500 582
rect 494 577 495 581
rect 499 577 500 581
rect 494 576 500 577
rect 582 581 588 582
rect 582 577 583 581
rect 587 577 588 581
rect 582 576 588 577
rect 670 581 676 582
rect 670 577 671 581
rect 675 577 676 581
rect 670 576 676 577
rect 758 581 764 582
rect 758 577 759 581
rect 763 577 764 581
rect 758 576 764 577
rect 846 581 852 582
rect 846 577 847 581
rect 851 577 852 581
rect 846 576 852 577
rect 934 581 940 582
rect 934 577 935 581
rect 939 577 940 581
rect 934 576 940 577
rect 1022 581 1028 582
rect 1022 577 1023 581
rect 1027 577 1028 581
rect 1022 576 1028 577
rect 110 569 116 570
rect 110 565 111 569
rect 115 565 116 569
rect 110 564 116 565
rect 1110 569 1116 570
rect 1110 565 1111 569
rect 1115 565 1116 569
rect 1110 564 1116 565
rect 582 563 588 564
rect 582 562 583 563
rect 549 560 583 562
rect 582 559 583 560
rect 587 559 588 563
rect 670 563 676 564
rect 670 562 671 563
rect 637 560 671 562
rect 582 558 588 559
rect 670 559 671 560
rect 675 559 676 563
rect 758 563 764 564
rect 758 562 759 563
rect 725 560 759 562
rect 670 558 676 559
rect 758 559 759 560
rect 763 559 764 563
rect 846 563 852 564
rect 846 562 847 563
rect 813 560 847 562
rect 758 558 764 559
rect 846 559 847 560
rect 851 559 852 563
rect 846 558 852 559
rect 922 563 928 564
rect 922 559 923 563
rect 927 562 928 563
rect 927 560 953 562
rect 927 559 928 560
rect 922 558 928 559
rect 110 551 116 552
rect 110 547 111 551
rect 115 547 116 551
rect 1022 551 1028 552
rect 897 548 910 550
rect 110 546 116 547
rect 906 547 912 548
rect 906 543 907 547
rect 911 543 912 547
rect 1022 547 1023 551
rect 1027 550 1028 551
rect 1110 551 1116 552
rect 1027 548 1033 550
rect 1027 547 1028 548
rect 1022 546 1028 547
rect 1110 547 1111 551
rect 1115 547 1116 551
rect 1110 546 1116 547
rect 906 542 912 543
rect 486 536 492 537
rect 486 532 487 536
rect 491 532 492 536
rect 486 531 492 532
rect 574 536 580 537
rect 574 532 575 536
rect 579 532 580 536
rect 574 531 580 532
rect 662 536 668 537
rect 662 532 663 536
rect 667 532 668 536
rect 662 531 668 532
rect 750 536 756 537
rect 750 532 751 536
rect 755 532 756 536
rect 750 531 756 532
rect 838 536 844 537
rect 838 532 839 536
rect 843 532 844 536
rect 838 531 844 532
rect 926 536 932 537
rect 926 532 927 536
rect 931 532 932 536
rect 926 531 932 532
rect 1014 536 1020 537
rect 1014 532 1015 536
rect 1019 532 1020 536
rect 1014 531 1020 532
rect 446 512 452 513
rect 446 508 447 512
rect 451 508 452 512
rect 446 507 452 508
rect 542 512 548 513
rect 542 508 543 512
rect 547 508 548 512
rect 542 507 548 508
rect 646 512 652 513
rect 646 508 647 512
rect 651 508 652 512
rect 646 507 652 508
rect 758 512 764 513
rect 758 508 759 512
rect 763 508 764 512
rect 758 507 764 508
rect 870 512 876 513
rect 870 508 871 512
rect 875 508 876 512
rect 870 507 876 508
rect 990 512 996 513
rect 990 508 991 512
rect 995 508 996 512
rect 990 507 996 508
rect 110 497 116 498
rect 110 493 111 497
rect 115 493 116 497
rect 110 492 116 493
rect 1110 497 1116 498
rect 1110 493 1111 497
rect 1115 493 1116 497
rect 1110 492 1116 493
rect 550 487 556 488
rect 550 483 551 487
rect 555 483 556 487
rect 998 487 1004 488
rect 550 482 556 483
rect 618 483 624 484
rect 618 482 619 483
rect 509 480 554 482
rect 605 480 619 482
rect 110 479 116 480
rect 110 475 111 479
rect 115 475 116 479
rect 618 479 619 480
rect 623 479 624 483
rect 714 483 720 484
rect 714 482 715 483
rect 709 480 715 482
rect 618 478 624 479
rect 714 479 715 480
rect 719 479 720 483
rect 714 478 720 479
rect 722 483 728 484
rect 722 479 723 483
rect 727 482 728 483
rect 839 483 845 484
rect 727 480 785 482
rect 727 479 728 480
rect 722 478 728 479
rect 839 479 840 483
rect 844 482 845 483
rect 998 483 999 487
rect 1003 483 1004 487
rect 998 482 1004 483
rect 844 480 897 482
rect 1000 480 1017 482
rect 844 479 845 480
rect 839 478 845 479
rect 1110 479 1116 480
rect 110 474 116 475
rect 1110 475 1111 479
rect 1115 475 1116 479
rect 1110 474 1116 475
rect 454 467 460 468
rect 454 463 455 467
rect 459 463 460 467
rect 454 462 460 463
rect 550 467 556 468
rect 550 463 551 467
rect 555 463 556 467
rect 550 462 556 463
rect 654 467 660 468
rect 654 463 655 467
rect 659 463 660 467
rect 654 462 660 463
rect 766 467 772 468
rect 766 463 767 467
rect 771 463 772 467
rect 766 462 772 463
rect 878 467 884 468
rect 878 463 879 467
rect 883 463 884 467
rect 878 462 884 463
rect 998 467 1004 468
rect 998 463 999 467
rect 1003 463 1004 467
rect 998 462 1004 463
rect 474 459 480 460
rect 474 455 475 459
rect 479 455 480 459
rect 474 454 480 455
rect 558 459 564 460
rect 558 455 559 459
rect 563 458 564 459
rect 898 459 904 460
rect 563 456 569 458
rect 563 455 564 456
rect 558 454 564 455
rect 714 455 720 456
rect 714 454 715 455
rect 296 452 446 454
rect 296 447 298 452
rect 444 450 446 452
rect 490 451 496 452
rect 490 450 491 451
rect 444 448 491 450
rect 414 447 420 448
rect 414 443 415 447
rect 419 446 420 447
rect 490 447 491 448
rect 495 447 496 451
rect 618 451 624 452
rect 490 446 496 447
rect 562 447 568 448
rect 419 444 425 446
rect 419 443 420 444
rect 414 442 420 443
rect 562 443 563 447
rect 567 443 568 447
rect 618 447 619 451
rect 623 450 624 451
rect 672 450 674 453
rect 623 448 674 450
rect 704 452 715 454
rect 623 447 624 448
rect 704 447 706 452
rect 714 451 715 452
rect 719 451 720 455
rect 839 455 845 456
rect 839 454 840 455
rect 714 450 720 451
rect 784 450 786 453
rect 804 452 840 454
rect 804 450 806 452
rect 839 451 840 452
rect 844 451 845 455
rect 898 455 899 459
rect 903 455 904 459
rect 898 454 904 455
rect 1018 459 1024 460
rect 1018 455 1019 459
rect 1023 455 1024 459
rect 1018 454 1024 455
rect 839 450 845 451
rect 784 448 806 450
rect 858 447 864 448
rect 618 446 624 447
rect 562 442 568 443
rect 858 443 859 447
rect 863 443 864 447
rect 858 442 864 443
rect 1006 447 1012 448
rect 1006 443 1007 447
rect 1011 446 1012 447
rect 1011 444 1017 446
rect 1011 443 1012 444
rect 1006 442 1012 443
rect 278 437 284 438
rect 278 433 279 437
rect 283 433 284 437
rect 278 432 284 433
rect 406 437 412 438
rect 406 433 407 437
rect 411 433 412 437
rect 406 432 412 433
rect 542 437 548 438
rect 542 433 543 437
rect 547 433 548 437
rect 542 432 548 433
rect 686 437 692 438
rect 686 433 687 437
rect 691 433 692 437
rect 686 432 692 433
rect 838 437 844 438
rect 838 433 839 437
rect 843 433 844 437
rect 838 432 844 433
rect 998 437 1004 438
rect 998 433 999 437
rect 1003 433 1004 437
rect 998 432 1004 433
rect 110 425 116 426
rect 110 421 111 425
rect 115 421 116 425
rect 1110 425 1116 426
rect 950 423 956 424
rect 950 422 951 423
rect 110 420 116 421
rect 893 420 951 422
rect 406 419 412 420
rect 406 418 407 419
rect 333 416 407 418
rect 406 415 407 416
rect 411 415 412 419
rect 406 414 412 415
rect 490 419 496 420
rect 490 415 491 419
rect 495 418 496 419
rect 610 419 616 420
rect 495 416 561 418
rect 495 415 496 416
rect 490 414 496 415
rect 610 415 611 419
rect 615 418 616 419
rect 950 419 951 420
rect 955 419 956 423
rect 1110 421 1111 425
rect 1115 421 1116 425
rect 1110 420 1116 421
rect 950 418 956 419
rect 615 416 705 418
rect 615 415 616 416
rect 610 414 616 415
rect 110 407 116 408
rect 110 403 111 407
rect 115 403 116 407
rect 502 407 508 408
rect 502 406 503 407
rect 457 404 503 406
rect 110 402 116 403
rect 502 403 503 404
rect 507 403 508 407
rect 502 402 508 403
rect 998 407 1004 408
rect 998 403 999 407
rect 1003 406 1004 407
rect 1110 407 1116 408
rect 1003 404 1009 406
rect 1003 403 1004 404
rect 998 402 1004 403
rect 1110 403 1111 407
rect 1115 403 1116 407
rect 1110 402 1116 403
rect 270 392 276 393
rect 270 388 271 392
rect 275 388 276 392
rect 270 387 276 388
rect 398 392 404 393
rect 398 388 399 392
rect 403 388 404 392
rect 398 387 404 388
rect 534 392 540 393
rect 534 388 535 392
rect 539 388 540 392
rect 534 387 540 388
rect 678 392 684 393
rect 678 388 679 392
rect 683 388 684 392
rect 678 387 684 388
rect 830 392 836 393
rect 830 388 831 392
rect 835 388 836 392
rect 830 387 836 388
rect 990 392 996 393
rect 990 388 991 392
rect 995 388 996 392
rect 990 387 996 388
rect 162 383 168 384
rect 134 380 140 381
rect 134 376 135 380
rect 139 376 140 380
rect 162 379 163 383
rect 167 382 168 383
rect 167 380 206 382
rect 167 379 168 380
rect 162 378 168 379
rect 134 375 140 376
rect 204 366 206 380
rect 286 380 292 381
rect 286 376 287 380
rect 291 376 292 380
rect 286 375 292 376
rect 478 380 484 381
rect 478 376 479 380
rect 483 376 484 380
rect 478 375 484 376
rect 670 380 676 381
rect 670 376 671 380
rect 675 376 676 380
rect 670 375 676 376
rect 870 380 876 381
rect 870 376 871 380
rect 875 376 876 380
rect 870 375 876 376
rect 858 367 864 368
rect 110 365 116 366
rect 110 361 111 365
rect 115 361 116 365
rect 204 364 305 366
rect 537 364 682 366
rect 110 360 116 361
rect 678 363 684 364
rect 678 359 679 363
rect 683 359 684 363
rect 858 363 859 367
rect 863 366 864 367
rect 863 364 889 366
rect 1110 365 1116 366
rect 863 363 864 364
rect 858 362 864 363
rect 1110 361 1111 365
rect 1115 361 1116 365
rect 1110 360 1116 361
rect 678 358 684 359
rect 142 355 148 356
rect 142 351 143 355
rect 147 351 148 355
rect 142 350 148 351
rect 558 351 564 352
rect 144 348 161 350
rect 110 347 116 348
rect 110 343 111 347
rect 115 343 116 347
rect 558 347 559 351
rect 563 350 564 351
rect 563 348 697 350
rect 563 347 564 348
rect 558 346 564 347
rect 1110 347 1116 348
rect 110 342 116 343
rect 1110 343 1111 347
rect 1115 343 1116 347
rect 1110 342 1116 343
rect 142 335 148 336
rect 142 331 143 335
rect 147 331 148 335
rect 142 330 148 331
rect 294 335 300 336
rect 294 331 295 335
rect 299 331 300 335
rect 294 330 300 331
rect 486 335 492 336
rect 486 331 487 335
rect 491 331 492 335
rect 486 330 492 331
rect 678 335 684 336
rect 678 331 679 335
rect 683 331 684 335
rect 678 330 684 331
rect 878 335 884 336
rect 878 331 879 335
rect 883 331 884 335
rect 878 330 884 331
rect 162 327 168 328
rect 162 323 163 327
rect 167 323 168 327
rect 162 322 168 323
rect 314 327 320 328
rect 314 323 315 327
rect 319 323 320 327
rect 314 322 320 323
rect 502 327 508 328
rect 502 323 503 327
rect 507 323 508 327
rect 502 322 508 323
rect 686 327 692 328
rect 686 323 687 327
rect 691 326 692 327
rect 894 327 900 328
rect 691 324 697 326
rect 691 323 692 324
rect 686 322 692 323
rect 894 323 895 327
rect 899 323 900 327
rect 894 322 900 323
rect 998 327 1004 328
rect 998 323 999 327
rect 1003 326 1004 327
rect 1003 324 1034 326
rect 1003 323 1004 324
rect 998 322 1004 323
rect 150 319 156 320
rect 150 315 151 319
rect 155 318 156 319
rect 462 319 468 320
rect 155 316 161 318
rect 155 315 156 316
rect 150 314 156 315
rect 286 315 292 316
rect 462 315 463 319
rect 467 318 468 319
rect 646 319 652 320
rect 467 316 473 318
rect 467 315 468 316
rect 286 311 287 315
rect 291 314 292 315
rect 296 314 298 315
rect 462 314 468 315
rect 646 315 647 319
rect 651 318 652 319
rect 842 319 848 320
rect 1032 319 1034 324
rect 651 316 657 318
rect 651 315 652 316
rect 646 314 652 315
rect 842 315 843 319
rect 847 315 848 319
rect 842 314 848 315
rect 291 312 298 314
rect 291 311 292 312
rect 286 310 292 311
rect 142 309 148 310
rect 142 305 143 309
rect 147 305 148 309
rect 142 304 148 305
rect 278 309 284 310
rect 278 305 279 309
rect 283 305 284 309
rect 278 304 284 305
rect 454 309 460 310
rect 454 305 455 309
rect 459 305 460 309
rect 454 304 460 305
rect 638 309 644 310
rect 638 305 639 309
rect 643 305 644 309
rect 638 304 644 305
rect 822 309 828 310
rect 822 305 823 309
rect 827 305 828 309
rect 822 304 828 305
rect 1014 309 1020 310
rect 1014 305 1015 309
rect 1019 305 1020 309
rect 1014 304 1020 305
rect 110 297 116 298
rect 110 293 111 297
rect 115 293 116 297
rect 1110 297 1116 298
rect 894 295 900 296
rect 894 294 895 295
rect 110 292 116 293
rect 877 292 895 294
rect 278 291 284 292
rect 278 290 279 291
rect 197 288 279 290
rect 278 287 279 288
rect 283 287 284 291
rect 454 291 460 292
rect 454 290 455 291
rect 333 288 455 290
rect 278 286 284 287
rect 454 287 455 288
rect 459 287 460 291
rect 638 291 644 292
rect 638 290 639 291
rect 509 288 639 290
rect 454 286 460 287
rect 638 287 639 288
rect 643 287 644 291
rect 894 291 895 292
rect 899 291 900 295
rect 1110 293 1111 297
rect 1115 293 1116 297
rect 1110 292 1116 293
rect 894 290 900 291
rect 638 286 644 287
rect 110 279 116 280
rect 110 275 111 279
rect 115 275 116 279
rect 110 274 116 275
rect 570 279 576 280
rect 570 275 571 279
rect 575 278 576 279
rect 938 279 944 280
rect 575 276 649 278
rect 575 275 576 276
rect 570 274 576 275
rect 938 275 939 279
rect 943 278 944 279
rect 1110 279 1116 280
rect 943 276 1025 278
rect 943 275 944 276
rect 938 274 944 275
rect 1110 275 1111 279
rect 1115 275 1116 279
rect 1110 274 1116 275
rect 134 264 140 265
rect 134 260 135 264
rect 139 260 140 264
rect 134 259 140 260
rect 270 264 276 265
rect 270 260 271 264
rect 275 260 276 264
rect 270 259 276 260
rect 446 264 452 265
rect 446 260 447 264
rect 451 260 452 264
rect 446 259 452 260
rect 630 264 636 265
rect 630 260 631 264
rect 635 260 636 264
rect 630 259 636 260
rect 814 264 820 265
rect 814 260 815 264
rect 819 260 820 264
rect 814 259 820 260
rect 1006 264 1012 265
rect 1006 260 1007 264
rect 1011 260 1012 264
rect 1006 259 1012 260
rect 294 244 300 245
rect 294 240 295 244
rect 299 240 300 244
rect 294 239 300 240
rect 422 244 428 245
rect 422 240 423 244
rect 427 240 428 244
rect 422 239 428 240
rect 542 244 548 245
rect 542 240 543 244
rect 547 240 548 244
rect 542 239 548 240
rect 662 244 668 245
rect 662 240 663 244
rect 667 240 668 244
rect 662 239 668 240
rect 782 244 788 245
rect 782 240 783 244
rect 787 240 788 244
rect 782 239 788 240
rect 910 244 916 245
rect 910 240 911 244
rect 915 240 916 244
rect 910 239 916 240
rect 1014 244 1020 245
rect 1014 240 1015 244
rect 1019 240 1020 244
rect 1014 239 1020 240
rect 110 229 116 230
rect 110 225 111 229
rect 115 225 116 229
rect 110 224 116 225
rect 1110 229 1116 230
rect 1110 225 1111 229
rect 1115 225 1116 229
rect 1110 224 1116 225
rect 362 215 368 216
rect 362 214 363 215
rect 357 212 363 214
rect 110 211 116 212
rect 110 207 111 211
rect 115 207 116 211
rect 362 211 363 212
rect 367 211 368 215
rect 362 210 368 211
rect 382 215 388 216
rect 382 211 383 215
rect 387 214 388 215
rect 506 215 512 216
rect 387 212 449 214
rect 387 211 388 212
rect 382 210 388 211
rect 506 211 507 215
rect 511 214 512 215
rect 746 215 752 216
rect 746 214 747 215
rect 511 212 569 214
rect 725 212 747 214
rect 511 211 512 212
rect 506 210 512 211
rect 746 211 747 212
rect 751 211 752 215
rect 850 215 856 216
rect 850 214 851 215
rect 845 212 851 214
rect 746 210 752 211
rect 850 211 851 212
rect 855 211 856 215
rect 986 215 992 216
rect 986 214 987 215
rect 973 212 987 214
rect 850 210 856 211
rect 986 211 987 212
rect 991 211 992 215
rect 1082 215 1088 216
rect 1082 214 1083 215
rect 1077 212 1083 214
rect 986 210 992 211
rect 1082 211 1083 212
rect 1087 211 1088 215
rect 1082 210 1088 211
rect 1110 211 1116 212
rect 110 206 116 207
rect 1110 207 1111 211
rect 1115 207 1116 211
rect 1110 206 1116 207
rect 302 199 308 200
rect 302 195 303 199
rect 307 195 308 199
rect 302 194 308 195
rect 430 199 436 200
rect 430 195 431 199
rect 435 195 436 199
rect 430 194 436 195
rect 550 199 556 200
rect 550 195 551 199
rect 555 195 556 199
rect 550 194 556 195
rect 670 199 676 200
rect 670 195 671 199
rect 675 195 676 199
rect 670 194 676 195
rect 790 199 796 200
rect 790 195 791 199
rect 795 195 796 199
rect 790 194 796 195
rect 918 199 924 200
rect 918 195 919 199
rect 923 195 924 199
rect 918 194 924 195
rect 1022 199 1028 200
rect 1022 195 1023 199
rect 1027 195 1028 199
rect 1022 194 1028 195
rect 570 191 576 192
rect 570 187 571 191
rect 575 187 576 191
rect 570 186 576 187
rect 938 191 944 192
rect 938 187 939 191
rect 943 187 944 191
rect 938 186 944 187
rect 320 182 322 185
rect 382 183 388 184
rect 382 182 383 183
rect 320 180 383 182
rect 382 179 383 180
rect 387 179 388 183
rect 448 182 450 185
rect 506 183 512 184
rect 506 182 507 183
rect 448 180 507 182
rect 382 178 388 179
rect 506 179 507 180
rect 511 179 512 183
rect 506 178 512 179
rect 362 175 368 176
rect 362 174 363 175
rect 336 172 363 174
rect 336 167 338 172
rect 362 171 363 172
rect 367 171 368 175
rect 688 174 690 185
rect 746 183 752 184
rect 746 179 747 183
rect 751 182 752 183
rect 808 182 810 185
rect 751 180 810 182
rect 986 183 992 184
rect 751 179 752 180
rect 746 178 752 179
rect 986 179 987 183
rect 991 182 992 183
rect 1040 182 1042 185
rect 991 180 1042 182
rect 991 179 992 180
rect 986 178 992 179
rect 826 175 832 176
rect 826 174 827 175
rect 688 172 827 174
rect 362 170 368 171
rect 826 171 827 172
rect 831 171 832 175
rect 1002 175 1008 176
rect 1002 174 1003 175
rect 826 170 832 171
rect 952 172 1003 174
rect 414 167 420 168
rect 414 163 415 167
rect 419 166 420 167
rect 502 167 508 168
rect 419 164 425 166
rect 419 163 420 164
rect 414 162 420 163
rect 502 163 503 167
rect 507 166 508 167
rect 590 167 596 168
rect 507 164 513 166
rect 507 163 508 164
rect 502 162 508 163
rect 590 163 591 167
rect 595 166 596 167
rect 678 167 684 168
rect 595 164 601 166
rect 595 163 596 164
rect 590 162 596 163
rect 678 163 679 167
rect 683 166 684 167
rect 766 167 772 168
rect 683 164 689 166
rect 683 163 684 164
rect 678 162 684 163
rect 766 163 767 167
rect 771 166 772 167
rect 854 167 860 168
rect 952 167 954 172
rect 1002 171 1003 172
rect 1007 171 1008 175
rect 1082 175 1088 176
rect 1082 174 1083 175
rect 1002 170 1008 171
rect 1040 172 1083 174
rect 1040 167 1042 172
rect 1082 171 1083 172
rect 1087 171 1088 175
rect 1082 170 1088 171
rect 771 164 777 166
rect 771 163 772 164
rect 766 162 772 163
rect 854 163 855 167
rect 859 166 860 167
rect 859 164 865 166
rect 859 163 860 164
rect 854 162 860 163
rect 318 157 324 158
rect 318 153 319 157
rect 323 153 324 157
rect 318 152 324 153
rect 406 157 412 158
rect 406 153 407 157
rect 411 153 412 157
rect 406 152 412 153
rect 494 157 500 158
rect 494 153 495 157
rect 499 153 500 157
rect 494 152 500 153
rect 582 157 588 158
rect 582 153 583 157
rect 587 153 588 157
rect 582 152 588 153
rect 670 157 676 158
rect 670 153 671 157
rect 675 153 676 157
rect 670 152 676 153
rect 758 157 764 158
rect 758 153 759 157
rect 763 153 764 157
rect 758 152 764 153
rect 846 157 852 158
rect 846 153 847 157
rect 851 153 852 157
rect 846 152 852 153
rect 934 157 940 158
rect 934 153 935 157
rect 939 153 940 157
rect 934 152 940 153
rect 1022 157 1028 158
rect 1022 153 1023 157
rect 1027 153 1028 157
rect 1022 152 1028 153
rect 110 145 116 146
rect 110 141 111 145
rect 115 141 116 145
rect 110 140 116 141
rect 1110 145 1116 146
rect 1110 141 1111 145
rect 1115 141 1116 145
rect 1110 140 1116 141
rect 406 139 412 140
rect 406 138 407 139
rect 373 136 407 138
rect 406 135 407 136
rect 411 135 412 139
rect 494 139 500 140
rect 494 138 495 139
rect 461 136 495 138
rect 406 134 412 135
rect 494 135 495 136
rect 499 135 500 139
rect 582 139 588 140
rect 582 138 583 139
rect 549 136 583 138
rect 494 134 500 135
rect 582 135 583 136
rect 587 135 588 139
rect 670 139 676 140
rect 670 138 671 139
rect 637 136 671 138
rect 582 134 588 135
rect 670 135 671 136
rect 675 135 676 139
rect 758 139 764 140
rect 758 138 759 139
rect 725 136 759 138
rect 670 134 676 135
rect 758 135 759 136
rect 763 135 764 139
rect 846 139 852 140
rect 846 138 847 139
rect 813 136 847 138
rect 758 134 764 135
rect 846 135 847 136
rect 851 135 852 139
rect 846 134 852 135
rect 1002 139 1008 140
rect 1002 135 1003 139
rect 1007 138 1008 139
rect 1007 136 1041 138
rect 1007 135 1008 136
rect 1002 134 1008 135
rect 110 127 116 128
rect 110 123 111 127
rect 115 123 116 127
rect 110 122 116 123
rect 826 127 832 128
rect 826 123 827 127
rect 831 126 832 127
rect 1110 127 1116 128
rect 831 124 857 126
rect 831 123 832 124
rect 826 122 832 123
rect 1110 123 1111 127
rect 1115 123 1116 127
rect 1110 122 1116 123
rect 310 112 316 113
rect 310 108 311 112
rect 315 108 316 112
rect 310 107 316 108
rect 398 112 404 113
rect 398 108 399 112
rect 403 108 404 112
rect 398 107 404 108
rect 486 112 492 113
rect 486 108 487 112
rect 491 108 492 112
rect 486 107 492 108
rect 574 112 580 113
rect 574 108 575 112
rect 579 108 580 112
rect 574 107 580 108
rect 662 112 668 113
rect 662 108 663 112
rect 667 108 668 112
rect 662 107 668 108
rect 750 112 756 113
rect 750 108 751 112
rect 755 108 756 112
rect 750 107 756 108
rect 838 112 844 113
rect 838 108 839 112
rect 843 108 844 112
rect 838 107 844 108
rect 926 112 932 113
rect 926 108 927 112
rect 931 108 932 112
rect 926 107 932 108
rect 1014 112 1020 113
rect 1014 108 1015 112
rect 1019 108 1020 112
rect 1014 107 1020 108
<< m3c >>
rect 135 1212 139 1216
rect 223 1212 227 1216
rect 311 1212 315 1216
rect 111 1197 115 1201
rect 1111 1197 1115 1201
rect 111 1179 115 1183
rect 143 1167 147 1171
rect 163 1159 167 1163
rect 203 1183 207 1187
rect 291 1183 295 1187
rect 1111 1179 1115 1183
rect 231 1167 235 1171
rect 319 1167 323 1171
rect 251 1159 255 1163
rect 411 1159 415 1163
rect 271 1151 275 1155
rect 359 1151 363 1155
rect 175 1141 179 1145
rect 263 1141 267 1145
rect 351 1141 355 1145
rect 439 1141 443 1145
rect 111 1129 115 1133
rect 259 1123 263 1127
rect 347 1123 351 1127
rect 411 1127 415 1131
rect 1111 1129 1115 1133
rect 111 1111 115 1115
rect 423 1111 427 1115
rect 1111 1111 1115 1115
rect 167 1096 171 1100
rect 255 1096 259 1100
rect 343 1096 347 1100
rect 431 1096 435 1100
rect 399 1084 403 1088
rect 487 1084 491 1088
rect 575 1084 579 1088
rect 663 1084 667 1088
rect 751 1084 755 1088
rect 839 1084 843 1088
rect 927 1084 931 1088
rect 955 1087 959 1091
rect 1015 1084 1019 1088
rect 111 1069 115 1073
rect 1111 1069 1115 1073
rect 495 1059 499 1063
rect 583 1059 587 1063
rect 671 1059 675 1063
rect 111 1051 115 1055
rect 743 1055 747 1059
rect 759 1059 763 1063
rect 935 1059 939 1063
rect 1023 1059 1027 1063
rect 1111 1051 1115 1055
rect 407 1039 411 1043
rect 495 1039 499 1043
rect 583 1039 587 1043
rect 671 1039 675 1043
rect 759 1039 763 1043
rect 847 1039 851 1043
rect 935 1039 939 1043
rect 1023 1039 1027 1043
rect 423 1031 427 1035
rect 503 1031 507 1035
rect 591 1031 595 1035
rect 679 1031 683 1035
rect 775 1031 779 1035
rect 855 1031 859 1035
rect 943 1031 947 1035
rect 1031 1031 1035 1035
rect 503 1023 507 1027
rect 415 1019 419 1023
rect 591 1023 595 1027
rect 767 1023 771 1027
rect 679 1019 683 1023
rect 863 1021 867 1025
rect 955 1021 959 1025
rect 1031 1023 1035 1027
rect 407 1013 411 1017
rect 495 1013 499 1017
rect 583 1013 587 1017
rect 671 1013 675 1017
rect 759 1013 763 1017
rect 847 1013 851 1017
rect 935 1013 939 1017
rect 1023 1013 1027 1017
rect 111 1001 115 1005
rect 1111 1001 1115 1005
rect 491 995 495 999
rect 579 995 583 999
rect 651 995 655 999
rect 739 995 743 999
rect 847 995 851 999
rect 1019 995 1023 999
rect 111 983 115 987
rect 671 983 675 987
rect 1023 983 1027 987
rect 1111 983 1115 987
rect 399 968 403 972
rect 487 968 491 972
rect 575 968 579 972
rect 663 968 667 972
rect 751 968 755 972
rect 839 968 843 972
rect 927 968 931 972
rect 1015 968 1019 972
rect 151 940 155 944
rect 271 940 275 944
rect 407 940 411 944
rect 551 940 555 944
rect 711 940 715 944
rect 871 940 875 944
rect 1015 940 1019 944
rect 111 925 115 929
rect 863 927 867 931
rect 1111 925 1115 929
rect 111 907 115 911
rect 371 911 375 915
rect 503 911 507 915
rect 655 911 659 915
rect 1083 911 1087 915
rect 1111 907 1115 911
rect 159 895 163 899
rect 279 895 283 899
rect 415 895 419 899
rect 559 895 563 899
rect 719 895 723 899
rect 879 895 883 899
rect 1023 895 1027 899
rect 1031 887 1035 891
rect 219 879 223 883
rect 371 879 375 883
rect 503 879 507 883
rect 655 879 659 883
rect 671 879 675 883
rect 755 879 759 883
rect 447 871 451 875
rect 931 879 935 883
rect 1083 879 1087 883
rect 639 871 643 875
rect 143 861 147 865
rect 271 861 275 865
rect 439 861 443 865
rect 631 861 635 865
rect 839 861 843 865
rect 1023 861 1027 865
rect 111 849 115 853
rect 219 847 223 851
rect 435 843 439 847
rect 627 843 631 847
rect 755 847 759 851
rect 1111 849 1115 853
rect 111 831 115 835
rect 739 831 743 835
rect 1023 831 1027 835
rect 1111 831 1115 835
rect 135 816 139 820
rect 263 816 267 820
rect 431 816 435 820
rect 623 816 627 820
rect 831 816 835 820
rect 1015 816 1019 820
rect 135 792 139 796
rect 239 792 243 796
rect 375 792 379 796
rect 527 792 531 796
rect 695 792 699 796
rect 863 792 867 796
rect 1015 792 1019 796
rect 111 777 115 781
rect 931 779 935 783
rect 1111 777 1115 781
rect 111 759 115 763
rect 211 763 215 767
rect 483 763 487 767
rect 675 763 679 767
rect 683 763 687 767
rect 1023 767 1027 771
rect 1111 759 1115 763
rect 143 747 147 751
rect 247 747 251 751
rect 383 747 387 751
rect 535 747 539 751
rect 703 747 707 751
rect 871 747 875 751
rect 1023 747 1027 751
rect 163 739 167 743
rect 211 731 215 735
rect 291 727 295 731
rect 431 735 435 739
rect 483 731 487 735
rect 583 735 587 739
rect 675 731 679 735
rect 751 735 755 739
rect 887 739 891 743
rect 1039 739 1043 743
rect 1031 727 1035 731
rect 271 717 275 721
rect 447 717 451 721
rect 639 717 643 721
rect 831 717 835 721
rect 1023 717 1027 721
rect 111 705 115 709
rect 431 703 435 707
rect 583 703 587 707
rect 751 703 755 707
rect 1111 705 1115 709
rect 111 687 115 691
rect 739 687 743 691
rect 1023 687 1027 691
rect 1111 687 1115 691
rect 263 672 267 676
rect 439 672 443 676
rect 631 672 635 676
rect 823 672 827 676
rect 1015 672 1019 676
rect 367 660 371 664
rect 463 660 467 664
rect 559 660 563 664
rect 663 660 667 664
rect 775 660 779 664
rect 895 660 899 664
rect 111 645 115 649
rect 887 647 891 651
rect 1111 645 1115 649
rect 111 627 115 631
rect 439 631 443 635
rect 535 631 539 635
rect 639 631 643 635
rect 747 631 751 635
rect 755 631 759 635
rect 1111 627 1115 631
rect 375 615 379 619
rect 471 615 475 619
rect 567 615 571 619
rect 671 615 675 619
rect 783 615 787 619
rect 903 615 907 619
rect 395 607 399 611
rect 923 607 927 611
rect 439 599 443 603
rect 535 599 539 603
rect 639 599 643 603
rect 747 599 751 603
rect 515 587 519 591
rect 591 587 595 591
rect 679 587 683 591
rect 767 587 771 591
rect 855 587 859 591
rect 951 587 955 591
rect 1031 587 1035 591
rect 495 577 499 581
rect 583 577 587 581
rect 671 577 675 581
rect 759 577 763 581
rect 847 577 851 581
rect 935 577 939 581
rect 1023 577 1027 581
rect 111 565 115 569
rect 1111 565 1115 569
rect 583 559 587 563
rect 671 559 675 563
rect 759 559 763 563
rect 847 559 851 563
rect 923 559 927 563
rect 111 547 115 551
rect 907 543 911 547
rect 1023 547 1027 551
rect 1111 547 1115 551
rect 487 532 491 536
rect 575 532 579 536
rect 663 532 667 536
rect 751 532 755 536
rect 839 532 843 536
rect 927 532 931 536
rect 1015 532 1019 536
rect 447 508 451 512
rect 543 508 547 512
rect 647 508 651 512
rect 759 508 763 512
rect 871 508 875 512
rect 991 508 995 512
rect 111 493 115 497
rect 1111 493 1115 497
rect 551 483 555 487
rect 111 475 115 479
rect 619 479 623 483
rect 715 479 719 483
rect 723 479 727 483
rect 999 483 1003 487
rect 1111 475 1115 479
rect 455 463 459 467
rect 551 463 555 467
rect 655 463 659 467
rect 767 463 771 467
rect 879 463 883 467
rect 999 463 1003 467
rect 475 455 479 459
rect 559 455 563 459
rect 415 443 419 447
rect 491 447 495 451
rect 563 443 567 447
rect 619 447 623 451
rect 715 451 719 455
rect 899 455 903 459
rect 1019 455 1023 459
rect 859 443 863 447
rect 1007 443 1011 447
rect 279 433 283 437
rect 407 433 411 437
rect 543 433 547 437
rect 687 433 691 437
rect 839 433 843 437
rect 999 433 1003 437
rect 111 421 115 425
rect 407 415 411 419
rect 491 415 495 419
rect 611 415 615 419
rect 951 419 955 423
rect 1111 421 1115 425
rect 111 403 115 407
rect 503 403 507 407
rect 999 403 1003 407
rect 1111 403 1115 407
rect 271 388 275 392
rect 399 388 403 392
rect 535 388 539 392
rect 679 388 683 392
rect 831 388 835 392
rect 991 388 995 392
rect 135 376 139 380
rect 163 379 167 383
rect 287 376 291 380
rect 479 376 483 380
rect 671 376 675 380
rect 871 376 875 380
rect 111 361 115 365
rect 679 359 683 363
rect 859 363 863 367
rect 1111 361 1115 365
rect 143 351 147 355
rect 111 343 115 347
rect 559 347 563 351
rect 1111 343 1115 347
rect 143 331 147 335
rect 295 331 299 335
rect 487 331 491 335
rect 679 331 683 335
rect 879 331 883 335
rect 163 323 167 327
rect 315 323 319 327
rect 503 323 507 327
rect 687 323 691 327
rect 895 323 899 327
rect 999 323 1003 327
rect 151 315 155 319
rect 463 315 467 319
rect 287 311 291 315
rect 647 315 651 319
rect 843 315 847 319
rect 143 305 147 309
rect 279 305 283 309
rect 455 305 459 309
rect 639 305 643 309
rect 823 305 827 309
rect 1015 305 1019 309
rect 111 293 115 297
rect 279 287 283 291
rect 455 287 459 291
rect 639 287 643 291
rect 895 291 899 295
rect 1111 293 1115 297
rect 111 275 115 279
rect 571 275 575 279
rect 939 275 943 279
rect 1111 275 1115 279
rect 135 260 139 264
rect 271 260 275 264
rect 447 260 451 264
rect 631 260 635 264
rect 815 260 819 264
rect 1007 260 1011 264
rect 295 240 299 244
rect 423 240 427 244
rect 543 240 547 244
rect 663 240 667 244
rect 783 240 787 244
rect 911 240 915 244
rect 1015 240 1019 244
rect 111 225 115 229
rect 1111 225 1115 229
rect 111 207 115 211
rect 363 211 367 215
rect 383 211 387 215
rect 507 211 511 215
rect 747 211 751 215
rect 851 211 855 215
rect 987 211 991 215
rect 1083 211 1087 215
rect 1111 207 1115 211
rect 303 195 307 199
rect 431 195 435 199
rect 551 195 555 199
rect 671 195 675 199
rect 791 195 795 199
rect 919 195 923 199
rect 1023 195 1027 199
rect 571 187 575 191
rect 939 187 943 191
rect 383 179 387 183
rect 507 179 511 183
rect 363 171 367 175
rect 747 179 751 183
rect 987 179 991 183
rect 827 171 831 175
rect 415 163 419 167
rect 503 163 507 167
rect 591 163 595 167
rect 679 163 683 167
rect 767 163 771 167
rect 1003 171 1007 175
rect 1083 171 1087 175
rect 855 163 859 167
rect 319 153 323 157
rect 407 153 411 157
rect 495 153 499 157
rect 583 153 587 157
rect 671 153 675 157
rect 759 153 763 157
rect 847 153 851 157
rect 935 153 939 157
rect 1023 153 1027 157
rect 111 141 115 145
rect 1111 141 1115 145
rect 407 135 411 139
rect 495 135 499 139
rect 583 135 587 139
rect 671 135 675 139
rect 759 135 763 139
rect 847 135 851 139
rect 1003 135 1007 139
rect 111 123 115 127
rect 827 123 831 127
rect 1111 123 1115 127
rect 311 108 315 112
rect 399 108 403 112
rect 487 108 491 112
rect 575 108 579 112
rect 663 108 667 112
rect 751 108 755 112
rect 839 108 843 112
rect 927 108 931 112
rect 1015 108 1019 112
<< m3 >>
rect 111 1222 115 1223
rect 111 1217 115 1218
rect 135 1222 139 1223
rect 135 1217 139 1218
rect 223 1222 227 1223
rect 223 1217 227 1218
rect 311 1222 315 1223
rect 311 1217 315 1218
rect 1111 1222 1115 1223
rect 1111 1217 1115 1218
rect 112 1202 114 1217
rect 134 1216 140 1217
rect 134 1212 135 1216
rect 139 1212 140 1216
rect 134 1211 140 1212
rect 222 1216 228 1217
rect 222 1212 223 1216
rect 227 1212 228 1216
rect 222 1211 228 1212
rect 310 1216 316 1217
rect 310 1212 311 1216
rect 315 1212 316 1216
rect 310 1211 316 1212
rect 1112 1202 1114 1217
rect 110 1201 116 1202
rect 110 1197 111 1201
rect 115 1197 116 1201
rect 110 1196 116 1197
rect 1110 1201 1116 1202
rect 1110 1197 1111 1201
rect 1115 1197 1116 1201
rect 1110 1196 1116 1197
rect 202 1187 208 1188
rect 110 1183 116 1184
rect 110 1179 111 1183
rect 115 1179 116 1183
rect 202 1183 203 1187
rect 207 1183 208 1187
rect 202 1182 208 1183
rect 290 1187 296 1188
rect 290 1183 291 1187
rect 295 1183 296 1187
rect 290 1182 296 1183
rect 1110 1183 1116 1184
rect 110 1178 116 1179
rect 112 1159 114 1178
rect 204 1173 206 1182
rect 292 1173 294 1182
rect 1110 1179 1111 1183
rect 1115 1179 1116 1183
rect 1110 1178 1116 1179
rect 163 1172 167 1173
rect 142 1171 148 1172
rect 142 1167 143 1171
rect 147 1167 148 1171
rect 163 1167 167 1168
rect 203 1172 207 1173
rect 251 1172 255 1173
rect 203 1167 207 1168
rect 230 1171 236 1172
rect 230 1167 231 1171
rect 235 1167 236 1171
rect 251 1167 255 1168
rect 291 1172 295 1173
rect 291 1167 295 1168
rect 318 1171 324 1172
rect 318 1167 319 1171
rect 323 1167 324 1171
rect 142 1166 148 1167
rect 144 1159 146 1166
rect 164 1164 166 1167
rect 230 1166 236 1167
rect 162 1163 168 1164
rect 162 1159 163 1163
rect 167 1159 168 1163
rect 232 1159 234 1166
rect 252 1164 254 1167
rect 318 1166 324 1167
rect 250 1163 256 1164
rect 250 1159 251 1163
rect 255 1159 256 1163
rect 320 1159 322 1166
rect 410 1163 416 1164
rect 410 1159 411 1163
rect 415 1159 416 1163
rect 1112 1159 1114 1178
rect 111 1158 115 1159
rect 111 1153 115 1154
rect 143 1158 147 1159
rect 162 1158 168 1159
rect 175 1158 179 1159
rect 143 1153 147 1154
rect 175 1153 179 1154
rect 231 1158 235 1159
rect 250 1158 256 1159
rect 263 1158 267 1159
rect 231 1153 235 1154
rect 319 1158 323 1159
rect 263 1153 267 1154
rect 270 1155 276 1156
rect 112 1134 114 1153
rect 176 1146 178 1153
rect 264 1146 266 1153
rect 270 1151 271 1155
rect 275 1151 276 1155
rect 319 1153 323 1154
rect 351 1158 355 1159
rect 410 1158 416 1159
rect 439 1158 443 1159
rect 351 1153 355 1154
rect 358 1155 364 1156
rect 270 1150 276 1151
rect 174 1145 180 1146
rect 174 1141 175 1145
rect 179 1141 180 1145
rect 174 1140 180 1141
rect 262 1145 268 1146
rect 262 1141 263 1145
rect 267 1141 268 1145
rect 262 1140 268 1141
rect 110 1133 116 1134
rect 110 1129 111 1133
rect 115 1129 116 1133
rect 110 1128 116 1129
rect 258 1127 264 1128
rect 258 1123 259 1127
rect 263 1123 264 1127
rect 272 1123 274 1150
rect 352 1146 354 1153
rect 358 1151 359 1155
rect 363 1151 364 1155
rect 358 1150 364 1151
rect 350 1145 356 1146
rect 350 1141 351 1145
rect 355 1141 356 1145
rect 350 1140 356 1141
rect 258 1122 274 1123
rect 346 1127 352 1128
rect 346 1123 347 1127
rect 351 1126 352 1127
rect 360 1126 362 1150
rect 412 1132 414 1158
rect 439 1153 443 1154
rect 1111 1158 1115 1159
rect 1111 1153 1115 1154
rect 440 1146 442 1153
rect 438 1145 444 1146
rect 438 1141 439 1145
rect 443 1141 444 1145
rect 438 1140 444 1141
rect 1112 1134 1114 1153
rect 1110 1133 1116 1134
rect 410 1131 416 1132
rect 410 1127 411 1131
rect 415 1127 416 1131
rect 1110 1129 1111 1133
rect 1115 1129 1116 1133
rect 1110 1128 1116 1129
rect 410 1126 416 1127
rect 351 1124 362 1126
rect 351 1123 352 1124
rect 346 1122 352 1123
rect 260 1121 274 1122
rect 110 1115 116 1116
rect 110 1111 111 1115
rect 115 1111 116 1115
rect 110 1110 116 1111
rect 422 1115 428 1116
rect 422 1111 423 1115
rect 427 1111 428 1115
rect 422 1110 428 1111
rect 1110 1115 1116 1116
rect 1110 1111 1111 1115
rect 1115 1111 1116 1115
rect 1110 1110 1116 1111
rect 112 1095 114 1110
rect 166 1100 172 1101
rect 166 1096 167 1100
rect 171 1096 172 1100
rect 166 1095 172 1096
rect 254 1100 260 1101
rect 254 1096 255 1100
rect 259 1096 260 1100
rect 254 1095 260 1096
rect 342 1100 348 1101
rect 342 1096 343 1100
rect 347 1096 348 1100
rect 342 1095 348 1096
rect 111 1094 115 1095
rect 111 1089 115 1090
rect 167 1094 171 1095
rect 167 1089 171 1090
rect 255 1094 259 1095
rect 255 1089 259 1090
rect 343 1094 347 1095
rect 343 1089 347 1090
rect 399 1094 403 1095
rect 399 1089 403 1090
rect 112 1074 114 1089
rect 398 1088 404 1089
rect 398 1084 399 1088
rect 403 1084 404 1088
rect 398 1083 404 1084
rect 110 1073 116 1074
rect 110 1069 111 1073
rect 115 1069 116 1073
rect 110 1068 116 1069
rect 110 1055 116 1056
rect 110 1051 111 1055
rect 115 1051 116 1055
rect 110 1050 116 1051
rect 112 1031 114 1050
rect 406 1043 412 1044
rect 406 1039 407 1043
rect 411 1039 412 1043
rect 406 1038 412 1039
rect 408 1031 410 1038
rect 424 1036 426 1110
rect 430 1100 436 1101
rect 430 1096 431 1100
rect 435 1096 436 1100
rect 430 1095 436 1096
rect 1112 1095 1114 1110
rect 431 1094 435 1095
rect 431 1089 435 1090
rect 487 1094 491 1095
rect 487 1089 491 1090
rect 575 1094 579 1095
rect 575 1089 579 1090
rect 663 1094 667 1095
rect 663 1089 667 1090
rect 751 1094 755 1095
rect 751 1089 755 1090
rect 839 1094 843 1095
rect 839 1089 843 1090
rect 927 1094 931 1095
rect 1015 1094 1019 1095
rect 927 1089 931 1090
rect 954 1091 960 1092
rect 486 1088 492 1089
rect 486 1084 487 1088
rect 491 1084 492 1088
rect 486 1083 492 1084
rect 574 1088 580 1089
rect 574 1084 575 1088
rect 579 1084 580 1088
rect 574 1083 580 1084
rect 662 1088 668 1089
rect 662 1084 663 1088
rect 667 1084 668 1088
rect 662 1083 668 1084
rect 750 1088 756 1089
rect 750 1084 751 1088
rect 755 1084 756 1088
rect 750 1083 756 1084
rect 838 1088 844 1089
rect 838 1084 839 1088
rect 843 1084 844 1088
rect 838 1083 844 1084
rect 926 1088 932 1089
rect 926 1084 927 1088
rect 931 1084 932 1088
rect 954 1087 955 1091
rect 959 1087 960 1091
rect 1015 1089 1019 1090
rect 1111 1094 1115 1095
rect 1111 1089 1115 1090
rect 954 1086 960 1087
rect 1014 1088 1020 1089
rect 926 1083 932 1084
rect 494 1063 500 1064
rect 494 1059 495 1063
rect 499 1059 500 1063
rect 494 1058 500 1059
rect 582 1063 588 1064
rect 582 1059 583 1063
rect 587 1059 588 1063
rect 582 1058 588 1059
rect 670 1063 676 1064
rect 670 1059 671 1063
rect 675 1059 676 1063
rect 758 1063 764 1064
rect 670 1058 676 1059
rect 742 1059 748 1060
rect 496 1051 498 1058
rect 584 1051 586 1058
rect 672 1051 674 1058
rect 742 1055 743 1059
rect 747 1055 748 1059
rect 758 1059 759 1063
rect 763 1059 764 1063
rect 758 1058 764 1059
rect 934 1063 940 1064
rect 934 1059 935 1063
rect 939 1062 940 1063
rect 939 1060 946 1062
rect 939 1059 940 1060
rect 934 1058 940 1059
rect 742 1054 748 1055
rect 496 1049 506 1051
rect 584 1049 594 1051
rect 672 1049 682 1051
rect 494 1043 500 1044
rect 494 1039 495 1043
rect 499 1039 500 1043
rect 494 1038 500 1039
rect 422 1035 428 1036
rect 422 1031 423 1035
rect 427 1031 428 1035
rect 496 1031 498 1038
rect 504 1036 506 1049
rect 582 1043 588 1044
rect 582 1039 583 1043
rect 587 1039 588 1043
rect 582 1038 588 1039
rect 502 1035 508 1036
rect 502 1031 503 1035
rect 507 1031 508 1035
rect 584 1031 586 1038
rect 592 1036 594 1049
rect 670 1043 676 1044
rect 670 1039 671 1043
rect 675 1039 676 1043
rect 670 1038 676 1039
rect 590 1035 596 1036
rect 590 1031 591 1035
rect 595 1031 596 1035
rect 672 1031 674 1038
rect 680 1036 682 1049
rect 744 1045 746 1054
rect 760 1051 762 1058
rect 760 1049 770 1051
rect 743 1044 747 1045
rect 743 1039 747 1040
rect 758 1043 764 1044
rect 758 1039 759 1043
rect 763 1039 764 1043
rect 758 1038 764 1039
rect 678 1035 684 1036
rect 678 1031 679 1035
rect 683 1031 684 1035
rect 760 1031 762 1038
rect 111 1030 115 1031
rect 111 1025 115 1026
rect 407 1030 411 1031
rect 422 1030 428 1031
rect 495 1030 499 1031
rect 502 1030 508 1031
rect 583 1030 587 1031
rect 590 1030 596 1031
rect 671 1030 675 1031
rect 678 1030 684 1031
rect 759 1030 763 1031
rect 407 1025 411 1026
rect 495 1025 499 1026
rect 502 1027 508 1028
rect 112 1006 114 1025
rect 408 1018 410 1025
rect 414 1023 420 1024
rect 414 1018 415 1023
rect 406 1017 412 1018
rect 406 1013 407 1017
rect 411 1013 412 1017
rect 419 1018 420 1023
rect 496 1018 498 1025
rect 502 1023 503 1027
rect 507 1023 508 1027
rect 583 1025 587 1026
rect 590 1027 596 1028
rect 502 1022 508 1023
rect 415 1015 419 1016
rect 494 1017 500 1018
rect 406 1012 412 1013
rect 494 1013 495 1017
rect 499 1013 500 1017
rect 494 1012 500 1013
rect 110 1005 116 1006
rect 110 1001 111 1005
rect 115 1001 116 1005
rect 110 1000 116 1001
rect 490 999 496 1000
rect 490 995 491 999
rect 495 998 496 999
rect 504 998 506 1022
rect 584 1018 586 1025
rect 590 1023 591 1027
rect 595 1023 596 1027
rect 671 1025 675 1026
rect 768 1028 770 1049
rect 775 1044 779 1045
rect 775 1039 779 1040
rect 846 1043 852 1044
rect 846 1039 847 1043
rect 851 1039 852 1043
rect 776 1036 778 1039
rect 846 1038 852 1039
rect 934 1043 940 1044
rect 934 1039 935 1043
rect 939 1039 940 1043
rect 934 1038 940 1039
rect 774 1035 780 1036
rect 774 1031 775 1035
rect 779 1031 780 1035
rect 848 1031 850 1038
rect 854 1035 860 1036
rect 854 1031 855 1035
rect 859 1031 860 1035
rect 936 1031 938 1038
rect 944 1036 946 1060
rect 942 1035 948 1036
rect 942 1031 943 1035
rect 947 1031 948 1035
rect 774 1030 780 1031
rect 847 1030 851 1031
rect 854 1030 860 1031
rect 935 1030 939 1031
rect 942 1030 948 1031
rect 759 1025 763 1026
rect 766 1027 772 1028
rect 590 1022 596 1023
rect 582 1017 588 1018
rect 582 1013 583 1017
rect 587 1013 588 1017
rect 582 1012 588 1013
rect 495 996 506 998
rect 578 999 584 1000
rect 495 995 496 996
rect 490 994 496 995
rect 578 995 579 999
rect 583 998 584 999
rect 592 998 594 1022
rect 651 1020 655 1021
rect 672 1018 674 1025
rect 678 1023 684 1024
rect 678 1018 679 1023
rect 651 1015 655 1016
rect 670 1017 676 1018
rect 652 1000 654 1015
rect 670 1013 671 1017
rect 675 1013 676 1017
rect 683 1018 684 1023
rect 739 1020 743 1021
rect 679 1015 683 1016
rect 760 1018 762 1025
rect 766 1023 767 1027
rect 771 1023 772 1027
rect 847 1025 851 1026
rect 766 1022 772 1023
rect 848 1018 850 1025
rect 739 1015 743 1016
rect 758 1017 764 1018
rect 670 1012 676 1013
rect 740 1000 742 1015
rect 758 1013 759 1017
rect 763 1013 764 1017
rect 758 1012 764 1013
rect 846 1017 852 1018
rect 846 1013 847 1017
rect 851 1013 852 1017
rect 846 1012 852 1013
rect 583 996 594 998
rect 650 999 656 1000
rect 583 995 584 996
rect 578 994 584 995
rect 650 995 651 999
rect 655 995 656 999
rect 650 994 656 995
rect 738 999 744 1000
rect 738 995 739 999
rect 743 995 744 999
rect 738 994 744 995
rect 846 999 852 1000
rect 846 995 847 999
rect 851 998 852 999
rect 856 998 858 1030
rect 956 1026 958 1086
rect 1014 1084 1015 1088
rect 1019 1084 1020 1088
rect 1014 1083 1020 1084
rect 1112 1074 1114 1089
rect 1110 1073 1116 1074
rect 1110 1069 1111 1073
rect 1115 1069 1116 1073
rect 1110 1068 1116 1069
rect 1022 1063 1028 1064
rect 1022 1059 1023 1063
rect 1027 1059 1028 1063
rect 1022 1058 1028 1059
rect 1024 1051 1026 1058
rect 1110 1055 1116 1056
rect 1110 1051 1111 1055
rect 1115 1051 1116 1055
rect 1024 1049 1034 1051
rect 1110 1050 1116 1051
rect 1022 1043 1028 1044
rect 1022 1039 1023 1043
rect 1027 1039 1028 1043
rect 1022 1038 1028 1039
rect 1024 1031 1026 1038
rect 1032 1036 1034 1049
rect 1030 1035 1036 1036
rect 1030 1031 1031 1035
rect 1035 1031 1036 1035
rect 1112 1031 1114 1050
rect 1023 1030 1027 1031
rect 1030 1030 1036 1031
rect 1111 1030 1115 1031
rect 862 1025 868 1026
rect 935 1025 939 1026
rect 954 1025 960 1026
rect 1023 1025 1027 1026
rect 1030 1027 1036 1028
rect 862 1021 863 1025
rect 867 1021 868 1025
rect 862 1020 868 1021
rect 851 996 858 998
rect 851 995 852 996
rect 846 994 852 995
rect 110 987 116 988
rect 110 983 111 987
rect 115 983 116 987
rect 110 982 116 983
rect 670 987 676 988
rect 670 983 671 987
rect 675 983 676 987
rect 670 982 676 983
rect 112 951 114 982
rect 398 972 404 973
rect 398 968 399 972
rect 403 968 404 972
rect 398 967 404 968
rect 486 972 492 973
rect 486 968 487 972
rect 491 968 492 972
rect 486 967 492 968
rect 574 972 580 973
rect 574 968 575 972
rect 579 968 580 972
rect 574 967 580 968
rect 662 972 668 973
rect 662 968 663 972
rect 667 968 668 972
rect 662 967 668 968
rect 400 951 402 967
rect 488 951 490 967
rect 576 951 578 967
rect 664 951 666 967
rect 111 950 115 951
rect 111 945 115 946
rect 151 950 155 951
rect 151 945 155 946
rect 271 950 275 951
rect 271 945 275 946
rect 399 950 403 951
rect 399 945 403 946
rect 407 950 411 951
rect 407 945 411 946
rect 487 950 491 951
rect 487 945 491 946
rect 551 950 555 951
rect 551 945 555 946
rect 575 950 579 951
rect 575 945 579 946
rect 663 950 667 951
rect 663 945 667 946
rect 112 930 114 945
rect 150 944 156 945
rect 150 940 151 944
rect 155 940 156 944
rect 150 939 156 940
rect 270 944 276 945
rect 270 940 271 944
rect 275 940 276 944
rect 270 939 276 940
rect 406 944 412 945
rect 406 940 407 944
rect 411 940 412 944
rect 406 939 412 940
rect 550 944 556 945
rect 550 940 551 944
rect 555 940 556 944
rect 550 939 556 940
rect 110 929 116 930
rect 110 925 111 929
rect 115 925 116 929
rect 110 924 116 925
rect 370 915 376 916
rect 110 911 116 912
rect 110 907 111 911
rect 115 907 116 911
rect 370 911 371 915
rect 375 911 376 915
rect 370 910 376 911
rect 502 915 508 916
rect 502 911 503 915
rect 507 911 508 915
rect 502 910 508 911
rect 654 915 660 916
rect 654 911 655 915
rect 659 911 660 915
rect 654 910 660 911
rect 110 906 116 907
rect 112 879 114 906
rect 158 899 164 900
rect 158 895 159 899
rect 163 895 164 899
rect 158 894 164 895
rect 278 899 284 900
rect 278 895 279 899
rect 283 895 284 899
rect 278 894 284 895
rect 160 879 162 894
rect 218 883 224 884
rect 218 879 219 883
rect 223 879 224 883
rect 280 879 282 894
rect 372 884 374 910
rect 414 899 420 900
rect 414 895 415 899
rect 419 895 420 899
rect 414 894 420 895
rect 370 883 376 884
rect 370 879 371 883
rect 375 879 376 883
rect 416 879 418 894
rect 504 884 506 910
rect 558 899 564 900
rect 558 895 559 899
rect 563 895 564 899
rect 558 894 564 895
rect 502 883 508 884
rect 502 879 503 883
rect 507 879 508 883
rect 560 879 562 894
rect 656 884 658 910
rect 672 884 674 982
rect 750 972 756 973
rect 750 968 751 972
rect 755 968 756 972
rect 750 967 756 968
rect 838 972 844 973
rect 838 968 839 972
rect 843 968 844 972
rect 838 967 844 968
rect 752 951 754 967
rect 840 951 842 967
rect 711 950 715 951
rect 711 945 715 946
rect 751 950 755 951
rect 751 945 755 946
rect 839 950 843 951
rect 839 945 843 946
rect 710 944 716 945
rect 710 940 711 944
rect 715 940 716 944
rect 710 939 716 940
rect 864 932 866 1020
rect 936 1018 938 1025
rect 954 1021 955 1025
rect 959 1021 960 1025
rect 954 1020 960 1021
rect 1024 1018 1026 1025
rect 1030 1023 1031 1027
rect 1035 1023 1036 1027
rect 1111 1025 1115 1026
rect 1030 1022 1036 1023
rect 934 1017 940 1018
rect 934 1013 935 1017
rect 939 1013 940 1017
rect 934 1012 940 1013
rect 1022 1017 1028 1018
rect 1022 1013 1023 1017
rect 1027 1013 1028 1017
rect 1022 1012 1028 1013
rect 1018 999 1024 1000
rect 1018 995 1019 999
rect 1023 998 1024 999
rect 1032 998 1034 1022
rect 1112 1006 1114 1025
rect 1110 1005 1116 1006
rect 1110 1001 1111 1005
rect 1115 1001 1116 1005
rect 1110 1000 1116 1001
rect 1023 996 1034 998
rect 1023 995 1024 996
rect 1018 994 1024 995
rect 1022 987 1028 988
rect 1022 983 1023 987
rect 1027 983 1028 987
rect 1022 982 1028 983
rect 1110 987 1116 988
rect 1110 983 1111 987
rect 1115 983 1116 987
rect 1110 982 1116 983
rect 926 972 932 973
rect 926 968 927 972
rect 931 968 932 972
rect 926 967 932 968
rect 1014 972 1020 973
rect 1014 968 1015 972
rect 1019 968 1020 972
rect 1014 967 1020 968
rect 928 951 930 967
rect 1016 951 1018 967
rect 871 950 875 951
rect 871 945 875 946
rect 927 950 931 951
rect 927 945 931 946
rect 1015 950 1019 951
rect 1015 945 1019 946
rect 870 944 876 945
rect 870 940 871 944
rect 875 940 876 944
rect 870 939 876 940
rect 1014 944 1020 945
rect 1014 940 1015 944
rect 1019 940 1020 944
rect 1014 939 1020 940
rect 862 931 868 932
rect 862 927 863 931
rect 867 927 868 931
rect 862 926 868 927
rect 1024 907 1026 982
rect 1112 951 1114 982
rect 1111 950 1115 951
rect 1111 945 1115 946
rect 1112 930 1114 945
rect 1110 929 1116 930
rect 1110 925 1111 929
rect 1115 925 1116 929
rect 1110 924 1116 925
rect 1082 915 1088 916
rect 1082 911 1083 915
rect 1087 911 1088 915
rect 1082 910 1088 911
rect 1110 911 1116 912
rect 1024 905 1034 907
rect 718 899 724 900
rect 718 895 719 899
rect 723 895 724 899
rect 718 894 724 895
rect 878 899 884 900
rect 878 895 879 899
rect 883 895 884 899
rect 878 894 884 895
rect 1022 899 1028 900
rect 1022 895 1023 899
rect 1027 895 1028 899
rect 1022 894 1028 895
rect 654 883 660 884
rect 654 879 655 883
rect 659 879 660 883
rect 111 878 115 879
rect 111 873 115 874
rect 143 878 147 879
rect 143 873 147 874
rect 159 878 163 879
rect 218 878 224 879
rect 271 878 275 879
rect 159 873 163 874
rect 112 854 114 873
rect 144 866 146 873
rect 142 865 148 866
rect 142 861 143 865
rect 147 861 148 865
rect 142 860 148 861
rect 110 853 116 854
rect 110 849 111 853
rect 115 849 116 853
rect 220 852 222 878
rect 271 873 275 874
rect 279 878 283 879
rect 370 878 376 879
rect 415 878 419 879
rect 279 873 283 874
rect 415 873 419 874
rect 439 878 443 879
rect 502 878 508 879
rect 559 878 563 879
rect 439 873 443 874
rect 446 875 452 876
rect 272 866 274 873
rect 440 866 442 873
rect 446 871 447 875
rect 451 871 452 875
rect 559 873 563 874
rect 631 878 635 879
rect 654 878 660 879
rect 670 883 676 884
rect 670 879 671 883
rect 675 879 676 883
rect 720 879 722 894
rect 754 883 760 884
rect 754 879 755 883
rect 759 879 760 883
rect 880 879 882 894
rect 930 883 936 884
rect 930 879 931 883
rect 935 879 936 883
rect 1024 879 1026 894
rect 1032 892 1034 905
rect 1030 891 1036 892
rect 1030 887 1031 891
rect 1035 887 1036 891
rect 1030 886 1036 887
rect 1084 884 1086 910
rect 1110 907 1111 911
rect 1115 907 1116 911
rect 1110 906 1116 907
rect 1082 883 1088 884
rect 1082 879 1083 883
rect 1087 879 1088 883
rect 1112 879 1114 906
rect 670 878 676 879
rect 719 878 723 879
rect 754 878 760 879
rect 839 878 843 879
rect 631 873 635 874
rect 638 875 644 876
rect 446 870 452 871
rect 270 865 276 866
rect 270 861 271 865
rect 275 861 276 865
rect 270 860 276 861
rect 438 865 444 866
rect 438 861 439 865
rect 443 861 444 865
rect 438 860 444 861
rect 110 848 116 849
rect 218 851 224 852
rect 218 847 219 851
rect 223 847 224 851
rect 218 846 224 847
rect 434 847 440 848
rect 434 843 435 847
rect 439 846 440 847
rect 448 846 450 870
rect 632 866 634 873
rect 638 871 639 875
rect 643 871 644 875
rect 719 873 723 874
rect 638 870 644 871
rect 630 865 636 866
rect 630 861 631 865
rect 635 861 636 865
rect 630 860 636 861
rect 439 844 450 846
rect 626 847 632 848
rect 439 843 440 844
rect 434 842 440 843
rect 626 843 627 847
rect 631 846 632 847
rect 640 846 642 870
rect 756 852 758 878
rect 839 873 843 874
rect 879 878 883 879
rect 930 878 936 879
rect 1023 878 1027 879
rect 1082 878 1088 879
rect 1111 878 1115 879
rect 879 873 883 874
rect 840 866 842 873
rect 838 865 844 866
rect 838 861 839 865
rect 843 861 844 865
rect 838 860 844 861
rect 754 851 760 852
rect 754 847 755 851
rect 759 847 760 851
rect 754 846 760 847
rect 631 844 642 846
rect 631 843 632 844
rect 626 842 632 843
rect 110 835 116 836
rect 110 831 111 835
rect 115 831 116 835
rect 110 830 116 831
rect 738 835 744 836
rect 738 831 739 835
rect 743 831 744 835
rect 738 830 744 831
rect 112 803 114 830
rect 134 820 140 821
rect 134 816 135 820
rect 139 816 140 820
rect 134 815 140 816
rect 262 820 268 821
rect 262 816 263 820
rect 267 816 268 820
rect 262 815 268 816
rect 430 820 436 821
rect 430 816 431 820
rect 435 816 436 820
rect 430 815 436 816
rect 622 820 628 821
rect 622 816 623 820
rect 627 816 628 820
rect 622 815 628 816
rect 136 803 138 815
rect 264 803 266 815
rect 432 803 434 815
rect 624 803 626 815
rect 111 802 115 803
rect 111 797 115 798
rect 135 802 139 803
rect 135 797 139 798
rect 239 802 243 803
rect 239 797 243 798
rect 263 802 267 803
rect 263 797 267 798
rect 375 802 379 803
rect 375 797 379 798
rect 431 802 435 803
rect 431 797 435 798
rect 527 802 531 803
rect 527 797 531 798
rect 623 802 627 803
rect 623 797 627 798
rect 695 802 699 803
rect 695 797 699 798
rect 112 782 114 797
rect 134 796 140 797
rect 134 792 135 796
rect 139 792 140 796
rect 134 791 140 792
rect 238 796 244 797
rect 238 792 239 796
rect 243 792 244 796
rect 238 791 244 792
rect 374 796 380 797
rect 374 792 375 796
rect 379 792 380 796
rect 374 791 380 792
rect 526 796 532 797
rect 526 792 527 796
rect 531 792 532 796
rect 526 791 532 792
rect 694 796 700 797
rect 694 792 695 796
rect 699 792 700 796
rect 694 791 700 792
rect 110 781 116 782
rect 110 777 111 781
rect 115 777 116 781
rect 110 776 116 777
rect 210 767 216 768
rect 163 764 167 765
rect 110 763 116 764
rect 110 759 111 763
rect 115 759 116 763
rect 210 763 211 767
rect 215 763 216 767
rect 210 762 216 763
rect 482 767 488 768
rect 482 763 483 767
rect 487 763 488 767
rect 482 762 488 763
rect 674 767 680 768
rect 674 763 675 767
rect 679 763 680 767
rect 674 762 680 763
rect 682 767 688 768
rect 682 763 683 767
rect 687 763 688 767
rect 740 765 742 830
rect 830 820 836 821
rect 830 816 831 820
rect 835 816 836 820
rect 830 815 836 816
rect 832 803 834 815
rect 831 802 835 803
rect 831 797 835 798
rect 863 802 867 803
rect 863 797 867 798
rect 862 796 868 797
rect 862 792 863 796
rect 867 792 868 796
rect 862 791 868 792
rect 932 784 934 878
rect 1023 873 1027 874
rect 1111 873 1115 874
rect 1024 866 1026 873
rect 1022 865 1028 866
rect 1022 861 1023 865
rect 1027 861 1028 865
rect 1022 860 1028 861
rect 1112 854 1114 873
rect 1110 853 1116 854
rect 1110 849 1111 853
rect 1115 849 1116 853
rect 1110 848 1116 849
rect 1022 835 1028 836
rect 1022 831 1023 835
rect 1027 831 1028 835
rect 1022 830 1028 831
rect 1110 835 1116 836
rect 1110 831 1111 835
rect 1115 831 1116 835
rect 1110 830 1116 831
rect 1014 820 1020 821
rect 1014 816 1015 820
rect 1019 816 1020 820
rect 1014 815 1020 816
rect 1016 803 1018 815
rect 1015 802 1019 803
rect 1015 797 1019 798
rect 1014 796 1020 797
rect 1014 792 1015 796
rect 1019 792 1020 796
rect 1014 791 1020 792
rect 1024 787 1026 830
rect 1112 803 1114 830
rect 1111 802 1115 803
rect 1111 797 1115 798
rect 1024 785 1042 787
rect 930 783 936 784
rect 930 779 931 783
rect 935 779 936 783
rect 930 778 936 779
rect 1022 771 1028 772
rect 1022 767 1023 771
rect 1027 767 1028 771
rect 1022 766 1028 767
rect 682 762 688 763
rect 739 764 743 765
rect 163 759 167 760
rect 110 758 116 759
rect 112 735 114 758
rect 142 751 148 752
rect 142 747 143 751
rect 147 747 148 751
rect 142 746 148 747
rect 144 735 146 746
rect 164 744 166 759
rect 162 743 168 744
rect 162 739 163 743
rect 167 739 168 743
rect 162 738 168 739
rect 212 736 214 762
rect 246 751 252 752
rect 246 747 247 751
rect 251 747 252 751
rect 382 751 388 752
rect 246 746 252 747
rect 291 748 295 749
rect 210 735 216 736
rect 248 735 250 746
rect 382 747 383 751
rect 387 747 388 751
rect 382 746 388 747
rect 291 743 295 744
rect 111 734 115 735
rect 111 729 115 730
rect 143 734 147 735
rect 210 731 211 735
rect 215 731 216 735
rect 210 730 216 731
rect 247 734 251 735
rect 143 729 147 730
rect 247 729 251 730
rect 271 734 275 735
rect 292 732 294 743
rect 384 735 386 746
rect 430 739 436 740
rect 430 735 431 739
rect 435 735 436 739
rect 484 736 486 762
rect 534 751 540 752
rect 534 747 535 751
rect 539 747 540 751
rect 534 746 540 747
rect 482 735 488 736
rect 536 735 538 746
rect 582 739 588 740
rect 582 735 583 739
rect 587 735 588 739
rect 676 736 678 762
rect 684 749 686 762
rect 1024 763 1026 766
rect 1024 761 1034 763
rect 739 759 743 760
rect 702 751 708 752
rect 683 748 687 749
rect 702 747 703 751
rect 707 747 708 751
rect 702 746 708 747
rect 870 751 876 752
rect 870 747 871 751
rect 875 747 876 751
rect 870 746 876 747
rect 1022 751 1028 752
rect 1022 747 1023 751
rect 1027 747 1028 751
rect 1022 746 1028 747
rect 683 743 687 744
rect 674 735 680 736
rect 704 735 706 746
rect 750 739 756 740
rect 750 735 751 739
rect 755 735 756 739
rect 872 735 874 746
rect 886 743 892 744
rect 886 739 887 743
rect 891 739 892 743
rect 886 738 892 739
rect 383 734 387 735
rect 430 734 436 735
rect 447 734 451 735
rect 271 729 275 730
rect 290 731 296 732
rect 112 710 114 729
rect 272 722 274 729
rect 290 727 291 731
rect 295 727 296 731
rect 383 729 387 730
rect 290 726 296 727
rect 270 721 276 722
rect 270 717 271 721
rect 275 717 276 721
rect 270 716 276 717
rect 110 709 116 710
rect 110 705 111 709
rect 115 705 116 709
rect 432 708 434 734
rect 482 731 483 735
rect 487 731 488 735
rect 482 730 488 731
rect 535 734 539 735
rect 582 734 588 735
rect 639 734 643 735
rect 447 729 451 730
rect 535 729 539 730
rect 448 722 450 729
rect 446 721 452 722
rect 446 717 447 721
rect 451 717 452 721
rect 446 716 452 717
rect 584 708 586 734
rect 674 731 675 735
rect 679 731 680 735
rect 674 730 680 731
rect 703 734 707 735
rect 750 734 756 735
rect 831 734 835 735
rect 639 729 643 730
rect 703 729 707 730
rect 640 722 642 729
rect 638 721 644 722
rect 638 717 639 721
rect 643 717 644 721
rect 638 716 644 717
rect 752 708 754 734
rect 831 729 835 730
rect 871 734 875 735
rect 871 729 875 730
rect 832 722 834 729
rect 830 721 836 722
rect 830 717 831 721
rect 835 717 836 721
rect 830 716 836 717
rect 110 704 116 705
rect 430 707 436 708
rect 430 703 431 707
rect 435 703 436 707
rect 430 702 436 703
rect 582 707 588 708
rect 582 703 583 707
rect 587 703 588 707
rect 582 702 588 703
rect 750 707 756 708
rect 750 703 751 707
rect 755 703 756 707
rect 750 702 756 703
rect 110 691 116 692
rect 110 687 111 691
rect 115 687 116 691
rect 110 686 116 687
rect 738 691 744 692
rect 738 687 739 691
rect 743 687 744 691
rect 738 686 744 687
rect 112 671 114 686
rect 262 676 268 677
rect 262 672 263 676
rect 267 672 268 676
rect 262 671 268 672
rect 438 676 444 677
rect 438 672 439 676
rect 443 672 444 676
rect 438 671 444 672
rect 630 676 636 677
rect 630 672 631 676
rect 635 672 636 676
rect 630 671 636 672
rect 111 670 115 671
rect 111 665 115 666
rect 263 670 267 671
rect 263 665 267 666
rect 367 670 371 671
rect 367 665 371 666
rect 439 670 443 671
rect 439 665 443 666
rect 463 670 467 671
rect 463 665 467 666
rect 559 670 563 671
rect 559 665 563 666
rect 631 670 635 671
rect 631 665 635 666
rect 663 670 667 671
rect 663 665 667 666
rect 112 650 114 665
rect 366 664 372 665
rect 366 660 367 664
rect 371 660 372 664
rect 366 659 372 660
rect 462 664 468 665
rect 462 660 463 664
rect 467 660 468 664
rect 462 659 468 660
rect 558 664 564 665
rect 558 660 559 664
rect 563 660 564 664
rect 558 659 564 660
rect 662 664 668 665
rect 662 660 663 664
rect 667 660 668 664
rect 662 659 668 660
rect 110 649 116 650
rect 110 645 111 649
rect 115 645 116 649
rect 110 644 116 645
rect 438 635 444 636
rect 110 631 116 632
rect 110 627 111 631
rect 115 627 116 631
rect 438 631 439 635
rect 443 631 444 635
rect 438 630 444 631
rect 534 635 540 636
rect 534 631 535 635
rect 539 631 540 635
rect 534 630 540 631
rect 638 635 644 636
rect 638 631 639 635
rect 643 631 644 635
rect 638 630 644 631
rect 110 626 116 627
rect 112 595 114 626
rect 395 620 399 621
rect 374 619 380 620
rect 374 615 375 619
rect 379 615 380 619
rect 395 615 399 616
rect 374 614 380 615
rect 376 595 378 614
rect 396 612 398 615
rect 394 611 400 612
rect 394 607 395 611
rect 399 607 400 611
rect 394 606 400 607
rect 440 604 442 630
rect 470 619 476 620
rect 470 615 471 619
rect 475 615 476 619
rect 470 614 476 615
rect 438 603 444 604
rect 438 599 439 603
rect 443 599 444 603
rect 438 598 444 599
rect 472 595 474 614
rect 515 604 519 605
rect 536 604 538 630
rect 566 619 572 620
rect 566 615 567 619
rect 571 615 572 619
rect 566 614 572 615
rect 515 599 519 600
rect 534 603 540 604
rect 534 599 535 603
rect 539 599 540 603
rect 111 594 115 595
rect 111 589 115 590
rect 375 594 379 595
rect 375 589 379 590
rect 471 594 475 595
rect 471 589 475 590
rect 495 594 499 595
rect 516 592 518 599
rect 534 598 540 599
rect 568 595 570 614
rect 640 604 642 630
rect 740 621 742 686
rect 822 676 828 677
rect 822 672 823 676
rect 827 672 828 676
rect 822 671 828 672
rect 775 670 779 671
rect 775 665 779 666
rect 823 670 827 671
rect 823 665 827 666
rect 774 664 780 665
rect 774 660 775 664
rect 779 660 780 664
rect 774 659 780 660
rect 888 652 890 738
rect 1024 735 1026 746
rect 1023 734 1027 735
rect 1032 732 1034 761
rect 1040 744 1042 785
rect 1112 782 1114 797
rect 1110 781 1116 782
rect 1110 777 1111 781
rect 1115 777 1116 781
rect 1110 776 1116 777
rect 1110 763 1116 764
rect 1110 759 1111 763
rect 1115 759 1116 763
rect 1110 758 1116 759
rect 1038 743 1044 744
rect 1038 739 1039 743
rect 1043 739 1044 743
rect 1038 738 1044 739
rect 1112 735 1114 758
rect 1111 734 1115 735
rect 1023 729 1027 730
rect 1030 731 1036 732
rect 1024 722 1026 729
rect 1030 727 1031 731
rect 1035 727 1036 731
rect 1111 729 1115 730
rect 1030 726 1036 727
rect 1022 721 1028 722
rect 1022 717 1023 721
rect 1027 717 1028 721
rect 1022 716 1028 717
rect 1112 710 1114 729
rect 1110 709 1116 710
rect 1110 705 1111 709
rect 1115 705 1116 709
rect 1110 704 1116 705
rect 1022 691 1028 692
rect 1022 687 1023 691
rect 1027 687 1028 691
rect 1022 686 1028 687
rect 1110 691 1116 692
rect 1110 687 1111 691
rect 1115 687 1116 691
rect 1110 686 1116 687
rect 1014 676 1020 677
rect 1014 672 1015 676
rect 1019 672 1020 676
rect 1014 671 1020 672
rect 895 670 899 671
rect 895 665 899 666
rect 1015 670 1019 671
rect 1015 665 1019 666
rect 894 664 900 665
rect 894 660 895 664
rect 899 660 900 664
rect 894 659 900 660
rect 886 651 892 652
rect 886 647 887 651
rect 891 647 892 651
rect 886 646 892 647
rect 746 635 752 636
rect 746 631 747 635
rect 751 631 752 635
rect 746 630 752 631
rect 754 635 760 636
rect 754 631 755 635
rect 759 631 760 635
rect 754 630 760 631
rect 739 620 743 621
rect 670 619 676 620
rect 670 615 671 619
rect 675 615 676 619
rect 739 615 743 616
rect 670 614 676 615
rect 638 603 644 604
rect 638 599 639 603
rect 643 599 644 603
rect 638 598 644 599
rect 672 595 674 614
rect 748 604 750 630
rect 756 605 758 630
rect 782 619 788 620
rect 782 615 783 619
rect 787 615 788 619
rect 782 614 788 615
rect 902 619 908 620
rect 902 615 903 619
rect 907 615 908 619
rect 902 614 908 615
rect 755 604 759 605
rect 746 603 752 604
rect 746 599 747 603
rect 751 599 752 603
rect 755 599 759 600
rect 746 598 752 599
rect 784 595 786 614
rect 904 595 906 614
rect 922 611 928 612
rect 922 607 923 611
rect 927 607 928 611
rect 922 606 928 607
rect 567 594 571 595
rect 495 589 499 590
rect 514 591 520 592
rect 112 570 114 589
rect 496 582 498 589
rect 514 587 515 591
rect 519 587 520 591
rect 567 589 571 590
rect 583 594 587 595
rect 671 594 675 595
rect 583 589 587 590
rect 590 591 596 592
rect 514 586 520 587
rect 584 582 586 589
rect 590 587 591 591
rect 595 587 596 591
rect 759 594 763 595
rect 671 589 675 590
rect 678 591 684 592
rect 590 586 596 587
rect 494 581 500 582
rect 494 577 495 581
rect 499 577 500 581
rect 494 576 500 577
rect 582 581 588 582
rect 582 577 583 581
rect 587 577 588 581
rect 582 576 588 577
rect 592 571 594 586
rect 672 582 674 589
rect 678 587 679 591
rect 683 587 684 591
rect 783 594 787 595
rect 759 589 763 590
rect 766 591 772 592
rect 678 586 684 587
rect 670 581 676 582
rect 670 577 671 581
rect 675 577 676 581
rect 670 576 676 577
rect 680 571 682 586
rect 760 582 762 589
rect 766 587 767 591
rect 771 587 772 591
rect 783 589 787 590
rect 847 594 851 595
rect 903 594 907 595
rect 847 589 851 590
rect 854 591 860 592
rect 766 586 772 587
rect 758 581 764 582
rect 758 577 759 581
rect 763 577 764 581
rect 758 576 764 577
rect 768 571 770 586
rect 848 582 850 589
rect 854 587 855 591
rect 859 587 860 591
rect 903 589 907 590
rect 854 586 860 587
rect 846 581 852 582
rect 846 577 847 581
rect 851 577 852 581
rect 846 576 852 577
rect 856 571 858 586
rect 110 569 116 570
rect 110 565 111 569
rect 115 565 116 569
rect 110 564 116 565
rect 584 569 594 571
rect 672 569 682 571
rect 760 569 770 571
rect 848 569 858 571
rect 584 564 586 569
rect 672 564 674 569
rect 760 564 762 569
rect 848 564 850 569
rect 924 564 926 606
rect 1024 603 1026 686
rect 1112 671 1114 686
rect 1111 670 1115 671
rect 1111 665 1115 666
rect 1112 650 1114 665
rect 1110 649 1116 650
rect 1110 645 1111 649
rect 1115 645 1116 649
rect 1110 644 1116 645
rect 1110 631 1116 632
rect 1110 627 1111 631
rect 1115 627 1116 631
rect 1110 626 1116 627
rect 1024 601 1034 603
rect 935 594 939 595
rect 1023 594 1027 595
rect 935 589 939 590
rect 950 591 956 592
rect 936 582 938 589
rect 950 587 951 591
rect 955 587 956 591
rect 1032 592 1034 601
rect 1112 595 1114 626
rect 1111 594 1115 595
rect 1023 589 1027 590
rect 1030 591 1036 592
rect 950 586 956 587
rect 934 581 940 582
rect 934 577 935 581
rect 939 577 940 581
rect 934 576 940 577
rect 582 563 588 564
rect 582 559 583 563
rect 587 559 588 563
rect 582 558 588 559
rect 670 563 676 564
rect 670 559 671 563
rect 675 559 676 563
rect 670 558 676 559
rect 758 563 764 564
rect 758 559 759 563
rect 763 559 764 563
rect 758 558 764 559
rect 846 563 852 564
rect 846 559 847 563
rect 851 559 852 563
rect 846 558 852 559
rect 922 563 928 564
rect 922 559 923 563
rect 927 559 928 563
rect 922 558 928 559
rect 110 551 116 552
rect 110 547 111 551
rect 115 547 116 551
rect 110 546 116 547
rect 906 547 912 548
rect 112 519 114 546
rect 906 543 907 547
rect 911 543 912 547
rect 906 542 912 543
rect 486 536 492 537
rect 486 532 487 536
rect 491 532 492 536
rect 486 531 492 532
rect 574 536 580 537
rect 574 532 575 536
rect 579 532 580 536
rect 574 531 580 532
rect 662 536 668 537
rect 662 532 663 536
rect 667 532 668 536
rect 662 531 668 532
rect 750 536 756 537
rect 750 532 751 536
rect 755 532 756 536
rect 750 531 756 532
rect 838 536 844 537
rect 838 532 839 536
rect 843 532 844 536
rect 838 531 844 532
rect 488 519 490 531
rect 576 519 578 531
rect 664 519 666 531
rect 752 519 754 531
rect 840 519 842 531
rect 111 518 115 519
rect 111 513 115 514
rect 447 518 451 519
rect 447 513 451 514
rect 487 518 491 519
rect 487 513 491 514
rect 543 518 547 519
rect 543 513 547 514
rect 575 518 579 519
rect 575 513 579 514
rect 647 518 651 519
rect 647 513 651 514
rect 663 518 667 519
rect 663 513 667 514
rect 751 518 755 519
rect 751 513 755 514
rect 759 518 763 519
rect 759 513 763 514
rect 839 518 843 519
rect 839 513 843 514
rect 871 518 875 519
rect 871 513 875 514
rect 112 498 114 513
rect 446 512 452 513
rect 446 508 447 512
rect 451 508 452 512
rect 446 507 452 508
rect 542 512 548 513
rect 542 508 543 512
rect 547 508 548 512
rect 542 507 548 508
rect 646 512 652 513
rect 646 508 647 512
rect 651 508 652 512
rect 646 507 652 508
rect 758 512 764 513
rect 758 508 759 512
rect 763 508 764 512
rect 758 507 764 508
rect 870 512 876 513
rect 870 508 871 512
rect 875 508 876 512
rect 870 507 876 508
rect 908 499 910 542
rect 926 536 932 537
rect 926 532 927 536
rect 931 532 932 536
rect 926 531 932 532
rect 928 519 930 531
rect 927 518 931 519
rect 927 513 931 514
rect 110 497 116 498
rect 110 493 111 497
rect 115 493 116 497
rect 110 492 116 493
rect 900 497 910 499
rect 550 487 556 488
rect 550 483 551 487
rect 555 483 556 487
rect 550 482 556 483
rect 618 483 624 484
rect 110 479 116 480
rect 110 475 111 479
rect 115 475 116 479
rect 110 474 116 475
rect 552 475 554 482
rect 618 479 619 483
rect 623 479 624 483
rect 618 478 624 479
rect 714 483 720 484
rect 714 479 715 483
rect 719 479 720 483
rect 714 478 720 479
rect 722 483 728 484
rect 722 479 723 483
rect 727 479 728 483
rect 722 478 728 479
rect 112 451 114 474
rect 552 473 562 475
rect 454 467 460 468
rect 454 463 455 467
rect 459 463 460 467
rect 454 462 460 463
rect 550 467 556 468
rect 550 463 551 467
rect 555 463 556 467
rect 550 462 556 463
rect 456 451 458 462
rect 475 460 479 461
rect 474 455 475 460
rect 479 455 480 460
rect 474 454 480 455
rect 490 451 496 452
rect 552 451 554 462
rect 560 460 562 473
rect 558 459 564 460
rect 558 455 559 459
rect 563 455 564 459
rect 558 454 564 455
rect 620 452 622 478
rect 654 467 660 468
rect 654 463 655 467
rect 659 463 660 467
rect 654 462 660 463
rect 618 451 624 452
rect 656 451 658 462
rect 716 456 718 478
rect 724 461 726 478
rect 766 467 772 468
rect 766 463 767 467
rect 771 463 772 467
rect 766 462 772 463
rect 878 467 884 468
rect 878 463 879 467
rect 883 463 884 467
rect 878 462 884 463
rect 723 460 727 461
rect 714 455 720 456
rect 723 455 727 456
rect 714 451 715 455
rect 719 451 720 455
rect 768 451 770 462
rect 880 451 882 462
rect 900 460 902 497
rect 898 459 904 460
rect 898 455 899 459
rect 903 455 904 459
rect 898 454 904 455
rect 111 450 115 451
rect 111 445 115 446
rect 279 450 283 451
rect 279 445 283 446
rect 407 450 411 451
rect 455 450 459 451
rect 407 445 411 446
rect 414 447 420 448
rect 112 426 114 445
rect 280 438 282 445
rect 408 438 410 445
rect 414 443 415 447
rect 419 443 420 447
rect 490 447 491 451
rect 495 447 496 451
rect 490 446 496 447
rect 543 450 547 451
rect 455 445 459 446
rect 414 442 420 443
rect 278 437 284 438
rect 278 433 279 437
rect 283 433 284 437
rect 278 432 284 433
rect 406 437 412 438
rect 406 433 407 437
rect 411 433 412 437
rect 406 432 412 433
rect 416 427 418 442
rect 110 425 116 426
rect 110 421 111 425
rect 115 421 116 425
rect 110 420 116 421
rect 408 425 418 427
rect 408 420 410 425
rect 492 420 494 446
rect 543 445 547 446
rect 551 450 555 451
rect 551 445 555 446
rect 562 447 568 448
rect 544 438 546 445
rect 562 443 563 447
rect 567 443 568 447
rect 618 447 619 451
rect 623 447 624 451
rect 618 446 624 447
rect 655 450 659 451
rect 655 445 659 446
rect 687 450 691 451
rect 714 450 720 451
rect 767 450 771 451
rect 687 445 691 446
rect 767 445 771 446
rect 839 450 843 451
rect 879 450 883 451
rect 839 445 843 446
rect 858 447 864 448
rect 562 442 568 443
rect 542 437 548 438
rect 564 437 566 442
rect 688 438 690 445
rect 840 438 842 445
rect 858 443 859 447
rect 863 443 864 447
rect 879 445 883 446
rect 858 442 864 443
rect 686 437 692 438
rect 542 433 543 437
rect 547 433 548 437
rect 542 432 548 433
rect 563 436 567 437
rect 563 431 567 432
rect 611 436 615 437
rect 686 433 687 437
rect 691 433 692 437
rect 686 432 692 433
rect 838 437 844 438
rect 838 433 839 437
rect 843 433 844 437
rect 838 432 844 433
rect 611 431 615 432
rect 612 420 614 431
rect 406 419 412 420
rect 406 415 407 419
rect 411 415 412 419
rect 406 414 412 415
rect 490 419 496 420
rect 490 415 491 419
rect 495 415 496 419
rect 490 414 496 415
rect 610 419 616 420
rect 610 415 611 419
rect 615 415 616 419
rect 610 414 616 415
rect 110 407 116 408
rect 110 403 111 407
rect 115 403 116 407
rect 110 402 116 403
rect 502 407 508 408
rect 502 403 503 407
rect 507 403 508 407
rect 502 402 508 403
rect 112 387 114 402
rect 270 392 276 393
rect 270 388 271 392
rect 275 388 276 392
rect 270 387 276 388
rect 398 392 404 393
rect 398 388 399 392
rect 403 388 404 392
rect 398 387 404 388
rect 111 386 115 387
rect 111 381 115 382
rect 135 386 139 387
rect 271 386 275 387
rect 135 381 139 382
rect 162 383 168 384
rect 112 366 114 381
rect 134 380 140 381
rect 134 376 135 380
rect 139 376 140 380
rect 162 379 163 383
rect 167 379 168 383
rect 271 381 275 382
rect 287 386 291 387
rect 287 381 291 382
rect 399 386 403 387
rect 399 381 403 382
rect 479 386 483 387
rect 479 381 483 382
rect 162 378 168 379
rect 286 380 292 381
rect 134 375 140 376
rect 110 365 116 366
rect 110 361 111 365
rect 115 361 116 365
rect 110 360 116 361
rect 142 355 148 356
rect 142 351 143 355
rect 147 351 148 355
rect 142 350 148 351
rect 110 347 116 348
rect 110 343 111 347
rect 115 343 116 347
rect 144 347 146 350
rect 144 345 154 347
rect 110 342 116 343
rect 112 323 114 342
rect 142 335 148 336
rect 142 331 143 335
rect 147 331 148 335
rect 142 330 148 331
rect 144 323 146 330
rect 111 322 115 323
rect 111 317 115 318
rect 143 322 147 323
rect 152 320 154 345
rect 164 328 166 378
rect 286 376 287 380
rect 291 376 292 380
rect 286 375 292 376
rect 478 380 484 381
rect 478 376 479 380
rect 483 376 484 380
rect 478 375 484 376
rect 294 335 300 336
rect 294 331 295 335
rect 299 331 300 335
rect 486 335 492 336
rect 294 330 300 331
rect 315 332 319 333
rect 162 327 168 328
rect 162 323 163 327
rect 167 323 168 327
rect 296 323 298 330
rect 486 331 487 335
rect 491 331 492 335
rect 486 330 492 331
rect 314 327 320 328
rect 314 323 315 327
rect 319 323 320 327
rect 488 323 490 330
rect 504 328 506 402
rect 534 392 540 393
rect 534 388 535 392
rect 539 388 540 392
rect 534 387 540 388
rect 678 392 684 393
rect 678 388 679 392
rect 683 388 684 392
rect 678 387 684 388
rect 830 392 836 393
rect 830 388 831 392
rect 835 388 836 392
rect 830 387 836 388
rect 535 386 539 387
rect 535 381 539 382
rect 671 386 675 387
rect 671 381 675 382
rect 679 386 683 387
rect 679 381 683 382
rect 831 386 835 387
rect 831 381 835 382
rect 670 380 676 381
rect 670 376 671 380
rect 675 376 676 380
rect 670 375 676 376
rect 860 368 862 442
rect 952 424 954 586
rect 1024 582 1026 589
rect 1030 587 1031 591
rect 1035 587 1036 591
rect 1111 589 1115 590
rect 1030 586 1036 587
rect 1022 581 1028 582
rect 1022 577 1023 581
rect 1027 577 1028 581
rect 1022 576 1028 577
rect 1112 570 1114 589
rect 1110 569 1116 570
rect 1110 565 1111 569
rect 1115 565 1116 569
rect 1110 564 1116 565
rect 1022 551 1028 552
rect 1022 547 1023 551
rect 1027 547 1028 551
rect 1022 546 1028 547
rect 1110 551 1116 552
rect 1110 547 1111 551
rect 1115 547 1116 551
rect 1110 546 1116 547
rect 1014 536 1020 537
rect 1014 532 1015 536
rect 1019 532 1020 536
rect 1014 531 1020 532
rect 1016 519 1018 531
rect 991 518 995 519
rect 991 513 995 514
rect 1015 518 1019 519
rect 1015 513 1019 514
rect 990 512 996 513
rect 990 508 991 512
rect 995 508 996 512
rect 990 507 996 508
rect 1024 499 1026 546
rect 1112 519 1114 546
rect 1111 518 1115 519
rect 1111 513 1115 514
rect 1020 497 1026 499
rect 1112 498 1114 513
rect 1110 497 1116 498
rect 998 487 1004 488
rect 998 483 999 487
rect 1003 483 1004 487
rect 998 482 1004 483
rect 1000 475 1002 482
rect 1000 473 1010 475
rect 998 467 1004 468
rect 998 463 999 467
rect 1003 463 1004 467
rect 998 462 1004 463
rect 1000 451 1002 462
rect 999 450 1003 451
rect 1008 448 1010 473
rect 1020 460 1022 497
rect 1110 493 1111 497
rect 1115 493 1116 497
rect 1110 492 1116 493
rect 1110 479 1116 480
rect 1110 475 1111 479
rect 1115 475 1116 479
rect 1110 474 1116 475
rect 1018 459 1024 460
rect 1018 455 1019 459
rect 1023 455 1024 459
rect 1018 454 1024 455
rect 1112 451 1114 474
rect 1111 450 1115 451
rect 999 445 1003 446
rect 1006 447 1012 448
rect 1000 438 1002 445
rect 1006 443 1007 447
rect 1011 443 1012 447
rect 1111 445 1115 446
rect 1006 442 1012 443
rect 998 437 1004 438
rect 998 433 999 437
rect 1003 433 1004 437
rect 998 432 1004 433
rect 1112 426 1114 445
rect 1110 425 1116 426
rect 950 423 956 424
rect 950 419 951 423
rect 955 419 956 423
rect 1110 421 1111 425
rect 1115 421 1116 425
rect 1110 420 1116 421
rect 950 418 956 419
rect 998 407 1004 408
rect 998 403 999 407
rect 1003 403 1004 407
rect 998 402 1004 403
rect 1110 407 1116 408
rect 1110 403 1111 407
rect 1115 403 1116 407
rect 1110 402 1116 403
rect 990 392 996 393
rect 990 388 991 392
rect 995 388 996 392
rect 990 387 996 388
rect 871 386 875 387
rect 871 381 875 382
rect 991 386 995 387
rect 991 381 995 382
rect 870 380 876 381
rect 870 376 871 380
rect 875 376 876 380
rect 870 375 876 376
rect 858 367 864 368
rect 678 363 684 364
rect 678 359 679 363
rect 683 359 684 363
rect 858 363 859 367
rect 863 363 864 367
rect 858 362 864 363
rect 678 358 684 359
rect 558 351 564 352
rect 558 347 559 351
rect 563 347 564 351
rect 558 346 564 347
rect 680 347 682 358
rect 560 333 562 346
rect 680 345 690 347
rect 678 335 684 336
rect 559 332 563 333
rect 678 331 679 335
rect 683 331 684 335
rect 678 330 684 331
rect 502 327 508 328
rect 559 327 563 328
rect 502 323 503 327
rect 507 323 508 327
rect 680 323 682 330
rect 688 328 690 345
rect 878 335 884 336
rect 878 331 879 335
rect 883 331 884 335
rect 878 330 884 331
rect 686 327 692 328
rect 686 323 687 327
rect 691 323 692 327
rect 880 323 882 330
rect 1000 328 1002 402
rect 1112 387 1114 402
rect 1111 386 1115 387
rect 1111 381 1115 382
rect 1112 366 1114 381
rect 1110 365 1116 366
rect 1110 361 1111 365
rect 1115 361 1116 365
rect 1110 360 1116 361
rect 1110 347 1116 348
rect 1110 343 1111 347
rect 1115 343 1116 347
rect 1110 342 1116 343
rect 894 327 900 328
rect 894 323 895 327
rect 899 323 900 327
rect 162 322 168 323
rect 279 322 283 323
rect 143 317 147 318
rect 150 319 156 320
rect 112 298 114 317
rect 144 310 146 317
rect 150 315 151 319
rect 155 315 156 319
rect 279 317 283 318
rect 295 322 299 323
rect 314 322 320 323
rect 455 322 459 323
rect 295 317 299 318
rect 487 322 491 323
rect 502 322 508 323
rect 639 322 643 323
rect 455 317 459 318
rect 462 319 468 320
rect 150 314 156 315
rect 280 310 282 317
rect 286 315 292 316
rect 286 311 287 315
rect 291 311 292 315
rect 286 310 292 311
rect 456 310 458 317
rect 462 315 463 319
rect 467 315 468 319
rect 487 317 491 318
rect 679 322 683 323
rect 686 322 692 323
rect 823 322 827 323
rect 639 317 643 318
rect 646 319 652 320
rect 462 314 468 315
rect 142 309 148 310
rect 142 305 143 309
rect 147 305 148 309
rect 142 304 148 305
rect 278 309 284 310
rect 278 305 279 309
rect 283 305 284 309
rect 278 304 284 305
rect 110 297 116 298
rect 110 293 111 297
rect 115 293 116 297
rect 110 292 116 293
rect 278 291 284 292
rect 288 291 290 310
rect 454 309 460 310
rect 454 305 455 309
rect 459 305 460 309
rect 454 304 460 305
rect 278 287 279 291
rect 283 289 290 291
rect 454 291 460 292
rect 464 291 466 314
rect 640 310 642 317
rect 646 315 647 319
rect 651 315 652 319
rect 679 317 683 318
rect 879 322 883 323
rect 894 322 900 323
rect 998 327 1004 328
rect 998 323 999 327
rect 1003 323 1004 327
rect 1112 323 1114 342
rect 998 322 1004 323
rect 1015 322 1019 323
rect 823 317 827 318
rect 842 319 848 320
rect 646 314 652 315
rect 638 309 644 310
rect 638 305 639 309
rect 643 305 644 309
rect 638 304 644 305
rect 283 287 284 289
rect 278 286 284 287
rect 454 287 455 291
rect 459 289 466 291
rect 638 291 644 292
rect 648 291 650 314
rect 824 310 826 317
rect 842 315 843 319
rect 847 315 848 319
rect 879 317 883 318
rect 842 314 848 315
rect 822 309 828 310
rect 822 305 823 309
rect 827 305 828 309
rect 822 304 828 305
rect 459 287 460 289
rect 454 286 460 287
rect 638 287 639 291
rect 643 289 650 291
rect 643 287 644 289
rect 638 286 644 287
rect 110 279 116 280
rect 110 275 111 279
rect 115 275 116 279
rect 110 274 116 275
rect 570 279 576 280
rect 570 275 571 279
rect 575 275 576 279
rect 570 274 576 275
rect 112 251 114 274
rect 134 264 140 265
rect 134 260 135 264
rect 139 260 140 264
rect 134 259 140 260
rect 270 264 276 265
rect 270 260 271 264
rect 275 260 276 264
rect 270 259 276 260
rect 446 264 452 265
rect 446 260 447 264
rect 451 260 452 264
rect 446 259 452 260
rect 136 251 138 259
rect 272 251 274 259
rect 448 251 450 259
rect 111 250 115 251
rect 111 245 115 246
rect 135 250 139 251
rect 135 245 139 246
rect 271 250 275 251
rect 271 245 275 246
rect 295 250 299 251
rect 295 245 299 246
rect 423 250 427 251
rect 423 245 427 246
rect 447 250 451 251
rect 447 245 451 246
rect 543 250 547 251
rect 543 245 547 246
rect 112 230 114 245
rect 294 244 300 245
rect 294 240 295 244
rect 299 240 300 244
rect 294 239 300 240
rect 422 244 428 245
rect 422 240 423 244
rect 427 240 428 244
rect 422 239 428 240
rect 542 244 548 245
rect 542 240 543 244
rect 547 240 548 244
rect 542 239 548 240
rect 110 229 116 230
rect 110 225 111 229
rect 115 225 116 229
rect 110 224 116 225
rect 362 215 368 216
rect 110 211 116 212
rect 110 207 111 211
rect 115 207 116 211
rect 362 211 363 215
rect 367 211 368 215
rect 362 210 368 211
rect 382 215 388 216
rect 382 211 383 215
rect 387 211 388 215
rect 382 210 388 211
rect 506 215 512 216
rect 506 211 507 215
rect 511 211 512 215
rect 506 210 512 211
rect 110 206 116 207
rect 112 171 114 206
rect 302 199 308 200
rect 302 195 303 199
rect 307 195 308 199
rect 302 194 308 195
rect 304 171 306 194
rect 364 176 366 210
rect 384 184 386 210
rect 430 199 436 200
rect 430 195 431 199
rect 435 195 436 199
rect 430 194 436 195
rect 382 183 388 184
rect 382 179 383 183
rect 387 179 388 183
rect 382 178 388 179
rect 362 175 368 176
rect 362 171 363 175
rect 367 171 368 175
rect 432 171 434 194
rect 508 184 510 210
rect 550 199 556 200
rect 550 195 551 199
rect 555 195 556 199
rect 550 194 556 195
rect 506 183 512 184
rect 506 179 507 183
rect 511 179 512 183
rect 506 178 512 179
rect 552 171 554 194
rect 572 192 574 274
rect 630 264 636 265
rect 630 260 631 264
rect 635 260 636 264
rect 630 259 636 260
rect 814 264 820 265
rect 814 260 815 264
rect 819 260 820 264
rect 814 259 820 260
rect 632 251 634 259
rect 816 251 818 259
rect 631 250 635 251
rect 631 245 635 246
rect 663 250 667 251
rect 663 245 667 246
rect 783 250 787 251
rect 783 245 787 246
rect 815 250 819 251
rect 815 245 819 246
rect 662 244 668 245
rect 662 240 663 244
rect 667 240 668 244
rect 662 239 668 240
rect 782 244 788 245
rect 782 240 783 244
rect 787 240 788 244
rect 782 239 788 240
rect 746 215 752 216
rect 746 211 747 215
rect 751 211 752 215
rect 844 214 846 314
rect 896 296 898 322
rect 1015 317 1019 318
rect 1111 322 1115 323
rect 1111 317 1115 318
rect 1016 310 1018 317
rect 1014 309 1020 310
rect 1014 305 1015 309
rect 1019 305 1020 309
rect 1014 304 1020 305
rect 1112 298 1114 317
rect 1110 297 1116 298
rect 894 295 900 296
rect 894 291 895 295
rect 899 291 900 295
rect 1110 293 1111 297
rect 1115 293 1116 297
rect 1110 292 1116 293
rect 894 290 900 291
rect 938 279 944 280
rect 938 275 939 279
rect 943 275 944 279
rect 938 274 944 275
rect 1110 279 1116 280
rect 1110 275 1111 279
rect 1115 275 1116 279
rect 1110 274 1116 275
rect 911 250 915 251
rect 911 245 915 246
rect 910 244 916 245
rect 910 240 911 244
rect 915 240 916 244
rect 910 239 916 240
rect 850 215 856 216
rect 850 214 851 215
rect 844 212 851 214
rect 746 210 752 211
rect 850 211 851 212
rect 855 211 856 215
rect 850 210 856 211
rect 670 199 676 200
rect 670 195 671 199
rect 675 195 676 199
rect 670 194 676 195
rect 570 191 576 192
rect 570 187 571 191
rect 575 187 576 191
rect 570 186 576 187
rect 672 171 674 194
rect 748 184 750 210
rect 790 199 796 200
rect 790 195 791 199
rect 795 195 796 199
rect 790 194 796 195
rect 918 199 924 200
rect 918 195 919 199
rect 923 195 924 199
rect 918 194 924 195
rect 746 183 752 184
rect 746 179 747 183
rect 751 179 752 183
rect 746 178 752 179
rect 792 171 794 194
rect 826 175 832 176
rect 826 171 827 175
rect 831 171 832 175
rect 920 171 922 194
rect 940 192 942 274
rect 1006 264 1012 265
rect 1006 260 1007 264
rect 1011 260 1012 264
rect 1006 259 1012 260
rect 1008 251 1010 259
rect 1112 251 1114 274
rect 1007 250 1011 251
rect 1007 245 1011 246
rect 1015 250 1019 251
rect 1015 245 1019 246
rect 1111 250 1115 251
rect 1111 245 1115 246
rect 1014 244 1020 245
rect 1014 240 1015 244
rect 1019 240 1020 244
rect 1014 239 1020 240
rect 1112 230 1114 245
rect 1110 229 1116 230
rect 1110 225 1111 229
rect 1115 225 1116 229
rect 1110 224 1116 225
rect 986 215 992 216
rect 986 211 987 215
rect 991 211 992 215
rect 986 210 992 211
rect 1082 215 1088 216
rect 1082 211 1083 215
rect 1087 211 1088 215
rect 1082 210 1088 211
rect 1110 211 1116 212
rect 938 191 944 192
rect 938 187 939 191
rect 943 187 944 191
rect 938 186 944 187
rect 988 184 990 210
rect 1022 199 1028 200
rect 1022 195 1023 199
rect 1027 195 1028 199
rect 1022 194 1028 195
rect 986 183 992 184
rect 986 179 987 183
rect 991 179 992 183
rect 986 178 992 179
rect 1002 175 1008 176
rect 1002 171 1003 175
rect 1007 171 1008 175
rect 1024 171 1026 194
rect 1084 176 1086 210
rect 1110 207 1111 211
rect 1115 207 1116 211
rect 1110 206 1116 207
rect 1082 175 1088 176
rect 1082 171 1083 175
rect 1087 171 1088 175
rect 1112 171 1114 206
rect 111 170 115 171
rect 111 165 115 166
rect 303 170 307 171
rect 303 165 307 166
rect 319 170 323 171
rect 362 170 368 171
rect 407 170 411 171
rect 319 165 323 166
rect 431 170 435 171
rect 407 165 411 166
rect 414 167 420 168
rect 112 146 114 165
rect 320 158 322 165
rect 408 158 410 165
rect 414 163 415 167
rect 419 163 420 167
rect 431 165 435 166
rect 495 170 499 171
rect 551 170 555 171
rect 495 165 499 166
rect 502 167 508 168
rect 414 162 420 163
rect 318 157 324 158
rect 318 153 319 157
rect 323 153 324 157
rect 318 152 324 153
rect 406 157 412 158
rect 406 153 407 157
rect 411 153 412 157
rect 406 152 412 153
rect 416 147 418 162
rect 496 158 498 165
rect 502 163 503 167
rect 507 163 508 167
rect 551 165 555 166
rect 583 170 587 171
rect 671 170 675 171
rect 583 165 587 166
rect 590 167 596 168
rect 502 162 508 163
rect 494 157 500 158
rect 494 153 495 157
rect 499 153 500 157
rect 494 152 500 153
rect 504 147 506 162
rect 584 158 586 165
rect 590 163 591 167
rect 595 163 596 167
rect 759 170 763 171
rect 671 165 675 166
rect 678 167 684 168
rect 590 162 596 163
rect 582 157 588 158
rect 582 153 583 157
rect 587 153 588 157
rect 582 152 588 153
rect 592 147 594 162
rect 672 158 674 165
rect 678 163 679 167
rect 683 163 684 167
rect 791 170 795 171
rect 826 170 832 171
rect 847 170 851 171
rect 759 165 763 166
rect 766 167 772 168
rect 678 162 684 163
rect 670 157 676 158
rect 670 153 671 157
rect 675 153 676 157
rect 670 152 676 153
rect 680 147 682 162
rect 760 158 762 165
rect 766 163 767 167
rect 771 163 772 167
rect 791 165 795 166
rect 766 162 772 163
rect 758 157 764 158
rect 758 153 759 157
rect 763 153 764 157
rect 758 152 764 153
rect 768 147 770 162
rect 110 145 116 146
rect 110 141 111 145
rect 115 141 116 145
rect 110 140 116 141
rect 408 145 418 147
rect 496 145 506 147
rect 584 145 594 147
rect 672 145 682 147
rect 760 145 770 147
rect 408 140 410 145
rect 496 140 498 145
rect 584 140 586 145
rect 672 140 674 145
rect 760 140 762 145
rect 406 139 412 140
rect 406 135 407 139
rect 411 135 412 139
rect 406 134 412 135
rect 494 139 500 140
rect 494 135 495 139
rect 499 135 500 139
rect 494 134 500 135
rect 582 139 588 140
rect 582 135 583 139
rect 587 135 588 139
rect 582 134 588 135
rect 670 139 676 140
rect 670 135 671 139
rect 675 135 676 139
rect 670 134 676 135
rect 758 139 764 140
rect 758 135 759 139
rect 763 135 764 139
rect 758 134 764 135
rect 828 128 830 170
rect 919 170 923 171
rect 847 165 851 166
rect 854 167 860 168
rect 848 158 850 165
rect 854 163 855 167
rect 859 163 860 167
rect 919 165 923 166
rect 935 170 939 171
rect 1002 170 1008 171
rect 1023 170 1027 171
rect 1082 170 1088 171
rect 1111 170 1115 171
rect 935 165 939 166
rect 854 162 860 163
rect 846 157 852 158
rect 846 153 847 157
rect 851 153 852 157
rect 846 152 852 153
rect 856 147 858 162
rect 936 158 938 165
rect 934 157 940 158
rect 934 153 935 157
rect 939 153 940 157
rect 934 152 940 153
rect 848 145 858 147
rect 848 140 850 145
rect 1004 140 1006 170
rect 1023 165 1027 166
rect 1111 165 1115 166
rect 1024 158 1026 165
rect 1022 157 1028 158
rect 1022 153 1023 157
rect 1027 153 1028 157
rect 1022 152 1028 153
rect 1112 146 1114 165
rect 1110 145 1116 146
rect 1110 141 1111 145
rect 1115 141 1116 145
rect 1110 140 1116 141
rect 846 139 852 140
rect 846 135 847 139
rect 851 135 852 139
rect 846 134 852 135
rect 1002 139 1008 140
rect 1002 135 1003 139
rect 1007 135 1008 139
rect 1002 134 1008 135
rect 110 127 116 128
rect 110 123 111 127
rect 115 123 116 127
rect 110 122 116 123
rect 826 127 832 128
rect 826 123 827 127
rect 831 123 832 127
rect 826 122 832 123
rect 1110 127 1116 128
rect 1110 123 1111 127
rect 1115 123 1116 127
rect 1110 122 1116 123
rect 112 107 114 122
rect 310 112 316 113
rect 310 108 311 112
rect 315 108 316 112
rect 310 107 316 108
rect 398 112 404 113
rect 398 108 399 112
rect 403 108 404 112
rect 398 107 404 108
rect 486 112 492 113
rect 486 108 487 112
rect 491 108 492 112
rect 486 107 492 108
rect 574 112 580 113
rect 574 108 575 112
rect 579 108 580 112
rect 574 107 580 108
rect 662 112 668 113
rect 662 108 663 112
rect 667 108 668 112
rect 662 107 668 108
rect 750 112 756 113
rect 750 108 751 112
rect 755 108 756 112
rect 750 107 756 108
rect 838 112 844 113
rect 838 108 839 112
rect 843 108 844 112
rect 838 107 844 108
rect 926 112 932 113
rect 926 108 927 112
rect 931 108 932 112
rect 926 107 932 108
rect 1014 112 1020 113
rect 1014 108 1015 112
rect 1019 108 1020 112
rect 1014 107 1020 108
rect 1112 107 1114 122
rect 111 106 115 107
rect 111 101 115 102
rect 311 106 315 107
rect 311 101 315 102
rect 399 106 403 107
rect 399 101 403 102
rect 487 106 491 107
rect 487 101 491 102
rect 575 106 579 107
rect 575 101 579 102
rect 663 106 667 107
rect 663 101 667 102
rect 751 106 755 107
rect 751 101 755 102
rect 839 106 843 107
rect 839 101 843 102
rect 927 106 931 107
rect 927 101 931 102
rect 1015 106 1019 107
rect 1015 101 1019 102
rect 1111 106 1115 107
rect 1111 101 1115 102
<< m4c >>
rect 111 1218 115 1222
rect 135 1218 139 1222
rect 223 1218 227 1222
rect 311 1218 315 1222
rect 1111 1218 1115 1222
rect 163 1168 167 1172
rect 203 1168 207 1172
rect 251 1168 255 1172
rect 291 1168 295 1172
rect 111 1154 115 1158
rect 143 1154 147 1158
rect 175 1154 179 1158
rect 231 1154 235 1158
rect 263 1154 267 1158
rect 319 1154 323 1158
rect 351 1154 355 1158
rect 439 1154 443 1158
rect 1111 1154 1115 1158
rect 111 1090 115 1094
rect 167 1090 171 1094
rect 255 1090 259 1094
rect 343 1090 347 1094
rect 399 1090 403 1094
rect 431 1090 435 1094
rect 487 1090 491 1094
rect 575 1090 579 1094
rect 663 1090 667 1094
rect 751 1090 755 1094
rect 839 1090 843 1094
rect 927 1090 931 1094
rect 1015 1090 1019 1094
rect 1111 1090 1115 1094
rect 743 1040 747 1044
rect 111 1026 115 1030
rect 407 1026 411 1030
rect 495 1026 499 1030
rect 415 1019 419 1020
rect 415 1016 419 1019
rect 583 1026 587 1030
rect 671 1026 675 1030
rect 759 1026 763 1030
rect 775 1040 779 1044
rect 651 1016 655 1020
rect 679 1019 683 1020
rect 679 1016 683 1019
rect 739 1016 743 1020
rect 847 1026 851 1030
rect 935 1026 939 1030
rect 1023 1026 1027 1030
rect 111 946 115 950
rect 151 946 155 950
rect 271 946 275 950
rect 399 946 403 950
rect 407 946 411 950
rect 487 946 491 950
rect 551 946 555 950
rect 575 946 579 950
rect 663 946 667 950
rect 711 946 715 950
rect 751 946 755 950
rect 839 946 843 950
rect 1111 1026 1115 1030
rect 871 946 875 950
rect 927 946 931 950
rect 1015 946 1019 950
rect 1111 946 1115 950
rect 111 874 115 878
rect 143 874 147 878
rect 159 874 163 878
rect 271 874 275 878
rect 279 874 283 878
rect 415 874 419 878
rect 439 874 443 878
rect 559 874 563 878
rect 631 874 635 878
rect 719 874 723 878
rect 839 874 843 878
rect 879 874 883 878
rect 111 798 115 802
rect 135 798 139 802
rect 239 798 243 802
rect 263 798 267 802
rect 375 798 379 802
rect 431 798 435 802
rect 527 798 531 802
rect 623 798 627 802
rect 695 798 699 802
rect 163 760 167 764
rect 831 798 835 802
rect 863 798 867 802
rect 1023 874 1027 878
rect 1111 874 1115 878
rect 1015 798 1019 802
rect 1111 798 1115 802
rect 291 744 295 748
rect 111 730 115 734
rect 143 730 147 734
rect 247 730 251 734
rect 271 730 275 734
rect 739 760 743 764
rect 683 744 687 748
rect 383 730 387 734
rect 447 730 451 734
rect 535 730 539 734
rect 639 730 643 734
rect 703 730 707 734
rect 831 730 835 734
rect 871 730 875 734
rect 111 666 115 670
rect 263 666 267 670
rect 367 666 371 670
rect 439 666 443 670
rect 463 666 467 670
rect 559 666 563 670
rect 631 666 635 670
rect 663 666 667 670
rect 395 616 399 620
rect 515 600 519 604
rect 111 590 115 594
rect 375 590 379 594
rect 471 590 475 594
rect 495 590 499 594
rect 775 666 779 670
rect 823 666 827 670
rect 1023 730 1027 734
rect 1111 730 1115 734
rect 895 666 899 670
rect 1015 666 1019 670
rect 739 616 743 620
rect 755 600 759 604
rect 567 590 571 594
rect 583 590 587 594
rect 671 590 675 594
rect 759 590 763 594
rect 783 590 787 594
rect 847 590 851 594
rect 903 590 907 594
rect 1111 666 1115 670
rect 935 590 939 594
rect 1023 590 1027 594
rect 111 514 115 518
rect 447 514 451 518
rect 487 514 491 518
rect 543 514 547 518
rect 575 514 579 518
rect 647 514 651 518
rect 663 514 667 518
rect 751 514 755 518
rect 759 514 763 518
rect 839 514 843 518
rect 871 514 875 518
rect 927 514 931 518
rect 475 459 479 460
rect 475 456 479 459
rect 723 456 727 460
rect 111 446 115 450
rect 279 446 283 450
rect 407 446 411 450
rect 455 446 459 450
rect 543 446 547 450
rect 551 446 555 450
rect 655 446 659 450
rect 687 446 691 450
rect 767 446 771 450
rect 839 446 843 450
rect 879 446 883 450
rect 563 432 567 436
rect 611 432 615 436
rect 111 382 115 386
rect 135 382 139 386
rect 271 382 275 386
rect 287 382 291 386
rect 399 382 403 386
rect 479 382 483 386
rect 111 318 115 322
rect 143 318 147 322
rect 315 328 319 332
rect 535 382 539 386
rect 671 382 675 386
rect 679 382 683 386
rect 831 382 835 386
rect 1111 590 1115 594
rect 991 514 995 518
rect 1015 514 1019 518
rect 1111 514 1115 518
rect 999 446 1003 450
rect 1111 446 1115 450
rect 871 382 875 386
rect 991 382 995 386
rect 559 328 563 332
rect 1111 382 1115 386
rect 279 318 283 322
rect 295 318 299 322
rect 455 318 459 322
rect 487 318 491 322
rect 639 318 643 322
rect 679 318 683 322
rect 823 318 827 322
rect 879 318 883 322
rect 111 246 115 250
rect 135 246 139 250
rect 271 246 275 250
rect 295 246 299 250
rect 423 246 427 250
rect 447 246 451 250
rect 543 246 547 250
rect 631 246 635 250
rect 663 246 667 250
rect 783 246 787 250
rect 815 246 819 250
rect 1015 318 1019 322
rect 1111 318 1115 322
rect 911 246 915 250
rect 1007 246 1011 250
rect 1015 246 1019 250
rect 1111 246 1115 250
rect 111 166 115 170
rect 303 166 307 170
rect 319 166 323 170
rect 407 166 411 170
rect 431 166 435 170
rect 495 166 499 170
rect 551 166 555 170
rect 583 166 587 170
rect 671 166 675 170
rect 759 166 763 170
rect 791 166 795 170
rect 847 166 851 170
rect 919 166 923 170
rect 935 166 939 170
rect 1023 166 1027 170
rect 1111 166 1115 170
rect 111 102 115 106
rect 311 102 315 106
rect 399 102 403 106
rect 487 102 491 106
rect 575 102 579 106
rect 663 102 667 106
rect 751 102 755 106
rect 839 102 843 106
rect 927 102 931 106
rect 1015 102 1019 106
rect 1111 102 1115 106
<< m4 >>
rect 84 1217 85 1223
rect 91 1222 1135 1223
rect 91 1218 111 1222
rect 115 1218 135 1222
rect 139 1218 223 1222
rect 227 1218 311 1222
rect 315 1218 1111 1222
rect 1115 1218 1135 1222
rect 91 1217 1135 1218
rect 1141 1217 1142 1223
rect 162 1172 168 1173
rect 202 1172 208 1173
rect 162 1168 163 1172
rect 167 1168 203 1172
rect 207 1168 208 1172
rect 162 1167 168 1168
rect 202 1167 208 1168
rect 250 1172 256 1173
rect 290 1172 296 1173
rect 250 1168 251 1172
rect 255 1168 291 1172
rect 295 1168 296 1172
rect 250 1167 256 1168
rect 290 1167 296 1168
rect 96 1153 97 1159
rect 103 1158 1147 1159
rect 103 1154 111 1158
rect 115 1154 143 1158
rect 147 1154 175 1158
rect 179 1154 231 1158
rect 235 1154 263 1158
rect 267 1154 319 1158
rect 323 1154 351 1158
rect 355 1154 439 1158
rect 443 1154 1111 1158
rect 1115 1154 1147 1158
rect 103 1153 1147 1154
rect 1153 1153 1154 1159
rect 84 1089 85 1095
rect 91 1094 1135 1095
rect 91 1090 111 1094
rect 115 1090 167 1094
rect 171 1090 255 1094
rect 259 1090 343 1094
rect 347 1090 399 1094
rect 403 1090 431 1094
rect 435 1090 487 1094
rect 491 1090 575 1094
rect 579 1090 663 1094
rect 667 1090 751 1094
rect 755 1090 839 1094
rect 843 1090 927 1094
rect 931 1090 1015 1094
rect 1019 1090 1111 1094
rect 1115 1090 1135 1094
rect 91 1089 1135 1090
rect 1141 1089 1142 1095
rect 742 1044 748 1045
rect 774 1044 780 1045
rect 742 1040 743 1044
rect 747 1040 775 1044
rect 779 1040 780 1044
rect 742 1039 748 1040
rect 774 1039 780 1040
rect 96 1025 97 1031
rect 103 1030 1147 1031
rect 103 1026 111 1030
rect 115 1026 407 1030
rect 411 1026 495 1030
rect 499 1026 583 1030
rect 587 1026 671 1030
rect 675 1026 759 1030
rect 763 1026 847 1030
rect 851 1026 935 1030
rect 939 1026 1023 1030
rect 1027 1026 1111 1030
rect 1115 1026 1147 1030
rect 103 1025 1147 1026
rect 1153 1025 1154 1031
rect 414 1020 420 1021
rect 650 1020 656 1021
rect 414 1016 415 1020
rect 419 1016 651 1020
rect 655 1016 656 1020
rect 414 1015 420 1016
rect 650 1015 656 1016
rect 678 1020 684 1021
rect 738 1020 744 1021
rect 678 1016 679 1020
rect 683 1016 739 1020
rect 743 1016 744 1020
rect 678 1015 684 1016
rect 738 1015 744 1016
rect 84 945 85 951
rect 91 950 1135 951
rect 91 946 111 950
rect 115 946 151 950
rect 155 946 271 950
rect 275 946 399 950
rect 403 946 407 950
rect 411 946 487 950
rect 491 946 551 950
rect 555 946 575 950
rect 579 946 663 950
rect 667 946 711 950
rect 715 946 751 950
rect 755 946 839 950
rect 843 946 871 950
rect 875 946 927 950
rect 931 946 1015 950
rect 1019 946 1111 950
rect 1115 946 1135 950
rect 91 945 1135 946
rect 1141 945 1142 951
rect 96 873 97 879
rect 103 878 1147 879
rect 103 874 111 878
rect 115 874 143 878
rect 147 874 159 878
rect 163 874 271 878
rect 275 874 279 878
rect 283 874 415 878
rect 419 874 439 878
rect 443 874 559 878
rect 563 874 631 878
rect 635 874 719 878
rect 723 874 839 878
rect 843 874 879 878
rect 883 874 1023 878
rect 1027 874 1111 878
rect 1115 874 1147 878
rect 103 873 1147 874
rect 1153 873 1154 879
rect 84 797 85 803
rect 91 802 1135 803
rect 91 798 111 802
rect 115 798 135 802
rect 139 798 239 802
rect 243 798 263 802
rect 267 798 375 802
rect 379 798 431 802
rect 435 798 527 802
rect 531 798 623 802
rect 627 798 695 802
rect 699 798 831 802
rect 835 798 863 802
rect 867 798 1015 802
rect 1019 798 1111 802
rect 1115 798 1135 802
rect 91 797 1135 798
rect 1141 797 1142 803
rect 162 764 168 765
rect 738 764 744 765
rect 162 760 163 764
rect 167 760 739 764
rect 743 760 744 764
rect 162 759 168 760
rect 738 759 744 760
rect 290 748 296 749
rect 682 748 688 749
rect 290 744 291 748
rect 295 744 683 748
rect 687 744 688 748
rect 290 743 296 744
rect 682 743 688 744
rect 96 729 97 735
rect 103 734 1147 735
rect 103 730 111 734
rect 115 730 143 734
rect 147 730 247 734
rect 251 730 271 734
rect 275 730 383 734
rect 387 730 447 734
rect 451 730 535 734
rect 539 730 639 734
rect 643 730 703 734
rect 707 730 831 734
rect 835 730 871 734
rect 875 730 1023 734
rect 1027 730 1111 734
rect 1115 730 1147 734
rect 103 729 1147 730
rect 1153 729 1154 735
rect 84 665 85 671
rect 91 670 1135 671
rect 91 666 111 670
rect 115 666 263 670
rect 267 666 367 670
rect 371 666 439 670
rect 443 666 463 670
rect 467 666 559 670
rect 563 666 631 670
rect 635 666 663 670
rect 667 666 775 670
rect 779 666 823 670
rect 827 666 895 670
rect 899 666 1015 670
rect 1019 666 1111 670
rect 1115 666 1135 670
rect 91 665 1135 666
rect 1141 665 1142 671
rect 394 620 400 621
rect 738 620 744 621
rect 394 616 395 620
rect 399 616 739 620
rect 743 616 744 620
rect 394 615 400 616
rect 738 615 744 616
rect 514 604 520 605
rect 754 604 760 605
rect 514 600 515 604
rect 519 600 755 604
rect 759 600 760 604
rect 514 599 520 600
rect 754 599 760 600
rect 96 589 97 595
rect 103 594 1147 595
rect 103 590 111 594
rect 115 590 375 594
rect 379 590 471 594
rect 475 590 495 594
rect 499 590 567 594
rect 571 590 583 594
rect 587 590 671 594
rect 675 590 759 594
rect 763 590 783 594
rect 787 590 847 594
rect 851 590 903 594
rect 907 590 935 594
rect 939 590 1023 594
rect 1027 590 1111 594
rect 1115 590 1147 594
rect 103 589 1147 590
rect 1153 589 1154 595
rect 84 513 85 519
rect 91 518 1135 519
rect 91 514 111 518
rect 115 514 447 518
rect 451 514 487 518
rect 491 514 543 518
rect 547 514 575 518
rect 579 514 647 518
rect 651 514 663 518
rect 667 514 751 518
rect 755 514 759 518
rect 763 514 839 518
rect 843 514 871 518
rect 875 514 927 518
rect 931 514 991 518
rect 995 514 1015 518
rect 1019 514 1111 518
rect 1115 514 1135 518
rect 91 513 1135 514
rect 1141 513 1142 519
rect 474 460 480 461
rect 722 460 728 461
rect 474 456 475 460
rect 479 456 723 460
rect 727 456 728 460
rect 474 455 480 456
rect 722 455 728 456
rect 96 445 97 451
rect 103 450 1147 451
rect 103 446 111 450
rect 115 446 279 450
rect 283 446 407 450
rect 411 446 455 450
rect 459 446 543 450
rect 547 446 551 450
rect 555 446 655 450
rect 659 446 687 450
rect 691 446 767 450
rect 771 446 839 450
rect 843 446 879 450
rect 883 446 999 450
rect 1003 446 1111 450
rect 1115 446 1147 450
rect 103 445 1147 446
rect 1153 445 1154 451
rect 562 436 568 437
rect 610 436 616 437
rect 562 432 563 436
rect 567 432 611 436
rect 615 432 616 436
rect 562 431 568 432
rect 610 431 616 432
rect 84 381 85 387
rect 91 386 1135 387
rect 91 382 111 386
rect 115 382 135 386
rect 139 382 271 386
rect 275 382 287 386
rect 291 382 399 386
rect 403 382 479 386
rect 483 382 535 386
rect 539 382 671 386
rect 675 382 679 386
rect 683 382 831 386
rect 835 382 871 386
rect 875 382 991 386
rect 995 382 1111 386
rect 1115 382 1135 386
rect 91 381 1135 382
rect 1141 381 1142 387
rect 314 332 320 333
rect 558 332 564 333
rect 314 328 315 332
rect 319 328 559 332
rect 563 328 564 332
rect 314 327 320 328
rect 558 327 564 328
rect 96 317 97 323
rect 103 322 1147 323
rect 103 318 111 322
rect 115 318 143 322
rect 147 318 279 322
rect 283 318 295 322
rect 299 318 455 322
rect 459 318 487 322
rect 491 318 639 322
rect 643 318 679 322
rect 683 318 823 322
rect 827 318 879 322
rect 883 318 1015 322
rect 1019 318 1111 322
rect 1115 318 1147 322
rect 103 317 1147 318
rect 1153 317 1154 323
rect 84 245 85 251
rect 91 250 1135 251
rect 91 246 111 250
rect 115 246 135 250
rect 139 246 271 250
rect 275 246 295 250
rect 299 246 423 250
rect 427 246 447 250
rect 451 246 543 250
rect 547 246 631 250
rect 635 246 663 250
rect 667 246 783 250
rect 787 246 815 250
rect 819 246 911 250
rect 915 246 1007 250
rect 1011 246 1015 250
rect 1019 246 1111 250
rect 1115 246 1135 250
rect 91 245 1135 246
rect 1141 245 1142 251
rect 96 165 97 171
rect 103 170 1147 171
rect 103 166 111 170
rect 115 166 303 170
rect 307 166 319 170
rect 323 166 407 170
rect 411 166 431 170
rect 435 166 495 170
rect 499 166 551 170
rect 555 166 583 170
rect 587 166 671 170
rect 675 166 759 170
rect 763 166 791 170
rect 795 166 847 170
rect 851 166 919 170
rect 923 166 935 170
rect 939 166 1023 170
rect 1027 166 1111 170
rect 1115 166 1147 170
rect 103 165 1147 166
rect 1153 165 1154 171
rect 84 101 85 107
rect 91 106 1135 107
rect 91 102 111 106
rect 115 102 311 106
rect 315 102 399 106
rect 403 102 487 106
rect 491 102 575 106
rect 579 102 663 106
rect 667 102 751 106
rect 755 102 839 106
rect 843 102 927 106
rect 931 102 1015 106
rect 1019 102 1111 106
rect 1115 102 1135 106
rect 91 101 1135 102
rect 1141 101 1142 107
<< m5c >>
rect 85 1217 91 1223
rect 1135 1217 1141 1223
rect 97 1153 103 1159
rect 1147 1153 1153 1159
rect 85 1089 91 1095
rect 1135 1089 1141 1095
rect 97 1025 103 1031
rect 1147 1025 1153 1031
rect 85 945 91 951
rect 1135 945 1141 951
rect 97 873 103 879
rect 1147 873 1153 879
rect 85 797 91 803
rect 1135 797 1141 803
rect 97 729 103 735
rect 1147 729 1153 735
rect 85 665 91 671
rect 1135 665 1141 671
rect 97 589 103 595
rect 1147 589 1153 595
rect 85 513 91 519
rect 1135 513 1141 519
rect 97 445 103 451
rect 1147 445 1153 451
rect 85 381 91 387
rect 1135 381 1141 387
rect 97 317 103 323
rect 1147 317 1153 323
rect 85 245 91 251
rect 1135 245 1141 251
rect 97 165 103 171
rect 1147 165 1153 171
rect 85 101 91 107
rect 1135 101 1141 107
<< m5 >>
rect 84 1223 92 1224
rect 84 1217 85 1223
rect 91 1217 92 1223
rect 84 1095 92 1217
rect 84 1089 85 1095
rect 91 1089 92 1095
rect 84 951 92 1089
rect 84 945 85 951
rect 91 945 92 951
rect 84 803 92 945
rect 84 797 85 803
rect 91 797 92 803
rect 84 671 92 797
rect 84 665 85 671
rect 91 665 92 671
rect 84 519 92 665
rect 84 513 85 519
rect 91 513 92 519
rect 84 387 92 513
rect 84 381 85 387
rect 91 381 92 387
rect 84 251 92 381
rect 84 245 85 251
rect 91 245 92 251
rect 84 107 92 245
rect 84 101 85 107
rect 91 101 92 107
rect 84 72 92 101
rect 96 1159 104 1224
rect 96 1153 97 1159
rect 103 1153 104 1159
rect 96 1031 104 1153
rect 96 1025 97 1031
rect 103 1025 104 1031
rect 96 879 104 1025
rect 96 873 97 879
rect 103 873 104 879
rect 96 735 104 873
rect 96 729 97 735
rect 103 729 104 735
rect 96 595 104 729
rect 96 589 97 595
rect 103 589 104 595
rect 96 451 104 589
rect 96 445 97 451
rect 103 445 104 451
rect 96 323 104 445
rect 96 317 97 323
rect 103 317 104 323
rect 96 171 104 317
rect 96 165 97 171
rect 103 165 104 171
rect 96 72 104 165
rect 1134 1223 1142 1224
rect 1134 1217 1135 1223
rect 1141 1217 1142 1223
rect 1134 1095 1142 1217
rect 1134 1089 1135 1095
rect 1141 1089 1142 1095
rect 1134 951 1142 1089
rect 1134 945 1135 951
rect 1141 945 1142 951
rect 1134 803 1142 945
rect 1134 797 1135 803
rect 1141 797 1142 803
rect 1134 671 1142 797
rect 1134 665 1135 671
rect 1141 665 1142 671
rect 1134 519 1142 665
rect 1134 513 1135 519
rect 1141 513 1142 519
rect 1134 387 1142 513
rect 1134 381 1135 387
rect 1141 381 1142 387
rect 1134 251 1142 381
rect 1134 245 1135 251
rect 1141 245 1142 251
rect 1134 107 1142 245
rect 1134 101 1135 107
rect 1141 101 1142 107
rect 1134 72 1142 101
rect 1146 1159 1154 1224
rect 1146 1153 1147 1159
rect 1153 1153 1154 1159
rect 1146 1031 1154 1153
rect 1146 1025 1147 1031
rect 1153 1025 1154 1031
rect 1146 879 1154 1025
rect 1146 873 1147 879
rect 1153 873 1154 879
rect 1146 735 1154 873
rect 1146 729 1147 735
rect 1153 729 1154 735
rect 1146 595 1154 729
rect 1146 589 1147 595
rect 1153 589 1154 595
rect 1146 451 1154 589
rect 1146 445 1147 451
rect 1153 445 1154 451
rect 1146 323 1154 445
rect 1146 317 1147 323
rect 1153 317 1154 323
rect 1146 171 1154 317
rect 1146 165 1147 171
rect 1153 165 1154 171
rect 1146 72 1154 165
use welltap_svt  __well_tap__0
timestamp 1731001260
transform 1 0 104 0 1 120
box 8 4 12 24
use circuitppnp  ppnps
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use circuitwell  npwells
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use welltap_svt  __well_tap__0
timestamp 1731001260
transform 1 0 104 0 1 120
box 8 4 12 24
use circuitppnp  ppnps
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use circuitwell  npwells
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use _0_0std_0_0cells_0_0MUX2X1  mux_566_6
timestamp 1731001260
transform 1 0 304 0 1 104
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_566_6
timestamp 1731001260
transform 1 0 304 0 1 104
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_567_6
timestamp 1731001260
transform 1 0 392 0 1 104
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_567_6
timestamp 1731001260
transform 1 0 392 0 1 104
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_568_6
timestamp 1731001260
transform 1 0 480 0 1 104
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_568_6
timestamp 1731001260
transform 1 0 480 0 1 104
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_569_6
timestamp 1731001260
transform 1 0 568 0 1 104
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_569_6
timestamp 1731001260
transform 1 0 568 0 1 104
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_570_6
timestamp 1731001260
transform 1 0 656 0 1 104
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_570_6
timestamp 1731001260
transform 1 0 656 0 1 104
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_571_6
timestamp 1731001260
transform 1 0 744 0 1 104
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_571_6
timestamp 1731001260
transform 1 0 744 0 1 104
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_572_6
timestamp 1731001260
transform 1 0 832 0 1 104
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_572_6
timestamp 1731001260
transform 1 0 832 0 1 104
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_599_6
timestamp 1731001260
transform 1 0 920 0 1 104
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_599_6
timestamp 1731001260
transform 1 0 920 0 1 104
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_598_6
timestamp 1731001260
transform 1 0 1008 0 1 104
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_598_6
timestamp 1731001260
transform 1 0 1008 0 1 104
box 8 2 80 63
use welltap_svt  __well_tap__1
timestamp 1731001260
transform 1 0 1104 0 1 120
box 8 4 12 24
use welltap_svt  __well_tap__1
timestamp 1731001260
transform 1 0 1104 0 1 120
box 8 4 12 24
use _0_0std_0_0cells_0_0MUX2X1  mux_565_6
timestamp 1731001260
transform 1 0 288 0 -1 248
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_565_6
timestamp 1731001260
transform 1 0 288 0 -1 248
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_564_6
timestamp 1731001260
transform 1 0 416 0 -1 248
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_564_6
timestamp 1731001260
transform 1 0 416 0 -1 248
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_563_6
timestamp 1731001260
transform 1 0 536 0 -1 248
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_563_6
timestamp 1731001260
transform 1 0 536 0 -1 248
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_573_6
timestamp 1731001260
transform 1 0 656 0 -1 248
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_573_6
timestamp 1731001260
transform 1 0 656 0 -1 248
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_574_6
timestamp 1731001260
transform 1 0 776 0 -1 248
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_574_6
timestamp 1731001260
transform 1 0 776 0 -1 248
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_596_6
timestamp 1731001260
transform 1 0 904 0 -1 248
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_596_6
timestamp 1731001260
transform 1 0 904 0 -1 248
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_597_6
timestamp 1731001260
transform 1 0 1008 0 -1 248
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_597_6
timestamp 1731001260
transform 1 0 1008 0 -1 248
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_559_6
timestamp 1731001260
transform 1 0 128 0 1 256
box 8 2 80 63
use welltap_svt  __well_tap__2
timestamp 1731001260
transform 1 0 104 0 -1 232
box 8 4 12 24
use _0_0std_0_0cells_0_0MUX2X1  mux_559_6
timestamp 1731001260
transform 1 0 128 0 1 256
box 8 2 80 63
use welltap_svt  __well_tap__2
timestamp 1731001260
transform 1 0 104 0 -1 232
box 8 4 12 24
use _0_0std_0_0cells_0_0MUX2X1  mux_560_6
timestamp 1731001260
transform 1 0 264 0 1 256
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_560_6
timestamp 1731001260
transform 1 0 264 0 1 256
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_561_6
timestamp 1731001260
transform 1 0 440 0 1 256
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_561_6
timestamp 1731001260
transform 1 0 440 0 1 256
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_562_6
timestamp 1731001260
transform 1 0 624 0 1 256
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_562_6
timestamp 1731001260
transform 1 0 624 0 1 256
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_575_6
timestamp 1731001260
transform 1 0 808 0 1 256
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_575_6
timestamp 1731001260
transform 1 0 808 0 1 256
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_595_6
timestamp 1731001260
transform 1 0 1000 0 1 256
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_595_6
timestamp 1731001260
transform 1 0 1000 0 1 256
box 8 2 80 63
use welltap_svt  __well_tap__3
timestamp 1731001260
transform 1 0 1104 0 -1 232
box 8 4 12 24
use welltap_svt  __well_tap__3
timestamp 1731001260
transform 1 0 1104 0 -1 232
box 8 4 12 24
use _0_0std_0_0cells_0_0MUX2X1  mux_558_6
timestamp 1731001260
transform 1 0 128 0 -1 384
box 8 2 80 63
use welltap_svt  __well_tap__4
timestamp 1731001260
transform 1 0 104 0 1 272
box 8 4 12 24
use _0_0std_0_0cells_0_0MUX2X1  mux_558_6
timestamp 1731001260
transform 1 0 128 0 -1 384
box 8 2 80 63
use welltap_svt  __well_tap__4
timestamp 1731001260
transform 1 0 104 0 1 272
box 8 4 12 24
use _0_0std_0_0cells_0_0MUX2X1  mux_557_6
timestamp 1731001260
transform 1 0 280 0 -1 384
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_557_6
timestamp 1731001260
transform 1 0 280 0 -1 384
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_555_6
timestamp 1731001260
transform 1 0 472 0 -1 384
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_555_6
timestamp 1731001260
transform 1 0 472 0 -1 384
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_556_6
timestamp 1731001260
transform 1 0 664 0 -1 384
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_556_6
timestamp 1731001260
transform 1 0 664 0 -1 384
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_576_6
timestamp 1731001260
transform 1 0 864 0 -1 384
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_576_6
timestamp 1731001260
transform 1 0 864 0 -1 384
box 8 2 80 63
use welltap_svt  __well_tap__5
timestamp 1731001260
transform 1 0 1104 0 1 272
box 8 4 12 24
use welltap_svt  __well_tap__5
timestamp 1731001260
transform 1 0 1104 0 1 272
box 8 4 12 24
use welltap_svt  __well_tap__6
timestamp 1731001260
transform 1 0 104 0 -1 368
box 8 4 12 24
use welltap_svt  __well_tap__8
timestamp 1731001260
transform 1 0 104 0 1 400
box 8 4 12 24
use welltap_svt  __well_tap__6
timestamp 1731001260
transform 1 0 104 0 -1 368
box 8 4 12 24
use welltap_svt  __well_tap__8
timestamp 1731001260
transform 1 0 104 0 1 400
box 8 4 12 24
use _0_0std_0_0cells_0_0MUX2X1  mux_553_6
timestamp 1731001260
transform 1 0 264 0 1 384
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_553_6
timestamp 1731001260
transform 1 0 264 0 1 384
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_554_6
timestamp 1731001260
transform 1 0 392 0 1 384
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_554_6
timestamp 1731001260
transform 1 0 392 0 1 384
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_552_6
timestamp 1731001260
transform 1 0 528 0 1 384
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_552_6
timestamp 1731001260
transform 1 0 528 0 1 384
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_551_6
timestamp 1731001260
transform 1 0 672 0 1 384
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_551_6
timestamp 1731001260
transform 1 0 672 0 1 384
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_577_6
timestamp 1731001260
transform 1 0 824 0 1 384
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_577_6
timestamp 1731001260
transform 1 0 824 0 1 384
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_594_6
timestamp 1731001260
transform 1 0 984 0 1 384
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_594_6
timestamp 1731001260
transform 1 0 984 0 1 384
box 8 2 80 63
use welltap_svt  __well_tap__7
timestamp 1731001260
transform 1 0 1104 0 -1 368
box 8 4 12 24
use welltap_svt  __well_tap__9
timestamp 1731001260
transform 1 0 1104 0 1 400
box 8 4 12 24
use welltap_svt  __well_tap__7
timestamp 1731001260
transform 1 0 1104 0 -1 368
box 8 4 12 24
use welltap_svt  __well_tap__9
timestamp 1731001260
transform 1 0 1104 0 1 400
box 8 4 12 24
use _0_0std_0_0cells_0_0MUX2X1  mux_548_6
timestamp 1731001260
transform 1 0 440 0 -1 516
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_548_6
timestamp 1731001260
transform 1 0 440 0 -1 516
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_549_6
timestamp 1731001260
transform 1 0 536 0 -1 516
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_549_6
timestamp 1731001260
transform 1 0 536 0 -1 516
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_550_6
timestamp 1731001260
transform 1 0 640 0 -1 516
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_550_6
timestamp 1731001260
transform 1 0 640 0 -1 516
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_547_6
timestamp 1731001260
transform 1 0 752 0 -1 516
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_547_6
timestamp 1731001260
transform 1 0 752 0 -1 516
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_546_6
timestamp 1731001260
transform 1 0 864 0 -1 516
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_546_6
timestamp 1731001260
transform 1 0 864 0 -1 516
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_593_6
timestamp 1731001260
transform 1 0 984 0 -1 516
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_593_6
timestamp 1731001260
transform 1 0 984 0 -1 516
box 8 2 80 63
use welltap_svt  __well_tap__10
timestamp 1731001260
transform 1 0 104 0 -1 500
box 8 4 12 24
use welltap_svt  __well_tap__10
timestamp 1731001260
transform 1 0 104 0 -1 500
box 8 4 12 24
use _0_0std_0_0cells_0_0MUX2X1  mux_541_6
timestamp 1731001260
transform 1 0 480 0 1 528
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_541_6
timestamp 1731001260
transform 1 0 480 0 1 528
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_542_6
timestamp 1731001260
transform 1 0 568 0 1 528
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_542_6
timestamp 1731001260
transform 1 0 568 0 1 528
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_543_6
timestamp 1731001260
transform 1 0 656 0 1 528
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_543_6
timestamp 1731001260
transform 1 0 656 0 1 528
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_544_6
timestamp 1731001260
transform 1 0 744 0 1 528
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_544_6
timestamp 1731001260
transform 1 0 744 0 1 528
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_545_6
timestamp 1731001260
transform 1 0 832 0 1 528
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_545_6
timestamp 1731001260
transform 1 0 832 0 1 528
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_578_6
timestamp 1731001260
transform 1 0 920 0 1 528
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_578_6
timestamp 1731001260
transform 1 0 920 0 1 528
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_592_6
timestamp 1731001260
transform 1 0 1008 0 1 528
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_592_6
timestamp 1731001260
transform 1 0 1008 0 1 528
box 8 2 80 63
use welltap_svt  __well_tap__11
timestamp 1731001260
transform 1 0 1104 0 -1 500
box 8 4 12 24
use welltap_svt  __well_tap__11
timestamp 1731001260
transform 1 0 1104 0 -1 500
box 8 4 12 24
use welltap_svt  __well_tap__12
timestamp 1731001260
transform 1 0 104 0 1 544
box 8 4 12 24
use welltap_svt  __well_tap__12
timestamp 1731001260
transform 1 0 104 0 1 544
box 8 4 12 24
use _0_0std_0_0cells_0_0MUX2X1  mux_536_6
timestamp 1731001260
transform 1 0 360 0 -1 668
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_536_6
timestamp 1731001260
transform 1 0 360 0 -1 668
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_537_6
timestamp 1731001260
transform 1 0 456 0 -1 668
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_537_6
timestamp 1731001260
transform 1 0 456 0 -1 668
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_538_6
timestamp 1731001260
transform 1 0 552 0 -1 668
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_538_6
timestamp 1731001260
transform 1 0 552 0 -1 668
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_539_6
timestamp 1731001260
transform 1 0 656 0 -1 668
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_539_6
timestamp 1731001260
transform 1 0 656 0 -1 668
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_540_6
timestamp 1731001260
transform 1 0 768 0 -1 668
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_540_6
timestamp 1731001260
transform 1 0 768 0 -1 668
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_579_6
timestamp 1731001260
transform 1 0 888 0 -1 668
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_579_6
timestamp 1731001260
transform 1 0 888 0 -1 668
box 8 2 80 63
use welltap_svt  __well_tap__13
timestamp 1731001260
transform 1 0 1104 0 1 544
box 8 4 12 24
use welltap_svt  __well_tap__13
timestamp 1731001260
transform 1 0 1104 0 1 544
box 8 4 12 24
use welltap_svt  __well_tap__14
timestamp 1731001260
transform 1 0 104 0 -1 652
box 8 4 12 24
use welltap_svt  __well_tap__14
timestamp 1731001260
transform 1 0 104 0 -1 652
box 8 4 12 24
use _0_0std_0_0cells_0_0MUX2X1  mux_532_6
timestamp 1731001260
transform 1 0 256 0 1 668
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_532_6
timestamp 1731001260
transform 1 0 256 0 1 668
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_533_6
timestamp 1731001260
transform 1 0 432 0 1 668
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_533_6
timestamp 1731001260
transform 1 0 432 0 1 668
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_534_6
timestamp 1731001260
transform 1 0 624 0 1 668
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_534_6
timestamp 1731001260
transform 1 0 624 0 1 668
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_535_6
timestamp 1731001260
transform 1 0 816 0 1 668
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_535_6
timestamp 1731001260
transform 1 0 816 0 1 668
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_591_6
timestamp 1731001260
transform 1 0 1008 0 1 668
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_591_6
timestamp 1731001260
transform 1 0 1008 0 1 668
box 8 2 80 63
use welltap_svt  __well_tap__15
timestamp 1731001260
transform 1 0 1104 0 -1 652
box 8 4 12 24
use welltap_svt  __well_tap__15
timestamp 1731001260
transform 1 0 1104 0 -1 652
box 8 4 12 24
use _0_0std_0_0cells_0_0MUX2X1  mux_527_6
timestamp 1731001260
transform 1 0 128 0 -1 800
box 8 2 80 63
use welltap_svt  __well_tap__16
timestamp 1731001260
transform 1 0 104 0 1 684
box 8 4 12 24
use _0_0std_0_0cells_0_0MUX2X1  mux_527_6
timestamp 1731001260
transform 1 0 128 0 -1 800
box 8 2 80 63
use welltap_svt  __well_tap__16
timestamp 1731001260
transform 1 0 104 0 1 684
box 8 4 12 24
use _0_0std_0_0cells_0_0MUX2X1  mux_528_6
timestamp 1731001260
transform 1 0 232 0 -1 800
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_528_6
timestamp 1731001260
transform 1 0 232 0 -1 800
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_529_6
timestamp 1731001260
transform 1 0 368 0 -1 800
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_529_6
timestamp 1731001260
transform 1 0 368 0 -1 800
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_530_6
timestamp 1731001260
transform 1 0 520 0 -1 800
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_530_6
timestamp 1731001260
transform 1 0 520 0 -1 800
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_531_6
timestamp 1731001260
transform 1 0 688 0 -1 800
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_531_6
timestamp 1731001260
transform 1 0 688 0 -1 800
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_580_6
timestamp 1731001260
transform 1 0 856 0 -1 800
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_580_6
timestamp 1731001260
transform 1 0 856 0 -1 800
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_590_6
timestamp 1731001260
transform 1 0 1008 0 -1 800
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_590_6
timestamp 1731001260
transform 1 0 1008 0 -1 800
box 8 2 80 63
use welltap_svt  __well_tap__17
timestamp 1731001260
transform 1 0 1104 0 1 684
box 8 4 12 24
use welltap_svt  __well_tap__17
timestamp 1731001260
transform 1 0 1104 0 1 684
box 8 4 12 24
use welltap_svt  __well_tap__18
timestamp 1731001260
transform 1 0 104 0 -1 784
box 8 4 12 24
use welltap_svt  __well_tap__18
timestamp 1731001260
transform 1 0 104 0 -1 784
box 8 4 12 24
use welltap_svt  __well_tap__19
timestamp 1731001260
transform 1 0 1104 0 -1 784
box 8 4 12 24
use welltap_svt  __well_tap__19
timestamp 1731001260
transform 1 0 1104 0 -1 784
box 8 4 12 24
use _0_0std_0_0cells_0_0MUX2X1  mux_522_6
timestamp 1731001260
transform 1 0 128 0 1 812
box 8 2 80 63
use welltap_svt  __well_tap__20
timestamp 1731001260
transform 1 0 104 0 1 828
box 8 4 12 24
use _0_0std_0_0cells_0_0MUX2X1  mux_522_6
timestamp 1731001260
transform 1 0 128 0 1 812
box 8 2 80 63
use welltap_svt  __well_tap__20
timestamp 1731001260
transform 1 0 104 0 1 828
box 8 4 12 24
use _0_0std_0_0cells_0_0MUX2X1  mux_523_6
timestamp 1731001260
transform 1 0 256 0 1 812
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_523_6
timestamp 1731001260
transform 1 0 256 0 1 812
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_524_6
timestamp 1731001260
transform 1 0 424 0 1 812
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_524_6
timestamp 1731001260
transform 1 0 424 0 1 812
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_525_6
timestamp 1731001260
transform 1 0 616 0 1 812
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_525_6
timestamp 1731001260
transform 1 0 616 0 1 812
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_526_6
timestamp 1731001260
transform 1 0 824 0 1 812
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_526_6
timestamp 1731001260
transform 1 0 824 0 1 812
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_589_6
timestamp 1731001260
transform 1 0 1008 0 1 812
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_589_6
timestamp 1731001260
transform 1 0 1008 0 1 812
box 8 2 80 63
use welltap_svt  __well_tap__21
timestamp 1731001260
transform 1 0 1104 0 1 828
box 8 4 12 24
use welltap_svt  __well_tap__21
timestamp 1731001260
transform 1 0 1104 0 1 828
box 8 4 12 24
use _0_0std_0_0cells_0_0MUX2X1  mux_521_6
timestamp 1731001260
transform 1 0 144 0 -1 948
box 8 2 80 63
use welltap_svt  __well_tap__22
timestamp 1731001260
transform 1 0 104 0 -1 932
box 8 4 12 24
use _0_0std_0_0cells_0_0MUX2X1  mux_521_6
timestamp 1731001260
transform 1 0 144 0 -1 948
box 8 2 80 63
use welltap_svt  __well_tap__22
timestamp 1731001260
transform 1 0 104 0 -1 932
box 8 4 12 24
use _0_0std_0_0cells_0_0MUX2X1  mux_520_6
timestamp 1731001260
transform 1 0 264 0 -1 948
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_520_6
timestamp 1731001260
transform 1 0 264 0 -1 948
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_519_6
timestamp 1731001260
transform 1 0 400 0 -1 948
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_519_6
timestamp 1731001260
transform 1 0 400 0 -1 948
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_518_6
timestamp 1731001260
transform 1 0 544 0 -1 948
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_518_6
timestamp 1731001260
transform 1 0 544 0 -1 948
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_517_6
timestamp 1731001260
transform 1 0 704 0 -1 948
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_517_6
timestamp 1731001260
transform 1 0 704 0 -1 948
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_581_6
timestamp 1731001260
transform 1 0 864 0 -1 948
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_581_6
timestamp 1731001260
transform 1 0 864 0 -1 948
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_588_6
timestamp 1731001260
transform 1 0 1008 0 -1 948
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_588_6
timestamp 1731001260
transform 1 0 1008 0 -1 948
box 8 2 80 63
use welltap_svt  __well_tap__23
timestamp 1731001260
transform 1 0 1104 0 -1 932
box 8 4 12 24
use welltap_svt  __well_tap__23
timestamp 1731001260
transform 1 0 1104 0 -1 932
box 8 4 12 24
use welltap_svt  __well_tap__24
timestamp 1731001260
transform 1 0 104 0 1 980
box 8 4 12 24
use welltap_svt  __well_tap__24
timestamp 1731001260
transform 1 0 104 0 1 980
box 8 4 12 24
use _0_0std_0_0cells_0_0MUX2X1  mux_514_6
timestamp 1731001260
transform 1 0 392 0 1 964
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_514_6
timestamp 1731001260
transform 1 0 392 0 1 964
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_515_6
timestamp 1731001260
transform 1 0 480 0 1 964
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_515_6
timestamp 1731001260
transform 1 0 480 0 1 964
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_516_6
timestamp 1731001260
transform 1 0 568 0 1 964
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_516_6
timestamp 1731001260
transform 1 0 568 0 1 964
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_513_6
timestamp 1731001260
transform 1 0 656 0 1 964
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_513_6
timestamp 1731001260
transform 1 0 656 0 1 964
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_512_6
timestamp 1731001260
transform 1 0 744 0 1 964
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_512_6
timestamp 1731001260
transform 1 0 744 0 1 964
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_582_6
timestamp 1731001260
transform 1 0 832 0 1 964
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_582_6
timestamp 1731001260
transform 1 0 832 0 1 964
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_586_6
timestamp 1731001260
transform 1 0 920 0 1 964
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_586_6
timestamp 1731001260
transform 1 0 920 0 1 964
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_587_6
timestamp 1731001260
transform 1 0 1008 0 1 964
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_587_6
timestamp 1731001260
transform 1 0 1008 0 1 964
box 8 2 80 63
use welltap_svt  __well_tap__25
timestamp 1731001260
transform 1 0 1104 0 1 980
box 8 4 12 24
use welltap_svt  __well_tap__25
timestamp 1731001260
transform 1 0 1104 0 1 980
box 8 4 12 24
use welltap_svt  __well_tap__26
timestamp 1731001260
transform 1 0 104 0 -1 1076
box 8 4 12 24
use welltap_svt  __well_tap__26
timestamp 1731001260
transform 1 0 104 0 -1 1076
box 8 4 12 24
use _0_0std_0_0cells_0_0MUX2X1  mux_57_6
timestamp 1731001260
transform 1 0 392 0 -1 1092
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_57_6
timestamp 1731001260
transform 1 0 392 0 -1 1092
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_58_6
timestamp 1731001260
transform 1 0 480 0 -1 1092
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_58_6
timestamp 1731001260
transform 1 0 480 0 -1 1092
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_59_6
timestamp 1731001260
transform 1 0 568 0 -1 1092
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_59_6
timestamp 1731001260
transform 1 0 568 0 -1 1092
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_510_6
timestamp 1731001260
transform 1 0 656 0 -1 1092
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_510_6
timestamp 1731001260
transform 1 0 656 0 -1 1092
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_511_6
timestamp 1731001260
transform 1 0 744 0 -1 1092
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_511_6
timestamp 1731001260
transform 1 0 744 0 -1 1092
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_583_6
timestamp 1731001260
transform 1 0 832 0 -1 1092
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_583_6
timestamp 1731001260
transform 1 0 832 0 -1 1092
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_584_6
timestamp 1731001260
transform 1 0 920 0 -1 1092
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_584_6
timestamp 1731001260
transform 1 0 920 0 -1 1092
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_585_6
timestamp 1731001260
transform 1 0 1008 0 -1 1092
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_585_6
timestamp 1731001260
transform 1 0 1008 0 -1 1092
box 8 2 80 63
use welltap_svt  __well_tap__27
timestamp 1731001260
transform 1 0 1104 0 -1 1076
box 8 4 12 24
use welltap_svt  __well_tap__27
timestamp 1731001260
transform 1 0 1104 0 -1 1076
box 8 4 12 24
use welltap_svt  __well_tap__28
timestamp 1731001260
transform 1 0 104 0 1 1108
box 8 4 12 24
use welltap_svt  __well_tap__28
timestamp 1731001260
transform 1 0 104 0 1 1108
box 8 4 12 24
use _0_0std_0_0cells_0_0MUX2X1  mux_53_6
timestamp 1731001260
transform 1 0 160 0 1 1092
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_53_6
timestamp 1731001260
transform 1 0 160 0 1 1092
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_54_6
timestamp 1731001260
transform 1 0 248 0 1 1092
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_54_6
timestamp 1731001260
transform 1 0 248 0 1 1092
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_55_6
timestamp 1731001260
transform 1 0 336 0 1 1092
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_55_6
timestamp 1731001260
transform 1 0 336 0 1 1092
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_56_6
timestamp 1731001260
transform 1 0 424 0 1 1092
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_56_6
timestamp 1731001260
transform 1 0 424 0 1 1092
box 8 2 80 63
use welltap_svt  __well_tap__29
timestamp 1731001260
transform 1 0 1104 0 1 1108
box 8 4 12 24
use welltap_svt  __well_tap__29
timestamp 1731001260
transform 1 0 1104 0 1 1108
box 8 4 12 24
use _0_0std_0_0cells_0_0MUX2X1  mux_52_6
timestamp 1731001260
transform 1 0 128 0 -1 1220
box 8 2 80 63
use welltap_svt  __well_tap__30
timestamp 1731001260
transform 1 0 104 0 -1 1204
box 8 4 12 24
use _0_0std_0_0cells_0_0MUX2X1  mux_52_6
timestamp 1731001260
transform 1 0 128 0 -1 1220
box 8 2 80 63
use welltap_svt  __well_tap__30
timestamp 1731001260
transform 1 0 104 0 -1 1204
box 8 4 12 24
use _0_0std_0_0cells_0_0MUX2X1  mux_51_6
timestamp 1731001260
transform 1 0 216 0 -1 1220
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_51_6
timestamp 1731001260
transform 1 0 216 0 -1 1220
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_50_6
timestamp 1731001260
transform 1 0 304 0 -1 1220
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_50_6
timestamp 1731001260
transform 1 0 304 0 -1 1220
box 8 2 80 63
use welltap_svt  __well_tap__31
timestamp 1731001260
transform 1 0 1104 0 -1 1204
box 8 4 12 24
use welltap_svt  __well_tap__31
timestamp 1731001260
transform 1 0 1104 0 -1 1204
box 8 4 12 24
<< end >>
