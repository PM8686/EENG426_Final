magic
tech sky130l
timestamp 1731220634
<< m1 >>
rect 1400 2119 1404 2135
rect 1448 2119 1452 2135
rect 1496 2119 1500 2135
rect 1552 2119 1556 2135
rect 1656 2119 1660 2135
rect 1864 2119 1868 2135
rect 1704 2011 1708 2027
rect 712 1967 716 1999
rect 2104 1991 2108 2027
rect 624 1939 628 1955
rect 688 1939 692 1955
rect 752 1939 756 1955
rect 808 1939 812 1955
rect 952 1939 956 1955
rect 1192 1903 1196 1919
rect 1568 1903 1572 1919
rect 1648 1903 1652 1919
rect 1816 1903 1820 1919
rect 1912 1903 1916 1919
rect 1536 1859 1540 1883
rect 368 1831 372 1847
rect 536 1831 540 1847
rect 584 1831 588 1847
rect 632 1831 636 1847
rect 680 1831 684 1847
rect 728 1831 732 1847
rect 248 1783 252 1799
rect 416 1783 420 1799
rect 1680 1795 1684 1811
rect 384 1719 388 1735
rect 512 1719 516 1735
rect 720 1719 724 1735
rect 400 1675 404 1691
rect 496 1675 500 1691
rect 2056 1691 2060 1707
rect 296 1607 300 1623
rect 376 1607 380 1623
rect 456 1607 460 1623
rect 992 1607 996 1623
rect 208 1567 212 1583
rect 216 1503 220 1563
rect 288 1531 292 1583
rect 336 1567 340 1583
rect 408 1567 412 1583
rect 632 1567 636 1583
rect 1496 1571 1500 1587
rect 1832 1571 1836 1587
rect 2104 1551 2108 1587
rect 1856 1531 1860 1547
rect 1944 1531 1948 1547
rect 264 1503 268 1519
rect 344 1503 348 1519
rect 424 1503 428 1519
rect 600 1503 604 1519
rect 688 1503 692 1519
rect 312 1463 316 1479
rect 1520 1467 1524 1483
rect 1656 1467 1660 1483
rect 1736 1467 1740 1483
rect 1808 1467 1812 1483
rect 1768 1423 1772 1439
rect 1840 1423 1844 1439
rect 368 1399 372 1415
rect 664 1399 668 1415
rect 816 1359 820 1375
rect 1032 1359 1036 1375
rect 1320 1355 1324 1419
rect 1752 1355 1756 1371
rect 1840 1355 1844 1371
rect 1192 1315 1196 1331
rect 1256 1315 1260 1331
rect 1440 1315 1444 1331
rect 1536 1315 1540 1331
rect 288 1287 292 1303
rect 424 1287 428 1303
rect 816 1287 820 1303
rect 896 1287 900 1303
rect 976 1287 980 1303
rect 288 1243 292 1259
rect 352 1243 356 1259
rect 1208 1251 1212 1267
rect 1264 1251 1268 1267
rect 1424 1251 1428 1267
rect 1512 1251 1516 1267
rect 1688 1251 1692 1267
rect 1776 1251 1780 1267
rect 1864 1251 1868 1267
rect 2104 1227 2108 1267
rect 584 1175 588 1191
rect 640 1175 644 1191
rect 704 1175 708 1191
rect 776 1175 780 1191
rect 848 1175 852 1191
rect 1192 1143 1196 1159
rect 1240 1143 1244 1159
rect 1384 1143 1388 1159
rect 1456 1143 1460 1159
rect 1592 1143 1596 1159
rect 1664 1143 1668 1159
rect 1744 1143 1748 1159
rect 1832 1143 1836 1159
rect 1248 1099 1252 1139
rect 232 1067 236 1083
rect 288 1067 292 1083
rect 352 1067 356 1083
rect 432 1067 436 1083
rect 512 1067 516 1083
rect 672 1067 676 1083
rect 744 1067 748 1083
rect 816 1067 820 1083
rect 664 1023 668 1039
rect 776 1023 780 1039
rect 832 1023 836 1039
rect 1696 1035 1700 1051
rect 1792 1035 1796 1051
rect 1440 991 1444 1007
rect 1744 991 1748 1015
rect 208 955 212 971
rect 616 955 620 971
rect 664 955 668 971
rect 720 955 724 971
rect 776 955 780 971
rect 1648 919 1652 935
rect 1720 919 1724 935
rect 336 843 340 859
rect 800 843 804 859
rect 864 843 868 859
rect 976 843 980 859
rect 2056 835 2060 915
rect 376 803 380 819
rect 896 803 900 819
rect 960 803 964 819
rect 1576 815 1580 831
rect 1664 815 1668 831
rect 1888 815 1892 831
rect 2104 795 2108 831
rect 1656 775 1660 791
rect 248 739 252 755
rect 312 739 316 755
rect 384 739 388 755
rect 672 739 676 755
rect 1400 735 1404 771
rect 272 699 276 715
rect 504 699 508 715
rect 768 699 772 719
rect 1488 707 1492 723
rect 1536 707 1540 723
rect 1584 707 1588 723
rect 1688 707 1692 723
rect 1800 707 1804 723
rect 2056 707 2060 723
rect 248 635 252 651
rect 432 635 436 651
rect 560 635 564 651
rect 792 635 796 651
rect 1312 603 1316 619
rect 1376 603 1380 619
rect 1528 603 1532 619
rect 1616 603 1620 619
rect 1704 603 1708 619
rect 568 587 572 603
rect 1392 559 1396 575
rect 1552 559 1556 575
rect 544 519 548 535
rect 592 519 596 535
rect 640 519 644 535
rect 736 519 740 535
rect 2040 491 2044 555
rect 360 403 364 419
rect 640 403 644 419
rect 712 403 716 419
rect 776 403 780 419
rect 840 403 844 419
rect 904 403 908 419
rect 1232 387 1236 403
rect 1288 387 1292 403
rect 1368 387 1372 403
rect 1448 387 1452 403
rect 1784 387 1788 403
rect 248 355 252 371
rect 304 355 308 371
rect 2104 363 2108 403
rect 1760 343 1764 359
rect 1832 343 1836 359
rect 576 287 580 303
rect 624 287 628 303
rect 672 287 676 303
rect 816 287 820 303
rect 864 287 868 303
rect 1544 271 1548 287
rect 1592 271 1596 287
rect 1648 271 1652 287
rect 1768 271 1772 287
rect 1960 231 1964 247
rect 280 163 284 179
rect 328 163 332 179
rect 376 163 380 179
rect 432 163 436 179
rect 1264 163 1268 179
rect 1328 163 1332 179
rect 1392 163 1396 179
rect 1464 163 1468 179
rect 1624 163 1628 179
rect 1696 163 1700 179
rect 1768 163 1772 179
rect 1912 163 1916 179
<< m2c >>
rect 1368 2199 1372 2203
rect 1408 2199 1412 2203
rect 1448 2199 1452 2203
rect 1488 2199 1492 2203
rect 1528 2199 1532 2203
rect 1568 2199 1572 2203
rect 1608 2199 1612 2203
rect 1648 2199 1652 2203
rect 1688 2199 1692 2203
rect 1728 2199 1732 2203
rect 1768 2199 1772 2203
rect 1808 2199 1812 2203
rect 1848 2199 1852 2203
rect 1368 2179 1372 2183
rect 1408 2179 1412 2183
rect 1448 2179 1452 2183
rect 1488 2179 1492 2183
rect 1528 2179 1532 2183
rect 1568 2179 1572 2183
rect 1608 2179 1612 2183
rect 1648 2179 1652 2183
rect 1688 2179 1692 2183
rect 1728 2179 1732 2183
rect 1768 2179 1772 2183
rect 1808 2179 1812 2183
rect 1848 2179 1852 2183
rect 1312 2135 1316 2139
rect 1352 2135 1356 2139
rect 1392 2135 1396 2139
rect 1400 2135 1404 2139
rect 1440 2135 1444 2139
rect 1448 2135 1452 2139
rect 1488 2135 1492 2139
rect 1496 2135 1500 2139
rect 1544 2135 1548 2139
rect 1552 2135 1556 2139
rect 1600 2135 1604 2139
rect 1648 2135 1652 2139
rect 1656 2135 1660 2139
rect 1696 2135 1700 2139
rect 1744 2135 1748 2139
rect 1800 2135 1804 2139
rect 1856 2135 1860 2139
rect 1864 2135 1868 2139
rect 1912 2135 1916 2139
rect 1312 2115 1316 2119
rect 1352 2115 1356 2119
rect 1392 2115 1396 2119
rect 1400 2115 1404 2119
rect 1440 2115 1444 2119
rect 1448 2115 1452 2119
rect 1488 2115 1492 2119
rect 1496 2115 1500 2119
rect 1544 2115 1548 2119
rect 1552 2115 1556 2119
rect 1600 2115 1604 2119
rect 1648 2115 1652 2119
rect 1656 2115 1660 2119
rect 1696 2115 1700 2119
rect 1744 2115 1748 2119
rect 1800 2115 1804 2119
rect 1856 2115 1860 2119
rect 1864 2115 1868 2119
rect 1912 2115 1916 2119
rect 1248 2091 1252 2095
rect 1304 2091 1308 2095
rect 1368 2091 1372 2095
rect 1448 2091 1452 2095
rect 1528 2091 1532 2095
rect 1608 2091 1612 2095
rect 1688 2091 1692 2095
rect 1768 2091 1772 2095
rect 1856 2091 1860 2095
rect 1944 2091 1948 2095
rect 2032 2091 2036 2095
rect 1248 2071 1252 2075
rect 1304 2071 1308 2075
rect 1368 2071 1372 2075
rect 1448 2071 1452 2075
rect 1528 2071 1532 2075
rect 1608 2071 1612 2075
rect 1688 2071 1692 2075
rect 1768 2071 1772 2075
rect 1856 2071 1860 2075
rect 1944 2071 1948 2075
rect 2032 2071 2036 2075
rect 2096 2071 2100 2075
rect 1208 2027 1212 2031
rect 1264 2027 1268 2031
rect 1336 2027 1340 2031
rect 1424 2027 1428 2031
rect 1512 2027 1516 2031
rect 1608 2027 1612 2031
rect 1696 2027 1700 2031
rect 1704 2027 1708 2031
rect 1784 2027 1788 2031
rect 1864 2027 1868 2031
rect 1944 2027 1948 2031
rect 2032 2027 2036 2031
rect 2096 2027 2100 2031
rect 2104 2027 2108 2031
rect 216 2019 220 2023
rect 256 2019 260 2023
rect 312 2019 316 2023
rect 376 2019 380 2023
rect 448 2019 452 2023
rect 520 2019 524 2023
rect 600 2019 604 2023
rect 672 2019 676 2023
rect 744 2019 748 2023
rect 808 2019 812 2023
rect 864 2019 868 2023
rect 920 2019 924 2023
rect 976 2019 980 2023
rect 1032 2019 1036 2023
rect 1072 2019 1076 2023
rect 1208 2007 1212 2011
rect 1264 2007 1268 2011
rect 1336 2007 1340 2011
rect 1424 2007 1428 2011
rect 1512 2007 1516 2011
rect 1608 2007 1612 2011
rect 1696 2007 1700 2011
rect 1704 2007 1708 2011
rect 1784 2007 1788 2011
rect 1864 2007 1868 2011
rect 1944 2007 1948 2011
rect 2032 2007 2036 2011
rect 2096 2007 2100 2011
rect 216 1999 220 2003
rect 256 1999 260 2003
rect 312 1999 316 2003
rect 376 1999 380 2003
rect 448 1999 452 2003
rect 520 1999 524 2003
rect 600 1999 604 2003
rect 672 1999 676 2003
rect 712 1999 716 2003
rect 744 1999 748 2003
rect 808 1999 812 2003
rect 864 1999 868 2003
rect 920 1999 924 2003
rect 976 1999 980 2003
rect 1032 1999 1036 2003
rect 1072 1999 1076 2003
rect 1328 1987 1332 1991
rect 1408 1987 1412 1991
rect 1488 1987 1492 1991
rect 1568 1987 1572 1991
rect 1640 1987 1644 1991
rect 1712 1987 1716 1991
rect 1776 1987 1780 1991
rect 1840 1987 1844 1991
rect 1904 1987 1908 1991
rect 1976 1987 1980 1991
rect 2048 1987 2052 1991
rect 2096 1987 2100 1991
rect 2104 1987 2108 1991
rect 1328 1967 1332 1971
rect 1408 1967 1412 1971
rect 1488 1967 1492 1971
rect 1568 1967 1572 1971
rect 1640 1967 1644 1971
rect 1712 1967 1716 1971
rect 1776 1967 1780 1971
rect 1840 1967 1844 1971
rect 1904 1967 1908 1971
rect 1976 1967 1980 1971
rect 2048 1967 2052 1971
rect 2096 1967 2100 1971
rect 712 1963 716 1967
rect 216 1955 220 1959
rect 272 1955 276 1959
rect 336 1955 340 1959
rect 400 1955 404 1959
rect 472 1955 476 1959
rect 544 1955 548 1959
rect 616 1955 620 1959
rect 624 1955 628 1959
rect 680 1955 684 1959
rect 688 1955 692 1959
rect 744 1955 748 1959
rect 752 1955 756 1959
rect 800 1955 804 1959
rect 808 1955 812 1959
rect 848 1955 852 1959
rect 896 1955 900 1959
rect 944 1955 948 1959
rect 952 1955 956 1959
rect 992 1955 996 1959
rect 1032 1955 1036 1959
rect 1072 1955 1076 1959
rect 216 1935 220 1939
rect 272 1935 276 1939
rect 336 1935 340 1939
rect 400 1935 404 1939
rect 472 1935 476 1939
rect 544 1935 548 1939
rect 616 1935 620 1939
rect 624 1935 628 1939
rect 680 1935 684 1939
rect 688 1935 692 1939
rect 744 1935 748 1939
rect 752 1935 756 1939
rect 800 1935 804 1939
rect 808 1935 812 1939
rect 848 1935 852 1939
rect 896 1935 900 1939
rect 944 1935 948 1939
rect 952 1935 956 1939
rect 992 1935 996 1939
rect 1032 1935 1036 1939
rect 1072 1935 1076 1939
rect 1184 1919 1188 1923
rect 1192 1919 1196 1923
rect 1248 1919 1252 1923
rect 1328 1919 1332 1923
rect 1408 1919 1412 1923
rect 1488 1919 1492 1923
rect 1560 1919 1564 1923
rect 1568 1919 1572 1923
rect 1640 1919 1644 1923
rect 1648 1919 1652 1923
rect 1720 1919 1724 1923
rect 1808 1919 1812 1923
rect 1816 1919 1820 1923
rect 1904 1919 1908 1923
rect 1912 1919 1916 1923
rect 2008 1919 2012 1923
rect 2096 1919 2100 1923
rect 160 1915 164 1919
rect 200 1915 204 1919
rect 256 1915 260 1919
rect 320 1915 324 1919
rect 392 1915 396 1919
rect 456 1915 460 1919
rect 520 1915 524 1919
rect 584 1915 588 1919
rect 640 1915 644 1919
rect 696 1915 700 1919
rect 752 1915 756 1919
rect 808 1915 812 1919
rect 872 1915 876 1919
rect 1184 1899 1188 1903
rect 1192 1899 1196 1903
rect 1248 1899 1252 1903
rect 1328 1899 1332 1903
rect 1408 1899 1412 1903
rect 1488 1899 1492 1903
rect 1560 1899 1564 1903
rect 1568 1899 1572 1903
rect 1640 1899 1644 1903
rect 1648 1899 1652 1903
rect 1720 1899 1724 1903
rect 1808 1899 1812 1903
rect 1816 1899 1820 1903
rect 1904 1899 1908 1903
rect 1912 1899 1916 1903
rect 2008 1899 2012 1903
rect 2096 1899 2100 1903
rect 160 1895 164 1899
rect 200 1895 204 1899
rect 256 1895 260 1899
rect 320 1895 324 1899
rect 392 1895 396 1899
rect 456 1895 460 1899
rect 520 1895 524 1899
rect 584 1895 588 1899
rect 640 1895 644 1899
rect 696 1895 700 1899
rect 752 1895 756 1899
rect 808 1895 812 1899
rect 872 1895 876 1899
rect 1536 1883 1540 1887
rect 1184 1875 1188 1879
rect 1224 1875 1228 1879
rect 1288 1875 1292 1879
rect 1352 1875 1356 1879
rect 1416 1875 1420 1879
rect 1472 1875 1476 1879
rect 1528 1875 1532 1879
rect 1584 1875 1588 1879
rect 1656 1875 1660 1879
rect 1736 1875 1740 1879
rect 1824 1875 1828 1879
rect 1920 1875 1924 1879
rect 2016 1875 2020 1879
rect 2096 1875 2100 1879
rect 1184 1855 1188 1859
rect 1224 1855 1228 1859
rect 1288 1855 1292 1859
rect 1352 1855 1356 1859
rect 1416 1855 1420 1859
rect 1472 1855 1476 1859
rect 1528 1855 1532 1859
rect 1536 1855 1540 1859
rect 1584 1855 1588 1859
rect 1656 1855 1660 1859
rect 1736 1855 1740 1859
rect 1824 1855 1828 1859
rect 1920 1855 1924 1859
rect 2016 1855 2020 1859
rect 2096 1855 2100 1859
rect 160 1847 164 1851
rect 224 1847 228 1851
rect 296 1847 300 1851
rect 360 1847 364 1851
rect 368 1847 372 1851
rect 424 1847 428 1851
rect 480 1847 484 1851
rect 528 1847 532 1851
rect 536 1847 540 1851
rect 576 1847 580 1851
rect 584 1847 588 1851
rect 624 1847 628 1851
rect 632 1847 636 1851
rect 672 1847 676 1851
rect 680 1847 684 1851
rect 720 1847 724 1851
rect 728 1847 732 1851
rect 776 1847 780 1851
rect 160 1827 164 1831
rect 224 1827 228 1831
rect 296 1827 300 1831
rect 360 1827 364 1831
rect 368 1827 372 1831
rect 424 1827 428 1831
rect 480 1827 484 1831
rect 528 1827 532 1831
rect 536 1827 540 1831
rect 576 1827 580 1831
rect 584 1827 588 1831
rect 624 1827 628 1831
rect 632 1827 636 1831
rect 672 1827 676 1831
rect 680 1827 684 1831
rect 720 1827 724 1831
rect 728 1827 732 1831
rect 776 1827 780 1831
rect 1184 1811 1188 1815
rect 1256 1811 1260 1815
rect 1328 1811 1332 1815
rect 1408 1811 1412 1815
rect 1488 1811 1492 1815
rect 1576 1811 1580 1815
rect 1672 1811 1676 1815
rect 1680 1811 1684 1815
rect 1776 1811 1780 1815
rect 1880 1811 1884 1815
rect 1992 1811 1996 1815
rect 2096 1811 2100 1815
rect 176 1799 180 1803
rect 240 1799 244 1803
rect 248 1799 252 1803
rect 296 1799 300 1803
rect 352 1799 356 1803
rect 408 1799 412 1803
rect 416 1799 420 1803
rect 456 1799 460 1803
rect 504 1799 508 1803
rect 552 1799 556 1803
rect 600 1799 604 1803
rect 648 1799 652 1803
rect 696 1799 700 1803
rect 752 1799 756 1803
rect 1184 1791 1188 1795
rect 1256 1791 1260 1795
rect 1328 1791 1332 1795
rect 1408 1791 1412 1795
rect 1488 1791 1492 1795
rect 1576 1791 1580 1795
rect 1672 1791 1676 1795
rect 1680 1791 1684 1795
rect 1776 1791 1780 1795
rect 1880 1791 1884 1795
rect 1992 1791 1996 1795
rect 2096 1791 2100 1795
rect 176 1779 180 1783
rect 240 1779 244 1783
rect 248 1779 252 1783
rect 296 1779 300 1783
rect 352 1779 356 1783
rect 408 1779 412 1783
rect 416 1779 420 1783
rect 456 1779 460 1783
rect 504 1779 508 1783
rect 552 1779 556 1783
rect 600 1779 604 1783
rect 648 1779 652 1783
rect 696 1779 700 1783
rect 752 1779 756 1783
rect 1216 1771 1220 1775
rect 1280 1771 1284 1775
rect 1344 1771 1348 1775
rect 1408 1771 1412 1775
rect 1480 1771 1484 1775
rect 1552 1773 1556 1777
rect 1632 1771 1636 1775
rect 1712 1771 1716 1775
rect 1792 1771 1796 1775
rect 1872 1771 1876 1775
rect 1952 1771 1956 1775
rect 2032 1771 2036 1775
rect 2096 1771 2100 1775
rect 1216 1751 1220 1755
rect 1280 1751 1284 1755
rect 1344 1751 1348 1755
rect 1408 1751 1412 1755
rect 1480 1751 1484 1755
rect 1552 1751 1556 1755
rect 1632 1751 1636 1755
rect 1712 1751 1716 1755
rect 1792 1751 1796 1755
rect 1872 1751 1876 1755
rect 1952 1751 1956 1755
rect 2032 1751 2036 1755
rect 2096 1751 2100 1755
rect 256 1735 260 1739
rect 320 1735 324 1739
rect 376 1735 380 1739
rect 384 1735 388 1739
rect 440 1735 444 1739
rect 504 1735 508 1739
rect 512 1735 516 1739
rect 568 1735 572 1739
rect 640 1735 644 1739
rect 712 1735 716 1739
rect 720 1735 724 1739
rect 784 1735 788 1739
rect 856 1735 860 1739
rect 936 1735 940 1739
rect 1016 1735 1020 1739
rect 256 1715 260 1719
rect 320 1715 324 1719
rect 376 1715 380 1719
rect 384 1715 388 1719
rect 440 1715 444 1719
rect 504 1715 508 1719
rect 512 1715 516 1719
rect 568 1715 572 1719
rect 640 1715 644 1719
rect 712 1715 716 1719
rect 720 1715 724 1719
rect 784 1715 788 1719
rect 856 1715 860 1719
rect 936 1715 940 1719
rect 1016 1715 1020 1719
rect 1272 1707 1276 1711
rect 1320 1707 1324 1711
rect 1368 1707 1372 1711
rect 1424 1707 1428 1711
rect 1488 1707 1492 1711
rect 1552 1707 1556 1711
rect 1624 1707 1628 1711
rect 1696 1707 1700 1711
rect 1768 1707 1772 1711
rect 1832 1707 1836 1711
rect 1904 1707 1908 1711
rect 1976 1707 1980 1711
rect 2048 1707 2052 1711
rect 2056 1707 2060 1711
rect 2096 1707 2100 1711
rect 160 1691 164 1695
rect 224 1691 228 1695
rect 304 1691 308 1695
rect 392 1691 396 1695
rect 400 1691 404 1695
rect 488 1691 492 1695
rect 496 1691 500 1695
rect 576 1691 580 1695
rect 664 1691 668 1695
rect 744 1691 748 1695
rect 816 1691 820 1695
rect 880 1691 884 1695
rect 944 1691 948 1695
rect 1008 1691 1012 1695
rect 1072 1691 1076 1695
rect 1272 1687 1276 1691
rect 1320 1687 1324 1691
rect 1368 1687 1372 1691
rect 1424 1687 1428 1691
rect 1488 1687 1492 1691
rect 1552 1687 1556 1691
rect 1624 1687 1628 1691
rect 1696 1687 1700 1691
rect 1768 1689 1772 1693
rect 1832 1687 1836 1691
rect 1904 1687 1908 1691
rect 1976 1687 1980 1691
rect 2048 1687 2052 1691
rect 2056 1687 2060 1691
rect 2096 1687 2100 1691
rect 160 1671 164 1675
rect 224 1671 228 1675
rect 304 1671 308 1675
rect 392 1671 396 1675
rect 400 1671 404 1675
rect 488 1671 492 1675
rect 496 1671 500 1675
rect 576 1671 580 1675
rect 664 1671 668 1675
rect 744 1671 748 1675
rect 816 1671 820 1675
rect 880 1671 884 1675
rect 944 1671 948 1675
rect 1008 1671 1012 1675
rect 1072 1671 1076 1675
rect 1288 1663 1292 1667
rect 1328 1663 1332 1667
rect 1368 1663 1372 1667
rect 1416 1663 1420 1667
rect 1472 1663 1476 1667
rect 1528 1665 1532 1669
rect 1592 1663 1596 1667
rect 1656 1663 1660 1667
rect 1720 1663 1724 1667
rect 1784 1663 1788 1667
rect 1856 1663 1860 1667
rect 1936 1663 1940 1667
rect 2024 1663 2028 1667
rect 2096 1663 2100 1667
rect 1288 1643 1292 1647
rect 1328 1643 1332 1647
rect 1368 1643 1372 1647
rect 1416 1643 1420 1647
rect 1472 1643 1476 1647
rect 1528 1643 1532 1647
rect 1592 1643 1596 1647
rect 1656 1643 1660 1647
rect 1720 1643 1724 1647
rect 1784 1643 1788 1647
rect 1856 1643 1860 1647
rect 1936 1643 1940 1647
rect 2024 1643 2028 1647
rect 2096 1643 2100 1647
rect 160 1623 164 1627
rect 208 1623 212 1627
rect 288 1623 292 1627
rect 296 1623 300 1627
rect 368 1623 372 1627
rect 376 1623 380 1627
rect 448 1623 452 1627
rect 456 1623 460 1627
rect 528 1623 532 1627
rect 608 1623 612 1627
rect 680 1623 684 1627
rect 752 1623 756 1627
rect 816 1623 820 1627
rect 872 1623 876 1627
rect 928 1623 932 1627
rect 984 1623 988 1627
rect 992 1623 996 1627
rect 1032 1623 1036 1627
rect 1072 1623 1076 1627
rect 160 1603 164 1607
rect 208 1603 212 1607
rect 288 1603 292 1607
rect 296 1603 300 1607
rect 368 1603 372 1607
rect 376 1603 380 1607
rect 448 1603 452 1607
rect 456 1603 460 1607
rect 528 1603 532 1607
rect 608 1603 612 1607
rect 680 1603 684 1607
rect 752 1603 756 1607
rect 816 1603 820 1607
rect 872 1603 876 1607
rect 928 1603 932 1607
rect 984 1603 988 1607
rect 992 1603 996 1607
rect 1032 1603 1036 1607
rect 1072 1603 1076 1607
rect 1184 1587 1188 1591
rect 1240 1587 1244 1591
rect 1328 1587 1332 1591
rect 1408 1587 1412 1591
rect 1488 1587 1492 1591
rect 1496 1587 1500 1591
rect 1568 1587 1572 1591
rect 1648 1587 1652 1591
rect 1736 1587 1740 1591
rect 1824 1587 1828 1591
rect 1832 1587 1836 1591
rect 1912 1587 1916 1591
rect 2008 1587 2012 1591
rect 2096 1587 2100 1591
rect 2104 1587 2108 1591
rect 160 1583 164 1587
rect 200 1583 204 1587
rect 208 1583 212 1587
rect 256 1583 260 1587
rect 288 1583 292 1587
rect 328 1583 332 1587
rect 336 1583 340 1587
rect 400 1583 404 1587
rect 408 1583 412 1587
rect 480 1583 484 1587
rect 552 1583 556 1587
rect 624 1583 628 1587
rect 632 1583 636 1587
rect 696 1583 700 1587
rect 768 1583 772 1587
rect 840 1583 844 1587
rect 912 1583 916 1587
rect 160 1563 164 1567
rect 200 1563 204 1567
rect 208 1563 212 1567
rect 216 1563 220 1567
rect 256 1563 260 1567
rect 160 1519 164 1523
rect 200 1519 204 1523
rect 1184 1567 1188 1571
rect 1240 1567 1244 1571
rect 1328 1567 1332 1571
rect 1408 1567 1412 1571
rect 1488 1567 1492 1571
rect 1496 1567 1500 1571
rect 1568 1567 1572 1571
rect 1648 1567 1652 1571
rect 1736 1567 1740 1571
rect 1824 1567 1828 1571
rect 1832 1567 1836 1571
rect 1912 1567 1916 1571
rect 2008 1567 2012 1571
rect 2096 1567 2100 1571
rect 328 1563 332 1567
rect 336 1563 340 1567
rect 400 1563 404 1567
rect 408 1563 412 1567
rect 480 1563 484 1567
rect 552 1563 556 1567
rect 624 1563 628 1567
rect 632 1563 636 1567
rect 696 1563 700 1567
rect 768 1563 772 1567
rect 840 1563 844 1567
rect 912 1563 916 1567
rect 1184 1547 1188 1551
rect 1224 1547 1228 1551
rect 1272 1547 1276 1551
rect 1344 1547 1348 1551
rect 1424 1547 1428 1551
rect 1504 1547 1508 1551
rect 1584 1547 1588 1551
rect 1672 1547 1676 1551
rect 1760 1547 1764 1551
rect 1848 1547 1852 1551
rect 1856 1547 1860 1551
rect 1936 1547 1940 1551
rect 1944 1547 1948 1551
rect 2024 1547 2028 1551
rect 2096 1547 2100 1551
rect 2104 1547 2108 1551
rect 288 1527 292 1531
rect 1184 1527 1188 1531
rect 1224 1527 1228 1531
rect 1272 1527 1276 1531
rect 1344 1527 1348 1531
rect 1424 1527 1428 1531
rect 1504 1527 1508 1531
rect 1584 1527 1588 1531
rect 1672 1527 1676 1531
rect 1760 1527 1764 1531
rect 1848 1527 1852 1531
rect 1856 1527 1860 1531
rect 1936 1527 1940 1531
rect 1944 1527 1948 1531
rect 2024 1527 2028 1531
rect 2096 1527 2100 1531
rect 256 1519 260 1523
rect 264 1519 268 1523
rect 336 1519 340 1523
rect 344 1519 348 1523
rect 416 1519 420 1523
rect 424 1519 428 1523
rect 504 1519 508 1523
rect 592 1519 596 1523
rect 600 1519 604 1523
rect 680 1519 684 1523
rect 688 1519 692 1523
rect 768 1519 772 1523
rect 848 1519 852 1523
rect 936 1519 940 1523
rect 1024 1519 1028 1523
rect 160 1499 164 1503
rect 200 1499 204 1503
rect 216 1499 220 1503
rect 256 1499 260 1503
rect 264 1499 268 1503
rect 336 1499 340 1503
rect 344 1499 348 1503
rect 416 1499 420 1503
rect 424 1499 428 1503
rect 504 1499 508 1503
rect 592 1499 596 1503
rect 600 1499 604 1503
rect 680 1499 684 1503
rect 688 1499 692 1503
rect 768 1499 772 1503
rect 848 1499 852 1503
rect 936 1499 940 1503
rect 1024 1499 1028 1503
rect 1184 1483 1188 1487
rect 1224 1483 1228 1487
rect 1264 1483 1268 1487
rect 1328 1483 1332 1487
rect 1400 1483 1404 1487
rect 1480 1483 1484 1487
rect 1520 1483 1524 1487
rect 1568 1483 1572 1487
rect 1648 1483 1652 1487
rect 1656 1483 1660 1487
rect 1728 1483 1732 1487
rect 1736 1483 1740 1487
rect 1800 1483 1804 1487
rect 1808 1483 1812 1487
rect 1872 1483 1876 1487
rect 1944 1483 1948 1487
rect 2016 1483 2020 1487
rect 2088 1483 2092 1487
rect 160 1479 164 1483
rect 224 1479 228 1483
rect 304 1479 308 1483
rect 312 1479 316 1483
rect 384 1479 388 1483
rect 464 1479 468 1483
rect 544 1479 548 1483
rect 624 1479 628 1483
rect 704 1479 708 1483
rect 792 1479 796 1483
rect 880 1479 884 1483
rect 968 1479 972 1483
rect 1056 1479 1060 1483
rect 1184 1463 1188 1467
rect 1224 1463 1228 1467
rect 1264 1463 1268 1467
rect 1328 1463 1332 1467
rect 1400 1463 1404 1467
rect 1480 1463 1484 1467
rect 1520 1463 1524 1467
rect 1568 1463 1572 1467
rect 1648 1463 1652 1467
rect 1656 1463 1660 1467
rect 1728 1463 1732 1467
rect 1736 1463 1740 1467
rect 1800 1463 1804 1467
rect 1808 1463 1812 1467
rect 1872 1463 1876 1467
rect 1944 1463 1948 1467
rect 2016 1463 2020 1467
rect 2088 1463 2092 1467
rect 160 1459 164 1463
rect 224 1459 228 1463
rect 304 1459 308 1463
rect 312 1459 316 1463
rect 384 1459 388 1463
rect 464 1459 468 1463
rect 544 1459 548 1463
rect 624 1459 628 1463
rect 704 1459 708 1463
rect 792 1459 796 1463
rect 880 1459 884 1463
rect 968 1459 972 1463
rect 1056 1459 1060 1463
rect 1304 1439 1308 1443
rect 1352 1439 1356 1443
rect 1408 1439 1412 1443
rect 1464 1439 1468 1443
rect 1520 1439 1524 1443
rect 1576 1439 1580 1443
rect 1632 1439 1636 1443
rect 1696 1439 1700 1443
rect 1760 1439 1764 1443
rect 1768 1439 1772 1443
rect 1832 1439 1836 1443
rect 1840 1439 1844 1443
rect 1912 1439 1916 1443
rect 2000 1439 2004 1443
rect 2088 1439 2092 1443
rect 1304 1419 1308 1423
rect 1320 1419 1324 1423
rect 1352 1419 1356 1423
rect 1408 1419 1412 1423
rect 1464 1419 1468 1423
rect 1520 1419 1524 1423
rect 1576 1419 1580 1423
rect 1632 1419 1636 1423
rect 1696 1419 1700 1423
rect 1760 1419 1764 1423
rect 1768 1419 1772 1423
rect 1832 1419 1836 1423
rect 1840 1419 1844 1423
rect 1912 1419 1916 1423
rect 2000 1419 2004 1423
rect 2088 1419 2092 1423
rect 160 1415 164 1419
rect 216 1415 220 1419
rect 288 1415 292 1419
rect 360 1415 364 1419
rect 368 1415 372 1419
rect 432 1415 436 1419
rect 504 1415 508 1419
rect 576 1415 580 1419
rect 656 1415 660 1419
rect 664 1415 668 1419
rect 736 1415 740 1419
rect 824 1415 828 1419
rect 912 1415 916 1419
rect 1000 1415 1004 1419
rect 1072 1415 1076 1419
rect 160 1395 164 1399
rect 216 1395 220 1399
rect 288 1395 292 1399
rect 360 1395 364 1399
rect 368 1395 372 1399
rect 432 1395 436 1399
rect 504 1395 508 1399
rect 576 1395 580 1399
rect 656 1395 660 1399
rect 664 1395 668 1399
rect 736 1395 740 1399
rect 824 1395 828 1399
rect 912 1395 916 1399
rect 1000 1395 1004 1399
rect 1072 1395 1076 1399
rect 160 1375 164 1379
rect 200 1375 204 1379
rect 264 1375 268 1379
rect 328 1375 332 1379
rect 392 1375 396 1379
rect 464 1375 468 1379
rect 528 1375 532 1379
rect 600 1375 604 1379
rect 672 1375 676 1379
rect 736 1375 740 1379
rect 808 1375 812 1379
rect 816 1375 820 1379
rect 880 1375 884 1379
rect 952 1375 956 1379
rect 1024 1375 1028 1379
rect 1032 1375 1036 1379
rect 1072 1375 1076 1379
rect 160 1355 164 1359
rect 200 1355 204 1359
rect 264 1355 268 1359
rect 328 1355 332 1359
rect 392 1355 396 1359
rect 464 1355 468 1359
rect 528 1355 532 1359
rect 600 1355 604 1359
rect 672 1355 676 1359
rect 736 1355 740 1359
rect 808 1355 812 1359
rect 816 1355 820 1359
rect 880 1355 884 1359
rect 952 1355 956 1359
rect 1024 1355 1028 1359
rect 1032 1355 1036 1359
rect 1072 1355 1076 1359
rect 1360 1371 1364 1375
rect 1400 1371 1404 1375
rect 1440 1371 1444 1375
rect 1480 1371 1484 1375
rect 1520 1371 1524 1375
rect 1560 1371 1564 1375
rect 1608 1371 1612 1375
rect 1672 1371 1676 1375
rect 1744 1371 1748 1375
rect 1752 1371 1756 1375
rect 1832 1371 1836 1375
rect 1840 1371 1844 1375
rect 1920 1371 1924 1375
rect 2016 1371 2020 1375
rect 2096 1371 2100 1375
rect 1320 1351 1324 1355
rect 1360 1351 1364 1355
rect 1400 1351 1404 1355
rect 1440 1351 1444 1355
rect 1480 1351 1484 1355
rect 1520 1351 1524 1355
rect 1560 1351 1564 1355
rect 1608 1351 1612 1355
rect 1672 1351 1676 1355
rect 1744 1351 1748 1355
rect 1752 1351 1756 1355
rect 1832 1351 1836 1355
rect 1840 1351 1844 1355
rect 1920 1351 1924 1355
rect 2016 1351 2020 1355
rect 2096 1351 2100 1355
rect 1184 1331 1188 1335
rect 1192 1331 1196 1335
rect 1248 1331 1252 1335
rect 1256 1331 1260 1335
rect 1336 1331 1340 1335
rect 1432 1331 1436 1335
rect 1440 1331 1444 1335
rect 1528 1331 1532 1335
rect 1536 1331 1540 1335
rect 1624 1331 1628 1335
rect 1704 1331 1708 1335
rect 1784 1331 1788 1335
rect 1856 1331 1860 1335
rect 1920 1331 1924 1335
rect 1984 1331 1988 1335
rect 2048 1331 2052 1335
rect 2096 1331 2100 1335
rect 1184 1311 1188 1315
rect 1192 1311 1196 1315
rect 1248 1311 1252 1315
rect 1256 1311 1260 1315
rect 1336 1311 1340 1315
rect 1432 1311 1436 1315
rect 1440 1311 1444 1315
rect 1528 1311 1532 1315
rect 1536 1311 1540 1315
rect 1624 1311 1628 1315
rect 1704 1311 1708 1315
rect 1784 1311 1788 1315
rect 1856 1311 1860 1315
rect 1920 1311 1924 1315
rect 1984 1311 1988 1315
rect 2048 1311 2052 1315
rect 2096 1311 2100 1315
rect 160 1303 164 1307
rect 200 1303 204 1307
rect 240 1303 244 1307
rect 280 1303 284 1307
rect 288 1303 292 1307
rect 344 1303 348 1307
rect 416 1303 420 1307
rect 424 1303 428 1307
rect 488 1303 492 1307
rect 568 1303 572 1307
rect 648 1303 652 1307
rect 728 1303 732 1307
rect 808 1303 812 1307
rect 816 1303 820 1307
rect 888 1303 892 1307
rect 896 1303 900 1307
rect 968 1303 972 1307
rect 976 1303 980 1307
rect 1048 1303 1052 1307
rect 160 1283 164 1287
rect 200 1283 204 1287
rect 240 1283 244 1287
rect 280 1283 284 1287
rect 288 1283 292 1287
rect 344 1283 348 1287
rect 416 1283 420 1287
rect 424 1283 428 1287
rect 488 1283 492 1287
rect 568 1283 572 1287
rect 648 1283 652 1287
rect 728 1283 732 1287
rect 808 1283 812 1287
rect 816 1283 820 1287
rect 888 1283 892 1287
rect 896 1283 900 1287
rect 968 1283 972 1287
rect 976 1283 980 1287
rect 1048 1283 1052 1287
rect 1200 1267 1204 1271
rect 1208 1267 1212 1271
rect 1256 1267 1260 1271
rect 1264 1267 1268 1271
rect 1328 1267 1332 1271
rect 1416 1267 1420 1271
rect 1424 1267 1428 1271
rect 1504 1267 1508 1271
rect 1512 1267 1516 1271
rect 1592 1267 1596 1271
rect 1680 1267 1684 1271
rect 1688 1267 1692 1271
rect 1768 1267 1772 1271
rect 1776 1267 1780 1271
rect 1856 1267 1860 1271
rect 1864 1267 1868 1271
rect 1944 1267 1948 1271
rect 2032 1267 2036 1271
rect 2096 1267 2100 1271
rect 2104 1267 2108 1271
rect 160 1259 164 1263
rect 200 1259 204 1263
rect 240 1259 244 1263
rect 280 1259 284 1263
rect 288 1259 292 1263
rect 344 1259 348 1263
rect 352 1259 356 1263
rect 424 1259 428 1263
rect 512 1259 516 1263
rect 608 1259 612 1263
rect 712 1259 716 1263
rect 824 1259 828 1263
rect 944 1259 948 1263
rect 1072 1259 1076 1263
rect 1200 1247 1204 1251
rect 1208 1247 1212 1251
rect 1256 1247 1260 1251
rect 1264 1247 1268 1251
rect 1328 1247 1332 1251
rect 1416 1247 1420 1251
rect 1424 1247 1428 1251
rect 1504 1247 1508 1251
rect 1512 1247 1516 1251
rect 1592 1247 1596 1251
rect 1680 1247 1684 1251
rect 1688 1247 1692 1251
rect 1768 1247 1772 1251
rect 1776 1247 1780 1251
rect 1856 1247 1860 1251
rect 1864 1247 1868 1251
rect 1944 1247 1948 1251
rect 2032 1247 2036 1251
rect 2096 1247 2100 1251
rect 160 1239 164 1243
rect 200 1239 204 1243
rect 240 1239 244 1243
rect 280 1239 284 1243
rect 288 1239 292 1243
rect 344 1239 348 1243
rect 352 1239 356 1243
rect 424 1239 428 1243
rect 512 1239 516 1243
rect 608 1239 612 1243
rect 712 1239 716 1243
rect 824 1239 828 1243
rect 944 1239 948 1243
rect 1072 1239 1076 1243
rect 1312 1223 1316 1227
rect 1352 1223 1356 1227
rect 1400 1223 1404 1227
rect 1456 1223 1460 1227
rect 1520 1223 1524 1227
rect 1584 1223 1588 1227
rect 1648 1223 1652 1227
rect 1704 1223 1708 1227
rect 1760 1223 1764 1227
rect 1816 1223 1820 1227
rect 1872 1223 1876 1227
rect 1928 1223 1932 1227
rect 1992 1223 1996 1227
rect 2056 1223 2060 1227
rect 2096 1223 2100 1227
rect 2104 1223 2108 1227
rect 1312 1203 1316 1207
rect 1352 1203 1356 1207
rect 1400 1203 1404 1207
rect 1456 1203 1460 1207
rect 1520 1203 1524 1207
rect 1584 1203 1588 1207
rect 1648 1203 1652 1207
rect 1704 1203 1708 1207
rect 1760 1203 1764 1207
rect 1816 1203 1820 1207
rect 1872 1203 1876 1207
rect 1928 1203 1932 1207
rect 1992 1203 1996 1207
rect 2056 1203 2060 1207
rect 2096 1203 2100 1207
rect 296 1191 300 1195
rect 336 1191 340 1195
rect 376 1191 380 1195
rect 424 1191 428 1195
rect 472 1191 476 1195
rect 520 1191 524 1195
rect 576 1191 580 1195
rect 584 1191 588 1195
rect 632 1191 636 1195
rect 640 1191 644 1195
rect 696 1191 700 1195
rect 704 1191 708 1195
rect 768 1191 772 1195
rect 776 1191 780 1195
rect 840 1191 844 1195
rect 848 1191 852 1195
rect 920 1191 924 1195
rect 1008 1191 1012 1195
rect 296 1171 300 1175
rect 336 1171 340 1175
rect 376 1171 380 1175
rect 424 1171 428 1175
rect 472 1171 476 1175
rect 520 1171 524 1175
rect 576 1171 580 1175
rect 584 1171 588 1175
rect 632 1171 636 1175
rect 640 1171 644 1175
rect 696 1171 700 1175
rect 704 1171 708 1175
rect 768 1171 772 1175
rect 776 1171 780 1175
rect 840 1171 844 1175
rect 848 1171 852 1175
rect 920 1171 924 1175
rect 1008 1171 1012 1175
rect 1184 1159 1188 1163
rect 1192 1159 1196 1163
rect 1232 1159 1236 1163
rect 1240 1159 1244 1163
rect 1304 1159 1308 1163
rect 1376 1159 1380 1163
rect 1384 1159 1388 1163
rect 1448 1159 1452 1163
rect 1456 1159 1460 1163
rect 1512 1159 1516 1163
rect 1584 1159 1588 1163
rect 1592 1159 1596 1163
rect 1656 1159 1660 1163
rect 1664 1159 1668 1163
rect 1736 1159 1740 1163
rect 1744 1159 1748 1163
rect 1824 1159 1828 1163
rect 1832 1159 1836 1163
rect 1912 1159 1916 1163
rect 2008 1159 2012 1163
rect 2096 1159 2100 1163
rect 424 1147 428 1151
rect 464 1147 468 1151
rect 504 1147 508 1151
rect 552 1147 556 1151
rect 600 1147 604 1151
rect 648 1147 652 1151
rect 696 1147 700 1151
rect 744 1147 748 1151
rect 800 1147 804 1151
rect 856 1147 860 1151
rect 912 1147 916 1151
rect 968 1147 972 1151
rect 1032 1147 1036 1151
rect 1072 1147 1076 1151
rect 1184 1139 1188 1143
rect 1192 1139 1196 1143
rect 1232 1139 1236 1143
rect 1240 1139 1244 1143
rect 1248 1139 1252 1143
rect 1304 1139 1308 1143
rect 1376 1139 1380 1143
rect 1384 1139 1388 1143
rect 1448 1139 1452 1143
rect 1456 1139 1460 1143
rect 1512 1139 1516 1143
rect 1584 1139 1588 1143
rect 1592 1139 1596 1143
rect 1656 1139 1660 1143
rect 1664 1139 1668 1143
rect 1736 1139 1740 1143
rect 1744 1139 1748 1143
rect 1824 1139 1828 1143
rect 1832 1139 1836 1143
rect 1912 1139 1916 1143
rect 2008 1139 2012 1143
rect 2096 1139 2100 1143
rect 424 1127 428 1131
rect 464 1127 468 1131
rect 504 1127 508 1131
rect 552 1127 556 1131
rect 600 1127 604 1131
rect 648 1127 652 1131
rect 696 1127 700 1131
rect 744 1127 748 1131
rect 800 1127 804 1131
rect 856 1127 860 1131
rect 912 1127 916 1131
rect 968 1127 972 1131
rect 1032 1127 1036 1131
rect 1072 1127 1076 1131
rect 1216 1115 1220 1119
rect 1296 1115 1300 1119
rect 1368 1115 1372 1119
rect 1440 1115 1444 1119
rect 1512 1115 1516 1119
rect 1592 1115 1596 1119
rect 1680 1115 1684 1119
rect 1776 1115 1780 1119
rect 1880 1115 1884 1119
rect 1984 1115 1988 1119
rect 2096 1115 2100 1119
rect 1216 1095 1220 1099
rect 1248 1095 1252 1099
rect 1296 1095 1300 1099
rect 1368 1095 1372 1099
rect 1440 1095 1444 1099
rect 1512 1095 1516 1099
rect 1592 1095 1596 1099
rect 1680 1095 1684 1099
rect 1776 1095 1780 1099
rect 1880 1095 1884 1099
rect 1984 1097 1988 1101
rect 2096 1095 2100 1099
rect 184 1083 188 1087
rect 224 1083 228 1087
rect 232 1083 236 1087
rect 280 1083 284 1087
rect 288 1083 292 1087
rect 344 1083 348 1087
rect 352 1083 356 1087
rect 424 1083 428 1087
rect 432 1083 436 1087
rect 504 1083 508 1087
rect 512 1083 516 1087
rect 584 1083 588 1087
rect 664 1083 668 1087
rect 672 1083 676 1087
rect 736 1083 740 1087
rect 744 1083 748 1087
rect 808 1083 812 1087
rect 816 1083 820 1087
rect 880 1083 884 1087
rect 952 1083 956 1087
rect 1024 1083 1028 1087
rect 1072 1083 1076 1087
rect 184 1063 188 1067
rect 224 1063 228 1067
rect 232 1063 236 1067
rect 280 1063 284 1067
rect 288 1063 292 1067
rect 344 1063 348 1067
rect 352 1063 356 1067
rect 424 1063 428 1067
rect 432 1063 436 1067
rect 504 1063 508 1067
rect 512 1063 516 1067
rect 584 1063 588 1067
rect 664 1063 668 1067
rect 672 1063 676 1067
rect 736 1063 740 1067
rect 744 1063 748 1067
rect 808 1063 812 1067
rect 816 1063 820 1067
rect 880 1063 884 1067
rect 952 1063 956 1067
rect 1024 1063 1028 1067
rect 1072 1063 1076 1067
rect 1184 1051 1188 1055
rect 1224 1051 1228 1055
rect 1272 1051 1276 1055
rect 1328 1051 1332 1055
rect 1376 1051 1380 1055
rect 1424 1051 1428 1055
rect 1480 1051 1484 1055
rect 1536 1051 1540 1055
rect 1608 1051 1612 1055
rect 1688 1051 1692 1055
rect 1696 1051 1700 1055
rect 1784 1051 1788 1055
rect 1792 1051 1796 1055
rect 1888 1051 1892 1055
rect 1992 1051 1996 1055
rect 2096 1051 2100 1055
rect 160 1039 164 1043
rect 200 1039 204 1043
rect 240 1039 244 1043
rect 280 1039 284 1043
rect 344 1039 348 1043
rect 408 1039 412 1043
rect 472 1039 476 1043
rect 536 1039 540 1043
rect 600 1039 604 1043
rect 656 1039 660 1043
rect 664 1039 668 1043
rect 712 1039 716 1043
rect 768 1039 772 1043
rect 776 1039 780 1043
rect 824 1039 828 1043
rect 832 1039 836 1043
rect 888 1039 892 1043
rect 1184 1031 1188 1035
rect 1224 1031 1228 1035
rect 1272 1031 1276 1035
rect 1328 1031 1332 1035
rect 1376 1031 1380 1035
rect 1424 1031 1428 1035
rect 1480 1031 1484 1035
rect 1536 1031 1540 1035
rect 1608 1031 1612 1035
rect 1688 1031 1692 1035
rect 1696 1031 1700 1035
rect 1784 1031 1788 1035
rect 1792 1031 1796 1035
rect 1888 1031 1892 1035
rect 1992 1031 1996 1035
rect 2096 1031 2100 1035
rect 160 1019 164 1023
rect 200 1019 204 1023
rect 240 1019 244 1023
rect 280 1019 284 1023
rect 344 1019 348 1023
rect 408 1019 412 1023
rect 472 1019 476 1023
rect 536 1019 540 1023
rect 600 1019 604 1023
rect 656 1019 660 1023
rect 664 1019 668 1023
rect 712 1019 716 1023
rect 768 1019 772 1023
rect 776 1019 780 1023
rect 824 1019 828 1023
rect 832 1019 836 1023
rect 888 1019 892 1023
rect 1744 1015 1748 1019
rect 1184 1007 1188 1011
rect 1224 1007 1228 1011
rect 1264 1007 1268 1011
rect 1320 1007 1324 1011
rect 1376 1007 1380 1011
rect 1432 1007 1436 1011
rect 1440 1007 1444 1011
rect 1488 1007 1492 1011
rect 1544 1007 1548 1011
rect 1600 1007 1604 1011
rect 1664 1009 1668 1013
rect 1736 1007 1740 1011
rect 1816 1007 1820 1011
rect 1904 1007 1908 1011
rect 1992 1007 1996 1011
rect 2088 1007 2092 1011
rect 1184 987 1188 991
rect 1224 987 1228 991
rect 1264 987 1268 991
rect 1320 987 1324 991
rect 1376 987 1380 991
rect 1432 987 1436 991
rect 1440 987 1444 991
rect 1488 987 1492 991
rect 1544 987 1548 991
rect 1600 987 1604 991
rect 1664 987 1668 991
rect 1736 987 1740 991
rect 1744 987 1748 991
rect 1816 987 1820 991
rect 1904 987 1908 991
rect 1992 987 1996 991
rect 2088 987 2092 991
rect 160 971 164 975
rect 200 971 204 975
rect 208 971 212 975
rect 248 971 252 975
rect 304 971 308 975
rect 368 971 372 975
rect 432 971 436 975
rect 496 971 500 975
rect 552 971 556 975
rect 608 971 612 975
rect 616 971 620 975
rect 656 971 660 975
rect 664 971 668 975
rect 712 971 716 975
rect 720 971 724 975
rect 768 971 772 975
rect 776 971 780 975
rect 824 971 828 975
rect 160 951 164 955
rect 200 951 204 955
rect 208 951 212 955
rect 248 951 252 955
rect 304 951 308 955
rect 368 951 372 955
rect 432 951 436 955
rect 496 951 500 955
rect 552 951 556 955
rect 608 951 612 955
rect 616 951 620 955
rect 656 951 660 955
rect 664 951 668 955
rect 712 951 716 955
rect 720 951 724 955
rect 768 951 772 955
rect 776 951 780 955
rect 824 951 828 955
rect 1184 935 1188 939
rect 1232 935 1236 939
rect 1312 935 1316 939
rect 1400 935 1404 939
rect 1480 935 1484 939
rect 1560 935 1564 939
rect 1640 935 1644 939
rect 1648 935 1652 939
rect 1712 935 1716 939
rect 1720 935 1724 939
rect 1776 935 1780 939
rect 1840 935 1844 939
rect 1904 935 1908 939
rect 1976 935 1980 939
rect 2048 935 2052 939
rect 2096 935 2100 939
rect 288 927 292 931
rect 328 927 332 931
rect 376 927 380 931
rect 424 927 428 931
rect 480 927 484 931
rect 536 927 540 931
rect 592 927 596 931
rect 648 927 652 931
rect 712 927 716 931
rect 776 927 780 931
rect 840 927 844 931
rect 904 927 908 931
rect 968 927 972 931
rect 1032 927 1036 931
rect 1072 927 1076 931
rect 1184 915 1188 919
rect 1232 915 1236 919
rect 1312 915 1316 919
rect 1400 915 1404 919
rect 1480 915 1484 919
rect 1560 915 1564 919
rect 1640 915 1644 919
rect 1648 915 1652 919
rect 1712 915 1716 919
rect 1720 915 1724 919
rect 1776 915 1780 919
rect 1840 915 1844 919
rect 1904 915 1908 919
rect 1976 915 1980 919
rect 2048 915 2052 919
rect 2056 915 2060 919
rect 2096 915 2100 919
rect 288 907 292 911
rect 328 907 332 911
rect 376 907 380 911
rect 424 907 428 911
rect 480 907 484 911
rect 536 907 540 911
rect 592 907 596 911
rect 648 907 652 911
rect 712 907 716 911
rect 776 907 780 911
rect 840 907 844 911
rect 904 907 908 911
rect 968 907 972 911
rect 1032 907 1036 911
rect 1072 907 1076 911
rect 1264 895 1268 899
rect 1344 895 1348 899
rect 1432 895 1436 899
rect 1520 895 1524 899
rect 1608 895 1612 899
rect 1688 895 1692 899
rect 1768 895 1772 899
rect 1840 895 1844 899
rect 1912 895 1916 899
rect 1976 895 1980 899
rect 2048 895 2052 899
rect 1264 875 1268 879
rect 1344 875 1348 879
rect 1432 875 1436 879
rect 1520 875 1524 879
rect 1608 875 1612 879
rect 1688 875 1692 879
rect 1768 875 1772 879
rect 1840 875 1844 879
rect 1912 875 1916 879
rect 1976 875 1980 879
rect 2048 875 2052 879
rect 328 859 332 863
rect 336 859 340 863
rect 376 859 380 863
rect 440 859 444 863
rect 504 859 508 863
rect 576 859 580 863
rect 648 859 652 863
rect 720 859 724 863
rect 792 859 796 863
rect 800 859 804 863
rect 856 859 860 863
rect 864 859 868 863
rect 912 859 916 863
rect 968 859 972 863
rect 976 859 980 863
rect 1032 859 1036 863
rect 1072 859 1076 863
rect 328 839 332 843
rect 336 839 340 843
rect 376 839 380 843
rect 440 839 444 843
rect 504 839 508 843
rect 576 839 580 843
rect 648 839 652 843
rect 720 839 724 843
rect 792 839 796 843
rect 800 839 804 843
rect 856 839 860 843
rect 864 839 868 843
rect 912 839 916 843
rect 968 839 972 843
rect 976 839 980 843
rect 1032 839 1036 843
rect 1072 839 1076 843
rect 2096 895 2100 899
rect 2096 875 2100 879
rect 1184 831 1188 835
rect 1272 831 1276 835
rect 1384 831 1388 835
rect 1480 831 1484 835
rect 1568 831 1572 835
rect 1576 831 1580 835
rect 1656 831 1660 835
rect 1664 831 1668 835
rect 1736 831 1740 835
rect 1808 831 1812 835
rect 1880 831 1884 835
rect 1888 831 1892 835
rect 1960 831 1964 835
rect 2040 831 2044 835
rect 2056 831 2060 835
rect 2096 831 2100 835
rect 2104 831 2108 835
rect 304 819 308 823
rect 368 819 372 823
rect 376 819 380 823
rect 440 819 444 823
rect 512 819 516 823
rect 592 819 596 823
rect 672 819 676 823
rect 752 819 756 823
rect 824 819 828 823
rect 888 819 892 823
rect 896 819 900 823
rect 952 819 956 823
rect 960 819 964 823
rect 1024 819 1028 823
rect 1072 819 1076 823
rect 1184 811 1188 815
rect 1272 811 1276 815
rect 1384 811 1388 815
rect 1480 811 1484 815
rect 1568 811 1572 815
rect 1576 811 1580 815
rect 1656 811 1660 815
rect 1664 811 1668 815
rect 1736 811 1740 815
rect 1808 811 1812 815
rect 1880 811 1884 815
rect 1888 811 1892 815
rect 1960 811 1964 815
rect 2040 811 2044 815
rect 2096 811 2100 815
rect 304 799 308 803
rect 368 799 372 803
rect 376 799 380 803
rect 440 799 444 803
rect 512 799 516 803
rect 592 799 596 803
rect 672 799 676 803
rect 752 799 756 803
rect 824 799 828 803
rect 888 799 892 803
rect 896 799 900 803
rect 952 799 956 803
rect 960 799 964 803
rect 1024 799 1028 803
rect 1072 799 1076 803
rect 1184 791 1188 795
rect 1304 791 1308 795
rect 1432 791 1436 795
rect 1544 791 1548 795
rect 1648 791 1652 795
rect 1656 791 1660 795
rect 1744 791 1748 795
rect 1840 791 1844 795
rect 1928 791 1932 795
rect 2024 791 2028 795
rect 2096 791 2100 795
rect 2104 791 2108 795
rect 1184 771 1188 775
rect 1304 771 1308 775
rect 1400 771 1404 775
rect 1432 771 1436 775
rect 1544 771 1548 775
rect 1648 771 1652 775
rect 1656 771 1660 775
rect 1744 771 1748 775
rect 1840 771 1844 775
rect 1928 771 1932 775
rect 2024 771 2028 775
rect 2096 771 2100 775
rect 240 755 244 759
rect 248 755 252 759
rect 304 755 308 759
rect 312 755 316 759
rect 376 755 380 759
rect 384 755 388 759
rect 448 755 452 759
rect 520 755 524 759
rect 592 755 596 759
rect 664 755 668 759
rect 672 755 676 759
rect 728 755 732 759
rect 784 755 788 759
rect 840 755 844 759
rect 888 755 892 759
rect 936 755 940 759
rect 984 755 988 759
rect 1032 755 1036 759
rect 1072 755 1076 759
rect 240 735 244 739
rect 248 735 252 739
rect 304 735 308 739
rect 312 735 316 739
rect 376 735 380 739
rect 384 735 388 739
rect 448 735 452 739
rect 520 735 524 739
rect 592 735 596 739
rect 664 735 668 739
rect 672 735 676 739
rect 728 735 732 739
rect 784 735 788 739
rect 840 735 844 739
rect 888 735 892 739
rect 936 735 940 739
rect 984 735 988 739
rect 1032 735 1036 739
rect 1072 735 1076 739
rect 1400 731 1404 735
rect 1360 723 1364 727
rect 1400 723 1404 727
rect 1440 723 1444 727
rect 1480 723 1484 727
rect 1488 723 1492 727
rect 1528 723 1532 727
rect 1536 723 1540 727
rect 1576 723 1580 727
rect 1584 723 1588 727
rect 1624 723 1628 727
rect 1680 723 1684 727
rect 1688 723 1692 727
rect 1736 723 1740 727
rect 1792 723 1796 727
rect 1800 723 1804 727
rect 1856 723 1860 727
rect 1920 723 1924 727
rect 1984 723 1988 727
rect 2048 723 2052 727
rect 2056 723 2060 727
rect 2096 723 2100 727
rect 768 719 772 723
rect 200 715 204 719
rect 264 715 268 719
rect 272 715 276 719
rect 336 715 340 719
rect 416 715 420 719
rect 496 715 500 719
rect 504 715 508 719
rect 568 715 572 719
rect 640 715 644 719
rect 704 715 708 719
rect 760 715 764 719
rect 824 715 828 719
rect 888 715 892 719
rect 952 715 956 719
rect 1360 703 1364 707
rect 1400 703 1404 707
rect 1440 703 1444 707
rect 1480 703 1484 707
rect 1488 703 1492 707
rect 1528 703 1532 707
rect 1536 703 1540 707
rect 1576 703 1580 707
rect 1584 703 1588 707
rect 1624 703 1628 707
rect 1680 703 1684 707
rect 1688 703 1692 707
rect 1736 703 1740 707
rect 1792 703 1796 707
rect 1800 703 1804 707
rect 1856 703 1860 707
rect 1920 703 1924 707
rect 1984 703 1988 707
rect 2048 703 2052 707
rect 2056 703 2060 707
rect 2096 703 2100 707
rect 200 695 204 699
rect 264 695 268 699
rect 272 695 276 699
rect 336 695 340 699
rect 416 695 420 699
rect 496 695 500 699
rect 504 695 508 699
rect 568 695 572 699
rect 640 695 644 699
rect 704 695 708 699
rect 760 695 764 699
rect 768 695 772 699
rect 824 695 828 699
rect 888 695 892 699
rect 952 695 956 699
rect 1272 683 1276 687
rect 1312 683 1316 687
rect 1360 683 1364 687
rect 1416 683 1420 687
rect 1472 683 1476 687
rect 1536 683 1540 687
rect 1608 683 1612 687
rect 1680 683 1684 687
rect 1760 683 1764 687
rect 1848 683 1852 687
rect 1936 683 1940 687
rect 2024 683 2028 687
rect 2096 683 2100 687
rect 1272 663 1276 667
rect 1312 663 1316 667
rect 1360 663 1364 667
rect 1416 663 1420 667
rect 1472 663 1476 667
rect 1536 663 1540 667
rect 1608 663 1612 667
rect 1680 663 1684 667
rect 1760 663 1764 667
rect 1848 663 1852 667
rect 1936 663 1940 667
rect 2024 663 2028 667
rect 2096 663 2100 667
rect 160 651 164 655
rect 200 651 204 655
rect 240 651 244 655
rect 248 651 252 655
rect 296 651 300 655
rect 360 651 364 655
rect 424 651 428 655
rect 432 651 436 655
rect 488 651 492 655
rect 552 651 556 655
rect 560 651 564 655
rect 616 651 620 655
rect 672 651 676 655
rect 728 651 732 655
rect 784 651 788 655
rect 792 651 796 655
rect 848 651 852 655
rect 160 631 164 635
rect 200 631 204 635
rect 240 631 244 635
rect 248 631 252 635
rect 296 631 300 635
rect 360 631 364 635
rect 424 631 428 635
rect 432 631 436 635
rect 488 631 492 635
rect 552 631 556 635
rect 560 631 564 635
rect 616 631 620 635
rect 672 631 676 635
rect 728 631 732 635
rect 784 631 788 635
rect 792 631 796 635
rect 848 631 852 635
rect 1184 619 1188 623
rect 1224 619 1228 623
rect 1264 619 1268 623
rect 1304 619 1308 623
rect 1312 619 1316 623
rect 1368 619 1372 623
rect 1376 619 1380 623
rect 1440 619 1444 623
rect 1520 619 1524 623
rect 1528 619 1532 623
rect 1608 619 1612 623
rect 1616 619 1620 623
rect 1696 619 1700 623
rect 1704 619 1708 623
rect 1784 619 1788 623
rect 1864 619 1868 623
rect 1944 619 1948 623
rect 2032 619 2036 623
rect 2096 619 2100 623
rect 160 603 164 607
rect 200 603 204 607
rect 240 603 244 607
rect 280 603 284 607
rect 328 603 332 607
rect 376 603 380 607
rect 424 603 428 607
rect 464 603 468 607
rect 512 603 516 607
rect 560 603 564 607
rect 568 603 572 607
rect 608 603 612 607
rect 656 603 660 607
rect 704 603 708 607
rect 752 603 756 607
rect 1184 599 1188 603
rect 1224 599 1228 603
rect 1264 599 1268 603
rect 1304 599 1308 603
rect 1312 599 1316 603
rect 1368 599 1372 603
rect 1376 599 1380 603
rect 1440 599 1444 603
rect 1520 599 1524 603
rect 1528 599 1532 603
rect 1608 599 1612 603
rect 1616 599 1620 603
rect 1696 599 1700 603
rect 1704 599 1708 603
rect 1784 599 1788 603
rect 1864 599 1868 603
rect 1944 599 1948 603
rect 2032 599 2036 603
rect 2096 599 2100 603
rect 160 583 164 587
rect 200 583 204 587
rect 240 583 244 587
rect 280 583 284 587
rect 328 583 332 587
rect 376 583 380 587
rect 424 583 428 587
rect 464 583 468 587
rect 512 583 516 587
rect 560 583 564 587
rect 568 583 572 587
rect 608 583 612 587
rect 656 583 660 587
rect 704 583 708 587
rect 752 583 756 587
rect 1184 575 1188 579
rect 1224 575 1228 579
rect 1264 575 1268 579
rect 1304 575 1308 579
rect 1344 575 1348 579
rect 1384 575 1388 579
rect 1392 575 1396 579
rect 1440 575 1444 579
rect 1512 575 1516 579
rect 1552 575 1556 579
rect 1592 575 1596 579
rect 1680 575 1684 579
rect 1776 575 1780 579
rect 1880 575 1884 579
rect 1992 575 1996 579
rect 2096 575 2100 579
rect 1184 555 1188 559
rect 1224 555 1228 559
rect 1264 555 1268 559
rect 1304 555 1308 559
rect 1344 555 1348 559
rect 1384 555 1388 559
rect 1392 555 1396 559
rect 1440 555 1444 559
rect 1512 555 1516 559
rect 1552 555 1556 559
rect 1592 555 1596 559
rect 1680 555 1684 559
rect 1776 555 1780 559
rect 1880 555 1884 559
rect 1992 555 1996 559
rect 2040 555 2044 559
rect 2096 555 2100 559
rect 160 535 164 539
rect 200 535 204 539
rect 248 535 252 539
rect 304 535 308 539
rect 352 535 356 539
rect 400 535 404 539
rect 448 535 452 539
rect 488 535 492 539
rect 536 535 540 539
rect 544 535 548 539
rect 584 535 588 539
rect 592 535 596 539
rect 632 535 636 539
rect 640 535 644 539
rect 680 535 684 539
rect 728 535 732 539
rect 736 535 740 539
rect 776 535 780 539
rect 160 515 164 519
rect 200 515 204 519
rect 248 515 252 519
rect 304 515 308 519
rect 352 515 356 519
rect 400 515 404 519
rect 448 515 452 519
rect 488 515 492 519
rect 536 515 540 519
rect 544 515 548 519
rect 584 515 588 519
rect 592 515 596 519
rect 632 515 636 519
rect 640 515 644 519
rect 680 515 684 519
rect 728 515 732 519
rect 736 515 740 519
rect 776 515 780 519
rect 1328 507 1332 511
rect 1368 507 1372 511
rect 1408 507 1412 511
rect 1448 507 1452 511
rect 1488 507 1492 511
rect 1528 507 1532 511
rect 1568 507 1572 511
rect 1616 507 1620 511
rect 1672 507 1676 511
rect 1728 507 1732 511
rect 1792 507 1796 511
rect 1864 507 1868 511
rect 1944 507 1948 511
rect 2032 507 2036 511
rect 2096 507 2100 511
rect 160 487 164 491
rect 200 487 204 491
rect 256 487 260 491
rect 320 487 324 491
rect 384 487 388 491
rect 448 487 452 491
rect 504 487 508 491
rect 560 487 564 491
rect 616 487 620 491
rect 664 487 668 491
rect 712 487 716 491
rect 760 487 764 491
rect 816 487 820 491
rect 872 487 876 491
rect 1328 487 1332 491
rect 1368 487 1372 491
rect 1408 487 1412 491
rect 1448 487 1452 491
rect 1488 487 1492 491
rect 1528 487 1532 491
rect 1568 487 1572 491
rect 1616 487 1620 491
rect 1672 487 1676 491
rect 1728 487 1732 491
rect 1792 487 1796 491
rect 1864 487 1868 491
rect 1944 487 1948 491
rect 2032 487 2036 491
rect 2040 487 2044 491
rect 2096 487 2100 491
rect 160 467 164 471
rect 200 467 204 471
rect 256 467 260 471
rect 320 467 324 471
rect 384 467 388 471
rect 448 467 452 471
rect 504 467 508 471
rect 560 469 564 473
rect 616 467 620 471
rect 664 467 668 471
rect 712 467 716 471
rect 760 467 764 471
rect 816 467 820 471
rect 872 467 876 471
rect 1320 467 1324 471
rect 1360 467 1364 471
rect 1400 467 1404 471
rect 1448 467 1452 471
rect 1496 467 1500 471
rect 1552 467 1556 471
rect 1608 467 1612 471
rect 1672 467 1676 471
rect 1744 467 1748 471
rect 1832 467 1836 471
rect 1920 467 1924 471
rect 2016 467 2020 471
rect 2096 467 2100 471
rect 1320 447 1324 451
rect 1360 447 1364 451
rect 1400 447 1404 451
rect 1448 447 1452 451
rect 1496 447 1500 451
rect 1552 447 1556 451
rect 1608 447 1612 451
rect 1672 447 1676 451
rect 1744 447 1748 451
rect 1832 447 1836 451
rect 1920 447 1924 451
rect 2016 447 2020 451
rect 2096 447 2100 451
rect 200 419 204 423
rect 240 419 244 423
rect 288 419 292 423
rect 352 419 356 423
rect 360 419 364 423
rect 416 419 420 423
rect 488 419 492 423
rect 560 419 564 423
rect 632 419 636 423
rect 640 419 644 423
rect 704 419 708 423
rect 712 419 716 423
rect 768 419 772 423
rect 776 419 780 423
rect 832 419 836 423
rect 840 419 844 423
rect 896 419 900 423
rect 904 419 908 423
rect 968 419 972 423
rect 1184 405 1188 409
rect 1224 403 1228 407
rect 1232 403 1236 407
rect 1280 403 1284 407
rect 1288 403 1292 407
rect 1360 403 1364 407
rect 1368 403 1372 407
rect 1440 403 1444 407
rect 1448 403 1452 407
rect 1528 403 1532 407
rect 1616 403 1620 407
rect 1696 403 1700 407
rect 1776 403 1780 407
rect 1784 403 1788 407
rect 1856 403 1860 407
rect 1936 403 1940 407
rect 2024 403 2028 407
rect 2096 403 2100 407
rect 2104 403 2108 407
rect 200 399 204 403
rect 240 399 244 403
rect 288 399 292 403
rect 352 399 356 403
rect 360 399 364 403
rect 416 399 420 403
rect 488 399 492 403
rect 560 399 564 403
rect 632 399 636 403
rect 640 399 644 403
rect 704 399 708 403
rect 712 399 716 403
rect 768 399 772 403
rect 776 399 780 403
rect 832 399 836 403
rect 840 399 844 403
rect 896 399 900 403
rect 904 399 908 403
rect 968 399 972 403
rect 1184 383 1188 387
rect 1224 383 1228 387
rect 1232 383 1236 387
rect 1280 383 1284 387
rect 1288 383 1292 387
rect 1360 383 1364 387
rect 1368 383 1372 387
rect 1440 383 1444 387
rect 1448 383 1452 387
rect 1528 383 1532 387
rect 1616 383 1620 387
rect 1696 383 1700 387
rect 1776 383 1780 387
rect 1784 383 1788 387
rect 1856 383 1860 387
rect 1936 383 1940 387
rect 2024 383 2028 387
rect 2096 383 2100 387
rect 200 371 204 375
rect 240 371 244 375
rect 248 371 252 375
rect 296 371 300 375
rect 304 371 308 375
rect 360 371 364 375
rect 432 371 436 375
rect 512 371 516 375
rect 592 371 596 375
rect 664 371 668 375
rect 736 371 740 375
rect 800 371 804 375
rect 864 371 868 375
rect 920 371 924 375
rect 976 371 980 375
rect 1032 371 1036 375
rect 1072 371 1076 375
rect 1184 359 1188 363
rect 1272 359 1276 363
rect 1384 359 1388 363
rect 1488 359 1492 363
rect 1584 359 1588 363
rect 1672 361 1676 365
rect 1752 359 1756 363
rect 1760 359 1764 363
rect 1824 359 1828 363
rect 1832 359 1836 363
rect 1888 359 1892 363
rect 1944 359 1948 363
rect 2000 359 2004 363
rect 2056 359 2060 363
rect 2096 359 2100 363
rect 2104 359 2108 363
rect 200 351 204 355
rect 240 351 244 355
rect 248 351 252 355
rect 296 351 300 355
rect 304 351 308 355
rect 360 351 364 355
rect 432 351 436 355
rect 512 351 516 355
rect 592 351 596 355
rect 664 351 668 355
rect 736 351 740 355
rect 800 351 804 355
rect 864 351 868 355
rect 920 351 924 355
rect 976 351 980 355
rect 1032 351 1036 355
rect 1072 351 1076 355
rect 1184 339 1188 343
rect 1272 339 1276 343
rect 1384 339 1388 343
rect 1488 339 1492 343
rect 1584 339 1588 343
rect 1672 339 1676 343
rect 1752 339 1756 343
rect 1760 339 1764 343
rect 1824 339 1828 343
rect 1832 339 1836 343
rect 1888 339 1892 343
rect 1944 339 1948 343
rect 2000 339 2004 343
rect 2056 339 2060 343
rect 2096 339 2100 343
rect 408 303 412 307
rect 448 303 452 307
rect 488 303 492 307
rect 528 303 532 307
rect 568 303 572 307
rect 576 303 580 307
rect 616 303 620 307
rect 624 303 628 307
rect 664 303 668 307
rect 672 303 676 307
rect 712 303 716 307
rect 760 303 764 307
rect 808 303 812 307
rect 816 303 820 307
rect 856 303 860 307
rect 864 303 868 307
rect 904 303 908 307
rect 952 303 956 307
rect 992 303 996 307
rect 1032 303 1036 307
rect 1072 303 1076 307
rect 1376 287 1380 291
rect 1416 287 1420 291
rect 1456 287 1460 291
rect 1496 287 1500 291
rect 1536 287 1540 291
rect 1544 287 1548 291
rect 1584 287 1588 291
rect 1592 287 1596 291
rect 1640 287 1644 291
rect 1648 287 1652 291
rect 1696 287 1700 291
rect 1760 287 1764 291
rect 1768 287 1772 291
rect 1832 287 1836 291
rect 1912 287 1916 291
rect 1992 287 1996 291
rect 2072 287 2076 291
rect 408 283 412 287
rect 448 283 452 287
rect 488 283 492 287
rect 528 283 532 287
rect 568 283 572 287
rect 576 283 580 287
rect 616 283 620 287
rect 624 283 628 287
rect 664 283 668 287
rect 672 283 676 287
rect 712 283 716 287
rect 760 283 764 287
rect 808 283 812 287
rect 816 283 820 287
rect 856 283 860 287
rect 864 283 868 287
rect 904 283 908 287
rect 952 283 956 287
rect 992 283 996 287
rect 1032 283 1036 287
rect 1072 283 1076 287
rect 1376 267 1380 271
rect 1416 267 1420 271
rect 1456 267 1460 271
rect 1496 267 1500 271
rect 1536 267 1540 271
rect 1544 267 1548 271
rect 1584 267 1588 271
rect 1592 267 1596 271
rect 1640 267 1644 271
rect 1648 267 1652 271
rect 1696 267 1700 271
rect 1760 267 1764 271
rect 1768 267 1772 271
rect 1832 267 1836 271
rect 1912 267 1916 271
rect 1992 267 1996 271
rect 2072 267 2076 271
rect 312 255 316 259
rect 352 255 356 259
rect 392 255 396 259
rect 440 255 444 259
rect 496 255 500 259
rect 560 255 564 259
rect 632 255 636 259
rect 704 255 708 259
rect 768 255 772 259
rect 832 255 836 259
rect 888 255 892 259
rect 952 255 956 259
rect 1016 255 1020 259
rect 1072 255 1076 259
rect 1288 247 1292 251
rect 1328 247 1332 251
rect 1368 247 1372 251
rect 1408 247 1412 251
rect 1448 247 1452 251
rect 1488 247 1492 251
rect 1528 247 1532 251
rect 1568 247 1572 251
rect 1624 247 1628 251
rect 1696 247 1700 251
rect 1784 247 1788 251
rect 1888 247 1892 251
rect 1960 247 1964 251
rect 2000 247 2004 251
rect 2096 247 2100 251
rect 312 235 316 239
rect 352 235 356 239
rect 392 235 396 239
rect 440 235 444 239
rect 496 235 500 239
rect 560 235 564 239
rect 632 235 636 239
rect 704 235 708 239
rect 768 235 772 239
rect 832 235 836 239
rect 888 235 892 239
rect 952 235 956 239
rect 1016 235 1020 239
rect 1072 235 1076 239
rect 1288 227 1292 231
rect 1328 227 1332 231
rect 1368 227 1372 231
rect 1408 227 1412 231
rect 1448 227 1452 231
rect 1488 227 1492 231
rect 1528 227 1532 231
rect 1568 227 1572 231
rect 1624 227 1628 231
rect 1696 227 1700 231
rect 1784 227 1788 231
rect 1888 227 1892 231
rect 1960 227 1964 231
rect 2000 227 2004 231
rect 2096 227 2100 231
rect 192 179 196 183
rect 232 179 236 183
rect 272 179 276 183
rect 280 179 284 183
rect 320 179 324 183
rect 328 179 332 183
rect 368 179 372 183
rect 376 179 380 183
rect 424 179 428 183
rect 432 179 436 183
rect 488 179 492 183
rect 552 179 556 183
rect 624 179 628 183
rect 696 179 700 183
rect 776 179 780 183
rect 856 179 860 183
rect 936 179 940 183
rect 1016 179 1020 183
rect 1072 179 1076 183
rect 1208 179 1212 183
rect 1256 179 1260 183
rect 1264 179 1268 183
rect 1320 179 1324 183
rect 1328 179 1332 183
rect 1384 179 1388 183
rect 1392 179 1396 183
rect 1456 179 1460 183
rect 1464 179 1468 183
rect 1536 179 1540 183
rect 1616 179 1620 183
rect 1624 179 1628 183
rect 1688 179 1692 183
rect 1696 179 1700 183
rect 1760 179 1764 183
rect 1768 179 1772 183
rect 1832 179 1836 183
rect 1904 179 1908 183
rect 1912 179 1916 183
rect 1976 179 1980 183
rect 2048 179 2052 183
rect 2096 179 2100 183
rect 192 159 196 163
rect 232 159 236 163
rect 272 159 276 163
rect 280 159 284 163
rect 320 159 324 163
rect 328 159 332 163
rect 368 159 372 163
rect 376 159 380 163
rect 424 159 428 163
rect 432 159 436 163
rect 488 159 492 163
rect 552 159 556 163
rect 624 159 628 163
rect 696 159 700 163
rect 776 159 780 163
rect 856 159 860 163
rect 936 159 940 163
rect 1016 159 1020 163
rect 1072 159 1076 163
rect 1208 159 1212 163
rect 1256 159 1260 163
rect 1264 159 1268 163
rect 1320 159 1324 163
rect 1328 159 1332 163
rect 1384 159 1388 163
rect 1392 159 1396 163
rect 1456 159 1460 163
rect 1464 159 1468 163
rect 1536 159 1540 163
rect 1616 159 1620 163
rect 1624 159 1628 163
rect 1688 159 1692 163
rect 1696 159 1700 163
rect 1760 159 1764 163
rect 1768 159 1772 163
rect 1832 159 1836 163
rect 1904 159 1908 163
rect 1912 159 1916 163
rect 1976 159 1980 163
rect 2048 159 2052 163
rect 2096 159 2100 163
rect 160 123 164 127
rect 200 123 204 127
rect 240 123 244 127
rect 280 123 284 127
rect 320 123 324 127
rect 360 123 364 127
rect 400 123 404 127
rect 440 123 444 127
rect 480 123 484 127
rect 520 123 524 127
rect 560 123 564 127
rect 600 123 604 127
rect 640 123 644 127
rect 680 123 684 127
rect 720 123 724 127
rect 760 123 764 127
rect 800 123 804 127
rect 840 123 844 127
rect 896 123 900 127
rect 960 123 964 127
rect 1024 123 1028 127
rect 1072 123 1076 127
rect 1184 115 1188 119
rect 1224 115 1228 119
rect 1264 115 1268 119
rect 1304 115 1308 119
rect 1344 115 1348 119
rect 1392 115 1396 119
rect 1456 115 1460 119
rect 1520 115 1524 119
rect 1584 115 1588 119
rect 1640 115 1644 119
rect 1696 115 1700 119
rect 1744 115 1748 119
rect 1792 115 1796 119
rect 1832 115 1836 119
rect 1880 115 1884 119
rect 1928 115 1932 119
rect 1976 115 1980 119
rect 2016 115 2020 119
rect 2056 115 2060 119
rect 2096 115 2100 119
rect 200 103 204 107
rect 240 103 244 107
rect 280 103 284 107
rect 320 103 324 107
rect 360 103 364 107
rect 400 103 404 107
rect 440 103 444 107
rect 480 103 484 107
rect 520 103 524 107
rect 560 103 564 107
rect 600 103 604 107
rect 640 103 644 107
rect 680 103 684 107
rect 720 103 724 107
rect 760 103 764 107
rect 800 103 804 107
rect 840 103 844 107
rect 896 103 900 107
rect 960 103 964 107
rect 1024 103 1028 107
rect 1072 103 1076 107
rect 1184 95 1188 99
rect 1224 95 1228 99
rect 1264 95 1268 99
rect 1304 95 1308 99
rect 1344 95 1348 99
rect 1392 95 1396 99
rect 1456 95 1460 99
rect 1520 95 1524 99
rect 1584 95 1588 99
rect 1640 95 1644 99
rect 1696 95 1700 99
rect 1744 95 1748 99
rect 1792 95 1796 99
rect 1832 95 1836 99
rect 1880 95 1884 99
rect 1928 95 1932 99
rect 1976 95 1980 99
rect 2016 95 2020 99
rect 2056 95 2060 99
rect 2096 95 2100 99
<< m2 >>
rect 1646 2211 1652 2212
rect 1646 2207 1647 2211
rect 1651 2210 1652 2211
rect 1651 2208 1850 2210
rect 1651 2207 1652 2208
rect 1646 2206 1652 2207
rect 1848 2204 1850 2208
rect 1367 2203 1373 2204
rect 1367 2199 1368 2203
rect 1372 2202 1373 2203
rect 1398 2203 1404 2204
rect 1398 2202 1399 2203
rect 1372 2200 1399 2202
rect 1372 2199 1373 2200
rect 1367 2198 1373 2199
rect 1398 2199 1399 2200
rect 1403 2199 1404 2203
rect 1398 2198 1404 2199
rect 1407 2203 1413 2204
rect 1407 2199 1408 2203
rect 1412 2202 1413 2203
rect 1438 2203 1444 2204
rect 1438 2202 1439 2203
rect 1412 2200 1439 2202
rect 1412 2199 1413 2200
rect 1407 2198 1413 2199
rect 1438 2199 1439 2200
rect 1443 2199 1444 2203
rect 1438 2198 1444 2199
rect 1447 2203 1453 2204
rect 1447 2199 1448 2203
rect 1452 2202 1453 2203
rect 1478 2203 1484 2204
rect 1478 2202 1479 2203
rect 1452 2200 1479 2202
rect 1452 2199 1453 2200
rect 1447 2198 1453 2199
rect 1478 2199 1479 2200
rect 1483 2199 1484 2203
rect 1478 2198 1484 2199
rect 1487 2203 1493 2204
rect 1487 2199 1488 2203
rect 1492 2202 1493 2203
rect 1518 2203 1524 2204
rect 1518 2202 1519 2203
rect 1492 2200 1519 2202
rect 1492 2199 1493 2200
rect 1487 2198 1493 2199
rect 1518 2199 1519 2200
rect 1523 2199 1524 2203
rect 1518 2198 1524 2199
rect 1527 2203 1533 2204
rect 1527 2199 1528 2203
rect 1532 2202 1533 2203
rect 1558 2203 1564 2204
rect 1558 2202 1559 2203
rect 1532 2200 1559 2202
rect 1532 2199 1533 2200
rect 1527 2198 1533 2199
rect 1558 2199 1559 2200
rect 1563 2199 1564 2203
rect 1558 2198 1564 2199
rect 1567 2203 1573 2204
rect 1567 2199 1568 2203
rect 1572 2202 1573 2203
rect 1598 2203 1604 2204
rect 1598 2202 1599 2203
rect 1572 2200 1599 2202
rect 1572 2199 1573 2200
rect 1567 2198 1573 2199
rect 1598 2199 1599 2200
rect 1603 2199 1604 2203
rect 1598 2198 1604 2199
rect 1607 2203 1613 2204
rect 1607 2199 1608 2203
rect 1612 2202 1613 2203
rect 1638 2203 1644 2204
rect 1638 2202 1639 2203
rect 1612 2200 1639 2202
rect 1612 2199 1613 2200
rect 1607 2198 1613 2199
rect 1638 2199 1639 2200
rect 1643 2199 1644 2203
rect 1638 2198 1644 2199
rect 1647 2203 1653 2204
rect 1647 2199 1648 2203
rect 1652 2202 1653 2203
rect 1678 2203 1684 2204
rect 1678 2202 1679 2203
rect 1652 2200 1679 2202
rect 1652 2199 1653 2200
rect 1647 2198 1653 2199
rect 1678 2199 1679 2200
rect 1683 2199 1684 2203
rect 1678 2198 1684 2199
rect 1687 2203 1693 2204
rect 1687 2199 1688 2203
rect 1692 2202 1693 2203
rect 1718 2203 1724 2204
rect 1718 2202 1719 2203
rect 1692 2200 1719 2202
rect 1692 2199 1693 2200
rect 1687 2198 1693 2199
rect 1718 2199 1719 2200
rect 1723 2199 1724 2203
rect 1718 2198 1724 2199
rect 1727 2203 1733 2204
rect 1727 2199 1728 2203
rect 1732 2202 1733 2203
rect 1758 2203 1764 2204
rect 1758 2202 1759 2203
rect 1732 2200 1759 2202
rect 1732 2199 1733 2200
rect 1727 2198 1733 2199
rect 1758 2199 1759 2200
rect 1763 2199 1764 2203
rect 1758 2198 1764 2199
rect 1767 2203 1773 2204
rect 1767 2199 1768 2203
rect 1772 2202 1773 2203
rect 1798 2203 1804 2204
rect 1798 2202 1799 2203
rect 1772 2200 1799 2202
rect 1772 2199 1773 2200
rect 1767 2198 1773 2199
rect 1798 2199 1799 2200
rect 1803 2199 1804 2203
rect 1798 2198 1804 2199
rect 1807 2203 1813 2204
rect 1807 2199 1808 2203
rect 1812 2202 1813 2203
rect 1838 2203 1844 2204
rect 1838 2202 1839 2203
rect 1812 2200 1839 2202
rect 1812 2199 1813 2200
rect 1807 2198 1813 2199
rect 1838 2199 1839 2200
rect 1843 2199 1844 2203
rect 1838 2198 1844 2199
rect 1847 2203 1853 2204
rect 1847 2199 1848 2203
rect 1852 2199 1853 2203
rect 1847 2198 1853 2199
rect 1342 2196 1348 2197
rect 1342 2192 1343 2196
rect 1347 2192 1348 2196
rect 1342 2191 1348 2192
rect 1382 2196 1388 2197
rect 1382 2192 1383 2196
rect 1387 2192 1388 2196
rect 1382 2191 1388 2192
rect 1422 2196 1428 2197
rect 1422 2192 1423 2196
rect 1427 2192 1428 2196
rect 1422 2191 1428 2192
rect 1462 2196 1468 2197
rect 1462 2192 1463 2196
rect 1467 2192 1468 2196
rect 1462 2191 1468 2192
rect 1502 2196 1508 2197
rect 1502 2192 1503 2196
rect 1507 2192 1508 2196
rect 1502 2191 1508 2192
rect 1542 2196 1548 2197
rect 1542 2192 1543 2196
rect 1547 2192 1548 2196
rect 1542 2191 1548 2192
rect 1582 2196 1588 2197
rect 1582 2192 1583 2196
rect 1587 2192 1588 2196
rect 1582 2191 1588 2192
rect 1622 2196 1628 2197
rect 1622 2192 1623 2196
rect 1627 2192 1628 2196
rect 1622 2191 1628 2192
rect 1662 2196 1668 2197
rect 1662 2192 1663 2196
rect 1667 2192 1668 2196
rect 1662 2191 1668 2192
rect 1702 2196 1708 2197
rect 1702 2192 1703 2196
rect 1707 2192 1708 2196
rect 1702 2191 1708 2192
rect 1742 2196 1748 2197
rect 1742 2192 1743 2196
rect 1747 2192 1748 2196
rect 1742 2191 1748 2192
rect 1782 2196 1788 2197
rect 1782 2192 1783 2196
rect 1787 2192 1788 2196
rect 1782 2191 1788 2192
rect 1822 2196 1828 2197
rect 1822 2192 1823 2196
rect 1827 2192 1828 2196
rect 1822 2191 1828 2192
rect 1134 2188 1140 2189
rect 1134 2184 1135 2188
rect 1139 2184 1140 2188
rect 2118 2188 2124 2189
rect 2118 2184 2119 2188
rect 2123 2184 2124 2188
rect 1134 2183 1140 2184
rect 1367 2183 1373 2184
rect 1367 2179 1368 2183
rect 1372 2182 1373 2183
rect 1390 2183 1396 2184
rect 1390 2182 1391 2183
rect 1372 2180 1391 2182
rect 1372 2179 1373 2180
rect 1367 2178 1373 2179
rect 1390 2179 1391 2180
rect 1395 2179 1396 2183
rect 1390 2178 1396 2179
rect 1398 2183 1404 2184
rect 1398 2179 1399 2183
rect 1403 2182 1404 2183
rect 1407 2183 1413 2184
rect 1407 2182 1408 2183
rect 1403 2180 1408 2182
rect 1403 2179 1404 2180
rect 1398 2178 1404 2179
rect 1407 2179 1408 2180
rect 1412 2179 1413 2183
rect 1407 2178 1413 2179
rect 1438 2183 1444 2184
rect 1438 2179 1439 2183
rect 1443 2182 1444 2183
rect 1447 2183 1453 2184
rect 1447 2182 1448 2183
rect 1443 2180 1448 2182
rect 1443 2179 1444 2180
rect 1438 2178 1444 2179
rect 1447 2179 1448 2180
rect 1452 2179 1453 2183
rect 1447 2178 1453 2179
rect 1478 2183 1484 2184
rect 1478 2179 1479 2183
rect 1483 2182 1484 2183
rect 1487 2183 1493 2184
rect 1487 2182 1488 2183
rect 1483 2180 1488 2182
rect 1483 2179 1484 2180
rect 1478 2178 1484 2179
rect 1487 2179 1488 2180
rect 1492 2179 1493 2183
rect 1487 2178 1493 2179
rect 1518 2183 1524 2184
rect 1518 2179 1519 2183
rect 1523 2182 1524 2183
rect 1527 2183 1533 2184
rect 1527 2182 1528 2183
rect 1523 2180 1528 2182
rect 1523 2179 1524 2180
rect 1518 2178 1524 2179
rect 1527 2179 1528 2180
rect 1532 2179 1533 2183
rect 1527 2178 1533 2179
rect 1558 2183 1564 2184
rect 1558 2179 1559 2183
rect 1563 2182 1564 2183
rect 1567 2183 1573 2184
rect 1567 2182 1568 2183
rect 1563 2180 1568 2182
rect 1563 2179 1564 2180
rect 1558 2178 1564 2179
rect 1567 2179 1568 2180
rect 1572 2179 1573 2183
rect 1567 2178 1573 2179
rect 1598 2183 1604 2184
rect 1598 2179 1599 2183
rect 1603 2182 1604 2183
rect 1607 2183 1613 2184
rect 1607 2182 1608 2183
rect 1603 2180 1608 2182
rect 1603 2179 1604 2180
rect 1598 2178 1604 2179
rect 1607 2179 1608 2180
rect 1612 2179 1613 2183
rect 1607 2178 1613 2179
rect 1638 2183 1644 2184
rect 1638 2179 1639 2183
rect 1643 2182 1644 2183
rect 1647 2183 1653 2184
rect 1647 2182 1648 2183
rect 1643 2180 1648 2182
rect 1643 2179 1644 2180
rect 1638 2178 1644 2179
rect 1647 2179 1648 2180
rect 1652 2179 1653 2183
rect 1647 2178 1653 2179
rect 1678 2183 1684 2184
rect 1678 2179 1679 2183
rect 1683 2182 1684 2183
rect 1687 2183 1693 2184
rect 1687 2182 1688 2183
rect 1683 2180 1688 2182
rect 1683 2179 1684 2180
rect 1678 2178 1684 2179
rect 1687 2179 1688 2180
rect 1692 2179 1693 2183
rect 1687 2178 1693 2179
rect 1718 2183 1724 2184
rect 1718 2179 1719 2183
rect 1723 2182 1724 2183
rect 1727 2183 1733 2184
rect 1727 2182 1728 2183
rect 1723 2180 1728 2182
rect 1723 2179 1724 2180
rect 1718 2178 1724 2179
rect 1727 2179 1728 2180
rect 1732 2179 1733 2183
rect 1727 2178 1733 2179
rect 1758 2183 1764 2184
rect 1758 2179 1759 2183
rect 1763 2182 1764 2183
rect 1767 2183 1773 2184
rect 1767 2182 1768 2183
rect 1763 2180 1768 2182
rect 1763 2179 1764 2180
rect 1758 2178 1764 2179
rect 1767 2179 1768 2180
rect 1772 2179 1773 2183
rect 1767 2178 1773 2179
rect 1798 2183 1804 2184
rect 1798 2179 1799 2183
rect 1803 2182 1804 2183
rect 1807 2183 1813 2184
rect 1807 2182 1808 2183
rect 1803 2180 1808 2182
rect 1803 2179 1804 2180
rect 1798 2178 1804 2179
rect 1807 2179 1808 2180
rect 1812 2179 1813 2183
rect 1807 2178 1813 2179
rect 1838 2183 1844 2184
rect 1838 2179 1839 2183
rect 1843 2182 1844 2183
rect 1847 2183 1853 2184
rect 2118 2183 2124 2184
rect 1847 2182 1848 2183
rect 1843 2180 1848 2182
rect 1843 2179 1844 2180
rect 1838 2178 1844 2179
rect 1847 2179 1848 2180
rect 1852 2179 1853 2183
rect 1847 2178 1853 2179
rect 1134 2171 1140 2172
rect 1134 2167 1135 2171
rect 1139 2167 1140 2171
rect 2118 2171 2124 2172
rect 1134 2166 1140 2167
rect 1342 2168 1348 2169
rect 1342 2164 1343 2168
rect 1347 2164 1348 2168
rect 1342 2163 1348 2164
rect 1382 2168 1388 2169
rect 1382 2164 1383 2168
rect 1387 2164 1388 2168
rect 1382 2163 1388 2164
rect 1422 2168 1428 2169
rect 1422 2164 1423 2168
rect 1427 2164 1428 2168
rect 1422 2163 1428 2164
rect 1462 2168 1468 2169
rect 1462 2164 1463 2168
rect 1467 2164 1468 2168
rect 1462 2163 1468 2164
rect 1502 2168 1508 2169
rect 1502 2164 1503 2168
rect 1507 2164 1508 2168
rect 1502 2163 1508 2164
rect 1542 2168 1548 2169
rect 1542 2164 1543 2168
rect 1547 2164 1548 2168
rect 1542 2163 1548 2164
rect 1582 2168 1588 2169
rect 1582 2164 1583 2168
rect 1587 2164 1588 2168
rect 1582 2163 1588 2164
rect 1622 2168 1628 2169
rect 1622 2164 1623 2168
rect 1627 2164 1628 2168
rect 1622 2163 1628 2164
rect 1662 2168 1668 2169
rect 1662 2164 1663 2168
rect 1667 2164 1668 2168
rect 1662 2163 1668 2164
rect 1702 2168 1708 2169
rect 1702 2164 1703 2168
rect 1707 2164 1708 2168
rect 1702 2163 1708 2164
rect 1742 2168 1748 2169
rect 1742 2164 1743 2168
rect 1747 2164 1748 2168
rect 1742 2163 1748 2164
rect 1782 2168 1788 2169
rect 1782 2164 1783 2168
rect 1787 2164 1788 2168
rect 1782 2163 1788 2164
rect 1822 2168 1828 2169
rect 1822 2164 1823 2168
rect 1827 2164 1828 2168
rect 2118 2167 2119 2171
rect 2123 2167 2124 2171
rect 2118 2166 2124 2167
rect 1822 2163 1828 2164
rect 1286 2156 1292 2157
rect 1134 2153 1140 2154
rect 1134 2149 1135 2153
rect 1139 2149 1140 2153
rect 1286 2152 1287 2156
rect 1291 2152 1292 2156
rect 1286 2151 1292 2152
rect 1326 2156 1332 2157
rect 1326 2152 1327 2156
rect 1331 2152 1332 2156
rect 1326 2151 1332 2152
rect 1366 2156 1372 2157
rect 1366 2152 1367 2156
rect 1371 2152 1372 2156
rect 1366 2151 1372 2152
rect 1414 2156 1420 2157
rect 1414 2152 1415 2156
rect 1419 2152 1420 2156
rect 1414 2151 1420 2152
rect 1462 2156 1468 2157
rect 1462 2152 1463 2156
rect 1467 2152 1468 2156
rect 1462 2151 1468 2152
rect 1518 2156 1524 2157
rect 1518 2152 1519 2156
rect 1523 2152 1524 2156
rect 1518 2151 1524 2152
rect 1574 2156 1580 2157
rect 1574 2152 1575 2156
rect 1579 2152 1580 2156
rect 1574 2151 1580 2152
rect 1622 2156 1628 2157
rect 1622 2152 1623 2156
rect 1627 2152 1628 2156
rect 1622 2151 1628 2152
rect 1670 2156 1676 2157
rect 1670 2152 1671 2156
rect 1675 2152 1676 2156
rect 1670 2151 1676 2152
rect 1718 2156 1724 2157
rect 1718 2152 1719 2156
rect 1723 2152 1724 2156
rect 1718 2151 1724 2152
rect 1774 2156 1780 2157
rect 1774 2152 1775 2156
rect 1779 2152 1780 2156
rect 1774 2151 1780 2152
rect 1830 2156 1836 2157
rect 1830 2152 1831 2156
rect 1835 2152 1836 2156
rect 1830 2151 1836 2152
rect 1886 2156 1892 2157
rect 1886 2152 1887 2156
rect 1891 2152 1892 2156
rect 1886 2151 1892 2152
rect 2118 2153 2124 2154
rect 1134 2148 1140 2149
rect 2118 2149 2119 2153
rect 2123 2149 2124 2153
rect 2118 2148 2124 2149
rect 1311 2139 1320 2140
rect 1134 2136 1140 2137
rect 1134 2132 1135 2136
rect 1139 2132 1140 2136
rect 1311 2135 1312 2139
rect 1319 2135 1320 2139
rect 1311 2134 1320 2135
rect 1334 2139 1340 2140
rect 1334 2135 1335 2139
rect 1339 2138 1340 2139
rect 1351 2139 1357 2140
rect 1351 2138 1352 2139
rect 1339 2136 1352 2138
rect 1339 2135 1340 2136
rect 1334 2134 1340 2135
rect 1351 2135 1352 2136
rect 1356 2135 1357 2139
rect 1351 2134 1357 2135
rect 1374 2139 1380 2140
rect 1374 2135 1375 2139
rect 1379 2138 1380 2139
rect 1391 2139 1397 2140
rect 1391 2138 1392 2139
rect 1379 2136 1392 2138
rect 1379 2135 1380 2136
rect 1374 2134 1380 2135
rect 1391 2135 1392 2136
rect 1396 2135 1397 2139
rect 1391 2134 1397 2135
rect 1399 2139 1405 2140
rect 1399 2135 1400 2139
rect 1404 2138 1405 2139
rect 1439 2139 1445 2140
rect 1439 2138 1440 2139
rect 1404 2136 1440 2138
rect 1404 2135 1405 2136
rect 1399 2134 1405 2135
rect 1439 2135 1440 2136
rect 1444 2135 1445 2139
rect 1439 2134 1445 2135
rect 1447 2139 1453 2140
rect 1447 2135 1448 2139
rect 1452 2138 1453 2139
rect 1487 2139 1493 2140
rect 1487 2138 1488 2139
rect 1452 2136 1488 2138
rect 1452 2135 1453 2136
rect 1447 2134 1453 2135
rect 1487 2135 1488 2136
rect 1492 2135 1493 2139
rect 1487 2134 1493 2135
rect 1495 2139 1501 2140
rect 1495 2135 1496 2139
rect 1500 2138 1501 2139
rect 1543 2139 1549 2140
rect 1543 2138 1544 2139
rect 1500 2136 1544 2138
rect 1500 2135 1501 2136
rect 1495 2134 1501 2135
rect 1543 2135 1544 2136
rect 1548 2135 1549 2139
rect 1543 2134 1549 2135
rect 1551 2139 1557 2140
rect 1551 2135 1552 2139
rect 1556 2138 1557 2139
rect 1599 2139 1605 2140
rect 1599 2138 1600 2139
rect 1556 2136 1600 2138
rect 1556 2135 1557 2136
rect 1551 2134 1557 2135
rect 1599 2135 1600 2136
rect 1604 2135 1605 2139
rect 1599 2134 1605 2135
rect 1646 2139 1653 2140
rect 1646 2135 1647 2139
rect 1652 2135 1653 2139
rect 1646 2134 1653 2135
rect 1655 2139 1661 2140
rect 1655 2135 1656 2139
rect 1660 2138 1661 2139
rect 1695 2139 1701 2140
rect 1695 2138 1696 2139
rect 1660 2136 1696 2138
rect 1660 2135 1661 2136
rect 1655 2134 1661 2135
rect 1695 2135 1696 2136
rect 1700 2135 1701 2139
rect 1695 2134 1701 2135
rect 1706 2139 1712 2140
rect 1706 2135 1707 2139
rect 1711 2138 1712 2139
rect 1743 2139 1749 2140
rect 1743 2138 1744 2139
rect 1711 2136 1744 2138
rect 1711 2135 1712 2136
rect 1706 2134 1712 2135
rect 1743 2135 1744 2136
rect 1748 2135 1749 2139
rect 1743 2134 1749 2135
rect 1754 2139 1760 2140
rect 1754 2135 1755 2139
rect 1759 2138 1760 2139
rect 1799 2139 1805 2140
rect 1799 2138 1800 2139
rect 1759 2136 1800 2138
rect 1759 2135 1760 2136
rect 1754 2134 1760 2135
rect 1799 2135 1800 2136
rect 1804 2135 1805 2139
rect 1799 2134 1805 2135
rect 1810 2139 1816 2140
rect 1810 2135 1811 2139
rect 1815 2138 1816 2139
rect 1855 2139 1861 2140
rect 1855 2138 1856 2139
rect 1815 2136 1856 2138
rect 1815 2135 1816 2136
rect 1810 2134 1816 2135
rect 1855 2135 1856 2136
rect 1860 2135 1861 2139
rect 1855 2134 1861 2135
rect 1863 2139 1869 2140
rect 1863 2135 1864 2139
rect 1868 2138 1869 2139
rect 1911 2139 1917 2140
rect 1911 2138 1912 2139
rect 1868 2136 1912 2138
rect 1868 2135 1869 2136
rect 1863 2134 1869 2135
rect 1911 2135 1912 2136
rect 1916 2135 1917 2139
rect 1911 2134 1917 2135
rect 2118 2136 2124 2137
rect 1134 2131 1140 2132
rect 2118 2132 2119 2136
rect 2123 2132 2124 2136
rect 2118 2131 2124 2132
rect 1286 2128 1292 2129
rect 1286 2124 1287 2128
rect 1291 2124 1292 2128
rect 1286 2123 1292 2124
rect 1326 2128 1332 2129
rect 1326 2124 1327 2128
rect 1331 2124 1332 2128
rect 1326 2123 1332 2124
rect 1366 2128 1372 2129
rect 1366 2124 1367 2128
rect 1371 2124 1372 2128
rect 1366 2123 1372 2124
rect 1414 2128 1420 2129
rect 1414 2124 1415 2128
rect 1419 2124 1420 2128
rect 1414 2123 1420 2124
rect 1462 2128 1468 2129
rect 1462 2124 1463 2128
rect 1467 2124 1468 2128
rect 1462 2123 1468 2124
rect 1518 2128 1524 2129
rect 1518 2124 1519 2128
rect 1523 2124 1524 2128
rect 1518 2123 1524 2124
rect 1574 2128 1580 2129
rect 1574 2124 1575 2128
rect 1579 2124 1580 2128
rect 1574 2123 1580 2124
rect 1622 2128 1628 2129
rect 1622 2124 1623 2128
rect 1627 2124 1628 2128
rect 1622 2123 1628 2124
rect 1670 2128 1676 2129
rect 1670 2124 1671 2128
rect 1675 2124 1676 2128
rect 1670 2123 1676 2124
rect 1718 2128 1724 2129
rect 1718 2124 1719 2128
rect 1723 2124 1724 2128
rect 1718 2123 1724 2124
rect 1774 2128 1780 2129
rect 1774 2124 1775 2128
rect 1779 2124 1780 2128
rect 1774 2123 1780 2124
rect 1830 2128 1836 2129
rect 1830 2124 1831 2128
rect 1835 2124 1836 2128
rect 1830 2123 1836 2124
rect 1886 2128 1892 2129
rect 1886 2124 1887 2128
rect 1891 2124 1892 2128
rect 1886 2123 1892 2124
rect 1311 2119 1317 2120
rect 1311 2115 1312 2119
rect 1316 2118 1317 2119
rect 1334 2119 1340 2120
rect 1334 2118 1335 2119
rect 1316 2116 1335 2118
rect 1316 2115 1317 2116
rect 1311 2114 1317 2115
rect 1334 2115 1335 2116
rect 1339 2115 1340 2119
rect 1334 2114 1340 2115
rect 1351 2119 1357 2120
rect 1351 2115 1352 2119
rect 1356 2118 1357 2119
rect 1374 2119 1380 2120
rect 1374 2118 1375 2119
rect 1356 2116 1375 2118
rect 1356 2115 1357 2116
rect 1351 2114 1357 2115
rect 1374 2115 1375 2116
rect 1379 2115 1380 2119
rect 1374 2114 1380 2115
rect 1391 2119 1397 2120
rect 1391 2115 1392 2119
rect 1396 2118 1397 2119
rect 1399 2119 1405 2120
rect 1399 2118 1400 2119
rect 1396 2116 1400 2118
rect 1396 2115 1397 2116
rect 1391 2114 1397 2115
rect 1399 2115 1400 2116
rect 1404 2115 1405 2119
rect 1399 2114 1405 2115
rect 1439 2119 1445 2120
rect 1439 2115 1440 2119
rect 1444 2118 1445 2119
rect 1447 2119 1453 2120
rect 1447 2118 1448 2119
rect 1444 2116 1448 2118
rect 1444 2115 1445 2116
rect 1439 2114 1445 2115
rect 1447 2115 1448 2116
rect 1452 2115 1453 2119
rect 1447 2114 1453 2115
rect 1487 2119 1493 2120
rect 1487 2115 1488 2119
rect 1492 2118 1493 2119
rect 1495 2119 1501 2120
rect 1495 2118 1496 2119
rect 1492 2116 1496 2118
rect 1492 2115 1493 2116
rect 1487 2114 1493 2115
rect 1495 2115 1496 2116
rect 1500 2115 1501 2119
rect 1495 2114 1501 2115
rect 1543 2119 1549 2120
rect 1543 2115 1544 2119
rect 1548 2118 1549 2119
rect 1551 2119 1557 2120
rect 1551 2118 1552 2119
rect 1548 2116 1552 2118
rect 1548 2115 1549 2116
rect 1543 2114 1549 2115
rect 1551 2115 1552 2116
rect 1556 2115 1557 2119
rect 1599 2119 1605 2120
rect 1599 2118 1600 2119
rect 1551 2114 1557 2115
rect 1560 2116 1600 2118
rect 1390 2111 1396 2112
rect 1390 2107 1391 2111
rect 1395 2110 1396 2111
rect 1560 2110 1562 2116
rect 1599 2115 1600 2116
rect 1604 2115 1605 2119
rect 1599 2114 1605 2115
rect 1647 2119 1653 2120
rect 1647 2115 1648 2119
rect 1652 2118 1653 2119
rect 1655 2119 1661 2120
rect 1655 2118 1656 2119
rect 1652 2116 1656 2118
rect 1652 2115 1653 2116
rect 1647 2114 1653 2115
rect 1655 2115 1656 2116
rect 1660 2115 1661 2119
rect 1655 2114 1661 2115
rect 1695 2119 1701 2120
rect 1695 2115 1696 2119
rect 1700 2118 1701 2119
rect 1706 2119 1712 2120
rect 1706 2118 1707 2119
rect 1700 2116 1707 2118
rect 1700 2115 1701 2116
rect 1695 2114 1701 2115
rect 1706 2115 1707 2116
rect 1711 2115 1712 2119
rect 1706 2114 1712 2115
rect 1743 2119 1749 2120
rect 1743 2115 1744 2119
rect 1748 2118 1749 2119
rect 1754 2119 1760 2120
rect 1754 2118 1755 2119
rect 1748 2116 1755 2118
rect 1748 2115 1749 2116
rect 1743 2114 1749 2115
rect 1754 2115 1755 2116
rect 1759 2115 1760 2119
rect 1754 2114 1760 2115
rect 1799 2119 1805 2120
rect 1799 2115 1800 2119
rect 1804 2118 1805 2119
rect 1810 2119 1816 2120
rect 1810 2118 1811 2119
rect 1804 2116 1811 2118
rect 1804 2115 1805 2116
rect 1799 2114 1805 2115
rect 1810 2115 1811 2116
rect 1815 2115 1816 2119
rect 1810 2114 1816 2115
rect 1855 2119 1861 2120
rect 1855 2115 1856 2119
rect 1860 2118 1861 2119
rect 1863 2119 1869 2120
rect 1863 2118 1864 2119
rect 1860 2116 1864 2118
rect 1860 2115 1861 2116
rect 1855 2114 1861 2115
rect 1863 2115 1864 2116
rect 1868 2115 1869 2119
rect 1911 2119 1917 2120
rect 1911 2118 1912 2119
rect 1863 2114 1869 2115
rect 1872 2116 1912 2118
rect 1395 2108 1562 2110
rect 1690 2111 1696 2112
rect 1395 2107 1396 2108
rect 1390 2106 1396 2107
rect 1690 2107 1691 2111
rect 1695 2110 1696 2111
rect 1872 2110 1874 2116
rect 1911 2115 1912 2116
rect 1916 2115 1917 2119
rect 1911 2114 1917 2115
rect 1695 2108 1874 2110
rect 1695 2107 1696 2108
rect 1690 2106 1696 2107
rect 1247 2095 1253 2096
rect 1247 2091 1248 2095
rect 1252 2094 1253 2095
rect 1294 2095 1300 2096
rect 1294 2094 1295 2095
rect 1252 2092 1295 2094
rect 1252 2091 1253 2092
rect 1247 2090 1253 2091
rect 1294 2091 1295 2092
rect 1299 2091 1300 2095
rect 1294 2090 1300 2091
rect 1303 2095 1309 2096
rect 1303 2091 1304 2095
rect 1308 2094 1309 2095
rect 1350 2095 1356 2096
rect 1350 2094 1351 2095
rect 1308 2092 1351 2094
rect 1308 2091 1309 2092
rect 1303 2090 1309 2091
rect 1350 2091 1351 2092
rect 1355 2091 1356 2095
rect 1350 2090 1356 2091
rect 1367 2095 1373 2096
rect 1367 2091 1368 2095
rect 1372 2094 1373 2095
rect 1438 2095 1444 2096
rect 1438 2094 1439 2095
rect 1372 2092 1439 2094
rect 1372 2091 1373 2092
rect 1367 2090 1373 2091
rect 1438 2091 1439 2092
rect 1443 2091 1444 2095
rect 1438 2090 1444 2091
rect 1447 2095 1453 2096
rect 1447 2091 1448 2095
rect 1452 2094 1453 2095
rect 1518 2095 1524 2096
rect 1518 2094 1519 2095
rect 1452 2092 1519 2094
rect 1452 2091 1453 2092
rect 1447 2090 1453 2091
rect 1518 2091 1519 2092
rect 1523 2091 1524 2095
rect 1518 2090 1524 2091
rect 1527 2095 1533 2096
rect 1527 2091 1528 2095
rect 1532 2094 1533 2095
rect 1598 2095 1604 2096
rect 1598 2094 1599 2095
rect 1532 2092 1599 2094
rect 1532 2091 1533 2092
rect 1527 2090 1533 2091
rect 1598 2091 1599 2092
rect 1603 2091 1604 2095
rect 1598 2090 1604 2091
rect 1606 2095 1613 2096
rect 1606 2091 1607 2095
rect 1612 2091 1613 2095
rect 1606 2090 1613 2091
rect 1687 2095 1693 2096
rect 1687 2091 1688 2095
rect 1692 2094 1693 2095
rect 1758 2095 1764 2096
rect 1758 2094 1759 2095
rect 1692 2092 1759 2094
rect 1692 2091 1693 2092
rect 1687 2090 1693 2091
rect 1758 2091 1759 2092
rect 1763 2091 1764 2095
rect 1758 2090 1764 2091
rect 1767 2095 1773 2096
rect 1767 2091 1768 2095
rect 1772 2094 1773 2095
rect 1846 2095 1852 2096
rect 1846 2094 1847 2095
rect 1772 2092 1847 2094
rect 1772 2091 1773 2092
rect 1767 2090 1773 2091
rect 1846 2091 1847 2092
rect 1851 2091 1852 2095
rect 1846 2090 1852 2091
rect 1855 2095 1861 2096
rect 1855 2091 1856 2095
rect 1860 2094 1861 2095
rect 1934 2095 1940 2096
rect 1934 2094 1935 2095
rect 1860 2092 1935 2094
rect 1860 2091 1861 2092
rect 1855 2090 1861 2091
rect 1934 2091 1935 2092
rect 1939 2091 1940 2095
rect 1934 2090 1940 2091
rect 1943 2095 1949 2096
rect 1943 2091 1944 2095
rect 1948 2094 1949 2095
rect 2022 2095 2028 2096
rect 2022 2094 2023 2095
rect 1948 2092 2023 2094
rect 1948 2091 1949 2092
rect 1943 2090 1949 2091
rect 2022 2091 2023 2092
rect 2027 2091 2028 2095
rect 2022 2090 2028 2091
rect 2030 2095 2037 2096
rect 2030 2091 2031 2095
rect 2036 2091 2037 2095
rect 2030 2090 2037 2091
rect 1222 2088 1228 2089
rect 1222 2084 1223 2088
rect 1227 2084 1228 2088
rect 1222 2083 1228 2084
rect 1278 2088 1284 2089
rect 1278 2084 1279 2088
rect 1283 2084 1284 2088
rect 1278 2083 1284 2084
rect 1342 2088 1348 2089
rect 1342 2084 1343 2088
rect 1347 2084 1348 2088
rect 1342 2083 1348 2084
rect 1422 2088 1428 2089
rect 1422 2084 1423 2088
rect 1427 2084 1428 2088
rect 1422 2083 1428 2084
rect 1502 2088 1508 2089
rect 1502 2084 1503 2088
rect 1507 2084 1508 2088
rect 1502 2083 1508 2084
rect 1582 2088 1588 2089
rect 1582 2084 1583 2088
rect 1587 2084 1588 2088
rect 1582 2083 1588 2084
rect 1662 2088 1668 2089
rect 1662 2084 1663 2088
rect 1667 2084 1668 2088
rect 1662 2083 1668 2084
rect 1742 2088 1748 2089
rect 1742 2084 1743 2088
rect 1747 2084 1748 2088
rect 1742 2083 1748 2084
rect 1830 2088 1836 2089
rect 1830 2084 1831 2088
rect 1835 2084 1836 2088
rect 1830 2083 1836 2084
rect 1918 2088 1924 2089
rect 1918 2084 1919 2088
rect 1923 2084 1924 2088
rect 1918 2083 1924 2084
rect 2006 2088 2012 2089
rect 2006 2084 2007 2088
rect 2011 2084 2012 2088
rect 2006 2083 2012 2084
rect 2070 2088 2076 2089
rect 2070 2084 2071 2088
rect 2075 2084 2076 2088
rect 2070 2083 2076 2084
rect 1134 2080 1140 2081
rect 1134 2076 1135 2080
rect 1139 2076 1140 2080
rect 2118 2080 2124 2081
rect 2118 2076 2119 2080
rect 2123 2076 2124 2080
rect 1134 2075 1140 2076
rect 1210 2075 1216 2076
rect 1210 2071 1211 2075
rect 1215 2074 1216 2075
rect 1247 2075 1253 2076
rect 1247 2074 1248 2075
rect 1215 2072 1248 2074
rect 1215 2071 1216 2072
rect 1210 2070 1216 2071
rect 1247 2071 1248 2072
rect 1252 2071 1253 2075
rect 1247 2070 1253 2071
rect 1294 2075 1300 2076
rect 1294 2071 1295 2075
rect 1299 2074 1300 2075
rect 1303 2075 1309 2076
rect 1303 2074 1304 2075
rect 1299 2072 1304 2074
rect 1299 2071 1300 2072
rect 1294 2070 1300 2071
rect 1303 2071 1304 2072
rect 1308 2071 1309 2075
rect 1303 2070 1309 2071
rect 1350 2075 1356 2076
rect 1350 2071 1351 2075
rect 1355 2074 1356 2075
rect 1367 2075 1373 2076
rect 1367 2074 1368 2075
rect 1355 2072 1368 2074
rect 1355 2071 1356 2072
rect 1350 2070 1356 2071
rect 1367 2071 1368 2072
rect 1372 2071 1373 2075
rect 1367 2070 1373 2071
rect 1438 2075 1444 2076
rect 1438 2071 1439 2075
rect 1443 2074 1444 2075
rect 1447 2075 1453 2076
rect 1447 2074 1448 2075
rect 1443 2072 1448 2074
rect 1443 2071 1444 2072
rect 1438 2070 1444 2071
rect 1447 2071 1448 2072
rect 1452 2071 1453 2075
rect 1447 2070 1453 2071
rect 1518 2075 1524 2076
rect 1518 2071 1519 2075
rect 1523 2074 1524 2075
rect 1527 2075 1533 2076
rect 1527 2074 1528 2075
rect 1523 2072 1528 2074
rect 1523 2071 1524 2072
rect 1518 2070 1524 2071
rect 1527 2071 1528 2072
rect 1532 2071 1533 2075
rect 1527 2070 1533 2071
rect 1598 2075 1604 2076
rect 1598 2071 1599 2075
rect 1603 2074 1604 2075
rect 1607 2075 1613 2076
rect 1607 2074 1608 2075
rect 1603 2072 1608 2074
rect 1603 2071 1604 2072
rect 1598 2070 1604 2071
rect 1607 2071 1608 2072
rect 1612 2071 1613 2075
rect 1607 2070 1613 2071
rect 1687 2075 1696 2076
rect 1687 2071 1688 2075
rect 1695 2071 1696 2075
rect 1687 2070 1696 2071
rect 1758 2075 1764 2076
rect 1758 2071 1759 2075
rect 1763 2074 1764 2075
rect 1767 2075 1773 2076
rect 1767 2074 1768 2075
rect 1763 2072 1768 2074
rect 1763 2071 1764 2072
rect 1758 2070 1764 2071
rect 1767 2071 1768 2072
rect 1772 2071 1773 2075
rect 1767 2070 1773 2071
rect 1846 2075 1852 2076
rect 1846 2071 1847 2075
rect 1851 2074 1852 2075
rect 1855 2075 1861 2076
rect 1855 2074 1856 2075
rect 1851 2072 1856 2074
rect 1851 2071 1852 2072
rect 1846 2070 1852 2071
rect 1855 2071 1856 2072
rect 1860 2071 1861 2075
rect 1855 2070 1861 2071
rect 1934 2075 1940 2076
rect 1934 2071 1935 2075
rect 1939 2074 1940 2075
rect 1943 2075 1949 2076
rect 1943 2074 1944 2075
rect 1939 2072 1944 2074
rect 1939 2071 1940 2072
rect 1934 2070 1940 2071
rect 1943 2071 1944 2072
rect 1948 2071 1949 2075
rect 1943 2070 1949 2071
rect 2022 2075 2028 2076
rect 2022 2071 2023 2075
rect 2027 2074 2028 2075
rect 2031 2075 2037 2076
rect 2031 2074 2032 2075
rect 2027 2072 2032 2074
rect 2027 2071 2028 2072
rect 2022 2070 2028 2071
rect 2031 2071 2032 2072
rect 2036 2071 2037 2075
rect 2031 2070 2037 2071
rect 2094 2075 2101 2076
rect 2118 2075 2124 2076
rect 2094 2071 2095 2075
rect 2100 2071 2101 2075
rect 2094 2070 2101 2071
rect 1134 2063 1140 2064
rect 1134 2059 1135 2063
rect 1139 2059 1140 2063
rect 2118 2063 2124 2064
rect 1134 2058 1140 2059
rect 1222 2060 1228 2061
rect 1222 2056 1223 2060
rect 1227 2056 1228 2060
rect 1222 2055 1228 2056
rect 1278 2060 1284 2061
rect 1278 2056 1279 2060
rect 1283 2056 1284 2060
rect 1278 2055 1284 2056
rect 1342 2060 1348 2061
rect 1342 2056 1343 2060
rect 1347 2056 1348 2060
rect 1342 2055 1348 2056
rect 1422 2060 1428 2061
rect 1422 2056 1423 2060
rect 1427 2056 1428 2060
rect 1422 2055 1428 2056
rect 1502 2060 1508 2061
rect 1502 2056 1503 2060
rect 1507 2056 1508 2060
rect 1502 2055 1508 2056
rect 1582 2060 1588 2061
rect 1582 2056 1583 2060
rect 1587 2056 1588 2060
rect 1582 2055 1588 2056
rect 1662 2060 1668 2061
rect 1662 2056 1663 2060
rect 1667 2056 1668 2060
rect 1662 2055 1668 2056
rect 1742 2060 1748 2061
rect 1742 2056 1743 2060
rect 1747 2056 1748 2060
rect 1742 2055 1748 2056
rect 1830 2060 1836 2061
rect 1830 2056 1831 2060
rect 1835 2056 1836 2060
rect 1830 2055 1836 2056
rect 1918 2060 1924 2061
rect 1918 2056 1919 2060
rect 1923 2056 1924 2060
rect 1918 2055 1924 2056
rect 2006 2060 2012 2061
rect 2006 2056 2007 2060
rect 2011 2056 2012 2060
rect 2006 2055 2012 2056
rect 2070 2060 2076 2061
rect 2070 2056 2071 2060
rect 2075 2056 2076 2060
rect 2118 2059 2119 2063
rect 2123 2059 2124 2063
rect 2118 2058 2124 2059
rect 2070 2055 2076 2056
rect 1182 2048 1188 2049
rect 1134 2045 1140 2046
rect 1134 2041 1135 2045
rect 1139 2041 1140 2045
rect 1182 2044 1183 2048
rect 1187 2044 1188 2048
rect 1182 2043 1188 2044
rect 1238 2048 1244 2049
rect 1238 2044 1239 2048
rect 1243 2044 1244 2048
rect 1238 2043 1244 2044
rect 1310 2048 1316 2049
rect 1310 2044 1311 2048
rect 1315 2044 1316 2048
rect 1310 2043 1316 2044
rect 1398 2048 1404 2049
rect 1398 2044 1399 2048
rect 1403 2044 1404 2048
rect 1398 2043 1404 2044
rect 1486 2048 1492 2049
rect 1486 2044 1487 2048
rect 1491 2044 1492 2048
rect 1486 2043 1492 2044
rect 1582 2048 1588 2049
rect 1582 2044 1583 2048
rect 1587 2044 1588 2048
rect 1582 2043 1588 2044
rect 1670 2048 1676 2049
rect 1670 2044 1671 2048
rect 1675 2044 1676 2048
rect 1670 2043 1676 2044
rect 1758 2048 1764 2049
rect 1758 2044 1759 2048
rect 1763 2044 1764 2048
rect 1758 2043 1764 2044
rect 1838 2048 1844 2049
rect 1838 2044 1839 2048
rect 1843 2044 1844 2048
rect 1838 2043 1844 2044
rect 1918 2048 1924 2049
rect 1918 2044 1919 2048
rect 1923 2044 1924 2048
rect 1918 2043 1924 2044
rect 2006 2048 2012 2049
rect 2006 2044 2007 2048
rect 2011 2044 2012 2048
rect 2006 2043 2012 2044
rect 2070 2048 2076 2049
rect 2070 2044 2071 2048
rect 2075 2044 2076 2048
rect 2070 2043 2076 2044
rect 2118 2045 2124 2046
rect 1134 2040 1140 2041
rect 2118 2041 2119 2045
rect 2123 2041 2124 2045
rect 2118 2040 2124 2041
rect 1862 2039 1868 2040
rect 1862 2038 1863 2039
rect 1696 2036 1863 2038
rect 1696 2032 1698 2036
rect 1862 2035 1863 2036
rect 1867 2035 1868 2039
rect 1862 2034 1868 2035
rect 1207 2031 1213 2032
rect 1134 2028 1140 2029
rect 1134 2024 1135 2028
rect 1139 2024 1140 2028
rect 1207 2027 1208 2031
rect 1212 2030 1213 2031
rect 1254 2031 1260 2032
rect 1254 2030 1255 2031
rect 1212 2028 1255 2030
rect 1212 2027 1213 2028
rect 1207 2026 1213 2027
rect 1254 2027 1255 2028
rect 1259 2027 1260 2031
rect 1254 2026 1260 2027
rect 1263 2031 1269 2032
rect 1263 2027 1264 2031
rect 1268 2030 1269 2031
rect 1326 2031 1332 2032
rect 1326 2030 1327 2031
rect 1268 2028 1327 2030
rect 1268 2027 1269 2028
rect 1263 2026 1269 2027
rect 1326 2027 1327 2028
rect 1331 2027 1332 2031
rect 1326 2026 1332 2027
rect 1335 2031 1341 2032
rect 1335 2027 1336 2031
rect 1340 2030 1341 2031
rect 1414 2031 1420 2032
rect 1414 2030 1415 2031
rect 1340 2028 1415 2030
rect 1340 2027 1341 2028
rect 1335 2026 1341 2027
rect 1414 2027 1415 2028
rect 1419 2027 1420 2031
rect 1414 2026 1420 2027
rect 1423 2031 1429 2032
rect 1423 2027 1424 2031
rect 1428 2030 1429 2031
rect 1502 2031 1508 2032
rect 1502 2030 1503 2031
rect 1428 2028 1503 2030
rect 1428 2027 1429 2028
rect 1423 2026 1429 2027
rect 1502 2027 1503 2028
rect 1507 2027 1508 2031
rect 1502 2026 1508 2027
rect 1511 2031 1517 2032
rect 1511 2027 1512 2031
rect 1516 2030 1517 2031
rect 1558 2031 1564 2032
rect 1558 2030 1559 2031
rect 1516 2028 1559 2030
rect 1516 2027 1517 2028
rect 1511 2026 1517 2027
rect 1558 2027 1559 2028
rect 1563 2027 1564 2031
rect 1558 2026 1564 2027
rect 1570 2031 1576 2032
rect 1570 2027 1571 2031
rect 1575 2030 1576 2031
rect 1607 2031 1613 2032
rect 1607 2030 1608 2031
rect 1575 2028 1608 2030
rect 1575 2027 1576 2028
rect 1570 2026 1576 2027
rect 1607 2027 1608 2028
rect 1612 2027 1613 2031
rect 1607 2026 1613 2027
rect 1695 2031 1701 2032
rect 1695 2027 1696 2031
rect 1700 2027 1701 2031
rect 1695 2026 1701 2027
rect 1703 2031 1709 2032
rect 1703 2027 1704 2031
rect 1708 2030 1709 2031
rect 1783 2031 1789 2032
rect 1783 2030 1784 2031
rect 1708 2028 1784 2030
rect 1708 2027 1709 2028
rect 1703 2026 1709 2027
rect 1783 2027 1784 2028
rect 1788 2027 1789 2031
rect 1783 2026 1789 2027
rect 1863 2031 1869 2032
rect 1863 2027 1864 2031
rect 1868 2030 1869 2031
rect 1934 2031 1940 2032
rect 1934 2030 1935 2031
rect 1868 2028 1935 2030
rect 1868 2027 1869 2028
rect 1863 2026 1869 2027
rect 1934 2027 1935 2028
rect 1939 2027 1940 2031
rect 1934 2026 1940 2027
rect 1943 2031 1949 2032
rect 1943 2027 1944 2031
rect 1948 2030 1949 2031
rect 2022 2031 2028 2032
rect 2022 2030 2023 2031
rect 1948 2028 2023 2030
rect 1948 2027 1949 2028
rect 1943 2026 1949 2027
rect 2022 2027 2023 2028
rect 2027 2027 2028 2031
rect 2022 2026 2028 2027
rect 2030 2031 2037 2032
rect 2030 2027 2031 2031
rect 2036 2027 2037 2031
rect 2030 2026 2037 2027
rect 2095 2031 2101 2032
rect 2095 2027 2096 2031
rect 2100 2030 2101 2031
rect 2103 2031 2109 2032
rect 2103 2030 2104 2031
rect 2100 2028 2104 2030
rect 2100 2027 2101 2028
rect 2095 2026 2101 2027
rect 2103 2027 2104 2028
rect 2108 2027 2109 2031
rect 2103 2026 2109 2027
rect 2118 2028 2124 2029
rect 215 2023 221 2024
rect 215 2019 216 2023
rect 220 2022 221 2023
rect 246 2023 252 2024
rect 246 2022 247 2023
rect 220 2020 247 2022
rect 220 2019 221 2020
rect 215 2018 221 2019
rect 246 2019 247 2020
rect 251 2019 252 2023
rect 246 2018 252 2019
rect 255 2023 261 2024
rect 255 2019 256 2023
rect 260 2022 261 2023
rect 302 2023 308 2024
rect 302 2022 303 2023
rect 260 2020 303 2022
rect 260 2019 261 2020
rect 255 2018 261 2019
rect 302 2019 303 2020
rect 307 2019 308 2023
rect 302 2018 308 2019
rect 311 2023 317 2024
rect 311 2019 312 2023
rect 316 2022 317 2023
rect 366 2023 372 2024
rect 366 2022 367 2023
rect 316 2020 367 2022
rect 316 2019 317 2020
rect 311 2018 317 2019
rect 366 2019 367 2020
rect 371 2019 372 2023
rect 366 2018 372 2019
rect 375 2023 381 2024
rect 375 2019 376 2023
rect 380 2022 381 2023
rect 438 2023 444 2024
rect 438 2022 439 2023
rect 380 2020 439 2022
rect 380 2019 381 2020
rect 375 2018 381 2019
rect 438 2019 439 2020
rect 443 2019 444 2023
rect 438 2018 444 2019
rect 447 2023 453 2024
rect 447 2019 448 2023
rect 452 2022 453 2023
rect 510 2023 516 2024
rect 510 2022 511 2023
rect 452 2020 511 2022
rect 452 2019 453 2020
rect 447 2018 453 2019
rect 510 2019 511 2020
rect 515 2019 516 2023
rect 510 2018 516 2019
rect 519 2023 525 2024
rect 519 2019 520 2023
rect 524 2022 525 2023
rect 538 2023 544 2024
rect 538 2022 539 2023
rect 524 2020 539 2022
rect 524 2019 525 2020
rect 519 2018 525 2019
rect 538 2019 539 2020
rect 543 2019 544 2023
rect 538 2018 544 2019
rect 546 2023 552 2024
rect 546 2019 547 2023
rect 551 2022 552 2023
rect 599 2023 605 2024
rect 599 2022 600 2023
rect 551 2020 600 2022
rect 551 2019 552 2020
rect 546 2018 552 2019
rect 599 2019 600 2020
rect 604 2019 605 2023
rect 599 2018 605 2019
rect 671 2023 677 2024
rect 671 2019 672 2023
rect 676 2022 677 2023
rect 734 2023 740 2024
rect 734 2022 735 2023
rect 676 2020 735 2022
rect 676 2019 677 2020
rect 671 2018 677 2019
rect 734 2019 735 2020
rect 739 2019 740 2023
rect 734 2018 740 2019
rect 743 2023 749 2024
rect 743 2019 744 2023
rect 748 2022 749 2023
rect 790 2023 796 2024
rect 790 2022 791 2023
rect 748 2020 791 2022
rect 748 2019 749 2020
rect 743 2018 749 2019
rect 790 2019 791 2020
rect 795 2019 796 2023
rect 790 2018 796 2019
rect 807 2023 813 2024
rect 807 2019 808 2023
rect 812 2022 813 2023
rect 854 2023 860 2024
rect 854 2022 855 2023
rect 812 2020 855 2022
rect 812 2019 813 2020
rect 807 2018 813 2019
rect 854 2019 855 2020
rect 859 2019 860 2023
rect 854 2018 860 2019
rect 863 2023 869 2024
rect 863 2019 864 2023
rect 868 2022 869 2023
rect 910 2023 916 2024
rect 910 2022 911 2023
rect 868 2020 911 2022
rect 868 2019 869 2020
rect 863 2018 869 2019
rect 910 2019 911 2020
rect 915 2019 916 2023
rect 910 2018 916 2019
rect 919 2023 925 2024
rect 919 2019 920 2023
rect 924 2022 925 2023
rect 966 2023 972 2024
rect 966 2022 967 2023
rect 924 2020 967 2022
rect 924 2019 925 2020
rect 919 2018 925 2019
rect 966 2019 967 2020
rect 971 2019 972 2023
rect 966 2018 972 2019
rect 975 2023 981 2024
rect 975 2019 976 2023
rect 980 2022 981 2023
rect 1022 2023 1028 2024
rect 1022 2022 1023 2023
rect 980 2020 1023 2022
rect 980 2019 981 2020
rect 975 2018 981 2019
rect 1022 2019 1023 2020
rect 1027 2019 1028 2023
rect 1022 2018 1028 2019
rect 1031 2023 1037 2024
rect 1031 2019 1032 2023
rect 1036 2022 1037 2023
rect 1062 2023 1068 2024
rect 1062 2022 1063 2023
rect 1036 2020 1063 2022
rect 1036 2019 1037 2020
rect 1031 2018 1037 2019
rect 1062 2019 1063 2020
rect 1067 2019 1068 2023
rect 1062 2018 1068 2019
rect 1070 2023 1077 2024
rect 1134 2023 1140 2024
rect 2118 2024 2119 2028
rect 2123 2024 2124 2028
rect 2118 2023 2124 2024
rect 1070 2019 1071 2023
rect 1076 2019 1077 2023
rect 1070 2018 1077 2019
rect 1182 2020 1188 2021
rect 190 2016 196 2017
rect 190 2012 191 2016
rect 195 2012 196 2016
rect 190 2011 196 2012
rect 230 2016 236 2017
rect 230 2012 231 2016
rect 235 2012 236 2016
rect 230 2011 236 2012
rect 286 2016 292 2017
rect 286 2012 287 2016
rect 291 2012 292 2016
rect 286 2011 292 2012
rect 350 2016 356 2017
rect 350 2012 351 2016
rect 355 2012 356 2016
rect 350 2011 356 2012
rect 422 2016 428 2017
rect 422 2012 423 2016
rect 427 2012 428 2016
rect 422 2011 428 2012
rect 494 2016 500 2017
rect 494 2012 495 2016
rect 499 2012 500 2016
rect 494 2011 500 2012
rect 574 2016 580 2017
rect 574 2012 575 2016
rect 579 2012 580 2016
rect 574 2011 580 2012
rect 646 2016 652 2017
rect 646 2012 647 2016
rect 651 2012 652 2016
rect 646 2011 652 2012
rect 718 2016 724 2017
rect 718 2012 719 2016
rect 723 2012 724 2016
rect 718 2011 724 2012
rect 782 2016 788 2017
rect 782 2012 783 2016
rect 787 2012 788 2016
rect 782 2011 788 2012
rect 838 2016 844 2017
rect 838 2012 839 2016
rect 843 2012 844 2016
rect 838 2011 844 2012
rect 894 2016 900 2017
rect 894 2012 895 2016
rect 899 2012 900 2016
rect 894 2011 900 2012
rect 950 2016 956 2017
rect 950 2012 951 2016
rect 955 2012 956 2016
rect 950 2011 956 2012
rect 1006 2016 1012 2017
rect 1006 2012 1007 2016
rect 1011 2012 1012 2016
rect 1006 2011 1012 2012
rect 1046 2016 1052 2017
rect 1046 2012 1047 2016
rect 1051 2012 1052 2016
rect 1182 2016 1183 2020
rect 1187 2016 1188 2020
rect 1182 2015 1188 2016
rect 1238 2020 1244 2021
rect 1238 2016 1239 2020
rect 1243 2016 1244 2020
rect 1238 2015 1244 2016
rect 1310 2020 1316 2021
rect 1310 2016 1311 2020
rect 1315 2016 1316 2020
rect 1310 2015 1316 2016
rect 1398 2020 1404 2021
rect 1398 2016 1399 2020
rect 1403 2016 1404 2020
rect 1398 2015 1404 2016
rect 1486 2020 1492 2021
rect 1486 2016 1487 2020
rect 1491 2016 1492 2020
rect 1486 2015 1492 2016
rect 1582 2020 1588 2021
rect 1582 2016 1583 2020
rect 1587 2016 1588 2020
rect 1582 2015 1588 2016
rect 1670 2020 1676 2021
rect 1670 2016 1671 2020
rect 1675 2016 1676 2020
rect 1670 2015 1676 2016
rect 1758 2020 1764 2021
rect 1758 2016 1759 2020
rect 1763 2016 1764 2020
rect 1758 2015 1764 2016
rect 1838 2020 1844 2021
rect 1838 2016 1839 2020
rect 1843 2016 1844 2020
rect 1838 2015 1844 2016
rect 1918 2020 1924 2021
rect 1918 2016 1919 2020
rect 1923 2016 1924 2020
rect 1918 2015 1924 2016
rect 2006 2020 2012 2021
rect 2006 2016 2007 2020
rect 2011 2016 2012 2020
rect 2006 2015 2012 2016
rect 2070 2020 2076 2021
rect 2070 2016 2071 2020
rect 2075 2016 2076 2020
rect 2070 2015 2076 2016
rect 1046 2011 1052 2012
rect 1207 2011 1216 2012
rect 110 2008 116 2009
rect 110 2004 111 2008
rect 115 2004 116 2008
rect 1094 2008 1100 2009
rect 1094 2004 1095 2008
rect 1099 2004 1100 2008
rect 1207 2007 1208 2011
rect 1215 2007 1216 2011
rect 1207 2006 1216 2007
rect 1254 2011 1260 2012
rect 1254 2007 1255 2011
rect 1259 2010 1260 2011
rect 1263 2011 1269 2012
rect 1263 2010 1264 2011
rect 1259 2008 1264 2010
rect 1259 2007 1260 2008
rect 1254 2006 1260 2007
rect 1263 2007 1264 2008
rect 1268 2007 1269 2011
rect 1263 2006 1269 2007
rect 1326 2011 1332 2012
rect 1326 2007 1327 2011
rect 1331 2010 1332 2011
rect 1335 2011 1341 2012
rect 1335 2010 1336 2011
rect 1331 2008 1336 2010
rect 1331 2007 1332 2008
rect 1326 2006 1332 2007
rect 1335 2007 1336 2008
rect 1340 2007 1341 2011
rect 1335 2006 1341 2007
rect 1414 2011 1420 2012
rect 1414 2007 1415 2011
rect 1419 2010 1420 2011
rect 1423 2011 1429 2012
rect 1423 2010 1424 2011
rect 1419 2008 1424 2010
rect 1419 2007 1420 2008
rect 1414 2006 1420 2007
rect 1423 2007 1424 2008
rect 1428 2007 1429 2011
rect 1423 2006 1429 2007
rect 1502 2011 1508 2012
rect 1502 2007 1503 2011
rect 1507 2010 1508 2011
rect 1511 2011 1517 2012
rect 1511 2010 1512 2011
rect 1507 2008 1512 2010
rect 1507 2007 1508 2008
rect 1502 2006 1508 2007
rect 1511 2007 1512 2008
rect 1516 2007 1517 2011
rect 1511 2006 1517 2007
rect 1558 2011 1564 2012
rect 1558 2007 1559 2011
rect 1563 2010 1564 2011
rect 1607 2011 1613 2012
rect 1607 2010 1608 2011
rect 1563 2008 1608 2010
rect 1563 2007 1564 2008
rect 1558 2006 1564 2007
rect 1607 2007 1608 2008
rect 1612 2007 1613 2011
rect 1607 2006 1613 2007
rect 1695 2011 1701 2012
rect 1695 2007 1696 2011
rect 1700 2010 1701 2011
rect 1703 2011 1709 2012
rect 1703 2010 1704 2011
rect 1700 2008 1704 2010
rect 1700 2007 1701 2008
rect 1695 2006 1701 2007
rect 1703 2007 1704 2008
rect 1708 2007 1709 2011
rect 1703 2006 1709 2007
rect 1783 2011 1789 2012
rect 1783 2007 1784 2011
rect 1788 2010 1789 2011
rect 1830 2011 1836 2012
rect 1830 2010 1831 2011
rect 1788 2008 1831 2010
rect 1788 2007 1789 2008
rect 1783 2006 1789 2007
rect 1830 2007 1831 2008
rect 1835 2007 1836 2011
rect 1830 2006 1836 2007
rect 1862 2011 1869 2012
rect 1862 2007 1863 2011
rect 1868 2007 1869 2011
rect 1862 2006 1869 2007
rect 1934 2011 1940 2012
rect 1934 2007 1935 2011
rect 1939 2010 1940 2011
rect 1943 2011 1949 2012
rect 1943 2010 1944 2011
rect 1939 2008 1944 2010
rect 1939 2007 1940 2008
rect 1934 2006 1940 2007
rect 1943 2007 1944 2008
rect 1948 2007 1949 2011
rect 1943 2006 1949 2007
rect 2022 2011 2028 2012
rect 2022 2007 2023 2011
rect 2027 2010 2028 2011
rect 2031 2011 2037 2012
rect 2031 2010 2032 2011
rect 2027 2008 2032 2010
rect 2027 2007 2028 2008
rect 2022 2006 2028 2007
rect 2031 2007 2032 2008
rect 2036 2007 2037 2011
rect 2031 2006 2037 2007
rect 2094 2011 2101 2012
rect 2094 2007 2095 2011
rect 2100 2007 2101 2011
rect 2094 2006 2101 2007
rect 110 2003 116 2004
rect 214 2003 221 2004
rect 214 1999 215 2003
rect 220 1999 221 2003
rect 214 1998 221 1999
rect 246 2003 252 2004
rect 246 1999 247 2003
rect 251 2002 252 2003
rect 255 2003 261 2004
rect 255 2002 256 2003
rect 251 2000 256 2002
rect 251 1999 252 2000
rect 246 1998 252 1999
rect 255 1999 256 2000
rect 260 1999 261 2003
rect 255 1998 261 1999
rect 302 2003 308 2004
rect 302 1999 303 2003
rect 307 2002 308 2003
rect 311 2003 317 2004
rect 311 2002 312 2003
rect 307 2000 312 2002
rect 307 1999 308 2000
rect 302 1998 308 1999
rect 311 1999 312 2000
rect 316 1999 317 2003
rect 311 1998 317 1999
rect 366 2003 372 2004
rect 366 1999 367 2003
rect 371 2002 372 2003
rect 375 2003 381 2004
rect 375 2002 376 2003
rect 371 2000 376 2002
rect 371 1999 372 2000
rect 366 1998 372 1999
rect 375 1999 376 2000
rect 380 1999 381 2003
rect 375 1998 381 1999
rect 438 2003 444 2004
rect 438 1999 439 2003
rect 443 2002 444 2003
rect 447 2003 453 2004
rect 447 2002 448 2003
rect 443 2000 448 2002
rect 443 1999 444 2000
rect 438 1998 444 1999
rect 447 1999 448 2000
rect 452 1999 453 2003
rect 447 1998 453 1999
rect 510 2003 516 2004
rect 510 1999 511 2003
rect 515 2002 516 2003
rect 519 2003 525 2004
rect 519 2002 520 2003
rect 515 2000 520 2002
rect 515 1999 516 2000
rect 510 1998 516 1999
rect 519 1999 520 2000
rect 524 1999 525 2003
rect 519 1998 525 1999
rect 538 2003 544 2004
rect 538 1999 539 2003
rect 543 2002 544 2003
rect 599 2003 605 2004
rect 599 2002 600 2003
rect 543 2000 600 2002
rect 543 1999 544 2000
rect 538 1998 544 1999
rect 599 1999 600 2000
rect 604 1999 605 2003
rect 599 1998 605 1999
rect 671 2003 677 2004
rect 671 1999 672 2003
rect 676 2002 677 2003
rect 711 2003 717 2004
rect 711 2002 712 2003
rect 676 2000 712 2002
rect 676 1999 677 2000
rect 671 1998 677 1999
rect 711 1999 712 2000
rect 716 1999 717 2003
rect 711 1998 717 1999
rect 734 2003 740 2004
rect 734 1999 735 2003
rect 739 2002 740 2003
rect 743 2003 749 2004
rect 743 2002 744 2003
rect 739 2000 744 2002
rect 739 1999 740 2000
rect 734 1998 740 1999
rect 743 1999 744 2000
rect 748 1999 749 2003
rect 743 1998 749 1999
rect 790 2003 796 2004
rect 790 1999 791 2003
rect 795 2002 796 2003
rect 807 2003 813 2004
rect 807 2002 808 2003
rect 795 2000 808 2002
rect 795 1999 796 2000
rect 790 1998 796 1999
rect 807 1999 808 2000
rect 812 1999 813 2003
rect 807 1998 813 1999
rect 854 2003 860 2004
rect 854 1999 855 2003
rect 859 2002 860 2003
rect 863 2003 869 2004
rect 863 2002 864 2003
rect 859 2000 864 2002
rect 859 1999 860 2000
rect 854 1998 860 1999
rect 863 1999 864 2000
rect 868 1999 869 2003
rect 863 1998 869 1999
rect 910 2003 916 2004
rect 910 1999 911 2003
rect 915 2002 916 2003
rect 919 2003 925 2004
rect 919 2002 920 2003
rect 915 2000 920 2002
rect 915 1999 916 2000
rect 910 1998 916 1999
rect 919 1999 920 2000
rect 924 1999 925 2003
rect 919 1998 925 1999
rect 966 2003 972 2004
rect 966 1999 967 2003
rect 971 2002 972 2003
rect 975 2003 981 2004
rect 975 2002 976 2003
rect 971 2000 976 2002
rect 971 1999 972 2000
rect 966 1998 972 1999
rect 975 1999 976 2000
rect 980 1999 981 2003
rect 975 1998 981 1999
rect 1022 2003 1028 2004
rect 1022 1999 1023 2003
rect 1027 2002 1028 2003
rect 1031 2003 1037 2004
rect 1031 2002 1032 2003
rect 1027 2000 1032 2002
rect 1027 1999 1028 2000
rect 1022 1998 1028 1999
rect 1031 1999 1032 2000
rect 1036 1999 1037 2003
rect 1031 1998 1037 1999
rect 1062 2003 1068 2004
rect 1062 1999 1063 2003
rect 1067 2002 1068 2003
rect 1071 2003 1077 2004
rect 1094 2003 1100 2004
rect 1071 2002 1072 2003
rect 1067 2000 1072 2002
rect 1067 1999 1068 2000
rect 1062 1998 1068 1999
rect 1071 1999 1072 2000
rect 1076 1999 1077 2003
rect 1071 1998 1077 1999
rect 110 1991 116 1992
rect 110 1987 111 1991
rect 115 1987 116 1991
rect 1094 1991 1100 1992
rect 110 1986 116 1987
rect 190 1988 196 1989
rect 190 1984 191 1988
rect 195 1984 196 1988
rect 190 1983 196 1984
rect 230 1988 236 1989
rect 230 1984 231 1988
rect 235 1984 236 1988
rect 230 1983 236 1984
rect 286 1988 292 1989
rect 286 1984 287 1988
rect 291 1984 292 1988
rect 286 1983 292 1984
rect 350 1988 356 1989
rect 350 1984 351 1988
rect 355 1984 356 1988
rect 350 1983 356 1984
rect 422 1988 428 1989
rect 422 1984 423 1988
rect 427 1984 428 1988
rect 422 1983 428 1984
rect 494 1988 500 1989
rect 494 1984 495 1988
rect 499 1984 500 1988
rect 494 1983 500 1984
rect 574 1988 580 1989
rect 574 1984 575 1988
rect 579 1984 580 1988
rect 574 1983 580 1984
rect 646 1988 652 1989
rect 646 1984 647 1988
rect 651 1984 652 1988
rect 646 1983 652 1984
rect 718 1988 724 1989
rect 718 1984 719 1988
rect 723 1984 724 1988
rect 718 1983 724 1984
rect 782 1988 788 1989
rect 782 1984 783 1988
rect 787 1984 788 1988
rect 782 1983 788 1984
rect 838 1988 844 1989
rect 838 1984 839 1988
rect 843 1984 844 1988
rect 838 1983 844 1984
rect 894 1988 900 1989
rect 894 1984 895 1988
rect 899 1984 900 1988
rect 894 1983 900 1984
rect 950 1988 956 1989
rect 950 1984 951 1988
rect 955 1984 956 1988
rect 950 1983 956 1984
rect 1006 1988 1012 1989
rect 1006 1984 1007 1988
rect 1011 1984 1012 1988
rect 1006 1983 1012 1984
rect 1046 1988 1052 1989
rect 1046 1984 1047 1988
rect 1051 1984 1052 1988
rect 1094 1987 1095 1991
rect 1099 1987 1100 1991
rect 1094 1986 1100 1987
rect 1327 1991 1333 1992
rect 1327 1987 1328 1991
rect 1332 1990 1333 1991
rect 1398 1991 1404 1992
rect 1398 1990 1399 1991
rect 1332 1988 1399 1990
rect 1332 1987 1333 1988
rect 1327 1986 1333 1987
rect 1398 1987 1399 1988
rect 1403 1987 1404 1991
rect 1398 1986 1404 1987
rect 1407 1991 1413 1992
rect 1407 1987 1408 1991
rect 1412 1990 1413 1991
rect 1478 1991 1484 1992
rect 1478 1990 1479 1991
rect 1412 1988 1479 1990
rect 1412 1987 1413 1988
rect 1407 1986 1413 1987
rect 1478 1987 1479 1988
rect 1483 1987 1484 1991
rect 1478 1986 1484 1987
rect 1487 1991 1493 1992
rect 1487 1987 1488 1991
rect 1492 1990 1493 1991
rect 1550 1991 1556 1992
rect 1550 1990 1551 1991
rect 1492 1988 1551 1990
rect 1492 1987 1493 1988
rect 1487 1986 1493 1987
rect 1550 1987 1551 1988
rect 1555 1987 1556 1991
rect 1550 1986 1556 1987
rect 1567 1991 1576 1992
rect 1567 1987 1568 1991
rect 1575 1987 1576 1991
rect 1567 1986 1576 1987
rect 1639 1991 1645 1992
rect 1639 1987 1640 1991
rect 1644 1990 1645 1991
rect 1694 1991 1700 1992
rect 1694 1990 1695 1991
rect 1644 1988 1695 1990
rect 1644 1987 1645 1988
rect 1639 1986 1645 1987
rect 1694 1987 1695 1988
rect 1699 1987 1700 1991
rect 1694 1986 1700 1987
rect 1711 1991 1717 1992
rect 1711 1987 1712 1991
rect 1716 1990 1717 1991
rect 1766 1991 1772 1992
rect 1766 1990 1767 1991
rect 1716 1988 1767 1990
rect 1716 1987 1717 1988
rect 1711 1986 1717 1987
rect 1766 1987 1767 1988
rect 1771 1987 1772 1991
rect 1766 1986 1772 1987
rect 1775 1991 1781 1992
rect 1775 1987 1776 1991
rect 1780 1990 1781 1991
rect 1806 1991 1812 1992
rect 1806 1990 1807 1991
rect 1780 1988 1807 1990
rect 1780 1987 1781 1988
rect 1775 1986 1781 1987
rect 1806 1987 1807 1988
rect 1811 1987 1812 1991
rect 1806 1986 1812 1987
rect 1839 1991 1845 1992
rect 1839 1987 1840 1991
rect 1844 1990 1845 1991
rect 1894 1991 1900 1992
rect 1894 1990 1895 1991
rect 1844 1988 1895 1990
rect 1844 1987 1845 1988
rect 1839 1986 1845 1987
rect 1894 1987 1895 1988
rect 1899 1987 1900 1991
rect 1894 1986 1900 1987
rect 1903 1991 1909 1992
rect 1903 1987 1904 1991
rect 1908 1990 1909 1991
rect 1966 1991 1972 1992
rect 1966 1990 1967 1991
rect 1908 1988 1967 1990
rect 1908 1987 1909 1988
rect 1903 1986 1909 1987
rect 1966 1987 1967 1988
rect 1971 1987 1972 1991
rect 1966 1986 1972 1987
rect 1974 1991 1981 1992
rect 1974 1987 1975 1991
rect 1980 1987 1981 1991
rect 1974 1986 1981 1987
rect 2047 1991 2053 1992
rect 2047 1987 2048 1991
rect 2052 1990 2053 1991
rect 2086 1991 2092 1992
rect 2086 1990 2087 1991
rect 2052 1988 2087 1990
rect 2052 1987 2053 1988
rect 2047 1986 2053 1987
rect 2086 1987 2087 1988
rect 2091 1987 2092 1991
rect 2086 1986 2092 1987
rect 2095 1991 2101 1992
rect 2095 1987 2096 1991
rect 2100 1990 2101 1991
rect 2103 1991 2109 1992
rect 2103 1990 2104 1991
rect 2100 1988 2104 1990
rect 2100 1987 2101 1988
rect 2095 1986 2101 1987
rect 2103 1987 2104 1988
rect 2108 1987 2109 1991
rect 2103 1986 2109 1987
rect 1046 1983 1052 1984
rect 1302 1984 1308 1985
rect 1302 1980 1303 1984
rect 1307 1980 1308 1984
rect 1302 1979 1308 1980
rect 1382 1984 1388 1985
rect 1382 1980 1383 1984
rect 1387 1980 1388 1984
rect 1382 1979 1388 1980
rect 1462 1984 1468 1985
rect 1462 1980 1463 1984
rect 1467 1980 1468 1984
rect 1462 1979 1468 1980
rect 1542 1984 1548 1985
rect 1542 1980 1543 1984
rect 1547 1980 1548 1984
rect 1542 1979 1548 1980
rect 1614 1984 1620 1985
rect 1614 1980 1615 1984
rect 1619 1980 1620 1984
rect 1614 1979 1620 1980
rect 1686 1984 1692 1985
rect 1686 1980 1687 1984
rect 1691 1980 1692 1984
rect 1686 1979 1692 1980
rect 1750 1984 1756 1985
rect 1750 1980 1751 1984
rect 1755 1980 1756 1984
rect 1750 1979 1756 1980
rect 1814 1984 1820 1985
rect 1814 1980 1815 1984
rect 1819 1980 1820 1984
rect 1814 1979 1820 1980
rect 1878 1984 1884 1985
rect 1878 1980 1879 1984
rect 1883 1980 1884 1984
rect 1878 1979 1884 1980
rect 1950 1984 1956 1985
rect 1950 1980 1951 1984
rect 1955 1980 1956 1984
rect 1950 1979 1956 1980
rect 2022 1984 2028 1985
rect 2022 1980 2023 1984
rect 2027 1980 2028 1984
rect 2022 1979 2028 1980
rect 2070 1984 2076 1985
rect 2070 1980 2071 1984
rect 2075 1980 2076 1984
rect 2070 1979 2076 1980
rect 190 1976 196 1977
rect 110 1973 116 1974
rect 110 1969 111 1973
rect 115 1969 116 1973
rect 190 1972 191 1976
rect 195 1972 196 1976
rect 190 1971 196 1972
rect 246 1976 252 1977
rect 246 1972 247 1976
rect 251 1972 252 1976
rect 246 1971 252 1972
rect 310 1976 316 1977
rect 310 1972 311 1976
rect 315 1972 316 1976
rect 310 1971 316 1972
rect 374 1976 380 1977
rect 374 1972 375 1976
rect 379 1972 380 1976
rect 374 1971 380 1972
rect 446 1976 452 1977
rect 446 1972 447 1976
rect 451 1972 452 1976
rect 446 1971 452 1972
rect 518 1976 524 1977
rect 518 1972 519 1976
rect 523 1972 524 1976
rect 518 1971 524 1972
rect 590 1976 596 1977
rect 590 1972 591 1976
rect 595 1972 596 1976
rect 590 1971 596 1972
rect 654 1976 660 1977
rect 654 1972 655 1976
rect 659 1972 660 1976
rect 654 1971 660 1972
rect 718 1976 724 1977
rect 718 1972 719 1976
rect 723 1972 724 1976
rect 718 1971 724 1972
rect 774 1976 780 1977
rect 774 1972 775 1976
rect 779 1972 780 1976
rect 774 1971 780 1972
rect 822 1976 828 1977
rect 822 1972 823 1976
rect 827 1972 828 1976
rect 822 1971 828 1972
rect 870 1976 876 1977
rect 870 1972 871 1976
rect 875 1972 876 1976
rect 870 1971 876 1972
rect 918 1976 924 1977
rect 918 1972 919 1976
rect 923 1972 924 1976
rect 918 1971 924 1972
rect 966 1976 972 1977
rect 966 1972 967 1976
rect 971 1972 972 1976
rect 966 1971 972 1972
rect 1006 1976 1012 1977
rect 1006 1972 1007 1976
rect 1011 1972 1012 1976
rect 1006 1971 1012 1972
rect 1046 1976 1052 1977
rect 1046 1972 1047 1976
rect 1051 1972 1052 1976
rect 1134 1976 1140 1977
rect 1046 1971 1052 1972
rect 1094 1973 1100 1974
rect 110 1968 116 1969
rect 1094 1969 1095 1973
rect 1099 1969 1100 1973
rect 1134 1972 1135 1976
rect 1139 1972 1140 1976
rect 2118 1976 2124 1977
rect 2118 1972 2119 1976
rect 2123 1972 2124 1976
rect 1134 1971 1140 1972
rect 1326 1971 1333 1972
rect 1094 1968 1100 1969
rect 711 1967 717 1968
rect 711 1963 712 1967
rect 716 1966 717 1967
rect 894 1967 900 1968
rect 894 1966 895 1967
rect 716 1964 895 1966
rect 716 1963 717 1964
rect 711 1962 717 1963
rect 894 1963 895 1964
rect 899 1963 900 1967
rect 1070 1967 1076 1968
rect 1070 1966 1071 1967
rect 894 1962 900 1963
rect 944 1964 1071 1966
rect 944 1960 946 1964
rect 1070 1963 1071 1964
rect 1075 1963 1076 1967
rect 1326 1967 1327 1971
rect 1332 1967 1333 1971
rect 1326 1966 1333 1967
rect 1398 1971 1404 1972
rect 1398 1967 1399 1971
rect 1403 1970 1404 1971
rect 1407 1971 1413 1972
rect 1407 1970 1408 1971
rect 1403 1968 1408 1970
rect 1403 1967 1404 1968
rect 1398 1966 1404 1967
rect 1407 1967 1408 1968
rect 1412 1967 1413 1971
rect 1407 1966 1413 1967
rect 1478 1971 1484 1972
rect 1478 1967 1479 1971
rect 1483 1970 1484 1971
rect 1487 1971 1493 1972
rect 1487 1970 1488 1971
rect 1483 1968 1488 1970
rect 1483 1967 1484 1968
rect 1478 1966 1484 1967
rect 1487 1967 1488 1968
rect 1492 1967 1493 1971
rect 1487 1966 1493 1967
rect 1550 1971 1556 1972
rect 1550 1967 1551 1971
rect 1555 1970 1556 1971
rect 1567 1971 1573 1972
rect 1567 1970 1568 1971
rect 1555 1968 1568 1970
rect 1555 1967 1556 1968
rect 1550 1966 1556 1967
rect 1567 1967 1568 1968
rect 1572 1967 1573 1971
rect 1567 1966 1573 1967
rect 1639 1971 1648 1972
rect 1639 1967 1640 1971
rect 1647 1967 1648 1971
rect 1639 1966 1648 1967
rect 1694 1971 1700 1972
rect 1694 1967 1695 1971
rect 1699 1970 1700 1971
rect 1711 1971 1717 1972
rect 1711 1970 1712 1971
rect 1699 1968 1712 1970
rect 1699 1967 1700 1968
rect 1694 1966 1700 1967
rect 1711 1967 1712 1968
rect 1716 1967 1717 1971
rect 1711 1966 1717 1967
rect 1766 1971 1772 1972
rect 1766 1967 1767 1971
rect 1771 1970 1772 1971
rect 1775 1971 1781 1972
rect 1775 1970 1776 1971
rect 1771 1968 1776 1970
rect 1771 1967 1772 1968
rect 1766 1966 1772 1967
rect 1775 1967 1776 1968
rect 1780 1967 1781 1971
rect 1775 1966 1781 1967
rect 1830 1971 1836 1972
rect 1830 1967 1831 1971
rect 1835 1970 1836 1971
rect 1839 1971 1845 1972
rect 1839 1970 1840 1971
rect 1835 1968 1840 1970
rect 1835 1967 1836 1968
rect 1830 1966 1836 1967
rect 1839 1967 1840 1968
rect 1844 1967 1845 1971
rect 1839 1966 1845 1967
rect 1894 1971 1900 1972
rect 1894 1967 1895 1971
rect 1899 1970 1900 1971
rect 1903 1971 1909 1972
rect 1903 1970 1904 1971
rect 1899 1968 1904 1970
rect 1899 1967 1900 1968
rect 1894 1966 1900 1967
rect 1903 1967 1904 1968
rect 1908 1967 1909 1971
rect 1903 1966 1909 1967
rect 1966 1971 1972 1972
rect 1966 1967 1967 1971
rect 1971 1970 1972 1971
rect 1975 1971 1981 1972
rect 1975 1970 1976 1971
rect 1971 1968 1976 1970
rect 1971 1967 1972 1968
rect 1966 1966 1972 1967
rect 1975 1967 1976 1968
rect 1980 1967 1981 1971
rect 1975 1966 1981 1967
rect 2047 1971 2053 1972
rect 2047 1967 2048 1971
rect 2052 1970 2053 1971
rect 2078 1971 2084 1972
rect 2078 1970 2079 1971
rect 2052 1968 2079 1970
rect 2052 1967 2053 1968
rect 2047 1966 2053 1967
rect 2078 1967 2079 1968
rect 2083 1967 2084 1971
rect 2078 1966 2084 1967
rect 2086 1971 2092 1972
rect 2086 1967 2087 1971
rect 2091 1970 2092 1971
rect 2095 1971 2101 1972
rect 2118 1971 2124 1972
rect 2095 1970 2096 1971
rect 2091 1968 2096 1970
rect 2091 1967 2092 1968
rect 2086 1966 2092 1967
rect 2095 1967 2096 1968
rect 2100 1967 2101 1971
rect 2095 1966 2101 1967
rect 1070 1962 1076 1963
rect 215 1959 221 1960
rect 110 1956 116 1957
rect 110 1952 111 1956
rect 115 1952 116 1956
rect 215 1955 216 1959
rect 220 1958 221 1959
rect 262 1959 268 1960
rect 262 1958 263 1959
rect 220 1956 263 1958
rect 220 1955 221 1956
rect 215 1954 221 1955
rect 262 1955 263 1956
rect 267 1955 268 1959
rect 262 1954 268 1955
rect 271 1959 277 1960
rect 271 1955 272 1959
rect 276 1958 277 1959
rect 326 1959 332 1960
rect 326 1958 327 1959
rect 276 1956 327 1958
rect 276 1955 277 1956
rect 271 1954 277 1955
rect 326 1955 327 1956
rect 331 1955 332 1959
rect 326 1954 332 1955
rect 334 1959 341 1960
rect 334 1955 335 1959
rect 340 1955 341 1959
rect 334 1954 341 1955
rect 399 1959 405 1960
rect 399 1955 400 1959
rect 404 1958 405 1959
rect 462 1959 468 1960
rect 462 1958 463 1959
rect 404 1956 463 1958
rect 404 1955 405 1956
rect 399 1954 405 1955
rect 462 1955 463 1956
rect 467 1955 468 1959
rect 462 1954 468 1955
rect 471 1959 477 1960
rect 471 1955 472 1959
rect 476 1958 477 1959
rect 534 1959 540 1960
rect 534 1958 535 1959
rect 476 1956 535 1958
rect 476 1955 477 1956
rect 471 1954 477 1955
rect 534 1955 535 1956
rect 539 1955 540 1959
rect 534 1954 540 1955
rect 543 1959 552 1960
rect 543 1955 544 1959
rect 551 1955 552 1959
rect 543 1954 552 1955
rect 606 1959 612 1960
rect 606 1955 607 1959
rect 611 1958 612 1959
rect 615 1959 621 1960
rect 615 1958 616 1959
rect 611 1956 616 1958
rect 611 1955 612 1956
rect 606 1954 612 1955
rect 615 1955 616 1956
rect 620 1955 621 1959
rect 615 1954 621 1955
rect 623 1959 629 1960
rect 623 1955 624 1959
rect 628 1958 629 1959
rect 679 1959 685 1960
rect 679 1958 680 1959
rect 628 1956 680 1958
rect 628 1955 629 1956
rect 623 1954 629 1955
rect 679 1955 680 1956
rect 684 1955 685 1959
rect 679 1954 685 1955
rect 687 1959 693 1960
rect 687 1955 688 1959
rect 692 1958 693 1959
rect 743 1959 749 1960
rect 743 1958 744 1959
rect 692 1956 744 1958
rect 692 1955 693 1956
rect 687 1954 693 1955
rect 743 1955 744 1956
rect 748 1955 749 1959
rect 743 1954 749 1955
rect 751 1959 757 1960
rect 751 1955 752 1959
rect 756 1958 757 1959
rect 799 1959 805 1960
rect 799 1958 800 1959
rect 756 1956 800 1958
rect 756 1955 757 1956
rect 751 1954 757 1955
rect 799 1955 800 1956
rect 804 1955 805 1959
rect 799 1954 805 1955
rect 807 1959 813 1960
rect 807 1955 808 1959
rect 812 1958 813 1959
rect 847 1959 853 1960
rect 847 1958 848 1959
rect 812 1956 848 1958
rect 812 1955 813 1956
rect 807 1954 813 1955
rect 847 1955 848 1956
rect 852 1955 853 1959
rect 847 1954 853 1955
rect 858 1959 864 1960
rect 858 1955 859 1959
rect 863 1958 864 1959
rect 895 1959 901 1960
rect 895 1958 896 1959
rect 863 1956 896 1958
rect 863 1955 864 1956
rect 858 1954 864 1955
rect 895 1955 896 1956
rect 900 1955 901 1959
rect 895 1954 901 1955
rect 943 1959 949 1960
rect 943 1955 944 1959
rect 948 1955 949 1959
rect 943 1954 949 1955
rect 951 1959 957 1960
rect 951 1955 952 1959
rect 956 1958 957 1959
rect 991 1959 997 1960
rect 991 1958 992 1959
rect 956 1956 992 1958
rect 956 1955 957 1956
rect 951 1954 957 1955
rect 991 1955 992 1956
rect 996 1955 997 1959
rect 991 1954 997 1955
rect 1014 1959 1020 1960
rect 1014 1955 1015 1959
rect 1019 1958 1020 1959
rect 1031 1959 1037 1960
rect 1031 1958 1032 1959
rect 1019 1956 1032 1958
rect 1019 1955 1020 1956
rect 1014 1954 1020 1955
rect 1031 1955 1032 1956
rect 1036 1955 1037 1959
rect 1031 1954 1037 1955
rect 1054 1959 1060 1960
rect 1054 1955 1055 1959
rect 1059 1958 1060 1959
rect 1071 1959 1077 1960
rect 1071 1958 1072 1959
rect 1059 1956 1072 1958
rect 1059 1955 1060 1956
rect 1054 1954 1060 1955
rect 1071 1955 1072 1956
rect 1076 1955 1077 1959
rect 1134 1959 1140 1960
rect 1071 1954 1077 1955
rect 1094 1956 1100 1957
rect 110 1951 116 1952
rect 1094 1952 1095 1956
rect 1099 1952 1100 1956
rect 1134 1955 1135 1959
rect 1139 1955 1140 1959
rect 2118 1959 2124 1960
rect 1134 1954 1140 1955
rect 1302 1956 1308 1957
rect 1094 1951 1100 1952
rect 1302 1952 1303 1956
rect 1307 1952 1308 1956
rect 1302 1951 1308 1952
rect 1382 1956 1388 1957
rect 1382 1952 1383 1956
rect 1387 1952 1388 1956
rect 1382 1951 1388 1952
rect 1462 1956 1468 1957
rect 1462 1952 1463 1956
rect 1467 1952 1468 1956
rect 1462 1951 1468 1952
rect 1542 1956 1548 1957
rect 1542 1952 1543 1956
rect 1547 1952 1548 1956
rect 1542 1951 1548 1952
rect 1614 1956 1620 1957
rect 1614 1952 1615 1956
rect 1619 1952 1620 1956
rect 1614 1951 1620 1952
rect 1686 1956 1692 1957
rect 1686 1952 1687 1956
rect 1691 1952 1692 1956
rect 1686 1951 1692 1952
rect 1750 1956 1756 1957
rect 1750 1952 1751 1956
rect 1755 1952 1756 1956
rect 1750 1951 1756 1952
rect 1814 1956 1820 1957
rect 1814 1952 1815 1956
rect 1819 1952 1820 1956
rect 1814 1951 1820 1952
rect 1878 1956 1884 1957
rect 1878 1952 1879 1956
rect 1883 1952 1884 1956
rect 1878 1951 1884 1952
rect 1950 1956 1956 1957
rect 1950 1952 1951 1956
rect 1955 1952 1956 1956
rect 1950 1951 1956 1952
rect 2022 1956 2028 1957
rect 2022 1952 2023 1956
rect 2027 1952 2028 1956
rect 2022 1951 2028 1952
rect 2070 1956 2076 1957
rect 2070 1952 2071 1956
rect 2075 1952 2076 1956
rect 2118 1955 2119 1959
rect 2123 1955 2124 1959
rect 2118 1954 2124 1955
rect 2070 1951 2076 1952
rect 190 1948 196 1949
rect 190 1944 191 1948
rect 195 1944 196 1948
rect 190 1943 196 1944
rect 246 1948 252 1949
rect 246 1944 247 1948
rect 251 1944 252 1948
rect 246 1943 252 1944
rect 310 1948 316 1949
rect 310 1944 311 1948
rect 315 1944 316 1948
rect 310 1943 316 1944
rect 374 1948 380 1949
rect 374 1944 375 1948
rect 379 1944 380 1948
rect 374 1943 380 1944
rect 446 1948 452 1949
rect 446 1944 447 1948
rect 451 1944 452 1948
rect 446 1943 452 1944
rect 518 1948 524 1949
rect 518 1944 519 1948
rect 523 1944 524 1948
rect 518 1943 524 1944
rect 590 1948 596 1949
rect 590 1944 591 1948
rect 595 1944 596 1948
rect 590 1943 596 1944
rect 654 1948 660 1949
rect 654 1944 655 1948
rect 659 1944 660 1948
rect 654 1943 660 1944
rect 718 1948 724 1949
rect 718 1944 719 1948
rect 723 1944 724 1948
rect 718 1943 724 1944
rect 774 1948 780 1949
rect 774 1944 775 1948
rect 779 1944 780 1948
rect 774 1943 780 1944
rect 822 1948 828 1949
rect 822 1944 823 1948
rect 827 1944 828 1948
rect 822 1943 828 1944
rect 870 1948 876 1949
rect 870 1944 871 1948
rect 875 1944 876 1948
rect 870 1943 876 1944
rect 918 1948 924 1949
rect 918 1944 919 1948
rect 923 1944 924 1948
rect 918 1943 924 1944
rect 966 1948 972 1949
rect 966 1944 967 1948
rect 971 1944 972 1948
rect 966 1943 972 1944
rect 1006 1948 1012 1949
rect 1006 1944 1007 1948
rect 1011 1944 1012 1948
rect 1006 1943 1012 1944
rect 1046 1948 1052 1949
rect 1046 1944 1047 1948
rect 1051 1944 1052 1948
rect 1046 1943 1052 1944
rect 1158 1940 1164 1941
rect 214 1939 221 1940
rect 214 1935 215 1939
rect 220 1935 221 1939
rect 214 1934 221 1935
rect 262 1939 268 1940
rect 262 1935 263 1939
rect 267 1938 268 1939
rect 271 1939 277 1940
rect 271 1938 272 1939
rect 267 1936 272 1938
rect 267 1935 268 1936
rect 262 1934 268 1935
rect 271 1935 272 1936
rect 276 1935 277 1939
rect 271 1934 277 1935
rect 326 1939 332 1940
rect 326 1935 327 1939
rect 331 1938 332 1939
rect 335 1939 341 1940
rect 335 1938 336 1939
rect 331 1936 336 1938
rect 331 1935 332 1936
rect 326 1934 332 1935
rect 335 1935 336 1936
rect 340 1935 341 1939
rect 335 1934 341 1935
rect 394 1939 405 1940
rect 394 1935 395 1939
rect 399 1935 400 1939
rect 404 1935 405 1939
rect 394 1934 405 1935
rect 462 1939 468 1940
rect 462 1935 463 1939
rect 467 1938 468 1939
rect 471 1939 477 1940
rect 471 1938 472 1939
rect 467 1936 472 1938
rect 467 1935 468 1936
rect 462 1934 468 1935
rect 471 1935 472 1936
rect 476 1935 477 1939
rect 471 1934 477 1935
rect 534 1939 540 1940
rect 534 1935 535 1939
rect 539 1938 540 1939
rect 543 1939 549 1940
rect 543 1938 544 1939
rect 539 1936 544 1938
rect 539 1935 540 1936
rect 534 1934 540 1935
rect 543 1935 544 1936
rect 548 1935 549 1939
rect 543 1934 549 1935
rect 615 1939 621 1940
rect 615 1935 616 1939
rect 620 1938 621 1939
rect 623 1939 629 1940
rect 623 1938 624 1939
rect 620 1936 624 1938
rect 620 1935 621 1936
rect 615 1934 621 1935
rect 623 1935 624 1936
rect 628 1935 629 1939
rect 623 1934 629 1935
rect 679 1939 685 1940
rect 679 1935 680 1939
rect 684 1938 685 1939
rect 687 1939 693 1940
rect 687 1938 688 1939
rect 684 1936 688 1938
rect 684 1935 685 1936
rect 679 1934 685 1935
rect 687 1935 688 1936
rect 692 1935 693 1939
rect 687 1934 693 1935
rect 743 1939 749 1940
rect 743 1935 744 1939
rect 748 1938 749 1939
rect 751 1939 757 1940
rect 751 1938 752 1939
rect 748 1936 752 1938
rect 748 1935 749 1936
rect 743 1934 749 1935
rect 751 1935 752 1936
rect 756 1935 757 1939
rect 751 1934 757 1935
rect 799 1939 805 1940
rect 799 1935 800 1939
rect 804 1938 805 1939
rect 807 1939 813 1940
rect 807 1938 808 1939
rect 804 1936 808 1938
rect 804 1935 805 1936
rect 799 1934 805 1935
rect 807 1935 808 1936
rect 812 1935 813 1939
rect 807 1934 813 1935
rect 847 1939 853 1940
rect 847 1935 848 1939
rect 852 1938 853 1939
rect 858 1939 864 1940
rect 858 1938 859 1939
rect 852 1936 859 1938
rect 852 1935 853 1936
rect 847 1934 853 1935
rect 858 1935 859 1936
rect 863 1935 864 1939
rect 858 1934 864 1935
rect 894 1939 901 1940
rect 894 1935 895 1939
rect 900 1935 901 1939
rect 894 1934 901 1935
rect 943 1939 949 1940
rect 943 1935 944 1939
rect 948 1938 949 1939
rect 951 1939 957 1940
rect 951 1938 952 1939
rect 948 1936 952 1938
rect 948 1935 949 1936
rect 943 1934 949 1935
rect 951 1935 952 1936
rect 956 1935 957 1939
rect 951 1934 957 1935
rect 991 1939 997 1940
rect 991 1935 992 1939
rect 996 1938 997 1939
rect 1014 1939 1020 1940
rect 1014 1938 1015 1939
rect 996 1936 1015 1938
rect 996 1935 997 1936
rect 991 1934 997 1935
rect 1014 1935 1015 1936
rect 1019 1935 1020 1939
rect 1014 1934 1020 1935
rect 1031 1939 1037 1940
rect 1031 1935 1032 1939
rect 1036 1938 1037 1939
rect 1054 1939 1060 1940
rect 1054 1938 1055 1939
rect 1036 1936 1055 1938
rect 1036 1935 1037 1936
rect 1031 1934 1037 1935
rect 1054 1935 1055 1936
rect 1059 1935 1060 1939
rect 1054 1934 1060 1935
rect 1071 1939 1077 1940
rect 1071 1935 1072 1939
rect 1076 1935 1077 1939
rect 1071 1934 1077 1935
rect 1134 1937 1140 1938
rect 606 1927 612 1928
rect 606 1923 607 1927
rect 611 1926 612 1927
rect 1073 1926 1075 1934
rect 1134 1933 1135 1937
rect 1139 1933 1140 1937
rect 1158 1936 1159 1940
rect 1163 1936 1164 1940
rect 1158 1935 1164 1936
rect 1222 1940 1228 1941
rect 1222 1936 1223 1940
rect 1227 1936 1228 1940
rect 1222 1935 1228 1936
rect 1302 1940 1308 1941
rect 1302 1936 1303 1940
rect 1307 1936 1308 1940
rect 1302 1935 1308 1936
rect 1382 1940 1388 1941
rect 1382 1936 1383 1940
rect 1387 1936 1388 1940
rect 1382 1935 1388 1936
rect 1462 1940 1468 1941
rect 1462 1936 1463 1940
rect 1467 1936 1468 1940
rect 1462 1935 1468 1936
rect 1534 1940 1540 1941
rect 1534 1936 1535 1940
rect 1539 1936 1540 1940
rect 1534 1935 1540 1936
rect 1614 1940 1620 1941
rect 1614 1936 1615 1940
rect 1619 1936 1620 1940
rect 1614 1935 1620 1936
rect 1694 1940 1700 1941
rect 1694 1936 1695 1940
rect 1699 1936 1700 1940
rect 1694 1935 1700 1936
rect 1782 1940 1788 1941
rect 1782 1936 1783 1940
rect 1787 1936 1788 1940
rect 1782 1935 1788 1936
rect 1878 1940 1884 1941
rect 1878 1936 1879 1940
rect 1883 1936 1884 1940
rect 1878 1935 1884 1936
rect 1982 1940 1988 1941
rect 1982 1936 1983 1940
rect 1987 1936 1988 1940
rect 1982 1935 1988 1936
rect 2070 1940 2076 1941
rect 2070 1936 2071 1940
rect 2075 1936 2076 1940
rect 2070 1935 2076 1936
rect 2118 1937 2124 1938
rect 1134 1932 1140 1933
rect 2118 1933 2119 1937
rect 2123 1933 2124 1937
rect 2118 1932 2124 1933
rect 2006 1931 2012 1932
rect 2006 1930 2007 1931
rect 1560 1928 2007 1930
rect 611 1924 866 1926
rect 1073 1924 1187 1926
rect 1560 1924 1562 1928
rect 2006 1927 2007 1928
rect 2011 1927 2012 1931
rect 2006 1926 2012 1927
rect 611 1923 612 1924
rect 606 1922 612 1923
rect 159 1919 165 1920
rect 159 1915 160 1919
rect 164 1918 165 1919
rect 190 1919 196 1920
rect 190 1918 191 1919
rect 164 1916 191 1918
rect 164 1915 165 1916
rect 159 1914 165 1915
rect 190 1915 191 1916
rect 195 1915 196 1919
rect 190 1914 196 1915
rect 199 1919 205 1920
rect 199 1915 200 1919
rect 204 1918 205 1919
rect 246 1919 252 1920
rect 246 1918 247 1919
rect 204 1916 247 1918
rect 204 1915 205 1916
rect 199 1914 205 1915
rect 246 1915 247 1916
rect 251 1915 252 1919
rect 246 1914 252 1915
rect 255 1919 261 1920
rect 255 1915 256 1919
rect 260 1918 261 1919
rect 286 1919 292 1920
rect 286 1918 287 1919
rect 260 1916 287 1918
rect 260 1915 261 1916
rect 255 1914 261 1915
rect 286 1915 287 1916
rect 291 1915 292 1919
rect 286 1914 292 1915
rect 319 1919 325 1920
rect 319 1915 320 1919
rect 324 1918 325 1919
rect 334 1919 340 1920
rect 334 1918 335 1919
rect 324 1916 335 1918
rect 324 1915 325 1916
rect 319 1914 325 1915
rect 334 1915 335 1916
rect 339 1915 340 1919
rect 334 1914 340 1915
rect 391 1919 397 1920
rect 391 1915 392 1919
rect 396 1918 397 1919
rect 438 1919 444 1920
rect 438 1918 439 1919
rect 396 1916 439 1918
rect 396 1915 397 1916
rect 391 1914 397 1915
rect 438 1915 439 1916
rect 443 1915 444 1919
rect 438 1914 444 1915
rect 455 1919 461 1920
rect 455 1915 456 1919
rect 460 1918 461 1919
rect 502 1919 508 1920
rect 502 1918 503 1919
rect 460 1916 503 1918
rect 460 1915 461 1916
rect 455 1914 461 1915
rect 502 1915 503 1916
rect 507 1915 508 1919
rect 502 1914 508 1915
rect 510 1919 516 1920
rect 510 1915 511 1919
rect 515 1918 516 1919
rect 519 1919 525 1920
rect 519 1918 520 1919
rect 515 1916 520 1918
rect 515 1915 516 1916
rect 510 1914 516 1915
rect 519 1915 520 1916
rect 524 1915 525 1919
rect 519 1914 525 1915
rect 583 1919 589 1920
rect 583 1915 584 1919
rect 588 1918 589 1919
rect 630 1919 636 1920
rect 630 1918 631 1919
rect 588 1916 631 1918
rect 588 1915 589 1916
rect 583 1914 589 1915
rect 630 1915 631 1916
rect 635 1915 636 1919
rect 630 1914 636 1915
rect 639 1919 645 1920
rect 639 1915 640 1919
rect 644 1918 645 1919
rect 686 1919 692 1920
rect 686 1918 687 1919
rect 644 1916 687 1918
rect 644 1915 645 1916
rect 639 1914 645 1915
rect 686 1915 687 1916
rect 691 1915 692 1919
rect 686 1914 692 1915
rect 695 1919 701 1920
rect 695 1915 696 1919
rect 700 1918 701 1919
rect 742 1919 748 1920
rect 742 1918 743 1919
rect 700 1916 743 1918
rect 700 1915 701 1916
rect 695 1914 701 1915
rect 742 1915 743 1916
rect 747 1915 748 1919
rect 742 1914 748 1915
rect 751 1919 757 1920
rect 751 1915 752 1919
rect 756 1918 757 1919
rect 798 1919 804 1920
rect 798 1918 799 1919
rect 756 1916 799 1918
rect 756 1915 757 1916
rect 751 1914 757 1915
rect 798 1915 799 1916
rect 803 1915 804 1919
rect 798 1914 804 1915
rect 807 1919 813 1920
rect 807 1915 808 1919
rect 812 1918 813 1919
rect 854 1919 860 1920
rect 854 1918 855 1919
rect 812 1916 855 1918
rect 812 1915 813 1916
rect 807 1914 813 1915
rect 854 1915 855 1916
rect 859 1915 860 1919
rect 864 1918 866 1924
rect 1183 1923 1189 1924
rect 1134 1920 1140 1921
rect 871 1919 877 1920
rect 871 1918 872 1919
rect 864 1916 872 1918
rect 854 1914 860 1915
rect 871 1915 872 1916
rect 876 1915 877 1919
rect 1134 1916 1135 1920
rect 1139 1916 1140 1920
rect 1183 1919 1184 1923
rect 1188 1919 1189 1923
rect 1183 1918 1189 1919
rect 1191 1923 1197 1924
rect 1191 1919 1192 1923
rect 1196 1922 1197 1923
rect 1247 1923 1253 1924
rect 1247 1922 1248 1923
rect 1196 1920 1248 1922
rect 1196 1919 1197 1920
rect 1191 1918 1197 1919
rect 1247 1919 1248 1920
rect 1252 1919 1253 1923
rect 1247 1918 1253 1919
rect 1327 1923 1333 1924
rect 1327 1919 1328 1923
rect 1332 1922 1333 1923
rect 1398 1923 1404 1924
rect 1398 1922 1399 1923
rect 1332 1920 1399 1922
rect 1332 1919 1333 1920
rect 1327 1918 1333 1919
rect 1398 1919 1399 1920
rect 1403 1919 1404 1923
rect 1398 1918 1404 1919
rect 1407 1923 1413 1924
rect 1407 1919 1408 1923
rect 1412 1922 1413 1923
rect 1446 1923 1452 1924
rect 1446 1922 1447 1923
rect 1412 1920 1447 1922
rect 1412 1919 1413 1920
rect 1407 1918 1413 1919
rect 1446 1919 1447 1920
rect 1451 1919 1452 1923
rect 1446 1918 1452 1919
rect 1474 1923 1480 1924
rect 1474 1919 1475 1923
rect 1479 1922 1480 1923
rect 1487 1923 1493 1924
rect 1487 1922 1488 1923
rect 1479 1920 1488 1922
rect 1479 1919 1480 1920
rect 1474 1918 1480 1919
rect 1487 1919 1488 1920
rect 1492 1919 1493 1923
rect 1487 1918 1493 1919
rect 1559 1923 1565 1924
rect 1559 1919 1560 1923
rect 1564 1919 1565 1923
rect 1559 1918 1565 1919
rect 1567 1923 1573 1924
rect 1567 1919 1568 1923
rect 1572 1922 1573 1923
rect 1639 1923 1645 1924
rect 1639 1922 1640 1923
rect 1572 1920 1640 1922
rect 1572 1919 1573 1920
rect 1567 1918 1573 1919
rect 1639 1919 1640 1920
rect 1644 1919 1645 1923
rect 1639 1918 1645 1919
rect 1647 1923 1653 1924
rect 1647 1919 1648 1923
rect 1652 1922 1653 1923
rect 1719 1923 1725 1924
rect 1719 1922 1720 1923
rect 1652 1920 1720 1922
rect 1652 1919 1653 1920
rect 1647 1918 1653 1919
rect 1719 1919 1720 1920
rect 1724 1919 1725 1923
rect 1719 1918 1725 1919
rect 1806 1923 1813 1924
rect 1806 1919 1807 1923
rect 1812 1919 1813 1923
rect 1806 1918 1813 1919
rect 1815 1923 1821 1924
rect 1815 1919 1816 1923
rect 1820 1922 1821 1923
rect 1903 1923 1909 1924
rect 1903 1922 1904 1923
rect 1820 1920 1904 1922
rect 1820 1919 1821 1920
rect 1815 1918 1821 1919
rect 1903 1919 1904 1920
rect 1908 1919 1909 1923
rect 1903 1918 1909 1919
rect 1911 1923 1917 1924
rect 1911 1919 1912 1923
rect 1916 1922 1917 1923
rect 2007 1923 2013 1924
rect 2007 1922 2008 1923
rect 1916 1920 2008 1922
rect 1916 1919 1917 1920
rect 1911 1918 1917 1919
rect 2007 1919 2008 1920
rect 2012 1919 2013 1923
rect 2007 1918 2013 1919
rect 2094 1923 2101 1924
rect 2094 1919 2095 1923
rect 2100 1919 2101 1923
rect 2094 1918 2101 1919
rect 2118 1920 2124 1921
rect 1134 1915 1140 1916
rect 2118 1916 2119 1920
rect 2123 1916 2124 1920
rect 2118 1915 2124 1916
rect 871 1914 877 1915
rect 134 1912 140 1913
rect 134 1908 135 1912
rect 139 1908 140 1912
rect 134 1907 140 1908
rect 174 1912 180 1913
rect 174 1908 175 1912
rect 179 1908 180 1912
rect 174 1907 180 1908
rect 230 1912 236 1913
rect 230 1908 231 1912
rect 235 1908 236 1912
rect 230 1907 236 1908
rect 294 1912 300 1913
rect 294 1908 295 1912
rect 299 1908 300 1912
rect 294 1907 300 1908
rect 366 1912 372 1913
rect 366 1908 367 1912
rect 371 1908 372 1912
rect 366 1907 372 1908
rect 430 1912 436 1913
rect 430 1908 431 1912
rect 435 1908 436 1912
rect 430 1907 436 1908
rect 494 1912 500 1913
rect 494 1908 495 1912
rect 499 1908 500 1912
rect 494 1907 500 1908
rect 558 1912 564 1913
rect 558 1908 559 1912
rect 563 1908 564 1912
rect 558 1907 564 1908
rect 614 1912 620 1913
rect 614 1908 615 1912
rect 619 1908 620 1912
rect 614 1907 620 1908
rect 670 1912 676 1913
rect 670 1908 671 1912
rect 675 1908 676 1912
rect 670 1907 676 1908
rect 726 1912 732 1913
rect 726 1908 727 1912
rect 731 1908 732 1912
rect 726 1907 732 1908
rect 782 1912 788 1913
rect 782 1908 783 1912
rect 787 1908 788 1912
rect 782 1907 788 1908
rect 846 1912 852 1913
rect 846 1908 847 1912
rect 851 1908 852 1912
rect 846 1907 852 1908
rect 1158 1912 1164 1913
rect 1158 1908 1159 1912
rect 1163 1908 1164 1912
rect 1158 1907 1164 1908
rect 1222 1912 1228 1913
rect 1222 1908 1223 1912
rect 1227 1908 1228 1912
rect 1222 1907 1228 1908
rect 1302 1912 1308 1913
rect 1302 1908 1303 1912
rect 1307 1908 1308 1912
rect 1302 1907 1308 1908
rect 1382 1912 1388 1913
rect 1382 1908 1383 1912
rect 1387 1908 1388 1912
rect 1382 1907 1388 1908
rect 1462 1912 1468 1913
rect 1462 1908 1463 1912
rect 1467 1908 1468 1912
rect 1462 1907 1468 1908
rect 1534 1912 1540 1913
rect 1534 1908 1535 1912
rect 1539 1908 1540 1912
rect 1534 1907 1540 1908
rect 1614 1912 1620 1913
rect 1614 1908 1615 1912
rect 1619 1908 1620 1912
rect 1614 1907 1620 1908
rect 1694 1912 1700 1913
rect 1694 1908 1695 1912
rect 1699 1908 1700 1912
rect 1694 1907 1700 1908
rect 1782 1912 1788 1913
rect 1782 1908 1783 1912
rect 1787 1908 1788 1912
rect 1782 1907 1788 1908
rect 1878 1912 1884 1913
rect 1878 1908 1879 1912
rect 1883 1908 1884 1912
rect 1878 1907 1884 1908
rect 1982 1912 1988 1913
rect 1982 1908 1983 1912
rect 1987 1908 1988 1912
rect 1982 1907 1988 1908
rect 2070 1912 2076 1913
rect 2070 1908 2071 1912
rect 2075 1908 2076 1912
rect 2070 1907 2076 1908
rect 110 1904 116 1905
rect 110 1900 111 1904
rect 115 1900 116 1904
rect 1094 1904 1100 1905
rect 1094 1900 1095 1904
rect 1099 1900 1100 1904
rect 110 1899 116 1900
rect 158 1899 165 1900
rect 158 1895 159 1899
rect 164 1895 165 1899
rect 158 1894 165 1895
rect 190 1899 196 1900
rect 190 1895 191 1899
rect 195 1898 196 1899
rect 199 1899 205 1900
rect 199 1898 200 1899
rect 195 1896 200 1898
rect 195 1895 196 1896
rect 190 1894 196 1895
rect 199 1895 200 1896
rect 204 1895 205 1899
rect 199 1894 205 1895
rect 246 1899 252 1900
rect 246 1895 247 1899
rect 251 1898 252 1899
rect 255 1899 261 1900
rect 255 1898 256 1899
rect 251 1896 256 1898
rect 251 1895 252 1896
rect 246 1894 252 1895
rect 255 1895 256 1896
rect 260 1895 261 1899
rect 255 1894 261 1895
rect 286 1899 292 1900
rect 286 1895 287 1899
rect 291 1898 292 1899
rect 319 1899 325 1900
rect 319 1898 320 1899
rect 291 1896 320 1898
rect 291 1895 292 1896
rect 286 1894 292 1895
rect 319 1895 320 1896
rect 324 1895 325 1899
rect 319 1894 325 1895
rect 391 1899 400 1900
rect 391 1895 392 1899
rect 399 1895 400 1899
rect 391 1894 400 1895
rect 438 1899 444 1900
rect 438 1895 439 1899
rect 443 1898 444 1899
rect 455 1899 461 1900
rect 455 1898 456 1899
rect 443 1896 456 1898
rect 443 1895 444 1896
rect 438 1894 444 1895
rect 455 1895 456 1896
rect 460 1895 461 1899
rect 455 1894 461 1895
rect 502 1899 508 1900
rect 502 1895 503 1899
rect 507 1898 508 1899
rect 519 1899 525 1900
rect 519 1898 520 1899
rect 507 1896 520 1898
rect 507 1895 508 1896
rect 502 1894 508 1895
rect 519 1895 520 1896
rect 524 1895 525 1899
rect 519 1894 525 1895
rect 583 1899 589 1900
rect 583 1895 584 1899
rect 588 1898 589 1899
rect 622 1899 628 1900
rect 622 1898 623 1899
rect 588 1896 623 1898
rect 588 1895 589 1896
rect 583 1894 589 1895
rect 622 1895 623 1896
rect 627 1895 628 1899
rect 622 1894 628 1895
rect 630 1899 636 1900
rect 630 1895 631 1899
rect 635 1898 636 1899
rect 639 1899 645 1900
rect 639 1898 640 1899
rect 635 1896 640 1898
rect 635 1895 636 1896
rect 630 1894 636 1895
rect 639 1895 640 1896
rect 644 1895 645 1899
rect 639 1894 645 1895
rect 686 1899 692 1900
rect 686 1895 687 1899
rect 691 1898 692 1899
rect 695 1899 701 1900
rect 695 1898 696 1899
rect 691 1896 696 1898
rect 691 1895 692 1896
rect 686 1894 692 1895
rect 695 1895 696 1896
rect 700 1895 701 1899
rect 695 1894 701 1895
rect 742 1899 748 1900
rect 742 1895 743 1899
rect 747 1898 748 1899
rect 751 1899 757 1900
rect 751 1898 752 1899
rect 747 1896 752 1898
rect 747 1895 748 1896
rect 742 1894 748 1895
rect 751 1895 752 1896
rect 756 1895 757 1899
rect 751 1894 757 1895
rect 798 1899 804 1900
rect 798 1895 799 1899
rect 803 1898 804 1899
rect 807 1899 813 1900
rect 807 1898 808 1899
rect 803 1896 808 1898
rect 803 1895 804 1896
rect 798 1894 804 1895
rect 807 1895 808 1896
rect 812 1895 813 1899
rect 807 1894 813 1895
rect 854 1899 860 1900
rect 854 1895 855 1899
rect 859 1898 860 1899
rect 871 1899 877 1900
rect 1094 1899 1100 1900
rect 1183 1903 1189 1904
rect 1183 1899 1184 1903
rect 1188 1902 1189 1903
rect 1191 1903 1197 1904
rect 1191 1902 1192 1903
rect 1188 1900 1192 1902
rect 1188 1899 1189 1900
rect 871 1898 872 1899
rect 859 1896 872 1898
rect 859 1895 860 1896
rect 854 1894 860 1895
rect 871 1895 872 1896
rect 876 1895 877 1899
rect 1183 1898 1189 1899
rect 1191 1899 1192 1900
rect 1196 1899 1197 1903
rect 1191 1898 1197 1899
rect 1206 1903 1212 1904
rect 1206 1899 1207 1903
rect 1211 1902 1212 1903
rect 1247 1903 1253 1904
rect 1247 1902 1248 1903
rect 1211 1900 1248 1902
rect 1211 1899 1212 1900
rect 1206 1898 1212 1899
rect 1247 1899 1248 1900
rect 1252 1899 1253 1903
rect 1247 1898 1253 1899
rect 1326 1903 1333 1904
rect 1326 1899 1327 1903
rect 1332 1899 1333 1903
rect 1326 1898 1333 1899
rect 1398 1903 1404 1904
rect 1398 1899 1399 1903
rect 1403 1902 1404 1903
rect 1407 1903 1413 1904
rect 1407 1902 1408 1903
rect 1403 1900 1408 1902
rect 1403 1899 1404 1900
rect 1398 1898 1404 1899
rect 1407 1899 1408 1900
rect 1412 1899 1413 1903
rect 1407 1898 1413 1899
rect 1446 1903 1452 1904
rect 1446 1899 1447 1903
rect 1451 1902 1452 1903
rect 1487 1903 1493 1904
rect 1487 1902 1488 1903
rect 1451 1900 1488 1902
rect 1451 1899 1452 1900
rect 1446 1898 1452 1899
rect 1487 1899 1488 1900
rect 1492 1899 1493 1903
rect 1487 1898 1493 1899
rect 1559 1903 1565 1904
rect 1559 1899 1560 1903
rect 1564 1902 1565 1903
rect 1567 1903 1573 1904
rect 1567 1902 1568 1903
rect 1564 1900 1568 1902
rect 1564 1899 1565 1900
rect 1559 1898 1565 1899
rect 1567 1899 1568 1900
rect 1572 1899 1573 1903
rect 1567 1898 1573 1899
rect 1639 1903 1645 1904
rect 1639 1899 1640 1903
rect 1644 1902 1645 1903
rect 1647 1903 1653 1904
rect 1647 1902 1648 1903
rect 1644 1900 1648 1902
rect 1644 1899 1645 1900
rect 1639 1898 1645 1899
rect 1647 1899 1648 1900
rect 1652 1899 1653 1903
rect 1647 1898 1653 1899
rect 1719 1903 1725 1904
rect 1719 1899 1720 1903
rect 1724 1902 1725 1903
rect 1734 1903 1740 1904
rect 1734 1902 1735 1903
rect 1724 1900 1735 1902
rect 1724 1899 1725 1900
rect 1719 1898 1725 1899
rect 1734 1899 1735 1900
rect 1739 1899 1740 1903
rect 1734 1898 1740 1899
rect 1807 1903 1813 1904
rect 1807 1899 1808 1903
rect 1812 1902 1813 1903
rect 1815 1903 1821 1904
rect 1815 1902 1816 1903
rect 1812 1900 1816 1902
rect 1812 1899 1813 1900
rect 1807 1898 1813 1899
rect 1815 1899 1816 1900
rect 1820 1899 1821 1903
rect 1815 1898 1821 1899
rect 1903 1903 1909 1904
rect 1903 1899 1904 1903
rect 1908 1902 1909 1903
rect 1911 1903 1917 1904
rect 1911 1902 1912 1903
rect 1908 1900 1912 1902
rect 1908 1899 1909 1900
rect 1903 1898 1909 1899
rect 1911 1899 1912 1900
rect 1916 1899 1917 1903
rect 1911 1898 1917 1899
rect 2006 1903 2013 1904
rect 2006 1899 2007 1903
rect 2012 1899 2013 1903
rect 2006 1898 2013 1899
rect 2078 1903 2084 1904
rect 2078 1899 2079 1903
rect 2083 1902 2084 1903
rect 2095 1903 2101 1904
rect 2095 1902 2096 1903
rect 2083 1900 2096 1902
rect 2083 1899 2084 1900
rect 2078 1898 2084 1899
rect 2095 1899 2096 1900
rect 2100 1899 2101 1903
rect 2095 1898 2101 1899
rect 871 1894 877 1895
rect 110 1887 116 1888
rect 110 1883 111 1887
rect 115 1883 116 1887
rect 1094 1887 1100 1888
rect 110 1882 116 1883
rect 134 1884 140 1885
rect 134 1880 135 1884
rect 139 1880 140 1884
rect 134 1879 140 1880
rect 174 1884 180 1885
rect 174 1880 175 1884
rect 179 1880 180 1884
rect 174 1879 180 1880
rect 230 1884 236 1885
rect 230 1880 231 1884
rect 235 1880 236 1884
rect 230 1879 236 1880
rect 294 1884 300 1885
rect 294 1880 295 1884
rect 299 1880 300 1884
rect 294 1879 300 1880
rect 366 1884 372 1885
rect 366 1880 367 1884
rect 371 1880 372 1884
rect 366 1879 372 1880
rect 430 1884 436 1885
rect 430 1880 431 1884
rect 435 1880 436 1884
rect 430 1879 436 1880
rect 494 1884 500 1885
rect 494 1880 495 1884
rect 499 1880 500 1884
rect 494 1879 500 1880
rect 558 1884 564 1885
rect 558 1880 559 1884
rect 563 1880 564 1884
rect 558 1879 564 1880
rect 614 1884 620 1885
rect 614 1880 615 1884
rect 619 1880 620 1884
rect 614 1879 620 1880
rect 670 1884 676 1885
rect 670 1880 671 1884
rect 675 1880 676 1884
rect 670 1879 676 1880
rect 726 1884 732 1885
rect 726 1880 727 1884
rect 731 1880 732 1884
rect 726 1879 732 1880
rect 782 1884 788 1885
rect 782 1880 783 1884
rect 787 1880 788 1884
rect 782 1879 788 1880
rect 846 1884 852 1885
rect 846 1880 847 1884
rect 851 1880 852 1884
rect 1094 1883 1095 1887
rect 1099 1883 1100 1887
rect 1094 1882 1100 1883
rect 1535 1887 1541 1888
rect 1535 1883 1536 1887
rect 1540 1886 1541 1887
rect 1540 1884 1922 1886
rect 1540 1883 1541 1884
rect 1535 1882 1541 1883
rect 1920 1880 1922 1884
rect 846 1879 852 1880
rect 1183 1879 1189 1880
rect 1183 1875 1184 1879
rect 1188 1878 1189 1879
rect 1214 1879 1220 1880
rect 1214 1878 1215 1879
rect 1188 1876 1215 1878
rect 1188 1875 1189 1876
rect 1183 1874 1189 1875
rect 1214 1875 1215 1876
rect 1219 1875 1220 1879
rect 1214 1874 1220 1875
rect 1223 1879 1229 1880
rect 1223 1875 1224 1879
rect 1228 1878 1229 1879
rect 1278 1879 1284 1880
rect 1278 1878 1279 1879
rect 1228 1876 1279 1878
rect 1228 1875 1229 1876
rect 1223 1874 1229 1875
rect 1278 1875 1279 1876
rect 1283 1875 1284 1879
rect 1278 1874 1284 1875
rect 1287 1879 1293 1880
rect 1287 1875 1288 1879
rect 1292 1878 1293 1879
rect 1318 1879 1324 1880
rect 1318 1878 1319 1879
rect 1292 1876 1319 1878
rect 1292 1875 1293 1876
rect 1287 1874 1293 1875
rect 1318 1875 1319 1876
rect 1323 1875 1324 1879
rect 1318 1874 1324 1875
rect 1351 1879 1357 1880
rect 1351 1875 1352 1879
rect 1356 1878 1357 1879
rect 1406 1879 1412 1880
rect 1406 1878 1407 1879
rect 1356 1876 1407 1878
rect 1356 1875 1357 1876
rect 1351 1874 1357 1875
rect 1406 1875 1407 1876
rect 1411 1875 1412 1879
rect 1406 1874 1412 1875
rect 1415 1879 1421 1880
rect 1415 1875 1416 1879
rect 1420 1878 1421 1879
rect 1462 1879 1468 1880
rect 1462 1878 1463 1879
rect 1420 1876 1463 1878
rect 1420 1875 1421 1876
rect 1415 1874 1421 1875
rect 1462 1875 1463 1876
rect 1467 1875 1468 1879
rect 1462 1874 1468 1875
rect 1471 1879 1480 1880
rect 1471 1875 1472 1879
rect 1479 1875 1480 1879
rect 1471 1874 1480 1875
rect 1527 1879 1533 1880
rect 1527 1875 1528 1879
rect 1532 1878 1533 1879
rect 1574 1879 1580 1880
rect 1574 1878 1575 1879
rect 1532 1876 1575 1878
rect 1532 1875 1533 1876
rect 1527 1874 1533 1875
rect 1574 1875 1575 1876
rect 1579 1875 1580 1879
rect 1574 1874 1580 1875
rect 1583 1879 1589 1880
rect 1583 1875 1584 1879
rect 1588 1878 1589 1879
rect 1646 1879 1652 1880
rect 1646 1878 1647 1879
rect 1588 1876 1647 1878
rect 1588 1875 1589 1876
rect 1583 1874 1589 1875
rect 1646 1875 1647 1876
rect 1651 1875 1652 1879
rect 1646 1874 1652 1875
rect 1655 1879 1661 1880
rect 1655 1875 1656 1879
rect 1660 1878 1661 1879
rect 1670 1879 1676 1880
rect 1670 1878 1671 1879
rect 1660 1876 1671 1878
rect 1660 1875 1661 1876
rect 1655 1874 1661 1875
rect 1670 1875 1671 1876
rect 1675 1875 1676 1879
rect 1670 1874 1676 1875
rect 1735 1879 1741 1880
rect 1735 1875 1736 1879
rect 1740 1878 1741 1879
rect 1814 1879 1820 1880
rect 1814 1878 1815 1879
rect 1740 1876 1815 1878
rect 1740 1875 1741 1876
rect 1735 1874 1741 1875
rect 1814 1875 1815 1876
rect 1819 1875 1820 1879
rect 1814 1874 1820 1875
rect 1823 1879 1829 1880
rect 1823 1875 1824 1879
rect 1828 1878 1829 1879
rect 1910 1879 1916 1880
rect 1910 1878 1911 1879
rect 1828 1876 1911 1878
rect 1828 1875 1829 1876
rect 1823 1874 1829 1875
rect 1910 1875 1911 1876
rect 1915 1875 1916 1879
rect 1910 1874 1916 1875
rect 1919 1879 1925 1880
rect 1919 1875 1920 1879
rect 1924 1875 1925 1879
rect 1919 1874 1925 1875
rect 2015 1879 2021 1880
rect 2015 1875 2016 1879
rect 2020 1878 2021 1879
rect 2086 1879 2092 1880
rect 2086 1878 2087 1879
rect 2020 1876 2087 1878
rect 2020 1875 2021 1876
rect 2015 1874 2021 1875
rect 2086 1875 2087 1876
rect 2091 1875 2092 1879
rect 2086 1874 2092 1875
rect 2094 1879 2101 1880
rect 2094 1875 2095 1879
rect 2100 1875 2101 1879
rect 2094 1874 2101 1875
rect 1158 1872 1164 1873
rect 134 1868 140 1869
rect 110 1865 116 1866
rect 110 1861 111 1865
rect 115 1861 116 1865
rect 134 1864 135 1868
rect 139 1864 140 1868
rect 134 1863 140 1864
rect 198 1868 204 1869
rect 198 1864 199 1868
rect 203 1864 204 1868
rect 198 1863 204 1864
rect 270 1868 276 1869
rect 270 1864 271 1868
rect 275 1864 276 1868
rect 270 1863 276 1864
rect 334 1868 340 1869
rect 334 1864 335 1868
rect 339 1864 340 1868
rect 334 1863 340 1864
rect 398 1868 404 1869
rect 398 1864 399 1868
rect 403 1864 404 1868
rect 398 1863 404 1864
rect 454 1868 460 1869
rect 454 1864 455 1868
rect 459 1864 460 1868
rect 454 1863 460 1864
rect 502 1868 508 1869
rect 502 1864 503 1868
rect 507 1864 508 1868
rect 502 1863 508 1864
rect 550 1868 556 1869
rect 550 1864 551 1868
rect 555 1864 556 1868
rect 550 1863 556 1864
rect 598 1868 604 1869
rect 598 1864 599 1868
rect 603 1864 604 1868
rect 598 1863 604 1864
rect 646 1868 652 1869
rect 646 1864 647 1868
rect 651 1864 652 1868
rect 646 1863 652 1864
rect 694 1868 700 1869
rect 694 1864 695 1868
rect 699 1864 700 1868
rect 694 1863 700 1864
rect 750 1868 756 1869
rect 750 1864 751 1868
rect 755 1864 756 1868
rect 1158 1868 1159 1872
rect 1163 1868 1164 1872
rect 1158 1867 1164 1868
rect 1198 1872 1204 1873
rect 1198 1868 1199 1872
rect 1203 1868 1204 1872
rect 1198 1867 1204 1868
rect 1262 1872 1268 1873
rect 1262 1868 1263 1872
rect 1267 1868 1268 1872
rect 1262 1867 1268 1868
rect 1326 1872 1332 1873
rect 1326 1868 1327 1872
rect 1331 1868 1332 1872
rect 1326 1867 1332 1868
rect 1390 1872 1396 1873
rect 1390 1868 1391 1872
rect 1395 1868 1396 1872
rect 1390 1867 1396 1868
rect 1446 1872 1452 1873
rect 1446 1868 1447 1872
rect 1451 1868 1452 1872
rect 1446 1867 1452 1868
rect 1502 1872 1508 1873
rect 1502 1868 1503 1872
rect 1507 1868 1508 1872
rect 1502 1867 1508 1868
rect 1558 1872 1564 1873
rect 1558 1868 1559 1872
rect 1563 1868 1564 1872
rect 1558 1867 1564 1868
rect 1630 1872 1636 1873
rect 1630 1868 1631 1872
rect 1635 1868 1636 1872
rect 1630 1867 1636 1868
rect 1710 1872 1716 1873
rect 1710 1868 1711 1872
rect 1715 1868 1716 1872
rect 1710 1867 1716 1868
rect 1798 1872 1804 1873
rect 1798 1868 1799 1872
rect 1803 1868 1804 1872
rect 1798 1867 1804 1868
rect 1894 1872 1900 1873
rect 1894 1868 1895 1872
rect 1899 1868 1900 1872
rect 1894 1867 1900 1868
rect 1990 1872 1996 1873
rect 1990 1868 1991 1872
rect 1995 1868 1996 1872
rect 1990 1867 1996 1868
rect 2070 1872 2076 1873
rect 2070 1868 2071 1872
rect 2075 1868 2076 1872
rect 2070 1867 2076 1868
rect 750 1863 756 1864
rect 1094 1865 1100 1866
rect 110 1860 116 1861
rect 1094 1861 1095 1865
rect 1099 1861 1100 1865
rect 1094 1860 1100 1861
rect 1134 1864 1140 1865
rect 1134 1860 1135 1864
rect 1139 1860 1140 1864
rect 2118 1864 2124 1865
rect 2118 1860 2119 1864
rect 2123 1860 2124 1864
rect 294 1859 300 1860
rect 294 1858 295 1859
rect 200 1856 295 1858
rect 159 1851 165 1852
rect 110 1848 116 1849
rect 110 1844 111 1848
rect 115 1844 116 1848
rect 159 1847 160 1851
rect 164 1850 165 1851
rect 200 1850 202 1856
rect 294 1855 295 1856
rect 299 1855 300 1859
rect 478 1859 484 1860
rect 1134 1859 1140 1860
rect 1183 1859 1189 1860
rect 478 1858 479 1859
rect 294 1854 300 1855
rect 360 1856 479 1858
rect 360 1852 362 1856
rect 478 1855 479 1856
rect 483 1855 484 1859
rect 478 1854 484 1855
rect 1183 1855 1184 1859
rect 1188 1858 1189 1859
rect 1206 1859 1212 1860
rect 1206 1858 1207 1859
rect 1188 1856 1207 1858
rect 1188 1855 1189 1856
rect 1183 1854 1189 1855
rect 1206 1855 1207 1856
rect 1211 1855 1212 1859
rect 1206 1854 1212 1855
rect 1214 1859 1220 1860
rect 1214 1855 1215 1859
rect 1219 1858 1220 1859
rect 1223 1859 1229 1860
rect 1223 1858 1224 1859
rect 1219 1856 1224 1858
rect 1219 1855 1220 1856
rect 1214 1854 1220 1855
rect 1223 1855 1224 1856
rect 1228 1855 1229 1859
rect 1223 1854 1229 1855
rect 1278 1859 1284 1860
rect 1278 1855 1279 1859
rect 1283 1858 1284 1859
rect 1287 1859 1293 1860
rect 1287 1858 1288 1859
rect 1283 1856 1288 1858
rect 1283 1855 1284 1856
rect 1278 1854 1284 1855
rect 1287 1855 1288 1856
rect 1292 1855 1293 1859
rect 1287 1854 1293 1855
rect 1351 1859 1357 1860
rect 1351 1855 1352 1859
rect 1356 1858 1357 1859
rect 1398 1859 1404 1860
rect 1398 1858 1399 1859
rect 1356 1856 1399 1858
rect 1356 1855 1357 1856
rect 1351 1854 1357 1855
rect 1398 1855 1399 1856
rect 1403 1855 1404 1859
rect 1398 1854 1404 1855
rect 1406 1859 1412 1860
rect 1406 1855 1407 1859
rect 1411 1858 1412 1859
rect 1415 1859 1421 1860
rect 1415 1858 1416 1859
rect 1411 1856 1416 1858
rect 1411 1855 1412 1856
rect 1406 1854 1412 1855
rect 1415 1855 1416 1856
rect 1420 1855 1421 1859
rect 1415 1854 1421 1855
rect 1462 1859 1468 1860
rect 1462 1855 1463 1859
rect 1467 1858 1468 1859
rect 1471 1859 1477 1860
rect 1471 1858 1472 1859
rect 1467 1856 1472 1858
rect 1467 1855 1468 1856
rect 1462 1854 1468 1855
rect 1471 1855 1472 1856
rect 1476 1855 1477 1859
rect 1471 1854 1477 1855
rect 1527 1859 1533 1860
rect 1527 1855 1528 1859
rect 1532 1858 1533 1859
rect 1535 1859 1541 1860
rect 1535 1858 1536 1859
rect 1532 1856 1536 1858
rect 1532 1855 1533 1856
rect 1527 1854 1533 1855
rect 1535 1855 1536 1856
rect 1540 1855 1541 1859
rect 1535 1854 1541 1855
rect 1574 1859 1580 1860
rect 1574 1855 1575 1859
rect 1579 1858 1580 1859
rect 1583 1859 1589 1860
rect 1583 1858 1584 1859
rect 1579 1856 1584 1858
rect 1579 1855 1580 1856
rect 1574 1854 1580 1855
rect 1583 1855 1584 1856
rect 1588 1855 1589 1859
rect 1583 1854 1589 1855
rect 1646 1859 1652 1860
rect 1646 1855 1647 1859
rect 1651 1858 1652 1859
rect 1655 1859 1661 1860
rect 1655 1858 1656 1859
rect 1651 1856 1656 1858
rect 1651 1855 1652 1856
rect 1646 1854 1652 1855
rect 1655 1855 1656 1856
rect 1660 1855 1661 1859
rect 1655 1854 1661 1855
rect 1734 1859 1741 1860
rect 1734 1855 1735 1859
rect 1740 1855 1741 1859
rect 1734 1854 1741 1855
rect 1814 1859 1820 1860
rect 1814 1855 1815 1859
rect 1819 1858 1820 1859
rect 1823 1859 1829 1860
rect 1823 1858 1824 1859
rect 1819 1856 1824 1858
rect 1819 1855 1820 1856
rect 1814 1854 1820 1855
rect 1823 1855 1824 1856
rect 1828 1855 1829 1859
rect 1823 1854 1829 1855
rect 1910 1859 1916 1860
rect 1910 1855 1911 1859
rect 1915 1858 1916 1859
rect 1919 1859 1925 1860
rect 1919 1858 1920 1859
rect 1915 1856 1920 1858
rect 1915 1855 1916 1856
rect 1910 1854 1916 1855
rect 1919 1855 1920 1856
rect 1924 1855 1925 1859
rect 1919 1854 1925 1855
rect 2015 1859 2021 1860
rect 2015 1855 2016 1859
rect 2020 1858 2021 1859
rect 2078 1859 2084 1860
rect 2078 1858 2079 1859
rect 2020 1856 2079 1858
rect 2020 1855 2021 1856
rect 2015 1854 2021 1855
rect 2078 1855 2079 1856
rect 2083 1855 2084 1859
rect 2078 1854 2084 1855
rect 2086 1859 2092 1860
rect 2086 1855 2087 1859
rect 2091 1858 2092 1859
rect 2095 1859 2101 1860
rect 2118 1859 2124 1860
rect 2095 1858 2096 1859
rect 2091 1856 2096 1858
rect 2091 1855 2092 1856
rect 2086 1854 2092 1855
rect 2095 1855 2096 1856
rect 2100 1855 2101 1859
rect 2095 1854 2101 1855
rect 164 1848 202 1850
rect 206 1851 212 1852
rect 164 1847 165 1848
rect 159 1846 165 1847
rect 206 1847 207 1851
rect 211 1850 212 1851
rect 223 1851 229 1852
rect 223 1850 224 1851
rect 211 1848 224 1850
rect 211 1847 212 1848
rect 206 1846 212 1847
rect 223 1847 224 1848
rect 228 1847 229 1851
rect 223 1846 229 1847
rect 234 1851 240 1852
rect 234 1847 235 1851
rect 239 1850 240 1851
rect 295 1851 301 1852
rect 295 1850 296 1851
rect 239 1848 296 1850
rect 239 1847 240 1848
rect 234 1846 240 1847
rect 295 1847 296 1848
rect 300 1847 301 1851
rect 295 1846 301 1847
rect 359 1851 365 1852
rect 359 1847 360 1851
rect 364 1847 365 1851
rect 359 1846 365 1847
rect 367 1851 373 1852
rect 367 1847 368 1851
rect 372 1850 373 1851
rect 423 1851 429 1852
rect 423 1850 424 1851
rect 372 1848 424 1850
rect 372 1847 373 1848
rect 367 1846 373 1847
rect 423 1847 424 1848
rect 428 1847 429 1851
rect 423 1846 429 1847
rect 479 1851 485 1852
rect 479 1847 480 1851
rect 484 1850 485 1851
rect 510 1851 516 1852
rect 510 1850 511 1851
rect 484 1848 511 1850
rect 484 1847 485 1848
rect 479 1846 485 1847
rect 510 1847 511 1848
rect 515 1847 516 1851
rect 510 1846 516 1847
rect 518 1851 524 1852
rect 518 1847 519 1851
rect 523 1850 524 1851
rect 527 1851 533 1852
rect 527 1850 528 1851
rect 523 1848 528 1850
rect 523 1847 524 1848
rect 518 1846 524 1847
rect 527 1847 528 1848
rect 532 1847 533 1851
rect 527 1846 533 1847
rect 535 1851 541 1852
rect 535 1847 536 1851
rect 540 1850 541 1851
rect 575 1851 581 1852
rect 575 1850 576 1851
rect 540 1848 576 1850
rect 540 1847 541 1848
rect 535 1846 541 1847
rect 575 1847 576 1848
rect 580 1847 581 1851
rect 575 1846 581 1847
rect 583 1851 589 1852
rect 583 1847 584 1851
rect 588 1850 589 1851
rect 623 1851 629 1852
rect 623 1850 624 1851
rect 588 1848 624 1850
rect 588 1847 589 1848
rect 583 1846 589 1847
rect 623 1847 624 1848
rect 628 1847 629 1851
rect 623 1846 629 1847
rect 631 1851 637 1852
rect 631 1847 632 1851
rect 636 1850 637 1851
rect 671 1851 677 1852
rect 671 1850 672 1851
rect 636 1848 672 1850
rect 636 1847 637 1848
rect 631 1846 637 1847
rect 671 1847 672 1848
rect 676 1847 677 1851
rect 671 1846 677 1847
rect 679 1851 685 1852
rect 679 1847 680 1851
rect 684 1850 685 1851
rect 719 1851 725 1852
rect 719 1850 720 1851
rect 684 1848 720 1850
rect 684 1847 685 1848
rect 679 1846 685 1847
rect 719 1847 720 1848
rect 724 1847 725 1851
rect 719 1846 725 1847
rect 727 1851 733 1852
rect 727 1847 728 1851
rect 732 1850 733 1851
rect 775 1851 781 1852
rect 775 1850 776 1851
rect 732 1848 776 1850
rect 732 1847 733 1848
rect 727 1846 733 1847
rect 775 1847 776 1848
rect 780 1847 781 1851
rect 775 1846 781 1847
rect 1094 1848 1100 1849
rect 110 1843 116 1844
rect 1094 1844 1095 1848
rect 1099 1844 1100 1848
rect 1094 1843 1100 1844
rect 1134 1847 1140 1848
rect 1134 1843 1135 1847
rect 1139 1843 1140 1847
rect 2118 1847 2124 1848
rect 1134 1842 1140 1843
rect 1158 1844 1164 1845
rect 134 1840 140 1841
rect 134 1836 135 1840
rect 139 1836 140 1840
rect 134 1835 140 1836
rect 198 1840 204 1841
rect 198 1836 199 1840
rect 203 1836 204 1840
rect 198 1835 204 1836
rect 270 1840 276 1841
rect 270 1836 271 1840
rect 275 1836 276 1840
rect 270 1835 276 1836
rect 334 1840 340 1841
rect 334 1836 335 1840
rect 339 1836 340 1840
rect 334 1835 340 1836
rect 398 1840 404 1841
rect 398 1836 399 1840
rect 403 1836 404 1840
rect 398 1835 404 1836
rect 454 1840 460 1841
rect 454 1836 455 1840
rect 459 1836 460 1840
rect 454 1835 460 1836
rect 502 1840 508 1841
rect 502 1836 503 1840
rect 507 1836 508 1840
rect 502 1835 508 1836
rect 550 1840 556 1841
rect 550 1836 551 1840
rect 555 1836 556 1840
rect 550 1835 556 1836
rect 598 1840 604 1841
rect 598 1836 599 1840
rect 603 1836 604 1840
rect 598 1835 604 1836
rect 646 1840 652 1841
rect 646 1836 647 1840
rect 651 1836 652 1840
rect 646 1835 652 1836
rect 694 1840 700 1841
rect 694 1836 695 1840
rect 699 1836 700 1840
rect 694 1835 700 1836
rect 750 1840 756 1841
rect 750 1836 751 1840
rect 755 1836 756 1840
rect 1158 1840 1159 1844
rect 1163 1840 1164 1844
rect 1158 1839 1164 1840
rect 1198 1844 1204 1845
rect 1198 1840 1199 1844
rect 1203 1840 1204 1844
rect 1198 1839 1204 1840
rect 1262 1844 1268 1845
rect 1262 1840 1263 1844
rect 1267 1840 1268 1844
rect 1262 1839 1268 1840
rect 1326 1844 1332 1845
rect 1326 1840 1327 1844
rect 1331 1840 1332 1844
rect 1326 1839 1332 1840
rect 1390 1844 1396 1845
rect 1390 1840 1391 1844
rect 1395 1840 1396 1844
rect 1390 1839 1396 1840
rect 1446 1844 1452 1845
rect 1446 1840 1447 1844
rect 1451 1840 1452 1844
rect 1446 1839 1452 1840
rect 1502 1844 1508 1845
rect 1502 1840 1503 1844
rect 1507 1840 1508 1844
rect 1502 1839 1508 1840
rect 1558 1844 1564 1845
rect 1558 1840 1559 1844
rect 1563 1840 1564 1844
rect 1558 1839 1564 1840
rect 1630 1844 1636 1845
rect 1630 1840 1631 1844
rect 1635 1840 1636 1844
rect 1630 1839 1636 1840
rect 1710 1844 1716 1845
rect 1710 1840 1711 1844
rect 1715 1840 1716 1844
rect 1710 1839 1716 1840
rect 1798 1844 1804 1845
rect 1798 1840 1799 1844
rect 1803 1840 1804 1844
rect 1798 1839 1804 1840
rect 1894 1844 1900 1845
rect 1894 1840 1895 1844
rect 1899 1840 1900 1844
rect 1894 1839 1900 1840
rect 1990 1844 1996 1845
rect 1990 1840 1991 1844
rect 1995 1840 1996 1844
rect 1990 1839 1996 1840
rect 2070 1844 2076 1845
rect 2070 1840 2071 1844
rect 2075 1840 2076 1844
rect 2118 1843 2119 1847
rect 2123 1843 2124 1847
rect 2118 1842 2124 1843
rect 2070 1839 2076 1840
rect 750 1835 756 1836
rect 1158 1832 1164 1833
rect 158 1831 165 1832
rect 158 1827 159 1831
rect 164 1827 165 1831
rect 158 1826 165 1827
rect 223 1831 229 1832
rect 223 1827 224 1831
rect 228 1830 229 1831
rect 234 1831 240 1832
rect 234 1830 235 1831
rect 228 1828 235 1830
rect 228 1827 229 1828
rect 223 1826 229 1827
rect 234 1827 235 1828
rect 239 1827 240 1831
rect 234 1826 240 1827
rect 294 1831 301 1832
rect 294 1827 295 1831
rect 300 1827 301 1831
rect 294 1826 301 1827
rect 359 1831 365 1832
rect 359 1827 360 1831
rect 364 1830 365 1831
rect 367 1831 373 1832
rect 367 1830 368 1831
rect 364 1828 368 1830
rect 364 1827 365 1828
rect 359 1826 365 1827
rect 367 1827 368 1828
rect 372 1827 373 1831
rect 367 1826 373 1827
rect 423 1831 429 1832
rect 423 1827 424 1831
rect 428 1830 429 1831
rect 438 1831 444 1832
rect 438 1830 439 1831
rect 428 1828 439 1830
rect 428 1827 429 1828
rect 423 1826 429 1827
rect 438 1827 439 1828
rect 443 1827 444 1831
rect 438 1826 444 1827
rect 478 1831 485 1832
rect 478 1827 479 1831
rect 484 1827 485 1831
rect 478 1826 485 1827
rect 527 1831 533 1832
rect 527 1827 528 1831
rect 532 1830 533 1831
rect 535 1831 541 1832
rect 535 1830 536 1831
rect 532 1828 536 1830
rect 532 1827 533 1828
rect 527 1826 533 1827
rect 535 1827 536 1828
rect 540 1827 541 1831
rect 535 1826 541 1827
rect 575 1831 581 1832
rect 575 1827 576 1831
rect 580 1830 581 1831
rect 583 1831 589 1832
rect 583 1830 584 1831
rect 580 1828 584 1830
rect 580 1827 581 1828
rect 575 1826 581 1827
rect 583 1827 584 1828
rect 588 1827 589 1831
rect 583 1826 589 1827
rect 623 1831 629 1832
rect 623 1827 624 1831
rect 628 1830 629 1831
rect 631 1831 637 1832
rect 631 1830 632 1831
rect 628 1828 632 1830
rect 628 1827 629 1828
rect 623 1826 629 1827
rect 631 1827 632 1828
rect 636 1827 637 1831
rect 631 1826 637 1827
rect 671 1831 677 1832
rect 671 1827 672 1831
rect 676 1830 677 1831
rect 679 1831 685 1832
rect 679 1830 680 1831
rect 676 1828 680 1830
rect 676 1827 677 1828
rect 671 1826 677 1827
rect 679 1827 680 1828
rect 684 1827 685 1831
rect 679 1826 685 1827
rect 719 1831 725 1832
rect 719 1827 720 1831
rect 724 1830 725 1831
rect 727 1831 733 1832
rect 727 1830 728 1831
rect 724 1828 728 1830
rect 724 1827 725 1828
rect 719 1826 725 1827
rect 727 1827 728 1828
rect 732 1827 733 1831
rect 775 1831 781 1832
rect 775 1830 776 1831
rect 727 1826 733 1827
rect 736 1828 776 1830
rect 622 1823 628 1824
rect 622 1819 623 1823
rect 627 1822 628 1823
rect 736 1822 738 1828
rect 775 1827 776 1828
rect 780 1827 781 1831
rect 775 1826 781 1827
rect 1134 1829 1140 1830
rect 1134 1825 1135 1829
rect 1139 1825 1140 1829
rect 1158 1828 1159 1832
rect 1163 1828 1164 1832
rect 1158 1827 1164 1828
rect 1230 1832 1236 1833
rect 1230 1828 1231 1832
rect 1235 1828 1236 1832
rect 1230 1827 1236 1828
rect 1302 1832 1308 1833
rect 1302 1828 1303 1832
rect 1307 1828 1308 1832
rect 1302 1827 1308 1828
rect 1382 1832 1388 1833
rect 1382 1828 1383 1832
rect 1387 1828 1388 1832
rect 1382 1827 1388 1828
rect 1462 1832 1468 1833
rect 1462 1828 1463 1832
rect 1467 1828 1468 1832
rect 1462 1827 1468 1828
rect 1550 1832 1556 1833
rect 1550 1828 1551 1832
rect 1555 1828 1556 1832
rect 1550 1827 1556 1828
rect 1646 1832 1652 1833
rect 1646 1828 1647 1832
rect 1651 1828 1652 1832
rect 1646 1827 1652 1828
rect 1750 1832 1756 1833
rect 1750 1828 1751 1832
rect 1755 1828 1756 1832
rect 1750 1827 1756 1828
rect 1854 1832 1860 1833
rect 1854 1828 1855 1832
rect 1859 1828 1860 1832
rect 1854 1827 1860 1828
rect 1966 1832 1972 1833
rect 1966 1828 1967 1832
rect 1971 1828 1972 1832
rect 1966 1827 1972 1828
rect 2070 1832 2076 1833
rect 2070 1828 2071 1832
rect 2075 1828 2076 1832
rect 2070 1827 2076 1828
rect 2118 1829 2124 1830
rect 1134 1824 1140 1825
rect 2118 1825 2119 1829
rect 2123 1825 2124 1829
rect 2118 1824 2124 1825
rect 627 1820 738 1822
rect 627 1819 628 1820
rect 622 1818 628 1819
rect 1183 1815 1189 1816
rect 1134 1812 1140 1813
rect 518 1811 524 1812
rect 518 1807 519 1811
rect 523 1810 524 1811
rect 523 1808 651 1810
rect 523 1807 524 1808
rect 518 1806 524 1807
rect 649 1804 651 1808
rect 1134 1808 1135 1812
rect 1139 1808 1140 1812
rect 1183 1811 1184 1815
rect 1188 1814 1189 1815
rect 1246 1815 1252 1816
rect 1246 1814 1247 1815
rect 1188 1812 1247 1814
rect 1188 1811 1189 1812
rect 1183 1810 1189 1811
rect 1246 1811 1247 1812
rect 1251 1811 1252 1815
rect 1246 1810 1252 1811
rect 1255 1815 1261 1816
rect 1255 1811 1256 1815
rect 1260 1814 1261 1815
rect 1310 1815 1316 1816
rect 1310 1814 1311 1815
rect 1260 1812 1311 1814
rect 1260 1811 1261 1812
rect 1255 1810 1261 1811
rect 1310 1811 1311 1812
rect 1315 1811 1316 1815
rect 1310 1810 1316 1811
rect 1318 1815 1324 1816
rect 1318 1811 1319 1815
rect 1323 1814 1324 1815
rect 1327 1815 1333 1816
rect 1327 1814 1328 1815
rect 1323 1812 1328 1814
rect 1323 1811 1324 1812
rect 1318 1810 1324 1811
rect 1327 1811 1328 1812
rect 1332 1811 1333 1815
rect 1327 1810 1333 1811
rect 1407 1815 1413 1816
rect 1407 1811 1408 1815
rect 1412 1814 1413 1815
rect 1478 1815 1484 1816
rect 1478 1814 1479 1815
rect 1412 1812 1479 1814
rect 1412 1811 1413 1812
rect 1407 1810 1413 1811
rect 1478 1811 1479 1812
rect 1483 1811 1484 1815
rect 1478 1810 1484 1811
rect 1487 1815 1493 1816
rect 1487 1811 1488 1815
rect 1492 1814 1493 1815
rect 1558 1815 1564 1816
rect 1558 1814 1559 1815
rect 1492 1812 1559 1814
rect 1492 1811 1493 1812
rect 1487 1810 1493 1811
rect 1558 1811 1559 1812
rect 1563 1811 1564 1815
rect 1558 1810 1564 1811
rect 1566 1815 1572 1816
rect 1566 1811 1567 1815
rect 1571 1814 1572 1815
rect 1575 1815 1581 1816
rect 1575 1814 1576 1815
rect 1571 1812 1576 1814
rect 1571 1811 1572 1812
rect 1566 1810 1572 1811
rect 1575 1811 1576 1812
rect 1580 1811 1581 1815
rect 1575 1810 1581 1811
rect 1670 1815 1677 1816
rect 1670 1811 1671 1815
rect 1676 1811 1677 1815
rect 1670 1810 1677 1811
rect 1679 1815 1685 1816
rect 1679 1811 1680 1815
rect 1684 1814 1685 1815
rect 1775 1815 1781 1816
rect 1775 1814 1776 1815
rect 1684 1812 1776 1814
rect 1684 1811 1685 1812
rect 1679 1810 1685 1811
rect 1775 1811 1776 1812
rect 1780 1811 1781 1815
rect 1775 1810 1781 1811
rect 1879 1815 1885 1816
rect 1879 1811 1880 1815
rect 1884 1814 1885 1815
rect 1950 1815 1956 1816
rect 1950 1814 1951 1815
rect 1884 1812 1951 1814
rect 1884 1811 1885 1812
rect 1879 1810 1885 1811
rect 1950 1811 1951 1812
rect 1955 1811 1956 1815
rect 1950 1810 1956 1811
rect 1958 1815 1964 1816
rect 1958 1811 1959 1815
rect 1963 1814 1964 1815
rect 1991 1815 1997 1816
rect 1991 1814 1992 1815
rect 1963 1812 1992 1814
rect 1963 1811 1964 1812
rect 1958 1810 1964 1811
rect 1991 1811 1992 1812
rect 1996 1811 1997 1815
rect 1991 1810 1997 1811
rect 2094 1815 2101 1816
rect 2094 1811 2095 1815
rect 2100 1811 2101 1815
rect 2094 1810 2101 1811
rect 2118 1812 2124 1813
rect 1134 1807 1140 1808
rect 2118 1808 2119 1812
rect 2123 1808 2124 1812
rect 2118 1807 2124 1808
rect 1158 1804 1164 1805
rect 175 1803 181 1804
rect 175 1799 176 1803
rect 180 1802 181 1803
rect 206 1803 212 1804
rect 206 1802 207 1803
rect 180 1800 207 1802
rect 180 1799 181 1800
rect 175 1798 181 1799
rect 206 1799 207 1800
rect 211 1799 212 1803
rect 206 1798 212 1799
rect 222 1803 228 1804
rect 222 1799 223 1803
rect 227 1802 228 1803
rect 239 1803 245 1804
rect 239 1802 240 1803
rect 227 1800 240 1802
rect 227 1799 228 1800
rect 222 1798 228 1799
rect 239 1799 240 1800
rect 244 1799 245 1803
rect 239 1798 245 1799
rect 247 1803 253 1804
rect 247 1799 248 1803
rect 252 1802 253 1803
rect 295 1803 301 1804
rect 295 1802 296 1803
rect 252 1800 296 1802
rect 252 1799 253 1800
rect 247 1798 253 1799
rect 295 1799 296 1800
rect 300 1799 301 1803
rect 295 1798 301 1799
rect 351 1803 357 1804
rect 351 1799 352 1803
rect 356 1802 357 1803
rect 374 1803 380 1804
rect 374 1802 375 1803
rect 356 1800 375 1802
rect 356 1799 357 1800
rect 351 1798 357 1799
rect 374 1799 375 1800
rect 379 1799 380 1803
rect 374 1798 380 1799
rect 390 1803 396 1804
rect 390 1799 391 1803
rect 395 1802 396 1803
rect 407 1803 413 1804
rect 407 1802 408 1803
rect 395 1800 408 1802
rect 395 1799 396 1800
rect 390 1798 396 1799
rect 407 1799 408 1800
rect 412 1799 413 1803
rect 407 1798 413 1799
rect 415 1803 421 1804
rect 415 1799 416 1803
rect 420 1802 421 1803
rect 455 1803 461 1804
rect 455 1802 456 1803
rect 420 1800 456 1802
rect 420 1799 421 1800
rect 415 1798 421 1799
rect 455 1799 456 1800
rect 460 1799 461 1803
rect 455 1798 461 1799
rect 503 1803 509 1804
rect 503 1799 504 1803
rect 508 1802 509 1803
rect 542 1803 548 1804
rect 542 1802 543 1803
rect 508 1800 543 1802
rect 508 1799 509 1800
rect 503 1798 509 1799
rect 542 1799 543 1800
rect 547 1799 548 1803
rect 542 1798 548 1799
rect 551 1803 557 1804
rect 551 1799 552 1803
rect 556 1802 557 1803
rect 590 1803 596 1804
rect 590 1802 591 1803
rect 556 1800 591 1802
rect 556 1799 557 1800
rect 551 1798 557 1799
rect 590 1799 591 1800
rect 595 1799 596 1803
rect 590 1798 596 1799
rect 599 1803 605 1804
rect 599 1799 600 1803
rect 604 1802 605 1803
rect 638 1803 644 1804
rect 638 1802 639 1803
rect 604 1800 639 1802
rect 604 1799 605 1800
rect 599 1798 605 1799
rect 638 1799 639 1800
rect 643 1799 644 1803
rect 638 1798 644 1799
rect 647 1803 653 1804
rect 647 1799 648 1803
rect 652 1799 653 1803
rect 695 1803 701 1804
rect 695 1802 696 1803
rect 647 1798 653 1799
rect 656 1800 696 1802
rect 150 1796 156 1797
rect 150 1792 151 1796
rect 155 1792 156 1796
rect 150 1791 156 1792
rect 214 1796 220 1797
rect 214 1792 215 1796
rect 219 1792 220 1796
rect 214 1791 220 1792
rect 270 1796 276 1797
rect 270 1792 271 1796
rect 275 1792 276 1796
rect 270 1791 276 1792
rect 326 1796 332 1797
rect 326 1792 327 1796
rect 331 1792 332 1796
rect 326 1791 332 1792
rect 382 1796 388 1797
rect 382 1792 383 1796
rect 387 1792 388 1796
rect 382 1791 388 1792
rect 430 1796 436 1797
rect 430 1792 431 1796
rect 435 1792 436 1796
rect 430 1791 436 1792
rect 478 1796 484 1797
rect 478 1792 479 1796
rect 483 1792 484 1796
rect 478 1791 484 1792
rect 526 1796 532 1797
rect 526 1792 527 1796
rect 531 1792 532 1796
rect 526 1791 532 1792
rect 574 1796 580 1797
rect 574 1792 575 1796
rect 579 1792 580 1796
rect 574 1791 580 1792
rect 622 1796 628 1797
rect 622 1792 623 1796
rect 627 1792 628 1796
rect 622 1791 628 1792
rect 656 1790 658 1800
rect 695 1799 696 1800
rect 700 1799 701 1803
rect 695 1798 701 1799
rect 718 1803 724 1804
rect 718 1799 719 1803
rect 723 1802 724 1803
rect 751 1803 757 1804
rect 751 1802 752 1803
rect 723 1800 752 1802
rect 723 1799 724 1800
rect 718 1798 724 1799
rect 751 1799 752 1800
rect 756 1799 757 1803
rect 1158 1800 1159 1804
rect 1163 1800 1164 1804
rect 1158 1799 1164 1800
rect 1230 1804 1236 1805
rect 1230 1800 1231 1804
rect 1235 1800 1236 1804
rect 1230 1799 1236 1800
rect 1302 1804 1308 1805
rect 1302 1800 1303 1804
rect 1307 1800 1308 1804
rect 1302 1799 1308 1800
rect 1382 1804 1388 1805
rect 1382 1800 1383 1804
rect 1387 1800 1388 1804
rect 1382 1799 1388 1800
rect 1462 1804 1468 1805
rect 1462 1800 1463 1804
rect 1467 1800 1468 1804
rect 1462 1799 1468 1800
rect 1550 1804 1556 1805
rect 1550 1800 1551 1804
rect 1555 1800 1556 1804
rect 1550 1799 1556 1800
rect 1646 1804 1652 1805
rect 1646 1800 1647 1804
rect 1651 1800 1652 1804
rect 1646 1799 1652 1800
rect 1750 1804 1756 1805
rect 1750 1800 1751 1804
rect 1755 1800 1756 1804
rect 1750 1799 1756 1800
rect 1854 1804 1860 1805
rect 1854 1800 1855 1804
rect 1859 1800 1860 1804
rect 1854 1799 1860 1800
rect 1966 1804 1972 1805
rect 1966 1800 1967 1804
rect 1971 1800 1972 1804
rect 1966 1799 1972 1800
rect 2070 1804 2076 1805
rect 2070 1800 2071 1804
rect 2075 1800 2076 1804
rect 2070 1799 2076 1800
rect 751 1798 757 1799
rect 670 1796 676 1797
rect 670 1792 671 1796
rect 675 1792 676 1796
rect 670 1791 676 1792
rect 726 1796 732 1797
rect 726 1792 727 1796
rect 731 1792 732 1796
rect 726 1791 732 1792
rect 1183 1795 1189 1796
rect 1183 1791 1184 1795
rect 1188 1794 1189 1795
rect 1214 1795 1220 1796
rect 1214 1794 1215 1795
rect 1188 1792 1215 1794
rect 1188 1791 1189 1792
rect 1183 1790 1189 1791
rect 1214 1791 1215 1792
rect 1219 1791 1220 1795
rect 1214 1790 1220 1791
rect 1246 1795 1252 1796
rect 1246 1791 1247 1795
rect 1251 1794 1252 1795
rect 1255 1795 1261 1796
rect 1255 1794 1256 1795
rect 1251 1792 1256 1794
rect 1251 1791 1252 1792
rect 1246 1790 1252 1791
rect 1255 1791 1256 1792
rect 1260 1791 1261 1795
rect 1255 1790 1261 1791
rect 1310 1795 1316 1796
rect 1310 1791 1311 1795
rect 1315 1794 1316 1795
rect 1327 1795 1333 1796
rect 1327 1794 1328 1795
rect 1315 1792 1328 1794
rect 1315 1791 1316 1792
rect 1310 1790 1316 1791
rect 1327 1791 1328 1792
rect 1332 1791 1333 1795
rect 1327 1790 1333 1791
rect 1398 1795 1404 1796
rect 1398 1791 1399 1795
rect 1403 1794 1404 1795
rect 1407 1795 1413 1796
rect 1407 1794 1408 1795
rect 1403 1792 1408 1794
rect 1403 1791 1404 1792
rect 1398 1790 1404 1791
rect 1407 1791 1408 1792
rect 1412 1791 1413 1795
rect 1407 1790 1413 1791
rect 1478 1795 1484 1796
rect 1478 1791 1479 1795
rect 1483 1794 1484 1795
rect 1487 1795 1493 1796
rect 1487 1794 1488 1795
rect 1483 1792 1488 1794
rect 1483 1791 1484 1792
rect 1478 1790 1484 1791
rect 1487 1791 1488 1792
rect 1492 1791 1493 1795
rect 1487 1790 1493 1791
rect 1558 1795 1564 1796
rect 1558 1791 1559 1795
rect 1563 1794 1564 1795
rect 1575 1795 1581 1796
rect 1575 1794 1576 1795
rect 1563 1792 1576 1794
rect 1563 1791 1564 1792
rect 1558 1790 1564 1791
rect 1575 1791 1576 1792
rect 1580 1791 1581 1795
rect 1575 1790 1581 1791
rect 1671 1795 1677 1796
rect 1671 1791 1672 1795
rect 1676 1794 1677 1795
rect 1679 1795 1685 1796
rect 1679 1794 1680 1795
rect 1676 1792 1680 1794
rect 1676 1791 1677 1792
rect 1671 1790 1677 1791
rect 1679 1791 1680 1792
rect 1684 1791 1685 1795
rect 1679 1790 1685 1791
rect 1714 1795 1720 1796
rect 1714 1791 1715 1795
rect 1719 1794 1720 1795
rect 1775 1795 1781 1796
rect 1775 1794 1776 1795
rect 1719 1792 1776 1794
rect 1719 1791 1720 1792
rect 1714 1790 1720 1791
rect 1775 1791 1776 1792
rect 1780 1791 1781 1795
rect 1775 1790 1781 1791
rect 1879 1795 1885 1796
rect 1879 1791 1880 1795
rect 1884 1794 1885 1795
rect 1958 1795 1964 1796
rect 1958 1794 1959 1795
rect 1884 1792 1959 1794
rect 1884 1791 1885 1792
rect 1879 1790 1885 1791
rect 1958 1791 1959 1792
rect 1963 1791 1964 1795
rect 1958 1790 1964 1791
rect 1991 1795 1997 1796
rect 1991 1791 1992 1795
rect 1996 1794 1997 1795
rect 2030 1795 2036 1796
rect 2030 1794 2031 1795
rect 1996 1792 2031 1794
rect 1996 1791 1997 1792
rect 1991 1790 1997 1791
rect 2030 1791 2031 1792
rect 2035 1791 2036 1795
rect 2030 1790 2036 1791
rect 2078 1795 2084 1796
rect 2078 1791 2079 1795
rect 2083 1794 2084 1795
rect 2095 1795 2101 1796
rect 2095 1794 2096 1795
rect 2083 1792 2096 1794
rect 2083 1791 2084 1792
rect 2078 1790 2084 1791
rect 2095 1791 2096 1792
rect 2100 1791 2101 1795
rect 2095 1790 2101 1791
rect 110 1788 116 1789
rect 110 1784 111 1788
rect 115 1784 116 1788
rect 536 1788 562 1790
rect 110 1783 116 1784
rect 175 1783 181 1784
rect 175 1779 176 1783
rect 180 1782 181 1783
rect 222 1783 228 1784
rect 222 1782 223 1783
rect 180 1780 223 1782
rect 180 1779 181 1780
rect 175 1778 181 1779
rect 222 1779 223 1780
rect 227 1779 228 1783
rect 222 1778 228 1779
rect 239 1783 245 1784
rect 239 1779 240 1783
rect 244 1782 245 1783
rect 247 1783 253 1784
rect 247 1782 248 1783
rect 244 1780 248 1782
rect 244 1779 245 1780
rect 239 1778 245 1779
rect 247 1779 248 1780
rect 252 1779 253 1783
rect 247 1778 253 1779
rect 258 1783 264 1784
rect 258 1779 259 1783
rect 263 1782 264 1783
rect 295 1783 301 1784
rect 295 1782 296 1783
rect 263 1780 296 1782
rect 263 1779 264 1780
rect 258 1778 264 1779
rect 295 1779 296 1780
rect 300 1779 301 1783
rect 295 1778 301 1779
rect 351 1783 357 1784
rect 351 1779 352 1783
rect 356 1782 357 1783
rect 390 1783 396 1784
rect 390 1782 391 1783
rect 356 1780 391 1782
rect 356 1779 357 1780
rect 351 1778 357 1779
rect 390 1779 391 1780
rect 395 1779 396 1783
rect 390 1778 396 1779
rect 407 1783 413 1784
rect 407 1779 408 1783
rect 412 1782 413 1783
rect 415 1783 421 1784
rect 415 1782 416 1783
rect 412 1780 416 1782
rect 412 1779 413 1780
rect 407 1778 413 1779
rect 415 1779 416 1780
rect 420 1779 421 1783
rect 415 1778 421 1779
rect 438 1783 444 1784
rect 438 1779 439 1783
rect 443 1782 444 1783
rect 455 1783 461 1784
rect 455 1782 456 1783
rect 443 1780 456 1782
rect 443 1779 444 1780
rect 438 1778 444 1779
rect 455 1779 456 1780
rect 460 1779 461 1783
rect 455 1778 461 1779
rect 503 1783 509 1784
rect 503 1779 504 1783
rect 508 1782 509 1783
rect 536 1782 538 1788
rect 560 1786 562 1788
rect 584 1788 610 1790
rect 584 1786 586 1788
rect 560 1784 586 1786
rect 608 1786 610 1788
rect 632 1788 658 1790
rect 1094 1788 1100 1789
rect 632 1786 634 1788
rect 608 1784 634 1786
rect 1094 1784 1095 1788
rect 1099 1784 1100 1788
rect 508 1780 538 1782
rect 542 1783 548 1784
rect 508 1779 509 1780
rect 503 1778 509 1779
rect 542 1779 543 1783
rect 547 1782 548 1783
rect 551 1783 557 1784
rect 551 1782 552 1783
rect 547 1780 552 1782
rect 547 1779 548 1780
rect 542 1778 548 1779
rect 551 1779 552 1780
rect 556 1779 557 1783
rect 551 1778 557 1779
rect 590 1783 596 1784
rect 590 1779 591 1783
rect 595 1782 596 1783
rect 599 1783 605 1784
rect 599 1782 600 1783
rect 595 1780 600 1782
rect 595 1779 596 1780
rect 590 1778 596 1779
rect 599 1779 600 1780
rect 604 1779 605 1783
rect 599 1778 605 1779
rect 638 1783 644 1784
rect 638 1779 639 1783
rect 643 1782 644 1783
rect 647 1783 653 1784
rect 647 1782 648 1783
rect 643 1780 648 1782
rect 643 1779 644 1780
rect 638 1778 644 1779
rect 647 1779 648 1780
rect 652 1779 653 1783
rect 647 1778 653 1779
rect 695 1783 701 1784
rect 695 1779 696 1783
rect 700 1782 701 1783
rect 718 1783 724 1784
rect 718 1782 719 1783
rect 700 1780 719 1782
rect 700 1779 701 1780
rect 695 1778 701 1779
rect 718 1779 719 1780
rect 723 1779 724 1783
rect 718 1778 724 1779
rect 751 1783 757 1784
rect 751 1779 752 1783
rect 756 1782 757 1783
rect 782 1783 788 1784
rect 1094 1783 1100 1784
rect 782 1782 783 1783
rect 756 1780 783 1782
rect 756 1779 757 1780
rect 751 1778 757 1779
rect 782 1779 783 1780
rect 787 1779 788 1783
rect 782 1778 788 1779
rect 1566 1779 1572 1780
rect 1566 1778 1567 1779
rect 1551 1777 1567 1778
rect 1215 1775 1221 1776
rect 110 1771 116 1772
rect 110 1767 111 1771
rect 115 1767 116 1771
rect 1094 1771 1100 1772
rect 110 1766 116 1767
rect 150 1768 156 1769
rect 150 1764 151 1768
rect 155 1764 156 1768
rect 150 1763 156 1764
rect 214 1768 220 1769
rect 214 1764 215 1768
rect 219 1764 220 1768
rect 214 1763 220 1764
rect 270 1768 276 1769
rect 270 1764 271 1768
rect 275 1764 276 1768
rect 270 1763 276 1764
rect 326 1768 332 1769
rect 326 1764 327 1768
rect 331 1764 332 1768
rect 326 1763 332 1764
rect 382 1768 388 1769
rect 382 1764 383 1768
rect 387 1764 388 1768
rect 382 1763 388 1764
rect 430 1768 436 1769
rect 430 1764 431 1768
rect 435 1764 436 1768
rect 430 1763 436 1764
rect 478 1768 484 1769
rect 478 1764 479 1768
rect 483 1764 484 1768
rect 478 1763 484 1764
rect 526 1768 532 1769
rect 526 1764 527 1768
rect 531 1764 532 1768
rect 526 1763 532 1764
rect 574 1768 580 1769
rect 574 1764 575 1768
rect 579 1764 580 1768
rect 574 1763 580 1764
rect 622 1768 628 1769
rect 622 1764 623 1768
rect 627 1764 628 1768
rect 622 1763 628 1764
rect 670 1768 676 1769
rect 670 1764 671 1768
rect 675 1764 676 1768
rect 670 1763 676 1764
rect 726 1768 732 1769
rect 726 1764 727 1768
rect 731 1764 732 1768
rect 1094 1767 1095 1771
rect 1099 1767 1100 1771
rect 1215 1771 1216 1775
rect 1220 1774 1221 1775
rect 1270 1775 1276 1776
rect 1270 1774 1271 1775
rect 1220 1772 1271 1774
rect 1220 1771 1221 1772
rect 1215 1770 1221 1771
rect 1270 1771 1271 1772
rect 1275 1771 1276 1775
rect 1270 1770 1276 1771
rect 1279 1775 1285 1776
rect 1279 1771 1280 1775
rect 1284 1774 1285 1775
rect 1334 1775 1340 1776
rect 1334 1774 1335 1775
rect 1284 1772 1335 1774
rect 1284 1771 1285 1772
rect 1279 1770 1285 1771
rect 1334 1771 1335 1772
rect 1339 1771 1340 1775
rect 1334 1770 1340 1771
rect 1343 1775 1349 1776
rect 1343 1771 1344 1775
rect 1348 1774 1349 1775
rect 1366 1775 1372 1776
rect 1366 1774 1367 1775
rect 1348 1772 1367 1774
rect 1348 1771 1349 1772
rect 1343 1770 1349 1771
rect 1366 1771 1367 1772
rect 1371 1771 1372 1775
rect 1366 1770 1372 1771
rect 1407 1775 1413 1776
rect 1407 1771 1408 1775
rect 1412 1774 1413 1775
rect 1470 1775 1476 1776
rect 1470 1774 1471 1775
rect 1412 1772 1471 1774
rect 1412 1771 1413 1772
rect 1407 1770 1413 1771
rect 1470 1771 1471 1772
rect 1475 1771 1476 1775
rect 1470 1770 1476 1771
rect 1479 1775 1485 1776
rect 1479 1771 1480 1775
rect 1484 1774 1485 1775
rect 1542 1775 1548 1776
rect 1542 1774 1543 1775
rect 1484 1772 1543 1774
rect 1484 1771 1485 1772
rect 1479 1770 1485 1771
rect 1542 1771 1543 1772
rect 1547 1771 1548 1775
rect 1551 1773 1552 1777
rect 1556 1776 1567 1777
rect 1556 1773 1557 1776
rect 1566 1775 1567 1776
rect 1571 1775 1572 1779
rect 1566 1774 1572 1775
rect 1631 1775 1637 1776
rect 1551 1772 1557 1773
rect 1542 1770 1548 1771
rect 1631 1771 1632 1775
rect 1636 1774 1637 1775
rect 1694 1775 1700 1776
rect 1694 1774 1695 1775
rect 1636 1772 1695 1774
rect 1636 1771 1637 1772
rect 1631 1770 1637 1771
rect 1694 1771 1695 1772
rect 1699 1771 1700 1775
rect 1694 1770 1700 1771
rect 1702 1775 1708 1776
rect 1702 1771 1703 1775
rect 1707 1774 1708 1775
rect 1711 1775 1717 1776
rect 1711 1774 1712 1775
rect 1707 1772 1712 1774
rect 1707 1771 1708 1772
rect 1702 1770 1708 1771
rect 1711 1771 1712 1772
rect 1716 1771 1717 1775
rect 1711 1770 1717 1771
rect 1791 1775 1797 1776
rect 1791 1771 1792 1775
rect 1796 1774 1797 1775
rect 1862 1775 1868 1776
rect 1862 1774 1863 1775
rect 1796 1772 1863 1774
rect 1796 1771 1797 1772
rect 1791 1770 1797 1771
rect 1862 1771 1863 1772
rect 1867 1771 1868 1775
rect 1862 1770 1868 1771
rect 1871 1775 1877 1776
rect 1871 1771 1872 1775
rect 1876 1774 1877 1775
rect 1942 1775 1948 1776
rect 1942 1774 1943 1775
rect 1876 1772 1943 1774
rect 1876 1771 1877 1772
rect 1871 1770 1877 1771
rect 1942 1771 1943 1772
rect 1947 1771 1948 1775
rect 1942 1770 1948 1771
rect 1950 1775 1957 1776
rect 1950 1771 1951 1775
rect 1956 1771 1957 1775
rect 1950 1770 1957 1771
rect 2014 1775 2020 1776
rect 2014 1771 2015 1775
rect 2019 1774 2020 1775
rect 2031 1775 2037 1776
rect 2031 1774 2032 1775
rect 2019 1772 2032 1774
rect 2019 1771 2020 1772
rect 2014 1770 2020 1771
rect 2031 1771 2032 1772
rect 2036 1771 2037 1775
rect 2031 1770 2037 1771
rect 2094 1775 2101 1776
rect 2094 1771 2095 1775
rect 2100 1771 2101 1775
rect 2094 1770 2101 1771
rect 1094 1766 1100 1767
rect 1190 1768 1196 1769
rect 726 1763 732 1764
rect 1190 1764 1191 1768
rect 1195 1764 1196 1768
rect 1190 1763 1196 1764
rect 1254 1768 1260 1769
rect 1254 1764 1255 1768
rect 1259 1764 1260 1768
rect 1254 1763 1260 1764
rect 1318 1768 1324 1769
rect 1318 1764 1319 1768
rect 1323 1764 1324 1768
rect 1318 1763 1324 1764
rect 1382 1768 1388 1769
rect 1382 1764 1383 1768
rect 1387 1764 1388 1768
rect 1382 1763 1388 1764
rect 1454 1768 1460 1769
rect 1454 1764 1455 1768
rect 1459 1764 1460 1768
rect 1454 1763 1460 1764
rect 1526 1768 1532 1769
rect 1526 1764 1527 1768
rect 1531 1764 1532 1768
rect 1526 1763 1532 1764
rect 1606 1768 1612 1769
rect 1606 1764 1607 1768
rect 1611 1764 1612 1768
rect 1606 1763 1612 1764
rect 1686 1768 1692 1769
rect 1686 1764 1687 1768
rect 1691 1764 1692 1768
rect 1686 1763 1692 1764
rect 1766 1768 1772 1769
rect 1766 1764 1767 1768
rect 1771 1764 1772 1768
rect 1766 1763 1772 1764
rect 1846 1768 1852 1769
rect 1846 1764 1847 1768
rect 1851 1764 1852 1768
rect 1846 1763 1852 1764
rect 1926 1768 1932 1769
rect 1926 1764 1927 1768
rect 1931 1764 1932 1768
rect 1926 1763 1932 1764
rect 2006 1768 2012 1769
rect 2006 1764 2007 1768
rect 2011 1764 2012 1768
rect 2006 1763 2012 1764
rect 2070 1768 2076 1769
rect 2070 1764 2071 1768
rect 2075 1764 2076 1768
rect 2070 1763 2076 1764
rect 1134 1760 1140 1761
rect 230 1756 236 1757
rect 110 1753 116 1754
rect 110 1749 111 1753
rect 115 1749 116 1753
rect 230 1752 231 1756
rect 235 1752 236 1756
rect 230 1751 236 1752
rect 294 1756 300 1757
rect 294 1752 295 1756
rect 299 1752 300 1756
rect 294 1751 300 1752
rect 350 1756 356 1757
rect 350 1752 351 1756
rect 355 1752 356 1756
rect 350 1751 356 1752
rect 414 1756 420 1757
rect 414 1752 415 1756
rect 419 1752 420 1756
rect 414 1751 420 1752
rect 478 1756 484 1757
rect 478 1752 479 1756
rect 483 1752 484 1756
rect 478 1751 484 1752
rect 542 1756 548 1757
rect 542 1752 543 1756
rect 547 1752 548 1756
rect 542 1751 548 1752
rect 614 1756 620 1757
rect 614 1752 615 1756
rect 619 1752 620 1756
rect 614 1751 620 1752
rect 686 1756 692 1757
rect 686 1752 687 1756
rect 691 1752 692 1756
rect 686 1751 692 1752
rect 758 1756 764 1757
rect 758 1752 759 1756
rect 763 1752 764 1756
rect 758 1751 764 1752
rect 830 1756 836 1757
rect 830 1752 831 1756
rect 835 1752 836 1756
rect 830 1751 836 1752
rect 910 1756 916 1757
rect 910 1752 911 1756
rect 915 1752 916 1756
rect 910 1751 916 1752
rect 990 1756 996 1757
rect 990 1752 991 1756
rect 995 1752 996 1756
rect 1134 1756 1135 1760
rect 1139 1756 1140 1760
rect 2118 1760 2124 1761
rect 2118 1756 2119 1760
rect 2123 1756 2124 1760
rect 1134 1755 1140 1756
rect 1214 1755 1221 1756
rect 990 1751 996 1752
rect 1094 1753 1100 1754
rect 110 1748 116 1749
rect 1094 1749 1095 1753
rect 1099 1749 1100 1753
rect 1214 1751 1215 1755
rect 1220 1751 1221 1755
rect 1214 1750 1221 1751
rect 1270 1755 1276 1756
rect 1270 1751 1271 1755
rect 1275 1754 1276 1755
rect 1279 1755 1285 1756
rect 1279 1754 1280 1755
rect 1275 1752 1280 1754
rect 1275 1751 1276 1752
rect 1270 1750 1276 1751
rect 1279 1751 1280 1752
rect 1284 1751 1285 1755
rect 1279 1750 1285 1751
rect 1334 1755 1340 1756
rect 1334 1751 1335 1755
rect 1339 1754 1340 1755
rect 1343 1755 1349 1756
rect 1343 1754 1344 1755
rect 1339 1752 1344 1754
rect 1339 1751 1340 1752
rect 1334 1750 1340 1751
rect 1343 1751 1344 1752
rect 1348 1751 1349 1755
rect 1343 1750 1349 1751
rect 1407 1755 1416 1756
rect 1407 1751 1408 1755
rect 1415 1751 1416 1755
rect 1407 1750 1416 1751
rect 1470 1755 1476 1756
rect 1470 1751 1471 1755
rect 1475 1754 1476 1755
rect 1479 1755 1485 1756
rect 1479 1754 1480 1755
rect 1475 1752 1480 1754
rect 1475 1751 1476 1752
rect 1470 1750 1476 1751
rect 1479 1751 1480 1752
rect 1484 1751 1485 1755
rect 1479 1750 1485 1751
rect 1542 1755 1548 1756
rect 1542 1751 1543 1755
rect 1547 1754 1548 1755
rect 1551 1755 1557 1756
rect 1551 1754 1552 1755
rect 1547 1752 1552 1754
rect 1547 1751 1548 1752
rect 1542 1750 1548 1751
rect 1551 1751 1552 1752
rect 1556 1751 1557 1755
rect 1551 1750 1557 1751
rect 1631 1755 1637 1756
rect 1631 1751 1632 1755
rect 1636 1754 1637 1755
rect 1702 1755 1708 1756
rect 1702 1754 1703 1755
rect 1636 1752 1703 1754
rect 1636 1751 1637 1752
rect 1631 1750 1637 1751
rect 1702 1751 1703 1752
rect 1707 1751 1708 1755
rect 1702 1750 1708 1751
rect 1711 1755 1720 1756
rect 1711 1751 1712 1755
rect 1719 1751 1720 1755
rect 1711 1750 1720 1751
rect 1782 1755 1788 1756
rect 1782 1751 1783 1755
rect 1787 1754 1788 1755
rect 1791 1755 1797 1756
rect 1791 1754 1792 1755
rect 1787 1752 1792 1754
rect 1787 1751 1788 1752
rect 1782 1750 1788 1751
rect 1791 1751 1792 1752
rect 1796 1751 1797 1755
rect 1791 1750 1797 1751
rect 1862 1755 1868 1756
rect 1862 1751 1863 1755
rect 1867 1754 1868 1755
rect 1871 1755 1877 1756
rect 1871 1754 1872 1755
rect 1867 1752 1872 1754
rect 1867 1751 1868 1752
rect 1862 1750 1868 1751
rect 1871 1751 1872 1752
rect 1876 1751 1877 1755
rect 1871 1750 1877 1751
rect 1942 1755 1948 1756
rect 1942 1751 1943 1755
rect 1947 1754 1948 1755
rect 1951 1755 1957 1756
rect 1951 1754 1952 1755
rect 1947 1752 1952 1754
rect 1947 1751 1948 1752
rect 1942 1750 1948 1751
rect 1951 1751 1952 1752
rect 1956 1751 1957 1755
rect 1951 1750 1957 1751
rect 2030 1755 2037 1756
rect 2030 1751 2031 1755
rect 2036 1751 2037 1755
rect 2030 1750 2037 1751
rect 2094 1755 2101 1756
rect 2118 1755 2124 1756
rect 2094 1751 2095 1755
rect 2100 1751 2101 1755
rect 2094 1750 2101 1751
rect 1094 1748 1100 1749
rect 1134 1743 1140 1744
rect 255 1739 261 1740
rect 110 1736 116 1737
rect 110 1732 111 1736
rect 115 1732 116 1736
rect 255 1735 256 1739
rect 260 1738 261 1739
rect 286 1739 292 1740
rect 286 1738 287 1739
rect 260 1736 287 1738
rect 260 1735 261 1736
rect 255 1734 261 1735
rect 286 1735 287 1736
rect 291 1735 292 1739
rect 286 1734 292 1735
rect 306 1739 312 1740
rect 306 1735 307 1739
rect 311 1738 312 1739
rect 319 1739 325 1740
rect 319 1738 320 1739
rect 311 1736 320 1738
rect 311 1735 312 1736
rect 306 1734 312 1735
rect 319 1735 320 1736
rect 324 1735 325 1739
rect 319 1734 325 1735
rect 374 1739 381 1740
rect 374 1735 375 1739
rect 380 1735 381 1739
rect 374 1734 381 1735
rect 383 1739 389 1740
rect 383 1735 384 1739
rect 388 1738 389 1739
rect 439 1739 445 1740
rect 439 1738 440 1739
rect 388 1736 440 1738
rect 388 1735 389 1736
rect 383 1734 389 1735
rect 439 1735 440 1736
rect 444 1735 445 1739
rect 439 1734 445 1735
rect 462 1739 468 1740
rect 462 1735 463 1739
rect 467 1738 468 1739
rect 503 1739 509 1740
rect 503 1738 504 1739
rect 467 1736 504 1738
rect 467 1735 468 1736
rect 462 1734 468 1735
rect 503 1735 504 1736
rect 508 1735 509 1739
rect 503 1734 509 1735
rect 511 1739 517 1740
rect 511 1735 512 1739
rect 516 1738 517 1739
rect 567 1739 573 1740
rect 567 1738 568 1739
rect 516 1736 568 1738
rect 516 1735 517 1736
rect 511 1734 517 1735
rect 567 1735 568 1736
rect 572 1735 573 1739
rect 567 1734 573 1735
rect 639 1739 645 1740
rect 639 1735 640 1739
rect 644 1738 645 1739
rect 662 1739 668 1740
rect 662 1738 663 1739
rect 644 1736 663 1738
rect 644 1735 645 1736
rect 639 1734 645 1735
rect 662 1735 663 1736
rect 667 1735 668 1739
rect 662 1734 668 1735
rect 674 1739 680 1740
rect 674 1735 675 1739
rect 679 1738 680 1739
rect 711 1739 717 1740
rect 711 1738 712 1739
rect 679 1736 712 1738
rect 679 1735 680 1736
rect 674 1734 680 1735
rect 711 1735 712 1736
rect 716 1735 717 1739
rect 711 1734 717 1735
rect 719 1739 725 1740
rect 719 1735 720 1739
rect 724 1738 725 1739
rect 783 1739 789 1740
rect 783 1738 784 1739
rect 724 1736 784 1738
rect 724 1735 725 1736
rect 719 1734 725 1735
rect 783 1735 784 1736
rect 788 1735 789 1739
rect 783 1734 789 1735
rect 855 1739 861 1740
rect 855 1735 856 1739
rect 860 1738 861 1739
rect 926 1739 932 1740
rect 926 1738 927 1739
rect 860 1736 927 1738
rect 860 1735 861 1736
rect 855 1734 861 1735
rect 926 1735 927 1736
rect 931 1735 932 1739
rect 926 1734 932 1735
rect 935 1739 941 1740
rect 935 1735 936 1739
rect 940 1738 941 1739
rect 1002 1739 1008 1740
rect 1002 1738 1003 1739
rect 940 1736 1003 1738
rect 940 1735 941 1736
rect 935 1734 941 1735
rect 1002 1735 1003 1736
rect 1007 1735 1008 1739
rect 1002 1734 1008 1735
rect 1010 1739 1021 1740
rect 1010 1735 1011 1739
rect 1015 1735 1016 1739
rect 1020 1735 1021 1739
rect 1134 1739 1135 1743
rect 1139 1739 1140 1743
rect 2118 1743 2124 1744
rect 1134 1738 1140 1739
rect 1190 1740 1196 1741
rect 1010 1734 1021 1735
rect 1094 1736 1100 1737
rect 110 1731 116 1732
rect 1094 1732 1095 1736
rect 1099 1732 1100 1736
rect 1190 1736 1191 1740
rect 1195 1736 1196 1740
rect 1190 1735 1196 1736
rect 1254 1740 1260 1741
rect 1254 1736 1255 1740
rect 1259 1736 1260 1740
rect 1254 1735 1260 1736
rect 1318 1740 1324 1741
rect 1318 1736 1319 1740
rect 1323 1736 1324 1740
rect 1318 1735 1324 1736
rect 1382 1740 1388 1741
rect 1382 1736 1383 1740
rect 1387 1736 1388 1740
rect 1382 1735 1388 1736
rect 1454 1740 1460 1741
rect 1454 1736 1455 1740
rect 1459 1736 1460 1740
rect 1454 1735 1460 1736
rect 1526 1740 1532 1741
rect 1526 1736 1527 1740
rect 1531 1736 1532 1740
rect 1526 1735 1532 1736
rect 1606 1740 1612 1741
rect 1606 1736 1607 1740
rect 1611 1736 1612 1740
rect 1606 1735 1612 1736
rect 1686 1740 1692 1741
rect 1686 1736 1687 1740
rect 1691 1736 1692 1740
rect 1686 1735 1692 1736
rect 1766 1740 1772 1741
rect 1766 1736 1767 1740
rect 1771 1736 1772 1740
rect 1766 1735 1772 1736
rect 1846 1740 1852 1741
rect 1846 1736 1847 1740
rect 1851 1736 1852 1740
rect 1846 1735 1852 1736
rect 1926 1740 1932 1741
rect 1926 1736 1927 1740
rect 1931 1736 1932 1740
rect 1926 1735 1932 1736
rect 2006 1740 2012 1741
rect 2006 1736 2007 1740
rect 2011 1736 2012 1740
rect 2006 1735 2012 1736
rect 2070 1740 2076 1741
rect 2070 1736 2071 1740
rect 2075 1736 2076 1740
rect 2118 1739 2119 1743
rect 2123 1739 2124 1743
rect 2118 1738 2124 1739
rect 2070 1735 2076 1736
rect 1094 1731 1100 1732
rect 230 1728 236 1729
rect 230 1724 231 1728
rect 235 1724 236 1728
rect 230 1723 236 1724
rect 294 1728 300 1729
rect 294 1724 295 1728
rect 299 1724 300 1728
rect 294 1723 300 1724
rect 350 1728 356 1729
rect 350 1724 351 1728
rect 355 1724 356 1728
rect 350 1723 356 1724
rect 414 1728 420 1729
rect 414 1724 415 1728
rect 419 1724 420 1728
rect 414 1723 420 1724
rect 478 1728 484 1729
rect 478 1724 479 1728
rect 483 1724 484 1728
rect 478 1723 484 1724
rect 542 1728 548 1729
rect 542 1724 543 1728
rect 547 1724 548 1728
rect 542 1723 548 1724
rect 614 1728 620 1729
rect 614 1724 615 1728
rect 619 1724 620 1728
rect 614 1723 620 1724
rect 686 1728 692 1729
rect 686 1724 687 1728
rect 691 1724 692 1728
rect 686 1723 692 1724
rect 758 1728 764 1729
rect 758 1724 759 1728
rect 763 1724 764 1728
rect 758 1723 764 1724
rect 830 1728 836 1729
rect 830 1724 831 1728
rect 835 1724 836 1728
rect 830 1723 836 1724
rect 910 1728 916 1729
rect 910 1724 911 1728
rect 915 1724 916 1728
rect 910 1723 916 1724
rect 990 1728 996 1729
rect 990 1724 991 1728
rect 995 1724 996 1728
rect 1246 1728 1252 1729
rect 990 1723 996 1724
rect 1134 1725 1140 1726
rect 1134 1721 1135 1725
rect 1139 1721 1140 1725
rect 1246 1724 1247 1728
rect 1251 1724 1252 1728
rect 1246 1723 1252 1724
rect 1294 1728 1300 1729
rect 1294 1724 1295 1728
rect 1299 1724 1300 1728
rect 1294 1723 1300 1724
rect 1342 1728 1348 1729
rect 1342 1724 1343 1728
rect 1347 1724 1348 1728
rect 1342 1723 1348 1724
rect 1398 1728 1404 1729
rect 1398 1724 1399 1728
rect 1403 1724 1404 1728
rect 1398 1723 1404 1724
rect 1462 1728 1468 1729
rect 1462 1724 1463 1728
rect 1467 1724 1468 1728
rect 1462 1723 1468 1724
rect 1526 1728 1532 1729
rect 1526 1724 1527 1728
rect 1531 1724 1532 1728
rect 1526 1723 1532 1724
rect 1598 1728 1604 1729
rect 1598 1724 1599 1728
rect 1603 1724 1604 1728
rect 1598 1723 1604 1724
rect 1670 1728 1676 1729
rect 1670 1724 1671 1728
rect 1675 1724 1676 1728
rect 1670 1723 1676 1724
rect 1742 1728 1748 1729
rect 1742 1724 1743 1728
rect 1747 1724 1748 1728
rect 1742 1723 1748 1724
rect 1806 1728 1812 1729
rect 1806 1724 1807 1728
rect 1811 1724 1812 1728
rect 1806 1723 1812 1724
rect 1878 1728 1884 1729
rect 1878 1724 1879 1728
rect 1883 1724 1884 1728
rect 1878 1723 1884 1724
rect 1950 1728 1956 1729
rect 1950 1724 1951 1728
rect 1955 1724 1956 1728
rect 1950 1723 1956 1724
rect 2022 1728 2028 1729
rect 2022 1724 2023 1728
rect 2027 1724 2028 1728
rect 2022 1723 2028 1724
rect 2070 1728 2076 1729
rect 2070 1724 2071 1728
rect 2075 1724 2076 1728
rect 2070 1723 2076 1724
rect 2118 1725 2124 1726
rect 1134 1720 1140 1721
rect 2118 1721 2119 1725
rect 2123 1721 2124 1725
rect 2118 1720 2124 1721
rect 255 1719 264 1720
rect 255 1715 256 1719
rect 263 1715 264 1719
rect 255 1714 264 1715
rect 286 1719 292 1720
rect 286 1715 287 1719
rect 291 1718 292 1719
rect 319 1719 325 1720
rect 319 1718 320 1719
rect 291 1716 320 1718
rect 291 1715 292 1716
rect 286 1714 292 1715
rect 319 1715 320 1716
rect 324 1715 325 1719
rect 319 1714 325 1715
rect 375 1719 381 1720
rect 375 1715 376 1719
rect 380 1718 381 1719
rect 383 1719 389 1720
rect 383 1718 384 1719
rect 380 1716 384 1718
rect 380 1715 381 1716
rect 375 1714 381 1715
rect 383 1715 384 1716
rect 388 1715 389 1719
rect 383 1714 389 1715
rect 439 1719 445 1720
rect 439 1715 440 1719
rect 444 1718 445 1719
rect 462 1719 468 1720
rect 462 1718 463 1719
rect 444 1716 463 1718
rect 444 1715 445 1716
rect 439 1714 445 1715
rect 462 1715 463 1716
rect 467 1715 468 1719
rect 462 1714 468 1715
rect 503 1719 509 1720
rect 503 1715 504 1719
rect 508 1718 509 1719
rect 511 1719 517 1720
rect 511 1718 512 1719
rect 508 1716 512 1718
rect 508 1715 509 1716
rect 503 1714 509 1715
rect 511 1715 512 1716
rect 516 1715 517 1719
rect 511 1714 517 1715
rect 567 1719 576 1720
rect 567 1715 568 1719
rect 575 1715 576 1719
rect 567 1714 576 1715
rect 639 1719 645 1720
rect 639 1715 640 1719
rect 644 1718 645 1719
rect 674 1719 680 1720
rect 674 1718 675 1719
rect 644 1716 675 1718
rect 644 1715 645 1716
rect 639 1714 645 1715
rect 674 1715 675 1716
rect 679 1715 680 1719
rect 674 1714 680 1715
rect 711 1719 717 1720
rect 711 1715 712 1719
rect 716 1718 717 1719
rect 719 1719 725 1720
rect 719 1718 720 1719
rect 716 1716 720 1718
rect 716 1715 717 1716
rect 711 1714 717 1715
rect 719 1715 720 1716
rect 724 1715 725 1719
rect 719 1714 725 1715
rect 782 1719 789 1720
rect 782 1715 783 1719
rect 788 1715 789 1719
rect 782 1714 789 1715
rect 798 1719 804 1720
rect 798 1715 799 1719
rect 803 1718 804 1719
rect 855 1719 861 1720
rect 855 1718 856 1719
rect 803 1716 856 1718
rect 803 1715 804 1716
rect 798 1714 804 1715
rect 855 1715 856 1716
rect 860 1715 861 1719
rect 855 1714 861 1715
rect 926 1719 932 1720
rect 926 1715 927 1719
rect 931 1718 932 1719
rect 935 1719 941 1720
rect 935 1718 936 1719
rect 931 1716 936 1718
rect 931 1715 932 1716
rect 926 1714 932 1715
rect 935 1715 936 1716
rect 940 1715 941 1719
rect 935 1714 941 1715
rect 1002 1719 1008 1720
rect 1002 1715 1003 1719
rect 1007 1718 1008 1719
rect 1015 1719 1021 1720
rect 1015 1718 1016 1719
rect 1007 1716 1016 1718
rect 1007 1715 1008 1716
rect 1002 1714 1008 1715
rect 1015 1715 1016 1716
rect 1020 1715 1021 1719
rect 1015 1714 1021 1715
rect 1271 1711 1277 1712
rect 1134 1708 1140 1709
rect 1134 1704 1135 1708
rect 1139 1704 1140 1708
rect 1271 1707 1272 1711
rect 1276 1710 1277 1711
rect 1310 1711 1316 1712
rect 1310 1710 1311 1711
rect 1276 1708 1311 1710
rect 1276 1707 1277 1708
rect 1271 1706 1277 1707
rect 1310 1707 1311 1708
rect 1315 1707 1316 1711
rect 1310 1706 1316 1707
rect 1319 1711 1325 1712
rect 1319 1707 1320 1711
rect 1324 1710 1325 1711
rect 1358 1711 1364 1712
rect 1358 1710 1359 1711
rect 1324 1708 1359 1710
rect 1324 1707 1325 1708
rect 1319 1706 1325 1707
rect 1358 1707 1359 1708
rect 1363 1707 1364 1711
rect 1358 1706 1364 1707
rect 1366 1711 1373 1712
rect 1366 1707 1367 1711
rect 1372 1707 1373 1711
rect 1366 1706 1373 1707
rect 1423 1711 1429 1712
rect 1423 1707 1424 1711
rect 1428 1710 1429 1711
rect 1478 1711 1484 1712
rect 1478 1710 1479 1711
rect 1428 1708 1479 1710
rect 1428 1707 1429 1708
rect 1423 1706 1429 1707
rect 1478 1707 1479 1708
rect 1483 1707 1484 1711
rect 1478 1706 1484 1707
rect 1487 1711 1493 1712
rect 1487 1707 1488 1711
rect 1492 1710 1493 1711
rect 1534 1711 1540 1712
rect 1534 1710 1535 1711
rect 1492 1708 1535 1710
rect 1492 1707 1493 1708
rect 1487 1706 1493 1707
rect 1534 1707 1535 1708
rect 1539 1707 1540 1711
rect 1534 1706 1540 1707
rect 1542 1711 1548 1712
rect 1542 1707 1543 1711
rect 1547 1710 1548 1711
rect 1551 1711 1557 1712
rect 1551 1710 1552 1711
rect 1547 1708 1552 1710
rect 1547 1707 1548 1708
rect 1542 1706 1548 1707
rect 1551 1707 1552 1708
rect 1556 1707 1557 1711
rect 1551 1706 1557 1707
rect 1623 1711 1629 1712
rect 1623 1707 1624 1711
rect 1628 1710 1629 1711
rect 1686 1711 1692 1712
rect 1686 1710 1687 1711
rect 1628 1708 1687 1710
rect 1628 1707 1629 1708
rect 1623 1706 1629 1707
rect 1686 1707 1687 1708
rect 1691 1707 1692 1711
rect 1686 1706 1692 1707
rect 1694 1711 1701 1712
rect 1694 1707 1695 1711
rect 1700 1707 1701 1711
rect 1694 1706 1701 1707
rect 1767 1711 1773 1712
rect 1767 1707 1768 1711
rect 1772 1710 1773 1711
rect 1814 1711 1820 1712
rect 1814 1710 1815 1711
rect 1772 1708 1815 1710
rect 1772 1707 1773 1708
rect 1767 1706 1773 1707
rect 1814 1707 1815 1708
rect 1819 1707 1820 1711
rect 1814 1706 1820 1707
rect 1831 1711 1837 1712
rect 1831 1707 1832 1711
rect 1836 1710 1837 1711
rect 1894 1711 1900 1712
rect 1894 1710 1895 1711
rect 1836 1708 1895 1710
rect 1836 1707 1837 1708
rect 1831 1706 1837 1707
rect 1894 1707 1895 1708
rect 1899 1707 1900 1711
rect 1894 1706 1900 1707
rect 1903 1711 1909 1712
rect 1903 1707 1904 1711
rect 1908 1710 1909 1711
rect 1934 1711 1940 1712
rect 1934 1710 1935 1711
rect 1908 1708 1935 1710
rect 1908 1707 1909 1708
rect 1903 1706 1909 1707
rect 1934 1707 1935 1708
rect 1939 1707 1940 1711
rect 1934 1706 1940 1707
rect 1975 1711 1981 1712
rect 1975 1707 1976 1711
rect 1980 1710 1981 1711
rect 2014 1711 2020 1712
rect 2014 1710 2015 1711
rect 1980 1708 2015 1710
rect 1980 1707 1981 1708
rect 1975 1706 1981 1707
rect 2014 1707 2015 1708
rect 2019 1707 2020 1711
rect 2014 1706 2020 1707
rect 2046 1711 2053 1712
rect 2046 1707 2047 1711
rect 2052 1707 2053 1711
rect 2046 1706 2053 1707
rect 2055 1711 2061 1712
rect 2055 1707 2056 1711
rect 2060 1710 2061 1711
rect 2095 1711 2101 1712
rect 2095 1710 2096 1711
rect 2060 1708 2096 1710
rect 2060 1707 2061 1708
rect 2055 1706 2061 1707
rect 2095 1707 2096 1708
rect 2100 1707 2101 1711
rect 2095 1706 2101 1707
rect 2118 1708 2124 1709
rect 1134 1703 1140 1704
rect 2118 1704 2119 1708
rect 2123 1704 2124 1708
rect 2118 1703 2124 1704
rect 1246 1700 1252 1701
rect 1246 1696 1247 1700
rect 1251 1696 1252 1700
rect 159 1695 165 1696
rect 159 1691 160 1695
rect 164 1694 165 1695
rect 206 1695 212 1696
rect 206 1694 207 1695
rect 164 1692 207 1694
rect 164 1691 165 1692
rect 159 1690 165 1691
rect 206 1691 207 1692
rect 211 1691 212 1695
rect 206 1690 212 1691
rect 223 1695 229 1696
rect 223 1691 224 1695
rect 228 1694 229 1695
rect 294 1695 300 1696
rect 294 1694 295 1695
rect 228 1692 295 1694
rect 228 1691 229 1692
rect 223 1690 229 1691
rect 294 1691 295 1692
rect 299 1691 300 1695
rect 294 1690 300 1691
rect 303 1695 312 1696
rect 303 1691 304 1695
rect 311 1691 312 1695
rect 303 1690 312 1691
rect 314 1695 320 1696
rect 314 1691 315 1695
rect 319 1694 320 1695
rect 391 1695 397 1696
rect 391 1694 392 1695
rect 319 1692 392 1694
rect 319 1691 320 1692
rect 314 1690 320 1691
rect 391 1691 392 1692
rect 396 1691 397 1695
rect 391 1690 397 1691
rect 399 1695 405 1696
rect 399 1691 400 1695
rect 404 1694 405 1695
rect 487 1695 493 1696
rect 487 1694 488 1695
rect 404 1692 488 1694
rect 404 1691 405 1692
rect 399 1690 405 1691
rect 487 1691 488 1692
rect 492 1691 493 1695
rect 487 1690 493 1691
rect 495 1695 501 1696
rect 495 1691 496 1695
rect 500 1694 501 1695
rect 575 1695 581 1696
rect 575 1694 576 1695
rect 500 1692 576 1694
rect 500 1691 501 1692
rect 495 1690 501 1691
rect 575 1691 576 1692
rect 580 1691 581 1695
rect 575 1690 581 1691
rect 662 1695 669 1696
rect 662 1691 663 1695
rect 668 1691 669 1695
rect 662 1690 669 1691
rect 743 1695 749 1696
rect 743 1691 744 1695
rect 748 1694 749 1695
rect 806 1695 812 1696
rect 806 1694 807 1695
rect 748 1692 807 1694
rect 748 1691 749 1692
rect 743 1690 749 1691
rect 806 1691 807 1692
rect 811 1691 812 1695
rect 806 1690 812 1691
rect 815 1695 821 1696
rect 815 1691 816 1695
rect 820 1694 821 1695
rect 862 1695 868 1696
rect 862 1694 863 1695
rect 820 1692 863 1694
rect 820 1691 821 1692
rect 815 1690 821 1691
rect 862 1691 863 1692
rect 867 1691 868 1695
rect 862 1690 868 1691
rect 870 1695 876 1696
rect 870 1691 871 1695
rect 875 1694 876 1695
rect 879 1695 885 1696
rect 879 1694 880 1695
rect 875 1692 880 1694
rect 875 1691 876 1692
rect 870 1690 876 1691
rect 879 1691 880 1692
rect 884 1691 885 1695
rect 879 1690 885 1691
rect 943 1695 949 1696
rect 943 1691 944 1695
rect 948 1694 949 1695
rect 998 1695 1004 1696
rect 998 1694 999 1695
rect 948 1692 999 1694
rect 948 1691 949 1692
rect 943 1690 949 1691
rect 998 1691 999 1692
rect 1003 1691 1004 1695
rect 998 1690 1004 1691
rect 1007 1695 1016 1696
rect 1007 1691 1008 1695
rect 1015 1691 1016 1695
rect 1071 1695 1077 1696
rect 1246 1695 1252 1696
rect 1294 1700 1300 1701
rect 1294 1696 1295 1700
rect 1299 1696 1300 1700
rect 1294 1695 1300 1696
rect 1342 1700 1348 1701
rect 1342 1696 1343 1700
rect 1347 1696 1348 1700
rect 1342 1695 1348 1696
rect 1398 1700 1404 1701
rect 1398 1696 1399 1700
rect 1403 1696 1404 1700
rect 1398 1695 1404 1696
rect 1462 1700 1468 1701
rect 1462 1696 1463 1700
rect 1467 1696 1468 1700
rect 1462 1695 1468 1696
rect 1526 1700 1532 1701
rect 1526 1696 1527 1700
rect 1531 1696 1532 1700
rect 1526 1695 1532 1696
rect 1598 1700 1604 1701
rect 1598 1696 1599 1700
rect 1603 1696 1604 1700
rect 1598 1695 1604 1696
rect 1670 1700 1676 1701
rect 1670 1696 1671 1700
rect 1675 1696 1676 1700
rect 1670 1695 1676 1696
rect 1742 1700 1748 1701
rect 1742 1696 1743 1700
rect 1747 1696 1748 1700
rect 1806 1700 1812 1701
rect 1806 1696 1807 1700
rect 1811 1696 1812 1700
rect 1742 1695 1748 1696
rect 1782 1695 1788 1696
rect 1806 1695 1812 1696
rect 1878 1700 1884 1701
rect 1878 1696 1879 1700
rect 1883 1696 1884 1700
rect 1878 1695 1884 1696
rect 1950 1700 1956 1701
rect 1950 1696 1951 1700
rect 1955 1696 1956 1700
rect 1950 1695 1956 1696
rect 2022 1700 2028 1701
rect 2022 1696 2023 1700
rect 2027 1696 2028 1700
rect 2022 1695 2028 1696
rect 2070 1700 2076 1701
rect 2070 1696 2071 1700
rect 2075 1696 2076 1700
rect 2070 1695 2076 1696
rect 1071 1694 1072 1695
rect 1007 1690 1016 1691
rect 1020 1692 1072 1694
rect 134 1688 140 1689
rect 134 1684 135 1688
rect 139 1684 140 1688
rect 134 1683 140 1684
rect 198 1688 204 1689
rect 198 1684 199 1688
rect 203 1684 204 1688
rect 198 1683 204 1684
rect 278 1688 284 1689
rect 278 1684 279 1688
rect 283 1684 284 1688
rect 278 1683 284 1684
rect 366 1688 372 1689
rect 366 1684 367 1688
rect 371 1684 372 1688
rect 366 1683 372 1684
rect 462 1688 468 1689
rect 462 1684 463 1688
rect 467 1684 468 1688
rect 462 1683 468 1684
rect 550 1688 556 1689
rect 550 1684 551 1688
rect 555 1684 556 1688
rect 550 1683 556 1684
rect 638 1688 644 1689
rect 638 1684 639 1688
rect 643 1684 644 1688
rect 638 1683 644 1684
rect 718 1688 724 1689
rect 718 1684 719 1688
rect 723 1684 724 1688
rect 718 1683 724 1684
rect 790 1688 796 1689
rect 790 1684 791 1688
rect 795 1684 796 1688
rect 790 1683 796 1684
rect 854 1688 860 1689
rect 854 1684 855 1688
rect 859 1684 860 1688
rect 854 1683 860 1684
rect 918 1688 924 1689
rect 918 1684 919 1688
rect 923 1684 924 1688
rect 918 1683 924 1684
rect 982 1688 988 1689
rect 982 1684 983 1688
rect 987 1684 988 1688
rect 982 1683 988 1684
rect 1020 1682 1022 1692
rect 1071 1691 1072 1692
rect 1076 1691 1077 1695
rect 1782 1694 1783 1695
rect 1767 1693 1783 1694
rect 1071 1690 1077 1691
rect 1271 1691 1277 1692
rect 1046 1688 1052 1689
rect 1046 1684 1047 1688
rect 1051 1684 1052 1688
rect 1271 1687 1272 1691
rect 1276 1690 1277 1691
rect 1286 1691 1292 1692
rect 1286 1690 1287 1691
rect 1276 1688 1287 1690
rect 1276 1687 1277 1688
rect 1271 1686 1277 1687
rect 1286 1687 1287 1688
rect 1291 1687 1292 1691
rect 1286 1686 1292 1687
rect 1310 1691 1316 1692
rect 1310 1687 1311 1691
rect 1315 1690 1316 1691
rect 1319 1691 1325 1692
rect 1319 1690 1320 1691
rect 1315 1688 1320 1690
rect 1315 1687 1316 1688
rect 1310 1686 1316 1687
rect 1319 1687 1320 1688
rect 1324 1687 1325 1691
rect 1319 1686 1325 1687
rect 1358 1691 1364 1692
rect 1358 1687 1359 1691
rect 1363 1690 1364 1691
rect 1367 1691 1373 1692
rect 1367 1690 1368 1691
rect 1363 1688 1368 1690
rect 1363 1687 1364 1688
rect 1358 1686 1364 1687
rect 1367 1687 1368 1688
rect 1372 1687 1373 1691
rect 1367 1686 1373 1687
rect 1410 1691 1416 1692
rect 1410 1687 1411 1691
rect 1415 1690 1416 1691
rect 1423 1691 1429 1692
rect 1423 1690 1424 1691
rect 1415 1688 1424 1690
rect 1415 1687 1416 1688
rect 1410 1686 1416 1687
rect 1423 1687 1424 1688
rect 1428 1687 1429 1691
rect 1423 1686 1429 1687
rect 1478 1691 1484 1692
rect 1478 1687 1479 1691
rect 1483 1690 1484 1691
rect 1487 1691 1493 1692
rect 1487 1690 1488 1691
rect 1483 1688 1488 1690
rect 1483 1687 1484 1688
rect 1478 1686 1484 1687
rect 1487 1687 1488 1688
rect 1492 1687 1493 1691
rect 1487 1686 1493 1687
rect 1534 1691 1540 1692
rect 1534 1687 1535 1691
rect 1539 1690 1540 1691
rect 1551 1691 1557 1692
rect 1551 1690 1552 1691
rect 1539 1688 1552 1690
rect 1539 1687 1540 1688
rect 1534 1686 1540 1687
rect 1551 1687 1552 1688
rect 1556 1687 1557 1691
rect 1551 1686 1557 1687
rect 1610 1691 1616 1692
rect 1610 1687 1611 1691
rect 1615 1690 1616 1691
rect 1623 1691 1629 1692
rect 1623 1690 1624 1691
rect 1615 1688 1624 1690
rect 1615 1687 1616 1688
rect 1610 1686 1616 1687
rect 1623 1687 1624 1688
rect 1628 1687 1629 1691
rect 1623 1686 1629 1687
rect 1686 1691 1692 1692
rect 1686 1687 1687 1691
rect 1691 1690 1692 1691
rect 1695 1691 1701 1692
rect 1695 1690 1696 1691
rect 1691 1688 1696 1690
rect 1691 1687 1692 1688
rect 1686 1686 1692 1687
rect 1695 1687 1696 1688
rect 1700 1687 1701 1691
rect 1767 1689 1768 1693
rect 1772 1692 1783 1693
rect 1772 1689 1773 1692
rect 1782 1691 1783 1692
rect 1787 1691 1788 1695
rect 1782 1690 1788 1691
rect 1814 1691 1820 1692
rect 1767 1688 1773 1689
rect 1695 1686 1701 1687
rect 1814 1687 1815 1691
rect 1819 1690 1820 1691
rect 1831 1691 1837 1692
rect 1831 1690 1832 1691
rect 1819 1688 1832 1690
rect 1819 1687 1820 1688
rect 1814 1686 1820 1687
rect 1831 1687 1832 1688
rect 1836 1687 1837 1691
rect 1831 1686 1837 1687
rect 1894 1691 1900 1692
rect 1894 1687 1895 1691
rect 1899 1690 1900 1691
rect 1903 1691 1909 1692
rect 1903 1690 1904 1691
rect 1899 1688 1904 1690
rect 1899 1687 1900 1688
rect 1894 1686 1900 1687
rect 1903 1687 1904 1688
rect 1908 1687 1909 1691
rect 1903 1686 1909 1687
rect 1975 1691 1981 1692
rect 1975 1687 1976 1691
rect 1980 1690 1981 1691
rect 1986 1691 1992 1692
rect 1986 1690 1987 1691
rect 1980 1688 1987 1690
rect 1980 1687 1981 1688
rect 1975 1686 1981 1687
rect 1986 1687 1987 1688
rect 1991 1687 1992 1691
rect 1986 1686 1992 1687
rect 2047 1691 2053 1692
rect 2047 1687 2048 1691
rect 2052 1690 2053 1691
rect 2055 1691 2061 1692
rect 2055 1690 2056 1691
rect 2052 1688 2056 1690
rect 2052 1687 2053 1688
rect 2047 1686 2053 1687
rect 2055 1687 2056 1688
rect 2060 1687 2061 1691
rect 2055 1686 2061 1687
rect 2094 1691 2101 1692
rect 2094 1687 2095 1691
rect 2100 1687 2101 1691
rect 2094 1686 2101 1687
rect 1046 1683 1052 1684
rect 110 1680 116 1681
rect 110 1676 111 1680
rect 115 1676 116 1680
rect 992 1680 1022 1682
rect 1094 1680 1100 1681
rect 110 1675 116 1676
rect 159 1675 165 1676
rect 159 1671 160 1675
rect 164 1674 165 1675
rect 190 1675 196 1676
rect 190 1674 191 1675
rect 164 1672 191 1674
rect 164 1671 165 1672
rect 159 1670 165 1671
rect 190 1671 191 1672
rect 195 1671 196 1675
rect 190 1670 196 1671
rect 206 1675 212 1676
rect 206 1671 207 1675
rect 211 1674 212 1675
rect 223 1675 229 1676
rect 223 1674 224 1675
rect 211 1672 224 1674
rect 211 1671 212 1672
rect 206 1670 212 1671
rect 223 1671 224 1672
rect 228 1671 229 1675
rect 223 1670 229 1671
rect 294 1675 300 1676
rect 294 1671 295 1675
rect 299 1674 300 1675
rect 303 1675 309 1676
rect 303 1674 304 1675
rect 299 1672 304 1674
rect 299 1671 300 1672
rect 294 1670 300 1671
rect 303 1671 304 1672
rect 308 1671 309 1675
rect 303 1670 309 1671
rect 391 1675 397 1676
rect 391 1671 392 1675
rect 396 1674 397 1675
rect 399 1675 405 1676
rect 399 1674 400 1675
rect 396 1672 400 1674
rect 396 1671 397 1672
rect 391 1670 397 1671
rect 399 1671 400 1672
rect 404 1671 405 1675
rect 399 1670 405 1671
rect 487 1675 493 1676
rect 487 1671 488 1675
rect 492 1674 493 1675
rect 495 1675 501 1676
rect 495 1674 496 1675
rect 492 1672 496 1674
rect 492 1671 493 1672
rect 487 1670 493 1671
rect 495 1671 496 1672
rect 500 1671 501 1675
rect 495 1670 501 1671
rect 570 1675 581 1676
rect 570 1671 571 1675
rect 575 1671 576 1675
rect 580 1671 581 1675
rect 570 1670 581 1671
rect 610 1675 616 1676
rect 610 1671 611 1675
rect 615 1674 616 1675
rect 663 1675 669 1676
rect 663 1674 664 1675
rect 615 1672 664 1674
rect 615 1671 616 1672
rect 610 1670 616 1671
rect 663 1671 664 1672
rect 668 1671 669 1675
rect 663 1670 669 1671
rect 743 1675 749 1676
rect 743 1671 744 1675
rect 748 1674 749 1675
rect 798 1675 804 1676
rect 798 1674 799 1675
rect 748 1672 799 1674
rect 748 1671 749 1672
rect 743 1670 749 1671
rect 798 1671 799 1672
rect 803 1671 804 1675
rect 798 1670 804 1671
rect 806 1675 812 1676
rect 806 1671 807 1675
rect 811 1674 812 1675
rect 815 1675 821 1676
rect 815 1674 816 1675
rect 811 1672 816 1674
rect 811 1671 812 1672
rect 806 1670 812 1671
rect 815 1671 816 1672
rect 820 1671 821 1675
rect 815 1670 821 1671
rect 862 1675 868 1676
rect 862 1671 863 1675
rect 867 1674 868 1675
rect 879 1675 885 1676
rect 879 1674 880 1675
rect 867 1672 880 1674
rect 867 1671 868 1672
rect 862 1670 868 1671
rect 879 1671 880 1672
rect 884 1671 885 1675
rect 879 1670 885 1671
rect 943 1675 949 1676
rect 943 1671 944 1675
rect 948 1674 949 1675
rect 992 1674 994 1680
rect 1094 1676 1095 1680
rect 1099 1676 1100 1680
rect 948 1672 994 1674
rect 998 1675 1004 1676
rect 948 1671 949 1672
rect 943 1670 949 1671
rect 998 1671 999 1675
rect 1003 1674 1004 1675
rect 1007 1675 1013 1676
rect 1007 1674 1008 1675
rect 1003 1672 1008 1674
rect 1003 1671 1004 1672
rect 998 1670 1004 1671
rect 1007 1671 1008 1672
rect 1012 1671 1013 1675
rect 1007 1670 1013 1671
rect 1034 1675 1040 1676
rect 1034 1671 1035 1675
rect 1039 1674 1040 1675
rect 1071 1675 1077 1676
rect 1094 1675 1100 1676
rect 1071 1674 1072 1675
rect 1039 1672 1072 1674
rect 1039 1671 1040 1672
rect 1034 1670 1040 1671
rect 1071 1671 1072 1672
rect 1076 1671 1077 1675
rect 1071 1670 1077 1671
rect 1542 1671 1548 1672
rect 1542 1670 1543 1671
rect 1527 1669 1543 1670
rect 1287 1667 1293 1668
rect 110 1663 116 1664
rect 110 1659 111 1663
rect 115 1659 116 1663
rect 1094 1663 1100 1664
rect 110 1658 116 1659
rect 134 1660 140 1661
rect 134 1656 135 1660
rect 139 1656 140 1660
rect 134 1655 140 1656
rect 198 1660 204 1661
rect 198 1656 199 1660
rect 203 1656 204 1660
rect 198 1655 204 1656
rect 278 1660 284 1661
rect 278 1656 279 1660
rect 283 1656 284 1660
rect 278 1655 284 1656
rect 366 1660 372 1661
rect 366 1656 367 1660
rect 371 1656 372 1660
rect 366 1655 372 1656
rect 462 1660 468 1661
rect 462 1656 463 1660
rect 467 1656 468 1660
rect 462 1655 468 1656
rect 550 1660 556 1661
rect 550 1656 551 1660
rect 555 1656 556 1660
rect 550 1655 556 1656
rect 638 1660 644 1661
rect 638 1656 639 1660
rect 643 1656 644 1660
rect 638 1655 644 1656
rect 718 1660 724 1661
rect 718 1656 719 1660
rect 723 1656 724 1660
rect 718 1655 724 1656
rect 790 1660 796 1661
rect 790 1656 791 1660
rect 795 1656 796 1660
rect 790 1655 796 1656
rect 854 1660 860 1661
rect 854 1656 855 1660
rect 859 1656 860 1660
rect 854 1655 860 1656
rect 918 1660 924 1661
rect 918 1656 919 1660
rect 923 1656 924 1660
rect 918 1655 924 1656
rect 982 1660 988 1661
rect 982 1656 983 1660
rect 987 1656 988 1660
rect 982 1655 988 1656
rect 1046 1660 1052 1661
rect 1046 1656 1047 1660
rect 1051 1656 1052 1660
rect 1094 1659 1095 1663
rect 1099 1659 1100 1663
rect 1287 1663 1288 1667
rect 1292 1666 1293 1667
rect 1318 1667 1324 1668
rect 1318 1666 1319 1667
rect 1292 1664 1319 1666
rect 1292 1663 1293 1664
rect 1287 1662 1293 1663
rect 1318 1663 1319 1664
rect 1323 1663 1324 1667
rect 1318 1662 1324 1663
rect 1327 1667 1333 1668
rect 1327 1663 1328 1667
rect 1332 1666 1333 1667
rect 1358 1667 1364 1668
rect 1358 1666 1359 1667
rect 1332 1664 1359 1666
rect 1332 1663 1333 1664
rect 1327 1662 1333 1663
rect 1358 1663 1359 1664
rect 1363 1663 1364 1667
rect 1358 1662 1364 1663
rect 1367 1667 1373 1668
rect 1367 1663 1368 1667
rect 1372 1666 1373 1667
rect 1406 1667 1412 1668
rect 1406 1666 1407 1667
rect 1372 1664 1407 1666
rect 1372 1663 1373 1664
rect 1367 1662 1373 1663
rect 1406 1663 1407 1664
rect 1411 1663 1412 1667
rect 1406 1662 1412 1663
rect 1415 1667 1421 1668
rect 1415 1663 1416 1667
rect 1420 1666 1421 1667
rect 1462 1667 1468 1668
rect 1462 1666 1463 1667
rect 1420 1664 1463 1666
rect 1420 1663 1421 1664
rect 1415 1662 1421 1663
rect 1462 1663 1463 1664
rect 1467 1663 1468 1667
rect 1462 1662 1468 1663
rect 1471 1667 1477 1668
rect 1471 1663 1472 1667
rect 1476 1666 1477 1667
rect 1518 1667 1524 1668
rect 1518 1666 1519 1667
rect 1476 1664 1519 1666
rect 1476 1663 1477 1664
rect 1471 1662 1477 1663
rect 1518 1663 1519 1664
rect 1523 1663 1524 1667
rect 1527 1665 1528 1669
rect 1532 1668 1543 1669
rect 1532 1665 1533 1668
rect 1542 1667 1543 1668
rect 1547 1667 1548 1671
rect 1542 1666 1548 1667
rect 1591 1667 1597 1668
rect 1527 1664 1533 1665
rect 1518 1662 1524 1663
rect 1591 1663 1592 1667
rect 1596 1666 1597 1667
rect 1642 1667 1648 1668
rect 1642 1666 1643 1667
rect 1596 1664 1643 1666
rect 1596 1663 1597 1664
rect 1591 1662 1597 1663
rect 1642 1663 1643 1664
rect 1647 1663 1648 1667
rect 1642 1662 1648 1663
rect 1650 1667 1661 1668
rect 1650 1663 1651 1667
rect 1655 1663 1656 1667
rect 1660 1663 1661 1667
rect 1650 1662 1661 1663
rect 1719 1667 1725 1668
rect 1719 1663 1720 1667
rect 1724 1666 1725 1667
rect 1774 1667 1780 1668
rect 1774 1666 1775 1667
rect 1724 1664 1775 1666
rect 1724 1663 1725 1664
rect 1719 1662 1725 1663
rect 1774 1663 1775 1664
rect 1779 1663 1780 1667
rect 1774 1662 1780 1663
rect 1783 1667 1789 1668
rect 1783 1663 1784 1667
rect 1788 1666 1789 1667
rect 1846 1667 1852 1668
rect 1846 1666 1847 1667
rect 1788 1664 1847 1666
rect 1788 1663 1789 1664
rect 1783 1662 1789 1663
rect 1846 1663 1847 1664
rect 1851 1663 1852 1667
rect 1846 1662 1852 1663
rect 1855 1667 1861 1668
rect 1855 1663 1856 1667
rect 1860 1666 1861 1667
rect 1926 1667 1932 1668
rect 1926 1666 1927 1667
rect 1860 1664 1927 1666
rect 1860 1663 1861 1664
rect 1855 1662 1861 1663
rect 1926 1663 1927 1664
rect 1931 1663 1932 1667
rect 1926 1662 1932 1663
rect 1934 1667 1941 1668
rect 1934 1663 1935 1667
rect 1940 1663 1941 1667
rect 1934 1662 1941 1663
rect 2010 1667 2016 1668
rect 2010 1663 2011 1667
rect 2015 1666 2016 1667
rect 2023 1667 2029 1668
rect 2023 1666 2024 1667
rect 2015 1664 2024 1666
rect 2015 1663 2016 1664
rect 2010 1662 2016 1663
rect 2023 1663 2024 1664
rect 2028 1663 2029 1667
rect 2023 1662 2029 1663
rect 2046 1667 2052 1668
rect 2046 1663 2047 1667
rect 2051 1666 2052 1667
rect 2095 1667 2101 1668
rect 2095 1666 2096 1667
rect 2051 1664 2096 1666
rect 2051 1663 2052 1664
rect 2046 1662 2052 1663
rect 2095 1663 2096 1664
rect 2100 1663 2101 1667
rect 2095 1662 2101 1663
rect 1094 1658 1100 1659
rect 1262 1660 1268 1661
rect 1046 1655 1052 1656
rect 1262 1656 1263 1660
rect 1267 1656 1268 1660
rect 1262 1655 1268 1656
rect 1302 1660 1308 1661
rect 1302 1656 1303 1660
rect 1307 1656 1308 1660
rect 1302 1655 1308 1656
rect 1342 1660 1348 1661
rect 1342 1656 1343 1660
rect 1347 1656 1348 1660
rect 1342 1655 1348 1656
rect 1390 1660 1396 1661
rect 1390 1656 1391 1660
rect 1395 1656 1396 1660
rect 1390 1655 1396 1656
rect 1446 1660 1452 1661
rect 1446 1656 1447 1660
rect 1451 1656 1452 1660
rect 1446 1655 1452 1656
rect 1502 1660 1508 1661
rect 1502 1656 1503 1660
rect 1507 1656 1508 1660
rect 1502 1655 1508 1656
rect 1566 1660 1572 1661
rect 1566 1656 1567 1660
rect 1571 1656 1572 1660
rect 1566 1655 1572 1656
rect 1630 1660 1636 1661
rect 1630 1656 1631 1660
rect 1635 1656 1636 1660
rect 1630 1655 1636 1656
rect 1694 1660 1700 1661
rect 1694 1656 1695 1660
rect 1699 1656 1700 1660
rect 1694 1655 1700 1656
rect 1758 1660 1764 1661
rect 1758 1656 1759 1660
rect 1763 1656 1764 1660
rect 1758 1655 1764 1656
rect 1830 1660 1836 1661
rect 1830 1656 1831 1660
rect 1835 1656 1836 1660
rect 1830 1655 1836 1656
rect 1910 1660 1916 1661
rect 1910 1656 1911 1660
rect 1915 1656 1916 1660
rect 1910 1655 1916 1656
rect 1998 1660 2004 1661
rect 1998 1656 1999 1660
rect 2003 1656 2004 1660
rect 1998 1655 2004 1656
rect 2070 1660 2076 1661
rect 2070 1656 2071 1660
rect 2075 1656 2076 1660
rect 2070 1655 2076 1656
rect 1134 1652 1140 1653
rect 1134 1648 1135 1652
rect 1139 1648 1140 1652
rect 2118 1652 2124 1653
rect 2118 1648 2119 1652
rect 2123 1648 2124 1652
rect 1134 1647 1140 1648
rect 1286 1647 1293 1648
rect 134 1644 140 1645
rect 110 1641 116 1642
rect 110 1637 111 1641
rect 115 1637 116 1641
rect 134 1640 135 1644
rect 139 1640 140 1644
rect 134 1639 140 1640
rect 182 1644 188 1645
rect 182 1640 183 1644
rect 187 1640 188 1644
rect 182 1639 188 1640
rect 262 1644 268 1645
rect 262 1640 263 1644
rect 267 1640 268 1644
rect 262 1639 268 1640
rect 342 1644 348 1645
rect 342 1640 343 1644
rect 347 1640 348 1644
rect 342 1639 348 1640
rect 422 1644 428 1645
rect 422 1640 423 1644
rect 427 1640 428 1644
rect 422 1639 428 1640
rect 502 1644 508 1645
rect 502 1640 503 1644
rect 507 1640 508 1644
rect 502 1639 508 1640
rect 582 1644 588 1645
rect 582 1640 583 1644
rect 587 1640 588 1644
rect 582 1639 588 1640
rect 654 1644 660 1645
rect 654 1640 655 1644
rect 659 1640 660 1644
rect 654 1639 660 1640
rect 726 1644 732 1645
rect 726 1640 727 1644
rect 731 1640 732 1644
rect 726 1639 732 1640
rect 790 1644 796 1645
rect 790 1640 791 1644
rect 795 1640 796 1644
rect 790 1639 796 1640
rect 846 1644 852 1645
rect 846 1640 847 1644
rect 851 1640 852 1644
rect 846 1639 852 1640
rect 902 1644 908 1645
rect 902 1640 903 1644
rect 907 1640 908 1644
rect 902 1639 908 1640
rect 958 1644 964 1645
rect 958 1640 959 1644
rect 963 1640 964 1644
rect 958 1639 964 1640
rect 1006 1644 1012 1645
rect 1006 1640 1007 1644
rect 1011 1640 1012 1644
rect 1006 1639 1012 1640
rect 1046 1644 1052 1645
rect 1046 1640 1047 1644
rect 1051 1640 1052 1644
rect 1286 1643 1287 1647
rect 1292 1643 1293 1647
rect 1286 1642 1293 1643
rect 1318 1647 1324 1648
rect 1318 1643 1319 1647
rect 1323 1646 1324 1647
rect 1327 1647 1333 1648
rect 1327 1646 1328 1647
rect 1323 1644 1328 1646
rect 1323 1643 1324 1644
rect 1318 1642 1324 1643
rect 1327 1643 1328 1644
rect 1332 1643 1333 1647
rect 1327 1642 1333 1643
rect 1358 1647 1364 1648
rect 1358 1643 1359 1647
rect 1363 1646 1364 1647
rect 1367 1647 1373 1648
rect 1367 1646 1368 1647
rect 1363 1644 1368 1646
rect 1363 1643 1364 1644
rect 1358 1642 1364 1643
rect 1367 1643 1368 1644
rect 1372 1643 1373 1647
rect 1367 1642 1373 1643
rect 1406 1647 1412 1648
rect 1406 1643 1407 1647
rect 1411 1646 1412 1647
rect 1415 1647 1421 1648
rect 1415 1646 1416 1647
rect 1411 1644 1416 1646
rect 1411 1643 1412 1644
rect 1406 1642 1412 1643
rect 1415 1643 1416 1644
rect 1420 1643 1421 1647
rect 1415 1642 1421 1643
rect 1462 1647 1468 1648
rect 1462 1643 1463 1647
rect 1467 1646 1468 1647
rect 1471 1647 1477 1648
rect 1471 1646 1472 1647
rect 1467 1644 1472 1646
rect 1467 1643 1468 1644
rect 1462 1642 1468 1643
rect 1471 1643 1472 1644
rect 1476 1643 1477 1647
rect 1471 1642 1477 1643
rect 1518 1647 1524 1648
rect 1518 1643 1519 1647
rect 1523 1646 1524 1647
rect 1527 1647 1533 1648
rect 1527 1646 1528 1647
rect 1523 1644 1528 1646
rect 1523 1643 1524 1644
rect 1518 1642 1524 1643
rect 1527 1643 1528 1644
rect 1532 1643 1533 1647
rect 1527 1642 1533 1643
rect 1591 1647 1597 1648
rect 1591 1643 1592 1647
rect 1596 1646 1597 1647
rect 1610 1647 1616 1648
rect 1610 1646 1611 1647
rect 1596 1644 1611 1646
rect 1596 1643 1597 1644
rect 1591 1642 1597 1643
rect 1610 1643 1611 1644
rect 1615 1643 1616 1647
rect 1610 1642 1616 1643
rect 1642 1647 1648 1648
rect 1642 1643 1643 1647
rect 1647 1646 1648 1647
rect 1655 1647 1661 1648
rect 1655 1646 1656 1647
rect 1647 1644 1656 1646
rect 1647 1643 1648 1644
rect 1642 1642 1648 1643
rect 1655 1643 1656 1644
rect 1660 1643 1661 1647
rect 1655 1642 1661 1643
rect 1719 1647 1725 1648
rect 1719 1643 1720 1647
rect 1724 1646 1725 1647
rect 1734 1647 1740 1648
rect 1734 1646 1735 1647
rect 1724 1644 1735 1646
rect 1724 1643 1725 1644
rect 1719 1642 1725 1643
rect 1734 1643 1735 1644
rect 1739 1643 1740 1647
rect 1734 1642 1740 1643
rect 1774 1647 1780 1648
rect 1774 1643 1775 1647
rect 1779 1646 1780 1647
rect 1783 1647 1789 1648
rect 1783 1646 1784 1647
rect 1779 1644 1784 1646
rect 1779 1643 1780 1644
rect 1774 1642 1780 1643
rect 1783 1643 1784 1644
rect 1788 1643 1789 1647
rect 1783 1642 1789 1643
rect 1846 1647 1852 1648
rect 1846 1643 1847 1647
rect 1851 1646 1852 1647
rect 1855 1647 1861 1648
rect 1855 1646 1856 1647
rect 1851 1644 1856 1646
rect 1851 1643 1852 1644
rect 1846 1642 1852 1643
rect 1855 1643 1856 1644
rect 1860 1643 1861 1647
rect 1855 1642 1861 1643
rect 1926 1647 1932 1648
rect 1926 1643 1927 1647
rect 1931 1646 1932 1647
rect 1935 1647 1941 1648
rect 1935 1646 1936 1647
rect 1931 1644 1936 1646
rect 1931 1643 1932 1644
rect 1926 1642 1932 1643
rect 1935 1643 1936 1644
rect 1940 1643 1941 1647
rect 1935 1642 1941 1643
rect 1986 1647 1992 1648
rect 1986 1643 1987 1647
rect 1991 1646 1992 1647
rect 2023 1647 2029 1648
rect 2023 1646 2024 1647
rect 1991 1644 2024 1646
rect 1991 1643 1992 1644
rect 1986 1642 1992 1643
rect 2023 1643 2024 1644
rect 2028 1643 2029 1647
rect 2023 1642 2029 1643
rect 2094 1647 2101 1648
rect 2118 1647 2124 1648
rect 2094 1643 2095 1647
rect 2100 1643 2101 1647
rect 2094 1642 2101 1643
rect 1046 1639 1052 1640
rect 1094 1641 1100 1642
rect 110 1636 116 1637
rect 1094 1637 1095 1641
rect 1099 1637 1100 1641
rect 1094 1636 1100 1637
rect 314 1635 320 1636
rect 314 1634 315 1635
rect 288 1632 315 1634
rect 288 1628 290 1632
rect 314 1631 315 1632
rect 319 1631 320 1635
rect 1134 1635 1140 1636
rect 314 1630 320 1631
rect 1114 1631 1120 1632
rect 1114 1630 1115 1631
rect 1073 1628 1115 1630
rect 158 1627 165 1628
rect 110 1624 116 1625
rect 110 1620 111 1624
rect 115 1620 116 1624
rect 158 1623 159 1627
rect 164 1623 165 1627
rect 158 1622 165 1623
rect 170 1627 176 1628
rect 170 1623 171 1627
rect 175 1626 176 1627
rect 207 1627 213 1628
rect 207 1626 208 1627
rect 175 1624 208 1626
rect 175 1623 176 1624
rect 170 1622 176 1623
rect 207 1623 208 1624
rect 212 1623 213 1627
rect 207 1622 213 1623
rect 287 1627 293 1628
rect 287 1623 288 1627
rect 292 1623 293 1627
rect 287 1622 293 1623
rect 295 1627 301 1628
rect 295 1623 296 1627
rect 300 1626 301 1627
rect 367 1627 373 1628
rect 367 1626 368 1627
rect 300 1624 368 1626
rect 300 1623 301 1624
rect 295 1622 301 1623
rect 367 1623 368 1624
rect 372 1623 373 1627
rect 367 1622 373 1623
rect 375 1627 381 1628
rect 375 1623 376 1627
rect 380 1626 381 1627
rect 447 1627 453 1628
rect 447 1626 448 1627
rect 380 1624 448 1626
rect 380 1623 381 1624
rect 375 1622 381 1623
rect 447 1623 448 1624
rect 452 1623 453 1627
rect 447 1622 453 1623
rect 455 1627 461 1628
rect 455 1623 456 1627
rect 460 1626 461 1627
rect 527 1627 533 1628
rect 527 1626 528 1627
rect 460 1624 528 1626
rect 460 1623 461 1624
rect 455 1622 461 1623
rect 527 1623 528 1624
rect 532 1623 533 1627
rect 527 1622 533 1623
rect 607 1627 613 1628
rect 607 1623 608 1627
rect 612 1626 613 1627
rect 670 1627 676 1628
rect 670 1626 671 1627
rect 612 1624 671 1626
rect 612 1623 613 1624
rect 607 1622 613 1623
rect 670 1623 671 1624
rect 675 1623 676 1627
rect 670 1622 676 1623
rect 679 1627 685 1628
rect 679 1623 680 1627
rect 684 1626 685 1627
rect 751 1627 757 1628
rect 684 1624 747 1626
rect 684 1623 685 1624
rect 679 1622 685 1623
rect 110 1619 116 1620
rect 745 1618 747 1624
rect 751 1623 752 1627
rect 756 1626 757 1627
rect 802 1627 808 1628
rect 802 1626 803 1627
rect 756 1624 803 1626
rect 756 1623 757 1624
rect 751 1622 757 1623
rect 802 1623 803 1624
rect 807 1623 808 1627
rect 802 1622 808 1623
rect 815 1627 821 1628
rect 815 1623 816 1627
rect 820 1626 821 1627
rect 862 1627 868 1628
rect 862 1626 863 1627
rect 820 1624 863 1626
rect 820 1623 821 1624
rect 815 1622 821 1623
rect 862 1623 863 1624
rect 867 1623 868 1627
rect 862 1622 868 1623
rect 870 1627 877 1628
rect 870 1623 871 1627
rect 876 1623 877 1627
rect 870 1622 877 1623
rect 927 1627 936 1628
rect 927 1623 928 1627
rect 935 1623 936 1627
rect 927 1622 936 1623
rect 938 1627 944 1628
rect 938 1623 939 1627
rect 943 1626 944 1627
rect 983 1627 989 1628
rect 983 1626 984 1627
rect 943 1624 984 1626
rect 943 1623 944 1624
rect 938 1622 944 1623
rect 983 1623 984 1624
rect 988 1623 989 1627
rect 983 1622 989 1623
rect 991 1627 997 1628
rect 991 1623 992 1627
rect 996 1626 997 1627
rect 1031 1627 1037 1628
rect 1031 1626 1032 1627
rect 996 1624 1032 1626
rect 996 1623 997 1624
rect 991 1622 997 1623
rect 1031 1623 1032 1624
rect 1036 1623 1037 1627
rect 1031 1622 1037 1623
rect 1071 1627 1077 1628
rect 1071 1623 1072 1627
rect 1076 1623 1077 1627
rect 1114 1627 1115 1628
rect 1119 1627 1120 1631
rect 1134 1631 1135 1635
rect 1139 1631 1140 1635
rect 2118 1635 2124 1636
rect 1134 1630 1140 1631
rect 1262 1632 1268 1633
rect 1262 1628 1263 1632
rect 1267 1628 1268 1632
rect 1262 1627 1268 1628
rect 1302 1632 1308 1633
rect 1302 1628 1303 1632
rect 1307 1628 1308 1632
rect 1302 1627 1308 1628
rect 1342 1632 1348 1633
rect 1342 1628 1343 1632
rect 1347 1628 1348 1632
rect 1342 1627 1348 1628
rect 1390 1632 1396 1633
rect 1390 1628 1391 1632
rect 1395 1628 1396 1632
rect 1390 1627 1396 1628
rect 1446 1632 1452 1633
rect 1446 1628 1447 1632
rect 1451 1628 1452 1632
rect 1446 1627 1452 1628
rect 1502 1632 1508 1633
rect 1502 1628 1503 1632
rect 1507 1628 1508 1632
rect 1502 1627 1508 1628
rect 1566 1632 1572 1633
rect 1566 1628 1567 1632
rect 1571 1628 1572 1632
rect 1566 1627 1572 1628
rect 1630 1632 1636 1633
rect 1630 1628 1631 1632
rect 1635 1628 1636 1632
rect 1630 1627 1636 1628
rect 1694 1632 1700 1633
rect 1694 1628 1695 1632
rect 1699 1628 1700 1632
rect 1694 1627 1700 1628
rect 1758 1632 1764 1633
rect 1758 1628 1759 1632
rect 1763 1628 1764 1632
rect 1758 1627 1764 1628
rect 1830 1632 1836 1633
rect 1830 1628 1831 1632
rect 1835 1628 1836 1632
rect 1830 1627 1836 1628
rect 1910 1632 1916 1633
rect 1910 1628 1911 1632
rect 1915 1628 1916 1632
rect 1910 1627 1916 1628
rect 1998 1632 2004 1633
rect 1998 1628 1999 1632
rect 2003 1628 2004 1632
rect 1998 1627 2004 1628
rect 2070 1632 2076 1633
rect 2070 1628 2071 1632
rect 2075 1628 2076 1632
rect 2118 1631 2119 1635
rect 2123 1631 2124 1635
rect 2118 1630 2124 1631
rect 2070 1627 2076 1628
rect 1114 1626 1120 1627
rect 1071 1622 1077 1623
rect 1094 1624 1100 1625
rect 1094 1620 1095 1624
rect 1099 1620 1100 1624
rect 778 1619 784 1620
rect 1094 1619 1100 1620
rect 778 1618 779 1619
rect 134 1616 140 1617
rect 134 1612 135 1616
rect 139 1612 140 1616
rect 134 1611 140 1612
rect 182 1616 188 1617
rect 182 1612 183 1616
rect 187 1612 188 1616
rect 182 1611 188 1612
rect 262 1616 268 1617
rect 262 1612 263 1616
rect 267 1612 268 1616
rect 262 1611 268 1612
rect 342 1616 348 1617
rect 342 1612 343 1616
rect 347 1612 348 1616
rect 342 1611 348 1612
rect 422 1616 428 1617
rect 422 1612 423 1616
rect 427 1612 428 1616
rect 422 1611 428 1612
rect 502 1616 508 1617
rect 502 1612 503 1616
rect 507 1612 508 1616
rect 502 1611 508 1612
rect 582 1616 588 1617
rect 582 1612 583 1616
rect 587 1612 588 1616
rect 582 1611 588 1612
rect 654 1616 660 1617
rect 654 1612 655 1616
rect 659 1612 660 1616
rect 654 1611 660 1612
rect 726 1616 732 1617
rect 745 1616 779 1618
rect 726 1612 727 1616
rect 731 1612 732 1616
rect 778 1615 779 1616
rect 783 1615 784 1619
rect 778 1614 784 1615
rect 790 1616 796 1617
rect 726 1611 732 1612
rect 790 1612 791 1616
rect 795 1612 796 1616
rect 790 1611 796 1612
rect 846 1616 852 1617
rect 846 1612 847 1616
rect 851 1612 852 1616
rect 846 1611 852 1612
rect 902 1616 908 1617
rect 902 1612 903 1616
rect 907 1612 908 1616
rect 902 1611 908 1612
rect 958 1616 964 1617
rect 958 1612 959 1616
rect 963 1612 964 1616
rect 958 1611 964 1612
rect 1006 1616 1012 1617
rect 1006 1612 1007 1616
rect 1011 1612 1012 1616
rect 1006 1611 1012 1612
rect 1046 1616 1052 1617
rect 1046 1612 1047 1616
rect 1051 1612 1052 1616
rect 1046 1611 1052 1612
rect 1158 1608 1164 1609
rect 159 1607 165 1608
rect 159 1603 160 1607
rect 164 1606 165 1607
rect 170 1607 176 1608
rect 170 1606 171 1607
rect 164 1604 171 1606
rect 164 1603 165 1604
rect 159 1602 165 1603
rect 170 1603 171 1604
rect 175 1603 176 1607
rect 170 1602 176 1603
rect 190 1607 196 1608
rect 190 1603 191 1607
rect 195 1606 196 1607
rect 207 1607 213 1608
rect 207 1606 208 1607
rect 195 1604 208 1606
rect 195 1603 196 1604
rect 190 1602 196 1603
rect 207 1603 208 1604
rect 212 1603 213 1607
rect 207 1602 213 1603
rect 287 1607 293 1608
rect 287 1603 288 1607
rect 292 1606 293 1607
rect 295 1607 301 1608
rect 295 1606 296 1607
rect 292 1604 296 1606
rect 292 1603 293 1604
rect 287 1602 293 1603
rect 295 1603 296 1604
rect 300 1603 301 1607
rect 295 1602 301 1603
rect 367 1607 373 1608
rect 367 1603 368 1607
rect 372 1606 373 1607
rect 375 1607 381 1608
rect 375 1606 376 1607
rect 372 1604 376 1606
rect 372 1603 373 1604
rect 367 1602 373 1603
rect 375 1603 376 1604
rect 380 1603 381 1607
rect 375 1602 381 1603
rect 447 1607 453 1608
rect 447 1603 448 1607
rect 452 1606 453 1607
rect 455 1607 461 1608
rect 455 1606 456 1607
rect 452 1604 456 1606
rect 452 1603 453 1604
rect 447 1602 453 1603
rect 455 1603 456 1604
rect 460 1603 461 1607
rect 455 1602 461 1603
rect 482 1607 488 1608
rect 482 1603 483 1607
rect 487 1606 488 1607
rect 527 1607 533 1608
rect 527 1606 528 1607
rect 487 1604 528 1606
rect 487 1603 488 1604
rect 482 1602 488 1603
rect 527 1603 528 1604
rect 532 1603 533 1607
rect 527 1602 533 1603
rect 607 1607 616 1608
rect 607 1603 608 1607
rect 615 1603 616 1607
rect 607 1602 616 1603
rect 670 1607 676 1608
rect 670 1603 671 1607
rect 675 1606 676 1607
rect 679 1607 685 1608
rect 679 1606 680 1607
rect 675 1604 680 1606
rect 675 1603 676 1604
rect 670 1602 676 1603
rect 679 1603 680 1604
rect 684 1603 685 1607
rect 679 1602 685 1603
rect 751 1607 757 1608
rect 751 1603 752 1607
rect 756 1606 757 1607
rect 766 1607 772 1608
rect 766 1606 767 1607
rect 756 1604 767 1606
rect 756 1603 757 1604
rect 751 1602 757 1603
rect 766 1603 767 1604
rect 771 1603 772 1607
rect 766 1602 772 1603
rect 802 1607 808 1608
rect 802 1603 803 1607
rect 807 1606 808 1607
rect 815 1607 821 1608
rect 815 1606 816 1607
rect 807 1604 816 1606
rect 807 1603 808 1604
rect 802 1602 808 1603
rect 815 1603 816 1604
rect 820 1603 821 1607
rect 815 1602 821 1603
rect 862 1607 868 1608
rect 862 1603 863 1607
rect 867 1606 868 1607
rect 871 1607 877 1608
rect 871 1606 872 1607
rect 867 1604 872 1606
rect 867 1603 868 1604
rect 862 1602 868 1603
rect 871 1603 872 1604
rect 876 1603 877 1607
rect 871 1602 877 1603
rect 927 1607 933 1608
rect 927 1603 928 1607
rect 932 1606 933 1607
rect 938 1607 944 1608
rect 938 1606 939 1607
rect 932 1604 939 1606
rect 932 1603 933 1604
rect 927 1602 933 1603
rect 938 1603 939 1604
rect 943 1603 944 1607
rect 938 1602 944 1603
rect 983 1607 989 1608
rect 983 1603 984 1607
rect 988 1606 989 1607
rect 991 1607 997 1608
rect 991 1606 992 1607
rect 988 1604 992 1606
rect 988 1603 989 1604
rect 983 1602 989 1603
rect 991 1603 992 1604
rect 996 1603 997 1607
rect 991 1602 997 1603
rect 1031 1607 1040 1608
rect 1031 1603 1032 1607
rect 1039 1603 1040 1607
rect 1031 1602 1040 1603
rect 1071 1607 1077 1608
rect 1071 1603 1072 1607
rect 1076 1603 1077 1607
rect 1071 1602 1077 1603
rect 1134 1605 1140 1606
rect 930 1599 936 1600
rect 930 1595 931 1599
rect 935 1598 936 1599
rect 1073 1598 1075 1602
rect 1134 1601 1135 1605
rect 1139 1601 1140 1605
rect 1158 1604 1159 1608
rect 1163 1604 1164 1608
rect 1158 1603 1164 1604
rect 1214 1608 1220 1609
rect 1214 1604 1215 1608
rect 1219 1604 1220 1608
rect 1214 1603 1220 1604
rect 1302 1608 1308 1609
rect 1302 1604 1303 1608
rect 1307 1604 1308 1608
rect 1302 1603 1308 1604
rect 1382 1608 1388 1609
rect 1382 1604 1383 1608
rect 1387 1604 1388 1608
rect 1382 1603 1388 1604
rect 1462 1608 1468 1609
rect 1462 1604 1463 1608
rect 1467 1604 1468 1608
rect 1462 1603 1468 1604
rect 1542 1608 1548 1609
rect 1542 1604 1543 1608
rect 1547 1604 1548 1608
rect 1542 1603 1548 1604
rect 1622 1608 1628 1609
rect 1622 1604 1623 1608
rect 1627 1604 1628 1608
rect 1622 1603 1628 1604
rect 1710 1608 1716 1609
rect 1710 1604 1711 1608
rect 1715 1604 1716 1608
rect 1710 1603 1716 1604
rect 1798 1608 1804 1609
rect 1798 1604 1799 1608
rect 1803 1604 1804 1608
rect 1798 1603 1804 1604
rect 1886 1608 1892 1609
rect 1886 1604 1887 1608
rect 1891 1604 1892 1608
rect 1886 1603 1892 1604
rect 1982 1608 1988 1609
rect 1982 1604 1983 1608
rect 1987 1604 1988 1608
rect 1982 1603 1988 1604
rect 2070 1608 2076 1609
rect 2070 1604 2071 1608
rect 2075 1604 2076 1608
rect 2070 1603 2076 1604
rect 2118 1605 2124 1606
rect 1134 1600 1140 1601
rect 2118 1601 2119 1605
rect 2123 1601 2124 1605
rect 2118 1600 2124 1601
rect 1614 1599 1620 1600
rect 1614 1598 1615 1599
rect 935 1596 1075 1598
rect 1488 1596 1615 1598
rect 935 1595 936 1596
rect 930 1594 936 1595
rect 1488 1592 1490 1596
rect 1614 1595 1615 1596
rect 1619 1595 1620 1599
rect 1614 1594 1620 1595
rect 1183 1591 1189 1592
rect 1134 1588 1140 1589
rect 158 1587 165 1588
rect 158 1583 159 1587
rect 164 1583 165 1587
rect 158 1582 165 1583
rect 182 1587 188 1588
rect 182 1583 183 1587
rect 187 1586 188 1587
rect 199 1587 205 1588
rect 199 1586 200 1587
rect 187 1584 200 1586
rect 187 1583 188 1584
rect 182 1582 188 1583
rect 199 1583 200 1584
rect 204 1583 205 1587
rect 199 1582 205 1583
rect 207 1587 213 1588
rect 207 1583 208 1587
rect 212 1586 213 1587
rect 255 1587 261 1588
rect 255 1586 256 1587
rect 212 1584 256 1586
rect 212 1583 213 1584
rect 207 1582 213 1583
rect 255 1583 256 1584
rect 260 1583 261 1587
rect 255 1582 261 1583
rect 287 1587 293 1588
rect 287 1583 288 1587
rect 292 1586 293 1587
rect 327 1587 333 1588
rect 327 1586 328 1587
rect 292 1584 328 1586
rect 292 1583 293 1584
rect 287 1582 293 1583
rect 327 1583 328 1584
rect 332 1583 333 1587
rect 327 1582 333 1583
rect 335 1587 341 1588
rect 335 1583 336 1587
rect 340 1586 341 1587
rect 399 1587 405 1588
rect 399 1586 400 1587
rect 340 1584 400 1586
rect 340 1583 341 1584
rect 335 1582 341 1583
rect 399 1583 400 1584
rect 404 1583 405 1587
rect 399 1582 405 1583
rect 407 1587 413 1588
rect 407 1583 408 1587
rect 412 1586 413 1587
rect 479 1587 485 1588
rect 479 1586 480 1587
rect 412 1584 480 1586
rect 412 1583 413 1584
rect 407 1582 413 1583
rect 479 1583 480 1584
rect 484 1583 485 1587
rect 479 1582 485 1583
rect 551 1587 557 1588
rect 551 1583 552 1587
rect 556 1586 557 1587
rect 590 1587 596 1588
rect 590 1586 591 1587
rect 556 1584 591 1586
rect 556 1583 557 1584
rect 551 1582 557 1583
rect 590 1583 591 1584
rect 595 1583 596 1587
rect 590 1582 596 1583
rect 606 1587 612 1588
rect 606 1583 607 1587
rect 611 1586 612 1587
rect 623 1587 629 1588
rect 623 1586 624 1587
rect 611 1584 624 1586
rect 611 1583 612 1584
rect 606 1582 612 1583
rect 623 1583 624 1584
rect 628 1583 629 1587
rect 623 1582 629 1583
rect 631 1587 637 1588
rect 631 1583 632 1587
rect 636 1586 637 1587
rect 695 1587 701 1588
rect 695 1586 696 1587
rect 636 1584 696 1586
rect 636 1583 637 1584
rect 631 1582 637 1583
rect 695 1583 696 1584
rect 700 1583 701 1587
rect 695 1582 701 1583
rect 706 1587 712 1588
rect 706 1583 707 1587
rect 711 1586 712 1587
rect 767 1587 773 1588
rect 767 1586 768 1587
rect 711 1584 768 1586
rect 711 1583 712 1584
rect 706 1582 712 1583
rect 767 1583 768 1584
rect 772 1583 773 1587
rect 767 1582 773 1583
rect 778 1587 784 1588
rect 778 1583 779 1587
rect 783 1586 784 1587
rect 839 1587 845 1588
rect 839 1586 840 1587
rect 783 1584 840 1586
rect 783 1583 784 1584
rect 778 1582 784 1583
rect 839 1583 840 1584
rect 844 1583 845 1587
rect 911 1587 917 1588
rect 911 1586 912 1587
rect 839 1582 845 1583
rect 848 1584 912 1586
rect 134 1580 140 1581
rect 134 1576 135 1580
rect 139 1576 140 1580
rect 134 1575 140 1576
rect 174 1580 180 1581
rect 174 1576 175 1580
rect 179 1576 180 1580
rect 174 1575 180 1576
rect 230 1580 236 1581
rect 230 1576 231 1580
rect 235 1576 236 1580
rect 230 1575 236 1576
rect 302 1580 308 1581
rect 302 1576 303 1580
rect 307 1576 308 1580
rect 302 1575 308 1576
rect 374 1580 380 1581
rect 374 1576 375 1580
rect 379 1576 380 1580
rect 374 1575 380 1576
rect 454 1580 460 1581
rect 454 1576 455 1580
rect 459 1576 460 1580
rect 454 1575 460 1576
rect 526 1580 532 1581
rect 526 1576 527 1580
rect 531 1576 532 1580
rect 526 1575 532 1576
rect 598 1580 604 1581
rect 598 1576 599 1580
rect 603 1576 604 1580
rect 598 1575 604 1576
rect 670 1580 676 1581
rect 670 1576 671 1580
rect 675 1576 676 1580
rect 670 1575 676 1576
rect 742 1580 748 1581
rect 742 1576 743 1580
rect 747 1576 748 1580
rect 742 1575 748 1576
rect 814 1580 820 1581
rect 814 1576 815 1580
rect 819 1576 820 1580
rect 814 1575 820 1576
rect 848 1574 850 1584
rect 911 1583 912 1584
rect 916 1583 917 1587
rect 1134 1584 1135 1588
rect 1139 1584 1140 1588
rect 1183 1587 1184 1591
rect 1188 1590 1189 1591
rect 1230 1591 1236 1592
rect 1230 1590 1231 1591
rect 1188 1588 1231 1590
rect 1188 1587 1189 1588
rect 1183 1586 1189 1587
rect 1230 1587 1231 1588
rect 1235 1587 1236 1591
rect 1230 1586 1236 1587
rect 1239 1591 1245 1592
rect 1239 1587 1240 1591
rect 1244 1590 1245 1591
rect 1318 1591 1324 1592
rect 1318 1590 1319 1591
rect 1244 1588 1319 1590
rect 1244 1587 1245 1588
rect 1239 1586 1245 1587
rect 1318 1587 1319 1588
rect 1323 1587 1324 1591
rect 1318 1586 1324 1587
rect 1327 1591 1333 1592
rect 1327 1587 1328 1591
rect 1332 1590 1333 1591
rect 1398 1591 1404 1592
rect 1398 1590 1399 1591
rect 1332 1588 1399 1590
rect 1332 1587 1333 1588
rect 1327 1586 1333 1587
rect 1398 1587 1399 1588
rect 1403 1587 1404 1591
rect 1398 1586 1404 1587
rect 1407 1591 1413 1592
rect 1407 1587 1408 1591
rect 1412 1590 1413 1591
rect 1487 1591 1493 1592
rect 1412 1588 1474 1590
rect 1412 1587 1413 1588
rect 1407 1586 1413 1587
rect 1134 1583 1140 1584
rect 911 1582 917 1583
rect 1472 1582 1474 1588
rect 1487 1587 1488 1591
rect 1492 1587 1493 1591
rect 1487 1586 1493 1587
rect 1495 1591 1501 1592
rect 1495 1587 1496 1591
rect 1500 1590 1501 1591
rect 1567 1591 1573 1592
rect 1567 1590 1568 1591
rect 1500 1588 1568 1590
rect 1500 1587 1501 1588
rect 1495 1586 1501 1587
rect 1567 1587 1568 1588
rect 1572 1587 1573 1591
rect 1567 1586 1573 1587
rect 1647 1591 1656 1592
rect 1647 1587 1648 1591
rect 1655 1587 1656 1591
rect 1647 1586 1656 1587
rect 1735 1591 1741 1592
rect 1735 1587 1736 1591
rect 1740 1590 1741 1591
rect 1774 1591 1780 1592
rect 1774 1590 1775 1591
rect 1740 1588 1775 1590
rect 1740 1587 1741 1588
rect 1735 1586 1741 1587
rect 1774 1587 1775 1588
rect 1779 1587 1780 1591
rect 1774 1586 1780 1587
rect 1782 1591 1788 1592
rect 1782 1587 1783 1591
rect 1787 1590 1788 1591
rect 1823 1591 1829 1592
rect 1823 1590 1824 1591
rect 1787 1588 1824 1590
rect 1787 1587 1788 1588
rect 1782 1586 1788 1587
rect 1823 1587 1824 1588
rect 1828 1587 1829 1591
rect 1823 1586 1829 1587
rect 1831 1591 1837 1592
rect 1831 1587 1832 1591
rect 1836 1590 1837 1591
rect 1911 1591 1917 1592
rect 1911 1590 1912 1591
rect 1836 1588 1912 1590
rect 1836 1587 1837 1588
rect 1831 1586 1837 1587
rect 1911 1587 1912 1588
rect 1916 1587 1917 1591
rect 1911 1586 1917 1587
rect 2007 1591 2016 1592
rect 2007 1587 2008 1591
rect 2015 1587 2016 1591
rect 2007 1586 2016 1587
rect 2095 1591 2101 1592
rect 2095 1587 2096 1591
rect 2100 1590 2101 1591
rect 2103 1591 2109 1592
rect 2103 1590 2104 1591
rect 2100 1588 2104 1590
rect 2100 1587 2101 1588
rect 2095 1586 2101 1587
rect 2103 1587 2104 1588
rect 2108 1587 2109 1591
rect 2103 1586 2109 1587
rect 2118 1588 2124 1589
rect 2118 1584 2119 1588
rect 2123 1584 2124 1588
rect 1502 1583 1508 1584
rect 2118 1583 2124 1584
rect 1502 1582 1503 1583
rect 886 1580 892 1581
rect 886 1576 887 1580
rect 891 1576 892 1580
rect 886 1575 892 1576
rect 1158 1580 1164 1581
rect 1158 1576 1159 1580
rect 1163 1576 1164 1580
rect 1158 1575 1164 1576
rect 1214 1580 1220 1581
rect 1214 1576 1215 1580
rect 1219 1576 1220 1580
rect 1214 1575 1220 1576
rect 1302 1580 1308 1581
rect 1302 1576 1303 1580
rect 1307 1576 1308 1580
rect 1302 1575 1308 1576
rect 1382 1580 1388 1581
rect 1382 1576 1383 1580
rect 1387 1576 1388 1580
rect 1382 1575 1388 1576
rect 1462 1580 1468 1581
rect 1472 1580 1503 1582
rect 1462 1576 1463 1580
rect 1467 1576 1468 1580
rect 1502 1579 1503 1580
rect 1507 1579 1508 1583
rect 1502 1578 1508 1579
rect 1542 1580 1548 1581
rect 1462 1575 1468 1576
rect 1542 1576 1543 1580
rect 1547 1576 1548 1580
rect 1542 1575 1548 1576
rect 1622 1580 1628 1581
rect 1622 1576 1623 1580
rect 1627 1576 1628 1580
rect 1622 1575 1628 1576
rect 1710 1580 1716 1581
rect 1710 1576 1711 1580
rect 1715 1576 1716 1580
rect 1710 1575 1716 1576
rect 1798 1580 1804 1581
rect 1798 1576 1799 1580
rect 1803 1576 1804 1580
rect 1798 1575 1804 1576
rect 1886 1580 1892 1581
rect 1886 1576 1887 1580
rect 1891 1576 1892 1580
rect 1886 1575 1892 1576
rect 1982 1580 1988 1581
rect 1982 1576 1983 1580
rect 1987 1576 1988 1580
rect 1982 1575 1988 1576
rect 2070 1580 2076 1581
rect 2070 1576 2071 1580
rect 2075 1576 2076 1580
rect 2070 1575 2076 1576
rect 110 1572 116 1573
rect 110 1568 111 1572
rect 115 1568 116 1572
rect 844 1572 850 1574
rect 1094 1572 1100 1573
rect 844 1568 846 1572
rect 1094 1568 1095 1572
rect 1099 1568 1100 1572
rect 110 1567 116 1568
rect 159 1567 165 1568
rect 159 1563 160 1567
rect 164 1566 165 1567
rect 182 1567 188 1568
rect 182 1566 183 1567
rect 164 1564 183 1566
rect 164 1563 165 1564
rect 159 1562 165 1563
rect 182 1563 183 1564
rect 187 1563 188 1567
rect 182 1562 188 1563
rect 199 1567 205 1568
rect 199 1563 200 1567
rect 204 1566 205 1567
rect 207 1567 213 1568
rect 207 1566 208 1567
rect 204 1564 208 1566
rect 204 1563 205 1564
rect 199 1562 205 1563
rect 207 1563 208 1564
rect 212 1563 213 1567
rect 207 1562 213 1563
rect 215 1567 221 1568
rect 215 1563 216 1567
rect 220 1566 221 1567
rect 255 1567 261 1568
rect 255 1566 256 1567
rect 220 1564 256 1566
rect 220 1563 221 1564
rect 215 1562 221 1563
rect 255 1563 256 1564
rect 260 1563 261 1567
rect 255 1562 261 1563
rect 327 1567 333 1568
rect 327 1563 328 1567
rect 332 1566 333 1567
rect 335 1567 341 1568
rect 335 1566 336 1567
rect 332 1564 336 1566
rect 332 1563 333 1564
rect 327 1562 333 1563
rect 335 1563 336 1564
rect 340 1563 341 1567
rect 335 1562 341 1563
rect 399 1567 405 1568
rect 399 1563 400 1567
rect 404 1566 405 1567
rect 407 1567 413 1568
rect 407 1566 408 1567
rect 404 1564 408 1566
rect 404 1563 405 1564
rect 399 1562 405 1563
rect 407 1563 408 1564
rect 412 1563 413 1567
rect 407 1562 413 1563
rect 479 1567 488 1568
rect 479 1563 480 1567
rect 487 1563 488 1567
rect 479 1562 488 1563
rect 551 1567 557 1568
rect 551 1563 552 1567
rect 556 1566 557 1567
rect 606 1567 612 1568
rect 606 1566 607 1567
rect 556 1564 607 1566
rect 556 1563 557 1564
rect 551 1562 557 1563
rect 606 1563 607 1564
rect 611 1563 612 1567
rect 606 1562 612 1563
rect 623 1567 629 1568
rect 623 1563 624 1567
rect 628 1566 629 1567
rect 631 1567 637 1568
rect 631 1566 632 1567
rect 628 1564 632 1566
rect 628 1563 629 1564
rect 623 1562 629 1563
rect 631 1563 632 1564
rect 636 1563 637 1567
rect 631 1562 637 1563
rect 695 1567 701 1568
rect 695 1563 696 1567
rect 700 1566 701 1567
rect 706 1567 712 1568
rect 706 1566 707 1567
rect 700 1564 707 1566
rect 700 1563 701 1564
rect 695 1562 701 1563
rect 706 1563 707 1564
rect 711 1563 712 1567
rect 706 1562 712 1563
rect 766 1567 773 1568
rect 766 1563 767 1567
rect 772 1563 773 1567
rect 766 1562 773 1563
rect 839 1567 846 1568
rect 839 1563 840 1567
rect 844 1564 846 1567
rect 850 1567 856 1568
rect 844 1563 845 1564
rect 839 1562 845 1563
rect 850 1563 851 1567
rect 855 1566 856 1567
rect 911 1567 917 1568
rect 1094 1567 1100 1568
rect 1114 1571 1120 1572
rect 1114 1567 1115 1571
rect 1119 1570 1120 1571
rect 1183 1571 1189 1572
rect 1183 1570 1184 1571
rect 1119 1568 1184 1570
rect 1119 1567 1120 1568
rect 911 1566 912 1567
rect 855 1564 912 1566
rect 855 1563 856 1564
rect 850 1562 856 1563
rect 911 1563 912 1564
rect 916 1563 917 1567
rect 1114 1566 1120 1567
rect 1183 1567 1184 1568
rect 1188 1567 1189 1571
rect 1183 1566 1189 1567
rect 1230 1571 1236 1572
rect 1230 1567 1231 1571
rect 1235 1570 1236 1571
rect 1239 1571 1245 1572
rect 1239 1570 1240 1571
rect 1235 1568 1240 1570
rect 1235 1567 1236 1568
rect 1230 1566 1236 1567
rect 1239 1567 1240 1568
rect 1244 1567 1245 1571
rect 1239 1566 1245 1567
rect 1318 1571 1324 1572
rect 1318 1567 1319 1571
rect 1323 1570 1324 1571
rect 1327 1571 1333 1572
rect 1327 1570 1328 1571
rect 1323 1568 1328 1570
rect 1323 1567 1324 1568
rect 1318 1566 1324 1567
rect 1327 1567 1328 1568
rect 1332 1567 1333 1571
rect 1327 1566 1333 1567
rect 1398 1571 1404 1572
rect 1398 1567 1399 1571
rect 1403 1570 1404 1571
rect 1407 1571 1413 1572
rect 1407 1570 1408 1571
rect 1403 1568 1408 1570
rect 1403 1567 1404 1568
rect 1398 1566 1404 1567
rect 1407 1567 1408 1568
rect 1412 1567 1413 1571
rect 1407 1566 1413 1567
rect 1487 1571 1493 1572
rect 1487 1567 1488 1571
rect 1492 1570 1493 1571
rect 1495 1571 1501 1572
rect 1495 1570 1496 1571
rect 1492 1568 1496 1570
rect 1492 1567 1493 1568
rect 1487 1566 1493 1567
rect 1495 1567 1496 1568
rect 1500 1567 1501 1571
rect 1495 1566 1501 1567
rect 1567 1571 1573 1572
rect 1567 1567 1568 1571
rect 1572 1570 1573 1571
rect 1582 1571 1588 1572
rect 1582 1570 1583 1571
rect 1572 1568 1583 1570
rect 1572 1567 1573 1568
rect 1567 1566 1573 1567
rect 1582 1567 1583 1568
rect 1587 1567 1588 1571
rect 1582 1566 1588 1567
rect 1614 1571 1620 1572
rect 1614 1567 1615 1571
rect 1619 1570 1620 1571
rect 1647 1571 1653 1572
rect 1647 1570 1648 1571
rect 1619 1568 1648 1570
rect 1619 1567 1620 1568
rect 1614 1566 1620 1567
rect 1647 1567 1648 1568
rect 1652 1567 1653 1571
rect 1647 1566 1653 1567
rect 1734 1571 1741 1572
rect 1734 1567 1735 1571
rect 1740 1567 1741 1571
rect 1734 1566 1741 1567
rect 1823 1571 1829 1572
rect 1823 1567 1824 1571
rect 1828 1570 1829 1571
rect 1831 1571 1837 1572
rect 1831 1570 1832 1571
rect 1828 1568 1832 1570
rect 1828 1567 1829 1568
rect 1823 1566 1829 1567
rect 1831 1567 1832 1568
rect 1836 1567 1837 1571
rect 1831 1566 1837 1567
rect 1911 1571 1917 1572
rect 1911 1567 1912 1571
rect 1916 1567 1917 1571
rect 1911 1566 1917 1567
rect 1946 1571 1952 1572
rect 1946 1567 1947 1571
rect 1951 1570 1952 1571
rect 2007 1571 2013 1572
rect 2007 1570 2008 1571
rect 1951 1568 2008 1570
rect 1951 1567 1952 1568
rect 1946 1566 1952 1567
rect 2007 1567 2008 1568
rect 2012 1567 2013 1571
rect 2007 1566 2013 1567
rect 2094 1571 2101 1572
rect 2094 1567 2095 1571
rect 2100 1567 2101 1571
rect 2094 1566 2101 1567
rect 911 1562 917 1563
rect 1774 1563 1780 1564
rect 1774 1559 1775 1563
rect 1779 1562 1780 1563
rect 1913 1562 1915 1566
rect 1779 1560 1915 1562
rect 1779 1559 1780 1560
rect 1774 1558 1780 1559
rect 110 1555 116 1556
rect 110 1551 111 1555
rect 115 1551 116 1555
rect 1094 1555 1100 1556
rect 110 1550 116 1551
rect 134 1552 140 1553
rect 134 1548 135 1552
rect 139 1548 140 1552
rect 134 1547 140 1548
rect 174 1552 180 1553
rect 174 1548 175 1552
rect 179 1548 180 1552
rect 174 1547 180 1548
rect 230 1552 236 1553
rect 230 1548 231 1552
rect 235 1548 236 1552
rect 230 1547 236 1548
rect 302 1552 308 1553
rect 302 1548 303 1552
rect 307 1548 308 1552
rect 302 1547 308 1548
rect 374 1552 380 1553
rect 374 1548 375 1552
rect 379 1548 380 1552
rect 374 1547 380 1548
rect 454 1552 460 1553
rect 454 1548 455 1552
rect 459 1548 460 1552
rect 454 1547 460 1548
rect 526 1552 532 1553
rect 526 1548 527 1552
rect 531 1548 532 1552
rect 526 1547 532 1548
rect 598 1552 604 1553
rect 598 1548 599 1552
rect 603 1548 604 1552
rect 598 1547 604 1548
rect 670 1552 676 1553
rect 670 1548 671 1552
rect 675 1548 676 1552
rect 670 1547 676 1548
rect 742 1552 748 1553
rect 742 1548 743 1552
rect 747 1548 748 1552
rect 742 1547 748 1548
rect 814 1552 820 1553
rect 814 1548 815 1552
rect 819 1548 820 1552
rect 814 1547 820 1548
rect 886 1552 892 1553
rect 886 1548 887 1552
rect 891 1548 892 1552
rect 1094 1551 1095 1555
rect 1099 1551 1100 1555
rect 1094 1550 1100 1551
rect 1183 1551 1189 1552
rect 886 1547 892 1548
rect 1183 1547 1184 1551
rect 1188 1550 1189 1551
rect 1214 1551 1220 1552
rect 1214 1550 1215 1551
rect 1188 1548 1215 1550
rect 1188 1547 1189 1548
rect 1183 1546 1189 1547
rect 1214 1547 1215 1548
rect 1219 1547 1220 1551
rect 1214 1546 1220 1547
rect 1223 1551 1229 1552
rect 1223 1547 1224 1551
rect 1228 1550 1229 1551
rect 1254 1551 1260 1552
rect 1254 1550 1255 1551
rect 1228 1548 1255 1550
rect 1228 1547 1229 1548
rect 1223 1546 1229 1547
rect 1254 1547 1255 1548
rect 1259 1547 1260 1551
rect 1254 1546 1260 1547
rect 1271 1551 1277 1552
rect 1271 1547 1272 1551
rect 1276 1550 1277 1551
rect 1334 1551 1340 1552
rect 1334 1550 1335 1551
rect 1276 1548 1335 1550
rect 1276 1547 1277 1548
rect 1271 1546 1277 1547
rect 1334 1547 1335 1548
rect 1339 1547 1340 1551
rect 1334 1546 1340 1547
rect 1343 1551 1349 1552
rect 1343 1547 1344 1551
rect 1348 1550 1349 1551
rect 1414 1551 1420 1552
rect 1414 1550 1415 1551
rect 1348 1548 1415 1550
rect 1348 1547 1349 1548
rect 1343 1546 1349 1547
rect 1414 1547 1415 1548
rect 1419 1547 1420 1551
rect 1414 1546 1420 1547
rect 1423 1551 1429 1552
rect 1423 1547 1424 1551
rect 1428 1550 1429 1551
rect 1494 1551 1500 1552
rect 1494 1550 1495 1551
rect 1428 1548 1495 1550
rect 1428 1547 1429 1548
rect 1423 1546 1429 1547
rect 1494 1547 1495 1548
rect 1499 1547 1500 1551
rect 1494 1546 1500 1547
rect 1502 1551 1509 1552
rect 1502 1547 1503 1551
rect 1508 1547 1509 1551
rect 1502 1546 1509 1547
rect 1583 1551 1589 1552
rect 1583 1547 1584 1551
rect 1588 1550 1589 1551
rect 1662 1551 1668 1552
rect 1662 1550 1663 1551
rect 1588 1548 1663 1550
rect 1588 1547 1589 1548
rect 1583 1546 1589 1547
rect 1662 1547 1663 1548
rect 1667 1547 1668 1551
rect 1662 1546 1668 1547
rect 1671 1551 1677 1552
rect 1671 1547 1672 1551
rect 1676 1550 1677 1551
rect 1750 1551 1756 1552
rect 1750 1550 1751 1551
rect 1676 1548 1751 1550
rect 1676 1547 1677 1548
rect 1671 1546 1677 1547
rect 1750 1547 1751 1548
rect 1755 1547 1756 1551
rect 1750 1546 1756 1547
rect 1759 1551 1765 1552
rect 1759 1547 1760 1551
rect 1764 1550 1765 1551
rect 1782 1551 1788 1552
rect 1782 1550 1783 1551
rect 1764 1548 1783 1550
rect 1764 1547 1765 1548
rect 1759 1546 1765 1547
rect 1782 1547 1783 1548
rect 1787 1547 1788 1551
rect 1782 1546 1788 1547
rect 1798 1551 1804 1552
rect 1798 1547 1799 1551
rect 1803 1550 1804 1551
rect 1847 1551 1853 1552
rect 1847 1550 1848 1551
rect 1803 1548 1848 1550
rect 1803 1547 1804 1548
rect 1798 1546 1804 1547
rect 1847 1547 1848 1548
rect 1852 1547 1853 1551
rect 1847 1546 1853 1547
rect 1855 1551 1861 1552
rect 1855 1547 1856 1551
rect 1860 1550 1861 1551
rect 1935 1551 1941 1552
rect 1935 1550 1936 1551
rect 1860 1548 1936 1550
rect 1860 1547 1861 1548
rect 1855 1546 1861 1547
rect 1935 1547 1936 1548
rect 1940 1547 1941 1551
rect 1935 1546 1941 1547
rect 1943 1551 1949 1552
rect 1943 1547 1944 1551
rect 1948 1550 1949 1551
rect 2023 1551 2029 1552
rect 2023 1550 2024 1551
rect 1948 1548 2024 1550
rect 1948 1547 1949 1548
rect 1943 1546 1949 1547
rect 2023 1547 2024 1548
rect 2028 1547 2029 1551
rect 2023 1546 2029 1547
rect 2095 1551 2101 1552
rect 2095 1547 2096 1551
rect 2100 1550 2101 1551
rect 2103 1551 2109 1552
rect 2103 1550 2104 1551
rect 2100 1548 2104 1550
rect 2100 1547 2101 1548
rect 2095 1546 2101 1547
rect 2103 1547 2104 1548
rect 2108 1547 2109 1551
rect 2103 1546 2109 1547
rect 1158 1544 1164 1545
rect 134 1540 140 1541
rect 110 1537 116 1538
rect 110 1533 111 1537
rect 115 1533 116 1537
rect 134 1536 135 1540
rect 139 1536 140 1540
rect 134 1535 140 1536
rect 174 1540 180 1541
rect 174 1536 175 1540
rect 179 1536 180 1540
rect 174 1535 180 1536
rect 230 1540 236 1541
rect 230 1536 231 1540
rect 235 1536 236 1540
rect 230 1535 236 1536
rect 310 1540 316 1541
rect 310 1536 311 1540
rect 315 1536 316 1540
rect 310 1535 316 1536
rect 390 1540 396 1541
rect 390 1536 391 1540
rect 395 1536 396 1540
rect 390 1535 396 1536
rect 478 1540 484 1541
rect 478 1536 479 1540
rect 483 1536 484 1540
rect 478 1535 484 1536
rect 566 1540 572 1541
rect 566 1536 567 1540
rect 571 1536 572 1540
rect 566 1535 572 1536
rect 654 1540 660 1541
rect 654 1536 655 1540
rect 659 1536 660 1540
rect 654 1535 660 1536
rect 742 1540 748 1541
rect 742 1536 743 1540
rect 747 1536 748 1540
rect 742 1535 748 1536
rect 822 1540 828 1541
rect 822 1536 823 1540
rect 827 1536 828 1540
rect 822 1535 828 1536
rect 910 1540 916 1541
rect 910 1536 911 1540
rect 915 1536 916 1540
rect 910 1535 916 1536
rect 998 1540 1004 1541
rect 998 1536 999 1540
rect 1003 1536 1004 1540
rect 1158 1540 1159 1544
rect 1163 1540 1164 1544
rect 1158 1539 1164 1540
rect 1198 1544 1204 1545
rect 1198 1540 1199 1544
rect 1203 1540 1204 1544
rect 1198 1539 1204 1540
rect 1246 1544 1252 1545
rect 1246 1540 1247 1544
rect 1251 1540 1252 1544
rect 1246 1539 1252 1540
rect 1318 1544 1324 1545
rect 1318 1540 1319 1544
rect 1323 1540 1324 1544
rect 1318 1539 1324 1540
rect 1398 1544 1404 1545
rect 1398 1540 1399 1544
rect 1403 1540 1404 1544
rect 1398 1539 1404 1540
rect 1478 1544 1484 1545
rect 1478 1540 1479 1544
rect 1483 1540 1484 1544
rect 1478 1539 1484 1540
rect 1558 1544 1564 1545
rect 1558 1540 1559 1544
rect 1563 1540 1564 1544
rect 1558 1539 1564 1540
rect 1646 1544 1652 1545
rect 1646 1540 1647 1544
rect 1651 1540 1652 1544
rect 1646 1539 1652 1540
rect 1734 1544 1740 1545
rect 1734 1540 1735 1544
rect 1739 1540 1740 1544
rect 1734 1539 1740 1540
rect 1822 1544 1828 1545
rect 1822 1540 1823 1544
rect 1827 1540 1828 1544
rect 1822 1539 1828 1540
rect 1910 1544 1916 1545
rect 1910 1540 1911 1544
rect 1915 1540 1916 1544
rect 1910 1539 1916 1540
rect 1998 1544 2004 1545
rect 1998 1540 1999 1544
rect 2003 1540 2004 1544
rect 1998 1539 2004 1540
rect 2070 1544 2076 1545
rect 2070 1540 2071 1544
rect 2075 1540 2076 1544
rect 2070 1539 2076 1540
rect 998 1535 1004 1536
rect 1094 1537 1100 1538
rect 110 1532 116 1533
rect 1094 1533 1095 1537
rect 1099 1533 1100 1537
rect 1094 1532 1100 1533
rect 1134 1536 1140 1537
rect 1134 1532 1135 1536
rect 1139 1532 1140 1536
rect 2118 1536 2124 1537
rect 2118 1532 2119 1536
rect 2123 1532 2124 1536
rect 287 1531 293 1532
rect 1134 1531 1140 1532
rect 1182 1531 1189 1532
rect 287 1530 288 1531
rect 257 1528 288 1530
rect 257 1524 259 1528
rect 287 1527 288 1528
rect 292 1527 293 1531
rect 287 1526 293 1527
rect 1182 1527 1183 1531
rect 1188 1527 1189 1531
rect 1182 1526 1189 1527
rect 1214 1531 1220 1532
rect 1214 1527 1215 1531
rect 1219 1530 1220 1531
rect 1223 1531 1229 1532
rect 1223 1530 1224 1531
rect 1219 1528 1224 1530
rect 1219 1527 1220 1528
rect 1214 1526 1220 1527
rect 1223 1527 1224 1528
rect 1228 1527 1229 1531
rect 1223 1526 1229 1527
rect 1254 1531 1260 1532
rect 1254 1527 1255 1531
rect 1259 1530 1260 1531
rect 1271 1531 1277 1532
rect 1271 1530 1272 1531
rect 1259 1528 1272 1530
rect 1259 1527 1260 1528
rect 1254 1526 1260 1527
rect 1271 1527 1272 1528
rect 1276 1527 1277 1531
rect 1271 1526 1277 1527
rect 1334 1531 1340 1532
rect 1334 1527 1335 1531
rect 1339 1530 1340 1531
rect 1343 1531 1349 1532
rect 1343 1530 1344 1531
rect 1339 1528 1344 1530
rect 1339 1527 1340 1528
rect 1334 1526 1340 1527
rect 1343 1527 1344 1528
rect 1348 1527 1349 1531
rect 1343 1526 1349 1527
rect 1414 1531 1420 1532
rect 1414 1527 1415 1531
rect 1419 1530 1420 1531
rect 1423 1531 1429 1532
rect 1423 1530 1424 1531
rect 1419 1528 1424 1530
rect 1419 1527 1420 1528
rect 1414 1526 1420 1527
rect 1423 1527 1424 1528
rect 1428 1527 1429 1531
rect 1423 1526 1429 1527
rect 1494 1531 1500 1532
rect 1494 1527 1495 1531
rect 1499 1530 1500 1531
rect 1503 1531 1509 1532
rect 1503 1530 1504 1531
rect 1499 1528 1504 1530
rect 1499 1527 1500 1528
rect 1494 1526 1500 1527
rect 1503 1527 1504 1528
rect 1508 1527 1509 1531
rect 1503 1526 1509 1527
rect 1582 1531 1589 1532
rect 1582 1527 1583 1531
rect 1588 1527 1589 1531
rect 1582 1526 1589 1527
rect 1662 1531 1668 1532
rect 1662 1527 1663 1531
rect 1667 1530 1668 1531
rect 1671 1531 1677 1532
rect 1671 1530 1672 1531
rect 1667 1528 1672 1530
rect 1667 1527 1668 1528
rect 1662 1526 1668 1527
rect 1671 1527 1672 1528
rect 1676 1527 1677 1531
rect 1671 1526 1677 1527
rect 1750 1531 1756 1532
rect 1750 1527 1751 1531
rect 1755 1530 1756 1531
rect 1759 1531 1765 1532
rect 1759 1530 1760 1531
rect 1755 1528 1760 1530
rect 1755 1527 1756 1528
rect 1750 1526 1756 1527
rect 1759 1527 1760 1528
rect 1764 1527 1765 1531
rect 1759 1526 1765 1527
rect 1847 1531 1853 1532
rect 1847 1527 1848 1531
rect 1852 1530 1853 1531
rect 1855 1531 1861 1532
rect 1855 1530 1856 1531
rect 1852 1528 1856 1530
rect 1852 1527 1853 1528
rect 1847 1526 1853 1527
rect 1855 1527 1856 1528
rect 1860 1527 1861 1531
rect 1855 1526 1861 1527
rect 1935 1531 1941 1532
rect 1935 1527 1936 1531
rect 1940 1530 1941 1531
rect 1943 1531 1949 1532
rect 1943 1530 1944 1531
rect 1940 1528 1944 1530
rect 1940 1527 1941 1528
rect 1935 1526 1941 1527
rect 1943 1527 1944 1528
rect 1948 1527 1949 1531
rect 1943 1526 1949 1527
rect 2018 1531 2029 1532
rect 2018 1527 2019 1531
rect 2023 1527 2024 1531
rect 2028 1527 2029 1531
rect 2018 1526 2029 1527
rect 2038 1531 2044 1532
rect 2038 1527 2039 1531
rect 2043 1530 2044 1531
rect 2095 1531 2101 1532
rect 2118 1531 2124 1532
rect 2095 1530 2096 1531
rect 2043 1528 2096 1530
rect 2043 1527 2044 1528
rect 2038 1526 2044 1527
rect 2095 1527 2096 1528
rect 2100 1527 2101 1531
rect 2095 1526 2101 1527
rect 159 1523 168 1524
rect 110 1520 116 1521
rect 110 1516 111 1520
rect 115 1516 116 1520
rect 159 1519 160 1523
rect 167 1519 168 1523
rect 159 1518 168 1519
rect 182 1523 188 1524
rect 182 1519 183 1523
rect 187 1522 188 1523
rect 199 1523 205 1524
rect 199 1522 200 1523
rect 187 1520 200 1522
rect 187 1519 188 1520
rect 182 1518 188 1519
rect 199 1519 200 1520
rect 204 1519 205 1523
rect 199 1518 205 1519
rect 255 1523 261 1524
rect 255 1519 256 1523
rect 260 1519 261 1523
rect 255 1518 261 1519
rect 263 1523 269 1524
rect 263 1519 264 1523
rect 268 1522 269 1523
rect 335 1523 341 1524
rect 335 1522 336 1523
rect 268 1520 336 1522
rect 268 1519 269 1520
rect 263 1518 269 1519
rect 335 1519 336 1520
rect 340 1519 341 1523
rect 335 1518 341 1519
rect 343 1523 349 1524
rect 343 1519 344 1523
rect 348 1522 349 1523
rect 415 1523 421 1524
rect 415 1522 416 1523
rect 348 1520 416 1522
rect 348 1519 349 1520
rect 343 1518 349 1519
rect 415 1519 416 1520
rect 420 1519 421 1523
rect 415 1518 421 1519
rect 423 1523 429 1524
rect 423 1519 424 1523
rect 428 1522 429 1523
rect 503 1523 509 1524
rect 503 1522 504 1523
rect 428 1520 504 1522
rect 428 1519 429 1520
rect 423 1518 429 1519
rect 503 1519 504 1520
rect 508 1519 509 1523
rect 503 1518 509 1519
rect 590 1523 597 1524
rect 590 1519 591 1523
rect 596 1519 597 1523
rect 590 1518 597 1519
rect 599 1523 605 1524
rect 599 1519 600 1523
rect 604 1522 605 1523
rect 679 1523 685 1524
rect 679 1522 680 1523
rect 604 1520 680 1522
rect 604 1519 605 1520
rect 599 1518 605 1519
rect 679 1519 680 1520
rect 684 1519 685 1523
rect 679 1518 685 1519
rect 687 1523 693 1524
rect 687 1519 688 1523
rect 692 1522 693 1523
rect 767 1523 773 1524
rect 767 1522 768 1523
rect 692 1520 768 1522
rect 692 1519 693 1520
rect 687 1518 693 1519
rect 767 1519 768 1520
rect 772 1519 773 1523
rect 767 1518 773 1519
rect 847 1523 853 1524
rect 847 1519 848 1523
rect 852 1522 853 1523
rect 926 1523 932 1524
rect 926 1522 927 1523
rect 852 1520 927 1522
rect 852 1519 853 1520
rect 847 1518 853 1519
rect 926 1519 927 1520
rect 931 1519 932 1523
rect 926 1518 932 1519
rect 935 1523 941 1524
rect 935 1519 936 1523
rect 940 1522 941 1523
rect 962 1523 968 1524
rect 962 1522 963 1523
rect 940 1520 963 1522
rect 940 1519 941 1520
rect 935 1518 941 1519
rect 962 1519 963 1520
rect 967 1519 968 1523
rect 962 1518 968 1519
rect 970 1523 976 1524
rect 970 1519 971 1523
rect 975 1522 976 1523
rect 1023 1523 1029 1524
rect 1023 1522 1024 1523
rect 975 1520 1024 1522
rect 975 1519 976 1520
rect 970 1518 976 1519
rect 1023 1519 1024 1520
rect 1028 1519 1029 1523
rect 1023 1518 1029 1519
rect 1094 1520 1100 1521
rect 110 1515 116 1516
rect 1094 1516 1095 1520
rect 1099 1516 1100 1520
rect 1094 1515 1100 1516
rect 1134 1519 1140 1520
rect 1134 1515 1135 1519
rect 1139 1515 1140 1519
rect 2118 1519 2124 1520
rect 1134 1514 1140 1515
rect 1158 1516 1164 1517
rect 134 1512 140 1513
rect 134 1508 135 1512
rect 139 1508 140 1512
rect 134 1507 140 1508
rect 174 1512 180 1513
rect 174 1508 175 1512
rect 179 1508 180 1512
rect 174 1507 180 1508
rect 230 1512 236 1513
rect 230 1508 231 1512
rect 235 1508 236 1512
rect 230 1507 236 1508
rect 310 1512 316 1513
rect 310 1508 311 1512
rect 315 1508 316 1512
rect 310 1507 316 1508
rect 390 1512 396 1513
rect 390 1508 391 1512
rect 395 1508 396 1512
rect 390 1507 396 1508
rect 478 1512 484 1513
rect 478 1508 479 1512
rect 483 1508 484 1512
rect 478 1507 484 1508
rect 566 1512 572 1513
rect 566 1508 567 1512
rect 571 1508 572 1512
rect 566 1507 572 1508
rect 654 1512 660 1513
rect 654 1508 655 1512
rect 659 1508 660 1512
rect 654 1507 660 1508
rect 742 1512 748 1513
rect 742 1508 743 1512
rect 747 1508 748 1512
rect 742 1507 748 1508
rect 822 1512 828 1513
rect 822 1508 823 1512
rect 827 1508 828 1512
rect 822 1507 828 1508
rect 910 1512 916 1513
rect 910 1508 911 1512
rect 915 1508 916 1512
rect 910 1507 916 1508
rect 998 1512 1004 1513
rect 998 1508 999 1512
rect 1003 1508 1004 1512
rect 1158 1512 1159 1516
rect 1163 1512 1164 1516
rect 1158 1511 1164 1512
rect 1198 1516 1204 1517
rect 1198 1512 1199 1516
rect 1203 1512 1204 1516
rect 1198 1511 1204 1512
rect 1246 1516 1252 1517
rect 1246 1512 1247 1516
rect 1251 1512 1252 1516
rect 1246 1511 1252 1512
rect 1318 1516 1324 1517
rect 1318 1512 1319 1516
rect 1323 1512 1324 1516
rect 1318 1511 1324 1512
rect 1398 1516 1404 1517
rect 1398 1512 1399 1516
rect 1403 1512 1404 1516
rect 1398 1511 1404 1512
rect 1478 1516 1484 1517
rect 1478 1512 1479 1516
rect 1483 1512 1484 1516
rect 1478 1511 1484 1512
rect 1558 1516 1564 1517
rect 1558 1512 1559 1516
rect 1563 1512 1564 1516
rect 1558 1511 1564 1512
rect 1646 1516 1652 1517
rect 1646 1512 1647 1516
rect 1651 1512 1652 1516
rect 1646 1511 1652 1512
rect 1734 1516 1740 1517
rect 1734 1512 1735 1516
rect 1739 1512 1740 1516
rect 1734 1511 1740 1512
rect 1822 1516 1828 1517
rect 1822 1512 1823 1516
rect 1827 1512 1828 1516
rect 1822 1511 1828 1512
rect 1910 1516 1916 1517
rect 1910 1512 1911 1516
rect 1915 1512 1916 1516
rect 1910 1511 1916 1512
rect 1998 1516 2004 1517
rect 1998 1512 1999 1516
rect 2003 1512 2004 1516
rect 1998 1511 2004 1512
rect 2070 1516 2076 1517
rect 2070 1512 2071 1516
rect 2075 1512 2076 1516
rect 2118 1515 2119 1519
rect 2123 1515 2124 1519
rect 2118 1514 2124 1515
rect 2070 1511 2076 1512
rect 998 1507 1004 1508
rect 1158 1504 1164 1505
rect 159 1503 165 1504
rect 159 1499 160 1503
rect 164 1502 165 1503
rect 182 1503 188 1504
rect 182 1502 183 1503
rect 164 1500 183 1502
rect 164 1499 165 1500
rect 159 1498 165 1499
rect 182 1499 183 1500
rect 187 1499 188 1503
rect 182 1498 188 1499
rect 199 1503 205 1504
rect 199 1499 200 1503
rect 204 1502 205 1503
rect 215 1503 221 1504
rect 215 1502 216 1503
rect 204 1500 216 1502
rect 204 1499 205 1500
rect 199 1498 205 1499
rect 215 1499 216 1500
rect 220 1499 221 1503
rect 215 1498 221 1499
rect 255 1503 261 1504
rect 255 1499 256 1503
rect 260 1502 261 1503
rect 263 1503 269 1504
rect 263 1502 264 1503
rect 260 1500 264 1502
rect 260 1499 261 1500
rect 255 1498 261 1499
rect 263 1499 264 1500
rect 268 1499 269 1503
rect 263 1498 269 1499
rect 335 1503 341 1504
rect 335 1499 336 1503
rect 340 1502 341 1503
rect 343 1503 349 1504
rect 343 1502 344 1503
rect 340 1500 344 1502
rect 340 1499 341 1500
rect 335 1498 341 1499
rect 343 1499 344 1500
rect 348 1499 349 1503
rect 343 1498 349 1499
rect 415 1503 421 1504
rect 415 1499 416 1503
rect 420 1502 421 1503
rect 423 1503 429 1504
rect 423 1502 424 1503
rect 420 1500 424 1502
rect 420 1499 421 1500
rect 415 1498 421 1499
rect 423 1499 424 1500
rect 428 1499 429 1503
rect 423 1498 429 1499
rect 434 1503 440 1504
rect 434 1499 435 1503
rect 439 1502 440 1503
rect 503 1503 509 1504
rect 503 1502 504 1503
rect 439 1500 504 1502
rect 439 1499 440 1500
rect 434 1498 440 1499
rect 503 1499 504 1500
rect 508 1499 509 1503
rect 503 1498 509 1499
rect 591 1503 597 1504
rect 591 1499 592 1503
rect 596 1502 597 1503
rect 599 1503 605 1504
rect 599 1502 600 1503
rect 596 1500 600 1502
rect 596 1499 597 1500
rect 591 1498 597 1499
rect 599 1499 600 1500
rect 604 1499 605 1503
rect 599 1498 605 1499
rect 679 1503 685 1504
rect 679 1499 680 1503
rect 684 1502 685 1503
rect 687 1503 693 1504
rect 687 1502 688 1503
rect 684 1500 688 1502
rect 684 1499 685 1500
rect 679 1498 685 1499
rect 687 1499 688 1500
rect 692 1499 693 1503
rect 687 1498 693 1499
rect 706 1503 712 1504
rect 706 1499 707 1503
rect 711 1502 712 1503
rect 767 1503 773 1504
rect 767 1502 768 1503
rect 711 1500 768 1502
rect 711 1499 712 1500
rect 706 1498 712 1499
rect 767 1499 768 1500
rect 772 1499 773 1503
rect 767 1498 773 1499
rect 847 1503 856 1504
rect 847 1499 848 1503
rect 855 1499 856 1503
rect 847 1498 856 1499
rect 926 1503 932 1504
rect 926 1499 927 1503
rect 931 1502 932 1503
rect 935 1503 941 1504
rect 935 1502 936 1503
rect 931 1500 936 1502
rect 931 1499 932 1500
rect 926 1498 932 1499
rect 935 1499 936 1500
rect 940 1499 941 1503
rect 935 1498 941 1499
rect 962 1503 968 1504
rect 962 1499 963 1503
rect 967 1502 968 1503
rect 1023 1503 1029 1504
rect 1023 1502 1024 1503
rect 967 1500 1024 1502
rect 967 1499 968 1500
rect 962 1498 968 1499
rect 1023 1499 1024 1500
rect 1028 1499 1029 1503
rect 1023 1498 1029 1499
rect 1134 1501 1140 1502
rect 1134 1497 1135 1501
rect 1139 1497 1140 1501
rect 1158 1500 1159 1504
rect 1163 1500 1164 1504
rect 1158 1499 1164 1500
rect 1198 1504 1204 1505
rect 1198 1500 1199 1504
rect 1203 1500 1204 1504
rect 1198 1499 1204 1500
rect 1238 1504 1244 1505
rect 1238 1500 1239 1504
rect 1243 1500 1244 1504
rect 1238 1499 1244 1500
rect 1302 1504 1308 1505
rect 1302 1500 1303 1504
rect 1307 1500 1308 1504
rect 1302 1499 1308 1500
rect 1374 1504 1380 1505
rect 1374 1500 1375 1504
rect 1379 1500 1380 1504
rect 1374 1499 1380 1500
rect 1454 1504 1460 1505
rect 1454 1500 1455 1504
rect 1459 1500 1460 1504
rect 1454 1499 1460 1500
rect 1542 1504 1548 1505
rect 1542 1500 1543 1504
rect 1547 1500 1548 1504
rect 1542 1499 1548 1500
rect 1622 1504 1628 1505
rect 1622 1500 1623 1504
rect 1627 1500 1628 1504
rect 1622 1499 1628 1500
rect 1702 1504 1708 1505
rect 1702 1500 1703 1504
rect 1707 1500 1708 1504
rect 1702 1499 1708 1500
rect 1774 1504 1780 1505
rect 1774 1500 1775 1504
rect 1779 1500 1780 1504
rect 1774 1499 1780 1500
rect 1846 1504 1852 1505
rect 1846 1500 1847 1504
rect 1851 1500 1852 1504
rect 1846 1499 1852 1500
rect 1918 1504 1924 1505
rect 1918 1500 1919 1504
rect 1923 1500 1924 1504
rect 1918 1499 1924 1500
rect 1990 1504 1996 1505
rect 1990 1500 1991 1504
rect 1995 1500 1996 1504
rect 1990 1499 1996 1500
rect 2062 1504 2068 1505
rect 2062 1500 2063 1504
rect 2067 1500 2068 1504
rect 2062 1499 2068 1500
rect 2118 1501 2124 1502
rect 1134 1496 1140 1497
rect 2118 1497 2119 1501
rect 2123 1497 2124 1501
rect 2118 1496 2124 1497
rect 1798 1495 1804 1496
rect 1798 1494 1799 1495
rect 1648 1492 1799 1494
rect 162 1491 168 1492
rect 162 1487 163 1491
rect 167 1490 168 1491
rect 167 1488 226 1490
rect 1648 1488 1650 1492
rect 1798 1491 1799 1492
rect 1803 1491 1804 1495
rect 1798 1490 1804 1491
rect 167 1487 168 1488
rect 162 1486 168 1487
rect 224 1484 226 1488
rect 1183 1487 1189 1488
rect 1134 1484 1140 1485
rect 159 1483 165 1484
rect 159 1479 160 1483
rect 164 1482 165 1483
rect 214 1483 220 1484
rect 214 1482 215 1483
rect 164 1480 215 1482
rect 164 1479 165 1480
rect 159 1478 165 1479
rect 214 1479 215 1480
rect 219 1479 220 1483
rect 214 1478 220 1479
rect 223 1483 229 1484
rect 223 1479 224 1483
rect 228 1479 229 1483
rect 223 1478 229 1479
rect 290 1483 296 1484
rect 290 1479 291 1483
rect 295 1482 296 1483
rect 303 1483 309 1484
rect 303 1482 304 1483
rect 295 1480 304 1482
rect 295 1479 296 1480
rect 290 1478 296 1479
rect 303 1479 304 1480
rect 308 1479 309 1483
rect 303 1478 309 1479
rect 311 1483 317 1484
rect 311 1479 312 1483
rect 316 1482 317 1483
rect 383 1483 389 1484
rect 383 1482 384 1483
rect 316 1480 384 1482
rect 316 1479 317 1480
rect 311 1478 317 1479
rect 383 1479 384 1480
rect 388 1479 389 1483
rect 383 1478 389 1479
rect 463 1483 469 1484
rect 463 1479 464 1483
rect 468 1482 469 1483
rect 534 1483 540 1484
rect 534 1482 535 1483
rect 468 1480 535 1482
rect 468 1479 469 1480
rect 463 1478 469 1479
rect 534 1479 535 1480
rect 539 1479 540 1483
rect 534 1478 540 1479
rect 543 1483 549 1484
rect 543 1479 544 1483
rect 548 1482 549 1483
rect 614 1483 620 1484
rect 614 1482 615 1483
rect 548 1480 615 1482
rect 548 1479 549 1480
rect 543 1478 549 1479
rect 614 1479 615 1480
rect 619 1479 620 1483
rect 614 1478 620 1479
rect 623 1483 629 1484
rect 623 1479 624 1483
rect 628 1482 629 1483
rect 654 1483 660 1484
rect 654 1482 655 1483
rect 628 1480 655 1482
rect 628 1479 629 1480
rect 623 1478 629 1479
rect 654 1479 655 1480
rect 659 1479 660 1483
rect 654 1478 660 1479
rect 703 1483 709 1484
rect 703 1479 704 1483
rect 708 1482 709 1483
rect 782 1483 788 1484
rect 782 1482 783 1483
rect 708 1480 783 1482
rect 708 1479 709 1480
rect 703 1478 709 1479
rect 782 1479 783 1480
rect 787 1479 788 1483
rect 782 1478 788 1479
rect 791 1483 797 1484
rect 791 1479 792 1483
rect 796 1482 797 1483
rect 818 1483 824 1484
rect 818 1482 819 1483
rect 796 1480 819 1482
rect 796 1479 797 1480
rect 791 1478 797 1479
rect 818 1479 819 1480
rect 823 1479 824 1483
rect 818 1478 824 1479
rect 826 1483 832 1484
rect 826 1479 827 1483
rect 831 1482 832 1483
rect 879 1483 885 1484
rect 879 1482 880 1483
rect 831 1480 880 1482
rect 831 1479 832 1480
rect 826 1478 832 1479
rect 879 1479 880 1480
rect 884 1479 885 1483
rect 879 1478 885 1479
rect 967 1483 976 1484
rect 967 1479 968 1483
rect 975 1479 976 1483
rect 967 1478 976 1479
rect 978 1483 984 1484
rect 978 1479 979 1483
rect 983 1482 984 1483
rect 1055 1483 1061 1484
rect 1055 1482 1056 1483
rect 983 1480 1056 1482
rect 983 1479 984 1480
rect 978 1478 984 1479
rect 1055 1479 1056 1480
rect 1060 1479 1061 1483
rect 1134 1480 1135 1484
rect 1139 1480 1140 1484
rect 1183 1483 1184 1487
rect 1188 1486 1189 1487
rect 1214 1487 1220 1488
rect 1214 1486 1215 1487
rect 1188 1484 1215 1486
rect 1188 1483 1189 1484
rect 1183 1482 1189 1483
rect 1214 1483 1215 1484
rect 1219 1483 1220 1487
rect 1214 1482 1220 1483
rect 1223 1487 1229 1488
rect 1223 1483 1224 1487
rect 1228 1486 1229 1487
rect 1254 1487 1260 1488
rect 1254 1486 1255 1487
rect 1228 1484 1255 1486
rect 1228 1483 1229 1484
rect 1223 1482 1229 1483
rect 1254 1483 1255 1484
rect 1259 1483 1260 1487
rect 1254 1482 1260 1483
rect 1263 1487 1269 1488
rect 1263 1483 1264 1487
rect 1268 1486 1269 1487
rect 1318 1487 1324 1488
rect 1318 1486 1319 1487
rect 1268 1484 1319 1486
rect 1268 1483 1269 1484
rect 1263 1482 1269 1483
rect 1318 1483 1319 1484
rect 1323 1483 1324 1487
rect 1318 1482 1324 1483
rect 1327 1487 1333 1488
rect 1327 1483 1328 1487
rect 1332 1486 1333 1487
rect 1390 1487 1396 1488
rect 1390 1486 1391 1487
rect 1332 1484 1391 1486
rect 1332 1483 1333 1484
rect 1327 1482 1333 1483
rect 1390 1483 1391 1484
rect 1395 1483 1396 1487
rect 1390 1482 1396 1483
rect 1399 1487 1405 1488
rect 1399 1483 1400 1487
rect 1404 1486 1405 1487
rect 1470 1487 1476 1488
rect 1470 1486 1471 1487
rect 1404 1484 1471 1486
rect 1404 1483 1405 1484
rect 1399 1482 1405 1483
rect 1470 1483 1471 1484
rect 1475 1483 1476 1487
rect 1470 1482 1476 1483
rect 1479 1487 1485 1488
rect 1479 1483 1480 1487
rect 1484 1486 1485 1487
rect 1519 1487 1525 1488
rect 1519 1486 1520 1487
rect 1484 1484 1520 1486
rect 1484 1483 1485 1484
rect 1479 1482 1485 1483
rect 1519 1483 1520 1484
rect 1524 1483 1525 1487
rect 1519 1482 1525 1483
rect 1534 1487 1540 1488
rect 1534 1483 1535 1487
rect 1539 1486 1540 1487
rect 1567 1487 1573 1488
rect 1567 1486 1568 1487
rect 1539 1484 1568 1486
rect 1539 1483 1540 1484
rect 1534 1482 1540 1483
rect 1567 1483 1568 1484
rect 1572 1483 1573 1487
rect 1567 1482 1573 1483
rect 1647 1487 1653 1488
rect 1647 1483 1648 1487
rect 1652 1483 1653 1487
rect 1647 1482 1653 1483
rect 1655 1487 1661 1488
rect 1655 1483 1656 1487
rect 1660 1486 1661 1487
rect 1727 1487 1733 1488
rect 1727 1486 1728 1487
rect 1660 1484 1728 1486
rect 1660 1483 1661 1484
rect 1655 1482 1661 1483
rect 1727 1483 1728 1484
rect 1732 1483 1733 1487
rect 1727 1482 1733 1483
rect 1735 1487 1741 1488
rect 1735 1483 1736 1487
rect 1740 1486 1741 1487
rect 1799 1487 1805 1488
rect 1799 1486 1800 1487
rect 1740 1484 1800 1486
rect 1740 1483 1741 1484
rect 1735 1482 1741 1483
rect 1799 1483 1800 1484
rect 1804 1483 1805 1487
rect 1799 1482 1805 1483
rect 1807 1487 1813 1488
rect 1807 1483 1808 1487
rect 1812 1486 1813 1487
rect 1871 1487 1877 1488
rect 1871 1486 1872 1487
rect 1812 1484 1872 1486
rect 1812 1483 1813 1484
rect 1807 1482 1813 1483
rect 1871 1483 1872 1484
rect 1876 1483 1877 1487
rect 1871 1482 1877 1483
rect 1943 1487 1952 1488
rect 1943 1483 1944 1487
rect 1951 1483 1952 1487
rect 1943 1482 1952 1483
rect 2015 1487 2021 1488
rect 2015 1483 2016 1487
rect 2020 1486 2021 1487
rect 2078 1487 2084 1488
rect 2078 1486 2079 1487
rect 2020 1484 2079 1486
rect 2020 1483 2021 1484
rect 2015 1482 2021 1483
rect 2078 1483 2079 1484
rect 2083 1483 2084 1487
rect 2078 1482 2084 1483
rect 2086 1487 2093 1488
rect 2086 1483 2087 1487
rect 2092 1483 2093 1487
rect 2086 1482 2093 1483
rect 2118 1484 2124 1485
rect 1134 1479 1140 1480
rect 2118 1480 2119 1484
rect 2123 1480 2124 1484
rect 2118 1479 2124 1480
rect 1055 1478 1061 1479
rect 134 1476 140 1477
rect 134 1472 135 1476
rect 139 1472 140 1476
rect 134 1471 140 1472
rect 198 1476 204 1477
rect 198 1472 199 1476
rect 203 1472 204 1476
rect 198 1471 204 1472
rect 278 1476 284 1477
rect 278 1472 279 1476
rect 283 1472 284 1476
rect 278 1471 284 1472
rect 358 1476 364 1477
rect 358 1472 359 1476
rect 363 1472 364 1476
rect 358 1471 364 1472
rect 438 1476 444 1477
rect 438 1472 439 1476
rect 443 1472 444 1476
rect 438 1471 444 1472
rect 518 1476 524 1477
rect 518 1472 519 1476
rect 523 1472 524 1476
rect 518 1471 524 1472
rect 598 1476 604 1477
rect 598 1472 599 1476
rect 603 1472 604 1476
rect 598 1471 604 1472
rect 678 1476 684 1477
rect 678 1472 679 1476
rect 683 1472 684 1476
rect 678 1471 684 1472
rect 766 1476 772 1477
rect 766 1472 767 1476
rect 771 1472 772 1476
rect 766 1471 772 1472
rect 854 1476 860 1477
rect 854 1472 855 1476
rect 859 1472 860 1476
rect 854 1471 860 1472
rect 942 1476 948 1477
rect 942 1472 943 1476
rect 947 1472 948 1476
rect 942 1471 948 1472
rect 1030 1476 1036 1477
rect 1030 1472 1031 1476
rect 1035 1472 1036 1476
rect 1030 1471 1036 1472
rect 1158 1476 1164 1477
rect 1158 1472 1159 1476
rect 1163 1472 1164 1476
rect 1158 1471 1164 1472
rect 1198 1476 1204 1477
rect 1198 1472 1199 1476
rect 1203 1472 1204 1476
rect 1198 1471 1204 1472
rect 1238 1476 1244 1477
rect 1238 1472 1239 1476
rect 1243 1472 1244 1476
rect 1238 1471 1244 1472
rect 1302 1476 1308 1477
rect 1302 1472 1303 1476
rect 1307 1472 1308 1476
rect 1302 1471 1308 1472
rect 1374 1476 1380 1477
rect 1374 1472 1375 1476
rect 1379 1472 1380 1476
rect 1374 1471 1380 1472
rect 1454 1476 1460 1477
rect 1454 1472 1455 1476
rect 1459 1472 1460 1476
rect 1454 1471 1460 1472
rect 1542 1476 1548 1477
rect 1542 1472 1543 1476
rect 1547 1472 1548 1476
rect 1542 1471 1548 1472
rect 1622 1476 1628 1477
rect 1622 1472 1623 1476
rect 1627 1472 1628 1476
rect 1622 1471 1628 1472
rect 1702 1476 1708 1477
rect 1702 1472 1703 1476
rect 1707 1472 1708 1476
rect 1702 1471 1708 1472
rect 1774 1476 1780 1477
rect 1774 1472 1775 1476
rect 1779 1472 1780 1476
rect 1774 1471 1780 1472
rect 1846 1476 1852 1477
rect 1846 1472 1847 1476
rect 1851 1472 1852 1476
rect 1846 1471 1852 1472
rect 1918 1476 1924 1477
rect 1918 1472 1919 1476
rect 1923 1472 1924 1476
rect 1918 1471 1924 1472
rect 1990 1476 1996 1477
rect 2062 1476 2068 1477
rect 1990 1472 1991 1476
rect 1995 1472 1996 1476
rect 2038 1475 2044 1476
rect 2038 1474 2039 1475
rect 1990 1471 1996 1472
rect 1999 1472 2039 1474
rect 110 1468 116 1469
rect 110 1464 111 1468
rect 115 1464 116 1468
rect 1094 1468 1100 1469
rect 1094 1464 1095 1468
rect 1099 1464 1100 1468
rect 110 1463 116 1464
rect 158 1463 165 1464
rect 158 1459 159 1463
rect 164 1459 165 1463
rect 158 1458 165 1459
rect 214 1463 220 1464
rect 214 1459 215 1463
rect 219 1462 220 1463
rect 223 1463 229 1464
rect 223 1462 224 1463
rect 219 1460 224 1462
rect 219 1459 220 1460
rect 214 1458 220 1459
rect 223 1459 224 1460
rect 228 1459 229 1463
rect 223 1458 229 1459
rect 303 1463 309 1464
rect 303 1459 304 1463
rect 308 1462 309 1463
rect 311 1463 317 1464
rect 311 1462 312 1463
rect 308 1460 312 1462
rect 308 1459 309 1460
rect 303 1458 309 1459
rect 311 1459 312 1460
rect 316 1459 317 1463
rect 311 1458 317 1459
rect 383 1463 389 1464
rect 383 1459 384 1463
rect 388 1462 389 1463
rect 430 1463 436 1464
rect 430 1462 431 1463
rect 388 1460 431 1462
rect 388 1459 389 1460
rect 383 1458 389 1459
rect 430 1459 431 1460
rect 435 1459 436 1463
rect 430 1458 436 1459
rect 446 1463 452 1464
rect 446 1459 447 1463
rect 451 1462 452 1463
rect 463 1463 469 1464
rect 463 1462 464 1463
rect 451 1460 464 1462
rect 451 1459 452 1460
rect 446 1458 452 1459
rect 463 1459 464 1460
rect 468 1459 469 1463
rect 463 1458 469 1459
rect 534 1463 540 1464
rect 534 1459 535 1463
rect 539 1462 540 1463
rect 543 1463 549 1464
rect 543 1462 544 1463
rect 539 1460 544 1462
rect 539 1459 540 1460
rect 534 1458 540 1459
rect 543 1459 544 1460
rect 548 1459 549 1463
rect 543 1458 549 1459
rect 614 1463 620 1464
rect 614 1459 615 1463
rect 619 1462 620 1463
rect 623 1463 629 1464
rect 623 1462 624 1463
rect 619 1460 624 1462
rect 619 1459 620 1460
rect 614 1458 620 1459
rect 623 1459 624 1460
rect 628 1459 629 1463
rect 623 1458 629 1459
rect 703 1463 712 1464
rect 703 1459 704 1463
rect 711 1459 712 1463
rect 703 1458 712 1459
rect 782 1463 788 1464
rect 782 1459 783 1463
rect 787 1462 788 1463
rect 791 1463 797 1464
rect 791 1462 792 1463
rect 787 1460 792 1462
rect 787 1459 788 1460
rect 782 1458 788 1459
rect 791 1459 792 1460
rect 796 1459 797 1463
rect 791 1458 797 1459
rect 818 1463 824 1464
rect 818 1459 819 1463
rect 823 1462 824 1463
rect 879 1463 885 1464
rect 879 1462 880 1463
rect 823 1460 880 1462
rect 823 1459 824 1460
rect 818 1458 824 1459
rect 879 1459 880 1460
rect 884 1459 885 1463
rect 879 1458 885 1459
rect 967 1463 973 1464
rect 967 1459 968 1463
rect 972 1462 973 1463
rect 978 1463 984 1464
rect 978 1462 979 1463
rect 972 1460 979 1462
rect 972 1459 973 1460
rect 967 1458 973 1459
rect 978 1459 979 1460
rect 983 1459 984 1463
rect 978 1458 984 1459
rect 1055 1463 1061 1464
rect 1055 1459 1056 1463
rect 1060 1462 1061 1463
rect 1070 1463 1076 1464
rect 1094 1463 1100 1464
rect 1182 1467 1189 1468
rect 1182 1463 1183 1467
rect 1188 1463 1189 1467
rect 1070 1462 1071 1463
rect 1060 1460 1071 1462
rect 1060 1459 1061 1460
rect 1055 1458 1061 1459
rect 1070 1459 1071 1460
rect 1075 1459 1076 1463
rect 1182 1462 1189 1463
rect 1214 1467 1220 1468
rect 1214 1463 1215 1467
rect 1219 1466 1220 1467
rect 1223 1467 1229 1468
rect 1223 1466 1224 1467
rect 1219 1464 1224 1466
rect 1219 1463 1220 1464
rect 1214 1462 1220 1463
rect 1223 1463 1224 1464
rect 1228 1463 1229 1467
rect 1223 1462 1229 1463
rect 1254 1467 1260 1468
rect 1254 1463 1255 1467
rect 1259 1466 1260 1467
rect 1263 1467 1269 1468
rect 1263 1466 1264 1467
rect 1259 1464 1264 1466
rect 1259 1463 1260 1464
rect 1254 1462 1260 1463
rect 1263 1463 1264 1464
rect 1268 1463 1269 1467
rect 1263 1462 1269 1463
rect 1318 1467 1324 1468
rect 1318 1463 1319 1467
rect 1323 1466 1324 1467
rect 1327 1467 1333 1468
rect 1327 1466 1328 1467
rect 1323 1464 1328 1466
rect 1323 1463 1324 1464
rect 1318 1462 1324 1463
rect 1327 1463 1328 1464
rect 1332 1463 1333 1467
rect 1327 1462 1333 1463
rect 1390 1467 1396 1468
rect 1390 1463 1391 1467
rect 1395 1466 1396 1467
rect 1399 1467 1405 1468
rect 1399 1466 1400 1467
rect 1395 1464 1400 1466
rect 1395 1463 1396 1464
rect 1390 1462 1396 1463
rect 1399 1463 1400 1464
rect 1404 1463 1405 1467
rect 1399 1462 1405 1463
rect 1470 1467 1476 1468
rect 1470 1463 1471 1467
rect 1475 1466 1476 1467
rect 1479 1467 1485 1468
rect 1479 1466 1480 1467
rect 1475 1464 1480 1466
rect 1475 1463 1476 1464
rect 1470 1462 1476 1463
rect 1479 1463 1480 1464
rect 1484 1463 1485 1467
rect 1479 1462 1485 1463
rect 1519 1467 1525 1468
rect 1519 1463 1520 1467
rect 1524 1466 1525 1467
rect 1567 1467 1573 1468
rect 1567 1466 1568 1467
rect 1524 1464 1568 1466
rect 1524 1463 1525 1464
rect 1519 1462 1525 1463
rect 1567 1463 1568 1464
rect 1572 1463 1573 1467
rect 1567 1462 1573 1463
rect 1647 1467 1653 1468
rect 1647 1463 1648 1467
rect 1652 1466 1653 1467
rect 1655 1467 1661 1468
rect 1655 1466 1656 1467
rect 1652 1464 1656 1466
rect 1652 1463 1653 1464
rect 1647 1462 1653 1463
rect 1655 1463 1656 1464
rect 1660 1463 1661 1467
rect 1655 1462 1661 1463
rect 1727 1467 1733 1468
rect 1727 1463 1728 1467
rect 1732 1466 1733 1467
rect 1735 1467 1741 1468
rect 1735 1466 1736 1467
rect 1732 1464 1736 1466
rect 1732 1463 1733 1464
rect 1727 1462 1733 1463
rect 1735 1463 1736 1464
rect 1740 1463 1741 1467
rect 1735 1462 1741 1463
rect 1799 1467 1805 1468
rect 1799 1463 1800 1467
rect 1804 1466 1805 1467
rect 1807 1467 1813 1468
rect 1807 1466 1808 1467
rect 1804 1464 1808 1466
rect 1804 1463 1805 1464
rect 1799 1462 1805 1463
rect 1807 1463 1808 1464
rect 1812 1463 1813 1467
rect 1807 1462 1813 1463
rect 1871 1467 1877 1468
rect 1871 1463 1872 1467
rect 1876 1466 1877 1467
rect 1910 1467 1916 1468
rect 1910 1466 1911 1467
rect 1876 1464 1911 1466
rect 1876 1463 1877 1464
rect 1871 1462 1877 1463
rect 1910 1463 1911 1464
rect 1915 1463 1916 1467
rect 1910 1462 1916 1463
rect 1943 1467 1949 1468
rect 1943 1463 1944 1467
rect 1948 1466 1949 1467
rect 1999 1466 2001 1472
rect 2038 1471 2039 1472
rect 2043 1471 2044 1475
rect 2062 1472 2063 1476
rect 2067 1472 2068 1476
rect 2062 1471 2068 1472
rect 2038 1470 2044 1471
rect 1948 1464 2001 1466
rect 2015 1467 2024 1468
rect 1948 1463 1949 1464
rect 1943 1462 1949 1463
rect 2015 1463 2016 1467
rect 2023 1463 2024 1467
rect 2015 1462 2024 1463
rect 2078 1467 2084 1468
rect 2078 1463 2079 1467
rect 2083 1466 2084 1467
rect 2087 1467 2093 1468
rect 2087 1466 2088 1467
rect 2083 1464 2088 1466
rect 2083 1463 2084 1464
rect 2078 1462 2084 1463
rect 2087 1463 2088 1464
rect 2092 1463 2093 1467
rect 2087 1462 2093 1463
rect 1070 1458 1076 1459
rect 110 1451 116 1452
rect 110 1447 111 1451
rect 115 1447 116 1451
rect 1094 1451 1100 1452
rect 110 1446 116 1447
rect 134 1448 140 1449
rect 134 1444 135 1448
rect 139 1444 140 1448
rect 134 1443 140 1444
rect 198 1448 204 1449
rect 198 1444 199 1448
rect 203 1444 204 1448
rect 198 1443 204 1444
rect 278 1448 284 1449
rect 278 1444 279 1448
rect 283 1444 284 1448
rect 278 1443 284 1444
rect 358 1448 364 1449
rect 358 1444 359 1448
rect 363 1444 364 1448
rect 358 1443 364 1444
rect 438 1448 444 1449
rect 438 1444 439 1448
rect 443 1444 444 1448
rect 438 1443 444 1444
rect 518 1448 524 1449
rect 518 1444 519 1448
rect 523 1444 524 1448
rect 518 1443 524 1444
rect 598 1448 604 1449
rect 598 1444 599 1448
rect 603 1444 604 1448
rect 598 1443 604 1444
rect 678 1448 684 1449
rect 678 1444 679 1448
rect 683 1444 684 1448
rect 678 1443 684 1444
rect 766 1448 772 1449
rect 766 1444 767 1448
rect 771 1444 772 1448
rect 766 1443 772 1444
rect 854 1448 860 1449
rect 854 1444 855 1448
rect 859 1444 860 1448
rect 854 1443 860 1444
rect 942 1448 948 1449
rect 942 1444 943 1448
rect 947 1444 948 1448
rect 942 1443 948 1444
rect 1030 1448 1036 1449
rect 1030 1444 1031 1448
rect 1035 1444 1036 1448
rect 1094 1447 1095 1451
rect 1099 1447 1100 1451
rect 1094 1446 1100 1447
rect 1578 1451 1584 1452
rect 1578 1447 1579 1451
rect 1583 1450 1584 1451
rect 1583 1448 1754 1450
rect 1583 1447 1584 1448
rect 1578 1446 1584 1447
rect 1030 1443 1036 1444
rect 1303 1443 1309 1444
rect 1303 1439 1304 1443
rect 1308 1442 1309 1443
rect 1342 1443 1348 1444
rect 1342 1442 1343 1443
rect 1308 1440 1343 1442
rect 1308 1439 1309 1440
rect 1303 1438 1309 1439
rect 1342 1439 1343 1440
rect 1347 1439 1348 1443
rect 1342 1438 1348 1439
rect 1351 1443 1357 1444
rect 1351 1439 1352 1443
rect 1356 1442 1357 1443
rect 1398 1443 1404 1444
rect 1398 1442 1399 1443
rect 1356 1440 1399 1442
rect 1356 1439 1357 1440
rect 1351 1438 1357 1439
rect 1398 1439 1399 1440
rect 1403 1439 1404 1443
rect 1398 1438 1404 1439
rect 1407 1443 1413 1444
rect 1407 1439 1408 1443
rect 1412 1442 1413 1443
rect 1446 1443 1452 1444
rect 1446 1442 1447 1443
rect 1412 1440 1447 1442
rect 1412 1439 1413 1440
rect 1407 1438 1413 1439
rect 1446 1439 1447 1440
rect 1451 1439 1452 1443
rect 1446 1438 1452 1439
rect 1463 1443 1469 1444
rect 1463 1439 1464 1443
rect 1468 1442 1469 1443
rect 1510 1443 1516 1444
rect 1510 1442 1511 1443
rect 1468 1440 1511 1442
rect 1468 1439 1469 1440
rect 1463 1438 1469 1439
rect 1510 1439 1511 1440
rect 1515 1439 1516 1443
rect 1510 1438 1516 1439
rect 1519 1443 1525 1444
rect 1519 1439 1520 1443
rect 1524 1442 1525 1443
rect 1534 1443 1540 1444
rect 1534 1442 1535 1443
rect 1524 1440 1535 1442
rect 1524 1439 1525 1440
rect 1519 1438 1525 1439
rect 1534 1439 1535 1440
rect 1539 1439 1540 1443
rect 1534 1438 1540 1439
rect 1575 1443 1581 1444
rect 1575 1439 1576 1443
rect 1580 1442 1581 1443
rect 1614 1443 1620 1444
rect 1614 1442 1615 1443
rect 1580 1440 1615 1442
rect 1580 1439 1581 1440
rect 1575 1438 1581 1439
rect 1614 1439 1615 1440
rect 1619 1439 1620 1443
rect 1614 1438 1620 1439
rect 1631 1443 1637 1444
rect 1631 1439 1632 1443
rect 1636 1442 1637 1443
rect 1686 1443 1692 1444
rect 1686 1442 1687 1443
rect 1636 1440 1687 1442
rect 1636 1439 1637 1440
rect 1631 1438 1637 1439
rect 1686 1439 1687 1440
rect 1691 1439 1692 1443
rect 1686 1438 1692 1439
rect 1695 1443 1701 1444
rect 1695 1439 1696 1443
rect 1700 1442 1701 1443
rect 1742 1443 1748 1444
rect 1742 1442 1743 1443
rect 1700 1440 1743 1442
rect 1700 1439 1701 1440
rect 1695 1438 1701 1439
rect 1742 1439 1743 1440
rect 1747 1439 1748 1443
rect 1752 1442 1754 1448
rect 1759 1443 1765 1444
rect 1759 1442 1760 1443
rect 1752 1440 1760 1442
rect 1742 1438 1748 1439
rect 1759 1439 1760 1440
rect 1764 1439 1765 1443
rect 1759 1438 1765 1439
rect 1767 1443 1773 1444
rect 1767 1439 1768 1443
rect 1772 1442 1773 1443
rect 1831 1443 1837 1444
rect 1831 1442 1832 1443
rect 1772 1440 1832 1442
rect 1772 1439 1773 1440
rect 1767 1438 1773 1439
rect 1831 1439 1832 1440
rect 1836 1439 1837 1443
rect 1831 1438 1837 1439
rect 1839 1443 1845 1444
rect 1839 1439 1840 1443
rect 1844 1442 1845 1443
rect 1911 1443 1917 1444
rect 1911 1442 1912 1443
rect 1844 1440 1912 1442
rect 1844 1439 1845 1440
rect 1839 1438 1845 1439
rect 1911 1439 1912 1440
rect 1916 1439 1917 1443
rect 1911 1438 1917 1439
rect 1999 1443 2005 1444
rect 1999 1439 2000 1443
rect 2004 1442 2005 1443
rect 2078 1443 2084 1444
rect 2078 1442 2079 1443
rect 2004 1440 2079 1442
rect 2004 1439 2005 1440
rect 1999 1438 2005 1439
rect 2078 1439 2079 1440
rect 2083 1439 2084 1443
rect 2078 1438 2084 1439
rect 2086 1443 2093 1444
rect 2086 1439 2087 1443
rect 2092 1439 2093 1443
rect 2086 1438 2093 1439
rect 134 1436 140 1437
rect 110 1433 116 1434
rect 110 1429 111 1433
rect 115 1429 116 1433
rect 134 1432 135 1436
rect 139 1432 140 1436
rect 134 1431 140 1432
rect 190 1436 196 1437
rect 190 1432 191 1436
rect 195 1432 196 1436
rect 190 1431 196 1432
rect 262 1436 268 1437
rect 262 1432 263 1436
rect 267 1432 268 1436
rect 262 1431 268 1432
rect 334 1436 340 1437
rect 334 1432 335 1436
rect 339 1432 340 1436
rect 334 1431 340 1432
rect 406 1436 412 1437
rect 406 1432 407 1436
rect 411 1432 412 1436
rect 406 1431 412 1432
rect 478 1436 484 1437
rect 478 1432 479 1436
rect 483 1432 484 1436
rect 478 1431 484 1432
rect 550 1436 556 1437
rect 550 1432 551 1436
rect 555 1432 556 1436
rect 550 1431 556 1432
rect 630 1436 636 1437
rect 630 1432 631 1436
rect 635 1432 636 1436
rect 630 1431 636 1432
rect 710 1436 716 1437
rect 710 1432 711 1436
rect 715 1432 716 1436
rect 710 1431 716 1432
rect 798 1436 804 1437
rect 798 1432 799 1436
rect 803 1432 804 1436
rect 798 1431 804 1432
rect 886 1436 892 1437
rect 886 1432 887 1436
rect 891 1432 892 1436
rect 886 1431 892 1432
rect 974 1436 980 1437
rect 974 1432 975 1436
rect 979 1432 980 1436
rect 974 1431 980 1432
rect 1046 1436 1052 1437
rect 1046 1432 1047 1436
rect 1051 1432 1052 1436
rect 1278 1436 1284 1437
rect 1046 1431 1052 1432
rect 1094 1433 1100 1434
rect 110 1428 116 1429
rect 1094 1429 1095 1433
rect 1099 1429 1100 1433
rect 1278 1432 1279 1436
rect 1283 1432 1284 1436
rect 1278 1431 1284 1432
rect 1326 1436 1332 1437
rect 1326 1432 1327 1436
rect 1331 1432 1332 1436
rect 1326 1431 1332 1432
rect 1382 1436 1388 1437
rect 1382 1432 1383 1436
rect 1387 1432 1388 1436
rect 1382 1431 1388 1432
rect 1438 1436 1444 1437
rect 1438 1432 1439 1436
rect 1443 1432 1444 1436
rect 1438 1431 1444 1432
rect 1494 1436 1500 1437
rect 1494 1432 1495 1436
rect 1499 1432 1500 1436
rect 1494 1431 1500 1432
rect 1550 1436 1556 1437
rect 1550 1432 1551 1436
rect 1555 1432 1556 1436
rect 1550 1431 1556 1432
rect 1606 1436 1612 1437
rect 1606 1432 1607 1436
rect 1611 1432 1612 1436
rect 1606 1431 1612 1432
rect 1670 1436 1676 1437
rect 1670 1432 1671 1436
rect 1675 1432 1676 1436
rect 1670 1431 1676 1432
rect 1734 1436 1740 1437
rect 1734 1432 1735 1436
rect 1739 1432 1740 1436
rect 1734 1431 1740 1432
rect 1806 1436 1812 1437
rect 1806 1432 1807 1436
rect 1811 1432 1812 1436
rect 1806 1431 1812 1432
rect 1886 1436 1892 1437
rect 1886 1432 1887 1436
rect 1891 1432 1892 1436
rect 1886 1431 1892 1432
rect 1974 1436 1980 1437
rect 1974 1432 1975 1436
rect 1979 1432 1980 1436
rect 1974 1431 1980 1432
rect 2062 1436 2068 1437
rect 2062 1432 2063 1436
rect 2067 1432 2068 1436
rect 2062 1431 2068 1432
rect 1094 1428 1100 1429
rect 1134 1428 1140 1429
rect 1134 1424 1135 1428
rect 1139 1424 1140 1428
rect 2118 1428 2124 1429
rect 2118 1424 2119 1428
rect 2123 1424 2124 1428
rect 1134 1423 1140 1424
rect 1303 1423 1309 1424
rect 150 1419 156 1420
rect 110 1416 116 1417
rect 110 1412 111 1416
rect 115 1412 116 1416
rect 150 1415 151 1419
rect 155 1418 156 1419
rect 159 1419 165 1420
rect 159 1418 160 1419
rect 155 1416 160 1418
rect 155 1415 156 1416
rect 150 1414 156 1415
rect 159 1415 160 1416
rect 164 1415 165 1419
rect 159 1414 165 1415
rect 215 1419 221 1420
rect 215 1415 216 1419
rect 220 1418 221 1419
rect 278 1419 284 1420
rect 278 1418 279 1419
rect 220 1416 279 1418
rect 220 1415 221 1416
rect 215 1414 221 1415
rect 278 1415 279 1416
rect 283 1415 284 1419
rect 278 1414 284 1415
rect 287 1419 296 1420
rect 287 1415 288 1419
rect 295 1415 296 1419
rect 287 1414 296 1415
rect 358 1419 365 1420
rect 358 1415 359 1419
rect 364 1415 365 1419
rect 358 1414 365 1415
rect 367 1419 373 1420
rect 367 1415 368 1419
rect 372 1418 373 1419
rect 431 1419 437 1420
rect 431 1418 432 1419
rect 372 1416 432 1418
rect 372 1415 373 1416
rect 367 1414 373 1415
rect 431 1415 432 1416
rect 436 1415 437 1419
rect 431 1414 437 1415
rect 503 1419 509 1420
rect 503 1415 504 1419
rect 508 1418 509 1419
rect 526 1419 532 1420
rect 526 1418 527 1419
rect 508 1416 527 1418
rect 508 1415 509 1416
rect 503 1414 509 1415
rect 526 1415 527 1416
rect 531 1415 532 1419
rect 526 1414 532 1415
rect 575 1419 581 1420
rect 575 1415 576 1419
rect 580 1418 581 1419
rect 654 1419 661 1420
rect 580 1416 651 1418
rect 580 1415 581 1416
rect 575 1414 581 1415
rect 110 1411 116 1412
rect 134 1408 140 1409
rect 134 1404 135 1408
rect 139 1404 140 1408
rect 134 1403 140 1404
rect 190 1408 196 1409
rect 190 1404 191 1408
rect 195 1404 196 1408
rect 190 1403 196 1404
rect 262 1408 268 1409
rect 262 1404 263 1408
rect 267 1404 268 1408
rect 262 1403 268 1404
rect 334 1408 340 1409
rect 334 1404 335 1408
rect 339 1404 340 1408
rect 334 1403 340 1404
rect 406 1408 412 1409
rect 406 1404 407 1408
rect 411 1404 412 1408
rect 406 1403 412 1404
rect 478 1408 484 1409
rect 478 1404 479 1408
rect 483 1404 484 1408
rect 478 1403 484 1404
rect 550 1408 556 1409
rect 550 1404 551 1408
rect 555 1404 556 1408
rect 550 1403 556 1404
rect 630 1408 636 1409
rect 630 1404 631 1408
rect 635 1404 636 1408
rect 649 1406 651 1416
rect 654 1415 655 1419
rect 660 1415 661 1419
rect 654 1414 661 1415
rect 663 1419 669 1420
rect 663 1415 664 1419
rect 668 1418 669 1419
rect 735 1419 741 1420
rect 735 1418 736 1419
rect 668 1416 736 1418
rect 668 1415 669 1416
rect 663 1414 669 1415
rect 735 1415 736 1416
rect 740 1415 741 1419
rect 735 1414 741 1415
rect 823 1419 832 1420
rect 823 1415 824 1419
rect 831 1415 832 1419
rect 823 1414 832 1415
rect 834 1419 840 1420
rect 834 1415 835 1419
rect 839 1418 840 1419
rect 911 1419 917 1420
rect 911 1418 912 1419
rect 839 1416 912 1418
rect 839 1415 840 1416
rect 834 1414 840 1415
rect 911 1415 912 1416
rect 916 1415 917 1419
rect 911 1414 917 1415
rect 999 1419 1005 1420
rect 999 1415 1000 1419
rect 1004 1418 1005 1419
rect 1022 1419 1028 1420
rect 1022 1418 1023 1419
rect 1004 1416 1023 1418
rect 1004 1415 1005 1416
rect 999 1414 1005 1415
rect 1022 1415 1023 1416
rect 1027 1415 1028 1419
rect 1022 1414 1028 1415
rect 1034 1419 1040 1420
rect 1034 1415 1035 1419
rect 1039 1418 1040 1419
rect 1071 1419 1077 1420
rect 1071 1418 1072 1419
rect 1039 1416 1072 1418
rect 1039 1415 1040 1416
rect 1034 1414 1040 1415
rect 1071 1415 1072 1416
rect 1076 1415 1077 1419
rect 1303 1419 1304 1423
rect 1308 1422 1309 1423
rect 1319 1423 1325 1424
rect 1319 1422 1320 1423
rect 1308 1420 1320 1422
rect 1308 1419 1309 1420
rect 1303 1418 1309 1419
rect 1319 1419 1320 1420
rect 1324 1419 1325 1423
rect 1319 1418 1325 1419
rect 1342 1423 1348 1424
rect 1342 1419 1343 1423
rect 1347 1422 1348 1423
rect 1351 1423 1357 1424
rect 1351 1422 1352 1423
rect 1347 1420 1352 1422
rect 1347 1419 1348 1420
rect 1342 1418 1348 1419
rect 1351 1419 1352 1420
rect 1356 1419 1357 1423
rect 1351 1418 1357 1419
rect 1398 1423 1404 1424
rect 1398 1419 1399 1423
rect 1403 1422 1404 1423
rect 1407 1423 1413 1424
rect 1407 1422 1408 1423
rect 1403 1420 1408 1422
rect 1403 1419 1404 1420
rect 1398 1418 1404 1419
rect 1407 1419 1408 1420
rect 1412 1419 1413 1423
rect 1407 1418 1413 1419
rect 1446 1423 1452 1424
rect 1446 1419 1447 1423
rect 1451 1422 1452 1423
rect 1463 1423 1469 1424
rect 1463 1422 1464 1423
rect 1451 1420 1464 1422
rect 1451 1419 1452 1420
rect 1446 1418 1452 1419
rect 1463 1419 1464 1420
rect 1468 1419 1469 1423
rect 1463 1418 1469 1419
rect 1510 1423 1516 1424
rect 1510 1419 1511 1423
rect 1515 1422 1516 1423
rect 1519 1423 1525 1424
rect 1519 1422 1520 1423
rect 1515 1420 1520 1422
rect 1515 1419 1516 1420
rect 1510 1418 1516 1419
rect 1519 1419 1520 1420
rect 1524 1419 1525 1423
rect 1519 1418 1525 1419
rect 1575 1423 1584 1424
rect 1575 1419 1576 1423
rect 1583 1419 1584 1423
rect 1575 1418 1584 1419
rect 1614 1423 1620 1424
rect 1614 1419 1615 1423
rect 1619 1422 1620 1423
rect 1631 1423 1637 1424
rect 1631 1422 1632 1423
rect 1619 1420 1632 1422
rect 1619 1419 1620 1420
rect 1614 1418 1620 1419
rect 1631 1419 1632 1420
rect 1636 1419 1637 1423
rect 1631 1418 1637 1419
rect 1686 1423 1692 1424
rect 1686 1419 1687 1423
rect 1691 1422 1692 1423
rect 1695 1423 1701 1424
rect 1695 1422 1696 1423
rect 1691 1420 1696 1422
rect 1691 1419 1692 1420
rect 1686 1418 1692 1419
rect 1695 1419 1696 1420
rect 1700 1419 1701 1423
rect 1695 1418 1701 1419
rect 1759 1423 1765 1424
rect 1759 1419 1760 1423
rect 1764 1422 1765 1423
rect 1767 1423 1773 1424
rect 1767 1422 1768 1423
rect 1764 1420 1768 1422
rect 1764 1419 1765 1420
rect 1759 1418 1765 1419
rect 1767 1419 1768 1420
rect 1772 1419 1773 1423
rect 1767 1418 1773 1419
rect 1831 1423 1837 1424
rect 1831 1419 1832 1423
rect 1836 1422 1837 1423
rect 1839 1423 1845 1424
rect 1839 1422 1840 1423
rect 1836 1420 1840 1422
rect 1836 1419 1837 1420
rect 1831 1418 1837 1419
rect 1839 1419 1840 1420
rect 1844 1419 1845 1423
rect 1839 1418 1845 1419
rect 1910 1423 1917 1424
rect 1910 1419 1911 1423
rect 1916 1419 1917 1423
rect 1910 1418 1917 1419
rect 1999 1423 2005 1424
rect 1999 1419 2000 1423
rect 2004 1422 2005 1423
rect 2014 1423 2020 1424
rect 2014 1422 2015 1423
rect 2004 1420 2015 1422
rect 2004 1419 2005 1420
rect 1999 1418 2005 1419
rect 2014 1419 2015 1420
rect 2019 1419 2020 1423
rect 2014 1418 2020 1419
rect 2078 1423 2084 1424
rect 2078 1419 2079 1423
rect 2083 1422 2084 1423
rect 2087 1423 2093 1424
rect 2118 1423 2124 1424
rect 2087 1422 2088 1423
rect 2083 1420 2088 1422
rect 2083 1419 2084 1420
rect 2078 1418 2084 1419
rect 2087 1419 2088 1420
rect 2092 1419 2093 1423
rect 2087 1418 2093 1419
rect 1071 1414 1077 1415
rect 1094 1416 1100 1417
rect 1094 1412 1095 1416
rect 1099 1412 1100 1416
rect 1094 1411 1100 1412
rect 1134 1411 1140 1412
rect 710 1408 716 1409
rect 649 1404 674 1406
rect 630 1403 636 1404
rect 158 1399 165 1400
rect 158 1395 159 1399
rect 164 1395 165 1399
rect 158 1394 165 1395
rect 202 1399 208 1400
rect 202 1395 203 1399
rect 207 1398 208 1399
rect 215 1399 221 1400
rect 215 1398 216 1399
rect 207 1396 216 1398
rect 207 1395 208 1396
rect 202 1394 208 1395
rect 215 1395 216 1396
rect 220 1395 221 1399
rect 215 1394 221 1395
rect 278 1399 284 1400
rect 278 1395 279 1399
rect 283 1398 284 1399
rect 287 1399 293 1400
rect 287 1398 288 1399
rect 283 1396 288 1398
rect 283 1395 284 1396
rect 278 1394 284 1395
rect 287 1395 288 1396
rect 292 1395 293 1399
rect 287 1394 293 1395
rect 359 1399 365 1400
rect 359 1395 360 1399
rect 364 1398 365 1399
rect 367 1399 373 1400
rect 367 1398 368 1399
rect 364 1396 368 1398
rect 364 1395 365 1396
rect 359 1394 365 1395
rect 367 1395 368 1396
rect 372 1395 373 1399
rect 367 1394 373 1395
rect 431 1399 437 1400
rect 431 1395 432 1399
rect 436 1398 437 1399
rect 446 1399 452 1400
rect 446 1398 447 1399
rect 436 1396 447 1398
rect 436 1395 437 1396
rect 431 1394 437 1395
rect 446 1395 447 1396
rect 451 1395 452 1399
rect 446 1394 452 1395
rect 503 1399 509 1400
rect 503 1395 504 1399
rect 508 1395 509 1399
rect 503 1394 509 1395
rect 575 1399 581 1400
rect 575 1395 576 1399
rect 580 1398 581 1399
rect 598 1399 604 1400
rect 598 1398 599 1399
rect 580 1396 599 1398
rect 580 1395 581 1396
rect 575 1394 581 1395
rect 598 1395 599 1396
rect 603 1395 604 1399
rect 598 1394 604 1395
rect 655 1399 661 1400
rect 655 1395 656 1399
rect 660 1398 661 1399
rect 663 1399 669 1400
rect 663 1398 664 1399
rect 660 1396 664 1398
rect 660 1395 661 1396
rect 655 1394 661 1395
rect 663 1395 664 1396
rect 668 1395 669 1399
rect 672 1398 674 1404
rect 710 1404 711 1408
rect 715 1404 716 1408
rect 710 1403 716 1404
rect 798 1408 804 1409
rect 798 1404 799 1408
rect 803 1404 804 1408
rect 798 1403 804 1404
rect 886 1408 892 1409
rect 886 1404 887 1408
rect 891 1404 892 1408
rect 886 1403 892 1404
rect 974 1408 980 1409
rect 974 1404 975 1408
rect 979 1404 980 1408
rect 974 1403 980 1404
rect 1046 1408 1052 1409
rect 1046 1404 1047 1408
rect 1051 1404 1052 1408
rect 1134 1407 1135 1411
rect 1139 1407 1140 1411
rect 2118 1411 2124 1412
rect 1134 1406 1140 1407
rect 1278 1408 1284 1409
rect 1046 1403 1052 1404
rect 1278 1404 1279 1408
rect 1283 1404 1284 1408
rect 1278 1403 1284 1404
rect 1326 1408 1332 1409
rect 1326 1404 1327 1408
rect 1331 1404 1332 1408
rect 1326 1403 1332 1404
rect 1382 1408 1388 1409
rect 1382 1404 1383 1408
rect 1387 1404 1388 1408
rect 1382 1403 1388 1404
rect 1438 1408 1444 1409
rect 1438 1404 1439 1408
rect 1443 1404 1444 1408
rect 1438 1403 1444 1404
rect 1494 1408 1500 1409
rect 1494 1404 1495 1408
rect 1499 1404 1500 1408
rect 1494 1403 1500 1404
rect 1550 1408 1556 1409
rect 1550 1404 1551 1408
rect 1555 1404 1556 1408
rect 1550 1403 1556 1404
rect 1606 1408 1612 1409
rect 1606 1404 1607 1408
rect 1611 1404 1612 1408
rect 1606 1403 1612 1404
rect 1670 1408 1676 1409
rect 1670 1404 1671 1408
rect 1675 1404 1676 1408
rect 1670 1403 1676 1404
rect 1734 1408 1740 1409
rect 1734 1404 1735 1408
rect 1739 1404 1740 1408
rect 1734 1403 1740 1404
rect 1806 1408 1812 1409
rect 1806 1404 1807 1408
rect 1811 1404 1812 1408
rect 1806 1403 1812 1404
rect 1886 1408 1892 1409
rect 1886 1404 1887 1408
rect 1891 1404 1892 1408
rect 1886 1403 1892 1404
rect 1974 1408 1980 1409
rect 1974 1404 1975 1408
rect 1979 1404 1980 1408
rect 1974 1403 1980 1404
rect 2062 1408 2068 1409
rect 2062 1404 2063 1408
rect 2067 1404 2068 1408
rect 2118 1407 2119 1411
rect 2123 1407 2124 1411
rect 2118 1406 2124 1407
rect 2062 1403 2068 1404
rect 735 1399 741 1400
rect 735 1398 736 1399
rect 672 1396 736 1398
rect 663 1394 669 1395
rect 735 1395 736 1396
rect 740 1395 741 1399
rect 735 1394 741 1395
rect 823 1399 829 1400
rect 823 1395 824 1399
rect 828 1398 829 1399
rect 834 1399 840 1400
rect 834 1398 835 1399
rect 828 1396 835 1398
rect 828 1395 829 1396
rect 823 1394 829 1395
rect 834 1395 835 1396
rect 839 1395 840 1399
rect 834 1394 840 1395
rect 911 1399 917 1400
rect 911 1395 912 1399
rect 916 1398 917 1399
rect 950 1399 956 1400
rect 950 1398 951 1399
rect 916 1396 951 1398
rect 916 1395 917 1396
rect 911 1394 917 1395
rect 950 1395 951 1396
rect 955 1395 956 1399
rect 950 1394 956 1395
rect 999 1399 1005 1400
rect 999 1395 1000 1399
rect 1004 1398 1005 1399
rect 1034 1399 1040 1400
rect 1034 1398 1035 1399
rect 1004 1396 1035 1398
rect 1004 1395 1005 1396
rect 999 1394 1005 1395
rect 1034 1395 1035 1396
rect 1039 1395 1040 1399
rect 1034 1394 1040 1395
rect 1070 1399 1077 1400
rect 1070 1395 1071 1399
rect 1076 1395 1077 1399
rect 1070 1394 1077 1395
rect 358 1391 364 1392
rect 358 1387 359 1391
rect 363 1390 364 1391
rect 505 1390 507 1394
rect 1334 1392 1340 1393
rect 363 1388 507 1390
rect 1134 1389 1140 1390
rect 363 1387 364 1388
rect 358 1386 364 1387
rect 1134 1385 1135 1389
rect 1139 1385 1140 1389
rect 1334 1388 1335 1392
rect 1339 1388 1340 1392
rect 1334 1387 1340 1388
rect 1374 1392 1380 1393
rect 1374 1388 1375 1392
rect 1379 1388 1380 1392
rect 1374 1387 1380 1388
rect 1414 1392 1420 1393
rect 1414 1388 1415 1392
rect 1419 1388 1420 1392
rect 1414 1387 1420 1388
rect 1454 1392 1460 1393
rect 1454 1388 1455 1392
rect 1459 1388 1460 1392
rect 1454 1387 1460 1388
rect 1494 1392 1500 1393
rect 1494 1388 1495 1392
rect 1499 1388 1500 1392
rect 1494 1387 1500 1388
rect 1534 1392 1540 1393
rect 1534 1388 1535 1392
rect 1539 1388 1540 1392
rect 1534 1387 1540 1388
rect 1582 1392 1588 1393
rect 1582 1388 1583 1392
rect 1587 1388 1588 1392
rect 1582 1387 1588 1388
rect 1646 1392 1652 1393
rect 1646 1388 1647 1392
rect 1651 1388 1652 1392
rect 1646 1387 1652 1388
rect 1718 1392 1724 1393
rect 1718 1388 1719 1392
rect 1723 1388 1724 1392
rect 1718 1387 1724 1388
rect 1806 1392 1812 1393
rect 1806 1388 1807 1392
rect 1811 1388 1812 1392
rect 1806 1387 1812 1388
rect 1894 1392 1900 1393
rect 1894 1388 1895 1392
rect 1899 1388 1900 1392
rect 1894 1387 1900 1388
rect 1990 1392 1996 1393
rect 1990 1388 1991 1392
rect 1995 1388 1996 1392
rect 1990 1387 1996 1388
rect 2070 1392 2076 1393
rect 2070 1388 2071 1392
rect 2075 1388 2076 1392
rect 2070 1387 2076 1388
rect 2118 1389 2124 1390
rect 1134 1384 1140 1385
rect 2118 1385 2119 1389
rect 2123 1385 2124 1389
rect 2118 1384 2124 1385
rect 1918 1383 1924 1384
rect 1918 1382 1919 1383
rect 1737 1380 1919 1382
rect 150 1379 156 1380
rect 150 1375 151 1379
rect 155 1378 156 1379
rect 159 1379 165 1380
rect 159 1378 160 1379
rect 155 1376 160 1378
rect 155 1375 156 1376
rect 150 1374 156 1375
rect 159 1375 160 1376
rect 164 1375 165 1379
rect 159 1374 165 1375
rect 199 1379 205 1380
rect 199 1375 200 1379
rect 204 1378 205 1379
rect 250 1379 256 1380
rect 250 1378 251 1379
rect 204 1376 251 1378
rect 204 1375 205 1376
rect 199 1374 205 1375
rect 250 1375 251 1376
rect 255 1375 256 1379
rect 250 1374 256 1375
rect 263 1379 269 1380
rect 263 1375 264 1379
rect 268 1378 269 1379
rect 327 1379 333 1380
rect 268 1376 321 1378
rect 268 1375 269 1376
rect 263 1374 269 1375
rect 134 1372 140 1373
rect 134 1368 135 1372
rect 139 1368 140 1372
rect 134 1367 140 1368
rect 174 1372 180 1373
rect 174 1368 175 1372
rect 179 1368 180 1372
rect 174 1367 180 1368
rect 238 1372 244 1373
rect 238 1368 239 1372
rect 243 1368 244 1372
rect 238 1367 244 1368
rect 302 1372 308 1373
rect 302 1368 303 1372
rect 307 1368 308 1372
rect 319 1370 321 1376
rect 327 1375 328 1379
rect 332 1378 333 1379
rect 382 1379 388 1380
rect 382 1378 383 1379
rect 332 1376 383 1378
rect 332 1375 333 1376
rect 327 1374 333 1375
rect 382 1375 383 1376
rect 387 1375 388 1379
rect 382 1374 388 1375
rect 391 1379 397 1380
rect 391 1375 392 1379
rect 396 1378 397 1379
rect 454 1379 460 1380
rect 454 1378 455 1379
rect 396 1376 455 1378
rect 396 1375 397 1376
rect 391 1374 397 1375
rect 454 1375 455 1376
rect 459 1375 460 1379
rect 454 1374 460 1375
rect 463 1379 469 1380
rect 463 1375 464 1379
rect 468 1378 469 1379
rect 510 1379 516 1380
rect 510 1378 511 1379
rect 468 1376 511 1378
rect 468 1375 469 1376
rect 463 1374 469 1375
rect 510 1375 511 1376
rect 515 1375 516 1379
rect 510 1374 516 1375
rect 526 1379 533 1380
rect 526 1375 527 1379
rect 532 1375 533 1379
rect 526 1374 533 1375
rect 599 1379 605 1380
rect 599 1375 600 1379
rect 604 1378 605 1379
rect 662 1379 668 1380
rect 662 1378 663 1379
rect 604 1376 663 1378
rect 604 1375 605 1376
rect 599 1374 605 1375
rect 662 1375 663 1376
rect 667 1375 668 1379
rect 662 1374 668 1375
rect 671 1379 677 1380
rect 671 1375 672 1379
rect 676 1378 677 1379
rect 718 1379 724 1380
rect 718 1378 719 1379
rect 676 1376 719 1378
rect 676 1375 677 1376
rect 671 1374 677 1375
rect 718 1375 719 1376
rect 723 1375 724 1379
rect 718 1374 724 1375
rect 730 1379 741 1380
rect 730 1375 731 1379
rect 735 1375 736 1379
rect 740 1375 741 1379
rect 730 1374 741 1375
rect 806 1379 813 1380
rect 806 1375 807 1379
rect 812 1375 813 1379
rect 806 1374 813 1375
rect 815 1379 821 1380
rect 815 1375 816 1379
rect 820 1378 821 1379
rect 879 1379 885 1380
rect 879 1378 880 1379
rect 820 1376 880 1378
rect 820 1375 821 1376
rect 815 1374 821 1375
rect 879 1375 880 1376
rect 884 1375 885 1379
rect 879 1374 885 1375
rect 890 1379 896 1380
rect 890 1375 891 1379
rect 895 1378 896 1379
rect 951 1379 957 1380
rect 951 1378 952 1379
rect 895 1376 952 1378
rect 895 1375 896 1376
rect 890 1374 896 1375
rect 951 1375 952 1376
rect 956 1375 957 1379
rect 951 1374 957 1375
rect 1022 1379 1029 1380
rect 1022 1375 1023 1379
rect 1028 1375 1029 1379
rect 1022 1374 1029 1375
rect 1031 1379 1037 1380
rect 1031 1375 1032 1379
rect 1036 1378 1037 1379
rect 1071 1379 1077 1380
rect 1071 1378 1072 1379
rect 1036 1376 1072 1378
rect 1036 1375 1037 1376
rect 1031 1374 1037 1375
rect 1071 1375 1072 1376
rect 1076 1375 1077 1379
rect 1071 1374 1077 1375
rect 1359 1375 1365 1376
rect 366 1372 372 1373
rect 358 1371 364 1372
rect 358 1370 359 1371
rect 319 1368 359 1370
rect 302 1367 308 1368
rect 358 1367 359 1368
rect 363 1367 364 1371
rect 366 1368 367 1372
rect 371 1368 372 1372
rect 366 1367 372 1368
rect 438 1372 444 1373
rect 438 1368 439 1372
rect 443 1368 444 1372
rect 438 1367 444 1368
rect 502 1372 508 1373
rect 502 1368 503 1372
rect 507 1368 508 1372
rect 502 1367 508 1368
rect 574 1372 580 1373
rect 574 1368 575 1372
rect 579 1368 580 1372
rect 574 1367 580 1368
rect 646 1372 652 1373
rect 646 1368 647 1372
rect 651 1368 652 1372
rect 646 1367 652 1368
rect 710 1372 716 1373
rect 710 1368 711 1372
rect 715 1368 716 1372
rect 710 1367 716 1368
rect 782 1372 788 1373
rect 782 1368 783 1372
rect 787 1368 788 1372
rect 782 1367 788 1368
rect 854 1372 860 1373
rect 854 1368 855 1372
rect 859 1368 860 1372
rect 854 1367 860 1368
rect 926 1372 932 1373
rect 926 1368 927 1372
rect 931 1368 932 1372
rect 926 1367 932 1368
rect 998 1372 1004 1373
rect 998 1368 999 1372
rect 1003 1368 1004 1372
rect 998 1367 1004 1368
rect 1046 1372 1052 1373
rect 1046 1368 1047 1372
rect 1051 1368 1052 1372
rect 1046 1367 1052 1368
rect 1134 1372 1140 1373
rect 1134 1368 1135 1372
rect 1139 1368 1140 1372
rect 1359 1371 1360 1375
rect 1364 1374 1365 1375
rect 1390 1375 1396 1376
rect 1390 1374 1391 1375
rect 1364 1372 1391 1374
rect 1364 1371 1365 1372
rect 1359 1370 1365 1371
rect 1390 1371 1391 1372
rect 1395 1371 1396 1375
rect 1390 1370 1396 1371
rect 1399 1375 1405 1376
rect 1399 1371 1400 1375
rect 1404 1374 1405 1375
rect 1422 1375 1428 1376
rect 1422 1374 1423 1375
rect 1404 1372 1423 1374
rect 1404 1371 1405 1372
rect 1399 1370 1405 1371
rect 1422 1371 1423 1372
rect 1427 1371 1428 1375
rect 1422 1370 1428 1371
rect 1430 1375 1436 1376
rect 1430 1371 1431 1375
rect 1435 1374 1436 1375
rect 1439 1375 1445 1376
rect 1439 1374 1440 1375
rect 1435 1372 1440 1374
rect 1435 1371 1436 1372
rect 1430 1370 1436 1371
rect 1439 1371 1440 1372
rect 1444 1371 1445 1375
rect 1439 1370 1445 1371
rect 1479 1375 1488 1376
rect 1479 1371 1480 1375
rect 1487 1371 1488 1375
rect 1479 1370 1488 1371
rect 1502 1375 1508 1376
rect 1502 1371 1503 1375
rect 1507 1374 1508 1375
rect 1519 1375 1525 1376
rect 1519 1374 1520 1375
rect 1507 1372 1520 1374
rect 1507 1371 1508 1372
rect 1502 1370 1508 1371
rect 1519 1371 1520 1372
rect 1524 1371 1525 1375
rect 1519 1370 1525 1371
rect 1542 1375 1548 1376
rect 1542 1371 1543 1375
rect 1547 1374 1548 1375
rect 1559 1375 1565 1376
rect 1559 1374 1560 1375
rect 1547 1372 1560 1374
rect 1547 1371 1548 1372
rect 1542 1370 1548 1371
rect 1559 1371 1560 1372
rect 1564 1371 1565 1375
rect 1559 1370 1565 1371
rect 1607 1375 1613 1376
rect 1607 1371 1608 1375
rect 1612 1374 1613 1375
rect 1662 1375 1668 1376
rect 1662 1374 1663 1375
rect 1612 1372 1663 1374
rect 1612 1371 1613 1372
rect 1607 1370 1613 1371
rect 1662 1371 1663 1372
rect 1667 1371 1668 1375
rect 1662 1370 1668 1371
rect 1671 1375 1677 1376
rect 1671 1371 1672 1375
rect 1676 1374 1677 1375
rect 1737 1374 1739 1380
rect 1918 1379 1919 1380
rect 1923 1379 1924 1383
rect 1918 1378 1924 1379
rect 1676 1372 1739 1374
rect 1742 1375 1749 1376
rect 1676 1371 1677 1372
rect 1671 1370 1677 1371
rect 1742 1371 1743 1375
rect 1748 1371 1749 1375
rect 1742 1370 1749 1371
rect 1751 1375 1757 1376
rect 1751 1371 1752 1375
rect 1756 1374 1757 1375
rect 1831 1375 1837 1376
rect 1831 1374 1832 1375
rect 1756 1372 1832 1374
rect 1756 1371 1757 1372
rect 1751 1370 1757 1371
rect 1831 1371 1832 1372
rect 1836 1371 1837 1375
rect 1831 1370 1837 1371
rect 1839 1375 1845 1376
rect 1839 1371 1840 1375
rect 1844 1374 1845 1375
rect 1919 1375 1925 1376
rect 1919 1374 1920 1375
rect 1844 1372 1920 1374
rect 1844 1371 1845 1372
rect 1839 1370 1845 1371
rect 1919 1371 1920 1372
rect 1924 1371 1925 1375
rect 1919 1370 1925 1371
rect 2015 1375 2021 1376
rect 2015 1371 2016 1375
rect 2020 1374 2021 1375
rect 2086 1375 2092 1376
rect 2086 1374 2087 1375
rect 2020 1372 2087 1374
rect 2020 1371 2021 1372
rect 2015 1370 2021 1371
rect 2086 1371 2087 1372
rect 2091 1371 2092 1375
rect 2086 1370 2092 1371
rect 2094 1375 2101 1376
rect 2094 1371 2095 1375
rect 2100 1371 2101 1375
rect 2094 1370 2101 1371
rect 2118 1372 2124 1373
rect 1134 1367 1140 1368
rect 2118 1368 2119 1372
rect 2123 1368 2124 1372
rect 2118 1367 2124 1368
rect 358 1366 364 1367
rect 110 1364 116 1365
rect 110 1360 111 1364
rect 115 1360 116 1364
rect 1094 1364 1100 1365
rect 1094 1360 1095 1364
rect 1099 1360 1100 1364
rect 110 1359 116 1360
rect 158 1359 165 1360
rect 158 1355 159 1359
rect 164 1355 165 1359
rect 158 1354 165 1355
rect 199 1359 208 1360
rect 199 1355 200 1359
rect 207 1355 208 1359
rect 199 1354 208 1355
rect 250 1359 256 1360
rect 250 1355 251 1359
rect 255 1358 256 1359
rect 263 1359 269 1360
rect 263 1358 264 1359
rect 255 1356 264 1358
rect 255 1355 256 1356
rect 250 1354 256 1355
rect 263 1355 264 1356
rect 268 1355 269 1359
rect 263 1354 269 1355
rect 327 1359 333 1360
rect 327 1355 328 1359
rect 332 1358 333 1359
rect 374 1359 380 1360
rect 374 1358 375 1359
rect 332 1356 375 1358
rect 332 1355 333 1356
rect 327 1354 333 1355
rect 374 1355 375 1356
rect 379 1355 380 1359
rect 374 1354 380 1355
rect 382 1359 388 1360
rect 382 1355 383 1359
rect 387 1358 388 1359
rect 391 1359 397 1360
rect 391 1358 392 1359
rect 387 1356 392 1358
rect 387 1355 388 1356
rect 382 1354 388 1355
rect 391 1355 392 1356
rect 396 1355 397 1359
rect 391 1354 397 1355
rect 454 1359 460 1360
rect 454 1355 455 1359
rect 459 1358 460 1359
rect 463 1359 469 1360
rect 463 1358 464 1359
rect 459 1356 464 1358
rect 459 1355 460 1356
rect 454 1354 460 1355
rect 463 1355 464 1356
rect 468 1355 469 1359
rect 463 1354 469 1355
rect 510 1359 516 1360
rect 510 1355 511 1359
rect 515 1358 516 1359
rect 527 1359 533 1360
rect 527 1358 528 1359
rect 515 1356 528 1358
rect 515 1355 516 1356
rect 510 1354 516 1355
rect 527 1355 528 1356
rect 532 1355 533 1359
rect 527 1354 533 1355
rect 598 1359 605 1360
rect 598 1355 599 1359
rect 604 1355 605 1359
rect 598 1354 605 1355
rect 662 1359 668 1360
rect 662 1355 663 1359
rect 667 1358 668 1359
rect 671 1359 677 1360
rect 671 1358 672 1359
rect 667 1356 672 1358
rect 667 1355 668 1356
rect 662 1354 668 1355
rect 671 1355 672 1356
rect 676 1355 677 1359
rect 671 1354 677 1355
rect 718 1359 724 1360
rect 718 1355 719 1359
rect 723 1358 724 1359
rect 735 1359 741 1360
rect 735 1358 736 1359
rect 723 1356 736 1358
rect 723 1355 724 1356
rect 718 1354 724 1355
rect 735 1355 736 1356
rect 740 1355 741 1359
rect 735 1354 741 1355
rect 807 1359 813 1360
rect 807 1355 808 1359
rect 812 1358 813 1359
rect 815 1359 821 1360
rect 815 1358 816 1359
rect 812 1356 816 1358
rect 812 1355 813 1356
rect 807 1354 813 1355
rect 815 1355 816 1356
rect 820 1355 821 1359
rect 815 1354 821 1355
rect 879 1359 885 1360
rect 879 1355 880 1359
rect 884 1358 885 1359
rect 890 1359 896 1360
rect 890 1358 891 1359
rect 884 1356 891 1358
rect 884 1355 885 1356
rect 879 1354 885 1355
rect 890 1355 891 1356
rect 895 1355 896 1359
rect 890 1354 896 1355
rect 950 1359 957 1360
rect 950 1355 951 1359
rect 956 1355 957 1359
rect 950 1354 957 1355
rect 1023 1359 1029 1360
rect 1023 1355 1024 1359
rect 1028 1358 1029 1359
rect 1031 1359 1037 1360
rect 1031 1358 1032 1359
rect 1028 1356 1032 1358
rect 1028 1355 1029 1356
rect 1023 1354 1029 1355
rect 1031 1355 1032 1356
rect 1036 1355 1037 1359
rect 1031 1354 1037 1355
rect 1071 1359 1077 1360
rect 1071 1355 1072 1359
rect 1076 1358 1077 1359
rect 1086 1359 1092 1360
rect 1094 1359 1100 1360
rect 1334 1364 1340 1365
rect 1334 1360 1335 1364
rect 1339 1360 1340 1364
rect 1334 1359 1340 1360
rect 1374 1364 1380 1365
rect 1374 1360 1375 1364
rect 1379 1360 1380 1364
rect 1374 1359 1380 1360
rect 1414 1364 1420 1365
rect 1414 1360 1415 1364
rect 1419 1360 1420 1364
rect 1414 1359 1420 1360
rect 1454 1364 1460 1365
rect 1454 1360 1455 1364
rect 1459 1360 1460 1364
rect 1454 1359 1460 1360
rect 1494 1364 1500 1365
rect 1494 1360 1495 1364
rect 1499 1360 1500 1364
rect 1494 1359 1500 1360
rect 1534 1364 1540 1365
rect 1534 1360 1535 1364
rect 1539 1360 1540 1364
rect 1534 1359 1540 1360
rect 1582 1364 1588 1365
rect 1582 1360 1583 1364
rect 1587 1360 1588 1364
rect 1582 1359 1588 1360
rect 1646 1364 1652 1365
rect 1646 1360 1647 1364
rect 1651 1360 1652 1364
rect 1646 1359 1652 1360
rect 1718 1364 1724 1365
rect 1718 1360 1719 1364
rect 1723 1360 1724 1364
rect 1718 1359 1724 1360
rect 1806 1364 1812 1365
rect 1806 1360 1807 1364
rect 1811 1360 1812 1364
rect 1806 1359 1812 1360
rect 1894 1364 1900 1365
rect 1894 1360 1895 1364
rect 1899 1360 1900 1364
rect 1894 1359 1900 1360
rect 1990 1364 1996 1365
rect 1990 1360 1991 1364
rect 1995 1360 1996 1364
rect 1990 1359 1996 1360
rect 2070 1364 2076 1365
rect 2070 1360 2071 1364
rect 2075 1360 2076 1364
rect 2070 1359 2076 1360
rect 1086 1358 1087 1359
rect 1076 1356 1087 1358
rect 1076 1355 1077 1356
rect 1071 1354 1077 1355
rect 1086 1355 1087 1356
rect 1091 1355 1092 1359
rect 1086 1354 1092 1355
rect 1319 1355 1325 1356
rect 1319 1351 1320 1355
rect 1324 1354 1325 1355
rect 1359 1355 1365 1356
rect 1359 1354 1360 1355
rect 1324 1352 1360 1354
rect 1324 1351 1325 1352
rect 1319 1350 1325 1351
rect 1359 1351 1360 1352
rect 1364 1351 1365 1355
rect 1359 1350 1365 1351
rect 1390 1355 1396 1356
rect 1390 1351 1391 1355
rect 1395 1354 1396 1355
rect 1399 1355 1405 1356
rect 1399 1354 1400 1355
rect 1395 1352 1400 1354
rect 1395 1351 1396 1352
rect 1390 1350 1396 1351
rect 1399 1351 1400 1352
rect 1404 1351 1405 1355
rect 1399 1350 1405 1351
rect 1422 1355 1428 1356
rect 1422 1351 1423 1355
rect 1427 1354 1428 1355
rect 1439 1355 1445 1356
rect 1439 1354 1440 1355
rect 1427 1352 1440 1354
rect 1427 1351 1428 1352
rect 1422 1350 1428 1351
rect 1439 1351 1440 1352
rect 1444 1351 1445 1355
rect 1439 1350 1445 1351
rect 1479 1355 1485 1356
rect 1479 1351 1480 1355
rect 1484 1354 1485 1355
rect 1502 1355 1508 1356
rect 1502 1354 1503 1355
rect 1484 1352 1503 1354
rect 1484 1351 1485 1352
rect 1479 1350 1485 1351
rect 1502 1351 1503 1352
rect 1507 1351 1508 1355
rect 1502 1350 1508 1351
rect 1519 1355 1525 1356
rect 1519 1351 1520 1355
rect 1524 1354 1525 1355
rect 1542 1355 1548 1356
rect 1542 1354 1543 1355
rect 1524 1352 1543 1354
rect 1524 1351 1525 1352
rect 1519 1350 1525 1351
rect 1542 1351 1543 1352
rect 1547 1351 1548 1355
rect 1542 1350 1548 1351
rect 1559 1355 1565 1356
rect 1559 1351 1560 1355
rect 1564 1354 1565 1355
rect 1590 1355 1596 1356
rect 1590 1354 1591 1355
rect 1564 1352 1591 1354
rect 1564 1351 1565 1352
rect 1559 1350 1565 1351
rect 1590 1351 1591 1352
rect 1595 1351 1596 1355
rect 1590 1350 1596 1351
rect 1607 1355 1613 1356
rect 1607 1351 1608 1355
rect 1612 1351 1613 1355
rect 1607 1350 1613 1351
rect 1662 1355 1668 1356
rect 1662 1351 1663 1355
rect 1667 1354 1668 1355
rect 1671 1355 1677 1356
rect 1671 1354 1672 1355
rect 1667 1352 1672 1354
rect 1667 1351 1668 1352
rect 1662 1350 1668 1351
rect 1671 1351 1672 1352
rect 1676 1351 1677 1355
rect 1671 1350 1677 1351
rect 1743 1355 1749 1356
rect 1743 1351 1744 1355
rect 1748 1354 1749 1355
rect 1751 1355 1757 1356
rect 1751 1354 1752 1355
rect 1748 1352 1752 1354
rect 1748 1351 1749 1352
rect 1743 1350 1749 1351
rect 1751 1351 1752 1352
rect 1756 1351 1757 1355
rect 1751 1350 1757 1351
rect 1831 1355 1837 1356
rect 1831 1351 1832 1355
rect 1836 1354 1837 1355
rect 1839 1355 1845 1356
rect 1839 1354 1840 1355
rect 1836 1352 1840 1354
rect 1836 1351 1837 1352
rect 1831 1350 1837 1351
rect 1839 1351 1840 1352
rect 1844 1351 1845 1355
rect 1839 1350 1845 1351
rect 1918 1355 1925 1356
rect 1918 1351 1919 1355
rect 1924 1351 1925 1355
rect 1918 1350 1925 1351
rect 2014 1355 2021 1356
rect 2014 1351 2015 1355
rect 2020 1351 2021 1355
rect 2014 1350 2021 1351
rect 2086 1355 2092 1356
rect 2086 1351 2087 1355
rect 2091 1354 2092 1355
rect 2095 1355 2101 1356
rect 2095 1354 2096 1355
rect 2091 1352 2096 1354
rect 2091 1351 2092 1352
rect 2086 1350 2092 1351
rect 2095 1351 2096 1352
rect 2100 1351 2101 1355
rect 2095 1350 2101 1351
rect 110 1347 116 1348
rect 110 1343 111 1347
rect 115 1343 116 1347
rect 1094 1347 1100 1348
rect 110 1342 116 1343
rect 134 1344 140 1345
rect 134 1340 135 1344
rect 139 1340 140 1344
rect 134 1339 140 1340
rect 174 1344 180 1345
rect 174 1340 175 1344
rect 179 1340 180 1344
rect 174 1339 180 1340
rect 238 1344 244 1345
rect 238 1340 239 1344
rect 243 1340 244 1344
rect 238 1339 244 1340
rect 302 1344 308 1345
rect 302 1340 303 1344
rect 307 1340 308 1344
rect 302 1339 308 1340
rect 366 1344 372 1345
rect 366 1340 367 1344
rect 371 1340 372 1344
rect 366 1339 372 1340
rect 438 1344 444 1345
rect 438 1340 439 1344
rect 443 1340 444 1344
rect 438 1339 444 1340
rect 502 1344 508 1345
rect 502 1340 503 1344
rect 507 1340 508 1344
rect 502 1339 508 1340
rect 574 1344 580 1345
rect 574 1340 575 1344
rect 579 1340 580 1344
rect 574 1339 580 1340
rect 646 1344 652 1345
rect 646 1340 647 1344
rect 651 1340 652 1344
rect 646 1339 652 1340
rect 710 1344 716 1345
rect 710 1340 711 1344
rect 715 1340 716 1344
rect 710 1339 716 1340
rect 782 1344 788 1345
rect 782 1340 783 1344
rect 787 1340 788 1344
rect 782 1339 788 1340
rect 854 1344 860 1345
rect 854 1340 855 1344
rect 859 1340 860 1344
rect 854 1339 860 1340
rect 926 1344 932 1345
rect 926 1340 927 1344
rect 931 1340 932 1344
rect 926 1339 932 1340
rect 998 1344 1004 1345
rect 998 1340 999 1344
rect 1003 1340 1004 1344
rect 998 1339 1004 1340
rect 1046 1344 1052 1345
rect 1046 1340 1047 1344
rect 1051 1340 1052 1344
rect 1094 1343 1095 1347
rect 1099 1343 1100 1347
rect 1094 1342 1100 1343
rect 1482 1347 1488 1348
rect 1482 1343 1483 1347
rect 1487 1346 1488 1347
rect 1609 1346 1611 1350
rect 1487 1344 1611 1346
rect 1487 1343 1488 1344
rect 1482 1342 1488 1343
rect 1046 1339 1052 1340
rect 1086 1335 1092 1336
rect 1086 1331 1087 1335
rect 1091 1334 1092 1335
rect 1183 1335 1189 1336
rect 1183 1334 1184 1335
rect 1091 1332 1184 1334
rect 1091 1331 1092 1332
rect 1086 1330 1092 1331
rect 1183 1331 1184 1332
rect 1188 1331 1189 1335
rect 1183 1330 1189 1331
rect 1191 1335 1197 1336
rect 1191 1331 1192 1335
rect 1196 1334 1197 1335
rect 1247 1335 1253 1336
rect 1247 1334 1248 1335
rect 1196 1332 1248 1334
rect 1196 1331 1197 1332
rect 1191 1330 1197 1331
rect 1247 1331 1248 1332
rect 1252 1331 1253 1335
rect 1247 1330 1253 1331
rect 1255 1335 1261 1336
rect 1255 1331 1256 1335
rect 1260 1334 1261 1335
rect 1335 1335 1341 1336
rect 1335 1334 1336 1335
rect 1260 1332 1336 1334
rect 1260 1331 1261 1332
rect 1255 1330 1261 1331
rect 1335 1331 1336 1332
rect 1340 1331 1341 1335
rect 1335 1330 1341 1331
rect 1430 1335 1437 1336
rect 1430 1331 1431 1335
rect 1436 1331 1437 1335
rect 1430 1330 1437 1331
rect 1439 1335 1445 1336
rect 1439 1331 1440 1335
rect 1444 1334 1445 1335
rect 1527 1335 1533 1336
rect 1527 1334 1528 1335
rect 1444 1332 1528 1334
rect 1444 1331 1445 1332
rect 1439 1330 1445 1331
rect 1527 1331 1528 1332
rect 1532 1331 1533 1335
rect 1527 1330 1533 1331
rect 1535 1335 1541 1336
rect 1535 1331 1536 1335
rect 1540 1334 1541 1335
rect 1623 1335 1629 1336
rect 1623 1334 1624 1335
rect 1540 1332 1624 1334
rect 1540 1331 1541 1332
rect 1535 1330 1541 1331
rect 1623 1331 1624 1332
rect 1628 1331 1629 1335
rect 1623 1330 1629 1331
rect 1703 1335 1709 1336
rect 1703 1331 1704 1335
rect 1708 1334 1709 1335
rect 1774 1335 1780 1336
rect 1774 1334 1775 1335
rect 1708 1332 1775 1334
rect 1708 1331 1709 1332
rect 1703 1330 1709 1331
rect 1774 1331 1775 1332
rect 1779 1331 1780 1335
rect 1774 1330 1780 1331
rect 1783 1335 1789 1336
rect 1783 1331 1784 1335
rect 1788 1334 1789 1335
rect 1846 1335 1852 1336
rect 1846 1334 1847 1335
rect 1788 1332 1847 1334
rect 1788 1331 1789 1332
rect 1783 1330 1789 1331
rect 1846 1331 1847 1332
rect 1851 1331 1852 1335
rect 1846 1330 1852 1331
rect 1855 1335 1861 1336
rect 1855 1331 1856 1335
rect 1860 1334 1861 1335
rect 1910 1335 1916 1336
rect 1910 1334 1911 1335
rect 1860 1332 1911 1334
rect 1860 1331 1861 1332
rect 1855 1330 1861 1331
rect 1910 1331 1911 1332
rect 1915 1331 1916 1335
rect 1910 1330 1916 1331
rect 1919 1335 1925 1336
rect 1919 1331 1920 1335
rect 1924 1334 1925 1335
rect 1974 1335 1980 1336
rect 1974 1334 1975 1335
rect 1924 1332 1975 1334
rect 1924 1331 1925 1332
rect 1919 1330 1925 1331
rect 1974 1331 1975 1332
rect 1979 1331 1980 1335
rect 1974 1330 1980 1331
rect 1983 1335 1989 1336
rect 1983 1331 1984 1335
rect 1988 1334 1989 1335
rect 2038 1335 2044 1336
rect 2038 1334 2039 1335
rect 1988 1332 2039 1334
rect 1988 1331 1989 1332
rect 1983 1330 1989 1331
rect 2038 1331 2039 1332
rect 2043 1331 2044 1335
rect 2038 1330 2044 1331
rect 2046 1335 2053 1336
rect 2046 1331 2047 1335
rect 2052 1331 2053 1335
rect 2046 1330 2053 1331
rect 2094 1335 2101 1336
rect 2094 1331 2095 1335
rect 2100 1331 2101 1335
rect 2094 1330 2101 1331
rect 1158 1328 1164 1329
rect 134 1324 140 1325
rect 110 1321 116 1322
rect 110 1317 111 1321
rect 115 1317 116 1321
rect 134 1320 135 1324
rect 139 1320 140 1324
rect 134 1319 140 1320
rect 174 1324 180 1325
rect 174 1320 175 1324
rect 179 1320 180 1324
rect 174 1319 180 1320
rect 214 1324 220 1325
rect 214 1320 215 1324
rect 219 1320 220 1324
rect 214 1319 220 1320
rect 254 1324 260 1325
rect 254 1320 255 1324
rect 259 1320 260 1324
rect 254 1319 260 1320
rect 318 1324 324 1325
rect 318 1320 319 1324
rect 323 1320 324 1324
rect 318 1319 324 1320
rect 390 1324 396 1325
rect 390 1320 391 1324
rect 395 1320 396 1324
rect 390 1319 396 1320
rect 462 1324 468 1325
rect 462 1320 463 1324
rect 467 1320 468 1324
rect 462 1319 468 1320
rect 542 1324 548 1325
rect 542 1320 543 1324
rect 547 1320 548 1324
rect 542 1319 548 1320
rect 622 1324 628 1325
rect 622 1320 623 1324
rect 627 1320 628 1324
rect 622 1319 628 1320
rect 702 1324 708 1325
rect 702 1320 703 1324
rect 707 1320 708 1324
rect 702 1319 708 1320
rect 782 1324 788 1325
rect 782 1320 783 1324
rect 787 1320 788 1324
rect 782 1319 788 1320
rect 862 1324 868 1325
rect 862 1320 863 1324
rect 867 1320 868 1324
rect 862 1319 868 1320
rect 942 1324 948 1325
rect 942 1320 943 1324
rect 947 1320 948 1324
rect 942 1319 948 1320
rect 1022 1324 1028 1325
rect 1022 1320 1023 1324
rect 1027 1320 1028 1324
rect 1158 1324 1159 1328
rect 1163 1324 1164 1328
rect 1158 1323 1164 1324
rect 1222 1328 1228 1329
rect 1222 1324 1223 1328
rect 1227 1324 1228 1328
rect 1222 1323 1228 1324
rect 1310 1328 1316 1329
rect 1310 1324 1311 1328
rect 1315 1324 1316 1328
rect 1310 1323 1316 1324
rect 1406 1328 1412 1329
rect 1406 1324 1407 1328
rect 1411 1324 1412 1328
rect 1406 1323 1412 1324
rect 1502 1328 1508 1329
rect 1502 1324 1503 1328
rect 1507 1324 1508 1328
rect 1502 1323 1508 1324
rect 1598 1328 1604 1329
rect 1598 1324 1599 1328
rect 1603 1324 1604 1328
rect 1598 1323 1604 1324
rect 1678 1328 1684 1329
rect 1678 1324 1679 1328
rect 1683 1324 1684 1328
rect 1678 1323 1684 1324
rect 1758 1328 1764 1329
rect 1758 1324 1759 1328
rect 1763 1324 1764 1328
rect 1758 1323 1764 1324
rect 1830 1328 1836 1329
rect 1830 1324 1831 1328
rect 1835 1324 1836 1328
rect 1830 1323 1836 1324
rect 1894 1328 1900 1329
rect 1894 1324 1895 1328
rect 1899 1324 1900 1328
rect 1894 1323 1900 1324
rect 1958 1328 1964 1329
rect 1958 1324 1959 1328
rect 1963 1324 1964 1328
rect 1958 1323 1964 1324
rect 2022 1328 2028 1329
rect 2022 1324 2023 1328
rect 2027 1324 2028 1328
rect 2022 1323 2028 1324
rect 2070 1328 2076 1329
rect 2070 1324 2071 1328
rect 2075 1324 2076 1328
rect 2070 1323 2076 1324
rect 1022 1319 1028 1320
rect 1094 1321 1100 1322
rect 110 1316 116 1317
rect 1094 1317 1095 1321
rect 1099 1317 1100 1321
rect 1094 1316 1100 1317
rect 1134 1320 1140 1321
rect 1134 1316 1135 1320
rect 1139 1316 1140 1320
rect 2118 1320 2124 1321
rect 2118 1316 2119 1320
rect 2123 1316 2124 1320
rect 342 1315 348 1316
rect 1134 1315 1140 1316
rect 1183 1315 1189 1316
rect 342 1314 343 1315
rect 272 1312 343 1314
rect 159 1307 165 1308
rect 110 1304 116 1305
rect 110 1300 111 1304
rect 115 1300 116 1304
rect 159 1303 160 1307
rect 164 1306 165 1307
rect 190 1307 196 1308
rect 190 1306 191 1307
rect 164 1304 191 1306
rect 164 1303 165 1304
rect 159 1302 165 1303
rect 190 1303 191 1304
rect 195 1303 196 1307
rect 190 1302 196 1303
rect 199 1307 205 1308
rect 199 1303 200 1307
rect 204 1306 205 1307
rect 230 1307 236 1308
rect 230 1306 231 1307
rect 204 1304 231 1306
rect 204 1303 205 1304
rect 199 1302 205 1303
rect 230 1303 231 1304
rect 235 1303 236 1307
rect 230 1302 236 1303
rect 239 1307 245 1308
rect 239 1303 240 1307
rect 244 1306 245 1307
rect 272 1306 274 1312
rect 342 1311 343 1312
rect 347 1311 348 1315
rect 342 1310 348 1311
rect 1183 1311 1184 1315
rect 1188 1314 1189 1315
rect 1191 1315 1197 1316
rect 1191 1314 1192 1315
rect 1188 1312 1192 1314
rect 1188 1311 1189 1312
rect 1183 1310 1189 1311
rect 1191 1311 1192 1312
rect 1196 1311 1197 1315
rect 1191 1310 1197 1311
rect 1247 1315 1253 1316
rect 1247 1311 1248 1315
rect 1252 1314 1253 1315
rect 1255 1315 1261 1316
rect 1255 1314 1256 1315
rect 1252 1312 1256 1314
rect 1252 1311 1253 1312
rect 1247 1310 1253 1311
rect 1255 1311 1256 1312
rect 1260 1311 1261 1315
rect 1255 1310 1261 1311
rect 1330 1315 1341 1316
rect 1330 1311 1331 1315
rect 1335 1311 1336 1315
rect 1340 1311 1341 1315
rect 1330 1310 1341 1311
rect 1431 1315 1437 1316
rect 1431 1311 1432 1315
rect 1436 1314 1437 1315
rect 1439 1315 1445 1316
rect 1439 1314 1440 1315
rect 1436 1312 1440 1314
rect 1436 1311 1437 1312
rect 1431 1310 1437 1311
rect 1439 1311 1440 1312
rect 1444 1311 1445 1315
rect 1439 1310 1445 1311
rect 1527 1315 1533 1316
rect 1527 1311 1528 1315
rect 1532 1314 1533 1315
rect 1535 1315 1541 1316
rect 1535 1314 1536 1315
rect 1532 1312 1536 1314
rect 1532 1311 1533 1312
rect 1527 1310 1533 1311
rect 1535 1311 1536 1312
rect 1540 1311 1541 1315
rect 1535 1310 1541 1311
rect 1590 1315 1596 1316
rect 1590 1311 1591 1315
rect 1595 1314 1596 1315
rect 1623 1315 1629 1316
rect 1623 1314 1624 1315
rect 1595 1312 1624 1314
rect 1595 1311 1596 1312
rect 1590 1310 1596 1311
rect 1623 1311 1624 1312
rect 1628 1311 1629 1315
rect 1623 1310 1629 1311
rect 1703 1315 1709 1316
rect 1703 1311 1704 1315
rect 1708 1314 1709 1315
rect 1766 1315 1772 1316
rect 1766 1314 1767 1315
rect 1708 1312 1767 1314
rect 1708 1311 1709 1312
rect 1703 1310 1709 1311
rect 1766 1311 1767 1312
rect 1771 1311 1772 1315
rect 1766 1310 1772 1311
rect 1774 1315 1780 1316
rect 1774 1311 1775 1315
rect 1779 1314 1780 1315
rect 1783 1315 1789 1316
rect 1783 1314 1784 1315
rect 1779 1312 1784 1314
rect 1779 1311 1780 1312
rect 1774 1310 1780 1311
rect 1783 1311 1784 1312
rect 1788 1311 1789 1315
rect 1783 1310 1789 1311
rect 1846 1315 1852 1316
rect 1846 1311 1847 1315
rect 1851 1314 1852 1315
rect 1855 1315 1861 1316
rect 1855 1314 1856 1315
rect 1851 1312 1856 1314
rect 1851 1311 1852 1312
rect 1846 1310 1852 1311
rect 1855 1311 1856 1312
rect 1860 1311 1861 1315
rect 1855 1310 1861 1311
rect 1910 1315 1916 1316
rect 1910 1311 1911 1315
rect 1915 1314 1916 1315
rect 1919 1315 1925 1316
rect 1919 1314 1920 1315
rect 1915 1312 1920 1314
rect 1915 1311 1916 1312
rect 1910 1310 1916 1311
rect 1919 1311 1920 1312
rect 1924 1311 1925 1315
rect 1919 1310 1925 1311
rect 1974 1315 1980 1316
rect 1974 1311 1975 1315
rect 1979 1314 1980 1315
rect 1983 1315 1989 1316
rect 1983 1314 1984 1315
rect 1979 1312 1984 1314
rect 1979 1311 1980 1312
rect 1974 1310 1980 1311
rect 1983 1311 1984 1312
rect 1988 1311 1989 1315
rect 1983 1310 1989 1311
rect 2038 1315 2044 1316
rect 2038 1311 2039 1315
rect 2043 1314 2044 1315
rect 2047 1315 2053 1316
rect 2047 1314 2048 1315
rect 2043 1312 2048 1314
rect 2043 1311 2044 1312
rect 2038 1310 2044 1311
rect 2047 1311 2048 1312
rect 2052 1311 2053 1315
rect 2047 1310 2053 1311
rect 2094 1315 2101 1316
rect 2118 1315 2124 1316
rect 2094 1311 2095 1315
rect 2100 1311 2101 1315
rect 2094 1310 2101 1311
rect 244 1304 274 1306
rect 278 1307 285 1308
rect 244 1303 245 1304
rect 239 1302 245 1303
rect 278 1303 279 1307
rect 284 1303 285 1307
rect 278 1302 285 1303
rect 287 1307 293 1308
rect 287 1303 288 1307
rect 292 1306 293 1307
rect 343 1307 349 1308
rect 343 1306 344 1307
rect 292 1304 344 1306
rect 292 1303 293 1304
rect 287 1302 293 1303
rect 343 1303 344 1304
rect 348 1303 349 1307
rect 343 1302 349 1303
rect 358 1307 364 1308
rect 358 1303 359 1307
rect 363 1306 364 1307
rect 415 1307 421 1308
rect 415 1306 416 1307
rect 363 1304 416 1306
rect 363 1303 364 1304
rect 358 1302 364 1303
rect 415 1303 416 1304
rect 420 1303 421 1307
rect 415 1302 421 1303
rect 423 1307 429 1308
rect 423 1303 424 1307
rect 428 1306 429 1307
rect 487 1307 493 1308
rect 487 1306 488 1307
rect 428 1304 488 1306
rect 428 1303 429 1304
rect 423 1302 429 1303
rect 487 1303 488 1304
rect 492 1303 493 1307
rect 487 1302 493 1303
rect 567 1307 573 1308
rect 567 1303 568 1307
rect 572 1306 573 1307
rect 638 1307 644 1308
rect 638 1306 639 1307
rect 572 1304 639 1306
rect 572 1303 573 1304
rect 567 1302 573 1303
rect 638 1303 639 1304
rect 643 1303 644 1307
rect 638 1302 644 1303
rect 647 1307 653 1308
rect 647 1303 648 1307
rect 652 1306 653 1307
rect 718 1307 724 1308
rect 718 1306 719 1307
rect 652 1304 719 1306
rect 652 1303 653 1304
rect 647 1302 653 1303
rect 718 1303 719 1304
rect 723 1303 724 1307
rect 718 1302 724 1303
rect 727 1307 736 1308
rect 727 1303 728 1307
rect 735 1303 736 1307
rect 727 1302 736 1303
rect 806 1307 813 1308
rect 806 1303 807 1307
rect 812 1303 813 1307
rect 806 1302 813 1303
rect 815 1307 821 1308
rect 815 1303 816 1307
rect 820 1306 821 1307
rect 887 1307 893 1308
rect 887 1306 888 1307
rect 820 1304 888 1306
rect 820 1303 821 1304
rect 815 1302 821 1303
rect 887 1303 888 1304
rect 892 1303 893 1307
rect 887 1302 893 1303
rect 895 1307 901 1308
rect 895 1303 896 1307
rect 900 1306 901 1307
rect 967 1307 973 1308
rect 967 1306 968 1307
rect 900 1304 968 1306
rect 900 1303 901 1304
rect 895 1302 901 1303
rect 967 1303 968 1304
rect 972 1303 973 1307
rect 967 1302 973 1303
rect 975 1307 981 1308
rect 975 1303 976 1307
rect 980 1306 981 1307
rect 1047 1307 1053 1308
rect 1047 1306 1048 1307
rect 980 1304 1048 1306
rect 980 1303 981 1304
rect 975 1302 981 1303
rect 1047 1303 1048 1304
rect 1052 1303 1053 1307
rect 1047 1302 1053 1303
rect 1094 1304 1100 1305
rect 110 1299 116 1300
rect 1094 1300 1095 1304
rect 1099 1300 1100 1304
rect 1094 1299 1100 1300
rect 1134 1303 1140 1304
rect 1134 1299 1135 1303
rect 1139 1299 1140 1303
rect 2118 1303 2124 1304
rect 1134 1298 1140 1299
rect 1158 1300 1164 1301
rect 134 1296 140 1297
rect 134 1292 135 1296
rect 139 1292 140 1296
rect 134 1291 140 1292
rect 174 1296 180 1297
rect 174 1292 175 1296
rect 179 1292 180 1296
rect 174 1291 180 1292
rect 214 1296 220 1297
rect 214 1292 215 1296
rect 219 1292 220 1296
rect 214 1291 220 1292
rect 254 1296 260 1297
rect 254 1292 255 1296
rect 259 1292 260 1296
rect 254 1291 260 1292
rect 318 1296 324 1297
rect 318 1292 319 1296
rect 323 1292 324 1296
rect 318 1291 324 1292
rect 390 1296 396 1297
rect 390 1292 391 1296
rect 395 1292 396 1296
rect 390 1291 396 1292
rect 462 1296 468 1297
rect 462 1292 463 1296
rect 467 1292 468 1296
rect 462 1291 468 1292
rect 542 1296 548 1297
rect 542 1292 543 1296
rect 547 1292 548 1296
rect 542 1291 548 1292
rect 622 1296 628 1297
rect 622 1292 623 1296
rect 627 1292 628 1296
rect 622 1291 628 1292
rect 702 1296 708 1297
rect 702 1292 703 1296
rect 707 1292 708 1296
rect 702 1291 708 1292
rect 782 1296 788 1297
rect 782 1292 783 1296
rect 787 1292 788 1296
rect 782 1291 788 1292
rect 862 1296 868 1297
rect 862 1292 863 1296
rect 867 1292 868 1296
rect 862 1291 868 1292
rect 942 1296 948 1297
rect 942 1292 943 1296
rect 947 1292 948 1296
rect 942 1291 948 1292
rect 1022 1296 1028 1297
rect 1022 1292 1023 1296
rect 1027 1292 1028 1296
rect 1158 1296 1159 1300
rect 1163 1296 1164 1300
rect 1158 1295 1164 1296
rect 1222 1300 1228 1301
rect 1222 1296 1223 1300
rect 1227 1296 1228 1300
rect 1222 1295 1228 1296
rect 1310 1300 1316 1301
rect 1310 1296 1311 1300
rect 1315 1296 1316 1300
rect 1310 1295 1316 1296
rect 1406 1300 1412 1301
rect 1406 1296 1407 1300
rect 1411 1296 1412 1300
rect 1406 1295 1412 1296
rect 1502 1300 1508 1301
rect 1502 1296 1503 1300
rect 1507 1296 1508 1300
rect 1502 1295 1508 1296
rect 1598 1300 1604 1301
rect 1598 1296 1599 1300
rect 1603 1296 1604 1300
rect 1598 1295 1604 1296
rect 1678 1300 1684 1301
rect 1678 1296 1679 1300
rect 1683 1296 1684 1300
rect 1678 1295 1684 1296
rect 1758 1300 1764 1301
rect 1758 1296 1759 1300
rect 1763 1296 1764 1300
rect 1758 1295 1764 1296
rect 1830 1300 1836 1301
rect 1830 1296 1831 1300
rect 1835 1296 1836 1300
rect 1830 1295 1836 1296
rect 1894 1300 1900 1301
rect 1894 1296 1895 1300
rect 1899 1296 1900 1300
rect 1894 1295 1900 1296
rect 1958 1300 1964 1301
rect 1958 1296 1959 1300
rect 1963 1296 1964 1300
rect 1958 1295 1964 1296
rect 2022 1300 2028 1301
rect 2022 1296 2023 1300
rect 2027 1296 2028 1300
rect 2022 1295 2028 1296
rect 2070 1300 2076 1301
rect 2070 1296 2071 1300
rect 2075 1296 2076 1300
rect 2118 1299 2119 1303
rect 2123 1299 2124 1303
rect 2118 1298 2124 1299
rect 2070 1295 2076 1296
rect 1022 1291 1028 1292
rect 1174 1288 1180 1289
rect 158 1287 165 1288
rect 158 1283 159 1287
rect 164 1283 165 1287
rect 158 1282 165 1283
rect 190 1287 196 1288
rect 190 1283 191 1287
rect 195 1286 196 1287
rect 199 1287 205 1288
rect 199 1286 200 1287
rect 195 1284 200 1286
rect 195 1283 196 1284
rect 190 1282 196 1283
rect 199 1283 200 1284
rect 204 1283 205 1287
rect 199 1282 205 1283
rect 230 1287 236 1288
rect 230 1283 231 1287
rect 235 1286 236 1287
rect 239 1287 245 1288
rect 239 1286 240 1287
rect 235 1284 240 1286
rect 235 1283 236 1284
rect 230 1282 236 1283
rect 239 1283 240 1284
rect 244 1283 245 1287
rect 239 1282 245 1283
rect 279 1287 285 1288
rect 279 1283 280 1287
rect 284 1286 285 1287
rect 287 1287 293 1288
rect 287 1286 288 1287
rect 284 1284 288 1286
rect 284 1283 285 1284
rect 279 1282 285 1283
rect 287 1283 288 1284
rect 292 1283 293 1287
rect 287 1282 293 1283
rect 342 1287 349 1288
rect 342 1283 343 1287
rect 348 1283 349 1287
rect 342 1282 349 1283
rect 415 1287 421 1288
rect 415 1283 416 1287
rect 420 1286 421 1287
rect 423 1287 429 1288
rect 423 1286 424 1287
rect 420 1284 424 1286
rect 420 1283 421 1284
rect 415 1282 421 1283
rect 423 1283 424 1284
rect 428 1283 429 1287
rect 487 1287 493 1288
rect 487 1286 488 1287
rect 423 1282 429 1283
rect 432 1284 488 1286
rect 374 1279 380 1280
rect 374 1275 375 1279
rect 379 1278 380 1279
rect 432 1278 434 1284
rect 487 1283 488 1284
rect 492 1283 493 1287
rect 487 1282 493 1283
rect 550 1287 556 1288
rect 550 1283 551 1287
rect 555 1286 556 1287
rect 567 1287 573 1288
rect 567 1286 568 1287
rect 555 1284 568 1286
rect 555 1283 556 1284
rect 550 1282 556 1283
rect 567 1283 568 1284
rect 572 1283 573 1287
rect 567 1282 573 1283
rect 638 1287 644 1288
rect 638 1283 639 1287
rect 643 1286 644 1287
rect 647 1287 653 1288
rect 647 1286 648 1287
rect 643 1284 648 1286
rect 643 1283 644 1284
rect 638 1282 644 1283
rect 647 1283 648 1284
rect 652 1283 653 1287
rect 647 1282 653 1283
rect 718 1287 724 1288
rect 718 1283 719 1287
rect 723 1286 724 1287
rect 727 1287 733 1288
rect 727 1286 728 1287
rect 723 1284 728 1286
rect 723 1283 724 1284
rect 718 1282 724 1283
rect 727 1283 728 1284
rect 732 1283 733 1287
rect 727 1282 733 1283
rect 807 1287 813 1288
rect 807 1283 808 1287
rect 812 1286 813 1287
rect 815 1287 821 1288
rect 815 1286 816 1287
rect 812 1284 816 1286
rect 812 1283 813 1284
rect 807 1282 813 1283
rect 815 1283 816 1284
rect 820 1283 821 1287
rect 815 1282 821 1283
rect 887 1287 893 1288
rect 887 1283 888 1287
rect 892 1286 893 1287
rect 895 1287 901 1288
rect 895 1286 896 1287
rect 892 1284 896 1286
rect 892 1283 893 1284
rect 887 1282 893 1283
rect 895 1283 896 1284
rect 900 1283 901 1287
rect 895 1282 901 1283
rect 967 1287 973 1288
rect 967 1283 968 1287
rect 972 1286 973 1287
rect 975 1287 981 1288
rect 975 1286 976 1287
rect 972 1284 976 1286
rect 972 1283 973 1284
rect 967 1282 973 1283
rect 975 1283 976 1284
rect 980 1283 981 1287
rect 975 1282 981 1283
rect 1047 1287 1053 1288
rect 1047 1283 1048 1287
rect 1052 1286 1053 1287
rect 1070 1287 1076 1288
rect 1070 1286 1071 1287
rect 1052 1284 1071 1286
rect 1052 1283 1053 1284
rect 1047 1282 1053 1283
rect 1070 1283 1071 1284
rect 1075 1283 1076 1287
rect 1070 1282 1076 1283
rect 1134 1285 1140 1286
rect 1134 1281 1135 1285
rect 1139 1281 1140 1285
rect 1174 1284 1175 1288
rect 1179 1284 1180 1288
rect 1174 1283 1180 1284
rect 1230 1288 1236 1289
rect 1230 1284 1231 1288
rect 1235 1284 1236 1288
rect 1230 1283 1236 1284
rect 1302 1288 1308 1289
rect 1302 1284 1303 1288
rect 1307 1284 1308 1288
rect 1302 1283 1308 1284
rect 1390 1288 1396 1289
rect 1390 1284 1391 1288
rect 1395 1284 1396 1288
rect 1390 1283 1396 1284
rect 1478 1288 1484 1289
rect 1478 1284 1479 1288
rect 1483 1284 1484 1288
rect 1478 1283 1484 1284
rect 1566 1288 1572 1289
rect 1566 1284 1567 1288
rect 1571 1284 1572 1288
rect 1566 1283 1572 1284
rect 1654 1288 1660 1289
rect 1654 1284 1655 1288
rect 1659 1284 1660 1288
rect 1654 1283 1660 1284
rect 1742 1288 1748 1289
rect 1742 1284 1743 1288
rect 1747 1284 1748 1288
rect 1742 1283 1748 1284
rect 1830 1288 1836 1289
rect 1830 1284 1831 1288
rect 1835 1284 1836 1288
rect 1830 1283 1836 1284
rect 1918 1288 1924 1289
rect 1918 1284 1919 1288
rect 1923 1284 1924 1288
rect 1918 1283 1924 1284
rect 2006 1288 2012 1289
rect 2006 1284 2007 1288
rect 2011 1284 2012 1288
rect 2006 1283 2012 1284
rect 2070 1288 2076 1289
rect 2070 1284 2071 1288
rect 2075 1284 2076 1288
rect 2070 1283 2076 1284
rect 2118 1285 2124 1286
rect 1134 1280 1140 1281
rect 2118 1281 2119 1285
rect 2123 1281 2124 1285
rect 2118 1280 2124 1281
rect 379 1276 434 1278
rect 379 1275 380 1276
rect 374 1274 380 1275
rect 278 1271 284 1272
rect 278 1270 279 1271
rect 260 1268 279 1270
rect 159 1263 165 1264
rect 159 1259 160 1263
rect 164 1262 165 1263
rect 190 1263 196 1264
rect 190 1262 191 1263
rect 164 1260 191 1262
rect 164 1259 165 1260
rect 159 1258 165 1259
rect 190 1259 191 1260
rect 195 1259 196 1263
rect 190 1258 196 1259
rect 199 1263 205 1264
rect 199 1259 200 1263
rect 204 1262 205 1263
rect 230 1263 236 1264
rect 230 1262 231 1263
rect 204 1260 231 1262
rect 204 1259 205 1260
rect 199 1258 205 1259
rect 230 1259 231 1260
rect 235 1259 236 1263
rect 230 1258 236 1259
rect 239 1263 245 1264
rect 239 1259 240 1263
rect 244 1262 245 1263
rect 260 1262 262 1268
rect 278 1267 279 1268
rect 283 1267 284 1271
rect 278 1266 284 1267
rect 574 1271 580 1272
rect 574 1267 575 1271
rect 579 1270 580 1271
rect 1198 1271 1205 1272
rect 579 1268 826 1270
rect 579 1267 580 1268
rect 574 1266 580 1267
rect 824 1264 826 1268
rect 1134 1268 1140 1269
rect 1134 1264 1135 1268
rect 1139 1264 1140 1268
rect 1198 1267 1199 1271
rect 1204 1267 1205 1271
rect 1198 1266 1205 1267
rect 1207 1271 1213 1272
rect 1207 1267 1208 1271
rect 1212 1270 1213 1271
rect 1255 1271 1261 1272
rect 1255 1270 1256 1271
rect 1212 1268 1256 1270
rect 1212 1267 1213 1268
rect 1207 1266 1213 1267
rect 1255 1267 1256 1268
rect 1260 1267 1261 1271
rect 1255 1266 1261 1267
rect 1263 1271 1269 1272
rect 1263 1267 1264 1271
rect 1268 1270 1269 1271
rect 1327 1271 1333 1272
rect 1327 1270 1328 1271
rect 1268 1268 1328 1270
rect 1268 1267 1269 1268
rect 1263 1266 1269 1267
rect 1327 1267 1328 1268
rect 1332 1267 1333 1271
rect 1327 1266 1333 1267
rect 1410 1271 1421 1272
rect 1410 1267 1411 1271
rect 1415 1267 1416 1271
rect 1420 1267 1421 1271
rect 1410 1266 1421 1267
rect 1423 1271 1429 1272
rect 1423 1267 1424 1271
rect 1428 1270 1429 1271
rect 1503 1271 1509 1272
rect 1503 1270 1504 1271
rect 1428 1268 1504 1270
rect 1428 1267 1429 1268
rect 1423 1266 1429 1267
rect 1503 1267 1504 1268
rect 1508 1267 1509 1271
rect 1503 1266 1509 1267
rect 1511 1271 1517 1272
rect 1511 1267 1512 1271
rect 1516 1270 1517 1271
rect 1591 1271 1597 1272
rect 1591 1270 1592 1271
rect 1516 1268 1592 1270
rect 1516 1267 1517 1268
rect 1511 1266 1517 1267
rect 1591 1267 1592 1268
rect 1596 1267 1597 1271
rect 1591 1266 1597 1267
rect 1670 1271 1676 1272
rect 1670 1267 1671 1271
rect 1675 1270 1676 1271
rect 1679 1271 1685 1272
rect 1679 1270 1680 1271
rect 1675 1268 1680 1270
rect 1675 1267 1676 1268
rect 1670 1266 1676 1267
rect 1679 1267 1680 1268
rect 1684 1267 1685 1271
rect 1679 1266 1685 1267
rect 1687 1271 1693 1272
rect 1687 1267 1688 1271
rect 1692 1270 1693 1271
rect 1767 1271 1773 1272
rect 1767 1270 1768 1271
rect 1692 1268 1768 1270
rect 1692 1267 1693 1268
rect 1687 1266 1693 1267
rect 1767 1267 1768 1268
rect 1772 1267 1773 1271
rect 1767 1266 1773 1267
rect 1775 1271 1781 1272
rect 1775 1267 1776 1271
rect 1780 1270 1781 1271
rect 1855 1271 1861 1272
rect 1855 1270 1856 1271
rect 1780 1268 1856 1270
rect 1780 1267 1781 1268
rect 1775 1266 1781 1267
rect 1855 1267 1856 1268
rect 1860 1267 1861 1271
rect 1855 1266 1861 1267
rect 1863 1271 1869 1272
rect 1863 1267 1864 1271
rect 1868 1270 1869 1271
rect 1943 1271 1949 1272
rect 1943 1270 1944 1271
rect 1868 1268 1944 1270
rect 1868 1267 1869 1268
rect 1863 1266 1869 1267
rect 1943 1267 1944 1268
rect 1948 1267 1949 1271
rect 1943 1266 1949 1267
rect 2031 1271 2037 1272
rect 2031 1267 2032 1271
rect 2036 1270 2037 1271
rect 2046 1271 2052 1272
rect 2046 1270 2047 1271
rect 2036 1268 2047 1270
rect 2036 1267 2037 1268
rect 2031 1266 2037 1267
rect 2046 1267 2047 1268
rect 2051 1267 2052 1271
rect 2046 1266 2052 1267
rect 2095 1271 2101 1272
rect 2095 1267 2096 1271
rect 2100 1270 2101 1271
rect 2103 1271 2109 1272
rect 2103 1270 2104 1271
rect 2100 1268 2104 1270
rect 2100 1267 2101 1268
rect 2095 1266 2101 1267
rect 2103 1267 2104 1268
rect 2108 1267 2109 1271
rect 2103 1266 2109 1267
rect 2118 1268 2124 1269
rect 279 1263 285 1264
rect 279 1262 280 1263
rect 244 1260 262 1262
rect 264 1260 280 1262
rect 244 1259 245 1260
rect 239 1258 245 1259
rect 134 1256 140 1257
rect 134 1252 135 1256
rect 139 1252 140 1256
rect 134 1251 140 1252
rect 174 1256 180 1257
rect 174 1252 175 1256
rect 179 1252 180 1256
rect 174 1251 180 1252
rect 214 1256 220 1257
rect 214 1252 215 1256
rect 219 1252 220 1256
rect 214 1251 220 1252
rect 254 1256 260 1257
rect 254 1252 255 1256
rect 259 1252 260 1256
rect 254 1251 260 1252
rect 110 1248 116 1249
rect 110 1244 111 1248
rect 115 1244 116 1248
rect 184 1248 210 1250
rect 110 1243 116 1244
rect 159 1243 165 1244
rect 159 1239 160 1243
rect 164 1242 165 1243
rect 184 1242 186 1248
rect 208 1246 210 1248
rect 224 1248 250 1250
rect 224 1246 226 1248
rect 208 1244 226 1246
rect 248 1246 250 1248
rect 264 1246 266 1260
rect 279 1259 280 1260
rect 284 1259 285 1263
rect 279 1258 285 1259
rect 287 1263 293 1264
rect 287 1259 288 1263
rect 292 1262 293 1263
rect 343 1263 349 1264
rect 343 1262 344 1263
rect 292 1260 344 1262
rect 292 1259 293 1260
rect 287 1258 293 1259
rect 343 1259 344 1260
rect 348 1259 349 1263
rect 343 1258 349 1259
rect 351 1263 357 1264
rect 351 1259 352 1263
rect 356 1262 357 1263
rect 423 1263 429 1264
rect 423 1262 424 1263
rect 356 1260 424 1262
rect 356 1259 357 1260
rect 351 1258 357 1259
rect 423 1259 424 1260
rect 428 1259 429 1263
rect 423 1258 429 1259
rect 511 1263 517 1264
rect 511 1259 512 1263
rect 516 1262 517 1263
rect 598 1263 604 1264
rect 598 1262 599 1263
rect 516 1260 599 1262
rect 516 1259 517 1260
rect 511 1258 517 1259
rect 598 1259 599 1260
rect 603 1259 604 1263
rect 598 1258 604 1259
rect 607 1263 613 1264
rect 607 1259 608 1263
rect 612 1262 613 1263
rect 702 1263 708 1264
rect 702 1262 703 1263
rect 612 1260 703 1262
rect 612 1259 613 1260
rect 607 1258 613 1259
rect 702 1259 703 1260
rect 707 1259 708 1263
rect 702 1258 708 1259
rect 711 1263 717 1264
rect 711 1259 712 1263
rect 716 1262 717 1263
rect 814 1263 820 1264
rect 814 1262 815 1263
rect 716 1260 815 1262
rect 716 1259 717 1260
rect 711 1258 717 1259
rect 814 1259 815 1260
rect 819 1259 820 1263
rect 814 1258 820 1259
rect 823 1263 829 1264
rect 823 1259 824 1263
rect 828 1259 829 1263
rect 823 1258 829 1259
rect 943 1263 949 1264
rect 943 1259 944 1263
rect 948 1262 949 1263
rect 1006 1263 1012 1264
rect 1006 1262 1007 1263
rect 948 1260 1007 1262
rect 948 1259 949 1260
rect 943 1258 949 1259
rect 1006 1259 1007 1260
rect 1011 1259 1012 1263
rect 1006 1258 1012 1259
rect 1014 1263 1020 1264
rect 1014 1259 1015 1263
rect 1019 1262 1020 1263
rect 1071 1263 1077 1264
rect 1134 1263 1140 1264
rect 2118 1264 2119 1268
rect 2123 1264 2124 1268
rect 2118 1263 2124 1264
rect 1071 1262 1072 1263
rect 1019 1260 1072 1262
rect 1019 1259 1020 1260
rect 1014 1258 1020 1259
rect 1071 1259 1072 1260
rect 1076 1259 1077 1263
rect 1071 1258 1077 1259
rect 1174 1260 1180 1261
rect 318 1256 324 1257
rect 318 1252 319 1256
rect 323 1252 324 1256
rect 318 1251 324 1252
rect 398 1256 404 1257
rect 398 1252 399 1256
rect 403 1252 404 1256
rect 398 1251 404 1252
rect 486 1256 492 1257
rect 486 1252 487 1256
rect 491 1252 492 1256
rect 486 1251 492 1252
rect 582 1256 588 1257
rect 582 1252 583 1256
rect 587 1252 588 1256
rect 582 1251 588 1252
rect 686 1256 692 1257
rect 686 1252 687 1256
rect 691 1252 692 1256
rect 686 1251 692 1252
rect 798 1256 804 1257
rect 798 1252 799 1256
rect 803 1252 804 1256
rect 798 1251 804 1252
rect 918 1256 924 1257
rect 918 1252 919 1256
rect 923 1252 924 1256
rect 918 1251 924 1252
rect 1046 1256 1052 1257
rect 1046 1252 1047 1256
rect 1051 1252 1052 1256
rect 1174 1256 1175 1260
rect 1179 1256 1180 1260
rect 1174 1255 1180 1256
rect 1230 1260 1236 1261
rect 1230 1256 1231 1260
rect 1235 1256 1236 1260
rect 1230 1255 1236 1256
rect 1302 1260 1308 1261
rect 1302 1256 1303 1260
rect 1307 1256 1308 1260
rect 1302 1255 1308 1256
rect 1390 1260 1396 1261
rect 1390 1256 1391 1260
rect 1395 1256 1396 1260
rect 1390 1255 1396 1256
rect 1478 1260 1484 1261
rect 1478 1256 1479 1260
rect 1483 1256 1484 1260
rect 1478 1255 1484 1256
rect 1566 1260 1572 1261
rect 1566 1256 1567 1260
rect 1571 1256 1572 1260
rect 1566 1255 1572 1256
rect 1654 1260 1660 1261
rect 1654 1256 1655 1260
rect 1659 1256 1660 1260
rect 1654 1255 1660 1256
rect 1742 1260 1748 1261
rect 1742 1256 1743 1260
rect 1747 1256 1748 1260
rect 1742 1255 1748 1256
rect 1830 1260 1836 1261
rect 1830 1256 1831 1260
rect 1835 1256 1836 1260
rect 1830 1255 1836 1256
rect 1918 1260 1924 1261
rect 1918 1256 1919 1260
rect 1923 1256 1924 1260
rect 1918 1255 1924 1256
rect 2006 1260 2012 1261
rect 2006 1256 2007 1260
rect 2011 1256 2012 1260
rect 2006 1255 2012 1256
rect 2070 1260 2076 1261
rect 2070 1256 2071 1260
rect 2075 1256 2076 1260
rect 2070 1255 2076 1256
rect 1046 1251 1052 1252
rect 1199 1251 1205 1252
rect 248 1244 266 1246
rect 1094 1248 1100 1249
rect 1094 1244 1095 1248
rect 1099 1244 1100 1248
rect 1199 1247 1200 1251
rect 1204 1250 1205 1251
rect 1207 1251 1213 1252
rect 1207 1250 1208 1251
rect 1204 1248 1208 1250
rect 1204 1247 1205 1248
rect 1199 1246 1205 1247
rect 1207 1247 1208 1248
rect 1212 1247 1213 1251
rect 1207 1246 1213 1247
rect 1255 1251 1261 1252
rect 1255 1247 1256 1251
rect 1260 1250 1261 1251
rect 1263 1251 1269 1252
rect 1263 1250 1264 1251
rect 1260 1248 1264 1250
rect 1260 1247 1261 1248
rect 1255 1246 1261 1247
rect 1263 1247 1264 1248
rect 1268 1247 1269 1251
rect 1263 1246 1269 1247
rect 1327 1251 1336 1252
rect 1327 1247 1328 1251
rect 1335 1247 1336 1251
rect 1327 1246 1336 1247
rect 1415 1251 1421 1252
rect 1415 1247 1416 1251
rect 1420 1250 1421 1251
rect 1423 1251 1429 1252
rect 1423 1250 1424 1251
rect 1420 1248 1424 1250
rect 1420 1247 1421 1248
rect 1415 1246 1421 1247
rect 1423 1247 1424 1248
rect 1428 1247 1429 1251
rect 1423 1246 1429 1247
rect 1503 1251 1509 1252
rect 1503 1247 1504 1251
rect 1508 1250 1509 1251
rect 1511 1251 1517 1252
rect 1511 1250 1512 1251
rect 1508 1248 1512 1250
rect 1508 1247 1509 1248
rect 1503 1246 1509 1247
rect 1511 1247 1512 1248
rect 1516 1247 1517 1251
rect 1511 1246 1517 1247
rect 1590 1251 1597 1252
rect 1590 1247 1591 1251
rect 1596 1247 1597 1251
rect 1590 1246 1597 1247
rect 1679 1251 1685 1252
rect 1679 1247 1680 1251
rect 1684 1250 1685 1251
rect 1687 1251 1693 1252
rect 1687 1250 1688 1251
rect 1684 1248 1688 1250
rect 1684 1247 1685 1248
rect 1679 1246 1685 1247
rect 1687 1247 1688 1248
rect 1692 1247 1693 1251
rect 1687 1246 1693 1247
rect 1767 1251 1773 1252
rect 1767 1247 1768 1251
rect 1772 1250 1773 1251
rect 1775 1251 1781 1252
rect 1775 1250 1776 1251
rect 1772 1248 1776 1250
rect 1772 1247 1773 1248
rect 1767 1246 1773 1247
rect 1775 1247 1776 1248
rect 1780 1247 1781 1251
rect 1775 1246 1781 1247
rect 1855 1251 1861 1252
rect 1855 1247 1856 1251
rect 1860 1250 1861 1251
rect 1863 1251 1869 1252
rect 1863 1250 1864 1251
rect 1860 1248 1864 1250
rect 1860 1247 1861 1248
rect 1855 1246 1861 1247
rect 1863 1247 1864 1248
rect 1868 1247 1869 1251
rect 1863 1246 1869 1247
rect 1943 1251 1949 1252
rect 1943 1247 1944 1251
rect 1948 1247 1949 1251
rect 1943 1246 1949 1247
rect 1994 1251 2000 1252
rect 1994 1247 1995 1251
rect 1999 1250 2000 1251
rect 2031 1251 2037 1252
rect 2031 1250 2032 1251
rect 1999 1248 2032 1250
rect 1999 1247 2000 1248
rect 1994 1246 2000 1247
rect 2031 1247 2032 1248
rect 2036 1247 2037 1251
rect 2031 1246 2037 1247
rect 2094 1251 2101 1252
rect 2094 1247 2095 1251
rect 2100 1247 2101 1251
rect 2094 1246 2101 1247
rect 164 1240 186 1242
rect 190 1243 196 1244
rect 164 1239 165 1240
rect 159 1238 165 1239
rect 190 1239 191 1243
rect 195 1242 196 1243
rect 199 1243 205 1244
rect 199 1242 200 1243
rect 195 1240 200 1242
rect 195 1239 196 1240
rect 190 1238 196 1239
rect 199 1239 200 1240
rect 204 1239 205 1243
rect 199 1238 205 1239
rect 230 1243 236 1244
rect 230 1239 231 1243
rect 235 1242 236 1243
rect 239 1243 245 1244
rect 239 1242 240 1243
rect 235 1240 240 1242
rect 235 1239 236 1240
rect 230 1238 236 1239
rect 239 1239 240 1240
rect 244 1239 245 1243
rect 239 1238 245 1239
rect 279 1243 285 1244
rect 279 1239 280 1243
rect 284 1242 285 1243
rect 287 1243 293 1244
rect 287 1242 288 1243
rect 284 1240 288 1242
rect 284 1239 285 1240
rect 279 1238 285 1239
rect 287 1239 288 1240
rect 292 1239 293 1243
rect 287 1238 293 1239
rect 343 1243 349 1244
rect 343 1239 344 1243
rect 348 1242 349 1243
rect 351 1243 357 1244
rect 351 1242 352 1243
rect 348 1240 352 1242
rect 348 1239 349 1240
rect 343 1238 349 1239
rect 351 1239 352 1240
rect 356 1239 357 1243
rect 351 1238 357 1239
rect 378 1243 384 1244
rect 378 1239 379 1243
rect 383 1242 384 1243
rect 423 1243 429 1244
rect 423 1242 424 1243
rect 383 1240 424 1242
rect 383 1239 384 1240
rect 378 1238 384 1239
rect 423 1239 424 1240
rect 428 1239 429 1243
rect 423 1238 429 1239
rect 511 1243 517 1244
rect 511 1239 512 1243
rect 516 1242 517 1243
rect 550 1243 556 1244
rect 550 1242 551 1243
rect 516 1240 551 1242
rect 516 1239 517 1240
rect 511 1238 517 1239
rect 550 1239 551 1240
rect 555 1239 556 1243
rect 550 1238 556 1239
rect 598 1243 604 1244
rect 598 1239 599 1243
rect 603 1242 604 1243
rect 607 1243 613 1244
rect 607 1242 608 1243
rect 603 1240 608 1242
rect 603 1239 604 1240
rect 598 1238 604 1239
rect 607 1239 608 1240
rect 612 1239 613 1243
rect 607 1238 613 1239
rect 702 1243 708 1244
rect 702 1239 703 1243
rect 707 1242 708 1243
rect 711 1243 717 1244
rect 711 1242 712 1243
rect 707 1240 712 1242
rect 707 1239 708 1240
rect 702 1238 708 1239
rect 711 1239 712 1240
rect 716 1239 717 1243
rect 711 1238 717 1239
rect 814 1243 820 1244
rect 814 1239 815 1243
rect 819 1242 820 1243
rect 823 1243 829 1244
rect 823 1242 824 1243
rect 819 1240 824 1242
rect 819 1239 820 1240
rect 814 1238 820 1239
rect 823 1239 824 1240
rect 828 1239 829 1243
rect 823 1238 829 1239
rect 943 1243 949 1244
rect 943 1239 944 1243
rect 948 1242 949 1243
rect 1014 1243 1020 1244
rect 1014 1242 1015 1243
rect 948 1240 1015 1242
rect 948 1239 949 1240
rect 943 1238 949 1239
rect 1014 1239 1015 1240
rect 1019 1239 1020 1243
rect 1014 1238 1020 1239
rect 1070 1243 1077 1244
rect 1094 1243 1100 1244
rect 1766 1243 1772 1244
rect 1070 1239 1071 1243
rect 1076 1239 1077 1243
rect 1070 1238 1077 1239
rect 1766 1239 1767 1243
rect 1771 1242 1772 1243
rect 1945 1242 1947 1246
rect 1771 1240 1947 1242
rect 1771 1239 1772 1240
rect 1766 1238 1772 1239
rect 1314 1235 1320 1236
rect 110 1231 116 1232
rect 110 1227 111 1231
rect 115 1227 116 1231
rect 1094 1231 1100 1232
rect 110 1226 116 1227
rect 134 1228 140 1229
rect 134 1224 135 1228
rect 139 1224 140 1228
rect 134 1223 140 1224
rect 174 1228 180 1229
rect 174 1224 175 1228
rect 179 1224 180 1228
rect 174 1223 180 1224
rect 214 1228 220 1229
rect 214 1224 215 1228
rect 219 1224 220 1228
rect 214 1223 220 1224
rect 254 1228 260 1229
rect 254 1224 255 1228
rect 259 1224 260 1228
rect 254 1223 260 1224
rect 318 1228 324 1229
rect 318 1224 319 1228
rect 323 1224 324 1228
rect 318 1223 324 1224
rect 398 1228 404 1229
rect 398 1224 399 1228
rect 403 1224 404 1228
rect 398 1223 404 1224
rect 486 1228 492 1229
rect 486 1224 487 1228
rect 491 1224 492 1228
rect 486 1223 492 1224
rect 582 1228 588 1229
rect 582 1224 583 1228
rect 587 1224 588 1228
rect 582 1223 588 1224
rect 686 1228 692 1229
rect 686 1224 687 1228
rect 691 1224 692 1228
rect 686 1223 692 1224
rect 798 1228 804 1229
rect 798 1224 799 1228
rect 803 1224 804 1228
rect 798 1223 804 1224
rect 918 1228 924 1229
rect 918 1224 919 1228
rect 923 1224 924 1228
rect 918 1223 924 1224
rect 1046 1228 1052 1229
rect 1046 1224 1047 1228
rect 1051 1224 1052 1228
rect 1094 1227 1095 1231
rect 1099 1227 1100 1231
rect 1314 1231 1315 1235
rect 1319 1234 1320 1235
rect 1458 1235 1464 1236
rect 1319 1232 1422 1234
rect 1319 1231 1320 1232
rect 1314 1230 1320 1231
rect 1094 1226 1100 1227
rect 1311 1227 1317 1228
rect 1046 1223 1052 1224
rect 1311 1223 1312 1227
rect 1316 1226 1317 1227
rect 1342 1227 1348 1228
rect 1342 1226 1343 1227
rect 1316 1224 1343 1226
rect 1316 1223 1317 1224
rect 1311 1222 1317 1223
rect 1342 1223 1343 1224
rect 1347 1223 1348 1227
rect 1342 1222 1348 1223
rect 1351 1227 1357 1228
rect 1351 1223 1352 1227
rect 1356 1226 1357 1227
rect 1390 1227 1396 1228
rect 1390 1226 1391 1227
rect 1356 1224 1391 1226
rect 1356 1223 1357 1224
rect 1351 1222 1357 1223
rect 1390 1223 1391 1224
rect 1395 1223 1396 1227
rect 1390 1222 1396 1223
rect 1399 1227 1405 1228
rect 1399 1223 1400 1227
rect 1404 1226 1405 1227
rect 1410 1227 1416 1228
rect 1410 1226 1411 1227
rect 1404 1224 1411 1226
rect 1404 1223 1405 1224
rect 1399 1222 1405 1223
rect 1410 1223 1411 1224
rect 1415 1223 1416 1227
rect 1420 1226 1422 1232
rect 1458 1231 1459 1235
rect 1463 1234 1464 1235
rect 1670 1235 1676 1236
rect 1463 1232 1587 1234
rect 1463 1231 1464 1232
rect 1458 1230 1464 1231
rect 1585 1228 1587 1232
rect 1670 1231 1671 1235
rect 1675 1234 1676 1235
rect 1675 1232 1930 1234
rect 1675 1231 1676 1232
rect 1670 1230 1676 1231
rect 1928 1228 1930 1232
rect 1455 1227 1461 1228
rect 1455 1226 1456 1227
rect 1420 1224 1456 1226
rect 1410 1222 1416 1223
rect 1455 1223 1456 1224
rect 1460 1223 1461 1227
rect 1455 1222 1461 1223
rect 1519 1227 1525 1228
rect 1519 1223 1520 1227
rect 1524 1226 1525 1227
rect 1574 1227 1580 1228
rect 1574 1226 1575 1227
rect 1524 1224 1575 1226
rect 1524 1223 1525 1224
rect 1519 1222 1525 1223
rect 1574 1223 1575 1224
rect 1579 1223 1580 1227
rect 1574 1222 1580 1223
rect 1583 1227 1589 1228
rect 1583 1223 1584 1227
rect 1588 1223 1589 1227
rect 1583 1222 1589 1223
rect 1647 1227 1653 1228
rect 1647 1223 1648 1227
rect 1652 1226 1653 1227
rect 1686 1227 1692 1228
rect 1686 1226 1687 1227
rect 1652 1224 1687 1226
rect 1652 1223 1653 1224
rect 1647 1222 1653 1223
rect 1686 1223 1687 1224
rect 1691 1223 1692 1227
rect 1686 1222 1692 1223
rect 1703 1227 1709 1228
rect 1703 1223 1704 1227
rect 1708 1226 1709 1227
rect 1750 1227 1756 1228
rect 1750 1226 1751 1227
rect 1708 1224 1751 1226
rect 1708 1223 1709 1224
rect 1703 1222 1709 1223
rect 1750 1223 1751 1224
rect 1755 1223 1756 1227
rect 1750 1222 1756 1223
rect 1759 1227 1765 1228
rect 1759 1223 1760 1227
rect 1764 1226 1765 1227
rect 1806 1227 1812 1228
rect 1806 1226 1807 1227
rect 1764 1224 1807 1226
rect 1764 1223 1765 1224
rect 1759 1222 1765 1223
rect 1806 1223 1807 1224
rect 1811 1223 1812 1227
rect 1806 1222 1812 1223
rect 1815 1227 1821 1228
rect 1815 1223 1816 1227
rect 1820 1226 1821 1227
rect 1854 1227 1860 1228
rect 1854 1226 1855 1227
rect 1820 1224 1855 1226
rect 1820 1223 1821 1224
rect 1815 1222 1821 1223
rect 1854 1223 1855 1224
rect 1859 1223 1860 1227
rect 1854 1222 1860 1223
rect 1871 1227 1877 1228
rect 1871 1223 1872 1227
rect 1876 1226 1877 1227
rect 1918 1227 1924 1228
rect 1918 1226 1919 1227
rect 1876 1224 1919 1226
rect 1876 1223 1877 1224
rect 1871 1222 1877 1223
rect 1918 1223 1919 1224
rect 1923 1223 1924 1227
rect 1918 1222 1924 1223
rect 1927 1227 1933 1228
rect 1927 1223 1928 1227
rect 1932 1223 1933 1227
rect 1927 1222 1933 1223
rect 1991 1227 1997 1228
rect 1991 1223 1992 1227
rect 1996 1226 1997 1227
rect 2006 1227 2012 1228
rect 2006 1226 2007 1227
rect 1996 1224 2007 1226
rect 1996 1223 1997 1224
rect 1991 1222 1997 1223
rect 2006 1223 2007 1224
rect 2011 1223 2012 1227
rect 2006 1222 2012 1223
rect 2055 1227 2061 1228
rect 2055 1223 2056 1227
rect 2060 1226 2061 1227
rect 2086 1227 2092 1228
rect 2086 1226 2087 1227
rect 2060 1224 2087 1226
rect 2060 1223 2061 1224
rect 2055 1222 2061 1223
rect 2086 1223 2087 1224
rect 2091 1223 2092 1227
rect 2086 1222 2092 1223
rect 2095 1227 2101 1228
rect 2095 1223 2096 1227
rect 2100 1226 2101 1227
rect 2103 1227 2109 1228
rect 2103 1226 2104 1227
rect 2100 1224 2104 1226
rect 2100 1223 2101 1224
rect 2095 1222 2101 1223
rect 2103 1223 2104 1224
rect 2108 1223 2109 1227
rect 2103 1222 2109 1223
rect 1286 1220 1292 1221
rect 1286 1216 1287 1220
rect 1291 1216 1292 1220
rect 1286 1215 1292 1216
rect 1326 1220 1332 1221
rect 1326 1216 1327 1220
rect 1331 1216 1332 1220
rect 1326 1215 1332 1216
rect 1374 1220 1380 1221
rect 1374 1216 1375 1220
rect 1379 1216 1380 1220
rect 1374 1215 1380 1216
rect 1430 1220 1436 1221
rect 1430 1216 1431 1220
rect 1435 1216 1436 1220
rect 1430 1215 1436 1216
rect 1494 1220 1500 1221
rect 1494 1216 1495 1220
rect 1499 1216 1500 1220
rect 1494 1215 1500 1216
rect 1558 1220 1564 1221
rect 1558 1216 1559 1220
rect 1563 1216 1564 1220
rect 1558 1215 1564 1216
rect 1622 1220 1628 1221
rect 1622 1216 1623 1220
rect 1627 1216 1628 1220
rect 1622 1215 1628 1216
rect 1678 1220 1684 1221
rect 1678 1216 1679 1220
rect 1683 1216 1684 1220
rect 1678 1215 1684 1216
rect 1734 1220 1740 1221
rect 1734 1216 1735 1220
rect 1739 1216 1740 1220
rect 1734 1215 1740 1216
rect 1790 1220 1796 1221
rect 1790 1216 1791 1220
rect 1795 1216 1796 1220
rect 1790 1215 1796 1216
rect 1846 1220 1852 1221
rect 1846 1216 1847 1220
rect 1851 1216 1852 1220
rect 1846 1215 1852 1216
rect 1902 1220 1908 1221
rect 1902 1216 1903 1220
rect 1907 1216 1908 1220
rect 1902 1215 1908 1216
rect 1966 1220 1972 1221
rect 1966 1216 1967 1220
rect 1971 1216 1972 1220
rect 1966 1215 1972 1216
rect 2030 1220 2036 1221
rect 2030 1216 2031 1220
rect 2035 1216 2036 1220
rect 2030 1215 2036 1216
rect 2070 1220 2076 1221
rect 2070 1216 2071 1220
rect 2075 1216 2076 1220
rect 2070 1215 2076 1216
rect 270 1212 276 1213
rect 110 1209 116 1210
rect 110 1205 111 1209
rect 115 1205 116 1209
rect 270 1208 271 1212
rect 275 1208 276 1212
rect 270 1207 276 1208
rect 310 1212 316 1213
rect 310 1208 311 1212
rect 315 1208 316 1212
rect 310 1207 316 1208
rect 350 1212 356 1213
rect 350 1208 351 1212
rect 355 1208 356 1212
rect 350 1207 356 1208
rect 398 1212 404 1213
rect 398 1208 399 1212
rect 403 1208 404 1212
rect 398 1207 404 1208
rect 446 1212 452 1213
rect 446 1208 447 1212
rect 451 1208 452 1212
rect 446 1207 452 1208
rect 494 1212 500 1213
rect 494 1208 495 1212
rect 499 1208 500 1212
rect 494 1207 500 1208
rect 550 1212 556 1213
rect 550 1208 551 1212
rect 555 1208 556 1212
rect 550 1207 556 1208
rect 606 1212 612 1213
rect 606 1208 607 1212
rect 611 1208 612 1212
rect 606 1207 612 1208
rect 670 1212 676 1213
rect 670 1208 671 1212
rect 675 1208 676 1212
rect 670 1207 676 1208
rect 742 1212 748 1213
rect 742 1208 743 1212
rect 747 1208 748 1212
rect 742 1207 748 1208
rect 814 1212 820 1213
rect 814 1208 815 1212
rect 819 1208 820 1212
rect 814 1207 820 1208
rect 894 1212 900 1213
rect 894 1208 895 1212
rect 899 1208 900 1212
rect 894 1207 900 1208
rect 982 1212 988 1213
rect 982 1208 983 1212
rect 987 1208 988 1212
rect 1134 1212 1140 1213
rect 982 1207 988 1208
rect 1094 1209 1100 1210
rect 110 1204 116 1205
rect 1094 1205 1095 1209
rect 1099 1205 1100 1209
rect 1134 1208 1135 1212
rect 1139 1208 1140 1212
rect 2118 1212 2124 1213
rect 2118 1208 2119 1212
rect 2123 1208 2124 1212
rect 1134 1207 1140 1208
rect 1311 1207 1320 1208
rect 1094 1204 1100 1205
rect 422 1203 428 1204
rect 422 1202 423 1203
rect 308 1200 423 1202
rect 295 1195 301 1196
rect 110 1192 116 1193
rect 110 1188 111 1192
rect 115 1188 116 1192
rect 295 1191 296 1195
rect 300 1194 301 1195
rect 308 1194 310 1200
rect 422 1199 423 1200
rect 427 1199 428 1203
rect 1311 1203 1312 1207
rect 1319 1203 1320 1207
rect 1311 1202 1320 1203
rect 1342 1207 1348 1208
rect 1342 1203 1343 1207
rect 1347 1206 1348 1207
rect 1351 1207 1357 1208
rect 1351 1206 1352 1207
rect 1347 1204 1352 1206
rect 1347 1203 1348 1204
rect 1342 1202 1348 1203
rect 1351 1203 1352 1204
rect 1356 1203 1357 1207
rect 1351 1202 1357 1203
rect 1390 1207 1396 1208
rect 1390 1203 1391 1207
rect 1395 1206 1396 1207
rect 1399 1207 1405 1208
rect 1399 1206 1400 1207
rect 1395 1204 1400 1206
rect 1395 1203 1396 1204
rect 1390 1202 1396 1203
rect 1399 1203 1400 1204
rect 1404 1203 1405 1207
rect 1399 1202 1405 1203
rect 1455 1207 1464 1208
rect 1455 1203 1456 1207
rect 1463 1203 1464 1207
rect 1455 1202 1464 1203
rect 1514 1207 1525 1208
rect 1514 1203 1515 1207
rect 1519 1203 1520 1207
rect 1524 1203 1525 1207
rect 1514 1202 1525 1203
rect 1574 1207 1580 1208
rect 1574 1203 1575 1207
rect 1579 1206 1580 1207
rect 1583 1207 1589 1208
rect 1583 1206 1584 1207
rect 1579 1204 1584 1206
rect 1579 1203 1580 1204
rect 1574 1202 1580 1203
rect 1583 1203 1584 1204
rect 1588 1203 1589 1207
rect 1583 1202 1589 1203
rect 1647 1207 1653 1208
rect 1647 1203 1648 1207
rect 1652 1206 1653 1207
rect 1670 1207 1676 1208
rect 1670 1206 1671 1207
rect 1652 1204 1671 1206
rect 1652 1203 1653 1204
rect 1647 1202 1653 1203
rect 1670 1203 1671 1204
rect 1675 1203 1676 1207
rect 1670 1202 1676 1203
rect 1686 1207 1692 1208
rect 1686 1203 1687 1207
rect 1691 1206 1692 1207
rect 1703 1207 1709 1208
rect 1703 1206 1704 1207
rect 1691 1204 1704 1206
rect 1691 1203 1692 1204
rect 1686 1202 1692 1203
rect 1703 1203 1704 1204
rect 1708 1203 1709 1207
rect 1703 1202 1709 1203
rect 1750 1207 1756 1208
rect 1750 1203 1751 1207
rect 1755 1206 1756 1207
rect 1759 1207 1765 1208
rect 1759 1206 1760 1207
rect 1755 1204 1760 1206
rect 1755 1203 1756 1204
rect 1750 1202 1756 1203
rect 1759 1203 1760 1204
rect 1764 1203 1765 1207
rect 1759 1202 1765 1203
rect 1806 1207 1812 1208
rect 1806 1203 1807 1207
rect 1811 1206 1812 1207
rect 1815 1207 1821 1208
rect 1815 1206 1816 1207
rect 1811 1204 1816 1206
rect 1811 1203 1812 1204
rect 1806 1202 1812 1203
rect 1815 1203 1816 1204
rect 1820 1203 1821 1207
rect 1815 1202 1821 1203
rect 1854 1207 1860 1208
rect 1854 1203 1855 1207
rect 1859 1206 1860 1207
rect 1871 1207 1877 1208
rect 1871 1206 1872 1207
rect 1859 1204 1872 1206
rect 1859 1203 1860 1204
rect 1854 1202 1860 1203
rect 1871 1203 1872 1204
rect 1876 1203 1877 1207
rect 1871 1202 1877 1203
rect 1918 1207 1924 1208
rect 1918 1203 1919 1207
rect 1923 1206 1924 1207
rect 1927 1207 1933 1208
rect 1927 1206 1928 1207
rect 1923 1204 1928 1206
rect 1923 1203 1924 1204
rect 1918 1202 1924 1203
rect 1927 1203 1928 1204
rect 1932 1203 1933 1207
rect 1927 1202 1933 1203
rect 1991 1207 2000 1208
rect 1991 1203 1992 1207
rect 1999 1203 2000 1207
rect 1991 1202 2000 1203
rect 2055 1207 2061 1208
rect 2055 1203 2056 1207
rect 2060 1206 2061 1207
rect 2078 1207 2084 1208
rect 2078 1206 2079 1207
rect 2060 1204 2079 1206
rect 2060 1203 2061 1204
rect 2055 1202 2061 1203
rect 2078 1203 2079 1204
rect 2083 1203 2084 1207
rect 2078 1202 2084 1203
rect 2086 1207 2092 1208
rect 2086 1203 2087 1207
rect 2091 1206 2092 1207
rect 2095 1207 2101 1208
rect 2118 1207 2124 1208
rect 2095 1206 2096 1207
rect 2091 1204 2096 1206
rect 2091 1203 2092 1204
rect 2086 1202 2092 1203
rect 2095 1203 2096 1204
rect 2100 1203 2101 1207
rect 2095 1202 2101 1203
rect 422 1198 428 1199
rect 300 1192 310 1194
rect 326 1195 332 1196
rect 300 1191 301 1192
rect 295 1190 301 1191
rect 326 1191 327 1195
rect 331 1194 332 1195
rect 335 1195 341 1196
rect 335 1194 336 1195
rect 331 1192 336 1194
rect 331 1191 332 1192
rect 326 1190 332 1191
rect 335 1191 336 1192
rect 340 1191 341 1195
rect 335 1190 341 1191
rect 358 1195 364 1196
rect 358 1191 359 1195
rect 363 1194 364 1195
rect 375 1195 381 1196
rect 375 1194 376 1195
rect 363 1192 376 1194
rect 363 1191 364 1192
rect 358 1190 364 1191
rect 375 1191 376 1192
rect 380 1191 381 1195
rect 375 1190 381 1191
rect 423 1195 429 1196
rect 423 1191 424 1195
rect 428 1194 429 1195
rect 462 1195 468 1196
rect 462 1194 463 1195
rect 428 1192 463 1194
rect 428 1191 429 1192
rect 423 1190 429 1191
rect 462 1191 463 1192
rect 467 1191 468 1195
rect 462 1190 468 1191
rect 471 1195 477 1196
rect 471 1191 472 1195
rect 476 1194 477 1195
rect 510 1195 516 1196
rect 510 1194 511 1195
rect 476 1192 511 1194
rect 476 1191 477 1192
rect 471 1190 477 1191
rect 510 1191 511 1192
rect 515 1191 516 1195
rect 510 1190 516 1191
rect 519 1195 525 1196
rect 519 1191 520 1195
rect 524 1194 525 1195
rect 566 1195 572 1196
rect 566 1194 567 1195
rect 524 1192 567 1194
rect 524 1191 525 1192
rect 519 1190 525 1191
rect 566 1191 567 1192
rect 571 1191 572 1195
rect 566 1190 572 1191
rect 574 1195 581 1196
rect 574 1191 575 1195
rect 580 1191 581 1195
rect 574 1190 581 1191
rect 583 1195 589 1196
rect 583 1191 584 1195
rect 588 1194 589 1195
rect 631 1195 637 1196
rect 631 1194 632 1195
rect 588 1192 632 1194
rect 588 1191 589 1192
rect 583 1190 589 1191
rect 631 1191 632 1192
rect 636 1191 637 1195
rect 631 1190 637 1191
rect 639 1195 645 1196
rect 639 1191 640 1195
rect 644 1194 645 1195
rect 695 1195 701 1196
rect 695 1194 696 1195
rect 644 1192 696 1194
rect 644 1191 645 1192
rect 639 1190 645 1191
rect 695 1191 696 1192
rect 700 1191 701 1195
rect 695 1190 701 1191
rect 703 1195 709 1196
rect 703 1191 704 1195
rect 708 1194 709 1195
rect 767 1195 773 1196
rect 767 1194 768 1195
rect 708 1192 768 1194
rect 708 1191 709 1192
rect 703 1190 709 1191
rect 767 1191 768 1192
rect 772 1191 773 1195
rect 767 1190 773 1191
rect 775 1195 781 1196
rect 775 1191 776 1195
rect 780 1194 781 1195
rect 839 1195 845 1196
rect 839 1194 840 1195
rect 780 1192 840 1194
rect 780 1191 781 1192
rect 775 1190 781 1191
rect 839 1191 840 1192
rect 844 1191 845 1195
rect 839 1190 845 1191
rect 847 1195 853 1196
rect 847 1191 848 1195
rect 852 1194 853 1195
rect 919 1195 925 1196
rect 919 1194 920 1195
rect 852 1192 920 1194
rect 852 1191 853 1192
rect 847 1190 853 1191
rect 919 1191 920 1192
rect 924 1191 925 1195
rect 919 1190 925 1191
rect 1006 1195 1013 1196
rect 1006 1191 1007 1195
rect 1012 1191 1013 1195
rect 1134 1195 1140 1196
rect 1006 1190 1013 1191
rect 1094 1192 1100 1193
rect 110 1187 116 1188
rect 1094 1188 1095 1192
rect 1099 1188 1100 1192
rect 1134 1191 1135 1195
rect 1139 1191 1140 1195
rect 2118 1195 2124 1196
rect 1134 1190 1140 1191
rect 1286 1192 1292 1193
rect 1094 1187 1100 1188
rect 1286 1188 1287 1192
rect 1291 1188 1292 1192
rect 1286 1187 1292 1188
rect 1326 1192 1332 1193
rect 1326 1188 1327 1192
rect 1331 1188 1332 1192
rect 1326 1187 1332 1188
rect 1374 1192 1380 1193
rect 1374 1188 1375 1192
rect 1379 1188 1380 1192
rect 1374 1187 1380 1188
rect 1430 1192 1436 1193
rect 1430 1188 1431 1192
rect 1435 1188 1436 1192
rect 1430 1187 1436 1188
rect 1494 1192 1500 1193
rect 1494 1188 1495 1192
rect 1499 1188 1500 1192
rect 1494 1187 1500 1188
rect 1558 1192 1564 1193
rect 1558 1188 1559 1192
rect 1563 1188 1564 1192
rect 1558 1187 1564 1188
rect 1622 1192 1628 1193
rect 1622 1188 1623 1192
rect 1627 1188 1628 1192
rect 1622 1187 1628 1188
rect 1678 1192 1684 1193
rect 1678 1188 1679 1192
rect 1683 1188 1684 1192
rect 1678 1187 1684 1188
rect 1734 1192 1740 1193
rect 1734 1188 1735 1192
rect 1739 1188 1740 1192
rect 1734 1187 1740 1188
rect 1790 1192 1796 1193
rect 1790 1188 1791 1192
rect 1795 1188 1796 1192
rect 1790 1187 1796 1188
rect 1846 1192 1852 1193
rect 1846 1188 1847 1192
rect 1851 1188 1852 1192
rect 1846 1187 1852 1188
rect 1902 1192 1908 1193
rect 1902 1188 1903 1192
rect 1907 1188 1908 1192
rect 1902 1187 1908 1188
rect 1966 1192 1972 1193
rect 1966 1188 1967 1192
rect 1971 1188 1972 1192
rect 1966 1187 1972 1188
rect 2030 1192 2036 1193
rect 2030 1188 2031 1192
rect 2035 1188 2036 1192
rect 2030 1187 2036 1188
rect 2070 1192 2076 1193
rect 2070 1188 2071 1192
rect 2075 1188 2076 1192
rect 2118 1191 2119 1195
rect 2123 1191 2124 1195
rect 2118 1190 2124 1191
rect 2070 1187 2076 1188
rect 270 1184 276 1185
rect 270 1180 271 1184
rect 275 1180 276 1184
rect 270 1179 276 1180
rect 310 1184 316 1185
rect 310 1180 311 1184
rect 315 1180 316 1184
rect 310 1179 316 1180
rect 350 1184 356 1185
rect 350 1180 351 1184
rect 355 1180 356 1184
rect 350 1179 356 1180
rect 398 1184 404 1185
rect 398 1180 399 1184
rect 403 1180 404 1184
rect 398 1179 404 1180
rect 446 1184 452 1185
rect 446 1180 447 1184
rect 451 1180 452 1184
rect 446 1179 452 1180
rect 494 1184 500 1185
rect 494 1180 495 1184
rect 499 1180 500 1184
rect 494 1179 500 1180
rect 550 1184 556 1185
rect 550 1180 551 1184
rect 555 1180 556 1184
rect 550 1179 556 1180
rect 606 1184 612 1185
rect 606 1180 607 1184
rect 611 1180 612 1184
rect 606 1179 612 1180
rect 670 1184 676 1185
rect 670 1180 671 1184
rect 675 1180 676 1184
rect 670 1179 676 1180
rect 742 1184 748 1185
rect 742 1180 743 1184
rect 747 1180 748 1184
rect 742 1179 748 1180
rect 814 1184 820 1185
rect 814 1180 815 1184
rect 819 1180 820 1184
rect 814 1179 820 1180
rect 894 1184 900 1185
rect 894 1180 895 1184
rect 899 1180 900 1184
rect 894 1179 900 1180
rect 982 1184 988 1185
rect 982 1180 983 1184
rect 987 1180 988 1184
rect 982 1179 988 1180
rect 1158 1180 1164 1181
rect 1134 1177 1140 1178
rect 295 1175 301 1176
rect 295 1171 296 1175
rect 300 1174 301 1175
rect 326 1175 332 1176
rect 326 1174 327 1175
rect 300 1172 327 1174
rect 300 1171 301 1172
rect 295 1170 301 1171
rect 326 1171 327 1172
rect 331 1171 332 1175
rect 326 1170 332 1171
rect 335 1175 341 1176
rect 335 1171 336 1175
rect 340 1174 341 1175
rect 358 1175 364 1176
rect 358 1174 359 1175
rect 340 1172 359 1174
rect 340 1171 341 1172
rect 335 1170 341 1171
rect 358 1171 359 1172
rect 363 1171 364 1175
rect 358 1170 364 1171
rect 375 1175 384 1176
rect 375 1171 376 1175
rect 383 1171 384 1175
rect 375 1170 384 1171
rect 422 1175 429 1176
rect 422 1171 423 1175
rect 428 1171 429 1175
rect 422 1170 429 1171
rect 462 1175 468 1176
rect 462 1171 463 1175
rect 467 1174 468 1175
rect 471 1175 477 1176
rect 471 1174 472 1175
rect 467 1172 472 1174
rect 467 1171 468 1172
rect 462 1170 468 1171
rect 471 1171 472 1172
rect 476 1171 477 1175
rect 471 1170 477 1171
rect 510 1175 516 1176
rect 510 1171 511 1175
rect 515 1174 516 1175
rect 519 1175 525 1176
rect 519 1174 520 1175
rect 515 1172 520 1174
rect 515 1171 516 1172
rect 510 1170 516 1171
rect 519 1171 520 1172
rect 524 1171 525 1175
rect 519 1170 525 1171
rect 575 1175 581 1176
rect 575 1171 576 1175
rect 580 1174 581 1175
rect 583 1175 589 1176
rect 583 1174 584 1175
rect 580 1172 584 1174
rect 580 1171 581 1172
rect 575 1170 581 1171
rect 583 1171 584 1172
rect 588 1171 589 1175
rect 583 1170 589 1171
rect 631 1175 637 1176
rect 631 1171 632 1175
rect 636 1174 637 1175
rect 639 1175 645 1176
rect 639 1174 640 1175
rect 636 1172 640 1174
rect 636 1171 637 1172
rect 631 1170 637 1171
rect 639 1171 640 1172
rect 644 1171 645 1175
rect 639 1170 645 1171
rect 695 1175 701 1176
rect 695 1171 696 1175
rect 700 1174 701 1175
rect 703 1175 709 1176
rect 703 1174 704 1175
rect 700 1172 704 1174
rect 700 1171 701 1172
rect 695 1170 701 1171
rect 703 1171 704 1172
rect 708 1171 709 1175
rect 703 1170 709 1171
rect 767 1175 773 1176
rect 767 1171 768 1175
rect 772 1174 773 1175
rect 775 1175 781 1176
rect 775 1174 776 1175
rect 772 1172 776 1174
rect 772 1171 773 1172
rect 767 1170 773 1171
rect 775 1171 776 1172
rect 780 1171 781 1175
rect 775 1170 781 1171
rect 839 1175 845 1176
rect 839 1171 840 1175
rect 844 1174 845 1175
rect 847 1175 853 1176
rect 847 1174 848 1175
rect 844 1172 848 1174
rect 844 1171 845 1172
rect 839 1170 845 1171
rect 847 1171 848 1172
rect 852 1171 853 1175
rect 847 1170 853 1171
rect 919 1175 925 1176
rect 919 1171 920 1175
rect 924 1171 925 1175
rect 919 1170 925 1171
rect 970 1175 976 1176
rect 970 1171 971 1175
rect 975 1174 976 1175
rect 1007 1175 1013 1176
rect 1007 1174 1008 1175
rect 975 1172 1008 1174
rect 975 1171 976 1172
rect 970 1170 976 1171
rect 1007 1171 1008 1172
rect 1012 1171 1013 1175
rect 1134 1173 1135 1177
rect 1139 1173 1140 1177
rect 1158 1176 1159 1180
rect 1163 1176 1164 1180
rect 1158 1175 1164 1176
rect 1206 1180 1212 1181
rect 1206 1176 1207 1180
rect 1211 1176 1212 1180
rect 1206 1175 1212 1176
rect 1278 1180 1284 1181
rect 1278 1176 1279 1180
rect 1283 1176 1284 1180
rect 1278 1175 1284 1176
rect 1350 1180 1356 1181
rect 1350 1176 1351 1180
rect 1355 1176 1356 1180
rect 1350 1175 1356 1176
rect 1422 1180 1428 1181
rect 1422 1176 1423 1180
rect 1427 1176 1428 1180
rect 1422 1175 1428 1176
rect 1486 1180 1492 1181
rect 1486 1176 1487 1180
rect 1491 1176 1492 1180
rect 1486 1175 1492 1176
rect 1558 1180 1564 1181
rect 1558 1176 1559 1180
rect 1563 1176 1564 1180
rect 1558 1175 1564 1176
rect 1630 1180 1636 1181
rect 1630 1176 1631 1180
rect 1635 1176 1636 1180
rect 1630 1175 1636 1176
rect 1710 1180 1716 1181
rect 1710 1176 1711 1180
rect 1715 1176 1716 1180
rect 1710 1175 1716 1176
rect 1798 1180 1804 1181
rect 1798 1176 1799 1180
rect 1803 1176 1804 1180
rect 1798 1175 1804 1176
rect 1886 1180 1892 1181
rect 1886 1176 1887 1180
rect 1891 1176 1892 1180
rect 1886 1175 1892 1176
rect 1982 1180 1988 1181
rect 1982 1176 1983 1180
rect 1987 1176 1988 1180
rect 1982 1175 1988 1176
rect 2070 1180 2076 1181
rect 2070 1176 2071 1180
rect 2075 1176 2076 1180
rect 2070 1175 2076 1176
rect 2118 1177 2124 1178
rect 1134 1172 1140 1173
rect 2118 1173 2119 1177
rect 2123 1173 2124 1177
rect 2118 1172 2124 1173
rect 1007 1170 1013 1171
rect 698 1167 704 1168
rect 698 1163 699 1167
rect 703 1166 704 1167
rect 921 1166 923 1170
rect 703 1164 923 1166
rect 703 1163 704 1164
rect 698 1162 704 1163
rect 1183 1163 1189 1164
rect 1183 1162 1184 1163
rect 1134 1160 1140 1161
rect 566 1159 572 1160
rect 566 1155 567 1159
rect 571 1158 572 1159
rect 662 1159 668 1160
rect 571 1156 642 1158
rect 571 1155 572 1156
rect 566 1154 572 1155
rect 423 1151 429 1152
rect 423 1147 424 1151
rect 428 1150 429 1151
rect 454 1151 460 1152
rect 454 1150 455 1151
rect 428 1148 455 1150
rect 428 1147 429 1148
rect 423 1146 429 1147
rect 454 1147 455 1148
rect 459 1147 460 1151
rect 454 1146 460 1147
rect 463 1151 469 1152
rect 463 1147 464 1151
rect 468 1150 469 1151
rect 494 1151 500 1152
rect 494 1150 495 1151
rect 468 1148 495 1150
rect 468 1147 469 1148
rect 463 1146 469 1147
rect 494 1147 495 1148
rect 499 1147 500 1151
rect 494 1146 500 1147
rect 503 1151 509 1152
rect 503 1147 504 1151
rect 508 1150 509 1151
rect 542 1151 548 1152
rect 542 1150 543 1151
rect 508 1148 543 1150
rect 508 1147 509 1148
rect 503 1146 509 1147
rect 542 1147 543 1148
rect 547 1147 548 1151
rect 542 1146 548 1147
rect 551 1151 557 1152
rect 551 1147 552 1151
rect 556 1150 557 1151
rect 590 1151 596 1152
rect 590 1150 591 1151
rect 556 1148 591 1150
rect 556 1147 557 1148
rect 551 1146 557 1147
rect 590 1147 591 1148
rect 595 1147 596 1151
rect 590 1146 596 1147
rect 599 1151 605 1152
rect 599 1147 600 1151
rect 604 1150 605 1151
rect 630 1151 636 1152
rect 630 1150 631 1151
rect 604 1148 631 1150
rect 604 1147 605 1148
rect 599 1146 605 1147
rect 630 1147 631 1148
rect 635 1147 636 1151
rect 640 1150 642 1156
rect 662 1155 663 1159
rect 667 1158 668 1159
rect 667 1156 914 1158
rect 667 1155 668 1156
rect 662 1154 668 1155
rect 912 1152 914 1156
rect 1134 1156 1135 1160
rect 1139 1156 1140 1160
rect 1134 1155 1140 1156
rect 1144 1160 1184 1162
rect 647 1151 653 1152
rect 647 1150 648 1151
rect 640 1148 648 1150
rect 630 1146 636 1147
rect 647 1147 648 1148
rect 652 1147 653 1151
rect 647 1146 653 1147
rect 695 1151 701 1152
rect 695 1147 696 1151
rect 700 1150 701 1151
rect 734 1151 740 1152
rect 734 1150 735 1151
rect 700 1148 735 1150
rect 700 1147 701 1148
rect 695 1146 701 1147
rect 734 1147 735 1148
rect 739 1147 740 1151
rect 734 1146 740 1147
rect 743 1151 749 1152
rect 743 1147 744 1151
rect 748 1150 749 1151
rect 790 1151 796 1152
rect 790 1150 791 1151
rect 748 1148 791 1150
rect 748 1147 749 1148
rect 743 1146 749 1147
rect 790 1147 791 1148
rect 795 1147 796 1151
rect 790 1146 796 1147
rect 799 1151 805 1152
rect 799 1147 800 1151
rect 804 1150 805 1151
rect 846 1151 852 1152
rect 846 1150 847 1151
rect 804 1148 847 1150
rect 804 1147 805 1148
rect 799 1146 805 1147
rect 846 1147 847 1148
rect 851 1147 852 1151
rect 846 1146 852 1147
rect 855 1151 861 1152
rect 855 1147 856 1151
rect 860 1150 861 1151
rect 902 1151 908 1152
rect 902 1150 903 1151
rect 860 1148 903 1150
rect 860 1147 861 1148
rect 855 1146 861 1147
rect 902 1147 903 1148
rect 907 1147 908 1151
rect 902 1146 908 1147
rect 911 1151 917 1152
rect 911 1147 912 1151
rect 916 1147 917 1151
rect 911 1146 917 1147
rect 967 1151 973 1152
rect 967 1147 968 1151
rect 972 1150 973 1151
rect 1022 1151 1028 1152
rect 1022 1150 1023 1151
rect 972 1148 1023 1150
rect 972 1147 973 1148
rect 967 1146 973 1147
rect 1022 1147 1023 1148
rect 1027 1147 1028 1151
rect 1022 1146 1028 1147
rect 1031 1151 1037 1152
rect 1031 1147 1032 1151
rect 1036 1150 1037 1151
rect 1062 1151 1068 1152
rect 1062 1150 1063 1151
rect 1036 1148 1063 1150
rect 1036 1147 1037 1148
rect 1031 1146 1037 1147
rect 1062 1147 1063 1148
rect 1067 1147 1068 1151
rect 1062 1146 1068 1147
rect 1071 1151 1077 1152
rect 1071 1147 1072 1151
rect 1076 1150 1077 1151
rect 1144 1150 1146 1160
rect 1183 1159 1184 1160
rect 1188 1159 1189 1163
rect 1183 1158 1189 1159
rect 1191 1163 1197 1164
rect 1191 1159 1192 1163
rect 1196 1162 1197 1163
rect 1231 1163 1237 1164
rect 1231 1162 1232 1163
rect 1196 1160 1232 1162
rect 1196 1159 1197 1160
rect 1191 1158 1197 1159
rect 1231 1159 1232 1160
rect 1236 1159 1237 1163
rect 1231 1158 1237 1159
rect 1239 1163 1245 1164
rect 1239 1159 1240 1163
rect 1244 1162 1245 1163
rect 1303 1163 1309 1164
rect 1303 1162 1304 1163
rect 1244 1160 1304 1162
rect 1244 1159 1245 1160
rect 1239 1158 1245 1159
rect 1303 1159 1304 1160
rect 1308 1159 1309 1163
rect 1303 1158 1309 1159
rect 1370 1163 1381 1164
rect 1370 1159 1371 1163
rect 1375 1159 1376 1163
rect 1380 1159 1381 1163
rect 1370 1158 1381 1159
rect 1383 1163 1389 1164
rect 1383 1159 1384 1163
rect 1388 1162 1389 1163
rect 1447 1163 1453 1164
rect 1447 1162 1448 1163
rect 1388 1160 1448 1162
rect 1388 1159 1389 1160
rect 1383 1158 1389 1159
rect 1447 1159 1448 1160
rect 1452 1159 1453 1163
rect 1447 1158 1453 1159
rect 1455 1163 1461 1164
rect 1455 1159 1456 1163
rect 1460 1162 1461 1163
rect 1511 1163 1517 1164
rect 1511 1162 1512 1163
rect 1460 1160 1512 1162
rect 1460 1159 1461 1160
rect 1455 1158 1461 1159
rect 1511 1159 1512 1160
rect 1516 1159 1517 1163
rect 1511 1158 1517 1159
rect 1582 1163 1589 1164
rect 1582 1159 1583 1163
rect 1588 1159 1589 1163
rect 1582 1158 1589 1159
rect 1591 1163 1597 1164
rect 1591 1159 1592 1163
rect 1596 1162 1597 1163
rect 1655 1163 1661 1164
rect 1655 1162 1656 1163
rect 1596 1160 1656 1162
rect 1596 1159 1597 1160
rect 1591 1158 1597 1159
rect 1655 1159 1656 1160
rect 1660 1159 1661 1163
rect 1655 1158 1661 1159
rect 1663 1163 1669 1164
rect 1663 1159 1664 1163
rect 1668 1162 1669 1163
rect 1735 1163 1741 1164
rect 1735 1162 1736 1163
rect 1668 1160 1736 1162
rect 1668 1159 1669 1160
rect 1663 1158 1669 1159
rect 1735 1159 1736 1160
rect 1740 1159 1741 1163
rect 1735 1158 1741 1159
rect 1743 1163 1749 1164
rect 1743 1159 1744 1163
rect 1748 1162 1749 1163
rect 1823 1163 1829 1164
rect 1823 1162 1824 1163
rect 1748 1160 1824 1162
rect 1748 1159 1749 1160
rect 1743 1158 1749 1159
rect 1823 1159 1824 1160
rect 1828 1159 1829 1163
rect 1823 1158 1829 1159
rect 1831 1163 1837 1164
rect 1831 1159 1832 1163
rect 1836 1162 1837 1163
rect 1911 1163 1917 1164
rect 1911 1162 1912 1163
rect 1836 1160 1912 1162
rect 1836 1159 1837 1160
rect 1831 1158 1837 1159
rect 1911 1159 1912 1160
rect 1916 1159 1917 1163
rect 1911 1158 1917 1159
rect 2006 1163 2013 1164
rect 2006 1159 2007 1163
rect 2012 1159 2013 1163
rect 2006 1158 2013 1159
rect 2094 1163 2101 1164
rect 2094 1159 2095 1163
rect 2100 1159 2101 1163
rect 2094 1158 2101 1159
rect 2118 1160 2124 1161
rect 2118 1156 2119 1160
rect 2123 1156 2124 1160
rect 2118 1155 2124 1156
rect 1076 1148 1146 1150
rect 1158 1152 1164 1153
rect 1158 1148 1159 1152
rect 1163 1148 1164 1152
rect 1076 1147 1077 1148
rect 1158 1147 1164 1148
rect 1206 1152 1212 1153
rect 1206 1148 1207 1152
rect 1211 1148 1212 1152
rect 1206 1147 1212 1148
rect 1278 1152 1284 1153
rect 1278 1148 1279 1152
rect 1283 1148 1284 1152
rect 1278 1147 1284 1148
rect 1350 1152 1356 1153
rect 1350 1148 1351 1152
rect 1355 1148 1356 1152
rect 1350 1147 1356 1148
rect 1422 1152 1428 1153
rect 1422 1148 1423 1152
rect 1427 1148 1428 1152
rect 1422 1147 1428 1148
rect 1486 1152 1492 1153
rect 1486 1148 1487 1152
rect 1491 1148 1492 1152
rect 1486 1147 1492 1148
rect 1558 1152 1564 1153
rect 1558 1148 1559 1152
rect 1563 1148 1564 1152
rect 1558 1147 1564 1148
rect 1630 1152 1636 1153
rect 1630 1148 1631 1152
rect 1635 1148 1636 1152
rect 1630 1147 1636 1148
rect 1710 1152 1716 1153
rect 1710 1148 1711 1152
rect 1715 1148 1716 1152
rect 1710 1147 1716 1148
rect 1798 1152 1804 1153
rect 1798 1148 1799 1152
rect 1803 1148 1804 1152
rect 1798 1147 1804 1148
rect 1886 1152 1892 1153
rect 1886 1148 1887 1152
rect 1891 1148 1892 1152
rect 1886 1147 1892 1148
rect 1982 1152 1988 1153
rect 1982 1148 1983 1152
rect 1987 1148 1988 1152
rect 1982 1147 1988 1148
rect 2070 1152 2076 1153
rect 2070 1148 2071 1152
rect 2075 1148 2076 1152
rect 2070 1147 2076 1148
rect 1071 1146 1077 1147
rect 398 1144 404 1145
rect 398 1140 399 1144
rect 403 1140 404 1144
rect 398 1139 404 1140
rect 438 1144 444 1145
rect 438 1140 439 1144
rect 443 1140 444 1144
rect 438 1139 444 1140
rect 478 1144 484 1145
rect 478 1140 479 1144
rect 483 1140 484 1144
rect 478 1139 484 1140
rect 526 1144 532 1145
rect 526 1140 527 1144
rect 531 1140 532 1144
rect 526 1139 532 1140
rect 574 1144 580 1145
rect 574 1140 575 1144
rect 579 1140 580 1144
rect 574 1139 580 1140
rect 622 1144 628 1145
rect 622 1140 623 1144
rect 627 1140 628 1144
rect 622 1139 628 1140
rect 670 1144 676 1145
rect 670 1140 671 1144
rect 675 1140 676 1144
rect 670 1139 676 1140
rect 718 1144 724 1145
rect 718 1140 719 1144
rect 723 1140 724 1144
rect 718 1139 724 1140
rect 774 1144 780 1145
rect 774 1140 775 1144
rect 779 1140 780 1144
rect 774 1139 780 1140
rect 830 1144 836 1145
rect 830 1140 831 1144
rect 835 1140 836 1144
rect 830 1139 836 1140
rect 886 1144 892 1145
rect 886 1140 887 1144
rect 891 1140 892 1144
rect 886 1139 892 1140
rect 942 1144 948 1145
rect 942 1140 943 1144
rect 947 1140 948 1144
rect 942 1139 948 1140
rect 1006 1144 1012 1145
rect 1006 1140 1007 1144
rect 1011 1140 1012 1144
rect 1006 1139 1012 1140
rect 1046 1144 1052 1145
rect 1046 1140 1047 1144
rect 1051 1140 1052 1144
rect 1046 1139 1052 1140
rect 1183 1143 1189 1144
rect 1183 1139 1184 1143
rect 1188 1142 1189 1143
rect 1191 1143 1197 1144
rect 1191 1142 1192 1143
rect 1188 1140 1192 1142
rect 1188 1139 1189 1140
rect 1183 1138 1189 1139
rect 1191 1139 1192 1140
rect 1196 1139 1197 1143
rect 1191 1138 1197 1139
rect 1231 1143 1237 1144
rect 1231 1139 1232 1143
rect 1236 1142 1237 1143
rect 1239 1143 1245 1144
rect 1239 1142 1240 1143
rect 1236 1140 1240 1142
rect 1236 1139 1237 1140
rect 1231 1138 1237 1139
rect 1239 1139 1240 1140
rect 1244 1139 1245 1143
rect 1239 1138 1245 1139
rect 1247 1143 1253 1144
rect 1247 1139 1248 1143
rect 1252 1142 1253 1143
rect 1303 1143 1309 1144
rect 1303 1142 1304 1143
rect 1252 1140 1304 1142
rect 1252 1139 1253 1140
rect 1247 1138 1253 1139
rect 1303 1139 1304 1140
rect 1308 1139 1309 1143
rect 1303 1138 1309 1139
rect 1375 1143 1381 1144
rect 1375 1139 1376 1143
rect 1380 1142 1381 1143
rect 1383 1143 1389 1144
rect 1383 1142 1384 1143
rect 1380 1140 1384 1142
rect 1380 1139 1381 1140
rect 1375 1138 1381 1139
rect 1383 1139 1384 1140
rect 1388 1139 1389 1143
rect 1383 1138 1389 1139
rect 1447 1143 1453 1144
rect 1447 1139 1448 1143
rect 1452 1142 1453 1143
rect 1455 1143 1461 1144
rect 1455 1142 1456 1143
rect 1452 1140 1456 1142
rect 1452 1139 1453 1140
rect 1447 1138 1453 1139
rect 1455 1139 1456 1140
rect 1460 1139 1461 1143
rect 1455 1138 1461 1139
rect 1511 1143 1520 1144
rect 1511 1139 1512 1143
rect 1519 1139 1520 1143
rect 1511 1138 1520 1139
rect 1583 1143 1589 1144
rect 1583 1139 1584 1143
rect 1588 1142 1589 1143
rect 1591 1143 1597 1144
rect 1591 1142 1592 1143
rect 1588 1140 1592 1142
rect 1588 1139 1589 1140
rect 1583 1138 1589 1139
rect 1591 1139 1592 1140
rect 1596 1139 1597 1143
rect 1591 1138 1597 1139
rect 1655 1143 1661 1144
rect 1655 1139 1656 1143
rect 1660 1142 1661 1143
rect 1663 1143 1669 1144
rect 1663 1142 1664 1143
rect 1660 1140 1664 1142
rect 1660 1139 1661 1140
rect 1655 1138 1661 1139
rect 1663 1139 1664 1140
rect 1668 1139 1669 1143
rect 1663 1138 1669 1139
rect 1735 1143 1741 1144
rect 1735 1139 1736 1143
rect 1740 1142 1741 1143
rect 1743 1143 1749 1144
rect 1743 1142 1744 1143
rect 1740 1140 1744 1142
rect 1740 1139 1741 1140
rect 1735 1138 1741 1139
rect 1743 1139 1744 1140
rect 1748 1139 1749 1143
rect 1743 1138 1749 1139
rect 1823 1143 1829 1144
rect 1823 1139 1824 1143
rect 1828 1142 1829 1143
rect 1831 1143 1837 1144
rect 1831 1142 1832 1143
rect 1828 1140 1832 1142
rect 1828 1139 1829 1140
rect 1823 1138 1829 1139
rect 1831 1139 1832 1140
rect 1836 1139 1837 1143
rect 1911 1143 1917 1144
rect 1911 1142 1912 1143
rect 1831 1138 1837 1139
rect 1840 1140 1912 1142
rect 110 1136 116 1137
rect 110 1132 111 1136
rect 115 1132 116 1136
rect 1094 1136 1100 1137
rect 1094 1132 1095 1136
rect 1099 1132 1100 1136
rect 110 1131 116 1132
rect 423 1131 432 1132
rect 423 1127 424 1131
rect 431 1127 432 1131
rect 423 1126 432 1127
rect 454 1131 460 1132
rect 454 1127 455 1131
rect 459 1130 460 1131
rect 463 1131 469 1132
rect 463 1130 464 1131
rect 459 1128 464 1130
rect 459 1127 460 1128
rect 454 1126 460 1127
rect 463 1127 464 1128
rect 468 1127 469 1131
rect 463 1126 469 1127
rect 494 1131 500 1132
rect 494 1127 495 1131
rect 499 1130 500 1131
rect 503 1131 509 1132
rect 503 1130 504 1131
rect 499 1128 504 1130
rect 499 1127 500 1128
rect 494 1126 500 1127
rect 503 1127 504 1128
rect 508 1127 509 1131
rect 503 1126 509 1127
rect 542 1131 548 1132
rect 542 1127 543 1131
rect 547 1130 548 1131
rect 551 1131 557 1132
rect 551 1130 552 1131
rect 547 1128 552 1130
rect 547 1127 548 1128
rect 542 1126 548 1127
rect 551 1127 552 1128
rect 556 1127 557 1131
rect 551 1126 557 1127
rect 590 1131 596 1132
rect 590 1127 591 1131
rect 595 1130 596 1131
rect 599 1131 605 1132
rect 599 1130 600 1131
rect 595 1128 600 1130
rect 595 1127 596 1128
rect 590 1126 596 1127
rect 599 1127 600 1128
rect 604 1127 605 1131
rect 599 1126 605 1127
rect 630 1131 636 1132
rect 630 1127 631 1131
rect 635 1130 636 1131
rect 647 1131 653 1132
rect 647 1130 648 1131
rect 635 1128 648 1130
rect 635 1127 636 1128
rect 630 1126 636 1127
rect 647 1127 648 1128
rect 652 1127 653 1131
rect 647 1126 653 1127
rect 695 1131 704 1132
rect 695 1127 696 1131
rect 703 1127 704 1131
rect 695 1126 704 1127
rect 734 1131 740 1132
rect 734 1127 735 1131
rect 739 1130 740 1131
rect 743 1131 749 1132
rect 743 1130 744 1131
rect 739 1128 744 1130
rect 739 1127 740 1128
rect 734 1126 740 1127
rect 743 1127 744 1128
rect 748 1127 749 1131
rect 743 1126 749 1127
rect 790 1131 796 1132
rect 790 1127 791 1131
rect 795 1130 796 1131
rect 799 1131 805 1132
rect 799 1130 800 1131
rect 795 1128 800 1130
rect 795 1127 796 1128
rect 790 1126 796 1127
rect 799 1127 800 1128
rect 804 1127 805 1131
rect 799 1126 805 1127
rect 846 1131 852 1132
rect 846 1127 847 1131
rect 851 1130 852 1131
rect 855 1131 861 1132
rect 855 1130 856 1131
rect 851 1128 856 1130
rect 851 1127 852 1128
rect 846 1126 852 1127
rect 855 1127 856 1128
rect 860 1127 861 1131
rect 855 1126 861 1127
rect 902 1131 908 1132
rect 902 1127 903 1131
rect 907 1130 908 1131
rect 911 1131 917 1132
rect 911 1130 912 1131
rect 907 1128 912 1130
rect 907 1127 908 1128
rect 902 1126 908 1127
rect 911 1127 912 1128
rect 916 1127 917 1131
rect 911 1126 917 1127
rect 967 1131 976 1132
rect 967 1127 968 1131
rect 975 1127 976 1131
rect 967 1126 976 1127
rect 1031 1131 1037 1132
rect 1031 1127 1032 1131
rect 1036 1130 1037 1131
rect 1054 1131 1060 1132
rect 1054 1130 1055 1131
rect 1036 1128 1055 1130
rect 1036 1127 1037 1128
rect 1031 1126 1037 1127
rect 1054 1127 1055 1128
rect 1059 1127 1060 1131
rect 1054 1126 1060 1127
rect 1062 1131 1068 1132
rect 1062 1127 1063 1131
rect 1067 1130 1068 1131
rect 1071 1131 1077 1132
rect 1094 1131 1100 1132
rect 1686 1135 1692 1136
rect 1686 1131 1687 1135
rect 1691 1134 1692 1135
rect 1840 1134 1842 1140
rect 1911 1139 1912 1140
rect 1916 1139 1917 1143
rect 1911 1138 1917 1139
rect 2002 1143 2013 1144
rect 2002 1139 2003 1143
rect 2007 1139 2008 1143
rect 2012 1139 2013 1143
rect 2002 1138 2013 1139
rect 2078 1143 2084 1144
rect 2078 1139 2079 1143
rect 2083 1142 2084 1143
rect 2095 1143 2101 1144
rect 2095 1142 2096 1143
rect 2083 1140 2096 1142
rect 2083 1139 2084 1140
rect 2078 1138 2084 1139
rect 2095 1139 2096 1140
rect 2100 1139 2101 1143
rect 2095 1138 2101 1139
rect 1691 1132 1842 1134
rect 1691 1131 1692 1132
rect 1071 1130 1072 1131
rect 1067 1128 1072 1130
rect 1067 1127 1068 1128
rect 1062 1126 1068 1127
rect 1071 1127 1072 1128
rect 1076 1127 1077 1131
rect 1686 1130 1692 1131
rect 1071 1126 1077 1127
rect 1582 1127 1588 1128
rect 1582 1123 1583 1127
rect 1587 1126 1588 1127
rect 1587 1124 1882 1126
rect 1587 1123 1588 1124
rect 1582 1122 1588 1123
rect 1880 1120 1882 1124
rect 110 1119 116 1120
rect 110 1115 111 1119
rect 115 1115 116 1119
rect 1094 1119 1100 1120
rect 110 1114 116 1115
rect 398 1116 404 1117
rect 398 1112 399 1116
rect 403 1112 404 1116
rect 398 1111 404 1112
rect 438 1116 444 1117
rect 438 1112 439 1116
rect 443 1112 444 1116
rect 438 1111 444 1112
rect 478 1116 484 1117
rect 478 1112 479 1116
rect 483 1112 484 1116
rect 478 1111 484 1112
rect 526 1116 532 1117
rect 526 1112 527 1116
rect 531 1112 532 1116
rect 526 1111 532 1112
rect 574 1116 580 1117
rect 574 1112 575 1116
rect 579 1112 580 1116
rect 574 1111 580 1112
rect 622 1116 628 1117
rect 622 1112 623 1116
rect 627 1112 628 1116
rect 622 1111 628 1112
rect 670 1116 676 1117
rect 670 1112 671 1116
rect 675 1112 676 1116
rect 670 1111 676 1112
rect 718 1116 724 1117
rect 718 1112 719 1116
rect 723 1112 724 1116
rect 718 1111 724 1112
rect 774 1116 780 1117
rect 774 1112 775 1116
rect 779 1112 780 1116
rect 774 1111 780 1112
rect 830 1116 836 1117
rect 830 1112 831 1116
rect 835 1112 836 1116
rect 830 1111 836 1112
rect 886 1116 892 1117
rect 886 1112 887 1116
rect 891 1112 892 1116
rect 886 1111 892 1112
rect 942 1116 948 1117
rect 942 1112 943 1116
rect 947 1112 948 1116
rect 942 1111 948 1112
rect 1006 1116 1012 1117
rect 1006 1112 1007 1116
rect 1011 1112 1012 1116
rect 1006 1111 1012 1112
rect 1046 1116 1052 1117
rect 1046 1112 1047 1116
rect 1051 1112 1052 1116
rect 1094 1115 1095 1119
rect 1099 1115 1100 1119
rect 1094 1114 1100 1115
rect 1215 1119 1221 1120
rect 1215 1115 1216 1119
rect 1220 1118 1221 1119
rect 1286 1119 1292 1120
rect 1286 1118 1287 1119
rect 1220 1116 1287 1118
rect 1220 1115 1221 1116
rect 1215 1114 1221 1115
rect 1286 1115 1287 1116
rect 1291 1115 1292 1119
rect 1286 1114 1292 1115
rect 1295 1119 1301 1120
rect 1295 1115 1296 1119
rect 1300 1118 1301 1119
rect 1326 1119 1332 1120
rect 1326 1118 1327 1119
rect 1300 1116 1327 1118
rect 1300 1115 1301 1116
rect 1295 1114 1301 1115
rect 1326 1115 1327 1116
rect 1331 1115 1332 1119
rect 1326 1114 1332 1115
rect 1367 1119 1376 1120
rect 1367 1115 1368 1119
rect 1375 1115 1376 1119
rect 1367 1114 1376 1115
rect 1439 1119 1445 1120
rect 1439 1115 1440 1119
rect 1444 1118 1445 1119
rect 1478 1119 1484 1120
rect 1478 1118 1479 1119
rect 1444 1116 1479 1118
rect 1444 1115 1445 1116
rect 1439 1114 1445 1115
rect 1478 1115 1479 1116
rect 1483 1115 1484 1119
rect 1478 1114 1484 1115
rect 1511 1119 1517 1120
rect 1511 1115 1512 1119
rect 1516 1118 1517 1119
rect 1582 1119 1588 1120
rect 1582 1118 1583 1119
rect 1516 1116 1583 1118
rect 1516 1115 1517 1116
rect 1511 1114 1517 1115
rect 1582 1115 1583 1116
rect 1587 1115 1588 1119
rect 1582 1114 1588 1115
rect 1591 1119 1597 1120
rect 1591 1115 1592 1119
rect 1596 1118 1597 1119
rect 1670 1119 1676 1120
rect 1670 1118 1671 1119
rect 1596 1116 1671 1118
rect 1596 1115 1597 1116
rect 1591 1114 1597 1115
rect 1670 1115 1671 1116
rect 1675 1115 1676 1119
rect 1670 1114 1676 1115
rect 1679 1119 1685 1120
rect 1679 1115 1680 1119
rect 1684 1118 1685 1119
rect 1766 1119 1772 1120
rect 1766 1118 1767 1119
rect 1684 1116 1767 1118
rect 1684 1115 1685 1116
rect 1679 1114 1685 1115
rect 1766 1115 1767 1116
rect 1771 1115 1772 1119
rect 1766 1114 1772 1115
rect 1775 1119 1781 1120
rect 1775 1115 1776 1119
rect 1780 1118 1781 1119
rect 1870 1119 1876 1120
rect 1870 1118 1871 1119
rect 1780 1116 1871 1118
rect 1780 1115 1781 1116
rect 1775 1114 1781 1115
rect 1870 1115 1871 1116
rect 1875 1115 1876 1119
rect 1870 1114 1876 1115
rect 1879 1119 1885 1120
rect 1879 1115 1880 1119
rect 1884 1115 1885 1119
rect 1879 1114 1885 1115
rect 1982 1119 1989 1120
rect 1982 1115 1983 1119
rect 1988 1115 1989 1119
rect 1982 1114 1989 1115
rect 2094 1119 2101 1120
rect 2094 1115 2095 1119
rect 2100 1115 2101 1119
rect 2094 1114 2101 1115
rect 1046 1111 1052 1112
rect 1190 1112 1196 1113
rect 1190 1108 1191 1112
rect 1195 1108 1196 1112
rect 1190 1107 1196 1108
rect 1270 1112 1276 1113
rect 1270 1108 1271 1112
rect 1275 1108 1276 1112
rect 1270 1107 1276 1108
rect 1342 1112 1348 1113
rect 1342 1108 1343 1112
rect 1347 1108 1348 1112
rect 1342 1107 1348 1108
rect 1414 1112 1420 1113
rect 1414 1108 1415 1112
rect 1419 1108 1420 1112
rect 1414 1107 1420 1108
rect 1486 1112 1492 1113
rect 1486 1108 1487 1112
rect 1491 1108 1492 1112
rect 1486 1107 1492 1108
rect 1566 1112 1572 1113
rect 1566 1108 1567 1112
rect 1571 1108 1572 1112
rect 1566 1107 1572 1108
rect 1654 1112 1660 1113
rect 1654 1108 1655 1112
rect 1659 1108 1660 1112
rect 1654 1107 1660 1108
rect 1750 1112 1756 1113
rect 1750 1108 1751 1112
rect 1755 1108 1756 1112
rect 1750 1107 1756 1108
rect 1854 1112 1860 1113
rect 1854 1108 1855 1112
rect 1859 1108 1860 1112
rect 1854 1107 1860 1108
rect 1958 1112 1964 1113
rect 1958 1108 1959 1112
rect 1963 1108 1964 1112
rect 1958 1107 1964 1108
rect 2070 1112 2076 1113
rect 2070 1108 2071 1112
rect 2075 1108 2076 1112
rect 2070 1107 2076 1108
rect 158 1104 164 1105
rect 110 1101 116 1102
rect 110 1097 111 1101
rect 115 1097 116 1101
rect 158 1100 159 1104
rect 163 1100 164 1104
rect 158 1099 164 1100
rect 198 1104 204 1105
rect 198 1100 199 1104
rect 203 1100 204 1104
rect 198 1099 204 1100
rect 254 1104 260 1105
rect 254 1100 255 1104
rect 259 1100 260 1104
rect 254 1099 260 1100
rect 318 1104 324 1105
rect 318 1100 319 1104
rect 323 1100 324 1104
rect 318 1099 324 1100
rect 398 1104 404 1105
rect 398 1100 399 1104
rect 403 1100 404 1104
rect 398 1099 404 1100
rect 478 1104 484 1105
rect 478 1100 479 1104
rect 483 1100 484 1104
rect 478 1099 484 1100
rect 558 1104 564 1105
rect 558 1100 559 1104
rect 563 1100 564 1104
rect 558 1099 564 1100
rect 638 1104 644 1105
rect 638 1100 639 1104
rect 643 1100 644 1104
rect 638 1099 644 1100
rect 710 1104 716 1105
rect 710 1100 711 1104
rect 715 1100 716 1104
rect 710 1099 716 1100
rect 782 1104 788 1105
rect 782 1100 783 1104
rect 787 1100 788 1104
rect 782 1099 788 1100
rect 854 1104 860 1105
rect 854 1100 855 1104
rect 859 1100 860 1104
rect 854 1099 860 1100
rect 926 1104 932 1105
rect 926 1100 927 1104
rect 931 1100 932 1104
rect 926 1099 932 1100
rect 998 1104 1004 1105
rect 998 1100 999 1104
rect 1003 1100 1004 1104
rect 998 1099 1004 1100
rect 1046 1104 1052 1105
rect 1046 1100 1047 1104
rect 1051 1100 1052 1104
rect 1134 1104 1140 1105
rect 2118 1104 2124 1105
rect 1046 1099 1052 1100
rect 1094 1101 1100 1102
rect 110 1096 116 1097
rect 1094 1097 1095 1101
rect 1099 1097 1100 1101
rect 1134 1100 1135 1104
rect 1139 1100 1140 1104
rect 2002 1103 2008 1104
rect 2002 1102 2003 1103
rect 1983 1101 2003 1102
rect 1134 1099 1140 1100
rect 1215 1099 1221 1100
rect 1094 1096 1100 1097
rect 1215 1095 1216 1099
rect 1220 1098 1221 1099
rect 1247 1099 1253 1100
rect 1247 1098 1248 1099
rect 1220 1096 1248 1098
rect 1220 1095 1221 1096
rect 1215 1094 1221 1095
rect 1247 1095 1248 1096
rect 1252 1095 1253 1099
rect 1247 1094 1253 1095
rect 1286 1099 1292 1100
rect 1286 1095 1287 1099
rect 1291 1098 1292 1099
rect 1295 1099 1301 1100
rect 1295 1098 1296 1099
rect 1291 1096 1296 1098
rect 1291 1095 1292 1096
rect 1286 1094 1292 1095
rect 1295 1095 1296 1096
rect 1300 1095 1301 1099
rect 1295 1094 1301 1095
rect 1367 1099 1376 1100
rect 1367 1095 1368 1099
rect 1375 1095 1376 1099
rect 1367 1094 1376 1095
rect 1439 1099 1445 1100
rect 1439 1095 1440 1099
rect 1444 1098 1445 1099
rect 1470 1099 1476 1100
rect 1470 1098 1471 1099
rect 1444 1096 1471 1098
rect 1444 1095 1445 1096
rect 1439 1094 1445 1095
rect 1470 1095 1471 1096
rect 1475 1095 1476 1099
rect 1470 1094 1476 1095
rect 1494 1099 1500 1100
rect 1494 1095 1495 1099
rect 1499 1098 1500 1099
rect 1511 1099 1517 1100
rect 1511 1098 1512 1099
rect 1499 1096 1512 1098
rect 1499 1095 1500 1096
rect 1494 1094 1500 1095
rect 1511 1095 1512 1096
rect 1516 1095 1517 1099
rect 1511 1094 1517 1095
rect 1582 1099 1588 1100
rect 1582 1095 1583 1099
rect 1587 1098 1588 1099
rect 1591 1099 1597 1100
rect 1591 1098 1592 1099
rect 1587 1096 1592 1098
rect 1587 1095 1588 1096
rect 1582 1094 1588 1095
rect 1591 1095 1592 1096
rect 1596 1095 1597 1099
rect 1591 1094 1597 1095
rect 1670 1099 1676 1100
rect 1670 1095 1671 1099
rect 1675 1098 1676 1099
rect 1679 1099 1685 1100
rect 1679 1098 1680 1099
rect 1675 1096 1680 1098
rect 1675 1095 1676 1096
rect 1670 1094 1676 1095
rect 1679 1095 1680 1096
rect 1684 1095 1685 1099
rect 1679 1094 1685 1095
rect 1766 1099 1772 1100
rect 1766 1095 1767 1099
rect 1771 1098 1772 1099
rect 1775 1099 1781 1100
rect 1775 1098 1776 1099
rect 1771 1096 1776 1098
rect 1771 1095 1772 1096
rect 1766 1094 1772 1095
rect 1775 1095 1776 1096
rect 1780 1095 1781 1099
rect 1775 1094 1781 1095
rect 1870 1099 1876 1100
rect 1870 1095 1871 1099
rect 1875 1098 1876 1099
rect 1879 1099 1885 1100
rect 1879 1098 1880 1099
rect 1875 1096 1880 1098
rect 1875 1095 1876 1096
rect 1870 1094 1876 1095
rect 1879 1095 1880 1096
rect 1884 1095 1885 1099
rect 1983 1097 1984 1101
rect 1988 1100 2003 1101
rect 1988 1097 1989 1100
rect 2002 1099 2003 1100
rect 2007 1099 2008 1103
rect 2118 1100 2119 1104
rect 2123 1100 2124 1104
rect 2002 1098 2008 1099
rect 2094 1099 2101 1100
rect 2118 1099 2124 1100
rect 1983 1096 1989 1097
rect 1879 1094 1885 1095
rect 2094 1095 2095 1099
rect 2100 1095 2101 1099
rect 2094 1094 2101 1095
rect 183 1087 192 1088
rect 110 1084 116 1085
rect 110 1080 111 1084
rect 115 1080 116 1084
rect 183 1083 184 1087
rect 191 1083 192 1087
rect 183 1082 192 1083
rect 206 1087 212 1088
rect 206 1083 207 1087
rect 211 1086 212 1087
rect 223 1087 229 1088
rect 223 1086 224 1087
rect 211 1084 224 1086
rect 211 1083 212 1084
rect 206 1082 212 1083
rect 223 1083 224 1084
rect 228 1083 229 1087
rect 223 1082 229 1083
rect 231 1087 237 1088
rect 231 1083 232 1087
rect 236 1086 237 1087
rect 279 1087 285 1088
rect 279 1086 280 1087
rect 236 1084 280 1086
rect 236 1083 237 1084
rect 231 1082 237 1083
rect 279 1083 280 1084
rect 284 1083 285 1087
rect 279 1082 285 1083
rect 287 1087 293 1088
rect 287 1083 288 1087
rect 292 1086 293 1087
rect 343 1087 349 1088
rect 343 1086 344 1087
rect 292 1084 344 1086
rect 292 1083 293 1084
rect 287 1082 293 1083
rect 343 1083 344 1084
rect 348 1083 349 1087
rect 343 1082 349 1083
rect 351 1087 357 1088
rect 351 1083 352 1087
rect 356 1086 357 1087
rect 423 1087 429 1088
rect 423 1086 424 1087
rect 356 1084 424 1086
rect 356 1083 357 1084
rect 351 1082 357 1083
rect 423 1083 424 1084
rect 428 1083 429 1087
rect 423 1082 429 1083
rect 431 1087 437 1088
rect 431 1083 432 1087
rect 436 1086 437 1087
rect 503 1087 509 1088
rect 503 1086 504 1087
rect 436 1084 504 1086
rect 436 1083 437 1084
rect 431 1082 437 1083
rect 503 1083 504 1084
rect 508 1083 509 1087
rect 503 1082 509 1083
rect 511 1087 517 1088
rect 511 1083 512 1087
rect 516 1086 517 1087
rect 583 1087 589 1088
rect 583 1086 584 1087
rect 516 1084 584 1086
rect 516 1083 517 1084
rect 511 1082 517 1083
rect 583 1083 584 1084
rect 588 1083 589 1087
rect 583 1082 589 1083
rect 662 1087 669 1088
rect 662 1083 663 1087
rect 668 1083 669 1087
rect 662 1082 669 1083
rect 671 1087 677 1088
rect 671 1083 672 1087
rect 676 1086 677 1087
rect 735 1087 741 1088
rect 735 1086 736 1087
rect 676 1084 736 1086
rect 676 1083 677 1084
rect 671 1082 677 1083
rect 735 1083 736 1084
rect 740 1083 741 1087
rect 735 1082 741 1083
rect 743 1087 749 1088
rect 743 1083 744 1087
rect 748 1086 749 1087
rect 807 1087 813 1088
rect 807 1086 808 1087
rect 748 1084 808 1086
rect 748 1083 749 1084
rect 743 1082 749 1083
rect 807 1083 808 1084
rect 812 1083 813 1087
rect 807 1082 813 1083
rect 815 1087 821 1088
rect 815 1083 816 1087
rect 820 1086 821 1087
rect 879 1087 885 1088
rect 879 1086 880 1087
rect 820 1084 880 1086
rect 820 1083 821 1084
rect 815 1082 821 1083
rect 879 1083 880 1084
rect 884 1083 885 1087
rect 879 1082 885 1083
rect 951 1087 957 1088
rect 951 1083 952 1087
rect 956 1086 957 1087
rect 1014 1087 1020 1088
rect 1014 1086 1015 1087
rect 956 1084 1015 1086
rect 956 1083 957 1084
rect 951 1082 957 1083
rect 1014 1083 1015 1084
rect 1019 1083 1020 1087
rect 1014 1082 1020 1083
rect 1022 1087 1029 1088
rect 1022 1083 1023 1087
rect 1028 1083 1029 1087
rect 1022 1082 1029 1083
rect 1071 1087 1077 1088
rect 1071 1083 1072 1087
rect 1076 1086 1077 1087
rect 1086 1087 1092 1088
rect 1086 1086 1087 1087
rect 1076 1084 1087 1086
rect 1076 1083 1077 1084
rect 1071 1082 1077 1083
rect 1086 1083 1087 1084
rect 1091 1083 1092 1087
rect 1134 1087 1140 1088
rect 1086 1082 1092 1083
rect 1094 1084 1100 1085
rect 110 1079 116 1080
rect 1094 1080 1095 1084
rect 1099 1080 1100 1084
rect 1134 1083 1135 1087
rect 1139 1083 1140 1087
rect 2118 1087 2124 1088
rect 1134 1082 1140 1083
rect 1190 1084 1196 1085
rect 1094 1079 1100 1080
rect 1190 1080 1191 1084
rect 1195 1080 1196 1084
rect 1190 1079 1196 1080
rect 1270 1084 1276 1085
rect 1270 1080 1271 1084
rect 1275 1080 1276 1084
rect 1270 1079 1276 1080
rect 1342 1084 1348 1085
rect 1342 1080 1343 1084
rect 1347 1080 1348 1084
rect 1342 1079 1348 1080
rect 1414 1084 1420 1085
rect 1414 1080 1415 1084
rect 1419 1080 1420 1084
rect 1414 1079 1420 1080
rect 1486 1084 1492 1085
rect 1486 1080 1487 1084
rect 1491 1080 1492 1084
rect 1486 1079 1492 1080
rect 1566 1084 1572 1085
rect 1566 1080 1567 1084
rect 1571 1080 1572 1084
rect 1566 1079 1572 1080
rect 1654 1084 1660 1085
rect 1654 1080 1655 1084
rect 1659 1080 1660 1084
rect 1654 1079 1660 1080
rect 1750 1084 1756 1085
rect 1750 1080 1751 1084
rect 1755 1080 1756 1084
rect 1750 1079 1756 1080
rect 1854 1084 1860 1085
rect 1854 1080 1855 1084
rect 1859 1080 1860 1084
rect 1854 1079 1860 1080
rect 1958 1084 1964 1085
rect 1958 1080 1959 1084
rect 1963 1080 1964 1084
rect 1958 1079 1964 1080
rect 2070 1084 2076 1085
rect 2070 1080 2071 1084
rect 2075 1080 2076 1084
rect 2118 1083 2119 1087
rect 2123 1083 2124 1087
rect 2118 1082 2124 1083
rect 2070 1079 2076 1080
rect 158 1076 164 1077
rect 158 1072 159 1076
rect 163 1072 164 1076
rect 158 1071 164 1072
rect 198 1076 204 1077
rect 198 1072 199 1076
rect 203 1072 204 1076
rect 198 1071 204 1072
rect 254 1076 260 1077
rect 254 1072 255 1076
rect 259 1072 260 1076
rect 254 1071 260 1072
rect 318 1076 324 1077
rect 318 1072 319 1076
rect 323 1072 324 1076
rect 318 1071 324 1072
rect 398 1076 404 1077
rect 398 1072 399 1076
rect 403 1072 404 1076
rect 398 1071 404 1072
rect 478 1076 484 1077
rect 478 1072 479 1076
rect 483 1072 484 1076
rect 478 1071 484 1072
rect 558 1076 564 1077
rect 558 1072 559 1076
rect 563 1072 564 1076
rect 558 1071 564 1072
rect 638 1076 644 1077
rect 638 1072 639 1076
rect 643 1072 644 1076
rect 638 1071 644 1072
rect 710 1076 716 1077
rect 710 1072 711 1076
rect 715 1072 716 1076
rect 710 1071 716 1072
rect 782 1076 788 1077
rect 782 1072 783 1076
rect 787 1072 788 1076
rect 782 1071 788 1072
rect 854 1076 860 1077
rect 854 1072 855 1076
rect 859 1072 860 1076
rect 854 1071 860 1072
rect 926 1076 932 1077
rect 926 1072 927 1076
rect 931 1072 932 1076
rect 926 1071 932 1072
rect 998 1076 1004 1077
rect 998 1072 999 1076
rect 1003 1072 1004 1076
rect 998 1071 1004 1072
rect 1046 1076 1052 1077
rect 1046 1072 1047 1076
rect 1051 1072 1052 1076
rect 1046 1071 1052 1072
rect 1158 1072 1164 1073
rect 1134 1069 1140 1070
rect 183 1067 189 1068
rect 183 1063 184 1067
rect 188 1066 189 1067
rect 206 1067 212 1068
rect 206 1066 207 1067
rect 188 1064 207 1066
rect 188 1063 189 1064
rect 183 1062 189 1063
rect 206 1063 207 1064
rect 211 1063 212 1067
rect 206 1062 212 1063
rect 223 1067 229 1068
rect 223 1063 224 1067
rect 228 1066 229 1067
rect 231 1067 237 1068
rect 231 1066 232 1067
rect 228 1064 232 1066
rect 228 1063 229 1064
rect 223 1062 229 1063
rect 231 1063 232 1064
rect 236 1063 237 1067
rect 231 1062 237 1063
rect 279 1067 285 1068
rect 279 1063 280 1067
rect 284 1066 285 1067
rect 287 1067 293 1068
rect 287 1066 288 1067
rect 284 1064 288 1066
rect 284 1063 285 1064
rect 279 1062 285 1063
rect 287 1063 288 1064
rect 292 1063 293 1067
rect 287 1062 293 1063
rect 343 1067 349 1068
rect 343 1063 344 1067
rect 348 1066 349 1067
rect 351 1067 357 1068
rect 351 1066 352 1067
rect 348 1064 352 1066
rect 348 1063 349 1064
rect 343 1062 349 1063
rect 351 1063 352 1064
rect 356 1063 357 1067
rect 351 1062 357 1063
rect 423 1067 429 1068
rect 423 1063 424 1067
rect 428 1066 429 1067
rect 431 1067 437 1068
rect 431 1066 432 1067
rect 428 1064 432 1066
rect 428 1063 429 1064
rect 423 1062 429 1063
rect 431 1063 432 1064
rect 436 1063 437 1067
rect 431 1062 437 1063
rect 503 1067 509 1068
rect 503 1063 504 1067
rect 508 1066 509 1067
rect 511 1067 517 1068
rect 511 1066 512 1067
rect 508 1064 512 1066
rect 508 1063 509 1064
rect 503 1062 509 1063
rect 511 1063 512 1064
rect 516 1063 517 1067
rect 511 1062 517 1063
rect 583 1067 589 1068
rect 583 1063 584 1067
rect 588 1063 589 1067
rect 583 1062 589 1063
rect 663 1067 669 1068
rect 663 1063 664 1067
rect 668 1066 669 1067
rect 671 1067 677 1068
rect 671 1066 672 1067
rect 668 1064 672 1066
rect 668 1063 669 1064
rect 663 1062 669 1063
rect 671 1063 672 1064
rect 676 1063 677 1067
rect 671 1062 677 1063
rect 735 1067 741 1068
rect 735 1063 736 1067
rect 740 1066 741 1067
rect 743 1067 749 1068
rect 743 1066 744 1067
rect 740 1064 744 1066
rect 740 1063 741 1064
rect 735 1062 741 1063
rect 743 1063 744 1064
rect 748 1063 749 1067
rect 743 1062 749 1063
rect 807 1067 813 1068
rect 807 1063 808 1067
rect 812 1066 813 1067
rect 815 1067 821 1068
rect 815 1066 816 1067
rect 812 1064 816 1066
rect 812 1063 813 1064
rect 807 1062 813 1063
rect 815 1063 816 1064
rect 820 1063 821 1067
rect 815 1062 821 1063
rect 879 1067 888 1068
rect 879 1063 880 1067
rect 887 1063 888 1067
rect 879 1062 888 1063
rect 951 1067 957 1068
rect 951 1063 952 1067
rect 956 1063 957 1067
rect 951 1062 957 1063
rect 1014 1067 1020 1068
rect 1014 1063 1015 1067
rect 1019 1066 1020 1067
rect 1023 1067 1029 1068
rect 1023 1066 1024 1067
rect 1019 1064 1024 1066
rect 1019 1063 1020 1064
rect 1014 1062 1020 1063
rect 1023 1063 1024 1064
rect 1028 1063 1029 1067
rect 1023 1062 1029 1063
rect 1054 1067 1060 1068
rect 1054 1063 1055 1067
rect 1059 1066 1060 1067
rect 1071 1067 1077 1068
rect 1071 1066 1072 1067
rect 1059 1064 1072 1066
rect 1059 1063 1060 1064
rect 1054 1062 1060 1063
rect 1071 1063 1072 1064
rect 1076 1063 1077 1067
rect 1134 1065 1135 1069
rect 1139 1065 1140 1069
rect 1158 1068 1159 1072
rect 1163 1068 1164 1072
rect 1158 1067 1164 1068
rect 1198 1072 1204 1073
rect 1198 1068 1199 1072
rect 1203 1068 1204 1072
rect 1198 1067 1204 1068
rect 1246 1072 1252 1073
rect 1246 1068 1247 1072
rect 1251 1068 1252 1072
rect 1246 1067 1252 1068
rect 1302 1072 1308 1073
rect 1302 1068 1303 1072
rect 1307 1068 1308 1072
rect 1302 1067 1308 1068
rect 1350 1072 1356 1073
rect 1350 1068 1351 1072
rect 1355 1068 1356 1072
rect 1350 1067 1356 1068
rect 1398 1072 1404 1073
rect 1398 1068 1399 1072
rect 1403 1068 1404 1072
rect 1398 1067 1404 1068
rect 1454 1072 1460 1073
rect 1454 1068 1455 1072
rect 1459 1068 1460 1072
rect 1454 1067 1460 1068
rect 1510 1072 1516 1073
rect 1510 1068 1511 1072
rect 1515 1068 1516 1072
rect 1510 1067 1516 1068
rect 1582 1072 1588 1073
rect 1582 1068 1583 1072
rect 1587 1068 1588 1072
rect 1582 1067 1588 1068
rect 1662 1072 1668 1073
rect 1662 1068 1663 1072
rect 1667 1068 1668 1072
rect 1662 1067 1668 1068
rect 1758 1072 1764 1073
rect 1758 1068 1759 1072
rect 1763 1068 1764 1072
rect 1758 1067 1764 1068
rect 1862 1072 1868 1073
rect 1862 1068 1863 1072
rect 1867 1068 1868 1072
rect 1862 1067 1868 1068
rect 1966 1072 1972 1073
rect 1966 1068 1967 1072
rect 1971 1068 1972 1072
rect 1966 1067 1972 1068
rect 2070 1072 2076 1073
rect 2070 1068 2071 1072
rect 2075 1068 2076 1072
rect 2070 1067 2076 1068
rect 2118 1069 2124 1070
rect 1134 1064 1140 1065
rect 2118 1065 2119 1069
rect 2123 1065 2124 1069
rect 2118 1064 2124 1065
rect 1071 1062 1077 1063
rect 1886 1063 1892 1064
rect 1886 1062 1887 1063
rect 166 1059 172 1060
rect 166 1055 167 1059
rect 171 1058 172 1059
rect 426 1059 432 1060
rect 171 1056 321 1058
rect 171 1055 172 1056
rect 166 1054 172 1055
rect 186 1051 192 1052
rect 186 1047 187 1051
rect 191 1050 192 1051
rect 319 1050 321 1056
rect 426 1055 427 1059
rect 431 1058 432 1059
rect 585 1058 587 1062
rect 431 1056 587 1058
rect 602 1059 608 1060
rect 431 1055 432 1056
rect 426 1054 432 1055
rect 602 1055 603 1059
rect 607 1058 608 1059
rect 953 1058 955 1062
rect 607 1056 955 1058
rect 1609 1060 1887 1062
rect 1609 1056 1611 1060
rect 1886 1059 1887 1060
rect 1891 1059 1892 1063
rect 1886 1058 1892 1059
rect 607 1055 608 1056
rect 602 1054 608 1055
rect 1183 1055 1189 1056
rect 1134 1052 1140 1053
rect 191 1048 282 1050
rect 319 1048 475 1050
rect 191 1047 192 1048
rect 186 1046 192 1047
rect 280 1044 282 1048
rect 473 1044 475 1048
rect 1134 1048 1135 1052
rect 1139 1048 1140 1052
rect 1183 1051 1184 1055
rect 1188 1054 1189 1055
rect 1214 1055 1220 1056
rect 1214 1054 1215 1055
rect 1188 1052 1215 1054
rect 1188 1051 1189 1052
rect 1183 1050 1189 1051
rect 1214 1051 1215 1052
rect 1219 1051 1220 1055
rect 1214 1050 1220 1051
rect 1222 1055 1229 1056
rect 1222 1051 1223 1055
rect 1228 1051 1229 1055
rect 1222 1050 1229 1051
rect 1271 1055 1277 1056
rect 1271 1051 1272 1055
rect 1276 1054 1277 1055
rect 1318 1055 1324 1056
rect 1318 1054 1319 1055
rect 1276 1052 1319 1054
rect 1276 1051 1277 1052
rect 1271 1050 1277 1051
rect 1318 1051 1319 1052
rect 1323 1051 1324 1055
rect 1318 1050 1324 1051
rect 1326 1055 1333 1056
rect 1326 1051 1327 1055
rect 1332 1051 1333 1055
rect 1326 1050 1333 1051
rect 1375 1055 1381 1056
rect 1375 1051 1376 1055
rect 1380 1054 1381 1055
rect 1414 1055 1420 1056
rect 1414 1054 1415 1055
rect 1380 1052 1415 1054
rect 1380 1051 1381 1052
rect 1375 1050 1381 1051
rect 1414 1051 1415 1052
rect 1419 1051 1420 1055
rect 1414 1050 1420 1051
rect 1423 1055 1432 1056
rect 1423 1051 1424 1055
rect 1431 1051 1432 1055
rect 1423 1050 1432 1051
rect 1478 1055 1485 1056
rect 1478 1051 1479 1055
rect 1484 1051 1485 1055
rect 1478 1050 1485 1051
rect 1535 1055 1541 1056
rect 1535 1051 1536 1055
rect 1540 1054 1541 1055
rect 1598 1055 1604 1056
rect 1598 1054 1599 1055
rect 1540 1052 1599 1054
rect 1540 1051 1541 1052
rect 1535 1050 1541 1051
rect 1598 1051 1599 1052
rect 1603 1051 1604 1055
rect 1598 1050 1604 1051
rect 1607 1055 1613 1056
rect 1607 1051 1608 1055
rect 1612 1051 1613 1055
rect 1607 1050 1613 1051
rect 1678 1055 1684 1056
rect 1678 1051 1679 1055
rect 1683 1054 1684 1055
rect 1687 1055 1693 1056
rect 1687 1054 1688 1055
rect 1683 1052 1688 1054
rect 1683 1051 1684 1052
rect 1678 1050 1684 1051
rect 1687 1051 1688 1052
rect 1692 1051 1693 1055
rect 1687 1050 1693 1051
rect 1695 1055 1701 1056
rect 1695 1051 1696 1055
rect 1700 1054 1701 1055
rect 1783 1055 1789 1056
rect 1783 1054 1784 1055
rect 1700 1052 1784 1054
rect 1700 1051 1701 1052
rect 1695 1050 1701 1051
rect 1783 1051 1784 1052
rect 1788 1051 1789 1055
rect 1783 1050 1789 1051
rect 1791 1055 1797 1056
rect 1791 1051 1792 1055
rect 1796 1054 1797 1055
rect 1887 1055 1893 1056
rect 1887 1054 1888 1055
rect 1796 1052 1888 1054
rect 1796 1051 1797 1052
rect 1791 1050 1797 1051
rect 1887 1051 1888 1052
rect 1892 1051 1893 1055
rect 1887 1050 1893 1051
rect 1990 1055 1997 1056
rect 1990 1051 1991 1055
rect 1996 1051 1997 1055
rect 1990 1050 1997 1051
rect 2046 1055 2052 1056
rect 2046 1051 2047 1055
rect 2051 1054 2052 1055
rect 2095 1055 2101 1056
rect 2095 1054 2096 1055
rect 2051 1052 2096 1054
rect 2051 1051 2052 1052
rect 2046 1050 2052 1051
rect 2095 1051 2096 1052
rect 2100 1051 2101 1055
rect 2095 1050 2101 1051
rect 2118 1052 2124 1053
rect 1134 1047 1140 1048
rect 2118 1048 2119 1052
rect 2123 1048 2124 1052
rect 2118 1047 2124 1048
rect 1158 1044 1164 1045
rect 159 1043 165 1044
rect 159 1039 160 1043
rect 164 1042 165 1043
rect 190 1043 196 1044
rect 190 1042 191 1043
rect 164 1040 191 1042
rect 164 1039 165 1040
rect 159 1038 165 1039
rect 190 1039 191 1040
rect 195 1039 196 1043
rect 190 1038 196 1039
rect 199 1043 205 1044
rect 199 1039 200 1043
rect 204 1042 205 1043
rect 230 1043 236 1044
rect 230 1042 231 1043
rect 204 1040 231 1042
rect 204 1039 205 1040
rect 199 1038 205 1039
rect 230 1039 231 1040
rect 235 1039 236 1043
rect 230 1038 236 1039
rect 239 1043 245 1044
rect 239 1039 240 1043
rect 244 1042 245 1043
rect 270 1043 276 1044
rect 270 1042 271 1043
rect 244 1040 271 1042
rect 244 1039 245 1040
rect 239 1038 245 1039
rect 270 1039 271 1040
rect 275 1039 276 1043
rect 270 1038 276 1039
rect 279 1043 285 1044
rect 279 1039 280 1043
rect 284 1039 285 1043
rect 279 1038 285 1039
rect 343 1043 349 1044
rect 343 1039 344 1043
rect 348 1042 349 1043
rect 398 1043 404 1044
rect 398 1042 399 1043
rect 348 1040 399 1042
rect 348 1039 349 1040
rect 343 1038 349 1039
rect 398 1039 399 1040
rect 403 1039 404 1043
rect 398 1038 404 1039
rect 407 1043 413 1044
rect 407 1039 408 1043
rect 412 1042 413 1043
rect 462 1043 468 1044
rect 462 1042 463 1043
rect 412 1040 463 1042
rect 412 1039 413 1040
rect 407 1038 413 1039
rect 462 1039 463 1040
rect 467 1039 468 1043
rect 462 1038 468 1039
rect 471 1043 477 1044
rect 471 1039 472 1043
rect 476 1039 477 1043
rect 471 1038 477 1039
rect 535 1043 541 1044
rect 535 1039 536 1043
rect 540 1042 541 1043
rect 546 1043 552 1044
rect 546 1042 547 1043
rect 540 1040 547 1042
rect 540 1039 541 1040
rect 535 1038 541 1039
rect 546 1039 547 1040
rect 551 1039 552 1043
rect 546 1038 552 1039
rect 554 1043 560 1044
rect 554 1039 555 1043
rect 559 1042 560 1043
rect 599 1043 605 1044
rect 599 1042 600 1043
rect 559 1040 600 1042
rect 559 1039 560 1040
rect 554 1038 560 1039
rect 599 1039 600 1040
rect 604 1039 605 1043
rect 599 1038 605 1039
rect 610 1043 616 1044
rect 610 1039 611 1043
rect 615 1042 616 1043
rect 655 1043 661 1044
rect 655 1042 656 1043
rect 615 1040 656 1042
rect 615 1039 616 1040
rect 610 1038 616 1039
rect 655 1039 656 1040
rect 660 1039 661 1043
rect 655 1038 661 1039
rect 663 1043 669 1044
rect 663 1039 664 1043
rect 668 1042 669 1043
rect 711 1043 717 1044
rect 711 1042 712 1043
rect 668 1040 712 1042
rect 668 1039 669 1040
rect 663 1038 669 1039
rect 711 1039 712 1040
rect 716 1039 717 1043
rect 711 1038 717 1039
rect 734 1043 740 1044
rect 734 1039 735 1043
rect 739 1042 740 1043
rect 767 1043 773 1044
rect 767 1042 768 1043
rect 739 1040 768 1042
rect 739 1039 740 1040
rect 734 1038 740 1039
rect 767 1039 768 1040
rect 772 1039 773 1043
rect 767 1038 773 1039
rect 775 1043 781 1044
rect 775 1039 776 1043
rect 780 1042 781 1043
rect 823 1043 829 1044
rect 823 1042 824 1043
rect 780 1040 824 1042
rect 780 1039 781 1040
rect 775 1038 781 1039
rect 823 1039 824 1040
rect 828 1039 829 1043
rect 823 1038 829 1039
rect 831 1043 837 1044
rect 831 1039 832 1043
rect 836 1042 837 1043
rect 887 1043 893 1044
rect 887 1042 888 1043
rect 836 1040 888 1042
rect 836 1039 837 1040
rect 831 1038 837 1039
rect 887 1039 888 1040
rect 892 1039 893 1043
rect 1158 1040 1159 1044
rect 1163 1040 1164 1044
rect 1158 1039 1164 1040
rect 1198 1044 1204 1045
rect 1198 1040 1199 1044
rect 1203 1040 1204 1044
rect 1198 1039 1204 1040
rect 1246 1044 1252 1045
rect 1246 1040 1247 1044
rect 1251 1040 1252 1044
rect 1246 1039 1252 1040
rect 1302 1044 1308 1045
rect 1302 1040 1303 1044
rect 1307 1040 1308 1044
rect 1302 1039 1308 1040
rect 1350 1044 1356 1045
rect 1350 1040 1351 1044
rect 1355 1040 1356 1044
rect 1350 1039 1356 1040
rect 1398 1044 1404 1045
rect 1398 1040 1399 1044
rect 1403 1040 1404 1044
rect 1398 1039 1404 1040
rect 1454 1044 1460 1045
rect 1510 1044 1516 1045
rect 1454 1040 1455 1044
rect 1459 1040 1460 1044
rect 1454 1039 1460 1040
rect 1470 1043 1476 1044
rect 1470 1039 1471 1043
rect 1475 1042 1476 1043
rect 1475 1040 1506 1042
rect 1475 1039 1476 1040
rect 887 1038 893 1039
rect 1470 1038 1476 1039
rect 134 1036 140 1037
rect 134 1032 135 1036
rect 139 1032 140 1036
rect 134 1031 140 1032
rect 174 1036 180 1037
rect 174 1032 175 1036
rect 179 1032 180 1036
rect 174 1031 180 1032
rect 214 1036 220 1037
rect 214 1032 215 1036
rect 219 1032 220 1036
rect 214 1031 220 1032
rect 254 1036 260 1037
rect 254 1032 255 1036
rect 259 1032 260 1036
rect 254 1031 260 1032
rect 318 1036 324 1037
rect 318 1032 319 1036
rect 323 1032 324 1036
rect 318 1031 324 1032
rect 382 1036 388 1037
rect 382 1032 383 1036
rect 387 1032 388 1036
rect 382 1031 388 1032
rect 446 1036 452 1037
rect 446 1032 447 1036
rect 451 1032 452 1036
rect 446 1031 452 1032
rect 510 1036 516 1037
rect 510 1032 511 1036
rect 515 1032 516 1036
rect 510 1031 516 1032
rect 574 1036 580 1037
rect 574 1032 575 1036
rect 579 1032 580 1036
rect 574 1031 580 1032
rect 630 1036 636 1037
rect 630 1032 631 1036
rect 635 1032 636 1036
rect 630 1031 636 1032
rect 686 1036 692 1037
rect 686 1032 687 1036
rect 691 1032 692 1036
rect 686 1031 692 1032
rect 742 1036 748 1037
rect 742 1032 743 1036
rect 747 1032 748 1036
rect 742 1031 748 1032
rect 798 1036 804 1037
rect 798 1032 799 1036
rect 803 1032 804 1036
rect 798 1031 804 1032
rect 862 1036 868 1037
rect 862 1032 863 1036
rect 867 1032 868 1036
rect 862 1031 868 1032
rect 1086 1035 1092 1036
rect 1086 1031 1087 1035
rect 1091 1034 1092 1035
rect 1183 1035 1189 1036
rect 1183 1034 1184 1035
rect 1091 1032 1184 1034
rect 1091 1031 1092 1032
rect 1086 1030 1092 1031
rect 1183 1031 1184 1032
rect 1188 1031 1189 1035
rect 1183 1030 1189 1031
rect 1214 1035 1220 1036
rect 1214 1031 1215 1035
rect 1219 1034 1220 1035
rect 1223 1035 1229 1036
rect 1223 1034 1224 1035
rect 1219 1032 1224 1034
rect 1219 1031 1220 1032
rect 1214 1030 1220 1031
rect 1223 1031 1224 1032
rect 1228 1031 1229 1035
rect 1223 1030 1229 1031
rect 1266 1035 1277 1036
rect 1266 1031 1267 1035
rect 1271 1031 1272 1035
rect 1276 1031 1277 1035
rect 1266 1030 1277 1031
rect 1318 1035 1324 1036
rect 1318 1031 1319 1035
rect 1323 1034 1324 1035
rect 1327 1035 1333 1036
rect 1327 1034 1328 1035
rect 1323 1032 1328 1034
rect 1323 1031 1324 1032
rect 1318 1030 1324 1031
rect 1327 1031 1328 1032
rect 1332 1031 1333 1035
rect 1327 1030 1333 1031
rect 1370 1035 1381 1036
rect 1370 1031 1371 1035
rect 1375 1031 1376 1035
rect 1380 1031 1381 1035
rect 1370 1030 1381 1031
rect 1414 1035 1420 1036
rect 1414 1031 1415 1035
rect 1419 1034 1420 1035
rect 1423 1035 1429 1036
rect 1423 1034 1424 1035
rect 1419 1032 1424 1034
rect 1419 1031 1420 1032
rect 1414 1030 1420 1031
rect 1423 1031 1424 1032
rect 1428 1031 1429 1035
rect 1423 1030 1429 1031
rect 1479 1035 1485 1036
rect 1479 1031 1480 1035
rect 1484 1034 1485 1035
rect 1494 1035 1500 1036
rect 1494 1034 1495 1035
rect 1484 1032 1495 1034
rect 1484 1031 1485 1032
rect 1479 1030 1485 1031
rect 1494 1031 1495 1032
rect 1499 1031 1500 1035
rect 1504 1034 1506 1040
rect 1510 1040 1511 1044
rect 1515 1040 1516 1044
rect 1510 1039 1516 1040
rect 1582 1044 1588 1045
rect 1582 1040 1583 1044
rect 1587 1040 1588 1044
rect 1582 1039 1588 1040
rect 1662 1044 1668 1045
rect 1662 1040 1663 1044
rect 1667 1040 1668 1044
rect 1662 1039 1668 1040
rect 1758 1044 1764 1045
rect 1758 1040 1759 1044
rect 1763 1040 1764 1044
rect 1758 1039 1764 1040
rect 1862 1044 1868 1045
rect 1862 1040 1863 1044
rect 1867 1040 1868 1044
rect 1862 1039 1868 1040
rect 1966 1044 1972 1045
rect 1966 1040 1967 1044
rect 1971 1040 1972 1044
rect 1966 1039 1972 1040
rect 2070 1044 2076 1045
rect 2070 1040 2071 1044
rect 2075 1040 2076 1044
rect 2070 1039 2076 1040
rect 1535 1035 1541 1036
rect 1535 1034 1536 1035
rect 1504 1032 1536 1034
rect 1494 1030 1500 1031
rect 1535 1031 1536 1032
rect 1540 1031 1541 1035
rect 1535 1030 1541 1031
rect 1598 1035 1604 1036
rect 1598 1031 1599 1035
rect 1603 1034 1604 1035
rect 1607 1035 1613 1036
rect 1607 1034 1608 1035
rect 1603 1032 1608 1034
rect 1603 1031 1604 1032
rect 1598 1030 1604 1031
rect 1607 1031 1608 1032
rect 1612 1031 1613 1035
rect 1607 1030 1613 1031
rect 1687 1035 1693 1036
rect 1687 1031 1688 1035
rect 1692 1034 1693 1035
rect 1695 1035 1701 1036
rect 1695 1034 1696 1035
rect 1692 1032 1696 1034
rect 1692 1031 1693 1032
rect 1687 1030 1693 1031
rect 1695 1031 1696 1032
rect 1700 1031 1701 1035
rect 1695 1030 1701 1031
rect 1783 1035 1789 1036
rect 1783 1031 1784 1035
rect 1788 1034 1789 1035
rect 1791 1035 1797 1036
rect 1791 1034 1792 1035
rect 1788 1032 1792 1034
rect 1788 1031 1789 1032
rect 1783 1030 1789 1031
rect 1791 1031 1792 1032
rect 1796 1031 1797 1035
rect 1791 1030 1797 1031
rect 1886 1035 1893 1036
rect 1886 1031 1887 1035
rect 1892 1031 1893 1035
rect 1886 1030 1893 1031
rect 1991 1035 1997 1036
rect 1991 1031 1992 1035
rect 1996 1034 1997 1035
rect 2046 1035 2052 1036
rect 2046 1034 2047 1035
rect 1996 1032 2047 1034
rect 1996 1031 1997 1032
rect 1991 1030 1997 1031
rect 2046 1031 2047 1032
rect 2051 1031 2052 1035
rect 2046 1030 2052 1031
rect 2094 1035 2101 1036
rect 2094 1031 2095 1035
rect 2100 1031 2101 1035
rect 2094 1030 2101 1031
rect 110 1028 116 1029
rect 110 1024 111 1028
rect 115 1024 116 1028
rect 1094 1028 1100 1029
rect 1094 1024 1095 1028
rect 1099 1024 1100 1028
rect 110 1023 116 1024
rect 159 1023 165 1024
rect 159 1019 160 1023
rect 164 1019 165 1023
rect 159 1018 165 1019
rect 190 1023 196 1024
rect 190 1019 191 1023
rect 195 1022 196 1023
rect 199 1023 205 1024
rect 199 1022 200 1023
rect 195 1020 200 1022
rect 195 1019 196 1020
rect 190 1018 196 1019
rect 199 1019 200 1020
rect 204 1019 205 1023
rect 199 1018 205 1019
rect 230 1023 236 1024
rect 230 1019 231 1023
rect 235 1022 236 1023
rect 239 1023 245 1024
rect 239 1022 240 1023
rect 235 1020 240 1022
rect 235 1019 236 1020
rect 230 1018 236 1019
rect 239 1019 240 1020
rect 244 1019 245 1023
rect 239 1018 245 1019
rect 270 1023 276 1024
rect 270 1019 271 1023
rect 275 1022 276 1023
rect 279 1023 285 1024
rect 279 1022 280 1023
rect 275 1020 280 1022
rect 275 1019 276 1020
rect 270 1018 276 1019
rect 279 1019 280 1020
rect 284 1019 285 1023
rect 279 1018 285 1019
rect 290 1023 296 1024
rect 290 1019 291 1023
rect 295 1022 296 1023
rect 343 1023 349 1024
rect 343 1022 344 1023
rect 295 1020 344 1022
rect 295 1019 296 1020
rect 290 1018 296 1019
rect 343 1019 344 1020
rect 348 1019 349 1023
rect 343 1018 349 1019
rect 398 1023 404 1024
rect 398 1019 399 1023
rect 403 1022 404 1023
rect 407 1023 413 1024
rect 407 1022 408 1023
rect 403 1020 408 1022
rect 403 1019 404 1020
rect 398 1018 404 1019
rect 407 1019 408 1020
rect 412 1019 413 1023
rect 407 1018 413 1019
rect 462 1023 468 1024
rect 462 1019 463 1023
rect 467 1022 468 1023
rect 471 1023 477 1024
rect 471 1022 472 1023
rect 467 1020 472 1022
rect 467 1019 468 1020
rect 462 1018 468 1019
rect 471 1019 472 1020
rect 476 1019 477 1023
rect 471 1018 477 1019
rect 535 1023 541 1024
rect 535 1019 536 1023
rect 540 1022 541 1023
rect 554 1023 560 1024
rect 554 1022 555 1023
rect 540 1020 555 1022
rect 540 1019 541 1020
rect 535 1018 541 1019
rect 554 1019 555 1020
rect 559 1019 560 1023
rect 554 1018 560 1019
rect 599 1023 608 1024
rect 599 1019 600 1023
rect 607 1019 608 1023
rect 599 1018 608 1019
rect 655 1023 661 1024
rect 655 1019 656 1023
rect 660 1022 661 1023
rect 663 1023 669 1024
rect 663 1022 664 1023
rect 660 1020 664 1022
rect 660 1019 661 1020
rect 655 1018 661 1019
rect 663 1019 664 1020
rect 668 1019 669 1023
rect 663 1018 669 1019
rect 711 1023 717 1024
rect 711 1019 712 1023
rect 716 1022 717 1023
rect 734 1023 740 1024
rect 734 1022 735 1023
rect 716 1020 735 1022
rect 716 1019 717 1020
rect 711 1018 717 1019
rect 734 1019 735 1020
rect 739 1019 740 1023
rect 734 1018 740 1019
rect 767 1023 773 1024
rect 767 1019 768 1023
rect 772 1022 773 1023
rect 775 1023 781 1024
rect 775 1022 776 1023
rect 772 1020 776 1022
rect 772 1019 773 1020
rect 767 1018 773 1019
rect 775 1019 776 1020
rect 780 1019 781 1023
rect 775 1018 781 1019
rect 823 1023 829 1024
rect 823 1019 824 1023
rect 828 1022 829 1023
rect 831 1023 837 1024
rect 831 1022 832 1023
rect 828 1020 832 1022
rect 828 1019 829 1020
rect 823 1018 829 1019
rect 831 1019 832 1020
rect 836 1019 837 1023
rect 831 1018 837 1019
rect 882 1023 893 1024
rect 1094 1023 1100 1024
rect 882 1019 883 1023
rect 887 1019 888 1023
rect 892 1019 893 1023
rect 882 1018 893 1019
rect 1743 1019 1749 1020
rect 1678 1015 1684 1016
rect 1678 1014 1679 1015
rect 1663 1013 1679 1014
rect 110 1011 116 1012
rect 110 1007 111 1011
rect 115 1007 116 1011
rect 1094 1011 1100 1012
rect 110 1006 116 1007
rect 134 1008 140 1009
rect 134 1004 135 1008
rect 139 1004 140 1008
rect 134 1003 140 1004
rect 174 1008 180 1009
rect 174 1004 175 1008
rect 179 1004 180 1008
rect 174 1003 180 1004
rect 214 1008 220 1009
rect 214 1004 215 1008
rect 219 1004 220 1008
rect 214 1003 220 1004
rect 254 1008 260 1009
rect 254 1004 255 1008
rect 259 1004 260 1008
rect 254 1003 260 1004
rect 318 1008 324 1009
rect 318 1004 319 1008
rect 323 1004 324 1008
rect 318 1003 324 1004
rect 382 1008 388 1009
rect 382 1004 383 1008
rect 387 1004 388 1008
rect 382 1003 388 1004
rect 446 1008 452 1009
rect 446 1004 447 1008
rect 451 1004 452 1008
rect 446 1003 452 1004
rect 510 1008 516 1009
rect 510 1004 511 1008
rect 515 1004 516 1008
rect 510 1003 516 1004
rect 574 1008 580 1009
rect 574 1004 575 1008
rect 579 1004 580 1008
rect 574 1003 580 1004
rect 630 1008 636 1009
rect 630 1004 631 1008
rect 635 1004 636 1008
rect 630 1003 636 1004
rect 686 1008 692 1009
rect 686 1004 687 1008
rect 691 1004 692 1008
rect 686 1003 692 1004
rect 742 1008 748 1009
rect 742 1004 743 1008
rect 747 1004 748 1008
rect 742 1003 748 1004
rect 798 1008 804 1009
rect 798 1004 799 1008
rect 803 1004 804 1008
rect 798 1003 804 1004
rect 862 1008 868 1009
rect 862 1004 863 1008
rect 867 1004 868 1008
rect 1094 1007 1095 1011
rect 1099 1007 1100 1011
rect 1094 1006 1100 1007
rect 1183 1011 1189 1012
rect 1183 1007 1184 1011
rect 1188 1010 1189 1011
rect 1214 1011 1220 1012
rect 1214 1010 1215 1011
rect 1188 1008 1215 1010
rect 1188 1007 1189 1008
rect 1183 1006 1189 1007
rect 1214 1007 1215 1008
rect 1219 1007 1220 1011
rect 1214 1006 1220 1007
rect 1222 1011 1229 1012
rect 1222 1007 1223 1011
rect 1228 1007 1229 1011
rect 1222 1006 1229 1007
rect 1263 1011 1269 1012
rect 1263 1007 1264 1011
rect 1268 1010 1269 1011
rect 1310 1011 1316 1012
rect 1310 1010 1311 1011
rect 1268 1008 1311 1010
rect 1268 1007 1269 1008
rect 1263 1006 1269 1007
rect 1310 1007 1311 1008
rect 1315 1007 1316 1011
rect 1310 1006 1316 1007
rect 1319 1011 1325 1012
rect 1319 1007 1320 1011
rect 1324 1010 1325 1011
rect 1358 1011 1364 1012
rect 1358 1010 1359 1011
rect 1324 1008 1359 1010
rect 1324 1007 1325 1008
rect 1319 1006 1325 1007
rect 1358 1007 1359 1008
rect 1363 1007 1364 1011
rect 1358 1006 1364 1007
rect 1375 1011 1381 1012
rect 1375 1007 1376 1011
rect 1380 1010 1381 1011
rect 1398 1011 1404 1012
rect 1398 1010 1399 1011
rect 1380 1008 1399 1010
rect 1380 1007 1381 1008
rect 1375 1006 1381 1007
rect 1398 1007 1399 1008
rect 1403 1007 1404 1011
rect 1398 1006 1404 1007
rect 1426 1011 1437 1012
rect 1426 1007 1427 1011
rect 1431 1007 1432 1011
rect 1436 1007 1437 1011
rect 1426 1006 1437 1007
rect 1439 1011 1445 1012
rect 1439 1007 1440 1011
rect 1444 1010 1445 1011
rect 1487 1011 1493 1012
rect 1487 1010 1488 1011
rect 1444 1008 1488 1010
rect 1444 1007 1445 1008
rect 1439 1006 1445 1007
rect 1487 1007 1488 1008
rect 1492 1007 1493 1011
rect 1487 1006 1493 1007
rect 1543 1011 1549 1012
rect 1543 1007 1544 1011
rect 1548 1010 1549 1011
rect 1590 1011 1596 1012
rect 1590 1010 1591 1011
rect 1548 1008 1591 1010
rect 1548 1007 1549 1008
rect 1543 1006 1549 1007
rect 1590 1007 1591 1008
rect 1595 1007 1596 1011
rect 1590 1006 1596 1007
rect 1599 1011 1605 1012
rect 1599 1007 1600 1011
rect 1604 1010 1605 1011
rect 1654 1011 1660 1012
rect 1654 1010 1655 1011
rect 1604 1008 1655 1010
rect 1604 1007 1605 1008
rect 1599 1006 1605 1007
rect 1654 1007 1655 1008
rect 1659 1007 1660 1011
rect 1663 1009 1664 1013
rect 1668 1012 1679 1013
rect 1668 1009 1669 1012
rect 1678 1011 1679 1012
rect 1683 1011 1684 1015
rect 1743 1015 1744 1019
rect 1748 1018 1749 1019
rect 1990 1019 1996 1020
rect 1748 1016 1906 1018
rect 1748 1015 1749 1016
rect 1743 1014 1749 1015
rect 1904 1012 1906 1016
rect 1990 1015 1991 1019
rect 1995 1018 1996 1019
rect 1995 1016 2001 1018
rect 1995 1015 1996 1016
rect 1990 1014 1996 1015
rect 1999 1014 2001 1016
rect 1999 1012 2046 1014
rect 1678 1010 1684 1011
rect 1735 1011 1741 1012
rect 1735 1010 1736 1011
rect 1663 1008 1669 1009
rect 1688 1008 1736 1010
rect 1654 1006 1660 1007
rect 862 1003 868 1004
rect 1158 1004 1164 1005
rect 1158 1000 1159 1004
rect 1163 1000 1164 1004
rect 1158 999 1164 1000
rect 1198 1004 1204 1005
rect 1198 1000 1199 1004
rect 1203 1000 1204 1004
rect 1198 999 1204 1000
rect 1238 1004 1244 1005
rect 1238 1000 1239 1004
rect 1243 1000 1244 1004
rect 1238 999 1244 1000
rect 1294 1004 1300 1005
rect 1294 1000 1295 1004
rect 1299 1000 1300 1004
rect 1294 999 1300 1000
rect 1350 1004 1356 1005
rect 1350 1000 1351 1004
rect 1355 1000 1356 1004
rect 1350 999 1356 1000
rect 1406 1004 1412 1005
rect 1406 1000 1407 1004
rect 1411 1000 1412 1004
rect 1406 999 1412 1000
rect 1462 1004 1468 1005
rect 1462 1000 1463 1004
rect 1467 1000 1468 1004
rect 1462 999 1468 1000
rect 1518 1004 1524 1005
rect 1518 1000 1519 1004
rect 1523 1000 1524 1004
rect 1518 999 1524 1000
rect 1574 1004 1580 1005
rect 1574 1000 1575 1004
rect 1579 1000 1580 1004
rect 1574 999 1580 1000
rect 1638 1004 1644 1005
rect 1638 1000 1639 1004
rect 1643 1000 1644 1004
rect 1688 1002 1690 1008
rect 1735 1007 1736 1008
rect 1740 1007 1741 1011
rect 1735 1006 1741 1007
rect 1815 1011 1821 1012
rect 1815 1007 1816 1011
rect 1820 1010 1821 1011
rect 1894 1011 1900 1012
rect 1894 1010 1895 1011
rect 1820 1008 1895 1010
rect 1820 1007 1821 1008
rect 1815 1006 1821 1007
rect 1894 1007 1895 1008
rect 1899 1007 1900 1011
rect 1894 1006 1900 1007
rect 1903 1011 1909 1012
rect 1903 1007 1904 1011
rect 1908 1007 1909 1011
rect 1903 1006 1909 1007
rect 1991 1011 1997 1012
rect 1991 1007 1992 1011
rect 1996 1010 1997 1011
rect 2044 1010 2046 1012
rect 2087 1011 2093 1012
rect 2087 1010 2088 1011
rect 1996 1008 2001 1010
rect 2044 1008 2088 1010
rect 1996 1007 1997 1008
rect 1991 1006 1997 1007
rect 1638 999 1644 1000
rect 1648 1000 1690 1002
rect 1710 1004 1716 1005
rect 1710 1000 1711 1004
rect 1715 1000 1716 1004
rect 1134 996 1140 997
rect 134 992 140 993
rect 110 989 116 990
rect 110 985 111 989
rect 115 985 116 989
rect 134 988 135 992
rect 139 988 140 992
rect 134 987 140 988
rect 174 992 180 993
rect 174 988 175 992
rect 179 988 180 992
rect 174 987 180 988
rect 222 992 228 993
rect 222 988 223 992
rect 227 988 228 992
rect 222 987 228 988
rect 278 992 284 993
rect 278 988 279 992
rect 283 988 284 992
rect 278 987 284 988
rect 342 992 348 993
rect 342 988 343 992
rect 347 988 348 992
rect 342 987 348 988
rect 406 992 412 993
rect 406 988 407 992
rect 411 988 412 992
rect 406 987 412 988
rect 470 992 476 993
rect 470 988 471 992
rect 475 988 476 992
rect 470 987 476 988
rect 526 992 532 993
rect 526 988 527 992
rect 531 988 532 992
rect 526 987 532 988
rect 582 992 588 993
rect 582 988 583 992
rect 587 988 588 992
rect 582 987 588 988
rect 630 992 636 993
rect 630 988 631 992
rect 635 988 636 992
rect 630 987 636 988
rect 686 992 692 993
rect 686 988 687 992
rect 691 988 692 992
rect 686 987 692 988
rect 742 992 748 993
rect 742 988 743 992
rect 747 988 748 992
rect 742 987 748 988
rect 798 992 804 993
rect 798 988 799 992
rect 803 988 804 992
rect 1134 992 1135 996
rect 1139 992 1140 996
rect 1585 996 1610 998
rect 1134 991 1140 992
rect 1183 991 1189 992
rect 798 987 804 988
rect 1094 989 1100 990
rect 110 984 116 985
rect 1094 985 1095 989
rect 1099 985 1100 989
rect 1183 987 1184 991
rect 1188 990 1189 991
rect 1206 991 1212 992
rect 1206 990 1207 991
rect 1188 988 1207 990
rect 1188 987 1189 988
rect 1183 986 1189 987
rect 1206 987 1207 988
rect 1211 987 1212 991
rect 1206 986 1212 987
rect 1214 991 1220 992
rect 1214 987 1215 991
rect 1219 990 1220 991
rect 1223 991 1229 992
rect 1223 990 1224 991
rect 1219 988 1224 990
rect 1219 987 1220 988
rect 1214 986 1220 987
rect 1223 987 1224 988
rect 1228 987 1229 991
rect 1223 986 1229 987
rect 1263 991 1272 992
rect 1263 987 1264 991
rect 1271 987 1272 991
rect 1263 986 1272 987
rect 1310 991 1316 992
rect 1310 987 1311 991
rect 1315 990 1316 991
rect 1319 991 1325 992
rect 1319 990 1320 991
rect 1315 988 1320 990
rect 1315 987 1316 988
rect 1310 986 1316 987
rect 1319 987 1320 988
rect 1324 987 1325 991
rect 1319 986 1325 987
rect 1358 991 1364 992
rect 1358 987 1359 991
rect 1363 990 1364 991
rect 1375 991 1381 992
rect 1375 990 1376 991
rect 1363 988 1376 990
rect 1363 987 1364 988
rect 1358 986 1364 987
rect 1375 987 1376 988
rect 1380 987 1381 991
rect 1375 986 1381 987
rect 1431 991 1437 992
rect 1431 987 1432 991
rect 1436 990 1437 991
rect 1439 991 1445 992
rect 1439 990 1440 991
rect 1436 988 1440 990
rect 1436 987 1437 988
rect 1431 986 1437 987
rect 1439 987 1440 988
rect 1444 987 1445 991
rect 1439 986 1445 987
rect 1482 991 1493 992
rect 1482 987 1483 991
rect 1487 987 1488 991
rect 1492 987 1493 991
rect 1482 986 1493 987
rect 1543 991 1549 992
rect 1543 987 1544 991
rect 1548 990 1549 991
rect 1585 990 1587 996
rect 1608 994 1610 996
rect 1648 994 1650 1000
rect 1710 999 1716 1000
rect 1790 1004 1796 1005
rect 1790 1000 1791 1004
rect 1795 1000 1796 1004
rect 1790 999 1796 1000
rect 1878 1004 1884 1005
rect 1878 1000 1879 1004
rect 1883 1000 1884 1004
rect 1878 999 1884 1000
rect 1966 1004 1972 1005
rect 1966 1000 1967 1004
rect 1971 1000 1972 1004
rect 1966 999 1972 1000
rect 1608 992 1650 994
rect 1548 988 1587 990
rect 1590 991 1596 992
rect 1548 987 1549 988
rect 1543 986 1549 987
rect 1590 987 1591 991
rect 1595 990 1596 991
rect 1599 991 1605 992
rect 1599 990 1600 991
rect 1595 988 1600 990
rect 1595 987 1596 988
rect 1590 986 1596 987
rect 1599 987 1600 988
rect 1604 987 1605 991
rect 1599 986 1605 987
rect 1654 991 1660 992
rect 1654 987 1655 991
rect 1659 990 1660 991
rect 1663 991 1669 992
rect 1663 990 1664 991
rect 1659 988 1664 990
rect 1659 987 1660 988
rect 1654 986 1660 987
rect 1663 987 1664 988
rect 1668 987 1669 991
rect 1663 986 1669 987
rect 1735 991 1741 992
rect 1735 987 1736 991
rect 1740 990 1741 991
rect 1743 991 1749 992
rect 1743 990 1744 991
rect 1740 988 1744 990
rect 1740 987 1741 988
rect 1735 986 1741 987
rect 1743 987 1744 988
rect 1748 987 1749 991
rect 1743 986 1749 987
rect 1778 991 1784 992
rect 1778 987 1779 991
rect 1783 990 1784 991
rect 1815 991 1821 992
rect 1815 990 1816 991
rect 1783 988 1816 990
rect 1783 987 1784 988
rect 1778 986 1784 987
rect 1815 987 1816 988
rect 1820 987 1821 991
rect 1815 986 1821 987
rect 1894 991 1900 992
rect 1894 987 1895 991
rect 1899 990 1900 991
rect 1903 991 1909 992
rect 1903 990 1904 991
rect 1899 988 1904 990
rect 1899 987 1900 988
rect 1894 986 1900 987
rect 1903 987 1904 988
rect 1908 987 1909 991
rect 1903 986 1909 987
rect 1982 991 1988 992
rect 1982 987 1983 991
rect 1987 990 1988 991
rect 1991 991 1997 992
rect 1991 990 1992 991
rect 1987 988 1992 990
rect 1987 987 1988 988
rect 1982 986 1988 987
rect 1991 987 1992 988
rect 1996 987 1997 991
rect 1999 990 2001 1008
rect 2087 1007 2088 1008
rect 2092 1007 2093 1011
rect 2087 1006 2093 1007
rect 2062 1004 2068 1005
rect 2062 1000 2063 1004
rect 2067 1000 2068 1004
rect 2062 999 2068 1000
rect 2118 996 2124 997
rect 2118 992 2119 996
rect 2123 992 2124 996
rect 2087 991 2093 992
rect 2118 991 2124 992
rect 2087 990 2088 991
rect 1999 988 2088 990
rect 1991 986 1997 987
rect 2087 987 2088 988
rect 2092 987 2093 991
rect 2087 986 2093 987
rect 1094 984 1100 985
rect 302 983 308 984
rect 302 982 303 983
rect 176 980 303 982
rect 159 975 165 976
rect 110 972 116 973
rect 110 968 111 972
rect 115 968 116 972
rect 159 971 160 975
rect 164 974 165 975
rect 176 974 178 980
rect 302 979 303 980
rect 307 979 308 983
rect 302 978 308 979
rect 1134 979 1140 980
rect 164 972 178 974
rect 182 975 188 976
rect 164 971 165 972
rect 159 970 165 971
rect 182 971 183 975
rect 187 974 188 975
rect 199 975 205 976
rect 199 974 200 975
rect 187 972 200 974
rect 187 971 188 972
rect 182 970 188 971
rect 199 971 200 972
rect 204 971 205 975
rect 199 970 205 971
rect 207 975 213 976
rect 207 971 208 975
rect 212 974 213 975
rect 247 975 253 976
rect 247 974 248 975
rect 212 972 248 974
rect 212 971 213 972
rect 207 970 213 971
rect 247 971 248 972
rect 252 971 253 975
rect 247 970 253 971
rect 303 975 309 976
rect 303 971 304 975
rect 308 974 309 975
rect 358 975 364 976
rect 358 974 359 975
rect 308 972 359 974
rect 308 971 309 972
rect 303 970 309 971
rect 358 971 359 972
rect 363 971 364 975
rect 358 970 364 971
rect 367 975 373 976
rect 367 971 368 975
rect 372 974 373 975
rect 418 975 424 976
rect 418 974 419 975
rect 372 972 419 974
rect 372 971 373 972
rect 367 970 373 971
rect 418 971 419 972
rect 423 971 424 975
rect 418 970 424 971
rect 426 975 437 976
rect 426 971 427 975
rect 431 971 432 975
rect 436 971 437 975
rect 426 970 437 971
rect 495 975 501 976
rect 495 971 496 975
rect 500 974 501 975
rect 538 975 544 976
rect 538 974 539 975
rect 500 972 539 974
rect 500 971 501 972
rect 495 970 501 971
rect 538 971 539 972
rect 543 971 544 975
rect 538 970 544 971
rect 546 975 557 976
rect 546 971 547 975
rect 551 971 552 975
rect 556 971 557 975
rect 546 970 557 971
rect 606 975 613 976
rect 606 971 607 975
rect 612 971 613 975
rect 606 970 613 971
rect 615 975 621 976
rect 615 971 616 975
rect 620 974 621 975
rect 655 975 661 976
rect 655 974 656 975
rect 620 972 656 974
rect 620 971 621 972
rect 615 970 621 971
rect 655 971 656 972
rect 660 971 661 975
rect 655 970 661 971
rect 663 975 669 976
rect 663 971 664 975
rect 668 974 669 975
rect 711 975 717 976
rect 711 974 712 975
rect 668 972 712 974
rect 668 971 669 972
rect 663 970 669 971
rect 711 971 712 972
rect 716 971 717 975
rect 711 970 717 971
rect 719 975 725 976
rect 719 971 720 975
rect 724 974 725 975
rect 767 975 773 976
rect 767 974 768 975
rect 724 972 768 974
rect 724 971 725 972
rect 719 970 725 971
rect 767 971 768 972
rect 772 971 773 975
rect 767 970 773 971
rect 775 975 781 976
rect 775 971 776 975
rect 780 974 781 975
rect 823 975 829 976
rect 823 974 824 975
rect 780 972 824 974
rect 780 971 781 972
rect 775 970 781 971
rect 823 971 824 972
rect 828 971 829 975
rect 1134 975 1135 979
rect 1139 975 1140 979
rect 2118 979 2124 980
rect 1134 974 1140 975
rect 1158 976 1164 977
rect 823 970 829 971
rect 1094 972 1100 973
rect 110 967 116 968
rect 1094 968 1095 972
rect 1099 968 1100 972
rect 1158 972 1159 976
rect 1163 972 1164 976
rect 1158 971 1164 972
rect 1198 976 1204 977
rect 1198 972 1199 976
rect 1203 972 1204 976
rect 1198 971 1204 972
rect 1238 976 1244 977
rect 1238 972 1239 976
rect 1243 972 1244 976
rect 1238 971 1244 972
rect 1294 976 1300 977
rect 1294 972 1295 976
rect 1299 972 1300 976
rect 1294 971 1300 972
rect 1350 976 1356 977
rect 1350 972 1351 976
rect 1355 972 1356 976
rect 1350 971 1356 972
rect 1406 976 1412 977
rect 1406 972 1407 976
rect 1411 972 1412 976
rect 1406 971 1412 972
rect 1462 976 1468 977
rect 1462 972 1463 976
rect 1467 972 1468 976
rect 1462 971 1468 972
rect 1518 976 1524 977
rect 1518 972 1519 976
rect 1523 972 1524 976
rect 1518 971 1524 972
rect 1574 976 1580 977
rect 1574 972 1575 976
rect 1579 972 1580 976
rect 1574 971 1580 972
rect 1638 976 1644 977
rect 1638 972 1639 976
rect 1643 972 1644 976
rect 1638 971 1644 972
rect 1710 976 1716 977
rect 1710 972 1711 976
rect 1715 972 1716 976
rect 1710 971 1716 972
rect 1790 976 1796 977
rect 1790 972 1791 976
rect 1795 972 1796 976
rect 1790 971 1796 972
rect 1878 976 1884 977
rect 1878 972 1879 976
rect 1883 972 1884 976
rect 1878 971 1884 972
rect 1966 976 1972 977
rect 1966 972 1967 976
rect 1971 972 1972 976
rect 1966 971 1972 972
rect 2062 976 2068 977
rect 2062 972 2063 976
rect 2067 972 2068 976
rect 2118 975 2119 979
rect 2123 975 2124 979
rect 2118 974 2124 975
rect 2062 971 2068 972
rect 1094 967 1100 968
rect 134 964 140 965
rect 134 960 135 964
rect 139 960 140 964
rect 134 959 140 960
rect 174 964 180 965
rect 174 960 175 964
rect 179 960 180 964
rect 174 959 180 960
rect 222 964 228 965
rect 222 960 223 964
rect 227 960 228 964
rect 222 959 228 960
rect 278 964 284 965
rect 278 960 279 964
rect 283 960 284 964
rect 278 959 284 960
rect 342 964 348 965
rect 342 960 343 964
rect 347 960 348 964
rect 342 959 348 960
rect 406 964 412 965
rect 406 960 407 964
rect 411 960 412 964
rect 406 959 412 960
rect 470 964 476 965
rect 470 960 471 964
rect 475 960 476 964
rect 470 959 476 960
rect 526 964 532 965
rect 526 960 527 964
rect 531 960 532 964
rect 526 959 532 960
rect 582 964 588 965
rect 582 960 583 964
rect 587 960 588 964
rect 582 959 588 960
rect 630 964 636 965
rect 630 960 631 964
rect 635 960 636 964
rect 630 959 636 960
rect 686 964 692 965
rect 686 960 687 964
rect 691 960 692 964
rect 686 959 692 960
rect 742 964 748 965
rect 742 960 743 964
rect 747 960 748 964
rect 742 959 748 960
rect 798 964 804 965
rect 798 960 799 964
rect 803 960 804 964
rect 798 959 804 960
rect 1158 956 1164 957
rect 159 955 165 956
rect 159 951 160 955
rect 164 954 165 955
rect 182 955 188 956
rect 182 954 183 955
rect 164 952 183 954
rect 164 951 165 952
rect 159 950 165 951
rect 182 951 183 952
rect 187 951 188 955
rect 182 950 188 951
rect 199 955 205 956
rect 199 951 200 955
rect 204 954 205 955
rect 207 955 213 956
rect 207 954 208 955
rect 204 952 208 954
rect 204 951 205 952
rect 199 950 205 951
rect 207 951 208 952
rect 212 951 213 955
rect 207 950 213 951
rect 247 955 253 956
rect 247 951 248 955
rect 252 954 253 955
rect 290 955 296 956
rect 290 954 291 955
rect 252 952 291 954
rect 252 951 253 952
rect 247 950 253 951
rect 290 951 291 952
rect 295 951 296 955
rect 290 950 296 951
rect 302 955 309 956
rect 302 951 303 955
rect 308 951 309 955
rect 302 950 309 951
rect 358 955 364 956
rect 358 951 359 955
rect 363 954 364 955
rect 367 955 373 956
rect 367 954 368 955
rect 363 952 368 954
rect 363 951 364 952
rect 358 950 364 951
rect 367 951 368 952
rect 372 951 373 955
rect 367 950 373 951
rect 418 955 424 956
rect 418 951 419 955
rect 423 954 424 955
rect 431 955 437 956
rect 431 954 432 955
rect 423 952 432 954
rect 423 951 424 952
rect 418 950 424 951
rect 431 951 432 952
rect 436 951 437 955
rect 431 950 437 951
rect 482 955 488 956
rect 482 951 483 955
rect 487 954 488 955
rect 495 955 501 956
rect 495 954 496 955
rect 487 952 496 954
rect 487 951 488 952
rect 482 950 488 951
rect 495 951 496 952
rect 500 951 501 955
rect 495 950 501 951
rect 538 955 544 956
rect 538 951 539 955
rect 543 954 544 955
rect 551 955 557 956
rect 551 954 552 955
rect 543 952 552 954
rect 543 951 544 952
rect 538 950 544 951
rect 551 951 552 952
rect 556 951 557 955
rect 551 950 557 951
rect 607 955 613 956
rect 607 951 608 955
rect 612 954 613 955
rect 615 955 621 956
rect 615 954 616 955
rect 612 952 616 954
rect 612 951 613 952
rect 607 950 613 951
rect 615 951 616 952
rect 620 951 621 955
rect 615 950 621 951
rect 655 955 661 956
rect 655 951 656 955
rect 660 954 661 955
rect 663 955 669 956
rect 663 954 664 955
rect 660 952 664 954
rect 660 951 661 952
rect 655 950 661 951
rect 663 951 664 952
rect 668 951 669 955
rect 663 950 669 951
rect 711 955 717 956
rect 711 951 712 955
rect 716 954 717 955
rect 719 955 725 956
rect 719 954 720 955
rect 716 952 720 954
rect 716 951 717 952
rect 711 950 717 951
rect 719 951 720 952
rect 724 951 725 955
rect 719 950 725 951
rect 767 955 773 956
rect 767 951 768 955
rect 772 954 773 955
rect 775 955 781 956
rect 775 954 776 955
rect 772 952 776 954
rect 772 951 773 952
rect 767 950 773 951
rect 775 951 776 952
rect 780 951 781 955
rect 823 955 829 956
rect 823 954 824 955
rect 775 950 781 951
rect 784 952 824 954
rect 714 947 720 948
rect 714 943 715 947
rect 719 946 720 947
rect 784 946 786 952
rect 823 951 824 952
rect 828 951 829 955
rect 823 950 829 951
rect 1134 953 1140 954
rect 1134 949 1135 953
rect 1139 949 1140 953
rect 1158 952 1159 956
rect 1163 952 1164 956
rect 1158 951 1164 952
rect 1206 956 1212 957
rect 1206 952 1207 956
rect 1211 952 1212 956
rect 1206 951 1212 952
rect 1286 956 1292 957
rect 1286 952 1287 956
rect 1291 952 1292 956
rect 1286 951 1292 952
rect 1374 956 1380 957
rect 1374 952 1375 956
rect 1379 952 1380 956
rect 1374 951 1380 952
rect 1454 956 1460 957
rect 1454 952 1455 956
rect 1459 952 1460 956
rect 1454 951 1460 952
rect 1534 956 1540 957
rect 1534 952 1535 956
rect 1539 952 1540 956
rect 1534 951 1540 952
rect 1614 956 1620 957
rect 1614 952 1615 956
rect 1619 952 1620 956
rect 1614 951 1620 952
rect 1686 956 1692 957
rect 1686 952 1687 956
rect 1691 952 1692 956
rect 1686 951 1692 952
rect 1750 956 1756 957
rect 1750 952 1751 956
rect 1755 952 1756 956
rect 1750 951 1756 952
rect 1814 956 1820 957
rect 1814 952 1815 956
rect 1819 952 1820 956
rect 1814 951 1820 952
rect 1878 956 1884 957
rect 1878 952 1879 956
rect 1883 952 1884 956
rect 1878 951 1884 952
rect 1950 956 1956 957
rect 1950 952 1951 956
rect 1955 952 1956 956
rect 1950 951 1956 952
rect 2022 956 2028 957
rect 2022 952 2023 956
rect 2027 952 2028 956
rect 2022 951 2028 952
rect 2070 956 2076 957
rect 2070 952 2071 956
rect 2075 952 2076 956
rect 2070 951 2076 952
rect 2118 953 2124 954
rect 1134 948 1140 949
rect 2118 949 2119 953
rect 2123 949 2124 953
rect 2118 948 2124 949
rect 1838 947 1844 948
rect 1838 946 1839 947
rect 719 944 786 946
rect 1640 944 1839 946
rect 719 943 720 944
rect 714 942 720 943
rect 1073 940 1187 942
rect 1640 940 1642 944
rect 1838 943 1839 944
rect 1843 943 1844 947
rect 1838 942 1844 943
rect 1073 932 1075 940
rect 1183 939 1189 940
rect 1134 936 1140 937
rect 1134 932 1135 936
rect 1139 932 1140 936
rect 1183 935 1184 939
rect 1188 935 1189 939
rect 1183 934 1189 935
rect 1214 939 1220 940
rect 1214 935 1215 939
rect 1219 938 1220 939
rect 1231 939 1237 940
rect 1231 938 1232 939
rect 1219 936 1232 938
rect 1219 935 1220 936
rect 1214 934 1220 935
rect 1231 935 1232 936
rect 1236 935 1237 939
rect 1231 934 1237 935
rect 1311 939 1317 940
rect 1311 935 1312 939
rect 1316 938 1317 939
rect 1390 939 1396 940
rect 1390 938 1391 939
rect 1316 936 1391 938
rect 1316 935 1317 936
rect 1311 934 1317 935
rect 1390 935 1391 936
rect 1395 935 1396 939
rect 1390 934 1396 935
rect 1398 939 1405 940
rect 1398 935 1399 939
rect 1404 935 1405 939
rect 1398 934 1405 935
rect 1479 939 1485 940
rect 1479 935 1480 939
rect 1484 938 1485 939
rect 1550 939 1556 940
rect 1550 938 1551 939
rect 1484 936 1551 938
rect 1484 935 1485 936
rect 1479 934 1485 935
rect 1550 935 1551 936
rect 1555 935 1556 939
rect 1550 934 1556 935
rect 1559 939 1565 940
rect 1559 935 1560 939
rect 1564 938 1565 939
rect 1606 939 1612 940
rect 1606 938 1607 939
rect 1564 936 1607 938
rect 1564 935 1565 936
rect 1559 934 1565 935
rect 1606 935 1607 936
rect 1611 935 1612 939
rect 1606 934 1612 935
rect 1639 939 1645 940
rect 1639 935 1640 939
rect 1644 935 1645 939
rect 1639 934 1645 935
rect 1647 939 1653 940
rect 1647 935 1648 939
rect 1652 938 1653 939
rect 1711 939 1717 940
rect 1711 938 1712 939
rect 1652 936 1712 938
rect 1652 935 1653 936
rect 1647 934 1653 935
rect 1711 935 1712 936
rect 1716 935 1717 939
rect 1711 934 1717 935
rect 1719 939 1725 940
rect 1719 935 1720 939
rect 1724 938 1725 939
rect 1775 939 1781 940
rect 1775 938 1776 939
rect 1724 936 1776 938
rect 1724 935 1725 936
rect 1719 934 1725 935
rect 1775 935 1776 936
rect 1780 935 1781 939
rect 1775 934 1781 935
rect 1839 939 1845 940
rect 1839 935 1840 939
rect 1844 938 1845 939
rect 1886 939 1892 940
rect 1886 938 1887 939
rect 1844 936 1887 938
rect 1844 935 1845 936
rect 1839 934 1845 935
rect 1886 935 1887 936
rect 1891 935 1892 939
rect 1886 934 1892 935
rect 1903 939 1909 940
rect 1903 935 1904 939
rect 1908 938 1909 939
rect 1966 939 1972 940
rect 1966 938 1967 939
rect 1908 936 1967 938
rect 1908 935 1909 936
rect 1903 934 1909 935
rect 1966 935 1967 936
rect 1971 935 1972 939
rect 1966 934 1972 935
rect 1975 939 1981 940
rect 1975 935 1976 939
rect 1980 938 1981 939
rect 2038 939 2044 940
rect 2038 938 2039 939
rect 1980 936 2039 938
rect 1980 935 1981 936
rect 1975 934 1981 935
rect 2038 935 2039 936
rect 2043 935 2044 939
rect 2038 934 2044 935
rect 2046 939 2053 940
rect 2046 935 2047 939
rect 2052 935 2053 939
rect 2046 934 2053 935
rect 2094 939 2101 940
rect 2094 935 2095 939
rect 2100 935 2101 939
rect 2094 934 2101 935
rect 2118 936 2124 937
rect 287 931 293 932
rect 287 927 288 931
rect 292 930 293 931
rect 318 931 324 932
rect 318 930 319 931
rect 292 928 319 930
rect 292 927 293 928
rect 287 926 293 927
rect 318 927 319 928
rect 323 927 324 931
rect 318 926 324 927
rect 327 931 333 932
rect 327 927 328 931
rect 332 930 333 931
rect 366 931 372 932
rect 366 930 367 931
rect 332 928 367 930
rect 332 927 333 928
rect 327 926 333 927
rect 366 927 367 928
rect 371 927 372 931
rect 366 926 372 927
rect 375 931 381 932
rect 375 927 376 931
rect 380 930 381 931
rect 414 931 420 932
rect 414 930 415 931
rect 380 928 415 930
rect 380 927 381 928
rect 375 926 381 927
rect 414 927 415 928
rect 419 927 420 931
rect 414 926 420 927
rect 423 931 432 932
rect 423 927 424 931
rect 431 927 432 931
rect 423 926 432 927
rect 479 931 485 932
rect 479 927 480 931
rect 484 930 485 931
rect 522 931 528 932
rect 522 930 523 931
rect 484 928 523 930
rect 484 927 485 928
rect 479 926 485 927
rect 522 927 523 928
rect 527 927 528 931
rect 522 926 528 927
rect 535 931 541 932
rect 535 927 536 931
rect 540 930 541 931
rect 574 931 580 932
rect 574 930 575 931
rect 540 928 575 930
rect 540 927 541 928
rect 535 926 541 927
rect 574 927 575 928
rect 579 927 580 931
rect 574 926 580 927
rect 591 931 597 932
rect 591 927 592 931
rect 596 930 597 931
rect 638 931 644 932
rect 638 930 639 931
rect 596 928 639 930
rect 596 927 597 928
rect 591 926 597 927
rect 638 927 639 928
rect 643 927 644 931
rect 638 926 644 927
rect 646 931 653 932
rect 646 927 647 931
rect 652 927 653 931
rect 646 926 653 927
rect 711 931 717 932
rect 711 927 712 931
rect 716 930 717 931
rect 766 931 772 932
rect 766 930 767 931
rect 716 928 767 930
rect 716 927 717 928
rect 711 926 717 927
rect 766 927 767 928
rect 771 927 772 931
rect 766 926 772 927
rect 775 931 781 932
rect 775 927 776 931
rect 780 930 781 931
rect 830 931 836 932
rect 830 930 831 931
rect 780 928 831 930
rect 780 927 781 928
rect 775 926 781 927
rect 830 927 831 928
rect 835 927 836 931
rect 830 926 836 927
rect 839 931 845 932
rect 839 927 840 931
rect 844 930 845 931
rect 894 931 900 932
rect 894 930 895 931
rect 844 928 895 930
rect 844 927 845 928
rect 839 926 845 927
rect 894 927 895 928
rect 899 927 900 931
rect 894 926 900 927
rect 903 931 909 932
rect 903 927 904 931
rect 908 930 909 931
rect 958 931 964 932
rect 958 930 959 931
rect 908 928 959 930
rect 908 927 909 928
rect 903 926 909 927
rect 958 927 959 928
rect 963 927 964 931
rect 958 926 964 927
rect 966 931 973 932
rect 966 927 967 931
rect 972 927 973 931
rect 966 926 973 927
rect 1031 931 1037 932
rect 1031 927 1032 931
rect 1036 930 1037 931
rect 1062 931 1068 932
rect 1062 930 1063 931
rect 1036 928 1063 930
rect 1036 927 1037 928
rect 1031 926 1037 927
rect 1062 927 1063 928
rect 1067 927 1068 931
rect 1062 926 1068 927
rect 1071 931 1077 932
rect 1134 931 1140 932
rect 2118 932 2119 936
rect 2123 932 2124 936
rect 2118 931 2124 932
rect 1071 927 1072 931
rect 1076 927 1077 931
rect 1071 926 1077 927
rect 1158 928 1164 929
rect 262 924 268 925
rect 262 920 263 924
rect 267 920 268 924
rect 262 919 268 920
rect 302 924 308 925
rect 302 920 303 924
rect 307 920 308 924
rect 302 919 308 920
rect 350 924 356 925
rect 350 920 351 924
rect 355 920 356 924
rect 350 919 356 920
rect 398 924 404 925
rect 398 920 399 924
rect 403 920 404 924
rect 398 919 404 920
rect 454 924 460 925
rect 454 920 455 924
rect 459 920 460 924
rect 454 919 460 920
rect 510 924 516 925
rect 510 920 511 924
rect 515 920 516 924
rect 510 919 516 920
rect 566 924 572 925
rect 566 920 567 924
rect 571 920 572 924
rect 566 919 572 920
rect 622 924 628 925
rect 622 920 623 924
rect 627 920 628 924
rect 622 919 628 920
rect 686 924 692 925
rect 686 920 687 924
rect 691 920 692 924
rect 686 919 692 920
rect 750 924 756 925
rect 750 920 751 924
rect 755 920 756 924
rect 750 919 756 920
rect 814 924 820 925
rect 814 920 815 924
rect 819 920 820 924
rect 814 919 820 920
rect 878 924 884 925
rect 878 920 879 924
rect 883 920 884 924
rect 878 919 884 920
rect 942 924 948 925
rect 942 920 943 924
rect 947 920 948 924
rect 942 919 948 920
rect 1006 924 1012 925
rect 1006 920 1007 924
rect 1011 920 1012 924
rect 1006 919 1012 920
rect 1046 924 1052 925
rect 1046 920 1047 924
rect 1051 920 1052 924
rect 1158 924 1159 928
rect 1163 924 1164 928
rect 1158 923 1164 924
rect 1206 928 1212 929
rect 1206 924 1207 928
rect 1211 924 1212 928
rect 1206 923 1212 924
rect 1286 928 1292 929
rect 1286 924 1287 928
rect 1291 924 1292 928
rect 1286 923 1292 924
rect 1374 928 1380 929
rect 1374 924 1375 928
rect 1379 924 1380 928
rect 1374 923 1380 924
rect 1454 928 1460 929
rect 1454 924 1455 928
rect 1459 924 1460 928
rect 1454 923 1460 924
rect 1534 928 1540 929
rect 1534 924 1535 928
rect 1539 924 1540 928
rect 1534 923 1540 924
rect 1614 928 1620 929
rect 1614 924 1615 928
rect 1619 924 1620 928
rect 1614 923 1620 924
rect 1686 928 1692 929
rect 1686 924 1687 928
rect 1691 924 1692 928
rect 1686 923 1692 924
rect 1750 928 1756 929
rect 1750 924 1751 928
rect 1755 924 1756 928
rect 1750 923 1756 924
rect 1814 928 1820 929
rect 1814 924 1815 928
rect 1819 924 1820 928
rect 1814 923 1820 924
rect 1878 928 1884 929
rect 1878 924 1879 928
rect 1883 924 1884 928
rect 1878 923 1884 924
rect 1950 928 1956 929
rect 1950 924 1951 928
rect 1955 924 1956 928
rect 1950 923 1956 924
rect 2022 928 2028 929
rect 2022 924 2023 928
rect 2027 924 2028 928
rect 2022 923 2028 924
rect 2070 928 2076 929
rect 2070 924 2071 928
rect 2075 924 2076 928
rect 2070 923 2076 924
rect 1046 919 1052 920
rect 1183 919 1189 920
rect 110 916 116 917
rect 110 912 111 916
rect 115 912 116 916
rect 1094 916 1100 917
rect 1094 912 1095 916
rect 1099 912 1100 916
rect 1183 915 1184 919
rect 1188 918 1189 919
rect 1214 919 1220 920
rect 1214 918 1215 919
rect 1188 916 1215 918
rect 1188 915 1189 916
rect 1183 914 1189 915
rect 1214 915 1215 916
rect 1219 915 1220 919
rect 1214 914 1220 915
rect 1222 919 1228 920
rect 1222 915 1223 919
rect 1227 918 1228 919
rect 1231 919 1237 920
rect 1231 918 1232 919
rect 1227 916 1232 918
rect 1227 915 1228 916
rect 1222 914 1228 915
rect 1231 915 1232 916
rect 1236 915 1237 919
rect 1231 914 1237 915
rect 1266 919 1272 920
rect 1266 915 1267 919
rect 1271 918 1272 919
rect 1311 919 1317 920
rect 1311 918 1312 919
rect 1271 916 1312 918
rect 1271 915 1272 916
rect 1266 914 1272 915
rect 1311 915 1312 916
rect 1316 915 1317 919
rect 1311 914 1317 915
rect 1390 919 1396 920
rect 1390 915 1391 919
rect 1395 918 1396 919
rect 1399 919 1405 920
rect 1399 918 1400 919
rect 1395 916 1400 918
rect 1395 915 1396 916
rect 1390 914 1396 915
rect 1399 915 1400 916
rect 1404 915 1405 919
rect 1399 914 1405 915
rect 1479 919 1488 920
rect 1479 915 1480 919
rect 1487 915 1488 919
rect 1479 914 1488 915
rect 1550 919 1556 920
rect 1550 915 1551 919
rect 1555 918 1556 919
rect 1559 919 1565 920
rect 1559 918 1560 919
rect 1555 916 1560 918
rect 1555 915 1556 916
rect 1550 914 1556 915
rect 1559 915 1560 916
rect 1564 915 1565 919
rect 1559 914 1565 915
rect 1639 919 1645 920
rect 1639 915 1640 919
rect 1644 918 1645 919
rect 1647 919 1653 920
rect 1647 918 1648 919
rect 1644 916 1648 918
rect 1644 915 1645 916
rect 1639 914 1645 915
rect 1647 915 1648 916
rect 1652 915 1653 919
rect 1647 914 1653 915
rect 1711 919 1717 920
rect 1711 915 1712 919
rect 1716 918 1717 919
rect 1719 919 1725 920
rect 1719 918 1720 919
rect 1716 916 1720 918
rect 1716 915 1717 916
rect 1711 914 1717 915
rect 1719 915 1720 916
rect 1724 915 1725 919
rect 1719 914 1725 915
rect 1775 919 1784 920
rect 1775 915 1776 919
rect 1783 915 1784 919
rect 1775 914 1784 915
rect 1838 919 1845 920
rect 1838 915 1839 919
rect 1844 915 1845 919
rect 1838 914 1845 915
rect 1886 919 1892 920
rect 1886 915 1887 919
rect 1891 918 1892 919
rect 1903 919 1909 920
rect 1903 918 1904 919
rect 1891 916 1904 918
rect 1891 915 1892 916
rect 1886 914 1892 915
rect 1903 915 1904 916
rect 1908 915 1909 919
rect 1903 914 1909 915
rect 1966 919 1972 920
rect 1966 915 1967 919
rect 1971 918 1972 919
rect 1975 919 1981 920
rect 1975 918 1976 919
rect 1971 916 1976 918
rect 1971 915 1972 916
rect 1966 914 1972 915
rect 1975 915 1976 916
rect 1980 915 1981 919
rect 1975 914 1981 915
rect 2038 919 2044 920
rect 2038 915 2039 919
rect 2043 918 2044 919
rect 2047 919 2053 920
rect 2047 918 2048 919
rect 2043 916 2048 918
rect 2043 915 2044 916
rect 2038 914 2044 915
rect 2047 915 2048 916
rect 2052 915 2053 919
rect 2047 914 2053 915
rect 2055 919 2061 920
rect 2055 915 2056 919
rect 2060 918 2061 919
rect 2095 919 2101 920
rect 2095 918 2096 919
rect 2060 916 2096 918
rect 2060 915 2061 916
rect 2055 914 2061 915
rect 2095 915 2096 916
rect 2100 915 2101 919
rect 2095 914 2101 915
rect 110 911 116 912
rect 287 911 296 912
rect 287 907 288 911
rect 295 907 296 911
rect 287 906 296 907
rect 318 911 324 912
rect 318 907 319 911
rect 323 910 324 911
rect 327 911 333 912
rect 327 910 328 911
rect 323 908 328 910
rect 323 907 324 908
rect 318 906 324 907
rect 327 907 328 908
rect 332 907 333 911
rect 327 906 333 907
rect 366 911 372 912
rect 366 907 367 911
rect 371 910 372 911
rect 375 911 381 912
rect 375 910 376 911
rect 371 908 376 910
rect 371 907 372 908
rect 366 906 372 907
rect 375 907 376 908
rect 380 907 381 911
rect 375 906 381 907
rect 414 911 420 912
rect 414 907 415 911
rect 419 910 420 911
rect 423 911 429 912
rect 423 910 424 911
rect 419 908 424 910
rect 419 907 420 908
rect 414 906 420 907
rect 423 907 424 908
rect 428 907 429 911
rect 423 906 429 907
rect 479 911 488 912
rect 479 907 480 911
rect 487 907 488 911
rect 479 906 488 907
rect 522 911 528 912
rect 522 907 523 911
rect 527 910 528 911
rect 535 911 541 912
rect 535 910 536 911
rect 527 908 536 910
rect 527 907 528 908
rect 522 906 528 907
rect 535 907 536 908
rect 540 907 541 911
rect 535 906 541 907
rect 574 911 580 912
rect 574 907 575 911
rect 579 910 580 911
rect 591 911 597 912
rect 591 910 592 911
rect 579 908 592 910
rect 579 907 580 908
rect 574 906 580 907
rect 591 907 592 908
rect 596 907 597 911
rect 591 906 597 907
rect 638 911 644 912
rect 638 907 639 911
rect 643 910 644 911
rect 647 911 653 912
rect 647 910 648 911
rect 643 908 648 910
rect 643 907 644 908
rect 638 906 644 907
rect 647 907 648 908
rect 652 907 653 911
rect 647 906 653 907
rect 711 911 720 912
rect 711 907 712 911
rect 719 907 720 911
rect 711 906 720 907
rect 766 911 772 912
rect 766 907 767 911
rect 771 910 772 911
rect 775 911 781 912
rect 775 910 776 911
rect 771 908 776 910
rect 771 907 772 908
rect 766 906 772 907
rect 775 907 776 908
rect 780 907 781 911
rect 775 906 781 907
rect 830 911 836 912
rect 830 907 831 911
rect 835 910 836 911
rect 839 911 845 912
rect 839 910 840 911
rect 835 908 840 910
rect 835 907 836 908
rect 830 906 836 907
rect 839 907 840 908
rect 844 907 845 911
rect 839 906 845 907
rect 894 911 900 912
rect 894 907 895 911
rect 899 910 900 911
rect 903 911 909 912
rect 903 910 904 911
rect 899 908 904 910
rect 899 907 900 908
rect 894 906 900 907
rect 903 907 904 908
rect 908 907 909 911
rect 903 906 909 907
rect 958 911 964 912
rect 958 907 959 911
rect 963 910 964 911
rect 967 911 973 912
rect 967 910 968 911
rect 963 908 968 910
rect 963 907 964 908
rect 958 906 964 907
rect 967 907 968 908
rect 972 907 973 911
rect 967 906 973 907
rect 1031 911 1037 912
rect 1031 907 1032 911
rect 1036 910 1037 911
rect 1054 911 1060 912
rect 1054 910 1055 911
rect 1036 908 1055 910
rect 1036 907 1037 908
rect 1031 906 1037 907
rect 1054 907 1055 908
rect 1059 907 1060 911
rect 1054 906 1060 907
rect 1062 911 1068 912
rect 1062 907 1063 911
rect 1067 910 1068 911
rect 1071 911 1077 912
rect 1094 911 1100 912
rect 1071 910 1072 911
rect 1067 908 1072 910
rect 1067 907 1068 908
rect 1062 906 1068 907
rect 1071 907 1072 908
rect 1076 907 1077 911
rect 1071 906 1077 907
rect 110 899 116 900
rect 110 895 111 899
rect 115 895 116 899
rect 1094 899 1100 900
rect 110 894 116 895
rect 262 896 268 897
rect 262 892 263 896
rect 267 892 268 896
rect 262 891 268 892
rect 302 896 308 897
rect 302 892 303 896
rect 307 892 308 896
rect 302 891 308 892
rect 350 896 356 897
rect 350 892 351 896
rect 355 892 356 896
rect 350 891 356 892
rect 398 896 404 897
rect 398 892 399 896
rect 403 892 404 896
rect 398 891 404 892
rect 454 896 460 897
rect 454 892 455 896
rect 459 892 460 896
rect 454 891 460 892
rect 510 896 516 897
rect 510 892 511 896
rect 515 892 516 896
rect 510 891 516 892
rect 566 896 572 897
rect 566 892 567 896
rect 571 892 572 896
rect 566 891 572 892
rect 622 896 628 897
rect 622 892 623 896
rect 627 892 628 896
rect 622 891 628 892
rect 686 896 692 897
rect 686 892 687 896
rect 691 892 692 896
rect 686 891 692 892
rect 750 896 756 897
rect 750 892 751 896
rect 755 892 756 896
rect 750 891 756 892
rect 814 896 820 897
rect 814 892 815 896
rect 819 892 820 896
rect 814 891 820 892
rect 878 896 884 897
rect 878 892 879 896
rect 883 892 884 896
rect 878 891 884 892
rect 942 896 948 897
rect 942 892 943 896
rect 947 892 948 896
rect 942 891 948 892
rect 1006 896 1012 897
rect 1006 892 1007 896
rect 1011 892 1012 896
rect 1006 891 1012 892
rect 1046 896 1052 897
rect 1046 892 1047 896
rect 1051 892 1052 896
rect 1094 895 1095 899
rect 1099 895 1100 899
rect 1094 894 1100 895
rect 1263 899 1269 900
rect 1263 895 1264 899
rect 1268 898 1269 899
rect 1334 899 1340 900
rect 1334 898 1335 899
rect 1268 896 1335 898
rect 1268 895 1269 896
rect 1263 894 1269 895
rect 1334 895 1335 896
rect 1339 895 1340 899
rect 1334 894 1340 895
rect 1343 899 1349 900
rect 1343 895 1344 899
rect 1348 898 1349 899
rect 1378 899 1384 900
rect 1378 898 1379 899
rect 1348 896 1379 898
rect 1348 895 1349 896
rect 1343 894 1349 895
rect 1378 895 1379 896
rect 1383 895 1384 899
rect 1378 894 1384 895
rect 1386 899 1392 900
rect 1386 895 1387 899
rect 1391 898 1392 899
rect 1431 899 1437 900
rect 1431 898 1432 899
rect 1391 896 1432 898
rect 1391 895 1392 896
rect 1386 894 1392 895
rect 1431 895 1432 896
rect 1436 895 1437 899
rect 1431 894 1437 895
rect 1519 899 1525 900
rect 1519 895 1520 899
rect 1524 898 1525 899
rect 1598 899 1604 900
rect 1598 898 1599 899
rect 1524 896 1599 898
rect 1524 895 1525 896
rect 1519 894 1525 895
rect 1598 895 1599 896
rect 1603 895 1604 899
rect 1598 894 1604 895
rect 1606 899 1613 900
rect 1606 895 1607 899
rect 1612 895 1613 899
rect 1606 894 1613 895
rect 1687 899 1693 900
rect 1687 895 1688 899
rect 1692 898 1693 899
rect 1758 899 1764 900
rect 1758 898 1759 899
rect 1692 896 1759 898
rect 1692 895 1693 896
rect 1687 894 1693 895
rect 1758 895 1759 896
rect 1763 895 1764 899
rect 1758 894 1764 895
rect 1767 899 1773 900
rect 1767 895 1768 899
rect 1772 898 1773 899
rect 1806 899 1812 900
rect 1806 898 1807 899
rect 1772 896 1807 898
rect 1772 895 1773 896
rect 1767 894 1773 895
rect 1806 895 1807 896
rect 1811 895 1812 899
rect 1806 894 1812 895
rect 1839 899 1845 900
rect 1839 895 1840 899
rect 1844 898 1845 899
rect 1902 899 1908 900
rect 1902 898 1903 899
rect 1844 896 1903 898
rect 1844 895 1845 896
rect 1839 894 1845 895
rect 1902 895 1903 896
rect 1907 895 1908 899
rect 1902 894 1908 895
rect 1911 899 1917 900
rect 1911 895 1912 899
rect 1916 898 1917 899
rect 1966 899 1972 900
rect 1966 898 1967 899
rect 1916 896 1967 898
rect 1916 895 1917 896
rect 1911 894 1917 895
rect 1966 895 1967 896
rect 1971 895 1972 899
rect 1966 894 1972 895
rect 1975 899 1981 900
rect 1975 895 1976 899
rect 1980 898 1981 899
rect 2038 899 2044 900
rect 2038 898 2039 899
rect 1980 896 2039 898
rect 1980 895 1981 896
rect 1975 894 1981 895
rect 2038 895 2039 896
rect 2043 895 2044 899
rect 2038 894 2044 895
rect 2046 899 2053 900
rect 2046 895 2047 899
rect 2052 895 2053 899
rect 2046 894 2053 895
rect 2094 899 2101 900
rect 2094 895 2095 899
rect 2100 895 2101 899
rect 2094 894 2101 895
rect 1046 891 1052 892
rect 1238 892 1244 893
rect 1238 888 1239 892
rect 1243 888 1244 892
rect 1238 887 1244 888
rect 1318 892 1324 893
rect 1318 888 1319 892
rect 1323 888 1324 892
rect 1318 887 1324 888
rect 1406 892 1412 893
rect 1406 888 1407 892
rect 1411 888 1412 892
rect 1406 887 1412 888
rect 1494 892 1500 893
rect 1494 888 1495 892
rect 1499 888 1500 892
rect 1494 887 1500 888
rect 1582 892 1588 893
rect 1582 888 1583 892
rect 1587 888 1588 892
rect 1582 887 1588 888
rect 1662 892 1668 893
rect 1662 888 1663 892
rect 1667 888 1668 892
rect 1662 887 1668 888
rect 1742 892 1748 893
rect 1742 888 1743 892
rect 1747 888 1748 892
rect 1742 887 1748 888
rect 1814 892 1820 893
rect 1814 888 1815 892
rect 1819 888 1820 892
rect 1814 887 1820 888
rect 1886 892 1892 893
rect 1886 888 1887 892
rect 1891 888 1892 892
rect 1886 887 1892 888
rect 1950 892 1956 893
rect 1950 888 1951 892
rect 1955 888 1956 892
rect 1950 887 1956 888
rect 2022 892 2028 893
rect 2022 888 2023 892
rect 2027 888 2028 892
rect 2022 887 2028 888
rect 2070 892 2076 893
rect 2070 888 2071 892
rect 2075 888 2076 892
rect 2070 887 2076 888
rect 1134 884 1140 885
rect 302 880 308 881
rect 110 877 116 878
rect 110 873 111 877
rect 115 873 116 877
rect 302 876 303 880
rect 307 876 308 880
rect 302 875 308 876
rect 350 880 356 881
rect 350 876 351 880
rect 355 876 356 880
rect 350 875 356 876
rect 414 880 420 881
rect 414 876 415 880
rect 419 876 420 880
rect 414 875 420 876
rect 478 880 484 881
rect 478 876 479 880
rect 483 876 484 880
rect 478 875 484 876
rect 550 880 556 881
rect 550 876 551 880
rect 555 876 556 880
rect 550 875 556 876
rect 622 880 628 881
rect 622 876 623 880
rect 627 876 628 880
rect 622 875 628 876
rect 694 880 700 881
rect 694 876 695 880
rect 699 876 700 880
rect 694 875 700 876
rect 766 880 772 881
rect 766 876 767 880
rect 771 876 772 880
rect 766 875 772 876
rect 830 880 836 881
rect 830 876 831 880
rect 835 876 836 880
rect 830 875 836 876
rect 886 880 892 881
rect 886 876 887 880
rect 891 876 892 880
rect 886 875 892 876
rect 942 880 948 881
rect 942 876 943 880
rect 947 876 948 880
rect 942 875 948 876
rect 1006 880 1012 881
rect 1006 876 1007 880
rect 1011 876 1012 880
rect 1006 875 1012 876
rect 1046 880 1052 881
rect 1046 876 1047 880
rect 1051 876 1052 880
rect 1134 880 1135 884
rect 1139 880 1140 884
rect 2118 884 2124 885
rect 2118 880 2119 884
rect 2123 880 2124 884
rect 1134 879 1140 880
rect 1263 879 1272 880
rect 1046 875 1052 876
rect 1094 877 1100 878
rect 110 872 116 873
rect 1094 873 1095 877
rect 1099 873 1100 877
rect 1263 875 1264 879
rect 1271 875 1272 879
rect 1263 874 1272 875
rect 1334 879 1340 880
rect 1334 875 1335 879
rect 1339 878 1340 879
rect 1343 879 1349 880
rect 1343 878 1344 879
rect 1339 876 1344 878
rect 1339 875 1340 876
rect 1334 874 1340 875
rect 1343 875 1344 876
rect 1348 875 1349 879
rect 1343 874 1349 875
rect 1378 879 1384 880
rect 1378 875 1379 879
rect 1383 878 1384 879
rect 1431 879 1437 880
rect 1431 878 1432 879
rect 1383 876 1432 878
rect 1383 875 1384 876
rect 1378 874 1384 875
rect 1431 875 1432 876
rect 1436 875 1437 879
rect 1431 874 1437 875
rect 1482 879 1488 880
rect 1482 875 1483 879
rect 1487 878 1488 879
rect 1519 879 1525 880
rect 1519 878 1520 879
rect 1487 876 1520 878
rect 1487 875 1488 876
rect 1482 874 1488 875
rect 1519 875 1520 876
rect 1524 875 1525 879
rect 1519 874 1525 875
rect 1598 879 1604 880
rect 1598 875 1599 879
rect 1603 878 1604 879
rect 1607 879 1613 880
rect 1607 878 1608 879
rect 1603 876 1608 878
rect 1603 875 1604 876
rect 1598 874 1604 875
rect 1607 875 1608 876
rect 1612 875 1613 879
rect 1607 874 1613 875
rect 1687 879 1693 880
rect 1687 875 1688 879
rect 1692 878 1693 879
rect 1734 879 1740 880
rect 1734 878 1735 879
rect 1692 876 1735 878
rect 1692 875 1693 876
rect 1687 874 1693 875
rect 1734 875 1735 876
rect 1739 875 1740 879
rect 1734 874 1740 875
rect 1758 879 1764 880
rect 1758 875 1759 879
rect 1763 878 1764 879
rect 1767 879 1773 880
rect 1767 878 1768 879
rect 1763 876 1768 878
rect 1763 875 1764 876
rect 1758 874 1764 875
rect 1767 875 1768 876
rect 1772 875 1773 879
rect 1767 874 1773 875
rect 1839 879 1845 880
rect 1839 875 1840 879
rect 1844 878 1845 879
rect 1894 879 1900 880
rect 1894 878 1895 879
rect 1844 876 1895 878
rect 1844 875 1845 876
rect 1839 874 1845 875
rect 1894 875 1895 876
rect 1899 875 1900 879
rect 1894 874 1900 875
rect 1902 879 1908 880
rect 1902 875 1903 879
rect 1907 878 1908 879
rect 1911 879 1917 880
rect 1911 878 1912 879
rect 1907 876 1912 878
rect 1907 875 1908 876
rect 1902 874 1908 875
rect 1911 875 1912 876
rect 1916 875 1917 879
rect 1911 874 1917 875
rect 1966 879 1972 880
rect 1966 875 1967 879
rect 1971 878 1972 879
rect 1975 879 1981 880
rect 1975 878 1976 879
rect 1971 876 1976 878
rect 1971 875 1972 876
rect 1966 874 1972 875
rect 1975 875 1976 876
rect 1980 875 1981 879
rect 1975 874 1981 875
rect 2038 879 2044 880
rect 2038 875 2039 879
rect 2043 878 2044 879
rect 2047 879 2053 880
rect 2047 878 2048 879
rect 2043 876 2048 878
rect 2043 875 2044 876
rect 2038 874 2044 875
rect 2047 875 2048 876
rect 2052 875 2053 879
rect 2047 874 2053 875
rect 2094 879 2101 880
rect 2118 879 2124 880
rect 2094 875 2095 879
rect 2100 875 2101 879
rect 2094 874 2101 875
rect 1094 872 1100 873
rect 966 871 972 872
rect 966 870 967 871
rect 724 868 967 870
rect 724 864 726 868
rect 966 867 967 868
rect 971 867 972 871
rect 966 866 972 867
rect 1134 867 1140 868
rect 310 863 316 864
rect 110 860 116 861
rect 110 856 111 860
rect 115 856 116 860
rect 310 859 311 863
rect 315 862 316 863
rect 327 863 333 864
rect 327 862 328 863
rect 315 860 328 862
rect 315 859 316 860
rect 310 858 316 859
rect 327 859 328 860
rect 332 859 333 863
rect 327 858 333 859
rect 335 863 341 864
rect 335 859 336 863
rect 340 862 341 863
rect 375 863 381 864
rect 375 862 376 863
rect 340 860 376 862
rect 340 859 341 860
rect 335 858 341 859
rect 375 859 376 860
rect 380 859 381 863
rect 439 863 445 864
rect 439 862 440 863
rect 375 858 381 859
rect 409 860 440 862
rect 110 855 116 856
rect 302 852 308 853
rect 302 848 303 852
rect 307 848 308 852
rect 302 847 308 848
rect 350 852 356 853
rect 350 848 351 852
rect 355 848 356 852
rect 350 847 356 848
rect 409 846 411 860
rect 439 859 440 860
rect 444 859 445 863
rect 439 858 445 859
rect 503 863 509 864
rect 503 859 504 863
rect 508 862 509 863
rect 566 863 572 864
rect 566 862 567 863
rect 508 860 567 862
rect 508 859 509 860
rect 503 858 509 859
rect 566 859 567 860
rect 571 859 572 863
rect 566 858 572 859
rect 575 863 581 864
rect 575 859 576 863
rect 580 862 581 863
rect 638 863 644 864
rect 638 862 639 863
rect 580 860 639 862
rect 580 859 581 860
rect 575 858 581 859
rect 638 859 639 860
rect 643 859 644 863
rect 638 858 644 859
rect 646 863 653 864
rect 646 859 647 863
rect 652 859 653 863
rect 646 858 653 859
rect 719 863 726 864
rect 719 859 720 863
rect 724 860 726 863
rect 730 863 736 864
rect 724 859 725 860
rect 719 858 725 859
rect 730 859 731 863
rect 735 862 736 863
rect 791 863 797 864
rect 791 862 792 863
rect 735 860 792 862
rect 735 859 736 860
rect 730 858 736 859
rect 791 859 792 860
rect 796 859 797 863
rect 791 858 797 859
rect 799 863 805 864
rect 799 859 800 863
rect 804 862 805 863
rect 855 863 861 864
rect 855 862 856 863
rect 804 860 856 862
rect 804 859 805 860
rect 799 858 805 859
rect 855 859 856 860
rect 860 859 861 863
rect 855 858 861 859
rect 863 863 869 864
rect 863 859 864 863
rect 868 862 869 863
rect 911 863 917 864
rect 911 862 912 863
rect 868 860 912 862
rect 868 859 869 860
rect 863 858 869 859
rect 911 859 912 860
rect 916 859 917 863
rect 911 858 917 859
rect 934 863 940 864
rect 934 859 935 863
rect 939 862 940 863
rect 967 863 973 864
rect 967 862 968 863
rect 939 860 968 862
rect 939 859 940 860
rect 934 858 940 859
rect 967 859 968 860
rect 972 859 973 863
rect 967 858 973 859
rect 975 863 981 864
rect 975 859 976 863
rect 980 862 981 863
rect 1031 863 1037 864
rect 1031 862 1032 863
rect 980 860 1032 862
rect 980 859 981 860
rect 975 858 981 859
rect 1031 859 1032 860
rect 1036 859 1037 863
rect 1031 858 1037 859
rect 1054 863 1060 864
rect 1054 859 1055 863
rect 1059 862 1060 863
rect 1071 863 1077 864
rect 1071 862 1072 863
rect 1059 860 1072 862
rect 1059 859 1060 860
rect 1054 858 1060 859
rect 1071 859 1072 860
rect 1076 859 1077 863
rect 1134 863 1135 867
rect 1139 863 1140 867
rect 2118 867 2124 868
rect 1134 862 1140 863
rect 1238 864 1244 865
rect 1071 858 1077 859
rect 1094 860 1100 861
rect 1094 856 1095 860
rect 1099 856 1100 860
rect 1238 860 1239 864
rect 1243 860 1244 864
rect 1238 859 1244 860
rect 1318 864 1324 865
rect 1318 860 1319 864
rect 1323 860 1324 864
rect 1318 859 1324 860
rect 1406 864 1412 865
rect 1406 860 1407 864
rect 1411 860 1412 864
rect 1406 859 1412 860
rect 1494 864 1500 865
rect 1494 860 1495 864
rect 1499 860 1500 864
rect 1494 859 1500 860
rect 1582 864 1588 865
rect 1582 860 1583 864
rect 1587 860 1588 864
rect 1582 859 1588 860
rect 1662 864 1668 865
rect 1662 860 1663 864
rect 1667 860 1668 864
rect 1662 859 1668 860
rect 1742 864 1748 865
rect 1742 860 1743 864
rect 1747 860 1748 864
rect 1742 859 1748 860
rect 1814 864 1820 865
rect 1814 860 1815 864
rect 1819 860 1820 864
rect 1814 859 1820 860
rect 1886 864 1892 865
rect 1886 860 1887 864
rect 1891 860 1892 864
rect 1886 859 1892 860
rect 1950 864 1956 865
rect 1950 860 1951 864
rect 1955 860 1956 864
rect 1950 859 1956 860
rect 2022 864 2028 865
rect 2022 860 2023 864
rect 2027 860 2028 864
rect 2022 859 2028 860
rect 2070 864 2076 865
rect 2070 860 2071 864
rect 2075 860 2076 864
rect 2118 863 2119 867
rect 2123 863 2124 867
rect 2118 862 2124 863
rect 2070 859 2076 860
rect 1094 855 1100 856
rect 414 852 420 853
rect 414 848 415 852
rect 419 848 420 852
rect 414 847 420 848
rect 478 852 484 853
rect 478 848 479 852
rect 483 848 484 852
rect 478 847 484 848
rect 550 852 556 853
rect 550 848 551 852
rect 555 848 556 852
rect 550 847 556 848
rect 622 852 628 853
rect 622 848 623 852
rect 627 848 628 852
rect 622 847 628 848
rect 694 852 700 853
rect 694 848 695 852
rect 699 848 700 852
rect 694 847 700 848
rect 766 852 772 853
rect 766 848 767 852
rect 771 848 772 852
rect 766 847 772 848
rect 830 852 836 853
rect 830 848 831 852
rect 835 848 836 852
rect 830 847 836 848
rect 886 852 892 853
rect 886 848 887 852
rect 891 848 892 852
rect 886 847 892 848
rect 942 852 948 853
rect 942 848 943 852
rect 947 848 948 852
rect 942 847 948 848
rect 1006 852 1012 853
rect 1006 848 1007 852
rect 1011 848 1012 852
rect 1006 847 1012 848
rect 1046 852 1052 853
rect 1046 848 1047 852
rect 1051 848 1052 852
rect 1158 852 1164 853
rect 1046 847 1052 848
rect 1134 849 1140 850
rect 377 844 411 846
rect 1134 845 1135 849
rect 1139 845 1140 849
rect 1158 848 1159 852
rect 1163 848 1164 852
rect 1158 847 1164 848
rect 1246 852 1252 853
rect 1246 848 1247 852
rect 1251 848 1252 852
rect 1246 847 1252 848
rect 1358 852 1364 853
rect 1358 848 1359 852
rect 1363 848 1364 852
rect 1358 847 1364 848
rect 1454 852 1460 853
rect 1454 848 1455 852
rect 1459 848 1460 852
rect 1454 847 1460 848
rect 1542 852 1548 853
rect 1542 848 1543 852
rect 1547 848 1548 852
rect 1542 847 1548 848
rect 1630 852 1636 853
rect 1630 848 1631 852
rect 1635 848 1636 852
rect 1630 847 1636 848
rect 1710 852 1716 853
rect 1710 848 1711 852
rect 1715 848 1716 852
rect 1710 847 1716 848
rect 1782 852 1788 853
rect 1782 848 1783 852
rect 1787 848 1788 852
rect 1782 847 1788 848
rect 1854 852 1860 853
rect 1854 848 1855 852
rect 1859 848 1860 852
rect 1854 847 1860 848
rect 1934 852 1940 853
rect 1934 848 1935 852
rect 1939 848 1940 852
rect 1934 847 1940 848
rect 2014 852 2020 853
rect 2014 848 2015 852
rect 2019 848 2020 852
rect 2014 847 2020 848
rect 2070 852 2076 853
rect 2070 848 2071 852
rect 2075 848 2076 852
rect 2070 847 2076 848
rect 2118 849 2124 850
rect 1134 844 1140 845
rect 2118 845 2119 849
rect 2123 845 2124 849
rect 2118 844 2124 845
rect 327 843 333 844
rect 327 839 328 843
rect 332 842 333 843
rect 335 843 341 844
rect 335 842 336 843
rect 332 840 336 842
rect 332 839 333 840
rect 327 838 333 839
rect 335 839 336 840
rect 340 839 341 843
rect 335 838 341 839
rect 375 843 381 844
rect 375 839 376 843
rect 380 839 381 843
rect 439 843 445 844
rect 439 842 440 843
rect 375 838 381 839
rect 384 840 440 842
rect 290 835 296 836
rect 290 831 291 835
rect 295 834 296 835
rect 384 834 386 840
rect 439 839 440 840
rect 444 839 445 843
rect 439 838 445 839
rect 503 843 512 844
rect 503 839 504 843
rect 511 839 512 843
rect 503 838 512 839
rect 566 843 572 844
rect 566 839 567 843
rect 571 842 572 843
rect 575 843 581 844
rect 575 842 576 843
rect 571 840 576 842
rect 571 839 572 840
rect 566 838 572 839
rect 575 839 576 840
rect 580 839 581 843
rect 575 838 581 839
rect 638 843 644 844
rect 638 839 639 843
rect 643 842 644 843
rect 647 843 653 844
rect 647 842 648 843
rect 643 840 648 842
rect 643 839 644 840
rect 638 838 644 839
rect 647 839 648 840
rect 652 839 653 843
rect 647 838 653 839
rect 719 843 725 844
rect 719 839 720 843
rect 724 842 725 843
rect 730 843 736 844
rect 730 842 731 843
rect 724 840 731 842
rect 724 839 725 840
rect 719 838 725 839
rect 730 839 731 840
rect 735 839 736 843
rect 730 838 736 839
rect 791 843 797 844
rect 791 839 792 843
rect 796 842 797 843
rect 799 843 805 844
rect 799 842 800 843
rect 796 840 800 842
rect 796 839 797 840
rect 791 838 797 839
rect 799 839 800 840
rect 804 839 805 843
rect 799 838 805 839
rect 855 843 861 844
rect 855 839 856 843
rect 860 842 861 843
rect 863 843 869 844
rect 863 842 864 843
rect 860 840 864 842
rect 860 839 861 840
rect 855 838 861 839
rect 863 839 864 840
rect 868 839 869 843
rect 911 843 917 844
rect 911 842 912 843
rect 863 838 869 839
rect 872 840 912 842
rect 295 832 386 834
rect 754 835 760 836
rect 295 831 296 832
rect 290 830 296 831
rect 754 831 755 835
rect 759 834 760 835
rect 872 834 874 840
rect 911 839 912 840
rect 916 839 917 843
rect 911 838 917 839
rect 967 843 973 844
rect 967 839 968 843
rect 972 842 973 843
rect 975 843 981 844
rect 975 842 976 843
rect 972 840 976 842
rect 972 839 973 840
rect 967 838 973 839
rect 975 839 976 840
rect 980 839 981 843
rect 975 838 981 839
rect 1031 843 1037 844
rect 1031 839 1032 843
rect 1036 842 1037 843
rect 1054 843 1060 844
rect 1054 842 1055 843
rect 1036 840 1055 842
rect 1036 839 1037 840
rect 1031 838 1037 839
rect 1054 839 1055 840
rect 1059 839 1060 843
rect 1054 838 1060 839
rect 1062 843 1068 844
rect 1062 839 1063 843
rect 1067 842 1068 843
rect 1071 843 1077 844
rect 1071 842 1072 843
rect 1067 840 1072 842
rect 1067 839 1068 840
rect 1062 838 1068 839
rect 1071 839 1072 840
rect 1076 839 1077 843
rect 1071 838 1077 839
rect 759 832 874 834
rect 1183 835 1189 836
rect 1134 832 1140 833
rect 759 831 760 832
rect 754 830 760 831
rect 934 831 940 832
rect 934 830 935 831
rect 880 828 935 830
rect 303 823 309 824
rect 303 819 304 823
rect 308 819 309 823
rect 303 818 309 819
rect 334 823 340 824
rect 334 819 335 823
rect 339 822 340 823
rect 367 823 373 824
rect 367 822 368 823
rect 339 820 368 822
rect 339 819 340 820
rect 334 818 340 819
rect 367 819 368 820
rect 372 819 373 823
rect 367 818 373 819
rect 375 823 381 824
rect 375 819 376 823
rect 380 822 381 823
rect 439 823 445 824
rect 439 822 440 823
rect 380 820 440 822
rect 380 819 381 820
rect 375 818 381 819
rect 439 819 440 820
rect 444 819 445 823
rect 439 818 445 819
rect 511 823 517 824
rect 511 819 512 823
rect 516 822 517 823
rect 582 823 588 824
rect 582 822 583 823
rect 516 820 583 822
rect 516 819 517 820
rect 511 818 517 819
rect 582 819 583 820
rect 587 819 588 823
rect 582 818 588 819
rect 591 823 597 824
rect 591 819 592 823
rect 596 822 597 823
rect 662 823 668 824
rect 662 822 663 823
rect 596 820 663 822
rect 596 819 597 820
rect 591 818 597 819
rect 662 819 663 820
rect 667 819 668 823
rect 662 818 668 819
rect 670 823 677 824
rect 670 819 671 823
rect 676 819 677 823
rect 670 818 677 819
rect 751 823 757 824
rect 751 819 752 823
rect 756 822 757 823
rect 814 823 820 824
rect 814 822 815 823
rect 756 820 815 822
rect 756 819 757 820
rect 751 818 757 819
rect 814 819 815 820
rect 819 819 820 823
rect 814 818 820 819
rect 823 823 829 824
rect 823 819 824 823
rect 828 822 829 823
rect 880 822 882 828
rect 934 827 935 828
rect 939 827 940 831
rect 1134 828 1135 832
rect 1139 828 1140 832
rect 1183 831 1184 835
rect 1188 834 1189 835
rect 1262 835 1268 836
rect 1262 834 1263 835
rect 1188 832 1263 834
rect 1188 831 1189 832
rect 1183 830 1189 831
rect 1262 831 1263 832
rect 1267 831 1268 835
rect 1262 830 1268 831
rect 1271 835 1277 836
rect 1271 831 1272 835
rect 1276 834 1277 835
rect 1374 835 1380 836
rect 1374 834 1375 835
rect 1276 832 1375 834
rect 1276 831 1277 832
rect 1271 830 1277 831
rect 1374 831 1375 832
rect 1379 831 1380 835
rect 1374 830 1380 831
rect 1383 835 1392 836
rect 1383 831 1384 835
rect 1391 831 1392 835
rect 1383 830 1392 831
rect 1462 835 1468 836
rect 1462 831 1463 835
rect 1467 834 1468 835
rect 1479 835 1485 836
rect 1479 834 1480 835
rect 1467 832 1480 834
rect 1467 831 1468 832
rect 1462 830 1468 831
rect 1479 831 1480 832
rect 1484 831 1485 835
rect 1479 830 1485 831
rect 1558 835 1564 836
rect 1558 831 1559 835
rect 1563 834 1564 835
rect 1567 835 1573 836
rect 1567 834 1568 835
rect 1563 832 1568 834
rect 1563 831 1564 832
rect 1558 830 1564 831
rect 1567 831 1568 832
rect 1572 831 1573 835
rect 1567 830 1573 831
rect 1575 835 1581 836
rect 1575 831 1576 835
rect 1580 834 1581 835
rect 1655 835 1661 836
rect 1655 834 1656 835
rect 1580 832 1656 834
rect 1580 831 1581 832
rect 1575 830 1581 831
rect 1655 831 1656 832
rect 1660 831 1661 835
rect 1655 830 1661 831
rect 1663 835 1669 836
rect 1663 831 1664 835
rect 1668 834 1669 835
rect 1735 835 1741 836
rect 1735 834 1736 835
rect 1668 832 1736 834
rect 1668 831 1669 832
rect 1663 830 1669 831
rect 1735 831 1736 832
rect 1740 831 1741 835
rect 1735 830 1741 831
rect 1806 835 1813 836
rect 1806 831 1807 835
rect 1812 831 1813 835
rect 1806 830 1813 831
rect 1818 835 1824 836
rect 1818 831 1819 835
rect 1823 834 1824 835
rect 1879 835 1885 836
rect 1879 834 1880 835
rect 1823 832 1880 834
rect 1823 831 1824 832
rect 1818 830 1824 831
rect 1879 831 1880 832
rect 1884 831 1885 835
rect 1879 830 1885 831
rect 1887 835 1893 836
rect 1887 831 1888 835
rect 1892 834 1893 835
rect 1959 835 1965 836
rect 1959 834 1960 835
rect 1892 832 1960 834
rect 1892 831 1893 832
rect 1887 830 1893 831
rect 1959 831 1960 832
rect 1964 831 1965 835
rect 1959 830 1965 831
rect 2039 835 2045 836
rect 2039 831 2040 835
rect 2044 834 2045 835
rect 2055 835 2061 836
rect 2055 834 2056 835
rect 2044 832 2056 834
rect 2044 831 2045 832
rect 2039 830 2045 831
rect 2055 831 2056 832
rect 2060 831 2061 835
rect 2055 830 2061 831
rect 2095 835 2101 836
rect 2095 831 2096 835
rect 2100 834 2101 835
rect 2103 835 2109 836
rect 2103 834 2104 835
rect 2100 832 2104 834
rect 2100 831 2101 832
rect 2095 830 2101 831
rect 2103 831 2104 832
rect 2108 831 2109 835
rect 2103 830 2109 831
rect 2118 832 2124 833
rect 1134 827 1140 828
rect 2118 828 2119 832
rect 2123 828 2124 832
rect 2118 827 2124 828
rect 934 826 940 827
rect 1158 824 1164 825
rect 828 820 882 822
rect 886 823 893 824
rect 828 819 829 820
rect 823 818 829 819
rect 886 819 887 823
rect 892 819 893 823
rect 886 818 893 819
rect 895 823 901 824
rect 895 819 896 823
rect 900 822 901 823
rect 951 823 957 824
rect 951 822 952 823
rect 900 820 952 822
rect 900 819 901 820
rect 895 818 901 819
rect 951 819 952 820
rect 956 819 957 823
rect 951 818 957 819
rect 959 823 965 824
rect 959 819 960 823
rect 964 822 965 823
rect 1023 823 1029 824
rect 1023 822 1024 823
rect 964 820 1024 822
rect 964 819 965 820
rect 959 818 965 819
rect 1023 819 1024 820
rect 1028 819 1029 823
rect 1023 818 1029 819
rect 1070 823 1077 824
rect 1070 819 1071 823
rect 1076 819 1077 823
rect 1158 820 1159 824
rect 1163 820 1164 824
rect 1158 819 1164 820
rect 1246 824 1252 825
rect 1246 820 1247 824
rect 1251 820 1252 824
rect 1246 819 1252 820
rect 1358 824 1364 825
rect 1358 820 1359 824
rect 1363 820 1364 824
rect 1358 819 1364 820
rect 1454 824 1460 825
rect 1454 820 1455 824
rect 1459 820 1460 824
rect 1454 819 1460 820
rect 1542 824 1548 825
rect 1542 820 1543 824
rect 1547 820 1548 824
rect 1542 819 1548 820
rect 1630 824 1636 825
rect 1630 820 1631 824
rect 1635 820 1636 824
rect 1630 819 1636 820
rect 1710 824 1716 825
rect 1710 820 1711 824
rect 1715 820 1716 824
rect 1710 819 1716 820
rect 1782 824 1788 825
rect 1782 820 1783 824
rect 1787 820 1788 824
rect 1782 819 1788 820
rect 1854 824 1860 825
rect 1854 820 1855 824
rect 1859 820 1860 824
rect 1854 819 1860 820
rect 1934 824 1940 825
rect 1934 820 1935 824
rect 1939 820 1940 824
rect 1934 819 1940 820
rect 2014 824 2020 825
rect 2014 820 2015 824
rect 2019 820 2020 824
rect 2014 819 2020 820
rect 2070 824 2076 825
rect 2070 820 2071 824
rect 2075 820 2076 824
rect 2070 819 2076 820
rect 1070 818 1077 819
rect 278 816 284 817
rect 278 812 279 816
rect 283 812 284 816
rect 278 811 284 812
rect 342 816 348 817
rect 342 812 343 816
rect 347 812 348 816
rect 342 811 348 812
rect 414 816 420 817
rect 414 812 415 816
rect 419 812 420 816
rect 414 811 420 812
rect 486 816 492 817
rect 486 812 487 816
rect 491 812 492 816
rect 486 811 492 812
rect 566 816 572 817
rect 566 812 567 816
rect 571 812 572 816
rect 566 811 572 812
rect 646 816 652 817
rect 646 812 647 816
rect 651 812 652 816
rect 646 811 652 812
rect 726 816 732 817
rect 726 812 727 816
rect 731 812 732 816
rect 726 811 732 812
rect 798 816 804 817
rect 798 812 799 816
rect 803 812 804 816
rect 798 811 804 812
rect 862 816 868 817
rect 862 812 863 816
rect 867 812 868 816
rect 862 811 868 812
rect 926 816 932 817
rect 926 812 927 816
rect 931 812 932 816
rect 926 811 932 812
rect 998 816 1004 817
rect 998 812 999 816
rect 1003 812 1004 816
rect 998 811 1004 812
rect 1046 816 1052 817
rect 1046 812 1047 816
rect 1051 812 1052 816
rect 1046 811 1052 812
rect 1182 815 1189 816
rect 1182 811 1183 815
rect 1188 811 1189 815
rect 1182 810 1189 811
rect 1262 815 1268 816
rect 1262 811 1263 815
rect 1267 814 1268 815
rect 1271 815 1277 816
rect 1271 814 1272 815
rect 1267 812 1272 814
rect 1267 811 1268 812
rect 1262 810 1268 811
rect 1271 811 1272 812
rect 1276 811 1277 815
rect 1271 810 1277 811
rect 1374 815 1380 816
rect 1374 811 1375 815
rect 1379 814 1380 815
rect 1383 815 1389 816
rect 1383 814 1384 815
rect 1379 812 1384 814
rect 1379 811 1380 812
rect 1374 810 1380 811
rect 1383 811 1384 812
rect 1388 811 1389 815
rect 1383 810 1389 811
rect 1479 815 1488 816
rect 1479 811 1480 815
rect 1487 811 1488 815
rect 1479 810 1488 811
rect 1567 815 1573 816
rect 1567 811 1568 815
rect 1572 814 1573 815
rect 1575 815 1581 816
rect 1575 814 1576 815
rect 1572 812 1576 814
rect 1572 811 1573 812
rect 1567 810 1573 811
rect 1575 811 1576 812
rect 1580 811 1581 815
rect 1575 810 1581 811
rect 1655 815 1661 816
rect 1655 811 1656 815
rect 1660 814 1661 815
rect 1663 815 1669 816
rect 1663 814 1664 815
rect 1660 812 1664 814
rect 1660 811 1661 812
rect 1655 810 1661 811
rect 1663 811 1664 812
rect 1668 811 1669 815
rect 1663 810 1669 811
rect 1734 815 1741 816
rect 1734 811 1735 815
rect 1740 811 1741 815
rect 1734 810 1741 811
rect 1807 815 1813 816
rect 1807 811 1808 815
rect 1812 814 1813 815
rect 1818 815 1824 816
rect 1818 814 1819 815
rect 1812 812 1819 814
rect 1812 811 1813 812
rect 1807 810 1813 811
rect 1818 811 1819 812
rect 1823 811 1824 815
rect 1818 810 1824 811
rect 1879 815 1885 816
rect 1879 811 1880 815
rect 1884 814 1885 815
rect 1887 815 1893 816
rect 1887 814 1888 815
rect 1884 812 1888 814
rect 1884 811 1885 812
rect 1879 810 1885 811
rect 1887 811 1888 812
rect 1892 811 1893 815
rect 1887 810 1893 811
rect 1910 815 1916 816
rect 1910 811 1911 815
rect 1915 814 1916 815
rect 1959 815 1965 816
rect 1959 814 1960 815
rect 1915 812 1960 814
rect 1915 811 1916 812
rect 1910 810 1916 811
rect 1959 811 1960 812
rect 1964 811 1965 815
rect 2039 815 2045 816
rect 2039 814 2040 815
rect 1959 810 1965 811
rect 1968 812 2040 814
rect 110 808 116 809
rect 110 804 111 808
rect 115 804 116 808
rect 1094 808 1100 809
rect 1094 804 1095 808
rect 1099 804 1100 808
rect 110 803 116 804
rect 303 803 309 804
rect 303 799 304 803
rect 308 802 309 803
rect 334 803 340 804
rect 334 802 335 803
rect 308 800 335 802
rect 308 799 309 800
rect 303 798 309 799
rect 334 799 335 800
rect 339 799 340 803
rect 334 798 340 799
rect 367 803 373 804
rect 367 799 368 803
rect 372 802 373 803
rect 375 803 381 804
rect 375 802 376 803
rect 372 800 376 802
rect 372 799 373 800
rect 367 798 373 799
rect 375 799 376 800
rect 380 799 381 803
rect 375 798 381 799
rect 439 803 448 804
rect 439 799 440 803
rect 447 799 448 803
rect 439 798 448 799
rect 506 803 517 804
rect 506 799 507 803
rect 511 799 512 803
rect 516 799 517 803
rect 506 798 517 799
rect 582 803 588 804
rect 582 799 583 803
rect 587 802 588 803
rect 591 803 597 804
rect 591 802 592 803
rect 587 800 592 802
rect 587 799 588 800
rect 582 798 588 799
rect 591 799 592 800
rect 596 799 597 803
rect 591 798 597 799
rect 662 803 668 804
rect 662 799 663 803
rect 667 802 668 803
rect 671 803 677 804
rect 671 802 672 803
rect 667 800 672 802
rect 667 799 668 800
rect 662 798 668 799
rect 671 799 672 800
rect 676 799 677 803
rect 671 798 677 799
rect 751 803 760 804
rect 751 799 752 803
rect 759 799 760 803
rect 751 798 760 799
rect 814 803 820 804
rect 814 799 815 803
rect 819 802 820 803
rect 823 803 829 804
rect 823 802 824 803
rect 819 800 824 802
rect 819 799 820 800
rect 814 798 820 799
rect 823 799 824 800
rect 828 799 829 803
rect 823 798 829 799
rect 887 803 893 804
rect 887 799 888 803
rect 892 802 893 803
rect 895 803 901 804
rect 895 802 896 803
rect 892 800 896 802
rect 892 799 893 800
rect 887 798 893 799
rect 895 799 896 800
rect 900 799 901 803
rect 895 798 901 799
rect 951 803 957 804
rect 951 799 952 803
rect 956 802 957 803
rect 959 803 965 804
rect 959 802 960 803
rect 956 800 960 802
rect 956 799 957 800
rect 951 798 957 799
rect 959 799 960 800
rect 964 799 965 803
rect 959 798 965 799
rect 1014 803 1020 804
rect 1014 799 1015 803
rect 1019 802 1020 803
rect 1023 803 1029 804
rect 1023 802 1024 803
rect 1019 800 1024 802
rect 1019 799 1020 800
rect 1014 798 1020 799
rect 1023 799 1024 800
rect 1028 799 1029 803
rect 1023 798 1029 799
rect 1071 803 1077 804
rect 1094 803 1100 804
rect 1894 807 1900 808
rect 1894 803 1895 807
rect 1899 806 1900 807
rect 1968 806 1970 812
rect 2039 811 2040 812
rect 2044 811 2045 815
rect 2039 810 2045 811
rect 2094 815 2101 816
rect 2094 811 2095 815
rect 2100 811 2101 815
rect 2094 810 2101 811
rect 1899 804 1970 806
rect 1899 803 1900 804
rect 1071 799 1072 803
rect 1076 799 1077 803
rect 1894 802 1900 803
rect 1071 798 1077 799
rect 1073 796 1187 798
rect 1183 795 1189 796
rect 110 791 116 792
rect 110 787 111 791
rect 115 787 116 791
rect 1094 791 1100 792
rect 110 786 116 787
rect 278 788 284 789
rect 278 784 279 788
rect 283 784 284 788
rect 278 783 284 784
rect 342 788 348 789
rect 342 784 343 788
rect 347 784 348 788
rect 342 783 348 784
rect 414 788 420 789
rect 414 784 415 788
rect 419 784 420 788
rect 414 783 420 784
rect 486 788 492 789
rect 486 784 487 788
rect 491 784 492 788
rect 486 783 492 784
rect 566 788 572 789
rect 566 784 567 788
rect 571 784 572 788
rect 566 783 572 784
rect 646 788 652 789
rect 646 784 647 788
rect 651 784 652 788
rect 646 783 652 784
rect 726 788 732 789
rect 726 784 727 788
rect 731 784 732 788
rect 726 783 732 784
rect 798 788 804 789
rect 798 784 799 788
rect 803 784 804 788
rect 798 783 804 784
rect 862 788 868 789
rect 862 784 863 788
rect 867 784 868 788
rect 862 783 868 784
rect 926 788 932 789
rect 926 784 927 788
rect 931 784 932 788
rect 926 783 932 784
rect 998 788 1004 789
rect 998 784 999 788
rect 1003 784 1004 788
rect 998 783 1004 784
rect 1046 788 1052 789
rect 1046 784 1047 788
rect 1051 784 1052 788
rect 1094 787 1095 791
rect 1099 787 1100 791
rect 1183 791 1184 795
rect 1188 791 1189 795
rect 1183 790 1189 791
rect 1303 795 1309 796
rect 1303 791 1304 795
rect 1308 794 1309 795
rect 1422 795 1428 796
rect 1422 794 1423 795
rect 1308 792 1423 794
rect 1308 791 1309 792
rect 1303 790 1309 791
rect 1422 791 1423 792
rect 1427 791 1428 795
rect 1422 790 1428 791
rect 1431 795 1437 796
rect 1431 791 1432 795
rect 1436 794 1437 795
rect 1462 795 1468 796
rect 1462 794 1463 795
rect 1436 792 1463 794
rect 1436 791 1437 792
rect 1431 790 1437 791
rect 1462 791 1463 792
rect 1467 791 1468 795
rect 1462 790 1468 791
rect 1543 795 1549 796
rect 1543 791 1544 795
rect 1548 794 1549 795
rect 1558 795 1564 796
rect 1558 794 1559 795
rect 1548 792 1559 794
rect 1548 791 1549 792
rect 1543 790 1549 791
rect 1558 791 1559 792
rect 1563 791 1564 795
rect 1558 790 1564 791
rect 1566 795 1572 796
rect 1566 791 1567 795
rect 1571 794 1572 795
rect 1647 795 1653 796
rect 1647 794 1648 795
rect 1571 792 1648 794
rect 1571 791 1572 792
rect 1566 790 1572 791
rect 1647 791 1648 792
rect 1652 791 1653 795
rect 1647 790 1653 791
rect 1655 795 1661 796
rect 1655 791 1656 795
rect 1660 794 1661 795
rect 1743 795 1749 796
rect 1743 794 1744 795
rect 1660 792 1744 794
rect 1660 791 1661 792
rect 1655 790 1661 791
rect 1743 791 1744 792
rect 1748 791 1749 795
rect 1743 790 1749 791
rect 1839 795 1845 796
rect 1839 791 1840 795
rect 1844 794 1845 795
rect 1918 795 1924 796
rect 1918 794 1919 795
rect 1844 792 1919 794
rect 1844 791 1845 792
rect 1839 790 1845 791
rect 1918 791 1919 792
rect 1923 791 1924 795
rect 1918 790 1924 791
rect 1927 795 1933 796
rect 1927 791 1928 795
rect 1932 794 1933 795
rect 1978 795 1984 796
rect 1978 794 1979 795
rect 1932 792 1979 794
rect 1932 791 1933 792
rect 1927 790 1933 791
rect 1978 791 1979 792
rect 1983 791 1984 795
rect 1978 790 1984 791
rect 1986 795 1992 796
rect 1986 791 1987 795
rect 1991 794 1992 795
rect 2023 795 2029 796
rect 2023 794 2024 795
rect 1991 792 2024 794
rect 1991 791 1992 792
rect 1986 790 1992 791
rect 2023 791 2024 792
rect 2028 791 2029 795
rect 2023 790 2029 791
rect 2095 795 2101 796
rect 2095 791 2096 795
rect 2100 794 2101 795
rect 2103 795 2109 796
rect 2103 794 2104 795
rect 2100 792 2104 794
rect 2100 791 2101 792
rect 2095 790 2101 791
rect 2103 791 2104 792
rect 2108 791 2109 795
rect 2103 790 2109 791
rect 1094 786 1100 787
rect 1158 788 1164 789
rect 1046 783 1052 784
rect 1158 784 1159 788
rect 1163 784 1164 788
rect 1158 783 1164 784
rect 1278 788 1284 789
rect 1278 784 1279 788
rect 1283 784 1284 788
rect 1278 783 1284 784
rect 1406 788 1412 789
rect 1406 784 1407 788
rect 1411 784 1412 788
rect 1406 783 1412 784
rect 1518 788 1524 789
rect 1518 784 1519 788
rect 1523 784 1524 788
rect 1518 783 1524 784
rect 1622 788 1628 789
rect 1622 784 1623 788
rect 1627 784 1628 788
rect 1622 783 1628 784
rect 1718 788 1724 789
rect 1718 784 1719 788
rect 1723 784 1724 788
rect 1718 783 1724 784
rect 1814 788 1820 789
rect 1814 784 1815 788
rect 1819 784 1820 788
rect 1814 783 1820 784
rect 1902 788 1908 789
rect 1902 784 1903 788
rect 1907 784 1908 788
rect 1902 783 1908 784
rect 1998 788 2004 789
rect 1998 784 1999 788
rect 2003 784 2004 788
rect 1998 783 2004 784
rect 2070 788 2076 789
rect 2070 784 2071 788
rect 2075 784 2076 788
rect 2070 783 2076 784
rect 1134 780 1140 781
rect 214 776 220 777
rect 110 773 116 774
rect 110 769 111 773
rect 115 769 116 773
rect 214 772 215 776
rect 219 772 220 776
rect 214 771 220 772
rect 278 776 284 777
rect 278 772 279 776
rect 283 772 284 776
rect 278 771 284 772
rect 350 776 356 777
rect 350 772 351 776
rect 355 772 356 776
rect 350 771 356 772
rect 422 776 428 777
rect 422 772 423 776
rect 427 772 428 776
rect 422 771 428 772
rect 494 776 500 777
rect 494 772 495 776
rect 499 772 500 776
rect 494 771 500 772
rect 566 776 572 777
rect 566 772 567 776
rect 571 772 572 776
rect 566 771 572 772
rect 638 776 644 777
rect 638 772 639 776
rect 643 772 644 776
rect 638 771 644 772
rect 702 776 708 777
rect 702 772 703 776
rect 707 772 708 776
rect 702 771 708 772
rect 758 776 764 777
rect 758 772 759 776
rect 763 772 764 776
rect 758 771 764 772
rect 814 776 820 777
rect 814 772 815 776
rect 819 772 820 776
rect 814 771 820 772
rect 862 776 868 777
rect 862 772 863 776
rect 867 772 868 776
rect 862 771 868 772
rect 910 776 916 777
rect 910 772 911 776
rect 915 772 916 776
rect 910 771 916 772
rect 958 776 964 777
rect 958 772 959 776
rect 963 772 964 776
rect 958 771 964 772
rect 1006 776 1012 777
rect 1006 772 1007 776
rect 1011 772 1012 776
rect 1006 771 1012 772
rect 1046 776 1052 777
rect 1046 772 1047 776
rect 1051 772 1052 776
rect 1134 776 1135 780
rect 1139 776 1140 780
rect 2118 780 2124 781
rect 2118 776 2119 780
rect 2123 776 2124 780
rect 1134 775 1140 776
rect 1182 775 1189 776
rect 1046 771 1052 772
rect 1094 773 1100 774
rect 110 768 116 769
rect 1094 769 1095 773
rect 1099 769 1100 773
rect 1182 771 1183 775
rect 1188 771 1189 775
rect 1182 770 1189 771
rect 1303 775 1309 776
rect 1303 771 1304 775
rect 1308 774 1309 775
rect 1399 775 1405 776
rect 1399 774 1400 775
rect 1308 772 1400 774
rect 1308 771 1309 772
rect 1303 770 1309 771
rect 1399 771 1400 772
rect 1404 771 1405 775
rect 1399 770 1405 771
rect 1422 775 1428 776
rect 1422 771 1423 775
rect 1427 774 1428 775
rect 1431 775 1437 776
rect 1431 774 1432 775
rect 1427 772 1432 774
rect 1427 771 1428 772
rect 1422 770 1428 771
rect 1431 771 1432 772
rect 1436 771 1437 775
rect 1431 770 1437 771
rect 1543 775 1549 776
rect 1543 771 1544 775
rect 1548 774 1549 775
rect 1566 775 1572 776
rect 1566 774 1567 775
rect 1548 772 1567 774
rect 1548 771 1549 772
rect 1543 770 1549 771
rect 1566 771 1567 772
rect 1571 771 1572 775
rect 1566 770 1572 771
rect 1647 775 1653 776
rect 1647 771 1648 775
rect 1652 774 1653 775
rect 1655 775 1661 776
rect 1655 774 1656 775
rect 1652 772 1656 774
rect 1652 771 1653 772
rect 1647 770 1653 771
rect 1655 771 1656 772
rect 1660 771 1661 775
rect 1655 770 1661 771
rect 1743 775 1749 776
rect 1743 771 1744 775
rect 1748 774 1749 775
rect 1822 775 1828 776
rect 1822 774 1823 775
rect 1748 772 1823 774
rect 1748 771 1749 772
rect 1743 770 1749 771
rect 1822 771 1823 772
rect 1827 771 1828 775
rect 1822 770 1828 771
rect 1839 775 1845 776
rect 1839 771 1840 775
rect 1844 774 1845 775
rect 1910 775 1916 776
rect 1910 774 1911 775
rect 1844 772 1911 774
rect 1844 771 1845 772
rect 1839 770 1845 771
rect 1910 771 1911 772
rect 1915 771 1916 775
rect 1910 770 1916 771
rect 1918 775 1924 776
rect 1918 771 1919 775
rect 1923 774 1924 775
rect 1927 775 1933 776
rect 1927 774 1928 775
rect 1923 772 1928 774
rect 1923 771 1924 772
rect 1918 770 1924 771
rect 1927 771 1928 772
rect 1932 771 1933 775
rect 1927 770 1933 771
rect 1978 775 1984 776
rect 1978 771 1979 775
rect 1983 774 1984 775
rect 2023 775 2029 776
rect 2023 774 2024 775
rect 1983 772 2024 774
rect 1983 771 1984 772
rect 1978 770 1984 771
rect 2023 771 2024 772
rect 2028 771 2029 775
rect 2023 770 2029 771
rect 2094 775 2101 776
rect 2118 775 2124 776
rect 2094 771 2095 775
rect 2100 771 2101 775
rect 2094 770 2101 771
rect 1094 768 1100 769
rect 670 767 676 768
rect 670 766 671 767
rect 633 764 671 766
rect 202 759 208 760
rect 110 756 116 757
rect 110 752 111 756
rect 115 752 116 756
rect 202 755 203 759
rect 207 758 208 759
rect 239 759 245 760
rect 239 758 240 759
rect 207 756 240 758
rect 207 755 208 756
rect 202 754 208 755
rect 239 755 240 756
rect 244 755 245 759
rect 239 754 245 755
rect 247 759 253 760
rect 247 755 248 759
rect 252 758 253 759
rect 303 759 309 760
rect 303 758 304 759
rect 252 756 304 758
rect 252 755 253 756
rect 247 754 253 755
rect 303 755 304 756
rect 308 755 309 759
rect 303 754 309 755
rect 311 759 317 760
rect 311 755 312 759
rect 316 758 317 759
rect 375 759 381 760
rect 375 758 376 759
rect 316 756 376 758
rect 316 755 317 756
rect 311 754 317 755
rect 375 755 376 756
rect 380 755 381 759
rect 375 754 381 755
rect 383 759 389 760
rect 383 755 384 759
rect 388 758 389 759
rect 447 759 453 760
rect 447 758 448 759
rect 388 756 448 758
rect 388 755 389 756
rect 383 754 389 755
rect 447 755 448 756
rect 452 755 453 759
rect 447 754 453 755
rect 519 759 525 760
rect 519 755 520 759
rect 524 758 525 759
rect 582 759 588 760
rect 582 758 583 759
rect 524 756 583 758
rect 524 755 525 756
rect 519 754 525 755
rect 582 755 583 756
rect 587 755 588 759
rect 582 754 588 755
rect 591 759 597 760
rect 591 755 592 759
rect 596 758 597 759
rect 633 758 635 764
rect 670 763 671 764
rect 675 763 676 767
rect 670 762 676 763
rect 886 767 892 768
rect 886 763 887 767
rect 891 766 892 767
rect 891 764 938 766
rect 891 763 892 764
rect 886 762 892 763
rect 936 760 938 764
rect 1134 763 1140 764
rect 596 756 635 758
rect 662 759 669 760
rect 596 755 597 756
rect 591 754 597 755
rect 662 755 663 759
rect 668 755 669 759
rect 662 754 669 755
rect 671 759 677 760
rect 671 755 672 759
rect 676 758 677 759
rect 727 759 733 760
rect 727 758 728 759
rect 676 756 728 758
rect 676 755 677 756
rect 671 754 677 755
rect 727 755 728 756
rect 732 755 733 759
rect 727 754 733 755
rect 750 759 756 760
rect 750 755 751 759
rect 755 758 756 759
rect 783 759 789 760
rect 783 758 784 759
rect 755 756 784 758
rect 755 755 756 756
rect 750 754 756 755
rect 783 755 784 756
rect 788 755 789 759
rect 783 754 789 755
rect 839 759 845 760
rect 839 755 840 759
rect 844 758 845 759
rect 878 759 884 760
rect 878 758 879 759
rect 844 756 879 758
rect 844 755 845 756
rect 839 754 845 755
rect 878 755 879 756
rect 883 755 884 759
rect 878 754 884 755
rect 887 759 893 760
rect 887 755 888 759
rect 892 758 893 759
rect 926 759 932 760
rect 926 758 927 759
rect 892 756 927 758
rect 892 755 893 756
rect 887 754 893 755
rect 926 755 927 756
rect 931 755 932 759
rect 926 754 932 755
rect 935 759 941 760
rect 935 755 936 759
rect 940 755 941 759
rect 935 754 941 755
rect 983 759 989 760
rect 983 755 984 759
rect 988 758 989 759
rect 1022 759 1028 760
rect 1022 758 1023 759
rect 988 756 1023 758
rect 988 755 989 756
rect 983 754 989 755
rect 1022 755 1023 756
rect 1027 755 1028 759
rect 1022 754 1028 755
rect 1031 759 1037 760
rect 1031 755 1032 759
rect 1036 758 1037 759
rect 1062 759 1068 760
rect 1062 758 1063 759
rect 1036 756 1063 758
rect 1036 755 1037 756
rect 1031 754 1037 755
rect 1062 755 1063 756
rect 1067 755 1068 759
rect 1062 754 1068 755
rect 1070 759 1077 760
rect 1070 755 1071 759
rect 1076 755 1077 759
rect 1134 759 1135 763
rect 1139 759 1140 763
rect 2118 763 2124 764
rect 1134 758 1140 759
rect 1158 760 1164 761
rect 1070 754 1077 755
rect 1094 756 1100 757
rect 110 751 116 752
rect 1094 752 1095 756
rect 1099 752 1100 756
rect 1158 756 1159 760
rect 1163 756 1164 760
rect 1158 755 1164 756
rect 1278 760 1284 761
rect 1278 756 1279 760
rect 1283 756 1284 760
rect 1278 755 1284 756
rect 1406 760 1412 761
rect 1406 756 1407 760
rect 1411 756 1412 760
rect 1406 755 1412 756
rect 1518 760 1524 761
rect 1518 756 1519 760
rect 1523 756 1524 760
rect 1518 755 1524 756
rect 1622 760 1628 761
rect 1622 756 1623 760
rect 1627 756 1628 760
rect 1622 755 1628 756
rect 1718 760 1724 761
rect 1718 756 1719 760
rect 1723 756 1724 760
rect 1718 755 1724 756
rect 1814 760 1820 761
rect 1814 756 1815 760
rect 1819 756 1820 760
rect 1814 755 1820 756
rect 1902 760 1908 761
rect 1902 756 1903 760
rect 1907 756 1908 760
rect 1902 755 1908 756
rect 1998 760 2004 761
rect 1998 756 1999 760
rect 2003 756 2004 760
rect 1998 755 2004 756
rect 2070 760 2076 761
rect 2070 756 2071 760
rect 2075 756 2076 760
rect 2118 759 2119 763
rect 2123 759 2124 763
rect 2118 758 2124 759
rect 2070 755 2076 756
rect 1094 751 1100 752
rect 214 748 220 749
rect 214 744 215 748
rect 219 744 220 748
rect 214 743 220 744
rect 278 748 284 749
rect 278 744 279 748
rect 283 744 284 748
rect 278 743 284 744
rect 350 748 356 749
rect 350 744 351 748
rect 355 744 356 748
rect 350 743 356 744
rect 422 748 428 749
rect 422 744 423 748
rect 427 744 428 748
rect 422 743 428 744
rect 494 748 500 749
rect 494 744 495 748
rect 499 744 500 748
rect 494 743 500 744
rect 566 748 572 749
rect 566 744 567 748
rect 571 744 572 748
rect 566 743 572 744
rect 638 748 644 749
rect 638 744 639 748
rect 643 744 644 748
rect 638 743 644 744
rect 702 748 708 749
rect 702 744 703 748
rect 707 744 708 748
rect 702 743 708 744
rect 758 748 764 749
rect 758 744 759 748
rect 763 744 764 748
rect 758 743 764 744
rect 814 748 820 749
rect 814 744 815 748
rect 819 744 820 748
rect 814 743 820 744
rect 862 748 868 749
rect 862 744 863 748
rect 867 744 868 748
rect 862 743 868 744
rect 910 748 916 749
rect 910 744 911 748
rect 915 744 916 748
rect 910 743 916 744
rect 958 748 964 749
rect 958 744 959 748
rect 963 744 964 748
rect 958 743 964 744
rect 1006 748 1012 749
rect 1006 744 1007 748
rect 1011 744 1012 748
rect 1006 743 1012 744
rect 1046 748 1052 749
rect 1046 744 1047 748
rect 1051 744 1052 748
rect 1046 743 1052 744
rect 1334 744 1340 745
rect 1134 741 1140 742
rect 239 739 245 740
rect 239 735 240 739
rect 244 738 245 739
rect 247 739 253 740
rect 247 738 248 739
rect 244 736 248 738
rect 244 735 245 736
rect 239 734 245 735
rect 247 735 248 736
rect 252 735 253 739
rect 247 734 253 735
rect 303 739 309 740
rect 303 735 304 739
rect 308 738 309 739
rect 311 739 317 740
rect 311 738 312 739
rect 308 736 312 738
rect 308 735 309 736
rect 303 734 309 735
rect 311 735 312 736
rect 316 735 317 739
rect 311 734 317 735
rect 375 739 381 740
rect 375 735 376 739
rect 380 738 381 739
rect 383 739 389 740
rect 383 738 384 739
rect 380 736 384 738
rect 380 735 381 736
rect 375 734 381 735
rect 383 735 384 736
rect 388 735 389 739
rect 383 734 389 735
rect 442 739 453 740
rect 442 735 443 739
rect 447 735 448 739
rect 452 735 453 739
rect 442 734 453 735
rect 519 739 525 740
rect 519 735 520 739
rect 524 738 525 739
rect 558 739 564 740
rect 558 738 559 739
rect 524 736 559 738
rect 524 735 525 736
rect 519 734 525 735
rect 558 735 559 736
rect 563 735 564 739
rect 558 734 564 735
rect 582 739 588 740
rect 582 735 583 739
rect 587 738 588 739
rect 591 739 597 740
rect 591 738 592 739
rect 587 736 592 738
rect 587 735 588 736
rect 582 734 588 735
rect 591 735 592 736
rect 596 735 597 739
rect 591 734 597 735
rect 663 739 669 740
rect 663 735 664 739
rect 668 738 669 739
rect 671 739 677 740
rect 671 738 672 739
rect 668 736 672 738
rect 668 735 669 736
rect 663 734 669 735
rect 671 735 672 736
rect 676 735 677 739
rect 671 734 677 735
rect 727 739 733 740
rect 727 735 728 739
rect 732 738 733 739
rect 750 739 756 740
rect 750 738 751 739
rect 732 736 751 738
rect 732 735 733 736
rect 727 734 733 735
rect 750 735 751 736
rect 755 735 756 739
rect 750 734 756 735
rect 783 739 789 740
rect 783 735 784 739
rect 788 738 789 739
rect 822 739 828 740
rect 822 738 823 739
rect 788 736 823 738
rect 788 735 789 736
rect 783 734 789 735
rect 822 735 823 736
rect 827 735 828 739
rect 822 734 828 735
rect 839 739 845 740
rect 839 735 840 739
rect 844 735 845 739
rect 839 734 845 735
rect 878 739 884 740
rect 878 735 879 739
rect 883 738 884 739
rect 887 739 893 740
rect 887 738 888 739
rect 883 736 888 738
rect 883 735 884 736
rect 878 734 884 735
rect 887 735 888 736
rect 892 735 893 739
rect 887 734 893 735
rect 926 739 932 740
rect 926 735 927 739
rect 931 738 932 739
rect 935 739 941 740
rect 935 738 936 739
rect 931 736 936 738
rect 931 735 932 736
rect 926 734 932 735
rect 935 735 936 736
rect 940 735 941 739
rect 935 734 941 735
rect 983 739 989 740
rect 983 735 984 739
rect 988 738 989 739
rect 1014 739 1020 740
rect 1014 738 1015 739
rect 988 736 1015 738
rect 988 735 989 736
rect 983 734 989 735
rect 1014 735 1015 736
rect 1019 735 1020 739
rect 1014 734 1020 735
rect 1022 739 1028 740
rect 1022 735 1023 739
rect 1027 738 1028 739
rect 1031 739 1037 740
rect 1031 738 1032 739
rect 1027 736 1032 738
rect 1027 735 1028 736
rect 1022 734 1028 735
rect 1031 735 1032 736
rect 1036 735 1037 739
rect 1031 734 1037 735
rect 1062 739 1068 740
rect 1062 735 1063 739
rect 1067 738 1068 739
rect 1071 739 1077 740
rect 1071 738 1072 739
rect 1067 736 1072 738
rect 1067 735 1068 736
rect 1062 734 1068 735
rect 1071 735 1072 736
rect 1076 735 1077 739
rect 1134 737 1135 741
rect 1139 737 1140 741
rect 1334 740 1335 744
rect 1339 740 1340 744
rect 1334 739 1340 740
rect 1374 744 1380 745
rect 1374 740 1375 744
rect 1379 740 1380 744
rect 1374 739 1380 740
rect 1414 744 1420 745
rect 1414 740 1415 744
rect 1419 740 1420 744
rect 1414 739 1420 740
rect 1454 744 1460 745
rect 1454 740 1455 744
rect 1459 740 1460 744
rect 1454 739 1460 740
rect 1502 744 1508 745
rect 1502 740 1503 744
rect 1507 740 1508 744
rect 1502 739 1508 740
rect 1550 744 1556 745
rect 1550 740 1551 744
rect 1555 740 1556 744
rect 1550 739 1556 740
rect 1598 744 1604 745
rect 1598 740 1599 744
rect 1603 740 1604 744
rect 1598 739 1604 740
rect 1654 744 1660 745
rect 1654 740 1655 744
rect 1659 740 1660 744
rect 1654 739 1660 740
rect 1710 744 1716 745
rect 1710 740 1711 744
rect 1715 740 1716 744
rect 1710 739 1716 740
rect 1766 744 1772 745
rect 1766 740 1767 744
rect 1771 740 1772 744
rect 1766 739 1772 740
rect 1830 744 1836 745
rect 1830 740 1831 744
rect 1835 740 1836 744
rect 1830 739 1836 740
rect 1894 744 1900 745
rect 1894 740 1895 744
rect 1899 740 1900 744
rect 1894 739 1900 740
rect 1958 744 1964 745
rect 1958 740 1959 744
rect 1963 740 1964 744
rect 1958 739 1964 740
rect 2022 744 2028 745
rect 2022 740 2023 744
rect 2027 740 2028 744
rect 2022 739 2028 740
rect 2070 744 2076 745
rect 2070 740 2071 744
rect 2075 740 2076 744
rect 2070 739 2076 740
rect 2118 741 2124 742
rect 1134 736 1140 737
rect 2118 737 2119 741
rect 2123 737 2124 741
rect 2118 736 2124 737
rect 1071 734 1077 735
rect 1399 735 1405 736
rect 662 731 668 732
rect 662 727 663 731
rect 667 730 668 731
rect 841 730 843 734
rect 1399 731 1400 735
rect 1404 734 1405 735
rect 1622 735 1628 736
rect 1622 734 1623 735
rect 1404 732 1623 734
rect 1404 731 1405 732
rect 1399 730 1405 731
rect 1622 731 1623 732
rect 1627 731 1628 735
rect 1622 730 1628 731
rect 667 728 843 730
rect 667 727 668 728
rect 662 726 668 727
rect 1359 727 1368 728
rect 769 724 955 726
rect 767 723 773 724
rect 199 719 208 720
rect 199 715 200 719
rect 207 715 208 719
rect 199 714 208 715
rect 210 719 216 720
rect 210 715 211 719
rect 215 718 216 719
rect 263 719 269 720
rect 263 718 264 719
rect 215 716 264 718
rect 215 715 216 716
rect 210 714 216 715
rect 263 715 264 716
rect 268 715 269 719
rect 263 714 269 715
rect 271 719 277 720
rect 271 715 272 719
rect 276 718 277 719
rect 335 719 341 720
rect 335 718 336 719
rect 276 716 336 718
rect 276 715 277 716
rect 271 714 277 715
rect 335 715 336 716
rect 340 715 341 719
rect 335 714 341 715
rect 415 719 424 720
rect 415 715 416 719
rect 423 715 424 719
rect 415 714 424 715
rect 426 719 432 720
rect 426 715 427 719
rect 431 718 432 719
rect 495 719 501 720
rect 495 718 496 719
rect 431 716 496 718
rect 431 715 432 716
rect 426 714 432 715
rect 495 715 496 716
rect 500 715 501 719
rect 495 714 501 715
rect 503 719 509 720
rect 503 715 504 719
rect 508 718 509 719
rect 567 719 573 720
rect 567 718 568 719
rect 508 716 568 718
rect 508 715 509 716
rect 503 714 509 715
rect 567 715 568 716
rect 572 715 573 719
rect 567 714 573 715
rect 639 719 645 720
rect 639 715 640 719
rect 644 718 645 719
rect 694 719 700 720
rect 694 718 695 719
rect 644 716 695 718
rect 644 715 645 716
rect 639 714 645 715
rect 694 715 695 716
rect 699 715 700 719
rect 694 714 700 715
rect 703 719 709 720
rect 703 715 704 719
rect 708 718 709 719
rect 726 719 732 720
rect 726 718 727 719
rect 708 716 727 718
rect 708 715 709 716
rect 703 714 709 715
rect 726 715 727 716
rect 731 715 732 719
rect 759 719 765 720
rect 759 718 760 719
rect 726 714 732 715
rect 744 716 760 718
rect 174 712 180 713
rect 174 708 175 712
rect 179 708 180 712
rect 174 707 180 708
rect 238 712 244 713
rect 238 708 239 712
rect 243 708 244 712
rect 238 707 244 708
rect 310 712 316 713
rect 310 708 311 712
rect 315 708 316 712
rect 310 707 316 708
rect 390 712 396 713
rect 390 708 391 712
rect 395 708 396 712
rect 390 707 396 708
rect 470 712 476 713
rect 470 708 471 712
rect 475 708 476 712
rect 470 707 476 708
rect 542 712 548 713
rect 542 708 543 712
rect 547 708 548 712
rect 542 707 548 708
rect 614 712 620 713
rect 614 708 615 712
rect 619 708 620 712
rect 614 707 620 708
rect 678 712 684 713
rect 678 708 679 712
rect 683 708 684 712
rect 678 707 684 708
rect 734 712 740 713
rect 734 708 735 712
rect 739 708 740 712
rect 734 707 740 708
rect 110 704 116 705
rect 110 700 111 704
rect 115 700 116 704
rect 688 704 714 706
rect 688 702 690 704
rect 641 700 690 702
rect 712 702 714 704
rect 744 702 746 716
rect 759 715 760 716
rect 764 715 765 719
rect 767 719 768 723
rect 772 719 773 723
rect 953 720 955 724
rect 1134 724 1140 725
rect 1134 720 1135 724
rect 1139 720 1140 724
rect 1359 723 1360 727
rect 1367 723 1368 727
rect 1359 722 1368 723
rect 1382 727 1388 728
rect 1382 723 1383 727
rect 1387 726 1388 727
rect 1399 727 1405 728
rect 1399 726 1400 727
rect 1387 724 1400 726
rect 1387 723 1388 724
rect 1382 722 1388 723
rect 1399 723 1400 724
rect 1404 723 1405 727
rect 1399 722 1405 723
rect 1422 727 1428 728
rect 1422 723 1423 727
rect 1427 726 1428 727
rect 1439 727 1445 728
rect 1439 726 1440 727
rect 1427 724 1440 726
rect 1427 723 1428 724
rect 1422 722 1428 723
rect 1439 723 1440 724
rect 1444 723 1445 727
rect 1439 722 1445 723
rect 1462 727 1468 728
rect 1462 723 1463 727
rect 1467 726 1468 727
rect 1479 727 1485 728
rect 1479 726 1480 727
rect 1467 724 1480 726
rect 1467 723 1468 724
rect 1462 722 1468 723
rect 1479 723 1480 724
rect 1484 723 1485 727
rect 1479 722 1485 723
rect 1487 727 1493 728
rect 1487 723 1488 727
rect 1492 726 1493 727
rect 1527 727 1533 728
rect 1527 726 1528 727
rect 1492 724 1528 726
rect 1492 723 1493 724
rect 1487 722 1493 723
rect 1527 723 1528 724
rect 1532 723 1533 727
rect 1527 722 1533 723
rect 1535 727 1541 728
rect 1535 723 1536 727
rect 1540 726 1541 727
rect 1575 727 1581 728
rect 1575 726 1576 727
rect 1540 724 1576 726
rect 1540 723 1541 724
rect 1535 722 1541 723
rect 1575 723 1576 724
rect 1580 723 1581 727
rect 1575 722 1581 723
rect 1583 727 1589 728
rect 1583 723 1584 727
rect 1588 726 1589 727
rect 1623 727 1629 728
rect 1623 726 1624 727
rect 1588 724 1624 726
rect 1588 723 1589 724
rect 1583 722 1589 723
rect 1623 723 1624 724
rect 1628 723 1629 727
rect 1623 722 1629 723
rect 1678 727 1685 728
rect 1678 723 1679 727
rect 1684 723 1685 727
rect 1678 722 1685 723
rect 1687 727 1693 728
rect 1687 723 1688 727
rect 1692 726 1693 727
rect 1735 727 1741 728
rect 1735 726 1736 727
rect 1692 724 1736 726
rect 1692 723 1693 724
rect 1687 722 1693 723
rect 1735 723 1736 724
rect 1740 723 1741 727
rect 1735 722 1741 723
rect 1758 727 1764 728
rect 1758 723 1759 727
rect 1763 726 1764 727
rect 1791 727 1797 728
rect 1791 726 1792 727
rect 1763 724 1792 726
rect 1763 723 1764 724
rect 1758 722 1764 723
rect 1791 723 1792 724
rect 1796 723 1797 727
rect 1791 722 1797 723
rect 1799 727 1805 728
rect 1799 723 1800 727
rect 1804 726 1805 727
rect 1855 727 1861 728
rect 1855 726 1856 727
rect 1804 724 1856 726
rect 1804 723 1805 724
rect 1799 722 1805 723
rect 1855 723 1856 724
rect 1860 723 1861 727
rect 1855 722 1861 723
rect 1919 727 1925 728
rect 1919 723 1920 727
rect 1924 726 1925 727
rect 1974 727 1980 728
rect 1974 726 1975 727
rect 1924 724 1975 726
rect 1924 723 1925 724
rect 1919 722 1925 723
rect 1974 723 1975 724
rect 1979 723 1980 727
rect 1974 722 1980 723
rect 1983 727 1992 728
rect 1983 723 1984 727
rect 1991 723 1992 727
rect 1983 722 1992 723
rect 2046 727 2053 728
rect 2046 723 2047 727
rect 2052 723 2053 727
rect 2046 722 2053 723
rect 2055 727 2061 728
rect 2055 723 2056 727
rect 2060 726 2061 727
rect 2095 727 2101 728
rect 2095 726 2096 727
rect 2060 724 2096 726
rect 2060 723 2061 724
rect 2055 722 2061 723
rect 2095 723 2096 724
rect 2100 723 2101 727
rect 2095 722 2101 723
rect 2118 724 2124 725
rect 767 718 773 719
rect 823 719 829 720
rect 759 714 765 715
rect 823 715 824 719
rect 828 718 829 719
rect 878 719 884 720
rect 878 718 879 719
rect 828 716 879 718
rect 828 715 829 716
rect 823 714 829 715
rect 878 715 879 716
rect 883 715 884 719
rect 878 714 884 715
rect 887 719 893 720
rect 887 715 888 719
rect 892 718 893 719
rect 942 719 948 720
rect 942 718 943 719
rect 892 716 943 718
rect 892 715 893 716
rect 887 714 893 715
rect 942 715 943 716
rect 947 715 948 719
rect 942 714 948 715
rect 951 719 957 720
rect 1134 719 1140 720
rect 2118 720 2119 724
rect 2123 720 2124 724
rect 2118 719 2124 720
rect 951 715 952 719
rect 956 715 957 719
rect 951 714 957 715
rect 1334 716 1340 717
rect 798 712 804 713
rect 798 708 799 712
rect 803 708 804 712
rect 798 707 804 708
rect 862 712 868 713
rect 862 708 863 712
rect 867 708 868 712
rect 862 707 868 708
rect 926 712 932 713
rect 926 708 927 712
rect 931 708 932 712
rect 1334 712 1335 716
rect 1339 712 1340 716
rect 1334 711 1340 712
rect 1374 716 1380 717
rect 1374 712 1375 716
rect 1379 712 1380 716
rect 1374 711 1380 712
rect 1414 716 1420 717
rect 1414 712 1415 716
rect 1419 712 1420 716
rect 1414 711 1420 712
rect 1454 716 1460 717
rect 1454 712 1455 716
rect 1459 712 1460 716
rect 1454 711 1460 712
rect 1502 716 1508 717
rect 1502 712 1503 716
rect 1507 712 1508 716
rect 1502 711 1508 712
rect 1550 716 1556 717
rect 1550 712 1551 716
rect 1555 712 1556 716
rect 1550 711 1556 712
rect 1598 716 1604 717
rect 1598 712 1599 716
rect 1603 712 1604 716
rect 1598 711 1604 712
rect 1654 716 1660 717
rect 1654 712 1655 716
rect 1659 712 1660 716
rect 1654 711 1660 712
rect 1710 716 1716 717
rect 1710 712 1711 716
rect 1715 712 1716 716
rect 1710 711 1716 712
rect 1766 716 1772 717
rect 1766 712 1767 716
rect 1771 712 1772 716
rect 1766 711 1772 712
rect 1830 716 1836 717
rect 1830 712 1831 716
rect 1835 712 1836 716
rect 1830 711 1836 712
rect 1894 716 1900 717
rect 1894 712 1895 716
rect 1899 712 1900 716
rect 1894 711 1900 712
rect 1958 716 1964 717
rect 1958 712 1959 716
rect 1963 712 1964 716
rect 1958 711 1964 712
rect 2022 716 2028 717
rect 2022 712 2023 716
rect 2027 712 2028 716
rect 2022 711 2028 712
rect 2070 716 2076 717
rect 2070 712 2071 716
rect 2075 712 2076 716
rect 2070 711 2076 712
rect 926 707 932 708
rect 1359 707 1365 708
rect 712 700 746 702
rect 1094 704 1100 705
rect 1094 700 1095 704
rect 1099 700 1100 704
rect 1359 703 1360 707
rect 1364 706 1365 707
rect 1382 707 1388 708
rect 1382 706 1383 707
rect 1364 704 1383 706
rect 1364 703 1365 704
rect 1359 702 1365 703
rect 1382 703 1383 704
rect 1387 703 1388 707
rect 1382 702 1388 703
rect 1399 707 1405 708
rect 1399 703 1400 707
rect 1404 706 1405 707
rect 1422 707 1428 708
rect 1422 706 1423 707
rect 1404 704 1423 706
rect 1404 703 1405 704
rect 1399 702 1405 703
rect 1422 703 1423 704
rect 1427 703 1428 707
rect 1422 702 1428 703
rect 1439 707 1445 708
rect 1439 703 1440 707
rect 1444 706 1445 707
rect 1462 707 1468 708
rect 1462 706 1463 707
rect 1444 704 1463 706
rect 1444 703 1445 704
rect 1439 702 1445 703
rect 1462 703 1463 704
rect 1467 703 1468 707
rect 1462 702 1468 703
rect 1479 707 1485 708
rect 1479 703 1480 707
rect 1484 706 1485 707
rect 1487 707 1493 708
rect 1487 706 1488 707
rect 1484 704 1488 706
rect 1484 703 1485 704
rect 1479 702 1485 703
rect 1487 703 1488 704
rect 1492 703 1493 707
rect 1487 702 1493 703
rect 1527 707 1533 708
rect 1527 703 1528 707
rect 1532 706 1533 707
rect 1535 707 1541 708
rect 1535 706 1536 707
rect 1532 704 1536 706
rect 1532 703 1533 704
rect 1527 702 1533 703
rect 1535 703 1536 704
rect 1540 703 1541 707
rect 1535 702 1541 703
rect 1575 707 1581 708
rect 1575 703 1576 707
rect 1580 706 1581 707
rect 1583 707 1589 708
rect 1583 706 1584 707
rect 1580 704 1584 706
rect 1580 703 1581 704
rect 1575 702 1581 703
rect 1583 703 1584 704
rect 1588 703 1589 707
rect 1583 702 1589 703
rect 1622 707 1629 708
rect 1622 703 1623 707
rect 1628 703 1629 707
rect 1622 702 1629 703
rect 1679 707 1685 708
rect 1679 703 1680 707
rect 1684 706 1685 707
rect 1687 707 1693 708
rect 1687 706 1688 707
rect 1684 704 1688 706
rect 1684 703 1685 704
rect 1679 702 1685 703
rect 1687 703 1688 704
rect 1692 703 1693 707
rect 1687 702 1693 703
rect 1735 707 1741 708
rect 1735 703 1736 707
rect 1740 706 1741 707
rect 1758 707 1764 708
rect 1758 706 1759 707
rect 1740 704 1759 706
rect 1740 703 1741 704
rect 1735 702 1741 703
rect 1758 703 1759 704
rect 1763 703 1764 707
rect 1758 702 1764 703
rect 1791 707 1797 708
rect 1791 703 1792 707
rect 1796 706 1797 707
rect 1799 707 1805 708
rect 1799 706 1800 707
rect 1796 704 1800 706
rect 1796 703 1797 704
rect 1791 702 1797 703
rect 1799 703 1800 704
rect 1804 703 1805 707
rect 1799 702 1805 703
rect 1822 707 1828 708
rect 1822 703 1823 707
rect 1827 706 1828 707
rect 1855 707 1861 708
rect 1855 706 1856 707
rect 1827 704 1856 706
rect 1827 703 1828 704
rect 1822 702 1828 703
rect 1855 703 1856 704
rect 1860 703 1861 707
rect 1855 702 1861 703
rect 1919 707 1925 708
rect 1919 703 1920 707
rect 1924 706 1925 707
rect 1934 707 1940 708
rect 1934 706 1935 707
rect 1924 704 1935 706
rect 1924 703 1925 704
rect 1919 702 1925 703
rect 1934 703 1935 704
rect 1939 703 1940 707
rect 1934 702 1940 703
rect 1974 707 1980 708
rect 1974 703 1975 707
rect 1979 706 1980 707
rect 1983 707 1989 708
rect 1983 706 1984 707
rect 1979 704 1984 706
rect 1979 703 1980 704
rect 1974 702 1980 703
rect 1983 703 1984 704
rect 1988 703 1989 707
rect 1983 702 1989 703
rect 2047 707 2053 708
rect 2047 703 2048 707
rect 2052 706 2053 707
rect 2055 707 2061 708
rect 2055 706 2056 707
rect 2052 704 2056 706
rect 2052 703 2053 704
rect 2047 702 2053 703
rect 2055 703 2056 704
rect 2060 703 2061 707
rect 2055 702 2061 703
rect 2094 707 2101 708
rect 2094 703 2095 707
rect 2100 703 2101 707
rect 2094 702 2101 703
rect 110 699 116 700
rect 199 699 205 700
rect 199 695 200 699
rect 204 698 205 699
rect 210 699 216 700
rect 210 698 211 699
rect 204 696 211 698
rect 204 695 205 696
rect 199 694 205 695
rect 210 695 211 696
rect 215 695 216 699
rect 210 694 216 695
rect 263 699 269 700
rect 263 695 264 699
rect 268 698 269 699
rect 271 699 277 700
rect 271 698 272 699
rect 268 696 272 698
rect 268 695 269 696
rect 263 694 269 695
rect 271 695 272 696
rect 276 695 277 699
rect 271 694 277 695
rect 298 699 304 700
rect 298 695 299 699
rect 303 698 304 699
rect 335 699 341 700
rect 335 698 336 699
rect 303 696 336 698
rect 303 695 304 696
rect 298 694 304 695
rect 335 695 336 696
rect 340 695 341 699
rect 335 694 341 695
rect 415 699 421 700
rect 415 695 416 699
rect 420 698 421 699
rect 426 699 432 700
rect 426 698 427 699
rect 420 696 427 698
rect 420 695 421 696
rect 415 694 421 695
rect 426 695 427 696
rect 431 695 432 699
rect 426 694 432 695
rect 495 699 501 700
rect 495 695 496 699
rect 500 698 501 699
rect 503 699 509 700
rect 503 698 504 699
rect 500 696 504 698
rect 500 695 501 696
rect 495 694 501 695
rect 503 695 504 696
rect 508 695 509 699
rect 503 694 509 695
rect 558 699 564 700
rect 558 695 559 699
rect 563 698 564 699
rect 567 699 573 700
rect 567 698 568 699
rect 563 696 568 698
rect 563 695 564 696
rect 558 694 564 695
rect 567 695 568 696
rect 572 695 573 699
rect 567 694 573 695
rect 639 699 645 700
rect 639 695 640 699
rect 644 695 645 699
rect 639 694 645 695
rect 694 699 700 700
rect 694 695 695 699
rect 699 698 700 699
rect 703 699 709 700
rect 703 698 704 699
rect 699 696 704 698
rect 699 695 700 696
rect 694 694 700 695
rect 703 695 704 696
rect 708 695 709 699
rect 703 694 709 695
rect 759 699 765 700
rect 759 695 760 699
rect 764 698 765 699
rect 767 699 773 700
rect 767 698 768 699
rect 764 696 768 698
rect 764 695 765 696
rect 759 694 765 695
rect 767 695 768 696
rect 772 695 773 699
rect 767 694 773 695
rect 822 699 829 700
rect 822 695 823 699
rect 828 695 829 699
rect 822 694 829 695
rect 878 699 884 700
rect 878 695 879 699
rect 883 698 884 699
rect 887 699 893 700
rect 887 698 888 699
rect 883 696 888 698
rect 883 695 884 696
rect 878 694 884 695
rect 887 695 888 696
rect 892 695 893 699
rect 887 694 893 695
rect 942 699 948 700
rect 942 695 943 699
rect 947 698 948 699
rect 951 699 957 700
rect 1094 699 1100 700
rect 951 698 952 699
rect 947 696 952 698
rect 947 695 948 696
rect 942 694 948 695
rect 951 695 952 696
rect 956 695 957 699
rect 951 694 957 695
rect 1362 695 1368 696
rect 1362 691 1363 695
rect 1367 694 1368 695
rect 1678 695 1684 696
rect 1367 692 1539 694
rect 1367 691 1368 692
rect 1362 690 1368 691
rect 1537 688 1539 692
rect 1678 691 1679 695
rect 1683 694 1684 695
rect 1946 695 1952 696
rect 1683 692 1851 694
rect 1683 691 1684 692
rect 1678 690 1684 691
rect 1849 688 1851 692
rect 1946 691 1947 695
rect 1951 694 1952 695
rect 1951 692 2001 694
rect 1951 691 1952 692
rect 1946 690 1952 691
rect 110 687 116 688
rect 110 683 111 687
rect 115 683 116 687
rect 1094 687 1100 688
rect 110 682 116 683
rect 174 684 180 685
rect 174 680 175 684
rect 179 680 180 684
rect 174 679 180 680
rect 238 684 244 685
rect 238 680 239 684
rect 243 680 244 684
rect 238 679 244 680
rect 310 684 316 685
rect 310 680 311 684
rect 315 680 316 684
rect 310 679 316 680
rect 390 684 396 685
rect 390 680 391 684
rect 395 680 396 684
rect 390 679 396 680
rect 470 684 476 685
rect 470 680 471 684
rect 475 680 476 684
rect 470 679 476 680
rect 542 684 548 685
rect 542 680 543 684
rect 547 680 548 684
rect 542 679 548 680
rect 614 684 620 685
rect 614 680 615 684
rect 619 680 620 684
rect 614 679 620 680
rect 678 684 684 685
rect 678 680 679 684
rect 683 680 684 684
rect 678 679 684 680
rect 734 684 740 685
rect 734 680 735 684
rect 739 680 740 684
rect 734 679 740 680
rect 798 684 804 685
rect 798 680 799 684
rect 803 680 804 684
rect 798 679 804 680
rect 862 684 868 685
rect 862 680 863 684
rect 867 680 868 684
rect 862 679 868 680
rect 926 684 932 685
rect 926 680 927 684
rect 931 680 932 684
rect 1094 683 1095 687
rect 1099 683 1100 687
rect 1094 682 1100 683
rect 1271 687 1277 688
rect 1271 683 1272 687
rect 1276 686 1277 687
rect 1302 687 1308 688
rect 1302 686 1303 687
rect 1276 684 1303 686
rect 1276 683 1277 684
rect 1271 682 1277 683
rect 1302 683 1303 684
rect 1307 683 1308 687
rect 1302 682 1308 683
rect 1311 687 1317 688
rect 1311 683 1312 687
rect 1316 686 1317 687
rect 1350 687 1356 688
rect 1350 686 1351 687
rect 1316 684 1351 686
rect 1316 683 1317 684
rect 1311 682 1317 683
rect 1350 683 1351 684
rect 1355 683 1356 687
rect 1350 682 1356 683
rect 1359 687 1365 688
rect 1359 683 1360 687
rect 1364 686 1365 687
rect 1406 687 1412 688
rect 1406 686 1407 687
rect 1364 684 1407 686
rect 1364 683 1365 684
rect 1359 682 1365 683
rect 1406 683 1407 684
rect 1411 683 1412 687
rect 1406 682 1412 683
rect 1415 687 1421 688
rect 1415 683 1416 687
rect 1420 686 1421 687
rect 1462 687 1468 688
rect 1462 686 1463 687
rect 1420 684 1463 686
rect 1420 683 1421 684
rect 1415 682 1421 683
rect 1462 683 1463 684
rect 1467 683 1468 687
rect 1462 682 1468 683
rect 1471 687 1477 688
rect 1471 683 1472 687
rect 1476 686 1477 687
rect 1526 687 1532 688
rect 1526 686 1527 687
rect 1476 684 1527 686
rect 1476 683 1477 684
rect 1471 682 1477 683
rect 1526 683 1527 684
rect 1531 683 1532 687
rect 1526 682 1532 683
rect 1535 687 1541 688
rect 1535 683 1536 687
rect 1540 683 1541 687
rect 1535 682 1541 683
rect 1607 687 1613 688
rect 1607 683 1608 687
rect 1612 686 1613 687
rect 1670 687 1676 688
rect 1670 686 1671 687
rect 1612 684 1671 686
rect 1612 683 1613 684
rect 1607 682 1613 683
rect 1670 683 1671 684
rect 1675 683 1676 687
rect 1670 682 1676 683
rect 1679 687 1685 688
rect 1679 683 1680 687
rect 1684 686 1685 687
rect 1718 687 1724 688
rect 1718 686 1719 687
rect 1684 684 1719 686
rect 1684 683 1685 684
rect 1679 682 1685 683
rect 1718 683 1719 684
rect 1723 683 1724 687
rect 1718 682 1724 683
rect 1759 687 1765 688
rect 1759 683 1760 687
rect 1764 686 1765 687
rect 1838 687 1844 688
rect 1838 686 1839 687
rect 1764 684 1839 686
rect 1764 683 1765 684
rect 1759 682 1765 683
rect 1838 683 1839 684
rect 1843 683 1844 687
rect 1838 682 1844 683
rect 1847 687 1853 688
rect 1847 683 1848 687
rect 1852 683 1853 687
rect 1847 682 1853 683
rect 1935 687 1941 688
rect 1935 683 1936 687
rect 1940 686 1941 687
rect 1999 686 2001 692
rect 2023 687 2029 688
rect 2023 686 2024 687
rect 1940 684 1982 686
rect 1999 684 2024 686
rect 1940 683 1941 684
rect 1935 682 1941 683
rect 926 679 932 680
rect 1246 680 1252 681
rect 1246 676 1247 680
rect 1251 676 1252 680
rect 1246 675 1252 676
rect 1286 680 1292 681
rect 1286 676 1287 680
rect 1291 676 1292 680
rect 1286 675 1292 676
rect 1334 680 1340 681
rect 1334 676 1335 680
rect 1339 676 1340 680
rect 1334 675 1340 676
rect 1390 680 1396 681
rect 1390 676 1391 680
rect 1395 676 1396 680
rect 1390 675 1396 676
rect 1446 680 1452 681
rect 1446 676 1447 680
rect 1451 676 1452 680
rect 1446 675 1452 676
rect 1510 680 1516 681
rect 1510 676 1511 680
rect 1515 676 1516 680
rect 1510 675 1516 676
rect 1582 680 1588 681
rect 1582 676 1583 680
rect 1587 676 1588 680
rect 1582 675 1588 676
rect 1654 680 1660 681
rect 1654 676 1655 680
rect 1659 676 1660 680
rect 1654 675 1660 676
rect 1734 680 1740 681
rect 1734 676 1735 680
rect 1739 676 1740 680
rect 1734 675 1740 676
rect 1822 680 1828 681
rect 1822 676 1823 680
rect 1827 676 1828 680
rect 1822 675 1828 676
rect 1910 680 1916 681
rect 1910 676 1911 680
rect 1915 676 1916 680
rect 1910 675 1916 676
rect 134 672 140 673
rect 110 669 116 670
rect 110 665 111 669
rect 115 665 116 669
rect 134 668 135 672
rect 139 668 140 672
rect 134 667 140 668
rect 174 672 180 673
rect 174 668 175 672
rect 179 668 180 672
rect 174 667 180 668
rect 214 672 220 673
rect 214 668 215 672
rect 219 668 220 672
rect 214 667 220 668
rect 270 672 276 673
rect 270 668 271 672
rect 275 668 276 672
rect 270 667 276 668
rect 334 672 340 673
rect 334 668 335 672
rect 339 668 340 672
rect 334 667 340 668
rect 398 672 404 673
rect 398 668 399 672
rect 403 668 404 672
rect 398 667 404 668
rect 462 672 468 673
rect 462 668 463 672
rect 467 668 468 672
rect 462 667 468 668
rect 526 672 532 673
rect 526 668 527 672
rect 531 668 532 672
rect 526 667 532 668
rect 590 672 596 673
rect 590 668 591 672
rect 595 668 596 672
rect 590 667 596 668
rect 646 672 652 673
rect 646 668 647 672
rect 651 668 652 672
rect 646 667 652 668
rect 702 672 708 673
rect 702 668 703 672
rect 707 668 708 672
rect 702 667 708 668
rect 758 672 764 673
rect 758 668 759 672
rect 763 668 764 672
rect 758 667 764 668
rect 822 672 828 673
rect 822 668 823 672
rect 827 668 828 672
rect 1134 672 1140 673
rect 822 667 828 668
rect 1094 669 1100 670
rect 110 664 116 665
rect 1094 665 1095 669
rect 1099 665 1100 669
rect 1134 668 1135 672
rect 1139 668 1140 672
rect 1134 667 1140 668
rect 1271 667 1277 668
rect 1094 664 1100 665
rect 846 663 852 664
rect 846 662 847 663
rect 673 660 847 662
rect 673 656 675 660
rect 846 659 847 660
rect 851 659 852 663
rect 1271 663 1272 667
rect 1276 666 1277 667
rect 1294 667 1300 668
rect 1294 666 1295 667
rect 1276 664 1295 666
rect 1276 663 1277 664
rect 1271 662 1277 663
rect 1294 663 1295 664
rect 1299 663 1300 667
rect 1294 662 1300 663
rect 1302 667 1308 668
rect 1302 663 1303 667
rect 1307 666 1308 667
rect 1311 667 1317 668
rect 1311 666 1312 667
rect 1307 664 1312 666
rect 1307 663 1308 664
rect 1302 662 1308 663
rect 1311 663 1312 664
rect 1316 663 1317 667
rect 1311 662 1317 663
rect 1350 667 1356 668
rect 1350 663 1351 667
rect 1355 666 1356 667
rect 1359 667 1365 668
rect 1359 666 1360 667
rect 1355 664 1360 666
rect 1355 663 1356 664
rect 1350 662 1356 663
rect 1359 663 1360 664
rect 1364 663 1365 667
rect 1359 662 1365 663
rect 1406 667 1412 668
rect 1406 663 1407 667
rect 1411 666 1412 667
rect 1415 667 1421 668
rect 1415 666 1416 667
rect 1411 664 1416 666
rect 1411 663 1412 664
rect 1406 662 1412 663
rect 1415 663 1416 664
rect 1420 663 1421 667
rect 1415 662 1421 663
rect 1462 667 1468 668
rect 1462 663 1463 667
rect 1467 666 1468 667
rect 1471 667 1477 668
rect 1471 666 1472 667
rect 1467 664 1472 666
rect 1467 663 1468 664
rect 1462 662 1468 663
rect 1471 663 1472 664
rect 1476 663 1477 667
rect 1471 662 1477 663
rect 1526 667 1532 668
rect 1526 663 1527 667
rect 1531 666 1532 667
rect 1535 667 1541 668
rect 1535 666 1536 667
rect 1531 664 1536 666
rect 1531 663 1532 664
rect 1526 662 1532 663
rect 1535 663 1536 664
rect 1540 663 1541 667
rect 1535 662 1541 663
rect 1607 667 1613 668
rect 1607 663 1608 667
rect 1612 666 1613 667
rect 1662 667 1668 668
rect 1662 666 1663 667
rect 1612 664 1663 666
rect 1612 663 1613 664
rect 1607 662 1613 663
rect 1662 663 1663 664
rect 1667 663 1668 667
rect 1662 662 1668 663
rect 1670 667 1676 668
rect 1670 663 1671 667
rect 1675 666 1676 667
rect 1679 667 1685 668
rect 1679 666 1680 667
rect 1675 664 1680 666
rect 1675 663 1676 664
rect 1670 662 1676 663
rect 1679 663 1680 664
rect 1684 663 1685 667
rect 1679 662 1685 663
rect 1718 667 1724 668
rect 1718 663 1719 667
rect 1723 666 1724 667
rect 1759 667 1765 668
rect 1759 666 1760 667
rect 1723 664 1760 666
rect 1723 663 1724 664
rect 1718 662 1724 663
rect 1759 663 1760 664
rect 1764 663 1765 667
rect 1759 662 1765 663
rect 1838 667 1844 668
rect 1838 663 1839 667
rect 1843 666 1844 667
rect 1847 667 1853 668
rect 1847 666 1848 667
rect 1843 664 1848 666
rect 1843 663 1844 664
rect 1838 662 1844 663
rect 1847 663 1848 664
rect 1852 663 1853 667
rect 1847 662 1853 663
rect 1934 667 1941 668
rect 1934 663 1935 667
rect 1940 663 1941 667
rect 1980 666 1982 684
rect 2023 683 2024 684
rect 2028 683 2029 687
rect 2023 682 2029 683
rect 2046 687 2052 688
rect 2046 683 2047 687
rect 2051 686 2052 687
rect 2095 687 2101 688
rect 2095 686 2096 687
rect 2051 684 2096 686
rect 2051 683 2052 684
rect 2046 682 2052 683
rect 2095 683 2096 684
rect 2100 683 2101 687
rect 2095 682 2101 683
rect 1998 680 2004 681
rect 1998 676 1999 680
rect 2003 676 2004 680
rect 1998 675 2004 676
rect 2070 680 2076 681
rect 2070 676 2071 680
rect 2075 676 2076 680
rect 2070 675 2076 676
rect 2118 672 2124 673
rect 2118 668 2119 672
rect 2123 668 2124 672
rect 2023 667 2029 668
rect 2023 666 2024 667
rect 1980 664 2024 666
rect 1934 662 1941 663
rect 2023 663 2024 664
rect 2028 663 2029 667
rect 2023 662 2029 663
rect 2094 667 2101 668
rect 2118 667 2124 668
rect 2094 663 2095 667
rect 2100 663 2101 667
rect 2094 662 2101 663
rect 846 658 852 659
rect 159 655 168 656
rect 110 652 116 653
rect 110 648 111 652
rect 115 648 116 652
rect 159 651 160 655
rect 167 651 168 655
rect 159 650 168 651
rect 182 655 188 656
rect 182 651 183 655
rect 187 654 188 655
rect 199 655 205 656
rect 199 654 200 655
rect 187 652 200 654
rect 187 651 188 652
rect 182 650 188 651
rect 199 651 200 652
rect 204 651 205 655
rect 199 650 205 651
rect 222 655 228 656
rect 222 651 223 655
rect 227 654 228 655
rect 239 655 245 656
rect 239 654 240 655
rect 227 652 240 654
rect 227 651 228 652
rect 222 650 228 651
rect 239 651 240 652
rect 244 651 245 655
rect 239 650 245 651
rect 247 655 253 656
rect 247 651 248 655
rect 252 654 253 655
rect 295 655 301 656
rect 295 654 296 655
rect 252 652 296 654
rect 252 651 253 652
rect 247 650 253 651
rect 295 651 296 652
rect 300 651 301 655
rect 295 650 301 651
rect 359 655 365 656
rect 359 651 360 655
rect 364 654 365 655
rect 418 655 429 656
rect 364 652 414 654
rect 364 651 365 652
rect 359 650 365 651
rect 110 647 116 648
rect 134 644 140 645
rect 134 640 135 644
rect 139 640 140 644
rect 134 639 140 640
rect 174 644 180 645
rect 174 640 175 644
rect 179 640 180 644
rect 174 639 180 640
rect 214 644 220 645
rect 214 640 215 644
rect 219 640 220 644
rect 214 639 220 640
rect 270 644 276 645
rect 270 640 271 644
rect 275 640 276 644
rect 270 639 276 640
rect 334 644 340 645
rect 334 640 335 644
rect 339 640 340 644
rect 334 639 340 640
rect 398 644 404 645
rect 398 640 399 644
rect 403 640 404 644
rect 412 642 414 652
rect 418 651 419 655
rect 423 651 424 655
rect 428 651 429 655
rect 418 650 429 651
rect 431 655 437 656
rect 431 651 432 655
rect 436 654 437 655
rect 487 655 493 656
rect 487 654 488 655
rect 436 652 488 654
rect 436 651 437 652
rect 431 650 437 651
rect 487 651 488 652
rect 492 651 493 655
rect 487 650 493 651
rect 550 655 557 656
rect 550 651 551 655
rect 556 651 557 655
rect 550 650 557 651
rect 559 655 565 656
rect 559 651 560 655
rect 564 654 565 655
rect 615 655 621 656
rect 615 654 616 655
rect 564 652 616 654
rect 564 651 565 652
rect 559 650 565 651
rect 615 651 616 652
rect 620 651 621 655
rect 615 650 621 651
rect 671 655 677 656
rect 671 651 672 655
rect 676 651 677 655
rect 671 650 677 651
rect 726 655 733 656
rect 726 651 727 655
rect 732 651 733 655
rect 726 650 733 651
rect 750 655 756 656
rect 750 651 751 655
rect 755 654 756 655
rect 783 655 789 656
rect 783 654 784 655
rect 755 652 784 654
rect 755 651 756 652
rect 750 650 756 651
rect 783 651 784 652
rect 788 651 789 655
rect 783 650 789 651
rect 791 655 797 656
rect 791 651 792 655
rect 796 654 797 655
rect 847 655 853 656
rect 847 654 848 655
rect 796 652 848 654
rect 796 651 797 652
rect 791 650 797 651
rect 847 651 848 652
rect 852 651 853 655
rect 1134 655 1140 656
rect 847 650 853 651
rect 1094 652 1100 653
rect 1094 648 1095 652
rect 1099 648 1100 652
rect 1134 651 1135 655
rect 1139 651 1140 655
rect 2118 655 2124 656
rect 1134 650 1140 651
rect 1246 652 1252 653
rect 1094 647 1100 648
rect 1246 648 1247 652
rect 1251 648 1252 652
rect 1246 647 1252 648
rect 1286 652 1292 653
rect 1286 648 1287 652
rect 1291 648 1292 652
rect 1286 647 1292 648
rect 1334 652 1340 653
rect 1334 648 1335 652
rect 1339 648 1340 652
rect 1334 647 1340 648
rect 1390 652 1396 653
rect 1390 648 1391 652
rect 1395 648 1396 652
rect 1390 647 1396 648
rect 1446 652 1452 653
rect 1446 648 1447 652
rect 1451 648 1452 652
rect 1446 647 1452 648
rect 1510 652 1516 653
rect 1510 648 1511 652
rect 1515 648 1516 652
rect 1510 647 1516 648
rect 1582 652 1588 653
rect 1582 648 1583 652
rect 1587 648 1588 652
rect 1582 647 1588 648
rect 1654 652 1660 653
rect 1654 648 1655 652
rect 1659 648 1660 652
rect 1654 647 1660 648
rect 1734 652 1740 653
rect 1734 648 1735 652
rect 1739 648 1740 652
rect 1734 647 1740 648
rect 1822 652 1828 653
rect 1822 648 1823 652
rect 1827 648 1828 652
rect 1822 647 1828 648
rect 1910 652 1916 653
rect 1910 648 1911 652
rect 1915 648 1916 652
rect 1910 647 1916 648
rect 1998 652 2004 653
rect 1998 648 1999 652
rect 2003 648 2004 652
rect 1998 647 2004 648
rect 2070 652 2076 653
rect 2070 648 2071 652
rect 2075 648 2076 652
rect 2118 651 2119 655
rect 2123 651 2124 655
rect 2118 650 2124 651
rect 2070 647 2076 648
rect 462 644 468 645
rect 412 640 442 642
rect 398 639 404 640
rect 159 635 165 636
rect 159 631 160 635
rect 164 634 165 635
rect 182 635 188 636
rect 182 634 183 635
rect 164 632 183 634
rect 164 631 165 632
rect 159 630 165 631
rect 182 631 183 632
rect 187 631 188 635
rect 182 630 188 631
rect 199 635 205 636
rect 199 631 200 635
rect 204 634 205 635
rect 222 635 228 636
rect 222 634 223 635
rect 204 632 223 634
rect 204 631 205 632
rect 199 630 205 631
rect 222 631 223 632
rect 227 631 228 635
rect 222 630 228 631
rect 239 635 245 636
rect 239 631 240 635
rect 244 634 245 635
rect 247 635 253 636
rect 247 634 248 635
rect 244 632 248 634
rect 244 631 245 632
rect 239 630 245 631
rect 247 631 248 632
rect 252 631 253 635
rect 247 630 253 631
rect 295 635 304 636
rect 295 631 296 635
rect 303 631 304 635
rect 295 630 304 631
rect 342 635 348 636
rect 342 631 343 635
rect 347 634 348 635
rect 359 635 365 636
rect 359 634 360 635
rect 347 632 360 634
rect 347 631 348 632
rect 342 630 348 631
rect 359 631 360 632
rect 364 631 365 635
rect 359 630 365 631
rect 423 635 429 636
rect 423 631 424 635
rect 428 634 429 635
rect 431 635 437 636
rect 431 634 432 635
rect 428 632 432 634
rect 428 631 429 632
rect 423 630 429 631
rect 431 631 432 632
rect 436 631 437 635
rect 440 634 442 640
rect 462 640 463 644
rect 467 640 468 644
rect 462 639 468 640
rect 526 644 532 645
rect 526 640 527 644
rect 531 640 532 644
rect 526 639 532 640
rect 590 644 596 645
rect 590 640 591 644
rect 595 640 596 644
rect 590 639 596 640
rect 646 644 652 645
rect 646 640 647 644
rect 651 640 652 644
rect 646 639 652 640
rect 702 644 708 645
rect 702 640 703 644
rect 707 640 708 644
rect 702 639 708 640
rect 758 644 764 645
rect 758 640 759 644
rect 763 640 764 644
rect 758 639 764 640
rect 822 644 828 645
rect 822 640 823 644
rect 827 640 828 644
rect 822 639 828 640
rect 1158 640 1164 641
rect 1134 637 1140 638
rect 487 635 493 636
rect 487 634 488 635
rect 440 632 488 634
rect 431 630 437 631
rect 487 631 488 632
rect 492 631 493 635
rect 487 630 493 631
rect 551 635 557 636
rect 551 631 552 635
rect 556 634 557 635
rect 559 635 565 636
rect 559 634 560 635
rect 556 632 560 634
rect 556 631 557 632
rect 551 630 557 631
rect 559 631 560 632
rect 564 631 565 635
rect 559 630 565 631
rect 615 635 621 636
rect 615 631 616 635
rect 620 634 621 635
rect 654 635 660 636
rect 654 634 655 635
rect 620 632 655 634
rect 620 631 621 632
rect 615 630 621 631
rect 654 631 655 632
rect 659 631 660 635
rect 654 630 660 631
rect 671 635 677 636
rect 671 631 672 635
rect 676 631 677 635
rect 671 630 677 631
rect 727 635 733 636
rect 727 631 728 635
rect 732 634 733 635
rect 750 635 756 636
rect 750 634 751 635
rect 732 632 751 634
rect 732 631 733 632
rect 727 630 733 631
rect 750 631 751 632
rect 755 631 756 635
rect 750 630 756 631
rect 783 635 789 636
rect 783 631 784 635
rect 788 634 789 635
rect 791 635 797 636
rect 791 634 792 635
rect 788 632 792 634
rect 788 631 789 632
rect 783 630 789 631
rect 791 631 792 632
rect 796 631 797 635
rect 791 630 797 631
rect 846 635 853 636
rect 846 631 847 635
rect 852 631 853 635
rect 1134 633 1135 637
rect 1139 633 1140 637
rect 1158 636 1159 640
rect 1163 636 1164 640
rect 1158 635 1164 636
rect 1198 640 1204 641
rect 1198 636 1199 640
rect 1203 636 1204 640
rect 1198 635 1204 636
rect 1238 640 1244 641
rect 1238 636 1239 640
rect 1243 636 1244 640
rect 1238 635 1244 636
rect 1278 640 1284 641
rect 1278 636 1279 640
rect 1283 636 1284 640
rect 1278 635 1284 636
rect 1342 640 1348 641
rect 1342 636 1343 640
rect 1347 636 1348 640
rect 1342 635 1348 636
rect 1414 640 1420 641
rect 1414 636 1415 640
rect 1419 636 1420 640
rect 1414 635 1420 636
rect 1494 640 1500 641
rect 1494 636 1495 640
rect 1499 636 1500 640
rect 1494 635 1500 636
rect 1582 640 1588 641
rect 1582 636 1583 640
rect 1587 636 1588 640
rect 1582 635 1588 636
rect 1670 640 1676 641
rect 1670 636 1671 640
rect 1675 636 1676 640
rect 1670 635 1676 636
rect 1758 640 1764 641
rect 1758 636 1759 640
rect 1763 636 1764 640
rect 1758 635 1764 636
rect 1838 640 1844 641
rect 1838 636 1839 640
rect 1843 636 1844 640
rect 1838 635 1844 636
rect 1918 640 1924 641
rect 1918 636 1919 640
rect 1923 636 1924 640
rect 1918 635 1924 636
rect 2006 640 2012 641
rect 2006 636 2007 640
rect 2011 636 2012 640
rect 2006 635 2012 636
rect 2070 640 2076 641
rect 2070 636 2071 640
rect 2075 636 2076 640
rect 2070 635 2076 636
rect 2118 637 2124 638
rect 1134 632 1140 633
rect 2118 633 2119 637
rect 2123 633 2124 637
rect 2118 632 2124 633
rect 846 630 853 631
rect 550 627 556 628
rect 550 623 551 627
rect 555 626 556 627
rect 673 626 675 630
rect 555 624 675 626
rect 555 623 556 624
rect 550 622 556 623
rect 1182 623 1189 624
rect 1134 620 1140 621
rect 1134 616 1135 620
rect 1139 616 1140 620
rect 1182 619 1183 623
rect 1188 619 1189 623
rect 1182 618 1189 619
rect 1206 623 1212 624
rect 1206 619 1207 623
rect 1211 622 1212 623
rect 1223 623 1229 624
rect 1223 622 1224 623
rect 1211 620 1224 622
rect 1211 619 1212 620
rect 1206 618 1212 619
rect 1223 619 1224 620
rect 1228 619 1229 623
rect 1223 618 1229 619
rect 1246 623 1252 624
rect 1246 619 1247 623
rect 1251 622 1252 623
rect 1263 623 1269 624
rect 1263 622 1264 623
rect 1251 620 1264 622
rect 1251 619 1252 620
rect 1246 618 1252 619
rect 1263 619 1264 620
rect 1268 619 1269 623
rect 1263 618 1269 619
rect 1286 623 1292 624
rect 1286 619 1287 623
rect 1291 622 1292 623
rect 1303 623 1309 624
rect 1303 622 1304 623
rect 1291 620 1304 622
rect 1291 619 1292 620
rect 1286 618 1292 619
rect 1303 619 1304 620
rect 1308 619 1309 623
rect 1303 618 1309 619
rect 1311 623 1317 624
rect 1311 619 1312 623
rect 1316 622 1317 623
rect 1367 623 1373 624
rect 1367 622 1368 623
rect 1316 620 1368 622
rect 1316 619 1317 620
rect 1311 618 1317 619
rect 1367 619 1368 620
rect 1372 619 1373 623
rect 1367 618 1373 619
rect 1375 623 1381 624
rect 1375 619 1376 623
rect 1380 622 1381 623
rect 1439 623 1445 624
rect 1439 622 1440 623
rect 1380 620 1440 622
rect 1380 619 1381 620
rect 1375 618 1381 619
rect 1439 619 1440 620
rect 1444 619 1445 623
rect 1439 618 1445 619
rect 1518 623 1525 624
rect 1518 619 1519 623
rect 1524 619 1525 623
rect 1518 618 1525 619
rect 1527 623 1533 624
rect 1527 619 1528 623
rect 1532 622 1533 623
rect 1607 623 1613 624
rect 1607 622 1608 623
rect 1532 620 1608 622
rect 1532 619 1533 620
rect 1527 618 1533 619
rect 1607 619 1608 620
rect 1612 619 1613 623
rect 1607 618 1613 619
rect 1615 623 1621 624
rect 1615 619 1616 623
rect 1620 622 1621 623
rect 1695 623 1701 624
rect 1695 622 1696 623
rect 1620 620 1696 622
rect 1620 619 1621 620
rect 1615 618 1621 619
rect 1695 619 1696 620
rect 1700 619 1701 623
rect 1695 618 1701 619
rect 1703 623 1709 624
rect 1703 619 1704 623
rect 1708 622 1709 623
rect 1783 623 1789 624
rect 1783 622 1784 623
rect 1708 620 1784 622
rect 1708 619 1709 620
rect 1703 618 1709 619
rect 1783 619 1784 620
rect 1788 619 1789 623
rect 1783 618 1789 619
rect 1863 623 1869 624
rect 1863 619 1864 623
rect 1868 622 1869 623
rect 1934 623 1940 624
rect 1934 622 1935 623
rect 1868 620 1935 622
rect 1868 619 1869 620
rect 1863 618 1869 619
rect 1934 619 1935 620
rect 1939 619 1940 623
rect 1934 618 1940 619
rect 1943 623 1952 624
rect 1943 619 1944 623
rect 1951 619 1952 623
rect 1943 618 1952 619
rect 2031 623 2037 624
rect 2031 619 2032 623
rect 2036 622 2037 623
rect 2046 623 2052 624
rect 2046 622 2047 623
rect 2036 620 2047 622
rect 2036 619 2037 620
rect 2031 618 2037 619
rect 2046 619 2047 620
rect 2051 619 2052 623
rect 2046 618 2052 619
rect 2054 623 2060 624
rect 2054 619 2055 623
rect 2059 622 2060 623
rect 2095 623 2101 624
rect 2095 622 2096 623
rect 2059 620 2096 622
rect 2059 619 2060 620
rect 2054 618 2060 619
rect 2095 619 2096 620
rect 2100 619 2101 623
rect 2095 618 2101 619
rect 2118 620 2124 621
rect 162 615 168 616
rect 162 611 163 615
rect 167 614 168 615
rect 610 615 616 616
rect 1134 615 1140 616
rect 2118 616 2119 620
rect 2123 616 2124 620
rect 2118 615 2124 616
rect 167 612 282 614
rect 167 611 168 612
rect 162 610 168 611
rect 280 608 282 612
rect 610 611 611 615
rect 615 614 616 615
rect 615 612 754 614
rect 615 611 616 612
rect 610 610 616 611
rect 752 608 754 612
rect 1158 612 1164 613
rect 1158 608 1159 612
rect 1163 608 1164 612
rect 159 607 165 608
rect 159 603 160 607
rect 164 606 165 607
rect 190 607 196 608
rect 190 606 191 607
rect 164 604 191 606
rect 164 603 165 604
rect 159 602 165 603
rect 190 603 191 604
rect 195 603 196 607
rect 190 602 196 603
rect 199 607 205 608
rect 199 603 200 607
rect 204 606 205 607
rect 230 607 236 608
rect 230 606 231 607
rect 204 604 231 606
rect 204 603 205 604
rect 199 602 205 603
rect 230 603 231 604
rect 235 603 236 607
rect 230 602 236 603
rect 239 607 245 608
rect 239 603 240 607
rect 244 606 245 607
rect 270 607 276 608
rect 270 606 271 607
rect 244 604 271 606
rect 244 603 245 604
rect 239 602 245 603
rect 270 603 271 604
rect 275 603 276 607
rect 270 602 276 603
rect 279 607 285 608
rect 279 603 280 607
rect 284 603 285 607
rect 279 602 285 603
rect 327 607 333 608
rect 327 603 328 607
rect 332 606 333 607
rect 366 607 372 608
rect 366 606 367 607
rect 332 604 367 606
rect 332 603 333 604
rect 327 602 333 603
rect 366 603 367 604
rect 371 603 372 607
rect 366 602 372 603
rect 375 607 381 608
rect 375 603 376 607
rect 380 606 381 607
rect 414 607 420 608
rect 414 606 415 607
rect 380 604 415 606
rect 380 603 381 604
rect 375 602 381 603
rect 414 603 415 604
rect 419 603 420 607
rect 414 602 420 603
rect 423 607 429 608
rect 423 603 424 607
rect 428 606 429 607
rect 446 607 452 608
rect 446 606 447 607
rect 428 604 447 606
rect 428 603 429 604
rect 423 602 429 603
rect 446 603 447 604
rect 451 603 452 607
rect 446 602 452 603
rect 463 607 469 608
rect 463 603 464 607
rect 468 606 469 607
rect 478 607 484 608
rect 478 606 479 607
rect 468 604 479 606
rect 468 603 469 604
rect 463 602 469 603
rect 478 603 479 604
rect 483 603 484 607
rect 478 602 484 603
rect 494 607 500 608
rect 494 603 495 607
rect 499 606 500 607
rect 511 607 517 608
rect 511 606 512 607
rect 499 604 512 606
rect 499 603 500 604
rect 494 602 500 603
rect 511 603 512 604
rect 516 603 517 607
rect 511 602 517 603
rect 526 607 532 608
rect 526 603 527 607
rect 531 606 532 607
rect 559 607 565 608
rect 559 606 560 607
rect 531 604 560 606
rect 531 603 532 604
rect 526 602 532 603
rect 559 603 560 604
rect 564 603 565 607
rect 559 602 565 603
rect 567 607 573 608
rect 567 603 568 607
rect 572 606 573 607
rect 607 607 613 608
rect 607 606 608 607
rect 572 604 608 606
rect 572 603 573 604
rect 567 602 573 603
rect 607 603 608 604
rect 612 603 613 607
rect 607 602 613 603
rect 655 607 661 608
rect 655 603 656 607
rect 660 606 661 607
rect 686 607 692 608
rect 686 606 687 607
rect 660 604 687 606
rect 660 603 661 604
rect 655 602 661 603
rect 686 603 687 604
rect 691 603 692 607
rect 686 602 692 603
rect 703 607 709 608
rect 703 603 704 607
rect 708 606 709 607
rect 742 607 748 608
rect 742 606 743 607
rect 708 604 743 606
rect 708 603 709 604
rect 703 602 709 603
rect 742 603 743 604
rect 747 603 748 607
rect 742 602 748 603
rect 751 607 757 608
rect 1158 607 1164 608
rect 1198 612 1204 613
rect 1198 608 1199 612
rect 1203 608 1204 612
rect 1198 607 1204 608
rect 1238 612 1244 613
rect 1238 608 1239 612
rect 1243 608 1244 612
rect 1238 607 1244 608
rect 1278 612 1284 613
rect 1278 608 1279 612
rect 1283 608 1284 612
rect 1278 607 1284 608
rect 1342 612 1348 613
rect 1342 608 1343 612
rect 1347 608 1348 612
rect 1342 607 1348 608
rect 1414 612 1420 613
rect 1414 608 1415 612
rect 1419 608 1420 612
rect 1414 607 1420 608
rect 1494 612 1500 613
rect 1494 608 1495 612
rect 1499 608 1500 612
rect 1494 607 1500 608
rect 1582 612 1588 613
rect 1582 608 1583 612
rect 1587 608 1588 612
rect 1582 607 1588 608
rect 1670 612 1676 613
rect 1670 608 1671 612
rect 1675 608 1676 612
rect 1670 607 1676 608
rect 1758 612 1764 613
rect 1758 608 1759 612
rect 1763 608 1764 612
rect 1758 607 1764 608
rect 1838 612 1844 613
rect 1838 608 1839 612
rect 1843 608 1844 612
rect 1838 607 1844 608
rect 1918 612 1924 613
rect 1918 608 1919 612
rect 1923 608 1924 612
rect 1918 607 1924 608
rect 2006 612 2012 613
rect 2006 608 2007 612
rect 2011 608 2012 612
rect 2006 607 2012 608
rect 2070 612 2076 613
rect 2070 608 2071 612
rect 2075 608 2076 612
rect 2070 607 2076 608
rect 751 603 752 607
rect 756 603 757 607
rect 751 602 757 603
rect 1183 603 1189 604
rect 134 600 140 601
rect 134 596 135 600
rect 139 596 140 600
rect 134 595 140 596
rect 174 600 180 601
rect 174 596 175 600
rect 179 596 180 600
rect 174 595 180 596
rect 214 600 220 601
rect 214 596 215 600
rect 219 596 220 600
rect 214 595 220 596
rect 254 600 260 601
rect 254 596 255 600
rect 259 596 260 600
rect 254 595 260 596
rect 302 600 308 601
rect 302 596 303 600
rect 307 596 308 600
rect 302 595 308 596
rect 350 600 356 601
rect 350 596 351 600
rect 355 596 356 600
rect 350 595 356 596
rect 398 600 404 601
rect 398 596 399 600
rect 403 596 404 600
rect 398 595 404 596
rect 438 600 444 601
rect 438 596 439 600
rect 443 596 444 600
rect 438 595 444 596
rect 486 600 492 601
rect 486 596 487 600
rect 491 596 492 600
rect 486 595 492 596
rect 534 600 540 601
rect 534 596 535 600
rect 539 596 540 600
rect 534 595 540 596
rect 582 600 588 601
rect 582 596 583 600
rect 587 596 588 600
rect 582 595 588 596
rect 630 600 636 601
rect 630 596 631 600
rect 635 596 636 600
rect 630 595 636 596
rect 678 600 684 601
rect 678 596 679 600
rect 683 596 684 600
rect 678 595 684 596
rect 726 600 732 601
rect 726 596 727 600
rect 731 596 732 600
rect 1183 599 1184 603
rect 1188 602 1189 603
rect 1206 603 1212 604
rect 1206 602 1207 603
rect 1188 600 1207 602
rect 1188 599 1189 600
rect 1183 598 1189 599
rect 1206 599 1207 600
rect 1211 599 1212 603
rect 1206 598 1212 599
rect 1223 603 1229 604
rect 1223 599 1224 603
rect 1228 602 1229 603
rect 1246 603 1252 604
rect 1246 602 1247 603
rect 1228 600 1247 602
rect 1228 599 1229 600
rect 1223 598 1229 599
rect 1246 599 1247 600
rect 1251 599 1252 603
rect 1246 598 1252 599
rect 1263 603 1269 604
rect 1263 599 1264 603
rect 1268 602 1269 603
rect 1286 603 1292 604
rect 1286 602 1287 603
rect 1268 600 1287 602
rect 1268 599 1269 600
rect 1263 598 1269 599
rect 1286 599 1287 600
rect 1291 599 1292 603
rect 1286 598 1292 599
rect 1303 603 1309 604
rect 1303 599 1304 603
rect 1308 602 1309 603
rect 1311 603 1317 604
rect 1311 602 1312 603
rect 1308 600 1312 602
rect 1308 599 1309 600
rect 1303 598 1309 599
rect 1311 599 1312 600
rect 1316 599 1317 603
rect 1311 598 1317 599
rect 1367 603 1373 604
rect 1367 599 1368 603
rect 1372 602 1373 603
rect 1375 603 1381 604
rect 1375 602 1376 603
rect 1372 600 1376 602
rect 1372 599 1373 600
rect 1367 598 1373 599
rect 1375 599 1376 600
rect 1380 599 1381 603
rect 1439 603 1445 604
rect 1439 602 1440 603
rect 1375 598 1381 599
rect 1384 600 1440 602
rect 726 595 732 596
rect 1294 595 1300 596
rect 110 592 116 593
rect 110 588 111 592
rect 115 588 116 592
rect 1094 592 1100 593
rect 1094 588 1095 592
rect 1099 588 1100 592
rect 1294 591 1295 595
rect 1299 594 1300 595
rect 1384 594 1386 600
rect 1439 599 1440 600
rect 1444 599 1445 603
rect 1439 598 1445 599
rect 1519 603 1525 604
rect 1519 599 1520 603
rect 1524 602 1525 603
rect 1527 603 1533 604
rect 1527 602 1528 603
rect 1524 600 1528 602
rect 1524 599 1525 600
rect 1519 598 1525 599
rect 1527 599 1528 600
rect 1532 599 1533 603
rect 1527 598 1533 599
rect 1607 603 1613 604
rect 1607 599 1608 603
rect 1612 602 1613 603
rect 1615 603 1621 604
rect 1615 602 1616 603
rect 1612 600 1616 602
rect 1612 599 1613 600
rect 1607 598 1613 599
rect 1615 599 1616 600
rect 1620 599 1621 603
rect 1615 598 1621 599
rect 1695 603 1701 604
rect 1695 599 1696 603
rect 1700 602 1701 603
rect 1703 603 1709 604
rect 1703 602 1704 603
rect 1700 600 1704 602
rect 1700 599 1701 600
rect 1695 598 1701 599
rect 1703 599 1704 600
rect 1708 599 1709 603
rect 1783 603 1789 604
rect 1783 602 1784 603
rect 1703 598 1709 599
rect 1712 600 1784 602
rect 1299 592 1386 594
rect 1662 595 1668 596
rect 1299 591 1300 592
rect 1294 590 1300 591
rect 1662 591 1663 595
rect 1667 594 1668 595
rect 1712 594 1714 600
rect 1783 599 1784 600
rect 1788 599 1789 603
rect 1783 598 1789 599
rect 1863 603 1869 604
rect 1863 599 1864 603
rect 1868 602 1869 603
rect 1878 603 1884 604
rect 1878 602 1879 603
rect 1868 600 1879 602
rect 1868 599 1869 600
rect 1863 598 1869 599
rect 1878 599 1879 600
rect 1883 599 1884 603
rect 1878 598 1884 599
rect 1934 603 1940 604
rect 1934 599 1935 603
rect 1939 602 1940 603
rect 1943 603 1949 604
rect 1943 602 1944 603
rect 1939 600 1944 602
rect 1939 599 1940 600
rect 1934 598 1940 599
rect 1943 599 1944 600
rect 1948 599 1949 603
rect 1943 598 1949 599
rect 2031 603 2037 604
rect 2031 599 2032 603
rect 2036 602 2037 603
rect 2054 603 2060 604
rect 2054 602 2055 603
rect 2036 600 2055 602
rect 2036 599 2037 600
rect 2031 598 2037 599
rect 2054 599 2055 600
rect 2059 599 2060 603
rect 2054 598 2060 599
rect 2094 603 2101 604
rect 2094 599 2095 603
rect 2100 599 2101 603
rect 2094 598 2101 599
rect 1667 592 1714 594
rect 1667 591 1668 592
rect 1662 590 1668 591
rect 110 587 116 588
rect 158 587 165 588
rect 158 583 159 587
rect 164 583 165 587
rect 158 582 165 583
rect 190 587 196 588
rect 190 583 191 587
rect 195 586 196 587
rect 199 587 205 588
rect 199 586 200 587
rect 195 584 200 586
rect 195 583 196 584
rect 190 582 196 583
rect 199 583 200 584
rect 204 583 205 587
rect 199 582 205 583
rect 230 587 236 588
rect 230 583 231 587
rect 235 586 236 587
rect 239 587 245 588
rect 239 586 240 587
rect 235 584 240 586
rect 235 583 236 584
rect 230 582 236 583
rect 239 583 240 584
rect 244 583 245 587
rect 239 582 245 583
rect 270 587 276 588
rect 270 583 271 587
rect 275 586 276 587
rect 279 587 285 588
rect 279 586 280 587
rect 275 584 280 586
rect 275 583 276 584
rect 270 582 276 583
rect 279 583 280 584
rect 284 583 285 587
rect 279 582 285 583
rect 327 587 333 588
rect 327 583 328 587
rect 332 586 333 587
rect 342 587 348 588
rect 342 586 343 587
rect 332 584 343 586
rect 332 583 333 584
rect 327 582 333 583
rect 342 583 343 584
rect 347 583 348 587
rect 342 582 348 583
rect 366 587 372 588
rect 366 583 367 587
rect 371 586 372 587
rect 375 587 381 588
rect 375 586 376 587
rect 371 584 376 586
rect 371 583 372 584
rect 366 582 372 583
rect 375 583 376 584
rect 380 583 381 587
rect 375 582 381 583
rect 414 587 420 588
rect 414 583 415 587
rect 419 586 420 587
rect 423 587 429 588
rect 423 586 424 587
rect 419 584 424 586
rect 419 583 420 584
rect 414 582 420 583
rect 423 583 424 584
rect 428 583 429 587
rect 423 582 429 583
rect 463 587 469 588
rect 463 583 464 587
rect 468 586 469 587
rect 494 587 500 588
rect 494 586 495 587
rect 468 584 495 586
rect 468 583 469 584
rect 463 582 469 583
rect 494 583 495 584
rect 499 583 500 587
rect 494 582 500 583
rect 511 587 517 588
rect 511 583 512 587
rect 516 586 517 587
rect 526 587 532 588
rect 526 586 527 587
rect 516 584 527 586
rect 516 583 517 584
rect 511 582 517 583
rect 526 583 527 584
rect 531 583 532 587
rect 526 582 532 583
rect 559 587 565 588
rect 559 583 560 587
rect 564 586 565 587
rect 567 587 573 588
rect 567 586 568 587
rect 564 584 568 586
rect 564 583 565 584
rect 559 582 565 583
rect 567 583 568 584
rect 572 583 573 587
rect 567 582 573 583
rect 607 587 616 588
rect 607 583 608 587
rect 615 583 616 587
rect 607 582 616 583
rect 654 587 661 588
rect 654 583 655 587
rect 660 583 661 587
rect 654 582 661 583
rect 686 587 692 588
rect 686 583 687 587
rect 691 586 692 587
rect 703 587 709 588
rect 703 586 704 587
rect 691 584 704 586
rect 691 583 692 584
rect 686 582 692 583
rect 703 583 704 584
rect 708 583 709 587
rect 703 582 709 583
rect 742 587 748 588
rect 742 583 743 587
rect 747 586 748 587
rect 751 587 757 588
rect 1094 587 1100 588
rect 1518 587 1524 588
rect 751 586 752 587
rect 747 584 752 586
rect 747 583 748 584
rect 742 582 748 583
rect 751 583 752 584
rect 756 583 757 587
rect 751 582 757 583
rect 1518 583 1519 587
rect 1523 586 1524 587
rect 1523 584 1778 586
rect 1523 583 1524 584
rect 1518 582 1524 583
rect 1776 580 1778 584
rect 1182 579 1189 580
rect 110 575 116 576
rect 110 571 111 575
rect 115 571 116 575
rect 1094 575 1100 576
rect 110 570 116 571
rect 134 572 140 573
rect 134 568 135 572
rect 139 568 140 572
rect 134 567 140 568
rect 174 572 180 573
rect 174 568 175 572
rect 179 568 180 572
rect 174 567 180 568
rect 214 572 220 573
rect 214 568 215 572
rect 219 568 220 572
rect 214 567 220 568
rect 254 572 260 573
rect 254 568 255 572
rect 259 568 260 572
rect 254 567 260 568
rect 302 572 308 573
rect 302 568 303 572
rect 307 568 308 572
rect 302 567 308 568
rect 350 572 356 573
rect 350 568 351 572
rect 355 568 356 572
rect 350 567 356 568
rect 398 572 404 573
rect 398 568 399 572
rect 403 568 404 572
rect 398 567 404 568
rect 438 572 444 573
rect 438 568 439 572
rect 443 568 444 572
rect 438 567 444 568
rect 486 572 492 573
rect 486 568 487 572
rect 491 568 492 572
rect 486 567 492 568
rect 534 572 540 573
rect 534 568 535 572
rect 539 568 540 572
rect 534 567 540 568
rect 582 572 588 573
rect 582 568 583 572
rect 587 568 588 572
rect 582 567 588 568
rect 630 572 636 573
rect 630 568 631 572
rect 635 568 636 572
rect 630 567 636 568
rect 678 572 684 573
rect 678 568 679 572
rect 683 568 684 572
rect 678 567 684 568
rect 726 572 732 573
rect 726 568 727 572
rect 731 568 732 572
rect 1094 571 1095 575
rect 1099 571 1100 575
rect 1182 575 1183 579
rect 1188 575 1189 579
rect 1182 574 1189 575
rect 1206 579 1212 580
rect 1206 575 1207 579
rect 1211 578 1212 579
rect 1223 579 1229 580
rect 1223 578 1224 579
rect 1211 576 1224 578
rect 1211 575 1212 576
rect 1206 574 1212 575
rect 1223 575 1224 576
rect 1228 575 1229 579
rect 1223 574 1229 575
rect 1246 579 1252 580
rect 1246 575 1247 579
rect 1251 578 1252 579
rect 1263 579 1269 580
rect 1263 578 1264 579
rect 1251 576 1264 578
rect 1251 575 1252 576
rect 1246 574 1252 575
rect 1263 575 1264 576
rect 1268 575 1269 579
rect 1263 574 1269 575
rect 1286 579 1292 580
rect 1286 575 1287 579
rect 1291 578 1292 579
rect 1303 579 1309 580
rect 1303 578 1304 579
rect 1291 576 1304 578
rect 1291 575 1292 576
rect 1286 574 1292 575
rect 1303 575 1304 576
rect 1308 575 1309 579
rect 1303 574 1309 575
rect 1326 579 1332 580
rect 1326 575 1327 579
rect 1331 578 1332 579
rect 1343 579 1349 580
rect 1343 578 1344 579
rect 1331 576 1344 578
rect 1331 575 1332 576
rect 1326 574 1332 575
rect 1343 575 1344 576
rect 1348 575 1349 579
rect 1343 574 1349 575
rect 1366 579 1372 580
rect 1366 575 1367 579
rect 1371 578 1372 579
rect 1383 579 1389 580
rect 1383 578 1384 579
rect 1371 576 1384 578
rect 1371 575 1372 576
rect 1366 574 1372 575
rect 1383 575 1384 576
rect 1388 575 1389 579
rect 1383 574 1389 575
rect 1391 579 1397 580
rect 1391 575 1392 579
rect 1396 578 1397 579
rect 1439 579 1445 580
rect 1439 578 1440 579
rect 1396 576 1440 578
rect 1396 575 1397 576
rect 1391 574 1397 575
rect 1439 575 1440 576
rect 1444 575 1445 579
rect 1439 574 1445 575
rect 1511 579 1517 580
rect 1511 575 1512 579
rect 1516 578 1517 579
rect 1551 579 1557 580
rect 1551 578 1552 579
rect 1516 576 1552 578
rect 1516 575 1517 576
rect 1511 574 1517 575
rect 1551 575 1552 576
rect 1556 575 1557 579
rect 1551 574 1557 575
rect 1591 579 1597 580
rect 1591 575 1592 579
rect 1596 578 1597 579
rect 1670 579 1676 580
rect 1670 578 1671 579
rect 1596 576 1671 578
rect 1596 575 1597 576
rect 1591 574 1597 575
rect 1670 575 1671 576
rect 1675 575 1676 579
rect 1670 574 1676 575
rect 1679 579 1685 580
rect 1679 575 1680 579
rect 1684 578 1685 579
rect 1766 579 1772 580
rect 1766 578 1767 579
rect 1684 576 1767 578
rect 1684 575 1685 576
rect 1679 574 1685 575
rect 1766 575 1767 576
rect 1771 575 1772 579
rect 1766 574 1772 575
rect 1775 579 1781 580
rect 1775 575 1776 579
rect 1780 575 1781 579
rect 1775 574 1781 575
rect 1879 579 1885 580
rect 1879 575 1880 579
rect 1884 578 1885 579
rect 1938 579 1944 580
rect 1938 578 1939 579
rect 1884 576 1939 578
rect 1884 575 1885 576
rect 1879 574 1885 575
rect 1938 575 1939 576
rect 1943 575 1944 579
rect 1938 574 1944 575
rect 1946 579 1952 580
rect 1946 575 1947 579
rect 1951 578 1952 579
rect 1991 579 1997 580
rect 1991 578 1992 579
rect 1951 576 1992 578
rect 1951 575 1952 576
rect 1946 574 1952 575
rect 1991 575 1992 576
rect 1996 575 1997 579
rect 1991 574 1997 575
rect 2046 579 2052 580
rect 2046 575 2047 579
rect 2051 578 2052 579
rect 2095 579 2101 580
rect 2095 578 2096 579
rect 2051 576 2096 578
rect 2051 575 2052 576
rect 2046 574 2052 575
rect 2095 575 2096 576
rect 2100 575 2101 579
rect 2095 574 2101 575
rect 1094 570 1100 571
rect 1158 572 1164 573
rect 726 567 732 568
rect 1158 568 1159 572
rect 1163 568 1164 572
rect 1158 567 1164 568
rect 1198 572 1204 573
rect 1198 568 1199 572
rect 1203 568 1204 572
rect 1198 567 1204 568
rect 1238 572 1244 573
rect 1238 568 1239 572
rect 1243 568 1244 572
rect 1238 567 1244 568
rect 1278 572 1284 573
rect 1278 568 1279 572
rect 1283 568 1284 572
rect 1278 567 1284 568
rect 1318 572 1324 573
rect 1318 568 1319 572
rect 1323 568 1324 572
rect 1318 567 1324 568
rect 1358 572 1364 573
rect 1358 568 1359 572
rect 1363 568 1364 572
rect 1358 567 1364 568
rect 1414 572 1420 573
rect 1414 568 1415 572
rect 1419 568 1420 572
rect 1414 567 1420 568
rect 1486 572 1492 573
rect 1486 568 1487 572
rect 1491 568 1492 572
rect 1486 567 1492 568
rect 1566 572 1572 573
rect 1566 568 1567 572
rect 1571 568 1572 572
rect 1566 567 1572 568
rect 1654 572 1660 573
rect 1654 568 1655 572
rect 1659 568 1660 572
rect 1654 567 1660 568
rect 1750 572 1756 573
rect 1750 568 1751 572
rect 1755 568 1756 572
rect 1750 567 1756 568
rect 1854 572 1860 573
rect 1854 568 1855 572
rect 1859 568 1860 572
rect 1854 567 1860 568
rect 1966 572 1972 573
rect 1966 568 1967 572
rect 1971 568 1972 572
rect 1966 567 1972 568
rect 2070 572 2076 573
rect 2070 568 2071 572
rect 2075 568 2076 572
rect 2070 567 2076 568
rect 1134 564 1140 565
rect 1134 560 1135 564
rect 1139 560 1140 564
rect 2118 564 2124 565
rect 2118 560 2119 564
rect 2123 560 2124 564
rect 1134 559 1140 560
rect 1183 559 1189 560
rect 134 556 140 557
rect 110 553 116 554
rect 110 549 111 553
rect 115 549 116 553
rect 134 552 135 556
rect 139 552 140 556
rect 134 551 140 552
rect 174 556 180 557
rect 174 552 175 556
rect 179 552 180 556
rect 174 551 180 552
rect 222 556 228 557
rect 222 552 223 556
rect 227 552 228 556
rect 222 551 228 552
rect 278 556 284 557
rect 278 552 279 556
rect 283 552 284 556
rect 278 551 284 552
rect 326 556 332 557
rect 326 552 327 556
rect 331 552 332 556
rect 326 551 332 552
rect 374 556 380 557
rect 374 552 375 556
rect 379 552 380 556
rect 374 551 380 552
rect 422 556 428 557
rect 422 552 423 556
rect 427 552 428 556
rect 422 551 428 552
rect 462 556 468 557
rect 462 552 463 556
rect 467 552 468 556
rect 462 551 468 552
rect 510 556 516 557
rect 510 552 511 556
rect 515 552 516 556
rect 510 551 516 552
rect 558 556 564 557
rect 558 552 559 556
rect 563 552 564 556
rect 558 551 564 552
rect 606 556 612 557
rect 606 552 607 556
rect 611 552 612 556
rect 606 551 612 552
rect 654 556 660 557
rect 654 552 655 556
rect 659 552 660 556
rect 654 551 660 552
rect 702 556 708 557
rect 702 552 703 556
rect 707 552 708 556
rect 702 551 708 552
rect 750 556 756 557
rect 750 552 751 556
rect 755 552 756 556
rect 1183 555 1184 559
rect 1188 558 1189 559
rect 1206 559 1212 560
rect 1206 558 1207 559
rect 1188 556 1207 558
rect 1188 555 1189 556
rect 1183 554 1189 555
rect 1206 555 1207 556
rect 1211 555 1212 559
rect 1206 554 1212 555
rect 1223 559 1229 560
rect 1223 555 1224 559
rect 1228 558 1229 559
rect 1246 559 1252 560
rect 1246 558 1247 559
rect 1228 556 1247 558
rect 1228 555 1229 556
rect 1223 554 1229 555
rect 1246 555 1247 556
rect 1251 555 1252 559
rect 1246 554 1252 555
rect 1263 559 1269 560
rect 1263 555 1264 559
rect 1268 558 1269 559
rect 1286 559 1292 560
rect 1286 558 1287 559
rect 1268 556 1287 558
rect 1268 555 1269 556
rect 1263 554 1269 555
rect 1286 555 1287 556
rect 1291 555 1292 559
rect 1286 554 1292 555
rect 1303 559 1309 560
rect 1303 555 1304 559
rect 1308 558 1309 559
rect 1326 559 1332 560
rect 1326 558 1327 559
rect 1308 556 1327 558
rect 1308 555 1309 556
rect 1303 554 1309 555
rect 1326 555 1327 556
rect 1331 555 1332 559
rect 1326 554 1332 555
rect 1343 559 1349 560
rect 1343 555 1344 559
rect 1348 558 1349 559
rect 1366 559 1372 560
rect 1366 558 1367 559
rect 1348 556 1367 558
rect 1348 555 1349 556
rect 1343 554 1349 555
rect 1366 555 1367 556
rect 1371 555 1372 559
rect 1366 554 1372 555
rect 1383 559 1389 560
rect 1383 555 1384 559
rect 1388 558 1389 559
rect 1391 559 1397 560
rect 1391 558 1392 559
rect 1388 556 1392 558
rect 1388 555 1389 556
rect 1383 554 1389 555
rect 1391 555 1392 556
rect 1396 555 1397 559
rect 1391 554 1397 555
rect 1430 559 1436 560
rect 1430 555 1431 559
rect 1435 558 1436 559
rect 1439 559 1445 560
rect 1439 558 1440 559
rect 1435 556 1440 558
rect 1435 555 1436 556
rect 1430 554 1436 555
rect 1439 555 1440 556
rect 1444 555 1445 559
rect 1439 554 1445 555
rect 1511 559 1517 560
rect 1511 555 1512 559
rect 1516 558 1517 559
rect 1534 559 1540 560
rect 1534 558 1535 559
rect 1516 556 1535 558
rect 1516 555 1517 556
rect 1511 554 1517 555
rect 1534 555 1535 556
rect 1539 555 1540 559
rect 1534 554 1540 555
rect 1551 559 1557 560
rect 1551 555 1552 559
rect 1556 558 1557 559
rect 1591 559 1597 560
rect 1591 558 1592 559
rect 1556 556 1592 558
rect 1556 555 1557 556
rect 1551 554 1557 555
rect 1591 555 1592 556
rect 1596 555 1597 559
rect 1591 554 1597 555
rect 1670 559 1676 560
rect 1670 555 1671 559
rect 1675 558 1676 559
rect 1679 559 1685 560
rect 1679 558 1680 559
rect 1675 556 1680 558
rect 1675 555 1676 556
rect 1670 554 1676 555
rect 1679 555 1680 556
rect 1684 555 1685 559
rect 1679 554 1685 555
rect 1766 559 1772 560
rect 1766 555 1767 559
rect 1771 558 1772 559
rect 1775 559 1781 560
rect 1775 558 1776 559
rect 1771 556 1776 558
rect 1771 555 1772 556
rect 1766 554 1772 555
rect 1775 555 1776 556
rect 1780 555 1781 559
rect 1775 554 1781 555
rect 1878 559 1885 560
rect 1878 555 1879 559
rect 1884 555 1885 559
rect 1878 554 1885 555
rect 1938 559 1944 560
rect 1938 555 1939 559
rect 1943 558 1944 559
rect 1991 559 1997 560
rect 1991 558 1992 559
rect 1943 556 1992 558
rect 1943 555 1944 556
rect 1938 554 1944 555
rect 1991 555 1992 556
rect 1996 555 1997 559
rect 1991 554 1997 555
rect 2039 559 2045 560
rect 2039 555 2040 559
rect 2044 558 2045 559
rect 2095 559 2101 560
rect 2118 559 2124 560
rect 2095 558 2096 559
rect 2044 556 2096 558
rect 2044 555 2045 556
rect 2039 554 2045 555
rect 2095 555 2096 556
rect 2100 555 2101 559
rect 2095 554 2101 555
rect 750 551 756 552
rect 1094 553 1100 554
rect 110 548 116 549
rect 1094 549 1095 553
rect 1099 549 1100 553
rect 1094 548 1100 549
rect 1134 547 1140 548
rect 1134 543 1135 547
rect 1139 543 1140 547
rect 2118 547 2124 548
rect 1134 542 1140 543
rect 1158 544 1164 545
rect 1158 540 1159 544
rect 1163 540 1164 544
rect 159 539 165 540
rect 110 536 116 537
rect 110 532 111 536
rect 115 532 116 536
rect 159 535 160 539
rect 164 538 165 539
rect 190 539 196 540
rect 190 538 191 539
rect 164 536 191 538
rect 164 535 165 536
rect 159 534 165 535
rect 190 535 191 536
rect 195 535 196 539
rect 190 534 196 535
rect 199 539 205 540
rect 199 535 200 539
rect 204 538 205 539
rect 238 539 244 540
rect 238 538 239 539
rect 204 536 239 538
rect 204 535 205 536
rect 199 534 205 535
rect 238 535 239 536
rect 243 535 244 539
rect 238 534 244 535
rect 247 539 253 540
rect 247 535 248 539
rect 252 538 253 539
rect 294 539 300 540
rect 294 538 295 539
rect 252 536 295 538
rect 252 535 253 536
rect 247 534 253 535
rect 294 535 295 536
rect 299 535 300 539
rect 294 534 300 535
rect 303 539 309 540
rect 303 535 304 539
rect 308 538 309 539
rect 318 539 324 540
rect 318 538 319 539
rect 308 536 319 538
rect 308 535 309 536
rect 303 534 309 535
rect 318 535 319 536
rect 323 535 324 539
rect 318 534 324 535
rect 351 539 357 540
rect 351 535 352 539
rect 356 538 357 539
rect 390 539 396 540
rect 390 538 391 539
rect 356 536 391 538
rect 356 535 357 536
rect 351 534 357 535
rect 390 535 391 536
rect 395 535 396 539
rect 390 534 396 535
rect 399 539 405 540
rect 399 535 400 539
rect 404 538 405 539
rect 438 539 444 540
rect 438 538 439 539
rect 404 536 439 538
rect 404 535 405 536
rect 399 534 405 535
rect 438 535 439 536
rect 443 535 444 539
rect 438 534 444 535
rect 446 539 453 540
rect 446 535 447 539
rect 452 535 453 539
rect 446 534 453 535
rect 478 539 484 540
rect 478 535 479 539
rect 483 538 484 539
rect 487 539 493 540
rect 487 538 488 539
rect 483 536 488 538
rect 483 535 484 536
rect 478 534 484 535
rect 487 535 488 536
rect 492 535 493 539
rect 487 534 493 535
rect 498 539 504 540
rect 498 535 499 539
rect 503 538 504 539
rect 535 539 541 540
rect 535 538 536 539
rect 503 536 536 538
rect 503 535 504 536
rect 498 534 504 535
rect 535 535 536 536
rect 540 535 541 539
rect 535 534 541 535
rect 543 539 549 540
rect 543 535 544 539
rect 548 538 549 539
rect 583 539 589 540
rect 583 538 584 539
rect 548 536 584 538
rect 548 535 549 536
rect 543 534 549 535
rect 583 535 584 536
rect 588 535 589 539
rect 583 534 589 535
rect 591 539 597 540
rect 591 535 592 539
rect 596 538 597 539
rect 631 539 637 540
rect 631 538 632 539
rect 596 536 632 538
rect 596 535 597 536
rect 591 534 597 535
rect 631 535 632 536
rect 636 535 637 539
rect 631 534 637 535
rect 639 539 645 540
rect 639 535 640 539
rect 644 538 645 539
rect 679 539 685 540
rect 679 538 680 539
rect 644 536 680 538
rect 644 535 645 536
rect 639 534 645 535
rect 679 535 680 536
rect 684 535 685 539
rect 679 534 685 535
rect 690 539 696 540
rect 690 535 691 539
rect 695 538 696 539
rect 727 539 733 540
rect 727 538 728 539
rect 695 536 728 538
rect 695 535 696 536
rect 690 534 696 535
rect 727 535 728 536
rect 732 535 733 539
rect 727 534 733 535
rect 735 539 741 540
rect 735 535 736 539
rect 740 538 741 539
rect 775 539 781 540
rect 1158 539 1164 540
rect 1198 544 1204 545
rect 1198 540 1199 544
rect 1203 540 1204 544
rect 1198 539 1204 540
rect 1238 544 1244 545
rect 1238 540 1239 544
rect 1243 540 1244 544
rect 1238 539 1244 540
rect 1278 544 1284 545
rect 1278 540 1279 544
rect 1283 540 1284 544
rect 1278 539 1284 540
rect 1318 544 1324 545
rect 1318 540 1319 544
rect 1323 540 1324 544
rect 1318 539 1324 540
rect 1358 544 1364 545
rect 1358 540 1359 544
rect 1363 540 1364 544
rect 1358 539 1364 540
rect 1414 544 1420 545
rect 1414 540 1415 544
rect 1419 540 1420 544
rect 1414 539 1420 540
rect 1486 544 1492 545
rect 1486 540 1487 544
rect 1491 540 1492 544
rect 1486 539 1492 540
rect 1566 544 1572 545
rect 1566 540 1567 544
rect 1571 540 1572 544
rect 1566 539 1572 540
rect 1654 544 1660 545
rect 1654 540 1655 544
rect 1659 540 1660 544
rect 1654 539 1660 540
rect 1750 544 1756 545
rect 1750 540 1751 544
rect 1755 540 1756 544
rect 1750 539 1756 540
rect 1854 544 1860 545
rect 1854 540 1855 544
rect 1859 540 1860 544
rect 1854 539 1860 540
rect 1966 544 1972 545
rect 1966 540 1967 544
rect 1971 540 1972 544
rect 1966 539 1972 540
rect 2070 544 2076 545
rect 2070 540 2071 544
rect 2075 540 2076 544
rect 2118 543 2119 547
rect 2123 543 2124 547
rect 2118 542 2124 543
rect 2070 539 2076 540
rect 775 538 776 539
rect 740 536 776 538
rect 740 535 741 536
rect 735 534 741 535
rect 775 535 776 536
rect 780 535 781 539
rect 775 534 781 535
rect 1094 536 1100 537
rect 110 531 116 532
rect 1094 532 1095 536
rect 1099 532 1100 536
rect 1094 531 1100 532
rect 134 528 140 529
rect 134 524 135 528
rect 139 524 140 528
rect 134 523 140 524
rect 174 528 180 529
rect 174 524 175 528
rect 179 524 180 528
rect 174 523 180 524
rect 222 528 228 529
rect 222 524 223 528
rect 227 524 228 528
rect 222 523 228 524
rect 278 528 284 529
rect 278 524 279 528
rect 283 524 284 528
rect 278 523 284 524
rect 326 528 332 529
rect 326 524 327 528
rect 331 524 332 528
rect 326 523 332 524
rect 374 528 380 529
rect 374 524 375 528
rect 379 524 380 528
rect 374 523 380 524
rect 422 528 428 529
rect 422 524 423 528
rect 427 524 428 528
rect 422 523 428 524
rect 462 528 468 529
rect 462 524 463 528
rect 467 524 468 528
rect 462 523 468 524
rect 510 528 516 529
rect 510 524 511 528
rect 515 524 516 528
rect 510 523 516 524
rect 558 528 564 529
rect 558 524 559 528
rect 563 524 564 528
rect 558 523 564 524
rect 606 528 612 529
rect 606 524 607 528
rect 611 524 612 528
rect 606 523 612 524
rect 654 528 660 529
rect 654 524 655 528
rect 659 524 660 528
rect 654 523 660 524
rect 702 528 708 529
rect 702 524 703 528
rect 707 524 708 528
rect 702 523 708 524
rect 750 528 756 529
rect 750 524 751 528
rect 755 524 756 528
rect 1302 528 1308 529
rect 750 523 756 524
rect 1134 525 1140 526
rect 1134 521 1135 525
rect 1139 521 1140 525
rect 1302 524 1303 528
rect 1307 524 1308 528
rect 1302 523 1308 524
rect 1342 528 1348 529
rect 1342 524 1343 528
rect 1347 524 1348 528
rect 1342 523 1348 524
rect 1382 528 1388 529
rect 1382 524 1383 528
rect 1387 524 1388 528
rect 1382 523 1388 524
rect 1422 528 1428 529
rect 1422 524 1423 528
rect 1427 524 1428 528
rect 1422 523 1428 524
rect 1462 528 1468 529
rect 1462 524 1463 528
rect 1467 524 1468 528
rect 1462 523 1468 524
rect 1502 528 1508 529
rect 1502 524 1503 528
rect 1507 524 1508 528
rect 1502 523 1508 524
rect 1542 528 1548 529
rect 1542 524 1543 528
rect 1547 524 1548 528
rect 1542 523 1548 524
rect 1590 528 1596 529
rect 1590 524 1591 528
rect 1595 524 1596 528
rect 1590 523 1596 524
rect 1646 528 1652 529
rect 1646 524 1647 528
rect 1651 524 1652 528
rect 1646 523 1652 524
rect 1702 528 1708 529
rect 1702 524 1703 528
rect 1707 524 1708 528
rect 1702 523 1708 524
rect 1766 528 1772 529
rect 1766 524 1767 528
rect 1771 524 1772 528
rect 1766 523 1772 524
rect 1838 528 1844 529
rect 1838 524 1839 528
rect 1843 524 1844 528
rect 1838 523 1844 524
rect 1918 528 1924 529
rect 1918 524 1919 528
rect 1923 524 1924 528
rect 1918 523 1924 524
rect 2006 528 2012 529
rect 2006 524 2007 528
rect 2011 524 2012 528
rect 2006 523 2012 524
rect 2070 528 2076 529
rect 2070 524 2071 528
rect 2075 524 2076 528
rect 2070 523 2076 524
rect 2118 525 2124 526
rect 1134 520 1140 521
rect 2118 521 2119 525
rect 2123 521 2124 525
rect 2118 520 2124 521
rect 158 519 165 520
rect 158 515 159 519
rect 164 515 165 519
rect 158 514 165 515
rect 190 519 196 520
rect 190 515 191 519
rect 195 518 196 519
rect 199 519 205 520
rect 199 518 200 519
rect 195 516 200 518
rect 195 515 196 516
rect 190 514 196 515
rect 199 515 200 516
rect 204 515 205 519
rect 199 514 205 515
rect 238 519 244 520
rect 238 515 239 519
rect 243 518 244 519
rect 247 519 253 520
rect 247 518 248 519
rect 243 516 248 518
rect 243 515 244 516
rect 238 514 244 515
rect 247 515 248 516
rect 252 515 253 519
rect 247 514 253 515
rect 294 519 300 520
rect 294 515 295 519
rect 299 518 300 519
rect 303 519 309 520
rect 303 518 304 519
rect 299 516 304 518
rect 299 515 300 516
rect 294 514 300 515
rect 303 515 304 516
rect 308 515 309 519
rect 303 514 309 515
rect 351 519 357 520
rect 351 515 352 519
rect 356 518 357 519
rect 382 519 388 520
rect 382 518 383 519
rect 356 516 383 518
rect 356 515 357 516
rect 351 514 357 515
rect 382 515 383 516
rect 387 515 388 519
rect 382 514 388 515
rect 390 519 396 520
rect 390 515 391 519
rect 395 518 396 519
rect 399 519 405 520
rect 399 518 400 519
rect 395 516 400 518
rect 395 515 396 516
rect 390 514 396 515
rect 399 515 400 516
rect 404 515 405 519
rect 399 514 405 515
rect 438 519 444 520
rect 438 515 439 519
rect 443 518 444 519
rect 447 519 453 520
rect 447 518 448 519
rect 443 516 448 518
rect 443 515 444 516
rect 438 514 444 515
rect 447 515 448 516
rect 452 515 453 519
rect 447 514 453 515
rect 487 519 493 520
rect 487 515 488 519
rect 492 518 493 519
rect 498 519 504 520
rect 498 518 499 519
rect 492 516 499 518
rect 492 515 493 516
rect 487 514 493 515
rect 498 515 499 516
rect 503 515 504 519
rect 498 514 504 515
rect 535 519 541 520
rect 535 515 536 519
rect 540 518 541 519
rect 543 519 549 520
rect 543 518 544 519
rect 540 516 544 518
rect 540 515 541 516
rect 535 514 541 515
rect 543 515 544 516
rect 548 515 549 519
rect 543 514 549 515
rect 583 519 589 520
rect 583 515 584 519
rect 588 518 589 519
rect 591 519 597 520
rect 591 518 592 519
rect 588 516 592 518
rect 588 515 589 516
rect 583 514 589 515
rect 591 515 592 516
rect 596 515 597 519
rect 591 514 597 515
rect 631 519 637 520
rect 631 515 632 519
rect 636 518 637 519
rect 639 519 645 520
rect 639 518 640 519
rect 636 516 640 518
rect 636 515 637 516
rect 631 514 637 515
rect 639 515 640 516
rect 644 515 645 519
rect 639 514 645 515
rect 679 519 685 520
rect 679 515 680 519
rect 684 518 685 519
rect 690 519 696 520
rect 690 518 691 519
rect 684 516 691 518
rect 684 515 685 516
rect 679 514 685 515
rect 690 515 691 516
rect 695 515 696 519
rect 690 514 696 515
rect 727 519 733 520
rect 727 515 728 519
rect 732 518 733 519
rect 735 519 741 520
rect 735 518 736 519
rect 732 516 736 518
rect 732 515 733 516
rect 727 514 733 515
rect 735 515 736 516
rect 740 515 741 519
rect 735 514 741 515
rect 775 519 781 520
rect 775 515 776 519
rect 780 515 781 519
rect 1446 519 1452 520
rect 1446 518 1447 519
rect 775 514 781 515
rect 1344 516 1447 518
rect 582 511 588 512
rect 582 507 583 511
rect 587 510 588 511
rect 777 510 779 514
rect 587 508 779 510
rect 1327 511 1333 512
rect 1134 508 1140 509
rect 587 507 588 508
rect 582 506 588 507
rect 1134 504 1135 508
rect 1139 504 1140 508
rect 1327 507 1328 511
rect 1332 510 1333 511
rect 1344 510 1346 516
rect 1446 515 1447 516
rect 1451 515 1452 519
rect 1446 514 1452 515
rect 1332 508 1346 510
rect 1350 511 1356 512
rect 1332 507 1333 508
rect 1327 506 1333 507
rect 1350 507 1351 511
rect 1355 510 1356 511
rect 1367 511 1373 512
rect 1367 510 1368 511
rect 1355 508 1368 510
rect 1355 507 1356 508
rect 1350 506 1356 507
rect 1367 507 1368 508
rect 1372 507 1373 511
rect 1367 506 1373 507
rect 1390 511 1396 512
rect 1390 507 1391 511
rect 1395 510 1396 511
rect 1407 511 1413 512
rect 1407 510 1408 511
rect 1395 508 1408 510
rect 1395 507 1396 508
rect 1390 506 1396 507
rect 1407 507 1408 508
rect 1412 507 1413 511
rect 1407 506 1413 507
rect 1447 511 1453 512
rect 1447 507 1448 511
rect 1452 510 1453 511
rect 1478 511 1484 512
rect 1478 510 1479 511
rect 1452 508 1479 510
rect 1452 507 1453 508
rect 1447 506 1453 507
rect 1478 507 1479 508
rect 1483 507 1484 511
rect 1478 506 1484 507
rect 1487 511 1493 512
rect 1487 507 1488 511
rect 1492 510 1493 511
rect 1518 511 1524 512
rect 1518 510 1519 511
rect 1492 508 1519 510
rect 1492 507 1493 508
rect 1487 506 1493 507
rect 1518 507 1519 508
rect 1523 507 1524 511
rect 1518 506 1524 507
rect 1527 511 1533 512
rect 1527 507 1528 511
rect 1532 510 1533 511
rect 1554 511 1560 512
rect 1532 508 1539 510
rect 1532 507 1533 508
rect 1527 506 1533 507
rect 1134 503 1140 504
rect 1302 500 1308 501
rect 1302 496 1303 500
rect 1307 496 1308 500
rect 1302 495 1308 496
rect 1342 500 1348 501
rect 1342 496 1343 500
rect 1347 496 1348 500
rect 1342 495 1348 496
rect 1382 500 1388 501
rect 1382 496 1383 500
rect 1387 496 1388 500
rect 1382 495 1388 496
rect 1422 500 1428 501
rect 1422 496 1423 500
rect 1427 496 1428 500
rect 1422 495 1428 496
rect 1462 500 1468 501
rect 1462 496 1463 500
rect 1467 496 1468 500
rect 1462 495 1468 496
rect 1502 500 1508 501
rect 1502 496 1503 500
rect 1507 496 1508 500
rect 1502 495 1508 496
rect 159 491 165 492
rect 159 487 160 491
rect 164 490 165 491
rect 190 491 196 492
rect 190 490 191 491
rect 164 488 191 490
rect 164 487 165 488
rect 159 486 165 487
rect 190 487 191 488
rect 195 487 196 491
rect 190 486 196 487
rect 199 491 205 492
rect 199 487 200 491
rect 204 490 205 491
rect 246 491 252 492
rect 246 490 247 491
rect 204 488 247 490
rect 204 487 205 488
rect 199 486 205 487
rect 246 487 247 488
rect 251 487 252 491
rect 246 486 252 487
rect 255 491 261 492
rect 255 487 256 491
rect 260 490 261 491
rect 286 491 292 492
rect 286 490 287 491
rect 260 488 287 490
rect 260 487 261 488
rect 255 486 261 487
rect 286 487 287 488
rect 291 487 292 491
rect 286 486 292 487
rect 318 491 325 492
rect 318 487 319 491
rect 324 487 325 491
rect 318 486 325 487
rect 383 491 389 492
rect 383 487 384 491
rect 388 490 389 491
rect 438 491 444 492
rect 438 490 439 491
rect 388 488 439 490
rect 388 487 389 488
rect 383 486 389 487
rect 438 487 439 488
rect 443 487 444 491
rect 438 486 444 487
rect 447 491 453 492
rect 447 487 448 491
rect 452 490 453 491
rect 494 491 500 492
rect 494 490 495 491
rect 452 488 495 490
rect 452 487 453 488
rect 447 486 453 487
rect 494 487 495 488
rect 499 487 500 491
rect 494 486 500 487
rect 503 491 509 492
rect 503 487 504 491
rect 508 490 509 491
rect 550 491 556 492
rect 550 490 551 491
rect 508 488 551 490
rect 508 487 509 488
rect 503 486 509 487
rect 550 487 551 488
rect 555 487 556 491
rect 550 486 556 487
rect 559 491 565 492
rect 559 487 560 491
rect 564 490 565 491
rect 598 491 604 492
rect 598 490 599 491
rect 564 488 599 490
rect 564 487 565 488
rect 559 486 565 487
rect 598 487 599 488
rect 603 487 604 491
rect 598 486 604 487
rect 615 491 621 492
rect 615 487 616 491
rect 620 490 621 491
rect 654 491 660 492
rect 654 490 655 491
rect 620 488 655 490
rect 620 487 621 488
rect 615 486 621 487
rect 654 487 655 488
rect 659 487 660 491
rect 654 486 660 487
rect 663 491 669 492
rect 663 487 664 491
rect 668 490 669 491
rect 702 491 708 492
rect 702 490 703 491
rect 668 488 703 490
rect 668 487 669 488
rect 663 486 669 487
rect 702 487 703 488
rect 707 487 708 491
rect 702 486 708 487
rect 711 491 717 492
rect 711 487 712 491
rect 716 490 717 491
rect 750 491 756 492
rect 750 490 751 491
rect 716 488 751 490
rect 716 487 717 488
rect 711 486 717 487
rect 750 487 751 488
rect 755 487 756 491
rect 750 486 756 487
rect 759 491 765 492
rect 759 487 760 491
rect 764 490 765 491
rect 806 491 812 492
rect 806 490 807 491
rect 764 488 807 490
rect 764 487 765 488
rect 759 486 765 487
rect 806 487 807 488
rect 811 487 812 491
rect 806 486 812 487
rect 815 491 821 492
rect 815 487 816 491
rect 820 490 821 491
rect 854 491 860 492
rect 854 490 855 491
rect 820 488 855 490
rect 820 487 821 488
rect 815 486 821 487
rect 854 487 855 488
rect 859 487 860 491
rect 854 486 860 487
rect 862 491 868 492
rect 862 487 863 491
rect 867 490 868 491
rect 871 491 877 492
rect 871 490 872 491
rect 867 488 872 490
rect 867 487 868 488
rect 862 486 868 487
rect 871 487 872 488
rect 876 487 877 491
rect 871 486 877 487
rect 1327 491 1333 492
rect 1327 487 1328 491
rect 1332 490 1333 491
rect 1350 491 1356 492
rect 1350 490 1351 491
rect 1332 488 1351 490
rect 1332 487 1333 488
rect 1327 486 1333 487
rect 1350 487 1351 488
rect 1355 487 1356 491
rect 1350 486 1356 487
rect 1367 491 1373 492
rect 1367 487 1368 491
rect 1372 490 1373 491
rect 1390 491 1396 492
rect 1390 490 1391 491
rect 1372 488 1391 490
rect 1372 487 1373 488
rect 1367 486 1373 487
rect 1390 487 1391 488
rect 1395 487 1396 491
rect 1390 486 1396 487
rect 1407 491 1413 492
rect 1407 487 1408 491
rect 1412 490 1413 491
rect 1430 491 1436 492
rect 1430 490 1431 491
rect 1412 488 1431 490
rect 1412 487 1413 488
rect 1407 486 1413 487
rect 1430 487 1431 488
rect 1435 487 1436 491
rect 1430 486 1436 487
rect 1446 491 1453 492
rect 1446 487 1447 491
rect 1452 487 1453 491
rect 1446 486 1453 487
rect 1478 491 1484 492
rect 1478 487 1479 491
rect 1483 490 1484 491
rect 1487 491 1493 492
rect 1487 490 1488 491
rect 1483 488 1488 490
rect 1483 487 1484 488
rect 1478 486 1484 487
rect 1487 487 1488 488
rect 1492 487 1493 491
rect 1487 486 1493 487
rect 1518 491 1524 492
rect 1518 487 1519 491
rect 1523 490 1524 491
rect 1527 491 1533 492
rect 1527 490 1528 491
rect 1523 488 1528 490
rect 1523 487 1524 488
rect 1518 486 1524 487
rect 1527 487 1528 488
rect 1532 487 1533 491
rect 1537 490 1539 508
rect 1554 507 1555 511
rect 1559 510 1560 511
rect 1567 511 1573 512
rect 1567 510 1568 511
rect 1559 508 1568 510
rect 1559 507 1560 508
rect 1554 506 1560 507
rect 1567 507 1568 508
rect 1572 507 1573 511
rect 1567 506 1573 507
rect 1615 511 1621 512
rect 1615 507 1616 511
rect 1620 510 1621 511
rect 1662 511 1668 512
rect 1662 510 1663 511
rect 1620 508 1663 510
rect 1620 507 1621 508
rect 1615 506 1621 507
rect 1662 507 1663 508
rect 1667 507 1668 511
rect 1662 506 1668 507
rect 1671 511 1677 512
rect 1671 507 1672 511
rect 1676 510 1677 511
rect 1718 511 1724 512
rect 1718 510 1719 511
rect 1676 508 1719 510
rect 1676 507 1677 508
rect 1671 506 1677 507
rect 1718 507 1719 508
rect 1723 507 1724 511
rect 1718 506 1724 507
rect 1727 511 1733 512
rect 1727 507 1728 511
rect 1732 510 1733 511
rect 1782 511 1788 512
rect 1782 510 1783 511
rect 1732 508 1783 510
rect 1732 507 1733 508
rect 1727 506 1733 507
rect 1782 507 1783 508
rect 1787 507 1788 511
rect 1782 506 1788 507
rect 1791 511 1797 512
rect 1791 507 1792 511
rect 1796 510 1797 511
rect 1846 511 1852 512
rect 1846 510 1847 511
rect 1796 508 1847 510
rect 1796 507 1797 508
rect 1791 506 1797 507
rect 1846 507 1847 508
rect 1851 507 1852 511
rect 1846 506 1852 507
rect 1863 511 1869 512
rect 1863 507 1864 511
rect 1868 510 1869 511
rect 1910 511 1916 512
rect 1910 510 1911 511
rect 1868 508 1911 510
rect 1868 507 1869 508
rect 1863 506 1869 507
rect 1910 507 1911 508
rect 1915 507 1916 511
rect 1910 506 1916 507
rect 1943 511 1952 512
rect 1943 507 1944 511
rect 1951 507 1952 511
rect 1943 506 1952 507
rect 2031 511 2037 512
rect 2031 507 2032 511
rect 2036 510 2037 511
rect 2078 511 2084 512
rect 2078 510 2079 511
rect 2036 508 2079 510
rect 2036 507 2037 508
rect 2031 506 2037 507
rect 2078 507 2079 508
rect 2083 507 2084 511
rect 2078 506 2084 507
rect 2094 511 2101 512
rect 2094 507 2095 511
rect 2100 507 2101 511
rect 2094 506 2101 507
rect 2118 508 2124 509
rect 2118 504 2119 508
rect 2123 504 2124 508
rect 2118 503 2124 504
rect 1542 500 1548 501
rect 1542 496 1543 500
rect 1547 496 1548 500
rect 1542 495 1548 496
rect 1590 500 1596 501
rect 1590 496 1591 500
rect 1595 496 1596 500
rect 1590 495 1596 496
rect 1646 500 1652 501
rect 1646 496 1647 500
rect 1651 496 1652 500
rect 1646 495 1652 496
rect 1702 500 1708 501
rect 1702 496 1703 500
rect 1707 496 1708 500
rect 1702 495 1708 496
rect 1766 500 1772 501
rect 1766 496 1767 500
rect 1771 496 1772 500
rect 1766 495 1772 496
rect 1838 500 1844 501
rect 1838 496 1839 500
rect 1843 496 1844 500
rect 1838 495 1844 496
rect 1918 500 1924 501
rect 1918 496 1919 500
rect 1923 496 1924 500
rect 1918 495 1924 496
rect 2006 500 2012 501
rect 2006 496 2007 500
rect 2011 496 2012 500
rect 2006 495 2012 496
rect 2070 500 2076 501
rect 2070 496 2071 500
rect 2075 496 2076 500
rect 2070 495 2076 496
rect 1567 491 1573 492
rect 1567 490 1568 491
rect 1537 488 1568 490
rect 1527 486 1533 487
rect 1567 487 1568 488
rect 1572 487 1573 491
rect 1615 491 1621 492
rect 1615 490 1616 491
rect 1567 486 1573 487
rect 1576 488 1616 490
rect 134 484 140 485
rect 134 480 135 484
rect 139 480 140 484
rect 134 479 140 480
rect 174 484 180 485
rect 174 480 175 484
rect 179 480 180 484
rect 174 479 180 480
rect 230 484 236 485
rect 230 480 231 484
rect 235 480 236 484
rect 230 479 236 480
rect 294 484 300 485
rect 294 480 295 484
rect 299 480 300 484
rect 294 479 300 480
rect 358 484 364 485
rect 358 480 359 484
rect 363 480 364 484
rect 358 479 364 480
rect 422 484 428 485
rect 422 480 423 484
rect 427 480 428 484
rect 422 479 428 480
rect 478 484 484 485
rect 478 480 479 484
rect 483 480 484 484
rect 478 479 484 480
rect 534 484 540 485
rect 534 480 535 484
rect 539 480 540 484
rect 534 479 540 480
rect 590 484 596 485
rect 590 480 591 484
rect 595 480 596 484
rect 590 479 596 480
rect 638 484 644 485
rect 638 480 639 484
rect 643 480 644 484
rect 638 479 644 480
rect 686 484 692 485
rect 686 480 687 484
rect 691 480 692 484
rect 686 479 692 480
rect 734 484 740 485
rect 734 480 735 484
rect 739 480 740 484
rect 734 479 740 480
rect 790 484 796 485
rect 790 480 791 484
rect 795 480 796 484
rect 790 479 796 480
rect 846 484 852 485
rect 846 480 847 484
rect 851 480 852 484
rect 846 479 852 480
rect 1534 483 1540 484
rect 1534 479 1535 483
rect 1539 482 1540 483
rect 1576 482 1578 488
rect 1615 487 1616 488
rect 1620 487 1621 491
rect 1615 486 1621 487
rect 1662 491 1668 492
rect 1662 487 1663 491
rect 1667 490 1668 491
rect 1671 491 1677 492
rect 1671 490 1672 491
rect 1667 488 1672 490
rect 1667 487 1668 488
rect 1662 486 1668 487
rect 1671 487 1672 488
rect 1676 487 1677 491
rect 1671 486 1677 487
rect 1718 491 1724 492
rect 1718 487 1719 491
rect 1723 490 1724 491
rect 1727 491 1733 492
rect 1727 490 1728 491
rect 1723 488 1728 490
rect 1723 487 1724 488
rect 1718 486 1724 487
rect 1727 487 1728 488
rect 1732 487 1733 491
rect 1727 486 1733 487
rect 1782 491 1788 492
rect 1782 487 1783 491
rect 1787 490 1788 491
rect 1791 491 1797 492
rect 1791 490 1792 491
rect 1787 488 1792 490
rect 1787 487 1788 488
rect 1782 486 1788 487
rect 1791 487 1792 488
rect 1796 487 1797 491
rect 1791 486 1797 487
rect 1846 491 1852 492
rect 1846 487 1847 491
rect 1851 490 1852 491
rect 1863 491 1869 492
rect 1863 490 1864 491
rect 1851 488 1864 490
rect 1851 487 1852 488
rect 1846 486 1852 487
rect 1863 487 1864 488
rect 1868 487 1869 491
rect 1863 486 1869 487
rect 1943 491 1949 492
rect 1943 487 1944 491
rect 1948 490 1949 491
rect 1998 491 2004 492
rect 1998 490 1999 491
rect 1948 488 1999 490
rect 1948 487 1949 488
rect 1943 486 1949 487
rect 1998 487 1999 488
rect 2003 487 2004 491
rect 1998 486 2004 487
rect 2031 491 2037 492
rect 2031 487 2032 491
rect 2036 490 2037 491
rect 2039 491 2045 492
rect 2039 490 2040 491
rect 2036 488 2040 490
rect 2036 487 2037 488
rect 2031 486 2037 487
rect 2039 487 2040 488
rect 2044 487 2045 491
rect 2039 486 2045 487
rect 2078 491 2084 492
rect 2078 487 2079 491
rect 2083 490 2084 491
rect 2095 491 2101 492
rect 2095 490 2096 491
rect 2083 488 2096 490
rect 2083 487 2084 488
rect 2078 486 2084 487
rect 2095 487 2096 488
rect 2100 487 2101 491
rect 2095 486 2101 487
rect 1539 480 1578 482
rect 1539 479 1540 480
rect 1534 478 1540 479
rect 110 476 116 477
rect 1094 476 1100 477
rect 110 472 111 476
rect 115 472 116 476
rect 582 475 588 476
rect 582 474 583 475
rect 559 473 583 474
rect 110 471 116 472
rect 159 471 165 472
rect 159 467 160 471
rect 164 470 165 471
rect 182 471 188 472
rect 182 470 183 471
rect 164 468 183 470
rect 164 467 165 468
rect 159 466 165 467
rect 182 467 183 468
rect 187 467 188 471
rect 182 466 188 467
rect 190 471 196 472
rect 190 467 191 471
rect 195 470 196 471
rect 199 471 205 472
rect 199 470 200 471
rect 195 468 200 470
rect 195 467 196 468
rect 190 466 196 467
rect 199 467 200 468
rect 204 467 205 471
rect 199 466 205 467
rect 246 471 252 472
rect 246 467 247 471
rect 251 470 252 471
rect 255 471 261 472
rect 255 470 256 471
rect 251 468 256 470
rect 251 467 252 468
rect 246 466 252 467
rect 255 467 256 468
rect 260 467 261 471
rect 255 466 261 467
rect 286 471 292 472
rect 286 467 287 471
rect 291 470 292 471
rect 319 471 325 472
rect 319 470 320 471
rect 291 468 320 470
rect 291 467 292 468
rect 286 466 292 467
rect 319 467 320 468
rect 324 467 325 471
rect 319 466 325 467
rect 382 471 389 472
rect 382 467 383 471
rect 388 467 389 471
rect 382 466 389 467
rect 438 471 444 472
rect 438 467 439 471
rect 443 470 444 471
rect 447 471 453 472
rect 447 470 448 471
rect 443 468 448 470
rect 443 467 444 468
rect 438 466 444 467
rect 447 467 448 468
rect 452 467 453 471
rect 447 466 453 467
rect 494 471 500 472
rect 494 467 495 471
rect 499 470 500 471
rect 503 471 509 472
rect 503 470 504 471
rect 499 468 504 470
rect 499 467 500 468
rect 494 466 500 467
rect 503 467 504 468
rect 508 467 509 471
rect 559 469 560 473
rect 564 472 583 473
rect 564 469 565 472
rect 582 471 583 472
rect 587 471 588 475
rect 1094 472 1095 476
rect 1099 472 1100 476
rect 582 470 588 471
rect 598 471 604 472
rect 559 468 565 469
rect 503 466 509 467
rect 598 467 599 471
rect 603 470 604 471
rect 615 471 621 472
rect 615 470 616 471
rect 603 468 616 470
rect 603 467 604 468
rect 598 466 604 467
rect 615 467 616 468
rect 620 467 621 471
rect 615 466 621 467
rect 654 471 660 472
rect 654 467 655 471
rect 659 470 660 471
rect 663 471 669 472
rect 663 470 664 471
rect 659 468 664 470
rect 659 467 660 468
rect 654 466 660 467
rect 663 467 664 468
rect 668 467 669 471
rect 663 466 669 467
rect 702 471 708 472
rect 702 467 703 471
rect 707 470 708 471
rect 711 471 717 472
rect 711 470 712 471
rect 707 468 712 470
rect 707 467 708 468
rect 702 466 708 467
rect 711 467 712 468
rect 716 467 717 471
rect 711 466 717 467
rect 750 471 756 472
rect 750 467 751 471
rect 755 470 756 471
rect 759 471 765 472
rect 759 470 760 471
rect 755 468 760 470
rect 755 467 756 468
rect 750 466 756 467
rect 759 467 760 468
rect 764 467 765 471
rect 759 466 765 467
rect 806 471 812 472
rect 806 467 807 471
rect 811 470 812 471
rect 815 471 821 472
rect 815 470 816 471
rect 811 468 816 470
rect 811 467 812 468
rect 806 466 812 467
rect 815 467 816 468
rect 820 467 821 471
rect 815 466 821 467
rect 854 471 860 472
rect 854 467 855 471
rect 859 470 860 471
rect 871 471 877 472
rect 1094 471 1100 472
rect 1319 471 1325 472
rect 871 470 872 471
rect 859 468 872 470
rect 859 467 860 468
rect 854 466 860 467
rect 871 467 872 468
rect 876 467 877 471
rect 871 466 877 467
rect 1319 467 1320 471
rect 1324 470 1325 471
rect 1350 471 1356 472
rect 1350 470 1351 471
rect 1324 468 1351 470
rect 1324 467 1325 468
rect 1319 466 1325 467
rect 1350 467 1351 468
rect 1355 467 1356 471
rect 1350 466 1356 467
rect 1359 471 1365 472
rect 1359 467 1360 471
rect 1364 470 1365 471
rect 1390 471 1396 472
rect 1390 470 1391 471
rect 1364 468 1391 470
rect 1364 467 1365 468
rect 1359 466 1365 467
rect 1390 467 1391 468
rect 1395 467 1396 471
rect 1390 466 1396 467
rect 1399 471 1405 472
rect 1399 467 1400 471
rect 1404 470 1405 471
rect 1438 471 1444 472
rect 1438 470 1439 471
rect 1404 468 1439 470
rect 1404 467 1405 468
rect 1399 466 1405 467
rect 1438 467 1439 468
rect 1443 467 1444 471
rect 1438 466 1444 467
rect 1447 471 1453 472
rect 1447 467 1448 471
rect 1452 470 1453 471
rect 1486 471 1492 472
rect 1486 470 1487 471
rect 1452 468 1487 470
rect 1452 467 1453 468
rect 1447 466 1453 467
rect 1486 467 1487 468
rect 1491 467 1492 471
rect 1486 466 1492 467
rect 1495 471 1501 472
rect 1495 467 1496 471
rect 1500 470 1501 471
rect 1542 471 1548 472
rect 1542 470 1543 471
rect 1500 468 1543 470
rect 1500 467 1501 468
rect 1495 466 1501 467
rect 1542 467 1543 468
rect 1547 467 1548 471
rect 1542 466 1548 467
rect 1551 471 1560 472
rect 1551 467 1552 471
rect 1559 467 1560 471
rect 1551 466 1560 467
rect 1607 471 1613 472
rect 1607 467 1608 471
rect 1612 470 1613 471
rect 1662 471 1668 472
rect 1662 470 1663 471
rect 1612 468 1663 470
rect 1612 467 1613 468
rect 1607 466 1613 467
rect 1662 467 1663 468
rect 1667 467 1668 471
rect 1662 466 1668 467
rect 1671 471 1677 472
rect 1671 467 1672 471
rect 1676 470 1677 471
rect 1734 471 1740 472
rect 1734 470 1735 471
rect 1676 468 1735 470
rect 1676 467 1677 468
rect 1671 466 1677 467
rect 1734 467 1735 468
rect 1739 467 1740 471
rect 1734 466 1740 467
rect 1743 471 1749 472
rect 1743 467 1744 471
rect 1748 470 1749 471
rect 1822 471 1828 472
rect 1822 470 1823 471
rect 1748 468 1823 470
rect 1748 467 1749 468
rect 1743 466 1749 467
rect 1822 467 1823 468
rect 1827 467 1828 471
rect 1822 466 1828 467
rect 1831 471 1837 472
rect 1831 467 1832 471
rect 1836 470 1837 471
rect 1902 471 1908 472
rect 1902 470 1903 471
rect 1836 468 1903 470
rect 1836 467 1837 468
rect 1831 466 1837 467
rect 1902 467 1903 468
rect 1907 467 1908 471
rect 1902 466 1908 467
rect 1910 471 1916 472
rect 1910 467 1911 471
rect 1915 470 1916 471
rect 1919 471 1925 472
rect 1919 470 1920 471
rect 1915 468 1920 470
rect 1915 467 1916 468
rect 1910 466 1916 467
rect 1919 467 1920 468
rect 1924 467 1925 471
rect 1919 466 1925 467
rect 2015 471 2024 472
rect 2015 467 2016 471
rect 2023 467 2024 471
rect 2015 466 2024 467
rect 2094 471 2101 472
rect 2094 467 2095 471
rect 2100 467 2101 471
rect 2094 466 2101 467
rect 1294 464 1300 465
rect 1294 460 1295 464
rect 1299 460 1300 464
rect 110 459 116 460
rect 110 455 111 459
rect 115 455 116 459
rect 1094 459 1100 460
rect 1294 459 1300 460
rect 1334 464 1340 465
rect 1334 460 1335 464
rect 1339 460 1340 464
rect 1334 459 1340 460
rect 1374 464 1380 465
rect 1374 460 1375 464
rect 1379 460 1380 464
rect 1374 459 1380 460
rect 1422 464 1428 465
rect 1422 460 1423 464
rect 1427 460 1428 464
rect 1422 459 1428 460
rect 1470 464 1476 465
rect 1470 460 1471 464
rect 1475 460 1476 464
rect 1470 459 1476 460
rect 1526 464 1532 465
rect 1526 460 1527 464
rect 1531 460 1532 464
rect 1526 459 1532 460
rect 1582 464 1588 465
rect 1582 460 1583 464
rect 1587 460 1588 464
rect 1582 459 1588 460
rect 1646 464 1652 465
rect 1646 460 1647 464
rect 1651 460 1652 464
rect 1646 459 1652 460
rect 1718 464 1724 465
rect 1718 460 1719 464
rect 1723 460 1724 464
rect 1718 459 1724 460
rect 1806 464 1812 465
rect 1806 460 1807 464
rect 1811 460 1812 464
rect 1806 459 1812 460
rect 1894 464 1900 465
rect 1894 460 1895 464
rect 1899 460 1900 464
rect 1894 459 1900 460
rect 1990 464 1996 465
rect 1990 460 1991 464
rect 1995 460 1996 464
rect 1990 459 1996 460
rect 2070 464 2076 465
rect 2070 460 2071 464
rect 2075 460 2076 464
rect 2070 459 2076 460
rect 110 454 116 455
rect 134 456 140 457
rect 134 452 135 456
rect 139 452 140 456
rect 134 451 140 452
rect 174 456 180 457
rect 174 452 175 456
rect 179 452 180 456
rect 174 451 180 452
rect 230 456 236 457
rect 230 452 231 456
rect 235 452 236 456
rect 230 451 236 452
rect 294 456 300 457
rect 294 452 295 456
rect 299 452 300 456
rect 294 451 300 452
rect 358 456 364 457
rect 358 452 359 456
rect 363 452 364 456
rect 358 451 364 452
rect 422 456 428 457
rect 422 452 423 456
rect 427 452 428 456
rect 422 451 428 452
rect 478 456 484 457
rect 478 452 479 456
rect 483 452 484 456
rect 478 451 484 452
rect 534 456 540 457
rect 534 452 535 456
rect 539 452 540 456
rect 534 451 540 452
rect 590 456 596 457
rect 590 452 591 456
rect 595 452 596 456
rect 590 451 596 452
rect 638 456 644 457
rect 638 452 639 456
rect 643 452 644 456
rect 638 451 644 452
rect 686 456 692 457
rect 686 452 687 456
rect 691 452 692 456
rect 686 451 692 452
rect 734 456 740 457
rect 734 452 735 456
rect 739 452 740 456
rect 734 451 740 452
rect 790 456 796 457
rect 790 452 791 456
rect 795 452 796 456
rect 790 451 796 452
rect 846 456 852 457
rect 846 452 847 456
rect 851 452 852 456
rect 1094 455 1095 459
rect 1099 455 1100 459
rect 1094 454 1100 455
rect 1134 456 1140 457
rect 846 451 852 452
rect 1134 452 1135 456
rect 1139 452 1140 456
rect 2118 456 2124 457
rect 2118 452 2119 456
rect 2123 452 2124 456
rect 1134 451 1140 452
rect 1319 451 1325 452
rect 1319 447 1320 451
rect 1324 450 1325 451
rect 1342 451 1348 452
rect 1342 450 1343 451
rect 1324 448 1343 450
rect 1324 447 1325 448
rect 1319 446 1325 447
rect 1342 447 1343 448
rect 1347 447 1348 451
rect 1342 446 1348 447
rect 1350 451 1356 452
rect 1350 447 1351 451
rect 1355 450 1356 451
rect 1359 451 1365 452
rect 1359 450 1360 451
rect 1355 448 1360 450
rect 1355 447 1356 448
rect 1350 446 1356 447
rect 1359 447 1360 448
rect 1364 447 1365 451
rect 1359 446 1365 447
rect 1390 451 1396 452
rect 1390 447 1391 451
rect 1395 450 1396 451
rect 1399 451 1405 452
rect 1399 450 1400 451
rect 1395 448 1400 450
rect 1395 447 1396 448
rect 1390 446 1396 447
rect 1399 447 1400 448
rect 1404 447 1405 451
rect 1399 446 1405 447
rect 1438 451 1444 452
rect 1438 447 1439 451
rect 1443 450 1444 451
rect 1447 451 1453 452
rect 1447 450 1448 451
rect 1443 448 1448 450
rect 1443 447 1444 448
rect 1438 446 1444 447
rect 1447 447 1448 448
rect 1452 447 1453 451
rect 1447 446 1453 447
rect 1486 451 1492 452
rect 1486 447 1487 451
rect 1491 450 1492 451
rect 1495 451 1501 452
rect 1495 450 1496 451
rect 1491 448 1496 450
rect 1491 447 1492 448
rect 1486 446 1492 447
rect 1495 447 1496 448
rect 1500 447 1501 451
rect 1495 446 1501 447
rect 1542 451 1548 452
rect 1542 447 1543 451
rect 1547 450 1548 451
rect 1551 451 1557 452
rect 1551 450 1552 451
rect 1547 448 1552 450
rect 1547 447 1548 448
rect 1542 446 1548 447
rect 1551 447 1552 448
rect 1556 447 1557 451
rect 1551 446 1557 447
rect 1607 451 1616 452
rect 1607 447 1608 451
rect 1615 447 1616 451
rect 1607 446 1616 447
rect 1662 451 1668 452
rect 1662 447 1663 451
rect 1667 450 1668 451
rect 1671 451 1677 452
rect 1671 450 1672 451
rect 1667 448 1672 450
rect 1667 447 1668 448
rect 1662 446 1668 447
rect 1671 447 1672 448
rect 1676 447 1677 451
rect 1671 446 1677 447
rect 1734 451 1740 452
rect 1734 447 1735 451
rect 1739 450 1740 451
rect 1743 451 1749 452
rect 1743 450 1744 451
rect 1739 448 1744 450
rect 1739 447 1740 448
rect 1734 446 1740 447
rect 1743 447 1744 448
rect 1748 447 1749 451
rect 1743 446 1749 447
rect 1822 451 1828 452
rect 1822 447 1823 451
rect 1827 450 1828 451
rect 1831 451 1837 452
rect 1831 450 1832 451
rect 1827 448 1832 450
rect 1827 447 1828 448
rect 1822 446 1828 447
rect 1831 447 1832 448
rect 1836 447 1837 451
rect 1831 446 1837 447
rect 1902 451 1908 452
rect 1902 447 1903 451
rect 1907 450 1908 451
rect 1919 451 1925 452
rect 1919 450 1920 451
rect 1907 448 1920 450
rect 1907 447 1908 448
rect 1902 446 1908 447
rect 1919 447 1920 448
rect 1924 447 1925 451
rect 1919 446 1925 447
rect 1998 451 2004 452
rect 1998 447 1999 451
rect 2003 450 2004 451
rect 2015 451 2021 452
rect 2015 450 2016 451
rect 2003 448 2016 450
rect 2003 447 2004 448
rect 1998 446 2004 447
rect 2015 447 2016 448
rect 2020 447 2021 451
rect 2015 446 2021 447
rect 2094 451 2101 452
rect 2118 451 2124 452
rect 2094 447 2095 451
rect 2100 447 2101 451
rect 2094 446 2101 447
rect 174 440 180 441
rect 110 437 116 438
rect 110 433 111 437
rect 115 433 116 437
rect 174 436 175 440
rect 179 436 180 440
rect 174 435 180 436
rect 214 440 220 441
rect 214 436 215 440
rect 219 436 220 440
rect 214 435 220 436
rect 262 440 268 441
rect 262 436 263 440
rect 267 436 268 440
rect 262 435 268 436
rect 326 440 332 441
rect 326 436 327 440
rect 331 436 332 440
rect 326 435 332 436
rect 390 440 396 441
rect 390 436 391 440
rect 395 436 396 440
rect 390 435 396 436
rect 462 440 468 441
rect 462 436 463 440
rect 467 436 468 440
rect 462 435 468 436
rect 534 440 540 441
rect 534 436 535 440
rect 539 436 540 440
rect 534 435 540 436
rect 606 440 612 441
rect 606 436 607 440
rect 611 436 612 440
rect 606 435 612 436
rect 678 440 684 441
rect 678 436 679 440
rect 683 436 684 440
rect 678 435 684 436
rect 742 440 748 441
rect 742 436 743 440
rect 747 436 748 440
rect 742 435 748 436
rect 806 440 812 441
rect 806 436 807 440
rect 811 436 812 440
rect 806 435 812 436
rect 870 440 876 441
rect 870 436 871 440
rect 875 436 876 440
rect 870 435 876 436
rect 942 440 948 441
rect 942 436 943 440
rect 947 436 948 440
rect 1134 439 1140 440
rect 942 435 948 436
rect 1094 437 1100 438
rect 110 432 116 433
rect 1094 433 1095 437
rect 1099 433 1100 437
rect 1134 435 1135 439
rect 1139 435 1140 439
rect 2118 439 2124 440
rect 1134 434 1140 435
rect 1294 436 1300 437
rect 1094 432 1100 433
rect 1294 432 1295 436
rect 1299 432 1300 436
rect 862 431 868 432
rect 1294 431 1300 432
rect 1334 436 1340 437
rect 1334 432 1335 436
rect 1339 432 1340 436
rect 1334 431 1340 432
rect 1374 436 1380 437
rect 1374 432 1375 436
rect 1379 432 1380 436
rect 1374 431 1380 432
rect 1422 436 1428 437
rect 1422 432 1423 436
rect 1427 432 1428 436
rect 1422 431 1428 432
rect 1470 436 1476 437
rect 1470 432 1471 436
rect 1475 432 1476 436
rect 1470 431 1476 432
rect 1526 436 1532 437
rect 1526 432 1527 436
rect 1531 432 1532 436
rect 1526 431 1532 432
rect 1582 436 1588 437
rect 1582 432 1583 436
rect 1587 432 1588 436
rect 1582 431 1588 432
rect 1646 436 1652 437
rect 1646 432 1647 436
rect 1651 432 1652 436
rect 1646 431 1652 432
rect 1718 436 1724 437
rect 1718 432 1719 436
rect 1723 432 1724 436
rect 1718 431 1724 432
rect 1806 436 1812 437
rect 1806 432 1807 436
rect 1811 432 1812 436
rect 1806 431 1812 432
rect 1894 436 1900 437
rect 1894 432 1895 436
rect 1899 432 1900 436
rect 1894 431 1900 432
rect 1990 436 1996 437
rect 1990 432 1991 436
rect 1995 432 1996 436
rect 1990 431 1996 432
rect 2070 436 2076 437
rect 2070 432 2071 436
rect 2075 432 2076 436
rect 2118 435 2119 439
rect 2123 435 2124 439
rect 2118 434 2124 435
rect 2070 431 2076 432
rect 862 430 863 431
rect 633 428 863 430
rect 633 424 635 428
rect 862 427 863 428
rect 867 427 868 431
rect 862 426 868 427
rect 1158 424 1164 425
rect 198 423 205 424
rect 110 420 116 421
rect 110 416 111 420
rect 115 416 116 420
rect 198 419 199 423
rect 204 419 205 423
rect 198 418 205 419
rect 222 423 228 424
rect 222 419 223 423
rect 227 422 228 423
rect 239 423 245 424
rect 239 422 240 423
rect 227 420 240 422
rect 227 419 228 420
rect 222 418 228 419
rect 239 419 240 420
rect 244 419 245 423
rect 239 418 245 419
rect 250 423 256 424
rect 250 419 251 423
rect 255 422 256 423
rect 287 423 293 424
rect 287 422 288 423
rect 255 420 288 422
rect 255 419 256 420
rect 250 418 256 419
rect 287 419 288 420
rect 292 419 293 423
rect 287 418 293 419
rect 350 423 357 424
rect 350 419 351 423
rect 356 419 357 423
rect 350 418 357 419
rect 359 423 365 424
rect 359 419 360 423
rect 364 422 365 423
rect 415 423 421 424
rect 415 422 416 423
rect 364 420 416 422
rect 364 419 365 420
rect 359 418 365 419
rect 415 419 416 420
rect 420 419 421 423
rect 415 418 421 419
rect 487 423 493 424
rect 487 419 488 423
rect 492 422 493 423
rect 550 423 556 424
rect 550 422 551 423
rect 492 420 551 422
rect 492 419 493 420
rect 487 418 493 419
rect 550 419 551 420
rect 555 419 556 423
rect 550 418 556 419
rect 558 423 565 424
rect 558 419 559 423
rect 564 419 565 423
rect 558 418 565 419
rect 631 423 637 424
rect 631 419 632 423
rect 636 419 637 423
rect 631 418 637 419
rect 639 423 645 424
rect 639 419 640 423
rect 644 422 645 423
rect 703 423 709 424
rect 703 422 704 423
rect 644 420 704 422
rect 644 419 645 420
rect 639 418 645 419
rect 703 419 704 420
rect 708 419 709 423
rect 703 418 709 419
rect 711 423 717 424
rect 711 419 712 423
rect 716 422 717 423
rect 767 423 773 424
rect 767 422 768 423
rect 716 420 768 422
rect 716 419 717 420
rect 711 418 717 419
rect 767 419 768 420
rect 772 419 773 423
rect 767 418 773 419
rect 775 423 781 424
rect 775 419 776 423
rect 780 422 781 423
rect 831 423 837 424
rect 831 422 832 423
rect 780 420 832 422
rect 780 419 781 420
rect 775 418 781 419
rect 831 419 832 420
rect 836 419 837 423
rect 831 418 837 419
rect 839 423 845 424
rect 839 419 840 423
rect 844 422 845 423
rect 895 423 901 424
rect 895 422 896 423
rect 844 420 896 422
rect 844 419 845 420
rect 839 418 845 419
rect 895 419 896 420
rect 900 419 901 423
rect 895 418 901 419
rect 903 423 909 424
rect 903 419 904 423
rect 908 422 909 423
rect 967 423 973 424
rect 967 422 968 423
rect 908 420 968 422
rect 908 419 909 420
rect 903 418 909 419
rect 967 419 968 420
rect 972 419 973 423
rect 1134 421 1140 422
rect 967 418 973 419
rect 1094 420 1100 421
rect 110 415 116 416
rect 1094 416 1095 420
rect 1099 416 1100 420
rect 1134 417 1135 421
rect 1139 417 1140 421
rect 1158 420 1159 424
rect 1163 420 1164 424
rect 1158 419 1164 420
rect 1198 424 1204 425
rect 1198 420 1199 424
rect 1203 420 1204 424
rect 1198 419 1204 420
rect 1254 424 1260 425
rect 1254 420 1255 424
rect 1259 420 1260 424
rect 1254 419 1260 420
rect 1334 424 1340 425
rect 1334 420 1335 424
rect 1339 420 1340 424
rect 1334 419 1340 420
rect 1414 424 1420 425
rect 1414 420 1415 424
rect 1419 420 1420 424
rect 1414 419 1420 420
rect 1502 424 1508 425
rect 1502 420 1503 424
rect 1507 420 1508 424
rect 1502 419 1508 420
rect 1590 424 1596 425
rect 1590 420 1591 424
rect 1595 420 1596 424
rect 1590 419 1596 420
rect 1670 424 1676 425
rect 1670 420 1671 424
rect 1675 420 1676 424
rect 1670 419 1676 420
rect 1750 424 1756 425
rect 1750 420 1751 424
rect 1755 420 1756 424
rect 1750 419 1756 420
rect 1830 424 1836 425
rect 1830 420 1831 424
rect 1835 420 1836 424
rect 1830 419 1836 420
rect 1910 424 1916 425
rect 1910 420 1911 424
rect 1915 420 1916 424
rect 1910 419 1916 420
rect 1998 424 2004 425
rect 1998 420 1999 424
rect 2003 420 2004 424
rect 1998 419 2004 420
rect 2070 424 2076 425
rect 2070 420 2071 424
rect 2075 420 2076 424
rect 2070 419 2076 420
rect 2118 421 2124 422
rect 1134 416 1140 417
rect 2118 417 2119 421
rect 2123 417 2124 421
rect 2118 416 2124 417
rect 1094 415 1100 416
rect 1486 415 1492 416
rect 1486 414 1487 415
rect 174 412 180 413
rect 174 408 175 412
rect 179 408 180 412
rect 174 407 180 408
rect 214 412 220 413
rect 214 408 215 412
rect 219 408 220 412
rect 214 407 220 408
rect 262 412 268 413
rect 262 408 263 412
rect 267 408 268 412
rect 262 407 268 408
rect 326 412 332 413
rect 326 408 327 412
rect 331 408 332 412
rect 326 407 332 408
rect 390 412 396 413
rect 390 408 391 412
rect 395 408 396 412
rect 390 407 396 408
rect 462 412 468 413
rect 462 408 463 412
rect 467 408 468 412
rect 462 407 468 408
rect 534 412 540 413
rect 534 408 535 412
rect 539 408 540 412
rect 534 407 540 408
rect 606 412 612 413
rect 606 408 607 412
rect 611 408 612 412
rect 606 407 612 408
rect 678 412 684 413
rect 678 408 679 412
rect 683 408 684 412
rect 678 407 684 408
rect 742 412 748 413
rect 742 408 743 412
rect 747 408 748 412
rect 742 407 748 408
rect 806 412 812 413
rect 806 408 807 412
rect 811 408 812 412
rect 806 407 812 408
rect 870 412 876 413
rect 870 408 871 412
rect 875 408 876 412
rect 870 407 876 408
rect 942 412 948 413
rect 942 408 943 412
rect 947 408 948 412
rect 1184 412 1487 414
rect 1184 410 1186 412
rect 1486 411 1487 412
rect 1491 411 1492 415
rect 1854 415 1860 416
rect 1854 414 1855 415
rect 1486 410 1492 411
rect 1681 412 1855 414
rect 942 407 948 408
rect 1183 409 1189 410
rect 1183 405 1184 409
rect 1188 405 1189 409
rect 1134 404 1140 405
rect 1183 404 1189 405
rect 1206 407 1212 408
rect 199 403 205 404
rect 199 399 200 403
rect 204 402 205 403
rect 222 403 228 404
rect 222 402 223 403
rect 204 400 223 402
rect 204 399 205 400
rect 199 398 205 399
rect 222 399 223 400
rect 227 399 228 403
rect 222 398 228 399
rect 239 403 245 404
rect 239 399 240 403
rect 244 402 245 403
rect 250 403 256 404
rect 250 402 251 403
rect 244 400 251 402
rect 244 399 245 400
rect 239 398 245 399
rect 250 399 251 400
rect 255 399 256 403
rect 287 403 293 404
rect 287 402 288 403
rect 250 398 256 399
rect 260 400 288 402
rect 182 395 188 396
rect 182 391 183 395
rect 187 394 188 395
rect 260 394 262 400
rect 287 399 288 400
rect 292 399 293 403
rect 287 398 293 399
rect 351 403 357 404
rect 351 399 352 403
rect 356 402 357 403
rect 359 403 365 404
rect 359 402 360 403
rect 356 400 360 402
rect 356 399 357 400
rect 351 398 357 399
rect 359 399 360 400
rect 364 399 365 403
rect 359 398 365 399
rect 415 403 421 404
rect 415 399 416 403
rect 420 402 421 403
rect 430 403 436 404
rect 430 402 431 403
rect 420 400 431 402
rect 420 399 421 400
rect 415 398 421 399
rect 430 399 431 400
rect 435 399 436 403
rect 430 398 436 399
rect 487 403 493 404
rect 487 399 488 403
rect 492 399 493 403
rect 487 398 493 399
rect 550 403 556 404
rect 550 399 551 403
rect 555 402 556 403
rect 559 403 565 404
rect 559 402 560 403
rect 555 400 560 402
rect 555 399 556 400
rect 550 398 556 399
rect 559 399 560 400
rect 564 399 565 403
rect 559 398 565 399
rect 631 403 637 404
rect 631 399 632 403
rect 636 402 637 403
rect 639 403 645 404
rect 639 402 640 403
rect 636 400 640 402
rect 636 399 637 400
rect 631 398 637 399
rect 639 399 640 400
rect 644 399 645 403
rect 639 398 645 399
rect 703 403 709 404
rect 703 399 704 403
rect 708 402 709 403
rect 711 403 717 404
rect 711 402 712 403
rect 708 400 712 402
rect 708 399 709 400
rect 703 398 709 399
rect 711 399 712 400
rect 716 399 717 403
rect 711 398 717 399
rect 767 403 773 404
rect 767 399 768 403
rect 772 402 773 403
rect 775 403 781 404
rect 775 402 776 403
rect 772 400 776 402
rect 772 399 773 400
rect 767 398 773 399
rect 775 399 776 400
rect 780 399 781 403
rect 775 398 781 399
rect 831 403 837 404
rect 831 399 832 403
rect 836 402 837 403
rect 839 403 845 404
rect 839 402 840 403
rect 836 400 840 402
rect 836 399 837 400
rect 831 398 837 399
rect 839 399 840 400
rect 844 399 845 403
rect 839 398 845 399
rect 895 403 901 404
rect 895 399 896 403
rect 900 402 901 403
rect 903 403 909 404
rect 903 402 904 403
rect 900 400 904 402
rect 900 399 901 400
rect 895 398 901 399
rect 903 399 904 400
rect 908 399 909 403
rect 903 398 909 399
rect 914 403 920 404
rect 914 399 915 403
rect 919 402 920 403
rect 967 403 973 404
rect 967 402 968 403
rect 919 400 968 402
rect 919 399 920 400
rect 914 398 920 399
rect 967 399 968 400
rect 972 399 973 403
rect 1134 400 1135 404
rect 1139 400 1140 404
rect 1206 403 1207 407
rect 1211 406 1212 407
rect 1223 407 1229 408
rect 1223 406 1224 407
rect 1211 404 1224 406
rect 1211 403 1212 404
rect 1206 402 1212 403
rect 1223 403 1224 404
rect 1228 403 1229 407
rect 1223 402 1229 403
rect 1231 407 1237 408
rect 1231 403 1232 407
rect 1236 406 1237 407
rect 1279 407 1285 408
rect 1279 406 1280 407
rect 1236 404 1280 406
rect 1236 403 1237 404
rect 1231 402 1237 403
rect 1279 403 1280 404
rect 1284 403 1285 407
rect 1279 402 1285 403
rect 1287 407 1293 408
rect 1287 403 1288 407
rect 1292 406 1293 407
rect 1359 407 1365 408
rect 1359 406 1360 407
rect 1292 404 1360 406
rect 1292 403 1293 404
rect 1287 402 1293 403
rect 1359 403 1360 404
rect 1364 403 1365 407
rect 1359 402 1365 403
rect 1367 407 1373 408
rect 1367 403 1368 407
rect 1372 406 1373 407
rect 1439 407 1445 408
rect 1439 406 1440 407
rect 1372 404 1440 406
rect 1372 403 1373 404
rect 1367 402 1373 403
rect 1439 403 1440 404
rect 1444 403 1445 407
rect 1439 402 1445 403
rect 1447 407 1453 408
rect 1447 403 1448 407
rect 1452 406 1453 407
rect 1527 407 1533 408
rect 1527 406 1528 407
rect 1452 404 1528 406
rect 1452 403 1453 404
rect 1447 402 1453 403
rect 1527 403 1528 404
rect 1532 403 1533 407
rect 1527 402 1533 403
rect 1615 407 1621 408
rect 1615 403 1616 407
rect 1620 406 1621 407
rect 1681 406 1683 412
rect 1854 411 1855 412
rect 1859 411 1860 415
rect 1854 410 1860 411
rect 1620 404 1683 406
rect 1686 407 1692 408
rect 1620 403 1621 404
rect 1615 402 1621 403
rect 1686 403 1687 407
rect 1691 406 1692 407
rect 1695 407 1701 408
rect 1695 406 1696 407
rect 1691 404 1696 406
rect 1691 403 1692 404
rect 1686 402 1692 403
rect 1695 403 1696 404
rect 1700 403 1701 407
rect 1695 402 1701 403
rect 1706 407 1712 408
rect 1706 403 1707 407
rect 1711 406 1712 407
rect 1775 407 1781 408
rect 1775 406 1776 407
rect 1711 404 1776 406
rect 1711 403 1712 404
rect 1706 402 1712 403
rect 1775 403 1776 404
rect 1780 403 1781 407
rect 1775 402 1781 403
rect 1783 407 1789 408
rect 1783 403 1784 407
rect 1788 406 1789 407
rect 1855 407 1861 408
rect 1855 406 1856 407
rect 1788 404 1856 406
rect 1788 403 1789 404
rect 1783 402 1789 403
rect 1855 403 1856 404
rect 1860 403 1861 407
rect 1855 402 1861 403
rect 1935 407 1941 408
rect 1935 403 1936 407
rect 1940 406 1941 407
rect 2010 407 2016 408
rect 2010 406 2011 407
rect 1940 404 2011 406
rect 1940 403 1941 404
rect 1935 402 1941 403
rect 2010 403 2011 404
rect 2015 403 2016 407
rect 2010 402 2016 403
rect 2018 407 2029 408
rect 2018 403 2019 407
rect 2023 403 2024 407
rect 2028 403 2029 407
rect 2018 402 2029 403
rect 2095 407 2101 408
rect 2095 403 2096 407
rect 2100 406 2101 407
rect 2103 407 2109 408
rect 2103 406 2104 407
rect 2100 404 2104 406
rect 2100 403 2101 404
rect 2095 402 2101 403
rect 2103 403 2104 404
rect 2108 403 2109 407
rect 2103 402 2109 403
rect 2118 404 2124 405
rect 1134 399 1140 400
rect 2118 400 2119 404
rect 2123 400 2124 404
rect 2118 399 2124 400
rect 967 398 973 399
rect 187 392 262 394
rect 350 395 356 396
rect 187 391 188 392
rect 182 390 188 391
rect 350 391 351 395
rect 355 394 356 395
rect 489 394 491 398
rect 355 392 491 394
rect 1158 396 1164 397
rect 1158 392 1159 396
rect 1163 392 1164 396
rect 355 391 356 392
rect 1158 391 1164 392
rect 1198 396 1204 397
rect 1198 392 1199 396
rect 1203 392 1204 396
rect 1198 391 1204 392
rect 1254 396 1260 397
rect 1254 392 1255 396
rect 1259 392 1260 396
rect 1254 391 1260 392
rect 1334 396 1340 397
rect 1334 392 1335 396
rect 1339 392 1340 396
rect 1334 391 1340 392
rect 1414 396 1420 397
rect 1414 392 1415 396
rect 1419 392 1420 396
rect 1414 391 1420 392
rect 1502 396 1508 397
rect 1502 392 1503 396
rect 1507 392 1508 396
rect 1502 391 1508 392
rect 1590 396 1596 397
rect 1590 392 1591 396
rect 1595 392 1596 396
rect 1590 391 1596 392
rect 1670 396 1676 397
rect 1670 392 1671 396
rect 1675 392 1676 396
rect 1670 391 1676 392
rect 1750 396 1756 397
rect 1750 392 1751 396
rect 1755 392 1756 396
rect 1750 391 1756 392
rect 1830 396 1836 397
rect 1830 392 1831 396
rect 1835 392 1836 396
rect 1830 391 1836 392
rect 1910 396 1916 397
rect 1910 392 1911 396
rect 1915 392 1916 396
rect 1910 391 1916 392
rect 1998 396 2004 397
rect 1998 392 1999 396
rect 2003 392 2004 396
rect 1998 391 2004 392
rect 2070 396 2076 397
rect 2070 392 2071 396
rect 2075 392 2076 396
rect 2070 391 2076 392
rect 350 390 356 391
rect 1183 387 1189 388
rect 362 383 368 384
rect 362 379 363 383
rect 367 382 368 383
rect 1183 383 1184 387
rect 1188 386 1189 387
rect 1206 387 1212 388
rect 1206 386 1207 387
rect 1188 384 1207 386
rect 1188 383 1189 384
rect 1183 382 1189 383
rect 1206 383 1207 384
rect 1211 383 1212 387
rect 1206 382 1212 383
rect 1223 387 1229 388
rect 1223 383 1224 387
rect 1228 386 1229 387
rect 1231 387 1237 388
rect 1231 386 1232 387
rect 1228 384 1232 386
rect 1228 383 1229 384
rect 1223 382 1229 383
rect 1231 383 1232 384
rect 1236 383 1237 387
rect 1231 382 1237 383
rect 1279 387 1285 388
rect 1279 383 1280 387
rect 1284 386 1285 387
rect 1287 387 1293 388
rect 1287 386 1288 387
rect 1284 384 1288 386
rect 1284 383 1285 384
rect 1279 382 1285 383
rect 1287 383 1288 384
rect 1292 383 1293 387
rect 1287 382 1293 383
rect 1359 387 1365 388
rect 1359 383 1360 387
rect 1364 386 1365 387
rect 1367 387 1373 388
rect 1367 386 1368 387
rect 1364 384 1368 386
rect 1364 383 1365 384
rect 1359 382 1365 383
rect 1367 383 1368 384
rect 1372 383 1373 387
rect 1367 382 1373 383
rect 1439 387 1445 388
rect 1439 383 1440 387
rect 1444 386 1445 387
rect 1447 387 1453 388
rect 1447 386 1448 387
rect 1444 384 1448 386
rect 1444 383 1445 384
rect 1439 382 1445 383
rect 1447 383 1448 384
rect 1452 383 1453 387
rect 1527 387 1533 388
rect 1527 386 1528 387
rect 1447 382 1453 383
rect 1519 384 1528 386
rect 367 380 594 382
rect 367 379 368 380
rect 362 378 368 379
rect 592 376 594 380
rect 1342 379 1348 380
rect 198 375 205 376
rect 198 371 199 375
rect 204 371 205 375
rect 198 370 205 371
rect 222 375 228 376
rect 222 371 223 375
rect 227 374 228 375
rect 239 375 245 376
rect 239 374 240 375
rect 227 372 240 374
rect 227 371 228 372
rect 222 370 228 371
rect 239 371 240 372
rect 244 371 245 375
rect 239 370 245 371
rect 247 375 253 376
rect 247 371 248 375
rect 252 374 253 375
rect 295 375 301 376
rect 295 374 296 375
rect 252 372 296 374
rect 252 371 253 372
rect 247 370 253 371
rect 295 371 296 372
rect 300 371 301 375
rect 295 370 301 371
rect 303 375 309 376
rect 303 371 304 375
rect 308 374 309 375
rect 359 375 365 376
rect 359 374 360 375
rect 308 372 360 374
rect 308 371 309 372
rect 303 370 309 371
rect 359 371 360 372
rect 364 371 365 375
rect 359 370 365 371
rect 431 375 437 376
rect 431 371 432 375
rect 436 374 437 375
rect 502 375 508 376
rect 502 374 503 375
rect 436 372 503 374
rect 436 371 437 372
rect 431 370 437 371
rect 502 371 503 372
rect 507 371 508 375
rect 502 370 508 371
rect 511 375 517 376
rect 511 371 512 375
rect 516 374 517 375
rect 582 375 588 376
rect 582 374 583 375
rect 516 372 583 374
rect 516 371 517 372
rect 511 370 517 371
rect 582 371 583 372
rect 587 371 588 375
rect 582 370 588 371
rect 591 375 597 376
rect 591 371 592 375
rect 596 371 597 375
rect 591 370 597 371
rect 663 375 669 376
rect 663 371 664 375
rect 668 374 669 375
rect 726 375 732 376
rect 726 374 727 375
rect 668 372 727 374
rect 668 371 669 372
rect 663 370 669 371
rect 726 371 727 372
rect 731 371 732 375
rect 726 370 732 371
rect 735 375 741 376
rect 735 371 736 375
rect 740 374 741 375
rect 790 375 796 376
rect 790 374 791 375
rect 740 372 791 374
rect 740 371 741 372
rect 735 370 741 371
rect 790 371 791 372
rect 795 371 796 375
rect 790 370 796 371
rect 799 375 805 376
rect 799 371 800 375
rect 804 374 805 375
rect 854 375 860 376
rect 854 374 855 375
rect 804 372 855 374
rect 804 371 805 372
rect 799 370 805 371
rect 854 371 855 372
rect 859 371 860 375
rect 854 370 860 371
rect 863 375 869 376
rect 863 371 864 375
rect 868 374 869 375
rect 886 375 892 376
rect 886 374 887 375
rect 868 372 887 374
rect 868 371 869 372
rect 863 370 869 371
rect 886 371 887 372
rect 891 371 892 375
rect 886 370 892 371
rect 919 375 925 376
rect 919 371 920 375
rect 924 374 925 375
rect 966 375 972 376
rect 966 374 967 375
rect 924 372 967 374
rect 924 371 925 372
rect 919 370 925 371
rect 966 371 967 372
rect 971 371 972 375
rect 966 370 972 371
rect 975 375 981 376
rect 975 371 976 375
rect 980 374 981 375
rect 1022 375 1028 376
rect 1022 374 1023 375
rect 980 372 1023 374
rect 980 371 981 372
rect 975 370 981 371
rect 1022 371 1023 372
rect 1027 371 1028 375
rect 1022 370 1028 371
rect 1030 375 1037 376
rect 1030 371 1031 375
rect 1036 371 1037 375
rect 1030 370 1037 371
rect 1071 375 1077 376
rect 1071 371 1072 375
rect 1076 374 1077 375
rect 1182 375 1188 376
rect 1182 374 1183 375
rect 1076 372 1183 374
rect 1076 371 1077 372
rect 1071 370 1077 371
rect 1182 371 1183 372
rect 1187 371 1188 375
rect 1342 375 1343 379
rect 1347 378 1348 379
rect 1519 378 1521 384
rect 1527 383 1528 384
rect 1532 383 1533 387
rect 1527 382 1533 383
rect 1610 387 1621 388
rect 1610 383 1611 387
rect 1615 383 1616 387
rect 1620 383 1621 387
rect 1610 382 1621 383
rect 1695 387 1701 388
rect 1695 383 1696 387
rect 1700 386 1701 387
rect 1706 387 1712 388
rect 1706 386 1707 387
rect 1700 384 1707 386
rect 1700 383 1701 384
rect 1695 382 1701 383
rect 1706 383 1707 384
rect 1711 383 1712 387
rect 1706 382 1712 383
rect 1775 387 1781 388
rect 1775 383 1776 387
rect 1780 386 1781 387
rect 1783 387 1789 388
rect 1783 386 1784 387
rect 1780 384 1784 386
rect 1780 383 1781 384
rect 1775 382 1781 383
rect 1783 383 1784 384
rect 1788 383 1789 387
rect 1783 382 1789 383
rect 1854 387 1861 388
rect 1854 383 1855 387
rect 1860 383 1861 387
rect 1854 382 1861 383
rect 1935 387 1944 388
rect 1935 383 1936 387
rect 1943 383 1944 387
rect 1935 382 1944 383
rect 2010 387 2016 388
rect 2010 383 2011 387
rect 2015 386 2016 387
rect 2023 387 2029 388
rect 2023 386 2024 387
rect 2015 384 2024 386
rect 2015 383 2016 384
rect 2010 382 2016 383
rect 2023 383 2024 384
rect 2028 383 2029 387
rect 2023 382 2029 383
rect 2094 387 2101 388
rect 2094 383 2095 387
rect 2100 383 2101 387
rect 2094 382 2101 383
rect 1347 376 1521 378
rect 1347 375 1348 376
rect 1342 374 1348 375
rect 1182 370 1188 371
rect 174 368 180 369
rect 174 364 175 368
rect 179 364 180 368
rect 174 363 180 364
rect 214 368 220 369
rect 214 364 215 368
rect 219 364 220 368
rect 214 363 220 364
rect 270 368 276 369
rect 270 364 271 368
rect 275 364 276 368
rect 270 363 276 364
rect 334 368 340 369
rect 334 364 335 368
rect 339 364 340 368
rect 334 363 340 364
rect 406 368 412 369
rect 406 364 407 368
rect 411 364 412 368
rect 406 363 412 364
rect 486 368 492 369
rect 486 364 487 368
rect 491 364 492 368
rect 486 363 492 364
rect 566 368 572 369
rect 566 364 567 368
rect 571 364 572 368
rect 566 363 572 364
rect 638 368 644 369
rect 638 364 639 368
rect 643 364 644 368
rect 638 363 644 364
rect 710 368 716 369
rect 710 364 711 368
rect 715 364 716 368
rect 710 363 716 364
rect 774 368 780 369
rect 774 364 775 368
rect 779 364 780 368
rect 774 363 780 364
rect 838 368 844 369
rect 838 364 839 368
rect 843 364 844 368
rect 838 363 844 364
rect 894 368 900 369
rect 894 364 895 368
rect 899 364 900 368
rect 894 363 900 364
rect 950 368 956 369
rect 950 364 951 368
rect 955 364 956 368
rect 950 363 956 364
rect 1006 368 1012 369
rect 1006 364 1007 368
rect 1011 364 1012 368
rect 1006 363 1012 364
rect 1046 368 1052 369
rect 1046 364 1047 368
rect 1051 364 1052 368
rect 1686 367 1692 368
rect 1686 366 1687 367
rect 1671 365 1687 366
rect 1046 363 1052 364
rect 1183 363 1189 364
rect 110 360 116 361
rect 110 356 111 360
rect 115 356 116 360
rect 1094 360 1100 361
rect 1094 356 1095 360
rect 1099 356 1100 360
rect 1183 359 1184 363
rect 1188 362 1189 363
rect 1262 363 1268 364
rect 1262 362 1263 363
rect 1188 360 1263 362
rect 1188 359 1189 360
rect 1183 358 1189 359
rect 1262 359 1263 360
rect 1267 359 1268 363
rect 1262 358 1268 359
rect 1271 363 1277 364
rect 1271 359 1272 363
rect 1276 362 1277 363
rect 1326 363 1332 364
rect 1326 362 1327 363
rect 1276 360 1327 362
rect 1276 359 1277 360
rect 1271 358 1277 359
rect 1326 359 1327 360
rect 1331 359 1332 363
rect 1326 358 1332 359
rect 1383 363 1389 364
rect 1383 359 1384 363
rect 1388 362 1389 363
rect 1478 363 1484 364
rect 1478 362 1479 363
rect 1388 360 1479 362
rect 1388 359 1389 360
rect 1383 358 1389 359
rect 1478 359 1479 360
rect 1483 359 1484 363
rect 1478 358 1484 359
rect 1486 363 1493 364
rect 1486 359 1487 363
rect 1492 359 1493 363
rect 1486 358 1493 359
rect 1583 363 1589 364
rect 1583 359 1584 363
rect 1588 362 1589 363
rect 1662 363 1668 364
rect 1662 362 1663 363
rect 1588 360 1663 362
rect 1588 359 1589 360
rect 1583 358 1589 359
rect 1662 359 1663 360
rect 1667 359 1668 363
rect 1671 361 1672 365
rect 1676 364 1687 365
rect 1676 361 1677 364
rect 1686 363 1687 364
rect 1691 363 1692 367
rect 1686 362 1692 363
rect 1751 363 1757 364
rect 1751 362 1752 363
rect 1671 360 1677 361
rect 1696 360 1752 362
rect 1662 358 1668 359
rect 110 355 116 356
rect 199 355 205 356
rect 199 351 200 355
rect 204 354 205 355
rect 222 355 228 356
rect 222 354 223 355
rect 204 352 223 354
rect 204 351 205 352
rect 199 350 205 351
rect 222 351 223 352
rect 227 351 228 355
rect 222 350 228 351
rect 239 355 245 356
rect 239 351 240 355
rect 244 354 245 355
rect 247 355 253 356
rect 247 354 248 355
rect 244 352 248 354
rect 244 351 245 352
rect 239 350 245 351
rect 247 351 248 352
rect 252 351 253 355
rect 247 350 253 351
rect 295 355 301 356
rect 295 351 296 355
rect 300 354 301 355
rect 303 355 309 356
rect 303 354 304 355
rect 300 352 304 354
rect 300 351 301 352
rect 295 350 301 351
rect 303 351 304 352
rect 308 351 309 355
rect 303 350 309 351
rect 359 355 368 356
rect 359 351 360 355
rect 367 351 368 355
rect 359 350 368 351
rect 430 355 437 356
rect 430 351 431 355
rect 436 351 437 355
rect 430 350 437 351
rect 502 355 508 356
rect 502 351 503 355
rect 507 354 508 355
rect 511 355 517 356
rect 511 354 512 355
rect 507 352 512 354
rect 507 351 508 352
rect 502 350 508 351
rect 511 351 512 352
rect 516 351 517 355
rect 511 350 517 351
rect 582 355 588 356
rect 582 351 583 355
rect 587 354 588 355
rect 591 355 597 356
rect 591 354 592 355
rect 587 352 592 354
rect 587 351 588 352
rect 582 350 588 351
rect 591 351 592 352
rect 596 351 597 355
rect 591 350 597 351
rect 663 355 672 356
rect 663 351 664 355
rect 671 351 672 355
rect 663 350 672 351
rect 726 355 732 356
rect 726 351 727 355
rect 731 354 732 355
rect 735 355 741 356
rect 735 354 736 355
rect 731 352 736 354
rect 731 351 732 352
rect 726 350 732 351
rect 735 351 736 352
rect 740 351 741 355
rect 735 350 741 351
rect 790 355 796 356
rect 790 351 791 355
rect 795 354 796 355
rect 799 355 805 356
rect 799 354 800 355
rect 795 352 800 354
rect 795 351 796 352
rect 790 350 796 351
rect 799 351 800 352
rect 804 351 805 355
rect 799 350 805 351
rect 854 355 860 356
rect 854 351 855 355
rect 859 354 860 355
rect 863 355 869 356
rect 863 354 864 355
rect 859 352 864 354
rect 859 351 860 352
rect 854 350 860 351
rect 863 351 864 352
rect 868 351 869 355
rect 863 350 869 351
rect 886 355 892 356
rect 886 351 887 355
rect 891 354 892 355
rect 919 355 925 356
rect 919 354 920 355
rect 891 352 920 354
rect 891 351 892 352
rect 886 350 892 351
rect 919 351 920 352
rect 924 351 925 355
rect 919 350 925 351
rect 966 355 972 356
rect 966 351 967 355
rect 971 354 972 355
rect 975 355 981 356
rect 975 354 976 355
rect 971 352 976 354
rect 971 351 972 352
rect 966 350 972 351
rect 975 351 976 352
rect 980 351 981 355
rect 975 350 981 351
rect 1022 355 1028 356
rect 1022 351 1023 355
rect 1027 354 1028 355
rect 1031 355 1037 356
rect 1031 354 1032 355
rect 1027 352 1032 354
rect 1027 351 1028 352
rect 1022 350 1028 351
rect 1031 351 1032 352
rect 1036 351 1037 355
rect 1031 350 1037 351
rect 1070 355 1077 356
rect 1094 355 1100 356
rect 1158 356 1164 357
rect 1070 351 1071 355
rect 1076 351 1077 355
rect 1158 352 1159 356
rect 1163 352 1164 356
rect 1158 351 1164 352
rect 1246 356 1252 357
rect 1246 352 1247 356
rect 1251 352 1252 356
rect 1246 351 1252 352
rect 1358 356 1364 357
rect 1358 352 1359 356
rect 1363 352 1364 356
rect 1358 351 1364 352
rect 1462 356 1468 357
rect 1462 352 1463 356
rect 1467 352 1468 356
rect 1462 351 1468 352
rect 1558 356 1564 357
rect 1558 352 1559 356
rect 1563 352 1564 356
rect 1558 351 1564 352
rect 1646 356 1652 357
rect 1646 352 1647 356
rect 1651 352 1652 356
rect 1696 354 1698 360
rect 1751 359 1752 360
rect 1756 359 1757 363
rect 1751 358 1757 359
rect 1759 363 1765 364
rect 1759 359 1760 363
rect 1764 362 1765 363
rect 1823 363 1829 364
rect 1823 362 1824 363
rect 1764 360 1824 362
rect 1764 359 1765 360
rect 1759 358 1765 359
rect 1823 359 1824 360
rect 1828 359 1829 363
rect 1823 358 1829 359
rect 1831 363 1837 364
rect 1831 359 1832 363
rect 1836 362 1837 363
rect 1887 363 1893 364
rect 1887 362 1888 363
rect 1836 360 1888 362
rect 1836 359 1837 360
rect 1831 358 1837 359
rect 1887 359 1888 360
rect 1892 359 1893 363
rect 1887 358 1893 359
rect 1943 363 1949 364
rect 1943 359 1944 363
rect 1948 362 1949 363
rect 1990 363 1996 364
rect 1990 362 1991 363
rect 1948 360 1991 362
rect 1948 359 1949 360
rect 1943 358 1949 359
rect 1990 359 1991 360
rect 1995 359 1996 363
rect 1990 358 1996 359
rect 1999 363 2005 364
rect 1999 359 2000 363
rect 2004 362 2005 363
rect 2046 363 2052 364
rect 2046 362 2047 363
rect 2004 360 2047 362
rect 2004 359 2005 360
rect 1999 358 2005 359
rect 2046 359 2047 360
rect 2051 359 2052 363
rect 2046 358 2052 359
rect 2055 363 2061 364
rect 2055 359 2056 363
rect 2060 362 2061 363
rect 2086 363 2092 364
rect 2086 362 2087 363
rect 2060 360 2087 362
rect 2060 359 2061 360
rect 2055 358 2061 359
rect 2086 359 2087 360
rect 2091 359 2092 363
rect 2086 358 2092 359
rect 2095 363 2101 364
rect 2095 359 2096 363
rect 2100 362 2101 363
rect 2103 363 2109 364
rect 2103 362 2104 363
rect 2100 360 2104 362
rect 2100 359 2101 360
rect 2095 358 2101 359
rect 2103 359 2104 360
rect 2108 359 2109 363
rect 2103 358 2109 359
rect 1646 351 1652 352
rect 1656 352 1698 354
rect 1726 356 1732 357
rect 1726 352 1727 356
rect 1731 352 1732 356
rect 1070 350 1077 351
rect 1134 348 1140 349
rect 1134 344 1135 348
rect 1139 344 1140 348
rect 110 343 116 344
rect 110 339 111 343
rect 115 339 116 343
rect 1094 343 1100 344
rect 1134 343 1140 344
rect 1182 343 1189 344
rect 110 338 116 339
rect 174 340 180 341
rect 174 336 175 340
rect 179 336 180 340
rect 174 335 180 336
rect 214 340 220 341
rect 214 336 215 340
rect 219 336 220 340
rect 214 335 220 336
rect 270 340 276 341
rect 270 336 271 340
rect 275 336 276 340
rect 270 335 276 336
rect 334 340 340 341
rect 334 336 335 340
rect 339 336 340 340
rect 334 335 340 336
rect 406 340 412 341
rect 406 336 407 340
rect 411 336 412 340
rect 406 335 412 336
rect 486 340 492 341
rect 486 336 487 340
rect 491 336 492 340
rect 486 335 492 336
rect 566 340 572 341
rect 566 336 567 340
rect 571 336 572 340
rect 566 335 572 336
rect 638 340 644 341
rect 638 336 639 340
rect 643 336 644 340
rect 638 335 644 336
rect 710 340 716 341
rect 710 336 711 340
rect 715 336 716 340
rect 710 335 716 336
rect 774 340 780 341
rect 774 336 775 340
rect 779 336 780 340
rect 774 335 780 336
rect 838 340 844 341
rect 838 336 839 340
rect 843 336 844 340
rect 838 335 844 336
rect 894 340 900 341
rect 894 336 895 340
rect 899 336 900 340
rect 894 335 900 336
rect 950 340 956 341
rect 950 336 951 340
rect 955 336 956 340
rect 950 335 956 336
rect 1006 340 1012 341
rect 1006 336 1007 340
rect 1011 336 1012 340
rect 1006 335 1012 336
rect 1046 340 1052 341
rect 1046 336 1047 340
rect 1051 336 1052 340
rect 1094 339 1095 343
rect 1099 339 1100 343
rect 1094 338 1100 339
rect 1182 339 1183 343
rect 1188 339 1189 343
rect 1182 338 1189 339
rect 1262 343 1268 344
rect 1262 339 1263 343
rect 1267 342 1268 343
rect 1271 343 1277 344
rect 1271 342 1272 343
rect 1267 340 1272 342
rect 1267 339 1268 340
rect 1262 338 1268 339
rect 1271 339 1272 340
rect 1276 339 1277 343
rect 1271 338 1277 339
rect 1326 343 1332 344
rect 1326 339 1327 343
rect 1331 342 1332 343
rect 1383 343 1389 344
rect 1383 342 1384 343
rect 1331 340 1384 342
rect 1331 339 1332 340
rect 1326 338 1332 339
rect 1383 339 1384 340
rect 1388 339 1389 343
rect 1383 338 1389 339
rect 1478 343 1484 344
rect 1478 339 1479 343
rect 1483 342 1484 343
rect 1487 343 1493 344
rect 1487 342 1488 343
rect 1483 340 1488 342
rect 1483 339 1484 340
rect 1478 338 1484 339
rect 1487 339 1488 340
rect 1492 339 1493 343
rect 1487 338 1493 339
rect 1583 343 1589 344
rect 1583 339 1584 343
rect 1588 342 1589 343
rect 1656 342 1658 352
rect 1726 351 1732 352
rect 1798 356 1804 357
rect 1798 352 1799 356
rect 1803 352 1804 356
rect 1798 351 1804 352
rect 1862 356 1868 357
rect 1862 352 1863 356
rect 1867 352 1868 356
rect 1862 351 1868 352
rect 1918 356 1924 357
rect 1918 352 1919 356
rect 1923 352 1924 356
rect 1918 351 1924 352
rect 1974 356 1980 357
rect 1974 352 1975 356
rect 1979 352 1980 356
rect 1974 351 1980 352
rect 2030 356 2036 357
rect 2030 352 2031 356
rect 2035 352 2036 356
rect 2030 351 2036 352
rect 2070 356 2076 357
rect 2070 352 2071 356
rect 2075 352 2076 356
rect 2070 351 2076 352
rect 2118 348 2124 349
rect 2118 344 2119 348
rect 2123 344 2124 348
rect 1588 340 1658 342
rect 1662 343 1668 344
rect 1588 339 1589 340
rect 1583 338 1589 339
rect 1662 339 1663 343
rect 1667 342 1668 343
rect 1671 343 1677 344
rect 1671 342 1672 343
rect 1667 340 1672 342
rect 1667 339 1668 340
rect 1662 338 1668 339
rect 1671 339 1672 340
rect 1676 339 1677 343
rect 1671 338 1677 339
rect 1751 343 1757 344
rect 1751 339 1752 343
rect 1756 342 1757 343
rect 1759 343 1765 344
rect 1759 342 1760 343
rect 1756 340 1760 342
rect 1756 339 1757 340
rect 1751 338 1757 339
rect 1759 339 1760 340
rect 1764 339 1765 343
rect 1759 338 1765 339
rect 1823 343 1829 344
rect 1823 339 1824 343
rect 1828 342 1829 343
rect 1831 343 1837 344
rect 1831 342 1832 343
rect 1828 340 1832 342
rect 1828 339 1829 340
rect 1823 338 1829 339
rect 1831 339 1832 340
rect 1836 339 1837 343
rect 1831 338 1837 339
rect 1887 343 1893 344
rect 1887 339 1888 343
rect 1892 342 1893 343
rect 1910 343 1916 344
rect 1910 342 1911 343
rect 1892 340 1911 342
rect 1892 339 1893 340
rect 1887 338 1893 339
rect 1910 339 1911 340
rect 1915 339 1916 343
rect 1910 338 1916 339
rect 1938 343 1949 344
rect 1938 339 1939 343
rect 1943 339 1944 343
rect 1948 339 1949 343
rect 1938 338 1949 339
rect 1990 343 1996 344
rect 1990 339 1991 343
rect 1995 342 1996 343
rect 1999 343 2005 344
rect 1999 342 2000 343
rect 1995 340 2000 342
rect 1995 339 1996 340
rect 1990 338 1996 339
rect 1999 339 2000 340
rect 2004 339 2005 343
rect 1999 338 2005 339
rect 2046 343 2052 344
rect 2046 339 2047 343
rect 2051 342 2052 343
rect 2055 343 2061 344
rect 2055 342 2056 343
rect 2051 340 2056 342
rect 2051 339 2052 340
rect 2046 338 2052 339
rect 2055 339 2056 340
rect 2060 339 2061 343
rect 2055 338 2061 339
rect 2086 343 2092 344
rect 2086 339 2087 343
rect 2091 342 2092 343
rect 2095 343 2101 344
rect 2118 343 2124 344
rect 2095 342 2096 343
rect 2091 340 2096 342
rect 2091 339 2092 340
rect 2086 338 2092 339
rect 2095 339 2096 340
rect 2100 339 2101 343
rect 2095 338 2101 339
rect 1046 335 1052 336
rect 1134 331 1140 332
rect 1134 327 1135 331
rect 1139 327 1140 331
rect 2118 331 2124 332
rect 1134 326 1140 327
rect 1158 328 1164 329
rect 382 324 388 325
rect 110 321 116 322
rect 110 317 111 321
rect 115 317 116 321
rect 382 320 383 324
rect 387 320 388 324
rect 382 319 388 320
rect 422 324 428 325
rect 422 320 423 324
rect 427 320 428 324
rect 422 319 428 320
rect 462 324 468 325
rect 462 320 463 324
rect 467 320 468 324
rect 462 319 468 320
rect 502 324 508 325
rect 502 320 503 324
rect 507 320 508 324
rect 502 319 508 320
rect 542 324 548 325
rect 542 320 543 324
rect 547 320 548 324
rect 542 319 548 320
rect 590 324 596 325
rect 590 320 591 324
rect 595 320 596 324
rect 590 319 596 320
rect 638 324 644 325
rect 638 320 639 324
rect 643 320 644 324
rect 638 319 644 320
rect 686 324 692 325
rect 686 320 687 324
rect 691 320 692 324
rect 686 319 692 320
rect 734 324 740 325
rect 734 320 735 324
rect 739 320 740 324
rect 734 319 740 320
rect 782 324 788 325
rect 782 320 783 324
rect 787 320 788 324
rect 782 319 788 320
rect 830 324 836 325
rect 830 320 831 324
rect 835 320 836 324
rect 830 319 836 320
rect 878 324 884 325
rect 878 320 879 324
rect 883 320 884 324
rect 878 319 884 320
rect 926 324 932 325
rect 926 320 927 324
rect 931 320 932 324
rect 926 319 932 320
rect 966 324 972 325
rect 966 320 967 324
rect 971 320 972 324
rect 966 319 972 320
rect 1006 324 1012 325
rect 1006 320 1007 324
rect 1011 320 1012 324
rect 1006 319 1012 320
rect 1046 324 1052 325
rect 1046 320 1047 324
rect 1051 320 1052 324
rect 1158 324 1159 328
rect 1163 324 1164 328
rect 1158 323 1164 324
rect 1246 328 1252 329
rect 1246 324 1247 328
rect 1251 324 1252 328
rect 1246 323 1252 324
rect 1358 328 1364 329
rect 1358 324 1359 328
rect 1363 324 1364 328
rect 1358 323 1364 324
rect 1462 328 1468 329
rect 1462 324 1463 328
rect 1467 324 1468 328
rect 1462 323 1468 324
rect 1558 328 1564 329
rect 1558 324 1559 328
rect 1563 324 1564 328
rect 1558 323 1564 324
rect 1646 328 1652 329
rect 1646 324 1647 328
rect 1651 324 1652 328
rect 1646 323 1652 324
rect 1726 328 1732 329
rect 1726 324 1727 328
rect 1731 324 1732 328
rect 1726 323 1732 324
rect 1798 328 1804 329
rect 1798 324 1799 328
rect 1803 324 1804 328
rect 1798 323 1804 324
rect 1862 328 1868 329
rect 1862 324 1863 328
rect 1867 324 1868 328
rect 1862 323 1868 324
rect 1918 328 1924 329
rect 1918 324 1919 328
rect 1923 324 1924 328
rect 1918 323 1924 324
rect 1974 328 1980 329
rect 1974 324 1975 328
rect 1979 324 1980 328
rect 1974 323 1980 324
rect 2030 328 2036 329
rect 2030 324 2031 328
rect 2035 324 2036 328
rect 2030 323 2036 324
rect 2070 328 2076 329
rect 2070 324 2071 328
rect 2075 324 2076 328
rect 2118 327 2119 331
rect 2123 327 2124 331
rect 2118 326 2124 327
rect 2070 323 2076 324
rect 1046 319 1052 320
rect 1094 321 1100 322
rect 110 316 116 317
rect 1094 317 1095 321
rect 1099 317 1100 321
rect 1094 316 1100 317
rect 1030 315 1036 316
rect 1030 314 1031 315
rect 953 312 1031 314
rect 953 308 955 312
rect 1030 311 1031 312
rect 1035 311 1036 315
rect 1030 310 1036 311
rect 1350 308 1356 309
rect 406 307 413 308
rect 110 304 116 305
rect 110 300 111 304
rect 115 300 116 304
rect 406 303 407 307
rect 412 303 413 307
rect 406 302 413 303
rect 430 307 436 308
rect 430 303 431 307
rect 435 306 436 307
rect 447 307 453 308
rect 447 306 448 307
rect 435 304 448 306
rect 435 303 436 304
rect 430 302 436 303
rect 447 303 448 304
rect 452 303 453 307
rect 447 302 453 303
rect 470 307 476 308
rect 470 303 471 307
rect 475 306 476 307
rect 487 307 493 308
rect 487 306 488 307
rect 475 304 488 306
rect 475 303 476 304
rect 470 302 476 303
rect 487 303 488 304
rect 492 303 493 307
rect 487 302 493 303
rect 510 307 516 308
rect 510 303 511 307
rect 515 306 516 307
rect 527 307 533 308
rect 527 306 528 307
rect 515 304 528 306
rect 515 303 516 304
rect 510 302 516 303
rect 527 303 528 304
rect 532 303 533 307
rect 527 302 533 303
rect 550 307 556 308
rect 550 303 551 307
rect 555 306 556 307
rect 567 307 573 308
rect 567 306 568 307
rect 555 304 568 306
rect 555 303 556 304
rect 550 302 556 303
rect 567 303 568 304
rect 572 303 573 307
rect 567 302 573 303
rect 575 307 581 308
rect 575 303 576 307
rect 580 306 581 307
rect 615 307 621 308
rect 615 306 616 307
rect 580 304 616 306
rect 580 303 581 304
rect 575 302 581 303
rect 615 303 616 304
rect 620 303 621 307
rect 615 302 621 303
rect 623 307 629 308
rect 623 303 624 307
rect 628 306 629 307
rect 663 307 669 308
rect 663 306 664 307
rect 628 304 664 306
rect 628 303 629 304
rect 623 302 629 303
rect 663 303 664 304
rect 668 303 669 307
rect 663 302 669 303
rect 671 307 677 308
rect 671 303 672 307
rect 676 306 677 307
rect 711 307 717 308
rect 711 306 712 307
rect 676 304 712 306
rect 676 303 677 304
rect 671 302 677 303
rect 711 303 712 304
rect 716 303 717 307
rect 711 302 717 303
rect 759 307 768 308
rect 759 303 760 307
rect 767 303 768 307
rect 759 302 768 303
rect 770 307 776 308
rect 770 303 771 307
rect 775 306 776 307
rect 807 307 813 308
rect 807 306 808 307
rect 775 304 808 306
rect 775 303 776 304
rect 770 302 776 303
rect 807 303 808 304
rect 812 303 813 307
rect 807 302 813 303
rect 815 307 821 308
rect 815 303 816 307
rect 820 306 821 307
rect 855 307 861 308
rect 855 306 856 307
rect 820 304 856 306
rect 820 303 821 304
rect 815 302 821 303
rect 855 303 856 304
rect 860 303 861 307
rect 855 302 861 303
rect 863 307 869 308
rect 863 303 864 307
rect 868 306 869 307
rect 903 307 909 308
rect 903 306 904 307
rect 868 304 904 306
rect 868 303 869 304
rect 863 302 869 303
rect 903 303 904 304
rect 908 303 909 307
rect 903 302 909 303
rect 951 307 957 308
rect 951 303 952 307
rect 956 303 957 307
rect 951 302 957 303
rect 974 307 980 308
rect 974 303 975 307
rect 979 306 980 307
rect 991 307 997 308
rect 991 306 992 307
rect 979 304 992 306
rect 979 303 980 304
rect 974 302 980 303
rect 991 303 992 304
rect 996 303 997 307
rect 991 302 997 303
rect 1014 307 1020 308
rect 1014 303 1015 307
rect 1019 306 1020 307
rect 1031 307 1037 308
rect 1031 306 1032 307
rect 1019 304 1032 306
rect 1019 303 1020 304
rect 1014 302 1020 303
rect 1031 303 1032 304
rect 1036 303 1037 307
rect 1031 302 1037 303
rect 1054 307 1060 308
rect 1054 303 1055 307
rect 1059 306 1060 307
rect 1071 307 1077 308
rect 1071 306 1072 307
rect 1059 304 1072 306
rect 1059 303 1060 304
rect 1054 302 1060 303
rect 1071 303 1072 304
rect 1076 303 1077 307
rect 1134 305 1140 306
rect 1071 302 1077 303
rect 1094 304 1100 305
rect 110 299 116 300
rect 1094 300 1095 304
rect 1099 300 1100 304
rect 1134 301 1135 305
rect 1139 301 1140 305
rect 1350 304 1351 308
rect 1355 304 1356 308
rect 1350 303 1356 304
rect 1390 308 1396 309
rect 1390 304 1391 308
rect 1395 304 1396 308
rect 1390 303 1396 304
rect 1430 308 1436 309
rect 1430 304 1431 308
rect 1435 304 1436 308
rect 1430 303 1436 304
rect 1470 308 1476 309
rect 1470 304 1471 308
rect 1475 304 1476 308
rect 1470 303 1476 304
rect 1510 308 1516 309
rect 1510 304 1511 308
rect 1515 304 1516 308
rect 1510 303 1516 304
rect 1558 308 1564 309
rect 1558 304 1559 308
rect 1563 304 1564 308
rect 1558 303 1564 304
rect 1614 308 1620 309
rect 1614 304 1615 308
rect 1619 304 1620 308
rect 1614 303 1620 304
rect 1670 308 1676 309
rect 1670 304 1671 308
rect 1675 304 1676 308
rect 1670 303 1676 304
rect 1734 308 1740 309
rect 1734 304 1735 308
rect 1739 304 1740 308
rect 1734 303 1740 304
rect 1806 308 1812 309
rect 1806 304 1807 308
rect 1811 304 1812 308
rect 1806 303 1812 304
rect 1886 308 1892 309
rect 1886 304 1887 308
rect 1891 304 1892 308
rect 1886 303 1892 304
rect 1966 308 1972 309
rect 1966 304 1967 308
rect 1971 304 1972 308
rect 1966 303 1972 304
rect 2046 308 2052 309
rect 2046 304 2047 308
rect 2051 304 2052 308
rect 2046 303 2052 304
rect 2118 305 2124 306
rect 1134 300 1140 301
rect 2118 301 2119 305
rect 2123 301 2124 305
rect 2118 300 2124 301
rect 1094 299 1100 300
rect 382 296 388 297
rect 382 292 383 296
rect 387 292 388 296
rect 382 291 388 292
rect 422 296 428 297
rect 422 292 423 296
rect 427 292 428 296
rect 422 291 428 292
rect 462 296 468 297
rect 462 292 463 296
rect 467 292 468 296
rect 462 291 468 292
rect 502 296 508 297
rect 502 292 503 296
rect 507 292 508 296
rect 502 291 508 292
rect 542 296 548 297
rect 542 292 543 296
rect 547 292 548 296
rect 542 291 548 292
rect 590 296 596 297
rect 590 292 591 296
rect 595 292 596 296
rect 590 291 596 292
rect 638 296 644 297
rect 638 292 639 296
rect 643 292 644 296
rect 638 291 644 292
rect 686 296 692 297
rect 686 292 687 296
rect 691 292 692 296
rect 686 291 692 292
rect 734 296 740 297
rect 734 292 735 296
rect 739 292 740 296
rect 734 291 740 292
rect 782 296 788 297
rect 782 292 783 296
rect 787 292 788 296
rect 782 291 788 292
rect 830 296 836 297
rect 830 292 831 296
rect 835 292 836 296
rect 830 291 836 292
rect 878 296 884 297
rect 878 292 879 296
rect 883 292 884 296
rect 878 291 884 292
rect 926 296 932 297
rect 926 292 927 296
rect 931 292 932 296
rect 926 291 932 292
rect 966 296 972 297
rect 966 292 967 296
rect 971 292 972 296
rect 966 291 972 292
rect 1006 296 1012 297
rect 1006 292 1007 296
rect 1011 292 1012 296
rect 1006 291 1012 292
rect 1046 296 1052 297
rect 1046 292 1047 296
rect 1051 292 1052 296
rect 1046 291 1052 292
rect 1374 291 1381 292
rect 1134 288 1140 289
rect 407 287 413 288
rect 407 283 408 287
rect 412 286 413 287
rect 430 287 436 288
rect 430 286 431 287
rect 412 284 431 286
rect 412 283 413 284
rect 407 282 413 283
rect 430 283 431 284
rect 435 283 436 287
rect 430 282 436 283
rect 447 287 453 288
rect 447 283 448 287
rect 452 286 453 287
rect 470 287 476 288
rect 470 286 471 287
rect 452 284 471 286
rect 452 283 453 284
rect 447 282 453 283
rect 470 283 471 284
rect 475 283 476 287
rect 470 282 476 283
rect 487 287 493 288
rect 487 283 488 287
rect 492 286 493 287
rect 510 287 516 288
rect 510 286 511 287
rect 492 284 511 286
rect 492 283 493 284
rect 487 282 493 283
rect 510 283 511 284
rect 515 283 516 287
rect 510 282 516 283
rect 527 287 533 288
rect 527 283 528 287
rect 532 286 533 287
rect 550 287 556 288
rect 550 286 551 287
rect 532 284 551 286
rect 532 283 533 284
rect 527 282 533 283
rect 550 283 551 284
rect 555 283 556 287
rect 550 282 556 283
rect 567 287 573 288
rect 567 283 568 287
rect 572 286 573 287
rect 575 287 581 288
rect 575 286 576 287
rect 572 284 576 286
rect 572 283 573 284
rect 567 282 573 283
rect 575 283 576 284
rect 580 283 581 287
rect 575 282 581 283
rect 615 287 621 288
rect 615 283 616 287
rect 620 286 621 287
rect 623 287 629 288
rect 623 286 624 287
rect 620 284 624 286
rect 620 283 621 284
rect 615 282 621 283
rect 623 283 624 284
rect 628 283 629 287
rect 623 282 629 283
rect 663 287 669 288
rect 663 283 664 287
rect 668 286 669 287
rect 671 287 677 288
rect 671 286 672 287
rect 668 284 672 286
rect 668 283 669 284
rect 663 282 669 283
rect 671 283 672 284
rect 676 283 677 287
rect 671 282 677 283
rect 706 287 717 288
rect 706 283 707 287
rect 711 283 712 287
rect 716 283 717 287
rect 706 282 717 283
rect 759 287 765 288
rect 759 283 760 287
rect 764 286 765 287
rect 770 287 776 288
rect 770 286 771 287
rect 764 284 771 286
rect 764 283 765 284
rect 759 282 765 283
rect 770 283 771 284
rect 775 283 776 287
rect 770 282 776 283
rect 807 287 813 288
rect 807 283 808 287
rect 812 286 813 287
rect 815 287 821 288
rect 815 286 816 287
rect 812 284 816 286
rect 812 283 813 284
rect 807 282 813 283
rect 815 283 816 284
rect 820 283 821 287
rect 815 282 821 283
rect 855 287 861 288
rect 855 283 856 287
rect 860 286 861 287
rect 863 287 869 288
rect 863 286 864 287
rect 860 284 864 286
rect 860 283 861 284
rect 855 282 861 283
rect 863 283 864 284
rect 868 283 869 287
rect 863 282 869 283
rect 886 287 892 288
rect 886 283 887 287
rect 891 286 892 287
rect 903 287 909 288
rect 903 286 904 287
rect 891 284 904 286
rect 891 283 892 284
rect 886 282 892 283
rect 903 283 904 284
rect 908 283 909 287
rect 903 282 909 283
rect 951 287 957 288
rect 951 283 952 287
rect 956 286 957 287
rect 974 287 980 288
rect 974 286 975 287
rect 956 284 975 286
rect 956 283 957 284
rect 951 282 957 283
rect 974 283 975 284
rect 979 283 980 287
rect 974 282 980 283
rect 991 287 997 288
rect 991 283 992 287
rect 996 286 997 287
rect 1014 287 1020 288
rect 1014 286 1015 287
rect 996 284 1015 286
rect 996 283 997 284
rect 991 282 997 283
rect 1014 283 1015 284
rect 1019 283 1020 287
rect 1014 282 1020 283
rect 1031 287 1037 288
rect 1031 283 1032 287
rect 1036 286 1037 287
rect 1054 287 1060 288
rect 1054 286 1055 287
rect 1036 284 1055 286
rect 1036 283 1037 284
rect 1031 282 1037 283
rect 1054 283 1055 284
rect 1059 283 1060 287
rect 1054 282 1060 283
rect 1070 287 1077 288
rect 1070 283 1071 287
rect 1076 283 1077 287
rect 1134 284 1135 288
rect 1139 284 1140 288
rect 1374 287 1375 291
rect 1380 287 1381 291
rect 1374 286 1381 287
rect 1398 291 1404 292
rect 1398 287 1399 291
rect 1403 290 1404 291
rect 1415 291 1421 292
rect 1415 290 1416 291
rect 1403 288 1416 290
rect 1403 287 1404 288
rect 1398 286 1404 287
rect 1415 287 1416 288
rect 1420 287 1421 291
rect 1415 286 1421 287
rect 1438 291 1444 292
rect 1438 287 1439 291
rect 1443 290 1444 291
rect 1455 291 1461 292
rect 1455 290 1456 291
rect 1443 288 1456 290
rect 1443 287 1444 288
rect 1438 286 1444 287
rect 1455 287 1456 288
rect 1460 287 1461 291
rect 1455 286 1461 287
rect 1478 291 1484 292
rect 1478 287 1479 291
rect 1483 290 1484 291
rect 1495 291 1501 292
rect 1495 290 1496 291
rect 1483 288 1496 290
rect 1483 287 1484 288
rect 1478 286 1484 287
rect 1495 287 1496 288
rect 1500 287 1501 291
rect 1495 286 1501 287
rect 1518 291 1524 292
rect 1518 287 1519 291
rect 1523 290 1524 291
rect 1535 291 1541 292
rect 1535 290 1536 291
rect 1523 288 1536 290
rect 1523 287 1524 288
rect 1518 286 1524 287
rect 1535 287 1536 288
rect 1540 287 1541 291
rect 1535 286 1541 287
rect 1543 291 1549 292
rect 1543 287 1544 291
rect 1548 290 1549 291
rect 1583 291 1589 292
rect 1583 290 1584 291
rect 1548 288 1584 290
rect 1548 287 1549 288
rect 1543 286 1549 287
rect 1583 287 1584 288
rect 1588 287 1589 291
rect 1583 286 1589 287
rect 1591 291 1597 292
rect 1591 287 1592 291
rect 1596 290 1597 291
rect 1639 291 1645 292
rect 1639 290 1640 291
rect 1596 288 1640 290
rect 1596 287 1597 288
rect 1591 286 1597 287
rect 1639 287 1640 288
rect 1644 287 1645 291
rect 1639 286 1645 287
rect 1647 291 1653 292
rect 1647 287 1648 291
rect 1652 290 1653 291
rect 1695 291 1701 292
rect 1695 290 1696 291
rect 1652 288 1696 290
rect 1652 287 1653 288
rect 1647 286 1653 287
rect 1695 287 1696 288
rect 1700 287 1701 291
rect 1695 286 1701 287
rect 1722 291 1728 292
rect 1722 287 1723 291
rect 1727 290 1728 291
rect 1759 291 1765 292
rect 1759 290 1760 291
rect 1727 288 1760 290
rect 1727 287 1728 288
rect 1722 286 1728 287
rect 1759 287 1760 288
rect 1764 287 1765 291
rect 1759 286 1765 287
rect 1767 291 1773 292
rect 1767 287 1768 291
rect 1772 290 1773 291
rect 1831 291 1837 292
rect 1831 290 1832 291
rect 1772 288 1832 290
rect 1772 287 1773 288
rect 1767 286 1773 287
rect 1831 287 1832 288
rect 1836 287 1837 291
rect 1831 286 1837 287
rect 1911 291 1917 292
rect 1911 287 1912 291
rect 1916 290 1917 291
rect 1982 291 1988 292
rect 1982 290 1983 291
rect 1916 288 1983 290
rect 1916 287 1917 288
rect 1911 286 1917 287
rect 1982 287 1983 288
rect 1987 287 1988 291
rect 1982 286 1988 287
rect 1991 291 1997 292
rect 1991 287 1992 291
rect 1996 290 1997 291
rect 2062 291 2068 292
rect 2062 290 2063 291
rect 1996 288 2063 290
rect 1996 287 1997 288
rect 1991 286 1997 287
rect 2062 287 2063 288
rect 2067 287 2068 291
rect 2062 286 2068 287
rect 2071 291 2077 292
rect 2071 287 2072 291
rect 2076 290 2077 291
rect 2094 291 2100 292
rect 2094 290 2095 291
rect 2076 288 2095 290
rect 2076 287 2077 288
rect 2071 286 2077 287
rect 2094 287 2095 288
rect 2099 287 2100 291
rect 2094 286 2100 287
rect 2118 288 2124 289
rect 1134 283 1140 284
rect 2118 284 2119 288
rect 2123 284 2124 288
rect 2118 283 2124 284
rect 1070 282 1077 283
rect 1350 280 1356 281
rect 1350 276 1351 280
rect 1355 276 1356 280
rect 1350 275 1356 276
rect 1390 280 1396 281
rect 1390 276 1391 280
rect 1395 276 1396 280
rect 1390 275 1396 276
rect 1430 280 1436 281
rect 1430 276 1431 280
rect 1435 276 1436 280
rect 1430 275 1436 276
rect 1470 280 1476 281
rect 1470 276 1471 280
rect 1475 276 1476 280
rect 1470 275 1476 276
rect 1510 280 1516 281
rect 1510 276 1511 280
rect 1515 276 1516 280
rect 1510 275 1516 276
rect 1558 280 1564 281
rect 1558 276 1559 280
rect 1563 276 1564 280
rect 1558 275 1564 276
rect 1614 280 1620 281
rect 1614 276 1615 280
rect 1619 276 1620 280
rect 1614 275 1620 276
rect 1670 280 1676 281
rect 1670 276 1671 280
rect 1675 276 1676 280
rect 1670 275 1676 276
rect 1734 280 1740 281
rect 1734 276 1735 280
rect 1739 276 1740 280
rect 1734 275 1740 276
rect 1806 280 1812 281
rect 1806 276 1807 280
rect 1811 276 1812 280
rect 1806 275 1812 276
rect 1886 280 1892 281
rect 1886 276 1887 280
rect 1891 276 1892 280
rect 1886 275 1892 276
rect 1966 280 1972 281
rect 1966 276 1967 280
rect 1971 276 1972 280
rect 1966 275 1972 276
rect 2046 280 2052 281
rect 2046 276 2047 280
rect 2051 276 2052 280
rect 2046 275 2052 276
rect 1375 271 1381 272
rect 406 267 412 268
rect 406 263 407 267
rect 411 266 412 267
rect 1375 267 1376 271
rect 1380 270 1381 271
rect 1398 271 1404 272
rect 1398 270 1399 271
rect 1380 268 1399 270
rect 1380 267 1381 268
rect 1375 266 1381 267
rect 1398 267 1399 268
rect 1403 267 1404 271
rect 1398 266 1404 267
rect 1415 271 1421 272
rect 1415 267 1416 271
rect 1420 270 1421 271
rect 1438 271 1444 272
rect 1438 270 1439 271
rect 1420 268 1439 270
rect 1420 267 1421 268
rect 1415 266 1421 267
rect 1438 267 1439 268
rect 1443 267 1444 271
rect 1438 266 1444 267
rect 1455 271 1461 272
rect 1455 267 1456 271
rect 1460 270 1461 271
rect 1478 271 1484 272
rect 1478 270 1479 271
rect 1460 268 1479 270
rect 1460 267 1461 268
rect 1455 266 1461 267
rect 1478 267 1479 268
rect 1483 267 1484 271
rect 1478 266 1484 267
rect 1495 271 1501 272
rect 1495 267 1496 271
rect 1500 270 1501 271
rect 1518 271 1524 272
rect 1518 270 1519 271
rect 1500 268 1519 270
rect 1500 267 1501 268
rect 1495 266 1501 267
rect 1518 267 1519 268
rect 1523 267 1524 271
rect 1518 266 1524 267
rect 1535 271 1541 272
rect 1535 267 1536 271
rect 1540 270 1541 271
rect 1543 271 1549 272
rect 1543 270 1544 271
rect 1540 268 1544 270
rect 1540 267 1541 268
rect 1535 266 1541 267
rect 1543 267 1544 268
rect 1548 267 1549 271
rect 1543 266 1549 267
rect 1583 271 1589 272
rect 1583 267 1584 271
rect 1588 270 1589 271
rect 1591 271 1597 272
rect 1591 270 1592 271
rect 1588 268 1592 270
rect 1588 267 1589 268
rect 1583 266 1589 267
rect 1591 267 1592 268
rect 1596 267 1597 271
rect 1591 266 1597 267
rect 1639 271 1645 272
rect 1639 267 1640 271
rect 1644 270 1645 271
rect 1647 271 1653 272
rect 1647 270 1648 271
rect 1644 268 1648 270
rect 1644 267 1645 268
rect 1639 266 1645 267
rect 1647 267 1648 268
rect 1652 267 1653 271
rect 1647 266 1653 267
rect 1695 271 1701 272
rect 1695 267 1696 271
rect 1700 270 1701 271
rect 1722 271 1728 272
rect 1722 270 1723 271
rect 1700 268 1723 270
rect 1700 267 1701 268
rect 1695 266 1701 267
rect 1722 267 1723 268
rect 1727 267 1728 271
rect 1722 266 1728 267
rect 1759 271 1765 272
rect 1759 267 1760 271
rect 1764 270 1765 271
rect 1767 271 1773 272
rect 1767 270 1768 271
rect 1764 268 1768 270
rect 1764 267 1765 268
rect 1759 266 1765 267
rect 1767 267 1768 268
rect 1772 267 1773 271
rect 1831 271 1837 272
rect 1831 270 1832 271
rect 1767 266 1773 267
rect 1776 268 1832 270
rect 411 264 634 266
rect 411 263 412 264
rect 406 262 412 263
rect 632 260 634 264
rect 1570 263 1576 264
rect 311 259 317 260
rect 311 255 312 259
rect 316 258 317 259
rect 342 259 348 260
rect 342 258 343 259
rect 316 256 343 258
rect 316 255 317 256
rect 311 254 317 255
rect 342 255 343 256
rect 347 255 348 259
rect 342 254 348 255
rect 351 259 357 260
rect 351 255 352 259
rect 356 258 357 259
rect 374 259 380 260
rect 374 258 375 259
rect 356 256 375 258
rect 356 255 357 256
rect 351 254 357 255
rect 374 255 375 256
rect 379 255 380 259
rect 374 254 380 255
rect 391 259 397 260
rect 391 255 392 259
rect 396 258 397 259
rect 430 259 436 260
rect 430 258 431 259
rect 396 256 431 258
rect 396 255 397 256
rect 391 254 397 255
rect 430 255 431 256
rect 435 255 436 259
rect 430 254 436 255
rect 439 259 445 260
rect 439 255 440 259
rect 444 258 445 259
rect 486 259 492 260
rect 486 258 487 259
rect 444 256 487 258
rect 444 255 445 256
rect 439 254 445 255
rect 486 255 487 256
rect 491 255 492 259
rect 486 254 492 255
rect 495 259 501 260
rect 495 255 496 259
rect 500 258 501 259
rect 550 259 556 260
rect 550 258 551 259
rect 500 256 551 258
rect 500 255 501 256
rect 495 254 501 255
rect 550 255 551 256
rect 555 255 556 259
rect 550 254 556 255
rect 559 259 565 260
rect 559 255 560 259
rect 564 258 565 259
rect 622 259 628 260
rect 622 258 623 259
rect 564 256 623 258
rect 564 255 565 256
rect 559 254 565 255
rect 622 255 623 256
rect 627 255 628 259
rect 622 254 628 255
rect 631 259 637 260
rect 631 255 632 259
rect 636 255 637 259
rect 631 254 637 255
rect 698 259 709 260
rect 698 255 699 259
rect 703 255 704 259
rect 708 255 709 259
rect 698 254 709 255
rect 762 259 773 260
rect 762 255 763 259
rect 767 255 768 259
rect 772 255 773 259
rect 831 259 837 260
rect 831 258 832 259
rect 762 254 773 255
rect 800 256 832 258
rect 286 252 292 253
rect 286 248 287 252
rect 291 248 292 252
rect 286 247 292 248
rect 326 252 332 253
rect 326 248 327 252
rect 331 248 332 252
rect 326 247 332 248
rect 366 252 372 253
rect 366 248 367 252
rect 371 248 372 252
rect 366 247 372 248
rect 414 252 420 253
rect 414 248 415 252
rect 419 248 420 252
rect 414 247 420 248
rect 470 252 476 253
rect 470 248 471 252
rect 475 248 476 252
rect 470 247 476 248
rect 534 252 540 253
rect 534 248 535 252
rect 539 248 540 252
rect 534 247 540 248
rect 606 252 612 253
rect 606 248 607 252
rect 611 248 612 252
rect 606 247 612 248
rect 678 252 684 253
rect 678 248 679 252
rect 683 248 684 252
rect 678 247 684 248
rect 742 252 748 253
rect 742 248 743 252
rect 747 248 748 252
rect 742 247 748 248
rect 800 246 802 256
rect 831 255 832 256
rect 836 255 837 259
rect 831 254 837 255
rect 887 259 893 260
rect 887 255 888 259
rect 892 258 893 259
rect 942 259 948 260
rect 942 258 943 259
rect 892 256 943 258
rect 892 255 893 256
rect 887 254 893 255
rect 942 255 943 256
rect 947 255 948 259
rect 942 254 948 255
rect 951 259 957 260
rect 951 255 952 259
rect 956 258 957 259
rect 1006 259 1012 260
rect 1006 258 1007 259
rect 956 256 1007 258
rect 956 255 957 256
rect 951 254 957 255
rect 1006 255 1007 256
rect 1011 255 1012 259
rect 1006 254 1012 255
rect 1015 259 1021 260
rect 1015 255 1016 259
rect 1020 258 1021 259
rect 1062 259 1068 260
rect 1062 258 1063 259
rect 1020 256 1063 258
rect 1020 255 1021 256
rect 1015 254 1021 255
rect 1062 255 1063 256
rect 1067 255 1068 259
rect 1062 254 1068 255
rect 1070 259 1077 260
rect 1070 255 1071 259
rect 1076 255 1077 259
rect 1070 254 1077 255
rect 1374 259 1380 260
rect 1374 255 1375 259
rect 1379 258 1380 259
rect 1570 259 1571 263
rect 1575 262 1576 263
rect 1776 262 1778 268
rect 1831 267 1832 268
rect 1836 267 1837 271
rect 1831 266 1837 267
rect 1910 271 1917 272
rect 1910 267 1911 271
rect 1916 267 1917 271
rect 1910 266 1917 267
rect 1982 271 1988 272
rect 1982 267 1983 271
rect 1987 270 1988 271
rect 1991 271 1997 272
rect 1991 270 1992 271
rect 1987 268 1992 270
rect 1987 267 1988 268
rect 1982 266 1988 267
rect 1991 267 1992 268
rect 1996 267 1997 271
rect 1991 266 1997 267
rect 2062 271 2068 272
rect 2062 267 2063 271
rect 2067 270 2068 271
rect 2071 271 2077 272
rect 2071 270 2072 271
rect 2067 268 2072 270
rect 2067 267 2068 268
rect 2062 266 2068 267
rect 2071 267 2072 268
rect 2076 267 2077 271
rect 2071 266 2077 267
rect 1575 260 1778 262
rect 1575 259 1576 260
rect 1570 258 1576 259
rect 1379 256 1530 258
rect 1379 255 1380 256
rect 1374 254 1380 255
rect 806 252 812 253
rect 806 248 807 252
rect 811 248 812 252
rect 806 247 812 248
rect 862 252 868 253
rect 862 248 863 252
rect 867 248 868 252
rect 862 247 868 248
rect 926 252 932 253
rect 926 248 927 252
rect 931 248 932 252
rect 926 247 932 248
rect 990 252 996 253
rect 990 248 991 252
rect 995 248 996 252
rect 990 247 996 248
rect 1046 252 1052 253
rect 1528 252 1530 256
rect 1046 248 1047 252
rect 1051 248 1052 252
rect 1046 247 1052 248
rect 1287 251 1293 252
rect 1287 247 1288 251
rect 1292 250 1293 251
rect 1318 251 1324 252
rect 1318 250 1319 251
rect 1292 248 1319 250
rect 1292 247 1293 248
rect 1287 246 1293 247
rect 1318 247 1319 248
rect 1323 247 1324 251
rect 1318 246 1324 247
rect 1327 251 1333 252
rect 1327 247 1328 251
rect 1332 250 1333 251
rect 1358 251 1364 252
rect 1358 250 1359 251
rect 1332 248 1359 250
rect 1332 247 1333 248
rect 1327 246 1333 247
rect 1358 247 1359 248
rect 1363 247 1364 251
rect 1358 246 1364 247
rect 1367 251 1373 252
rect 1367 247 1368 251
rect 1372 250 1373 251
rect 1398 251 1404 252
rect 1398 250 1399 251
rect 1372 248 1399 250
rect 1372 247 1373 248
rect 1367 246 1373 247
rect 1398 247 1399 248
rect 1403 247 1404 251
rect 1398 246 1404 247
rect 1407 251 1413 252
rect 1407 247 1408 251
rect 1412 250 1413 251
rect 1438 251 1444 252
rect 1438 250 1439 251
rect 1412 248 1439 250
rect 1412 247 1413 248
rect 1407 246 1413 247
rect 1438 247 1439 248
rect 1443 247 1444 251
rect 1438 246 1444 247
rect 1447 251 1453 252
rect 1447 247 1448 251
rect 1452 250 1453 251
rect 1478 251 1484 252
rect 1478 250 1479 251
rect 1452 248 1479 250
rect 1452 247 1453 248
rect 1447 246 1453 247
rect 1478 247 1479 248
rect 1483 247 1484 251
rect 1478 246 1484 247
rect 1487 251 1493 252
rect 1487 247 1488 251
rect 1492 250 1493 251
rect 1518 251 1524 252
rect 1518 250 1519 251
rect 1492 248 1519 250
rect 1492 247 1493 248
rect 1487 246 1493 247
rect 1518 247 1519 248
rect 1523 247 1524 251
rect 1518 246 1524 247
rect 1527 251 1533 252
rect 1527 247 1528 251
rect 1532 247 1533 251
rect 1527 246 1533 247
rect 1567 251 1573 252
rect 1567 247 1568 251
rect 1572 250 1573 251
rect 1614 251 1620 252
rect 1614 250 1615 251
rect 1572 248 1615 250
rect 1572 247 1573 248
rect 1567 246 1573 247
rect 1614 247 1615 248
rect 1619 247 1620 251
rect 1614 246 1620 247
rect 1623 251 1629 252
rect 1623 247 1624 251
rect 1628 250 1629 251
rect 1686 251 1692 252
rect 1686 250 1687 251
rect 1628 248 1687 250
rect 1628 247 1629 248
rect 1623 246 1629 247
rect 1686 247 1687 248
rect 1691 247 1692 251
rect 1686 246 1692 247
rect 1695 251 1701 252
rect 1695 247 1696 251
rect 1700 250 1701 251
rect 1774 251 1780 252
rect 1774 250 1775 251
rect 1700 248 1775 250
rect 1700 247 1701 248
rect 1695 246 1701 247
rect 1774 247 1775 248
rect 1779 247 1780 251
rect 1774 246 1780 247
rect 1783 251 1789 252
rect 1783 247 1784 251
rect 1788 250 1789 251
rect 1878 251 1884 252
rect 1878 250 1879 251
rect 1788 248 1879 250
rect 1788 247 1789 248
rect 1783 246 1789 247
rect 1878 247 1879 248
rect 1883 247 1884 251
rect 1878 246 1884 247
rect 1887 251 1893 252
rect 1887 247 1888 251
rect 1892 250 1893 251
rect 1959 251 1965 252
rect 1959 250 1960 251
rect 1892 248 1960 250
rect 1892 247 1893 248
rect 1887 246 1893 247
rect 1959 247 1960 248
rect 1964 247 1965 251
rect 1959 246 1965 247
rect 1998 251 2005 252
rect 1998 247 1999 251
rect 2004 247 2005 251
rect 1998 246 2005 247
rect 2094 251 2101 252
rect 2094 247 2095 251
rect 2100 247 2101 251
rect 2094 246 2101 247
rect 110 244 116 245
rect 110 240 111 244
rect 115 240 116 244
rect 772 244 802 246
rect 1094 244 1100 245
rect 772 240 774 244
rect 1094 240 1095 244
rect 1099 240 1100 244
rect 110 239 116 240
rect 311 239 317 240
rect 311 235 312 239
rect 316 238 317 239
rect 334 239 340 240
rect 334 238 335 239
rect 316 236 335 238
rect 316 235 317 236
rect 311 234 317 235
rect 334 235 335 236
rect 339 235 340 239
rect 334 234 340 235
rect 342 239 348 240
rect 342 235 343 239
rect 347 238 348 239
rect 351 239 357 240
rect 351 238 352 239
rect 347 236 352 238
rect 347 235 348 236
rect 342 234 348 235
rect 351 235 352 236
rect 356 235 357 239
rect 351 234 357 235
rect 374 239 380 240
rect 374 235 375 239
rect 379 238 380 239
rect 391 239 397 240
rect 391 238 392 239
rect 379 236 392 238
rect 379 235 380 236
rect 374 234 380 235
rect 391 235 392 236
rect 396 235 397 239
rect 391 234 397 235
rect 430 239 436 240
rect 430 235 431 239
rect 435 238 436 239
rect 439 239 445 240
rect 439 238 440 239
rect 435 236 440 238
rect 435 235 436 236
rect 430 234 436 235
rect 439 235 440 236
rect 444 235 445 239
rect 439 234 445 235
rect 486 239 492 240
rect 486 235 487 239
rect 491 238 492 239
rect 495 239 501 240
rect 495 238 496 239
rect 491 236 496 238
rect 491 235 492 236
rect 486 234 492 235
rect 495 235 496 236
rect 500 235 501 239
rect 495 234 501 235
rect 550 239 556 240
rect 550 235 551 239
rect 555 238 556 239
rect 559 239 565 240
rect 559 238 560 239
rect 555 236 560 238
rect 555 235 556 236
rect 550 234 556 235
rect 559 235 560 236
rect 564 235 565 239
rect 559 234 565 235
rect 622 239 628 240
rect 622 235 623 239
rect 627 238 628 239
rect 631 239 637 240
rect 631 238 632 239
rect 627 236 632 238
rect 627 235 628 236
rect 622 234 628 235
rect 631 235 632 236
rect 636 235 637 239
rect 631 234 637 235
rect 703 239 712 240
rect 703 235 704 239
rect 711 235 712 239
rect 703 234 712 235
rect 767 239 774 240
rect 767 235 768 239
rect 772 236 774 239
rect 778 239 784 240
rect 772 235 773 236
rect 767 234 773 235
rect 778 235 779 239
rect 783 238 784 239
rect 831 239 837 240
rect 831 238 832 239
rect 783 236 832 238
rect 783 235 784 236
rect 778 234 784 235
rect 831 235 832 236
rect 836 235 837 239
rect 831 234 837 235
rect 886 239 893 240
rect 886 235 887 239
rect 892 235 893 239
rect 886 234 893 235
rect 942 239 948 240
rect 942 235 943 239
rect 947 238 948 239
rect 951 239 957 240
rect 951 238 952 239
rect 947 236 952 238
rect 947 235 948 236
rect 942 234 948 235
rect 951 235 952 236
rect 956 235 957 239
rect 951 234 957 235
rect 1006 239 1012 240
rect 1006 235 1007 239
rect 1011 238 1012 239
rect 1015 239 1021 240
rect 1015 238 1016 239
rect 1011 236 1016 238
rect 1011 235 1012 236
rect 1006 234 1012 235
rect 1015 235 1016 236
rect 1020 235 1021 239
rect 1015 234 1021 235
rect 1062 239 1068 240
rect 1062 235 1063 239
rect 1067 238 1068 239
rect 1071 239 1077 240
rect 1094 239 1100 240
rect 1262 244 1268 245
rect 1262 240 1263 244
rect 1267 240 1268 244
rect 1262 239 1268 240
rect 1302 244 1308 245
rect 1302 240 1303 244
rect 1307 240 1308 244
rect 1302 239 1308 240
rect 1342 244 1348 245
rect 1342 240 1343 244
rect 1347 240 1348 244
rect 1342 239 1348 240
rect 1382 244 1388 245
rect 1382 240 1383 244
rect 1387 240 1388 244
rect 1382 239 1388 240
rect 1422 244 1428 245
rect 1422 240 1423 244
rect 1427 240 1428 244
rect 1422 239 1428 240
rect 1462 244 1468 245
rect 1462 240 1463 244
rect 1467 240 1468 244
rect 1462 239 1468 240
rect 1502 244 1508 245
rect 1502 240 1503 244
rect 1507 240 1508 244
rect 1502 239 1508 240
rect 1542 244 1548 245
rect 1542 240 1543 244
rect 1547 240 1548 244
rect 1542 239 1548 240
rect 1598 244 1604 245
rect 1598 240 1599 244
rect 1603 240 1604 244
rect 1598 239 1604 240
rect 1670 244 1676 245
rect 1670 240 1671 244
rect 1675 240 1676 244
rect 1670 239 1676 240
rect 1758 244 1764 245
rect 1758 240 1759 244
rect 1763 240 1764 244
rect 1758 239 1764 240
rect 1862 244 1868 245
rect 1862 240 1863 244
rect 1867 240 1868 244
rect 1862 239 1868 240
rect 1974 244 1980 245
rect 1974 240 1975 244
rect 1979 240 1980 244
rect 1974 239 1980 240
rect 2070 244 2076 245
rect 2070 240 2071 244
rect 2075 240 2076 244
rect 2070 239 2076 240
rect 1071 238 1072 239
rect 1067 236 1072 238
rect 1067 235 1068 236
rect 1062 234 1068 235
rect 1071 235 1072 236
rect 1076 235 1077 239
rect 1071 234 1077 235
rect 1134 236 1140 237
rect 1134 232 1135 236
rect 1139 232 1140 236
rect 2118 236 2124 237
rect 2118 232 2119 236
rect 2123 232 2124 236
rect 1134 231 1140 232
rect 1287 231 1293 232
rect 110 227 116 228
rect 110 223 111 227
rect 115 223 116 227
rect 1094 227 1100 228
rect 110 222 116 223
rect 286 224 292 225
rect 286 220 287 224
rect 291 220 292 224
rect 286 219 292 220
rect 326 224 332 225
rect 326 220 327 224
rect 331 220 332 224
rect 326 219 332 220
rect 366 224 372 225
rect 366 220 367 224
rect 371 220 372 224
rect 366 219 372 220
rect 414 224 420 225
rect 414 220 415 224
rect 419 220 420 224
rect 414 219 420 220
rect 470 224 476 225
rect 470 220 471 224
rect 475 220 476 224
rect 470 219 476 220
rect 534 224 540 225
rect 534 220 535 224
rect 539 220 540 224
rect 534 219 540 220
rect 606 224 612 225
rect 606 220 607 224
rect 611 220 612 224
rect 606 219 612 220
rect 678 224 684 225
rect 678 220 679 224
rect 683 220 684 224
rect 678 219 684 220
rect 742 224 748 225
rect 742 220 743 224
rect 747 220 748 224
rect 742 219 748 220
rect 806 224 812 225
rect 806 220 807 224
rect 811 220 812 224
rect 806 219 812 220
rect 862 224 868 225
rect 862 220 863 224
rect 867 220 868 224
rect 862 219 868 220
rect 926 224 932 225
rect 926 220 927 224
rect 931 220 932 224
rect 926 219 932 220
rect 990 224 996 225
rect 990 220 991 224
rect 995 220 996 224
rect 990 219 996 220
rect 1046 224 1052 225
rect 1046 220 1047 224
rect 1051 220 1052 224
rect 1094 223 1095 227
rect 1099 223 1100 227
rect 1287 227 1288 231
rect 1292 230 1293 231
rect 1310 231 1316 232
rect 1310 230 1311 231
rect 1292 228 1311 230
rect 1292 227 1293 228
rect 1287 226 1293 227
rect 1310 227 1311 228
rect 1315 227 1316 231
rect 1310 226 1316 227
rect 1318 231 1324 232
rect 1318 227 1319 231
rect 1323 230 1324 231
rect 1327 231 1333 232
rect 1327 230 1328 231
rect 1323 228 1328 230
rect 1323 227 1324 228
rect 1318 226 1324 227
rect 1327 227 1328 228
rect 1332 227 1333 231
rect 1327 226 1333 227
rect 1358 231 1364 232
rect 1358 227 1359 231
rect 1363 230 1364 231
rect 1367 231 1373 232
rect 1367 230 1368 231
rect 1363 228 1368 230
rect 1363 227 1364 228
rect 1358 226 1364 227
rect 1367 227 1368 228
rect 1372 227 1373 231
rect 1367 226 1373 227
rect 1398 231 1404 232
rect 1398 227 1399 231
rect 1403 230 1404 231
rect 1407 231 1413 232
rect 1407 230 1408 231
rect 1403 228 1408 230
rect 1403 227 1404 228
rect 1398 226 1404 227
rect 1407 227 1408 228
rect 1412 227 1413 231
rect 1407 226 1413 227
rect 1438 231 1444 232
rect 1438 227 1439 231
rect 1443 230 1444 231
rect 1447 231 1453 232
rect 1447 230 1448 231
rect 1443 228 1448 230
rect 1443 227 1444 228
rect 1438 226 1444 227
rect 1447 227 1448 228
rect 1452 227 1453 231
rect 1447 226 1453 227
rect 1478 231 1484 232
rect 1478 227 1479 231
rect 1483 230 1484 231
rect 1487 231 1493 232
rect 1487 230 1488 231
rect 1483 228 1488 230
rect 1483 227 1484 228
rect 1478 226 1484 227
rect 1487 227 1488 228
rect 1492 227 1493 231
rect 1487 226 1493 227
rect 1518 231 1524 232
rect 1518 227 1519 231
rect 1523 230 1524 231
rect 1527 231 1533 232
rect 1527 230 1528 231
rect 1523 228 1528 230
rect 1523 227 1524 228
rect 1518 226 1524 227
rect 1527 227 1528 228
rect 1532 227 1533 231
rect 1527 226 1533 227
rect 1567 231 1576 232
rect 1567 227 1568 231
rect 1575 227 1576 231
rect 1567 226 1576 227
rect 1614 231 1620 232
rect 1614 227 1615 231
rect 1619 230 1620 231
rect 1623 231 1629 232
rect 1623 230 1624 231
rect 1619 228 1624 230
rect 1619 227 1620 228
rect 1614 226 1620 227
rect 1623 227 1624 228
rect 1628 227 1629 231
rect 1623 226 1629 227
rect 1686 231 1692 232
rect 1686 227 1687 231
rect 1691 230 1692 231
rect 1695 231 1701 232
rect 1695 230 1696 231
rect 1691 228 1696 230
rect 1691 227 1692 228
rect 1686 226 1692 227
rect 1695 227 1696 228
rect 1700 227 1701 231
rect 1695 226 1701 227
rect 1774 231 1780 232
rect 1774 227 1775 231
rect 1779 230 1780 231
rect 1783 231 1789 232
rect 1783 230 1784 231
rect 1779 228 1784 230
rect 1779 227 1780 228
rect 1774 226 1780 227
rect 1783 227 1784 228
rect 1788 227 1789 231
rect 1783 226 1789 227
rect 1878 231 1884 232
rect 1878 227 1879 231
rect 1883 230 1884 231
rect 1887 231 1893 232
rect 1887 230 1888 231
rect 1883 228 1888 230
rect 1883 227 1884 228
rect 1878 226 1884 227
rect 1887 227 1888 228
rect 1892 227 1893 231
rect 1887 226 1893 227
rect 1959 231 1965 232
rect 1959 227 1960 231
rect 1964 230 1965 231
rect 1999 231 2005 232
rect 1999 230 2000 231
rect 1964 228 2000 230
rect 1964 227 1965 228
rect 1959 226 1965 227
rect 1999 227 2000 228
rect 2004 227 2005 231
rect 1999 226 2005 227
rect 2062 231 2068 232
rect 2062 227 2063 231
rect 2067 230 2068 231
rect 2095 231 2101 232
rect 2118 231 2124 232
rect 2095 230 2096 231
rect 2067 228 2096 230
rect 2067 227 2068 228
rect 2062 226 2068 227
rect 2095 227 2096 228
rect 2100 227 2101 231
rect 2095 226 2101 227
rect 1094 222 1100 223
rect 1046 219 1052 220
rect 1134 219 1140 220
rect 1134 215 1135 219
rect 1139 215 1140 219
rect 2118 219 2124 220
rect 1134 214 1140 215
rect 1262 216 1268 217
rect 1262 212 1263 216
rect 1267 212 1268 216
rect 1262 211 1268 212
rect 1302 216 1308 217
rect 1302 212 1303 216
rect 1307 212 1308 216
rect 1302 211 1308 212
rect 1342 216 1348 217
rect 1342 212 1343 216
rect 1347 212 1348 216
rect 1342 211 1348 212
rect 1382 216 1388 217
rect 1382 212 1383 216
rect 1387 212 1388 216
rect 1382 211 1388 212
rect 1422 216 1428 217
rect 1422 212 1423 216
rect 1427 212 1428 216
rect 1422 211 1428 212
rect 1462 216 1468 217
rect 1462 212 1463 216
rect 1467 212 1468 216
rect 1462 211 1468 212
rect 1502 216 1508 217
rect 1502 212 1503 216
rect 1507 212 1508 216
rect 1502 211 1508 212
rect 1542 216 1548 217
rect 1542 212 1543 216
rect 1547 212 1548 216
rect 1542 211 1548 212
rect 1598 216 1604 217
rect 1598 212 1599 216
rect 1603 212 1604 216
rect 1598 211 1604 212
rect 1670 216 1676 217
rect 1670 212 1671 216
rect 1675 212 1676 216
rect 1670 211 1676 212
rect 1758 216 1764 217
rect 1758 212 1759 216
rect 1763 212 1764 216
rect 1758 211 1764 212
rect 1862 216 1868 217
rect 1862 212 1863 216
rect 1867 212 1868 216
rect 1862 211 1868 212
rect 1974 216 1980 217
rect 1974 212 1975 216
rect 1979 212 1980 216
rect 1974 211 1980 212
rect 2070 216 2076 217
rect 2070 212 2071 216
rect 2075 212 2076 216
rect 2118 215 2119 219
rect 2123 215 2124 219
rect 2118 214 2124 215
rect 2070 211 2076 212
rect 1614 207 1620 208
rect 1614 203 1615 207
rect 1619 206 1620 207
rect 1998 207 2004 208
rect 1998 206 1999 207
rect 1619 204 1999 206
rect 1619 203 1620 204
rect 1614 202 1620 203
rect 1998 203 1999 204
rect 2003 203 2004 207
rect 1998 202 2004 203
rect 166 200 172 201
rect 110 197 116 198
rect 110 193 111 197
rect 115 193 116 197
rect 166 196 167 200
rect 171 196 172 200
rect 166 195 172 196
rect 206 200 212 201
rect 206 196 207 200
rect 211 196 212 200
rect 206 195 212 196
rect 246 200 252 201
rect 246 196 247 200
rect 251 196 252 200
rect 246 195 252 196
rect 294 200 300 201
rect 294 196 295 200
rect 299 196 300 200
rect 294 195 300 196
rect 342 200 348 201
rect 342 196 343 200
rect 347 196 348 200
rect 342 195 348 196
rect 398 200 404 201
rect 398 196 399 200
rect 403 196 404 200
rect 398 195 404 196
rect 462 200 468 201
rect 462 196 463 200
rect 467 196 468 200
rect 462 195 468 196
rect 526 200 532 201
rect 526 196 527 200
rect 531 196 532 200
rect 526 195 532 196
rect 598 200 604 201
rect 598 196 599 200
rect 603 196 604 200
rect 598 195 604 196
rect 670 200 676 201
rect 670 196 671 200
rect 675 196 676 200
rect 670 195 676 196
rect 750 200 756 201
rect 750 196 751 200
rect 755 196 756 200
rect 750 195 756 196
rect 830 200 836 201
rect 830 196 831 200
rect 835 196 836 200
rect 830 195 836 196
rect 910 200 916 201
rect 910 196 911 200
rect 915 196 916 200
rect 910 195 916 196
rect 990 200 996 201
rect 990 196 991 200
rect 995 196 996 200
rect 990 195 996 196
rect 1046 200 1052 201
rect 1046 196 1047 200
rect 1051 196 1052 200
rect 1182 200 1188 201
rect 1046 195 1052 196
rect 1094 197 1100 198
rect 110 192 116 193
rect 1094 193 1095 197
rect 1099 193 1100 197
rect 1094 192 1100 193
rect 1134 197 1140 198
rect 1134 193 1135 197
rect 1139 193 1140 197
rect 1182 196 1183 200
rect 1187 196 1188 200
rect 1182 195 1188 196
rect 1230 200 1236 201
rect 1230 196 1231 200
rect 1235 196 1236 200
rect 1230 195 1236 196
rect 1294 200 1300 201
rect 1294 196 1295 200
rect 1299 196 1300 200
rect 1294 195 1300 196
rect 1358 200 1364 201
rect 1358 196 1359 200
rect 1363 196 1364 200
rect 1358 195 1364 196
rect 1430 200 1436 201
rect 1430 196 1431 200
rect 1435 196 1436 200
rect 1430 195 1436 196
rect 1510 200 1516 201
rect 1510 196 1511 200
rect 1515 196 1516 200
rect 1510 195 1516 196
rect 1590 200 1596 201
rect 1590 196 1591 200
rect 1595 196 1596 200
rect 1590 195 1596 196
rect 1662 200 1668 201
rect 1662 196 1663 200
rect 1667 196 1668 200
rect 1662 195 1668 196
rect 1734 200 1740 201
rect 1734 196 1735 200
rect 1739 196 1740 200
rect 1734 195 1740 196
rect 1806 200 1812 201
rect 1806 196 1807 200
rect 1811 196 1812 200
rect 1806 195 1812 196
rect 1878 200 1884 201
rect 1878 196 1879 200
rect 1883 196 1884 200
rect 1878 195 1884 196
rect 1950 200 1956 201
rect 1950 196 1951 200
rect 1955 196 1956 200
rect 1950 195 1956 196
rect 2022 200 2028 201
rect 2022 196 2023 200
rect 2027 196 2028 200
rect 2022 195 2028 196
rect 2070 200 2076 201
rect 2070 196 2071 200
rect 2075 196 2076 200
rect 2070 195 2076 196
rect 2118 197 2124 198
rect 1134 192 1140 193
rect 2118 193 2119 197
rect 2123 193 2124 197
rect 2118 192 2124 193
rect 1974 191 1980 192
rect 1974 190 1975 191
rect 1904 188 1975 190
rect 1904 184 1906 188
rect 1974 187 1975 188
rect 1979 187 1980 191
rect 1974 186 1980 187
rect 191 183 200 184
rect 110 180 116 181
rect 110 176 111 180
rect 115 176 116 180
rect 191 179 192 183
rect 199 179 200 183
rect 191 178 200 179
rect 214 183 220 184
rect 214 179 215 183
rect 219 182 220 183
rect 231 183 237 184
rect 231 182 232 183
rect 219 180 232 182
rect 219 179 220 180
rect 214 178 220 179
rect 231 179 232 180
rect 236 179 237 183
rect 231 178 237 179
rect 254 183 260 184
rect 254 179 255 183
rect 259 182 260 183
rect 271 183 277 184
rect 271 182 272 183
rect 259 180 272 182
rect 259 179 260 180
rect 254 178 260 179
rect 271 179 272 180
rect 276 179 277 183
rect 271 178 277 179
rect 279 183 285 184
rect 279 179 280 183
rect 284 182 285 183
rect 319 183 325 184
rect 319 182 320 183
rect 284 180 320 182
rect 284 179 285 180
rect 279 178 285 179
rect 319 179 320 180
rect 324 179 325 183
rect 319 178 325 179
rect 327 183 333 184
rect 327 179 328 183
rect 332 182 333 183
rect 367 183 373 184
rect 367 182 368 183
rect 332 180 368 182
rect 332 179 333 180
rect 327 178 333 179
rect 367 179 368 180
rect 372 179 373 183
rect 367 178 373 179
rect 375 183 381 184
rect 375 179 376 183
rect 380 182 381 183
rect 423 183 429 184
rect 423 182 424 183
rect 380 180 424 182
rect 380 179 381 180
rect 375 178 381 179
rect 423 179 424 180
rect 428 179 429 183
rect 423 178 429 179
rect 431 183 437 184
rect 431 179 432 183
rect 436 182 437 183
rect 487 183 493 184
rect 487 182 488 183
rect 436 180 488 182
rect 436 179 437 180
rect 431 178 437 179
rect 487 179 488 180
rect 492 179 493 183
rect 487 178 493 179
rect 551 183 557 184
rect 551 179 552 183
rect 556 182 557 183
rect 614 183 620 184
rect 614 182 615 183
rect 556 180 615 182
rect 556 179 557 180
rect 551 178 557 179
rect 614 179 615 180
rect 619 179 620 183
rect 614 178 620 179
rect 623 183 629 184
rect 623 179 624 183
rect 628 182 629 183
rect 678 183 684 184
rect 678 182 679 183
rect 628 180 679 182
rect 628 179 629 180
rect 623 178 629 179
rect 678 179 679 180
rect 683 179 684 183
rect 678 178 684 179
rect 695 183 704 184
rect 695 179 696 183
rect 703 179 704 183
rect 695 178 704 179
rect 775 183 781 184
rect 775 179 776 183
rect 780 182 781 183
rect 846 183 852 184
rect 846 182 847 183
rect 780 180 847 182
rect 780 179 781 180
rect 775 178 781 179
rect 846 179 847 180
rect 851 179 852 183
rect 846 178 852 179
rect 855 183 861 184
rect 855 179 856 183
rect 860 182 861 183
rect 926 183 932 184
rect 926 182 927 183
rect 860 180 927 182
rect 860 179 861 180
rect 855 178 861 179
rect 926 179 927 180
rect 931 179 932 183
rect 926 178 932 179
rect 935 183 941 184
rect 935 179 936 183
rect 940 182 941 183
rect 958 183 964 184
rect 958 182 959 183
rect 940 180 959 182
rect 940 179 941 180
rect 935 178 941 179
rect 958 179 959 180
rect 963 179 964 183
rect 958 178 964 179
rect 1015 183 1021 184
rect 1015 179 1016 183
rect 1020 182 1021 183
rect 1062 183 1068 184
rect 1062 182 1063 183
rect 1020 180 1063 182
rect 1020 179 1021 180
rect 1015 178 1021 179
rect 1062 179 1063 180
rect 1067 179 1068 183
rect 1062 178 1068 179
rect 1070 183 1077 184
rect 1070 179 1071 183
rect 1076 179 1077 183
rect 1207 183 1216 184
rect 1070 178 1077 179
rect 1094 180 1100 181
rect 110 175 116 176
rect 1094 176 1095 180
rect 1099 176 1100 180
rect 1094 175 1100 176
rect 1134 180 1140 181
rect 1134 176 1135 180
rect 1139 176 1140 180
rect 1207 179 1208 183
rect 1215 179 1216 183
rect 1207 178 1216 179
rect 1218 183 1224 184
rect 1218 179 1219 183
rect 1223 182 1224 183
rect 1255 183 1261 184
rect 1255 182 1256 183
rect 1223 180 1256 182
rect 1223 179 1224 180
rect 1218 178 1224 179
rect 1255 179 1256 180
rect 1260 179 1261 183
rect 1255 178 1261 179
rect 1263 183 1269 184
rect 1263 179 1264 183
rect 1268 182 1269 183
rect 1319 183 1325 184
rect 1319 182 1320 183
rect 1268 180 1320 182
rect 1268 179 1269 180
rect 1263 178 1269 179
rect 1319 179 1320 180
rect 1324 179 1325 183
rect 1319 178 1325 179
rect 1327 183 1333 184
rect 1327 179 1328 183
rect 1332 182 1333 183
rect 1383 183 1389 184
rect 1383 182 1384 183
rect 1332 180 1384 182
rect 1332 179 1333 180
rect 1327 178 1333 179
rect 1383 179 1384 180
rect 1388 179 1389 183
rect 1383 178 1389 179
rect 1391 183 1397 184
rect 1391 179 1392 183
rect 1396 182 1397 183
rect 1455 183 1461 184
rect 1455 182 1456 183
rect 1396 180 1456 182
rect 1396 179 1397 180
rect 1391 178 1397 179
rect 1455 179 1456 180
rect 1460 179 1461 183
rect 1455 178 1461 179
rect 1463 183 1469 184
rect 1463 179 1464 183
rect 1468 182 1469 183
rect 1535 183 1541 184
rect 1535 182 1536 183
rect 1468 180 1536 182
rect 1468 179 1469 180
rect 1463 178 1469 179
rect 1535 179 1536 180
rect 1540 179 1541 183
rect 1535 178 1541 179
rect 1614 183 1621 184
rect 1614 179 1615 183
rect 1620 179 1621 183
rect 1614 178 1621 179
rect 1623 183 1629 184
rect 1623 179 1624 183
rect 1628 182 1629 183
rect 1687 183 1693 184
rect 1687 182 1688 183
rect 1628 180 1688 182
rect 1628 179 1629 180
rect 1623 178 1629 179
rect 1687 179 1688 180
rect 1692 179 1693 183
rect 1687 178 1693 179
rect 1695 183 1701 184
rect 1695 179 1696 183
rect 1700 182 1701 183
rect 1759 183 1765 184
rect 1759 182 1760 183
rect 1700 180 1760 182
rect 1700 179 1701 180
rect 1695 178 1701 179
rect 1759 179 1760 180
rect 1764 179 1765 183
rect 1759 178 1765 179
rect 1767 183 1773 184
rect 1767 179 1768 183
rect 1772 182 1773 183
rect 1831 183 1837 184
rect 1831 182 1832 183
rect 1772 180 1832 182
rect 1772 179 1773 180
rect 1767 178 1773 179
rect 1831 179 1832 180
rect 1836 179 1837 183
rect 1831 178 1837 179
rect 1903 183 1909 184
rect 1903 179 1904 183
rect 1908 179 1909 183
rect 1903 178 1909 179
rect 1911 183 1917 184
rect 1911 179 1912 183
rect 1916 182 1917 183
rect 1975 183 1981 184
rect 1975 182 1976 183
rect 1916 180 1976 182
rect 1916 179 1917 180
rect 1911 178 1917 179
rect 1975 179 1976 180
rect 1980 179 1981 183
rect 1975 178 1981 179
rect 2047 183 2053 184
rect 2047 179 2048 183
rect 2052 182 2053 183
rect 2086 183 2092 184
rect 2086 182 2087 183
rect 2052 180 2087 182
rect 2052 179 2053 180
rect 2047 178 2053 179
rect 2086 179 2087 180
rect 2091 179 2092 183
rect 2086 178 2092 179
rect 2094 183 2101 184
rect 2094 179 2095 183
rect 2100 179 2101 183
rect 2094 178 2101 179
rect 2118 180 2124 181
rect 1134 175 1140 176
rect 2118 176 2119 180
rect 2123 176 2124 180
rect 2118 175 2124 176
rect 166 172 172 173
rect 166 168 167 172
rect 171 168 172 172
rect 166 167 172 168
rect 206 172 212 173
rect 206 168 207 172
rect 211 168 212 172
rect 206 167 212 168
rect 246 172 252 173
rect 246 168 247 172
rect 251 168 252 172
rect 246 167 252 168
rect 294 172 300 173
rect 294 168 295 172
rect 299 168 300 172
rect 294 167 300 168
rect 342 172 348 173
rect 342 168 343 172
rect 347 168 348 172
rect 342 167 348 168
rect 398 172 404 173
rect 398 168 399 172
rect 403 168 404 172
rect 398 167 404 168
rect 462 172 468 173
rect 462 168 463 172
rect 467 168 468 172
rect 462 167 468 168
rect 526 172 532 173
rect 526 168 527 172
rect 531 168 532 172
rect 526 167 532 168
rect 598 172 604 173
rect 598 168 599 172
rect 603 168 604 172
rect 598 167 604 168
rect 670 172 676 173
rect 670 168 671 172
rect 675 168 676 172
rect 670 167 676 168
rect 750 172 756 173
rect 750 168 751 172
rect 755 168 756 172
rect 750 167 756 168
rect 830 172 836 173
rect 830 168 831 172
rect 835 168 836 172
rect 830 167 836 168
rect 910 172 916 173
rect 910 168 911 172
rect 915 168 916 172
rect 910 167 916 168
rect 990 172 996 173
rect 990 168 991 172
rect 995 168 996 172
rect 990 167 996 168
rect 1046 172 1052 173
rect 1046 168 1047 172
rect 1051 168 1052 172
rect 1046 167 1052 168
rect 1182 172 1188 173
rect 1182 168 1183 172
rect 1187 168 1188 172
rect 1182 167 1188 168
rect 1230 172 1236 173
rect 1230 168 1231 172
rect 1235 168 1236 172
rect 1230 167 1236 168
rect 1294 172 1300 173
rect 1294 168 1295 172
rect 1299 168 1300 172
rect 1294 167 1300 168
rect 1358 172 1364 173
rect 1358 168 1359 172
rect 1363 168 1364 172
rect 1358 167 1364 168
rect 1430 172 1436 173
rect 1430 168 1431 172
rect 1435 168 1436 172
rect 1430 167 1436 168
rect 1510 172 1516 173
rect 1510 168 1511 172
rect 1515 168 1516 172
rect 1510 167 1516 168
rect 1590 172 1596 173
rect 1590 168 1591 172
rect 1595 168 1596 172
rect 1590 167 1596 168
rect 1662 172 1668 173
rect 1662 168 1663 172
rect 1667 168 1668 172
rect 1662 167 1668 168
rect 1734 172 1740 173
rect 1734 168 1735 172
rect 1739 168 1740 172
rect 1734 167 1740 168
rect 1806 172 1812 173
rect 1806 168 1807 172
rect 1811 168 1812 172
rect 1806 167 1812 168
rect 1878 172 1884 173
rect 1878 168 1879 172
rect 1883 168 1884 172
rect 1878 167 1884 168
rect 1950 172 1956 173
rect 1950 168 1951 172
rect 1955 168 1956 172
rect 1950 167 1956 168
rect 2022 172 2028 173
rect 2022 168 2023 172
rect 2027 168 2028 172
rect 2022 167 2028 168
rect 2070 172 2076 173
rect 2070 168 2071 172
rect 2075 168 2076 172
rect 2070 167 2076 168
rect 191 163 197 164
rect 191 159 192 163
rect 196 162 197 163
rect 214 163 220 164
rect 214 162 215 163
rect 196 160 215 162
rect 196 159 197 160
rect 191 158 197 159
rect 214 159 215 160
rect 219 159 220 163
rect 214 158 220 159
rect 231 163 237 164
rect 231 159 232 163
rect 236 162 237 163
rect 254 163 260 164
rect 254 162 255 163
rect 236 160 255 162
rect 236 159 237 160
rect 231 158 237 159
rect 254 159 255 160
rect 259 159 260 163
rect 254 158 260 159
rect 271 163 277 164
rect 271 159 272 163
rect 276 162 277 163
rect 279 163 285 164
rect 279 162 280 163
rect 276 160 280 162
rect 276 159 277 160
rect 271 158 277 159
rect 279 159 280 160
rect 284 159 285 163
rect 279 158 285 159
rect 319 163 325 164
rect 319 159 320 163
rect 324 162 325 163
rect 327 163 333 164
rect 327 162 328 163
rect 324 160 328 162
rect 324 159 325 160
rect 319 158 325 159
rect 327 159 328 160
rect 332 159 333 163
rect 327 158 333 159
rect 367 163 373 164
rect 367 159 368 163
rect 372 162 373 163
rect 375 163 381 164
rect 375 162 376 163
rect 372 160 376 162
rect 372 159 373 160
rect 367 158 373 159
rect 375 159 376 160
rect 380 159 381 163
rect 375 158 381 159
rect 423 163 429 164
rect 423 159 424 163
rect 428 162 429 163
rect 431 163 437 164
rect 431 162 432 163
rect 428 160 432 162
rect 428 159 429 160
rect 423 158 429 159
rect 431 159 432 160
rect 436 159 437 163
rect 487 163 493 164
rect 487 162 488 163
rect 431 158 437 159
rect 440 160 488 162
rect 334 155 340 156
rect 334 151 335 155
rect 339 154 340 155
rect 440 154 442 160
rect 487 159 488 160
rect 492 159 493 163
rect 487 158 493 159
rect 551 163 560 164
rect 551 159 552 163
rect 559 159 560 163
rect 551 158 560 159
rect 614 163 620 164
rect 614 159 615 163
rect 619 162 620 163
rect 623 163 629 164
rect 623 162 624 163
rect 619 160 624 162
rect 619 159 620 160
rect 614 158 620 159
rect 623 159 624 160
rect 628 159 629 163
rect 623 158 629 159
rect 678 163 684 164
rect 678 159 679 163
rect 683 162 684 163
rect 695 163 701 164
rect 695 162 696 163
rect 683 160 696 162
rect 683 159 684 160
rect 678 158 684 159
rect 695 159 696 160
rect 700 159 701 163
rect 695 158 701 159
rect 775 163 784 164
rect 775 159 776 163
rect 783 159 784 163
rect 775 158 784 159
rect 846 163 852 164
rect 846 159 847 163
rect 851 162 852 163
rect 855 163 861 164
rect 855 162 856 163
rect 851 160 856 162
rect 851 159 852 160
rect 846 158 852 159
rect 855 159 856 160
rect 860 159 861 163
rect 855 158 861 159
rect 926 163 932 164
rect 926 159 927 163
rect 931 162 932 163
rect 935 163 941 164
rect 935 162 936 163
rect 931 160 936 162
rect 931 159 932 160
rect 926 158 932 159
rect 935 159 936 160
rect 940 159 941 163
rect 935 158 941 159
rect 1015 163 1024 164
rect 1015 159 1016 163
rect 1023 159 1024 163
rect 1015 158 1024 159
rect 1062 163 1068 164
rect 1062 159 1063 163
rect 1067 162 1068 163
rect 1071 163 1077 164
rect 1071 162 1072 163
rect 1067 160 1072 162
rect 1067 159 1068 160
rect 1062 158 1068 159
rect 1071 159 1072 160
rect 1076 159 1077 163
rect 1071 158 1077 159
rect 1207 163 1213 164
rect 1207 159 1208 163
rect 1212 162 1213 163
rect 1218 163 1224 164
rect 1218 162 1219 163
rect 1212 160 1219 162
rect 1212 159 1213 160
rect 1207 158 1213 159
rect 1218 159 1219 160
rect 1223 159 1224 163
rect 1218 158 1224 159
rect 1255 163 1261 164
rect 1255 159 1256 163
rect 1260 162 1261 163
rect 1263 163 1269 164
rect 1263 162 1264 163
rect 1260 160 1264 162
rect 1260 159 1261 160
rect 1255 158 1261 159
rect 1263 159 1264 160
rect 1268 159 1269 163
rect 1263 158 1269 159
rect 1319 163 1325 164
rect 1319 159 1320 163
rect 1324 162 1325 163
rect 1327 163 1333 164
rect 1327 162 1328 163
rect 1324 160 1328 162
rect 1324 159 1325 160
rect 1319 158 1325 159
rect 1327 159 1328 160
rect 1332 159 1333 163
rect 1327 158 1333 159
rect 1383 163 1389 164
rect 1383 159 1384 163
rect 1388 162 1389 163
rect 1391 163 1397 164
rect 1391 162 1392 163
rect 1388 160 1392 162
rect 1388 159 1389 160
rect 1383 158 1389 159
rect 1391 159 1392 160
rect 1396 159 1397 163
rect 1391 158 1397 159
rect 1455 163 1461 164
rect 1455 159 1456 163
rect 1460 162 1461 163
rect 1463 163 1469 164
rect 1463 162 1464 163
rect 1460 160 1464 162
rect 1460 159 1461 160
rect 1455 158 1461 159
rect 1463 159 1464 160
rect 1468 159 1469 163
rect 1535 163 1541 164
rect 1535 162 1536 163
rect 1463 158 1469 159
rect 1472 160 1536 162
rect 339 152 442 154
rect 1310 155 1316 156
rect 339 151 340 152
rect 334 150 340 151
rect 1310 151 1311 155
rect 1315 154 1316 155
rect 1472 154 1474 160
rect 1535 159 1536 160
rect 1540 159 1541 163
rect 1535 158 1541 159
rect 1615 163 1621 164
rect 1615 159 1616 163
rect 1620 162 1621 163
rect 1623 163 1629 164
rect 1623 162 1624 163
rect 1620 160 1624 162
rect 1620 159 1621 160
rect 1615 158 1621 159
rect 1623 159 1624 160
rect 1628 159 1629 163
rect 1623 158 1629 159
rect 1687 163 1693 164
rect 1687 159 1688 163
rect 1692 162 1693 163
rect 1695 163 1701 164
rect 1695 162 1696 163
rect 1692 160 1696 162
rect 1692 159 1693 160
rect 1687 158 1693 159
rect 1695 159 1696 160
rect 1700 159 1701 163
rect 1695 158 1701 159
rect 1759 163 1765 164
rect 1759 159 1760 163
rect 1764 162 1765 163
rect 1767 163 1773 164
rect 1767 162 1768 163
rect 1764 160 1768 162
rect 1764 159 1765 160
rect 1759 158 1765 159
rect 1767 159 1768 160
rect 1772 159 1773 163
rect 1831 163 1837 164
rect 1831 162 1832 163
rect 1767 158 1773 159
rect 1776 160 1832 162
rect 1315 152 1474 154
rect 1598 155 1604 156
rect 1315 151 1316 152
rect 1310 150 1316 151
rect 1598 151 1599 155
rect 1603 154 1604 155
rect 1776 154 1778 160
rect 1831 159 1832 160
rect 1836 159 1837 163
rect 1831 158 1837 159
rect 1903 163 1909 164
rect 1903 159 1904 163
rect 1908 162 1909 163
rect 1911 163 1917 164
rect 1911 162 1912 163
rect 1908 160 1912 162
rect 1908 159 1909 160
rect 1903 158 1909 159
rect 1911 159 1912 160
rect 1916 159 1917 163
rect 1911 158 1917 159
rect 1975 163 1981 164
rect 1975 159 1976 163
rect 1980 162 1981 163
rect 2014 163 2020 164
rect 2014 162 2015 163
rect 1980 160 2015 162
rect 1980 159 1981 160
rect 1975 158 1981 159
rect 2014 159 2015 160
rect 2019 159 2020 163
rect 2014 158 2020 159
rect 2047 163 2053 164
rect 2047 159 2048 163
rect 2052 162 2053 163
rect 2062 163 2068 164
rect 2062 162 2063 163
rect 2052 160 2063 162
rect 2052 159 2053 160
rect 2047 158 2053 159
rect 2062 159 2063 160
rect 2067 159 2068 163
rect 2062 158 2068 159
rect 2086 163 2092 164
rect 2086 159 2087 163
rect 2091 162 2092 163
rect 2095 163 2101 164
rect 2095 162 2096 163
rect 2091 160 2096 162
rect 2091 159 2092 160
rect 2086 158 2092 159
rect 2095 159 2096 160
rect 2100 159 2101 163
rect 2095 158 2101 159
rect 1603 152 1778 154
rect 1603 151 1604 152
rect 1598 150 1604 151
rect 194 135 200 136
rect 194 131 195 135
rect 199 134 200 135
rect 199 132 522 134
rect 199 131 200 132
rect 194 130 200 131
rect 520 128 522 132
rect 159 127 165 128
rect 159 123 160 127
rect 164 126 165 127
rect 190 127 196 128
rect 190 126 191 127
rect 164 124 191 126
rect 164 123 165 124
rect 159 122 165 123
rect 190 123 191 124
rect 195 123 196 127
rect 190 122 196 123
rect 199 127 205 128
rect 199 123 200 127
rect 204 126 205 127
rect 230 127 236 128
rect 230 126 231 127
rect 204 124 231 126
rect 204 123 205 124
rect 199 122 205 123
rect 230 123 231 124
rect 235 123 236 127
rect 230 122 236 123
rect 239 127 245 128
rect 239 123 240 127
rect 244 126 245 127
rect 270 127 276 128
rect 270 126 271 127
rect 244 124 271 126
rect 244 123 245 124
rect 239 122 245 123
rect 270 123 271 124
rect 275 123 276 127
rect 270 122 276 123
rect 279 127 285 128
rect 279 123 280 127
rect 284 126 285 127
rect 302 127 308 128
rect 302 126 303 127
rect 284 124 303 126
rect 284 123 285 124
rect 279 122 285 123
rect 302 123 303 124
rect 307 123 308 127
rect 302 122 308 123
rect 319 127 325 128
rect 319 123 320 127
rect 324 126 325 127
rect 350 127 356 128
rect 350 126 351 127
rect 324 124 351 126
rect 324 123 325 124
rect 319 122 325 123
rect 350 123 351 124
rect 355 123 356 127
rect 350 122 356 123
rect 359 127 365 128
rect 359 123 360 127
rect 364 126 365 127
rect 390 127 396 128
rect 390 126 391 127
rect 364 124 391 126
rect 364 123 365 124
rect 359 122 365 123
rect 390 123 391 124
rect 395 123 396 127
rect 390 122 396 123
rect 399 127 405 128
rect 399 123 400 127
rect 404 126 405 127
rect 430 127 436 128
rect 430 126 431 127
rect 404 124 431 126
rect 404 123 405 124
rect 399 122 405 123
rect 430 123 431 124
rect 435 123 436 127
rect 430 122 436 123
rect 439 127 445 128
rect 439 123 440 127
rect 444 126 445 127
rect 470 127 476 128
rect 470 126 471 127
rect 444 124 471 126
rect 444 123 445 124
rect 439 122 445 123
rect 470 123 471 124
rect 475 123 476 127
rect 470 122 476 123
rect 479 127 485 128
rect 479 123 480 127
rect 484 126 485 127
rect 510 127 516 128
rect 510 126 511 127
rect 484 124 511 126
rect 484 123 485 124
rect 479 122 485 123
rect 510 123 511 124
rect 515 123 516 127
rect 510 122 516 123
rect 519 127 525 128
rect 519 123 520 127
rect 524 123 525 127
rect 519 122 525 123
rect 559 127 565 128
rect 559 123 560 127
rect 564 126 565 127
rect 590 127 596 128
rect 590 126 591 127
rect 564 124 591 126
rect 564 123 565 124
rect 559 122 565 123
rect 590 123 591 124
rect 595 123 596 127
rect 590 122 596 123
rect 599 127 605 128
rect 599 123 600 127
rect 604 126 605 127
rect 630 127 636 128
rect 630 126 631 127
rect 604 124 631 126
rect 604 123 605 124
rect 599 122 605 123
rect 630 123 631 124
rect 635 123 636 127
rect 630 122 636 123
rect 639 127 645 128
rect 639 123 640 127
rect 644 126 645 127
rect 670 127 676 128
rect 670 126 671 127
rect 644 124 671 126
rect 644 123 645 124
rect 639 122 645 123
rect 670 123 671 124
rect 675 123 676 127
rect 670 122 676 123
rect 679 127 685 128
rect 679 123 680 127
rect 684 126 685 127
rect 710 127 716 128
rect 710 126 711 127
rect 684 124 711 126
rect 684 123 685 124
rect 679 122 685 123
rect 710 123 711 124
rect 715 123 716 127
rect 710 122 716 123
rect 719 127 725 128
rect 719 123 720 127
rect 724 126 725 127
rect 750 127 756 128
rect 750 126 751 127
rect 724 124 751 126
rect 724 123 725 124
rect 719 122 725 123
rect 750 123 751 124
rect 755 123 756 127
rect 750 122 756 123
rect 759 127 765 128
rect 759 123 760 127
rect 764 126 765 127
rect 790 127 796 128
rect 790 126 791 127
rect 764 124 791 126
rect 764 123 765 124
rect 759 122 765 123
rect 790 123 791 124
rect 795 123 796 127
rect 790 122 796 123
rect 799 127 805 128
rect 799 123 800 127
rect 804 126 805 127
rect 830 127 836 128
rect 830 126 831 127
rect 804 124 831 126
rect 804 123 805 124
rect 799 122 805 123
rect 830 123 831 124
rect 835 123 836 127
rect 830 122 836 123
rect 839 127 845 128
rect 839 123 840 127
rect 844 126 845 127
rect 886 127 892 128
rect 886 126 887 127
rect 844 124 887 126
rect 844 123 845 124
rect 839 122 845 123
rect 886 123 887 124
rect 891 123 892 127
rect 886 122 892 123
rect 895 127 901 128
rect 895 123 896 127
rect 900 126 901 127
rect 942 127 948 128
rect 942 126 943 127
rect 900 124 943 126
rect 900 123 901 124
rect 895 122 901 123
rect 942 123 943 124
rect 947 123 948 127
rect 942 122 948 123
rect 958 127 965 128
rect 958 123 959 127
rect 964 123 965 127
rect 958 122 965 123
rect 1023 127 1029 128
rect 1023 123 1024 127
rect 1028 126 1029 127
rect 1062 127 1068 128
rect 1062 126 1063 127
rect 1028 124 1063 126
rect 1028 123 1029 124
rect 1023 122 1029 123
rect 1062 123 1063 124
rect 1067 123 1068 127
rect 1062 122 1068 123
rect 1071 127 1077 128
rect 1071 123 1072 127
rect 1076 126 1077 127
rect 1174 127 1180 128
rect 1174 126 1175 127
rect 1076 124 1175 126
rect 1076 123 1077 124
rect 1071 122 1077 123
rect 1174 123 1175 124
rect 1179 123 1180 127
rect 1174 122 1180 123
rect 1210 127 1216 128
rect 1210 123 1211 127
rect 1215 126 1216 127
rect 1215 124 1514 126
rect 1215 123 1216 124
rect 1210 122 1216 123
rect 134 120 140 121
rect 134 116 135 120
rect 139 116 140 120
rect 134 115 140 116
rect 174 120 180 121
rect 174 116 175 120
rect 179 116 180 120
rect 174 115 180 116
rect 214 120 220 121
rect 214 116 215 120
rect 219 116 220 120
rect 214 115 220 116
rect 254 120 260 121
rect 254 116 255 120
rect 259 116 260 120
rect 254 115 260 116
rect 294 120 300 121
rect 294 116 295 120
rect 299 116 300 120
rect 294 115 300 116
rect 334 120 340 121
rect 334 116 335 120
rect 339 116 340 120
rect 334 115 340 116
rect 374 120 380 121
rect 374 116 375 120
rect 379 116 380 120
rect 374 115 380 116
rect 414 120 420 121
rect 414 116 415 120
rect 419 116 420 120
rect 414 115 420 116
rect 454 120 460 121
rect 454 116 455 120
rect 459 116 460 120
rect 454 115 460 116
rect 494 120 500 121
rect 494 116 495 120
rect 499 116 500 120
rect 494 115 500 116
rect 534 120 540 121
rect 534 116 535 120
rect 539 116 540 120
rect 534 115 540 116
rect 574 120 580 121
rect 574 116 575 120
rect 579 116 580 120
rect 574 115 580 116
rect 614 120 620 121
rect 614 116 615 120
rect 619 116 620 120
rect 614 115 620 116
rect 654 120 660 121
rect 654 116 655 120
rect 659 116 660 120
rect 654 115 660 116
rect 694 120 700 121
rect 694 116 695 120
rect 699 116 700 120
rect 694 115 700 116
rect 734 120 740 121
rect 734 116 735 120
rect 739 116 740 120
rect 734 115 740 116
rect 774 120 780 121
rect 774 116 775 120
rect 779 116 780 120
rect 774 115 780 116
rect 814 120 820 121
rect 814 116 815 120
rect 819 116 820 120
rect 814 115 820 116
rect 870 120 876 121
rect 870 116 871 120
rect 875 116 876 120
rect 870 115 876 116
rect 934 120 940 121
rect 934 116 935 120
rect 939 116 940 120
rect 934 115 940 116
rect 998 120 1004 121
rect 998 116 999 120
rect 1003 116 1004 120
rect 998 115 1004 116
rect 1046 120 1052 121
rect 1046 116 1047 120
rect 1051 116 1052 120
rect 1046 115 1052 116
rect 1183 119 1189 120
rect 1183 115 1184 119
rect 1188 118 1189 119
rect 1214 119 1220 120
rect 1214 118 1215 119
rect 1188 116 1215 118
rect 1188 115 1189 116
rect 1183 114 1189 115
rect 1214 115 1215 116
rect 1219 115 1220 119
rect 1214 114 1220 115
rect 1223 119 1229 120
rect 1223 115 1224 119
rect 1228 118 1229 119
rect 1254 119 1260 120
rect 1254 118 1255 119
rect 1228 116 1255 118
rect 1228 115 1229 116
rect 1223 114 1229 115
rect 1254 115 1255 116
rect 1259 115 1260 119
rect 1254 114 1260 115
rect 1263 119 1269 120
rect 1263 115 1264 119
rect 1268 118 1269 119
rect 1294 119 1300 120
rect 1294 118 1295 119
rect 1268 116 1295 118
rect 1268 115 1269 116
rect 1263 114 1269 115
rect 1294 115 1295 116
rect 1299 115 1300 119
rect 1294 114 1300 115
rect 1303 119 1309 120
rect 1303 115 1304 119
rect 1308 118 1309 119
rect 1334 119 1340 120
rect 1334 118 1335 119
rect 1308 116 1335 118
rect 1308 115 1309 116
rect 1303 114 1309 115
rect 1334 115 1335 116
rect 1339 115 1340 119
rect 1334 114 1340 115
rect 1343 119 1349 120
rect 1343 115 1344 119
rect 1348 118 1349 119
rect 1382 119 1388 120
rect 1382 118 1383 119
rect 1348 116 1383 118
rect 1348 115 1349 116
rect 1343 114 1349 115
rect 1382 115 1383 116
rect 1387 115 1388 119
rect 1382 114 1388 115
rect 1391 119 1397 120
rect 1391 115 1392 119
rect 1396 118 1397 119
rect 1446 119 1452 120
rect 1446 118 1447 119
rect 1396 116 1447 118
rect 1396 115 1397 116
rect 1391 114 1397 115
rect 1446 115 1447 116
rect 1451 115 1452 119
rect 1446 114 1452 115
rect 1455 119 1461 120
rect 1455 115 1456 119
rect 1460 118 1461 119
rect 1502 119 1508 120
rect 1502 118 1503 119
rect 1460 116 1503 118
rect 1460 115 1461 116
rect 1455 114 1461 115
rect 1502 115 1503 116
rect 1507 115 1508 119
rect 1512 118 1514 124
rect 1519 119 1525 120
rect 1519 118 1520 119
rect 1512 116 1520 118
rect 1502 114 1508 115
rect 1519 115 1520 116
rect 1524 115 1525 119
rect 1519 114 1525 115
rect 1583 119 1589 120
rect 1583 115 1584 119
rect 1588 118 1589 119
rect 1630 119 1636 120
rect 1630 118 1631 119
rect 1588 116 1631 118
rect 1588 115 1589 116
rect 1583 114 1589 115
rect 1630 115 1631 116
rect 1635 115 1636 119
rect 1630 114 1636 115
rect 1639 119 1645 120
rect 1639 115 1640 119
rect 1644 118 1645 119
rect 1686 119 1692 120
rect 1686 118 1687 119
rect 1644 116 1687 118
rect 1644 115 1645 116
rect 1639 114 1645 115
rect 1686 115 1687 116
rect 1691 115 1692 119
rect 1686 114 1692 115
rect 1695 119 1701 120
rect 1695 115 1696 119
rect 1700 118 1701 119
rect 1734 119 1740 120
rect 1734 118 1735 119
rect 1700 116 1735 118
rect 1700 115 1701 116
rect 1695 114 1701 115
rect 1734 115 1735 116
rect 1739 115 1740 119
rect 1734 114 1740 115
rect 1743 119 1749 120
rect 1743 115 1744 119
rect 1748 118 1749 119
rect 1782 119 1788 120
rect 1782 118 1783 119
rect 1748 116 1783 118
rect 1748 115 1749 116
rect 1743 114 1749 115
rect 1782 115 1783 116
rect 1787 115 1788 119
rect 1782 114 1788 115
rect 1791 119 1797 120
rect 1791 115 1792 119
rect 1796 118 1797 119
rect 1822 119 1828 120
rect 1822 118 1823 119
rect 1796 116 1823 118
rect 1796 115 1797 116
rect 1791 114 1797 115
rect 1822 115 1823 116
rect 1827 115 1828 119
rect 1822 114 1828 115
rect 1831 119 1837 120
rect 1831 115 1832 119
rect 1836 118 1837 119
rect 1870 119 1876 120
rect 1870 118 1871 119
rect 1836 116 1871 118
rect 1836 115 1837 116
rect 1831 114 1837 115
rect 1870 115 1871 116
rect 1875 115 1876 119
rect 1870 114 1876 115
rect 1879 119 1885 120
rect 1879 115 1880 119
rect 1884 118 1885 119
rect 1918 119 1924 120
rect 1918 118 1919 119
rect 1884 116 1919 118
rect 1884 115 1885 116
rect 1879 114 1885 115
rect 1918 115 1919 116
rect 1923 115 1924 119
rect 1918 114 1924 115
rect 1927 119 1933 120
rect 1927 115 1928 119
rect 1932 118 1933 119
rect 1966 119 1972 120
rect 1966 118 1967 119
rect 1932 116 1967 118
rect 1932 115 1933 116
rect 1927 114 1933 115
rect 1966 115 1967 116
rect 1971 115 1972 119
rect 1966 114 1972 115
rect 1974 119 1981 120
rect 1974 115 1975 119
rect 1980 115 1981 119
rect 1974 114 1981 115
rect 2015 119 2021 120
rect 2015 115 2016 119
rect 2020 118 2021 119
rect 2046 119 2052 120
rect 2046 118 2047 119
rect 2020 116 2047 118
rect 2020 115 2021 116
rect 2015 114 2021 115
rect 2046 115 2047 116
rect 2051 115 2052 119
rect 2046 114 2052 115
rect 2055 119 2061 120
rect 2055 115 2056 119
rect 2060 118 2061 119
rect 2086 119 2092 120
rect 2086 118 2087 119
rect 2060 116 2087 118
rect 2060 115 2061 116
rect 2055 114 2061 115
rect 2086 115 2087 116
rect 2091 115 2092 119
rect 2086 114 2092 115
rect 2094 119 2101 120
rect 2094 115 2095 119
rect 2100 115 2101 119
rect 2094 114 2101 115
rect 110 112 116 113
rect 110 108 111 112
rect 115 108 116 112
rect 1094 112 1100 113
rect 1094 108 1095 112
rect 1099 108 1100 112
rect 110 107 116 108
rect 190 107 196 108
rect 190 103 191 107
rect 195 106 196 107
rect 199 107 205 108
rect 199 106 200 107
rect 195 104 200 106
rect 195 103 196 104
rect 190 102 196 103
rect 199 103 200 104
rect 204 103 205 107
rect 199 102 205 103
rect 230 107 236 108
rect 230 103 231 107
rect 235 106 236 107
rect 239 107 245 108
rect 239 106 240 107
rect 235 104 240 106
rect 235 103 236 104
rect 230 102 236 103
rect 239 103 240 104
rect 244 103 245 107
rect 239 102 245 103
rect 270 107 276 108
rect 270 103 271 107
rect 275 106 276 107
rect 279 107 285 108
rect 279 106 280 107
rect 275 104 280 106
rect 275 103 276 104
rect 270 102 276 103
rect 279 103 280 104
rect 284 103 285 107
rect 279 102 285 103
rect 302 107 308 108
rect 302 103 303 107
rect 307 106 308 107
rect 319 107 325 108
rect 319 106 320 107
rect 307 104 320 106
rect 307 103 308 104
rect 302 102 308 103
rect 319 103 320 104
rect 324 103 325 107
rect 319 102 325 103
rect 350 107 356 108
rect 350 103 351 107
rect 355 106 356 107
rect 359 107 365 108
rect 359 106 360 107
rect 355 104 360 106
rect 355 103 356 104
rect 350 102 356 103
rect 359 103 360 104
rect 364 103 365 107
rect 359 102 365 103
rect 390 107 396 108
rect 390 103 391 107
rect 395 106 396 107
rect 399 107 405 108
rect 399 106 400 107
rect 395 104 400 106
rect 395 103 396 104
rect 390 102 396 103
rect 399 103 400 104
rect 404 103 405 107
rect 399 102 405 103
rect 430 107 436 108
rect 430 103 431 107
rect 435 106 436 107
rect 439 107 445 108
rect 439 106 440 107
rect 435 104 440 106
rect 435 103 436 104
rect 430 102 436 103
rect 439 103 440 104
rect 444 103 445 107
rect 439 102 445 103
rect 470 107 476 108
rect 470 103 471 107
rect 475 106 476 107
rect 479 107 485 108
rect 479 106 480 107
rect 475 104 480 106
rect 475 103 476 104
rect 470 102 476 103
rect 479 103 480 104
rect 484 103 485 107
rect 479 102 485 103
rect 510 107 516 108
rect 510 103 511 107
rect 515 106 516 107
rect 519 107 525 108
rect 519 106 520 107
rect 515 104 520 106
rect 515 103 516 104
rect 510 102 516 103
rect 519 103 520 104
rect 524 103 525 107
rect 519 102 525 103
rect 554 107 565 108
rect 554 103 555 107
rect 559 103 560 107
rect 564 103 565 107
rect 554 102 565 103
rect 590 107 596 108
rect 590 103 591 107
rect 595 106 596 107
rect 599 107 605 108
rect 599 106 600 107
rect 595 104 600 106
rect 595 103 596 104
rect 590 102 596 103
rect 599 103 600 104
rect 604 103 605 107
rect 599 102 605 103
rect 630 107 636 108
rect 630 103 631 107
rect 635 106 636 107
rect 639 107 645 108
rect 639 106 640 107
rect 635 104 640 106
rect 635 103 636 104
rect 630 102 636 103
rect 639 103 640 104
rect 644 103 645 107
rect 639 102 645 103
rect 670 107 676 108
rect 670 103 671 107
rect 675 106 676 107
rect 679 107 685 108
rect 679 106 680 107
rect 675 104 680 106
rect 675 103 676 104
rect 670 102 676 103
rect 679 103 680 104
rect 684 103 685 107
rect 679 102 685 103
rect 710 107 716 108
rect 710 103 711 107
rect 715 106 716 107
rect 719 107 725 108
rect 719 106 720 107
rect 715 104 720 106
rect 715 103 716 104
rect 710 102 716 103
rect 719 103 720 104
rect 724 103 725 107
rect 719 102 725 103
rect 750 107 756 108
rect 750 103 751 107
rect 755 106 756 107
rect 759 107 765 108
rect 759 106 760 107
rect 755 104 760 106
rect 755 103 756 104
rect 750 102 756 103
rect 759 103 760 104
rect 764 103 765 107
rect 759 102 765 103
rect 790 107 796 108
rect 790 103 791 107
rect 795 106 796 107
rect 799 107 805 108
rect 799 106 800 107
rect 795 104 800 106
rect 795 103 796 104
rect 790 102 796 103
rect 799 103 800 104
rect 804 103 805 107
rect 799 102 805 103
rect 830 107 836 108
rect 830 103 831 107
rect 835 106 836 107
rect 839 107 845 108
rect 839 106 840 107
rect 835 104 840 106
rect 835 103 836 104
rect 830 102 836 103
rect 839 103 840 104
rect 844 103 845 107
rect 839 102 845 103
rect 886 107 892 108
rect 886 103 887 107
rect 891 106 892 107
rect 895 107 901 108
rect 895 106 896 107
rect 891 104 896 106
rect 891 103 892 104
rect 886 102 892 103
rect 895 103 896 104
rect 900 103 901 107
rect 895 102 901 103
rect 942 107 948 108
rect 942 103 943 107
rect 947 106 948 107
rect 959 107 965 108
rect 959 106 960 107
rect 947 104 960 106
rect 947 103 948 104
rect 942 102 948 103
rect 959 103 960 104
rect 964 103 965 107
rect 959 102 965 103
rect 1018 107 1029 108
rect 1018 103 1019 107
rect 1023 103 1024 107
rect 1028 103 1029 107
rect 1018 102 1029 103
rect 1062 107 1068 108
rect 1062 103 1063 107
rect 1067 106 1068 107
rect 1071 107 1077 108
rect 1094 107 1100 108
rect 1158 112 1164 113
rect 1158 108 1159 112
rect 1163 108 1164 112
rect 1158 107 1164 108
rect 1198 112 1204 113
rect 1198 108 1199 112
rect 1203 108 1204 112
rect 1198 107 1204 108
rect 1238 112 1244 113
rect 1238 108 1239 112
rect 1243 108 1244 112
rect 1238 107 1244 108
rect 1278 112 1284 113
rect 1278 108 1279 112
rect 1283 108 1284 112
rect 1278 107 1284 108
rect 1318 112 1324 113
rect 1318 108 1319 112
rect 1323 108 1324 112
rect 1318 107 1324 108
rect 1366 112 1372 113
rect 1366 108 1367 112
rect 1371 108 1372 112
rect 1366 107 1372 108
rect 1430 112 1436 113
rect 1430 108 1431 112
rect 1435 108 1436 112
rect 1430 107 1436 108
rect 1494 112 1500 113
rect 1494 108 1495 112
rect 1499 108 1500 112
rect 1494 107 1500 108
rect 1558 112 1564 113
rect 1558 108 1559 112
rect 1563 108 1564 112
rect 1558 107 1564 108
rect 1614 112 1620 113
rect 1614 108 1615 112
rect 1619 108 1620 112
rect 1614 107 1620 108
rect 1670 112 1676 113
rect 1670 108 1671 112
rect 1675 108 1676 112
rect 1670 107 1676 108
rect 1718 112 1724 113
rect 1718 108 1719 112
rect 1723 108 1724 112
rect 1718 107 1724 108
rect 1766 112 1772 113
rect 1766 108 1767 112
rect 1771 108 1772 112
rect 1766 107 1772 108
rect 1806 112 1812 113
rect 1806 108 1807 112
rect 1811 108 1812 112
rect 1806 107 1812 108
rect 1854 112 1860 113
rect 1854 108 1855 112
rect 1859 108 1860 112
rect 1854 107 1860 108
rect 1902 112 1908 113
rect 1902 108 1903 112
rect 1907 108 1908 112
rect 1902 107 1908 108
rect 1950 112 1956 113
rect 1950 108 1951 112
rect 1955 108 1956 112
rect 1950 107 1956 108
rect 1990 112 1996 113
rect 1990 108 1991 112
rect 1995 108 1996 112
rect 1990 107 1996 108
rect 2030 112 2036 113
rect 2030 108 2031 112
rect 2035 108 2036 112
rect 2030 107 2036 108
rect 2070 112 2076 113
rect 2070 108 2071 112
rect 2075 108 2076 112
rect 2070 107 2076 108
rect 1071 106 1072 107
rect 1067 104 1072 106
rect 1067 103 1068 104
rect 1062 102 1068 103
rect 1071 103 1072 104
rect 1076 103 1077 107
rect 1071 102 1077 103
rect 1134 104 1140 105
rect 1134 100 1135 104
rect 1139 100 1140 104
rect 2118 104 2124 105
rect 2118 100 2119 104
rect 2123 100 2124 104
rect 1134 99 1140 100
rect 1174 99 1180 100
rect 110 95 116 96
rect 110 91 111 95
rect 115 91 116 95
rect 1094 95 1100 96
rect 110 90 116 91
rect 134 92 140 93
rect 134 88 135 92
rect 139 88 140 92
rect 134 87 140 88
rect 174 92 180 93
rect 174 88 175 92
rect 179 88 180 92
rect 174 87 180 88
rect 214 92 220 93
rect 214 88 215 92
rect 219 88 220 92
rect 214 87 220 88
rect 254 92 260 93
rect 254 88 255 92
rect 259 88 260 92
rect 254 87 260 88
rect 294 92 300 93
rect 294 88 295 92
rect 299 88 300 92
rect 294 87 300 88
rect 334 92 340 93
rect 334 88 335 92
rect 339 88 340 92
rect 334 87 340 88
rect 374 92 380 93
rect 374 88 375 92
rect 379 88 380 92
rect 374 87 380 88
rect 414 92 420 93
rect 414 88 415 92
rect 419 88 420 92
rect 414 87 420 88
rect 454 92 460 93
rect 454 88 455 92
rect 459 88 460 92
rect 454 87 460 88
rect 494 92 500 93
rect 494 88 495 92
rect 499 88 500 92
rect 494 87 500 88
rect 534 92 540 93
rect 534 88 535 92
rect 539 88 540 92
rect 534 87 540 88
rect 574 92 580 93
rect 574 88 575 92
rect 579 88 580 92
rect 574 87 580 88
rect 614 92 620 93
rect 614 88 615 92
rect 619 88 620 92
rect 614 87 620 88
rect 654 92 660 93
rect 654 88 655 92
rect 659 88 660 92
rect 654 87 660 88
rect 694 92 700 93
rect 694 88 695 92
rect 699 88 700 92
rect 694 87 700 88
rect 734 92 740 93
rect 734 88 735 92
rect 739 88 740 92
rect 734 87 740 88
rect 774 92 780 93
rect 774 88 775 92
rect 779 88 780 92
rect 774 87 780 88
rect 814 92 820 93
rect 814 88 815 92
rect 819 88 820 92
rect 814 87 820 88
rect 870 92 876 93
rect 870 88 871 92
rect 875 88 876 92
rect 870 87 876 88
rect 934 92 940 93
rect 934 88 935 92
rect 939 88 940 92
rect 934 87 940 88
rect 998 92 1004 93
rect 998 88 999 92
rect 1003 88 1004 92
rect 998 87 1004 88
rect 1046 92 1052 93
rect 1046 88 1047 92
rect 1051 88 1052 92
rect 1094 91 1095 95
rect 1099 91 1100 95
rect 1174 95 1175 99
rect 1179 98 1180 99
rect 1183 99 1189 100
rect 1183 98 1184 99
rect 1179 96 1184 98
rect 1179 95 1180 96
rect 1174 94 1180 95
rect 1183 95 1184 96
rect 1188 95 1189 99
rect 1183 94 1189 95
rect 1214 99 1220 100
rect 1214 95 1215 99
rect 1219 98 1220 99
rect 1223 99 1229 100
rect 1223 98 1224 99
rect 1219 96 1224 98
rect 1219 95 1220 96
rect 1214 94 1220 95
rect 1223 95 1224 96
rect 1228 95 1229 99
rect 1223 94 1229 95
rect 1254 99 1260 100
rect 1254 95 1255 99
rect 1259 98 1260 99
rect 1263 99 1269 100
rect 1263 98 1264 99
rect 1259 96 1264 98
rect 1259 95 1260 96
rect 1254 94 1260 95
rect 1263 95 1264 96
rect 1268 95 1269 99
rect 1263 94 1269 95
rect 1294 99 1300 100
rect 1294 95 1295 99
rect 1299 98 1300 99
rect 1303 99 1309 100
rect 1303 98 1304 99
rect 1299 96 1304 98
rect 1299 95 1300 96
rect 1294 94 1300 95
rect 1303 95 1304 96
rect 1308 95 1309 99
rect 1303 94 1309 95
rect 1334 99 1340 100
rect 1334 95 1335 99
rect 1339 98 1340 99
rect 1343 99 1349 100
rect 1343 98 1344 99
rect 1339 96 1344 98
rect 1339 95 1340 96
rect 1334 94 1340 95
rect 1343 95 1344 96
rect 1348 95 1349 99
rect 1343 94 1349 95
rect 1382 99 1388 100
rect 1382 95 1383 99
rect 1387 98 1388 99
rect 1391 99 1397 100
rect 1391 98 1392 99
rect 1387 96 1392 98
rect 1387 95 1388 96
rect 1382 94 1388 95
rect 1391 95 1392 96
rect 1396 95 1397 99
rect 1391 94 1397 95
rect 1446 99 1452 100
rect 1446 95 1447 99
rect 1451 98 1452 99
rect 1455 99 1461 100
rect 1455 98 1456 99
rect 1451 96 1456 98
rect 1451 95 1452 96
rect 1446 94 1452 95
rect 1455 95 1456 96
rect 1460 95 1461 99
rect 1455 94 1461 95
rect 1502 99 1508 100
rect 1502 95 1503 99
rect 1507 98 1508 99
rect 1519 99 1525 100
rect 1519 98 1520 99
rect 1507 96 1520 98
rect 1507 95 1508 96
rect 1502 94 1508 95
rect 1519 95 1520 96
rect 1524 95 1525 99
rect 1519 94 1525 95
rect 1583 99 1589 100
rect 1583 95 1584 99
rect 1588 98 1589 99
rect 1598 99 1604 100
rect 1598 98 1599 99
rect 1588 96 1599 98
rect 1588 95 1589 96
rect 1583 94 1589 95
rect 1598 95 1599 96
rect 1603 95 1604 99
rect 1598 94 1604 95
rect 1630 99 1636 100
rect 1630 95 1631 99
rect 1635 98 1636 99
rect 1639 99 1645 100
rect 1639 98 1640 99
rect 1635 96 1640 98
rect 1635 95 1636 96
rect 1630 94 1636 95
rect 1639 95 1640 96
rect 1644 95 1645 99
rect 1639 94 1645 95
rect 1686 99 1692 100
rect 1686 95 1687 99
rect 1691 98 1692 99
rect 1695 99 1701 100
rect 1695 98 1696 99
rect 1691 96 1696 98
rect 1691 95 1692 96
rect 1686 94 1692 95
rect 1695 95 1696 96
rect 1700 95 1701 99
rect 1695 94 1701 95
rect 1734 99 1740 100
rect 1734 95 1735 99
rect 1739 98 1740 99
rect 1743 99 1749 100
rect 1743 98 1744 99
rect 1739 96 1744 98
rect 1739 95 1740 96
rect 1734 94 1740 95
rect 1743 95 1744 96
rect 1748 95 1749 99
rect 1743 94 1749 95
rect 1782 99 1788 100
rect 1782 95 1783 99
rect 1787 98 1788 99
rect 1791 99 1797 100
rect 1791 98 1792 99
rect 1787 96 1792 98
rect 1787 95 1788 96
rect 1782 94 1788 95
rect 1791 95 1792 96
rect 1796 95 1797 99
rect 1791 94 1797 95
rect 1822 99 1828 100
rect 1822 95 1823 99
rect 1827 98 1828 99
rect 1831 99 1837 100
rect 1831 98 1832 99
rect 1827 96 1832 98
rect 1827 95 1828 96
rect 1822 94 1828 95
rect 1831 95 1832 96
rect 1836 95 1837 99
rect 1831 94 1837 95
rect 1870 99 1876 100
rect 1870 95 1871 99
rect 1875 98 1876 99
rect 1879 99 1885 100
rect 1879 98 1880 99
rect 1875 96 1880 98
rect 1875 95 1876 96
rect 1870 94 1876 95
rect 1879 95 1880 96
rect 1884 95 1885 99
rect 1879 94 1885 95
rect 1918 99 1924 100
rect 1918 95 1919 99
rect 1923 98 1924 99
rect 1927 99 1933 100
rect 1927 98 1928 99
rect 1923 96 1928 98
rect 1923 95 1924 96
rect 1918 94 1924 95
rect 1927 95 1928 96
rect 1932 95 1933 99
rect 1927 94 1933 95
rect 1966 99 1972 100
rect 1966 95 1967 99
rect 1971 98 1972 99
rect 1975 99 1981 100
rect 1975 98 1976 99
rect 1971 96 1976 98
rect 1971 95 1972 96
rect 1966 94 1972 95
rect 1975 95 1976 96
rect 1980 95 1981 99
rect 1975 94 1981 95
rect 2014 99 2021 100
rect 2014 95 2015 99
rect 2020 95 2021 99
rect 2014 94 2021 95
rect 2046 99 2052 100
rect 2046 95 2047 99
rect 2051 98 2052 99
rect 2055 99 2061 100
rect 2055 98 2056 99
rect 2051 96 2056 98
rect 2051 95 2052 96
rect 2046 94 2052 95
rect 2055 95 2056 96
rect 2060 95 2061 99
rect 2055 94 2061 95
rect 2086 99 2092 100
rect 2086 95 2087 99
rect 2091 98 2092 99
rect 2095 99 2101 100
rect 2118 99 2124 100
rect 2095 98 2096 99
rect 2091 96 2096 98
rect 2091 95 2092 96
rect 2086 94 2092 95
rect 2095 95 2096 96
rect 2100 95 2101 99
rect 2095 94 2101 95
rect 1094 90 1100 91
rect 1046 87 1052 88
rect 1134 87 1140 88
rect 1134 83 1135 87
rect 1139 83 1140 87
rect 2118 87 2124 88
rect 1134 82 1140 83
rect 1158 84 1164 85
rect 1158 80 1159 84
rect 1163 80 1164 84
rect 1158 79 1164 80
rect 1198 84 1204 85
rect 1198 80 1199 84
rect 1203 80 1204 84
rect 1198 79 1204 80
rect 1238 84 1244 85
rect 1238 80 1239 84
rect 1243 80 1244 84
rect 1238 79 1244 80
rect 1278 84 1284 85
rect 1278 80 1279 84
rect 1283 80 1284 84
rect 1278 79 1284 80
rect 1318 84 1324 85
rect 1318 80 1319 84
rect 1323 80 1324 84
rect 1318 79 1324 80
rect 1366 84 1372 85
rect 1366 80 1367 84
rect 1371 80 1372 84
rect 1366 79 1372 80
rect 1430 84 1436 85
rect 1430 80 1431 84
rect 1435 80 1436 84
rect 1430 79 1436 80
rect 1494 84 1500 85
rect 1494 80 1495 84
rect 1499 80 1500 84
rect 1494 79 1500 80
rect 1558 84 1564 85
rect 1558 80 1559 84
rect 1563 80 1564 84
rect 1558 79 1564 80
rect 1614 84 1620 85
rect 1614 80 1615 84
rect 1619 80 1620 84
rect 1614 79 1620 80
rect 1670 84 1676 85
rect 1670 80 1671 84
rect 1675 80 1676 84
rect 1670 79 1676 80
rect 1718 84 1724 85
rect 1718 80 1719 84
rect 1723 80 1724 84
rect 1718 79 1724 80
rect 1766 84 1772 85
rect 1766 80 1767 84
rect 1771 80 1772 84
rect 1766 79 1772 80
rect 1806 84 1812 85
rect 1806 80 1807 84
rect 1811 80 1812 84
rect 1806 79 1812 80
rect 1854 84 1860 85
rect 1854 80 1855 84
rect 1859 80 1860 84
rect 1854 79 1860 80
rect 1902 84 1908 85
rect 1902 80 1903 84
rect 1907 80 1908 84
rect 1902 79 1908 80
rect 1950 84 1956 85
rect 1950 80 1951 84
rect 1955 80 1956 84
rect 1950 79 1956 80
rect 1990 84 1996 85
rect 1990 80 1991 84
rect 1995 80 1996 84
rect 1990 79 1996 80
rect 2030 84 2036 85
rect 2030 80 2031 84
rect 2035 80 2036 84
rect 2030 79 2036 80
rect 2070 84 2076 85
rect 2070 80 2071 84
rect 2075 80 2076 84
rect 2118 83 2119 87
rect 2123 83 2124 87
rect 2118 82 2124 83
rect 2070 79 2076 80
<< m3c >>
rect 1647 2207 1651 2211
rect 1399 2199 1403 2203
rect 1439 2199 1443 2203
rect 1479 2199 1483 2203
rect 1519 2199 1523 2203
rect 1559 2199 1563 2203
rect 1599 2199 1603 2203
rect 1639 2199 1643 2203
rect 1679 2199 1683 2203
rect 1719 2199 1723 2203
rect 1759 2199 1763 2203
rect 1799 2199 1803 2203
rect 1839 2199 1843 2203
rect 1343 2192 1347 2196
rect 1383 2192 1387 2196
rect 1423 2192 1427 2196
rect 1463 2192 1467 2196
rect 1503 2192 1507 2196
rect 1543 2192 1547 2196
rect 1583 2192 1587 2196
rect 1623 2192 1627 2196
rect 1663 2192 1667 2196
rect 1703 2192 1707 2196
rect 1743 2192 1747 2196
rect 1783 2192 1787 2196
rect 1823 2192 1827 2196
rect 1135 2184 1139 2188
rect 2119 2184 2123 2188
rect 1391 2179 1395 2183
rect 1399 2179 1403 2183
rect 1439 2179 1443 2183
rect 1479 2179 1483 2183
rect 1519 2179 1523 2183
rect 1559 2179 1563 2183
rect 1599 2179 1603 2183
rect 1639 2179 1643 2183
rect 1679 2179 1683 2183
rect 1719 2179 1723 2183
rect 1759 2179 1763 2183
rect 1799 2179 1803 2183
rect 1839 2179 1843 2183
rect 1135 2167 1139 2171
rect 1343 2164 1347 2168
rect 1383 2164 1387 2168
rect 1423 2164 1427 2168
rect 1463 2164 1467 2168
rect 1503 2164 1507 2168
rect 1543 2164 1547 2168
rect 1583 2164 1587 2168
rect 1623 2164 1627 2168
rect 1663 2164 1667 2168
rect 1703 2164 1707 2168
rect 1743 2164 1747 2168
rect 1783 2164 1787 2168
rect 1823 2164 1827 2168
rect 2119 2167 2123 2171
rect 1135 2149 1139 2153
rect 1287 2152 1291 2156
rect 1327 2152 1331 2156
rect 1367 2152 1371 2156
rect 1415 2152 1419 2156
rect 1463 2152 1467 2156
rect 1519 2152 1523 2156
rect 1575 2152 1579 2156
rect 1623 2152 1627 2156
rect 1671 2152 1675 2156
rect 1719 2152 1723 2156
rect 1775 2152 1779 2156
rect 1831 2152 1835 2156
rect 1887 2152 1891 2156
rect 2119 2149 2123 2153
rect 1135 2132 1139 2136
rect 1315 2135 1316 2139
rect 1316 2135 1319 2139
rect 1335 2135 1339 2139
rect 1375 2135 1379 2139
rect 1647 2135 1648 2139
rect 1648 2135 1651 2139
rect 1707 2135 1711 2139
rect 1755 2135 1759 2139
rect 1811 2135 1815 2139
rect 2119 2132 2123 2136
rect 1287 2124 1291 2128
rect 1327 2124 1331 2128
rect 1367 2124 1371 2128
rect 1415 2124 1419 2128
rect 1463 2124 1467 2128
rect 1519 2124 1523 2128
rect 1575 2124 1579 2128
rect 1623 2124 1627 2128
rect 1671 2124 1675 2128
rect 1719 2124 1723 2128
rect 1775 2124 1779 2128
rect 1831 2124 1835 2128
rect 1887 2124 1891 2128
rect 1335 2115 1339 2119
rect 1375 2115 1379 2119
rect 1391 2107 1395 2111
rect 1707 2115 1711 2119
rect 1755 2115 1759 2119
rect 1811 2115 1815 2119
rect 1691 2107 1695 2111
rect 1295 2091 1299 2095
rect 1351 2091 1355 2095
rect 1439 2091 1443 2095
rect 1519 2091 1523 2095
rect 1599 2091 1603 2095
rect 1607 2091 1608 2095
rect 1608 2091 1611 2095
rect 1759 2091 1763 2095
rect 1847 2091 1851 2095
rect 1935 2091 1939 2095
rect 2023 2091 2027 2095
rect 2031 2091 2032 2095
rect 2032 2091 2035 2095
rect 1223 2084 1227 2088
rect 1279 2084 1283 2088
rect 1343 2084 1347 2088
rect 1423 2084 1427 2088
rect 1503 2084 1507 2088
rect 1583 2084 1587 2088
rect 1663 2084 1667 2088
rect 1743 2084 1747 2088
rect 1831 2084 1835 2088
rect 1919 2084 1923 2088
rect 2007 2084 2011 2088
rect 2071 2084 2075 2088
rect 1135 2076 1139 2080
rect 2119 2076 2123 2080
rect 1211 2071 1215 2075
rect 1295 2071 1299 2075
rect 1351 2071 1355 2075
rect 1439 2071 1443 2075
rect 1519 2071 1523 2075
rect 1599 2071 1603 2075
rect 1691 2071 1692 2075
rect 1692 2071 1695 2075
rect 1759 2071 1763 2075
rect 1847 2071 1851 2075
rect 1935 2071 1939 2075
rect 2023 2071 2027 2075
rect 2095 2071 2096 2075
rect 2096 2071 2099 2075
rect 1135 2059 1139 2063
rect 1223 2056 1227 2060
rect 1279 2056 1283 2060
rect 1343 2056 1347 2060
rect 1423 2056 1427 2060
rect 1503 2056 1507 2060
rect 1583 2056 1587 2060
rect 1663 2056 1667 2060
rect 1743 2056 1747 2060
rect 1831 2056 1835 2060
rect 1919 2056 1923 2060
rect 2007 2056 2011 2060
rect 2071 2056 2075 2060
rect 2119 2059 2123 2063
rect 1135 2041 1139 2045
rect 1183 2044 1187 2048
rect 1239 2044 1243 2048
rect 1311 2044 1315 2048
rect 1399 2044 1403 2048
rect 1487 2044 1491 2048
rect 1583 2044 1587 2048
rect 1671 2044 1675 2048
rect 1759 2044 1763 2048
rect 1839 2044 1843 2048
rect 1919 2044 1923 2048
rect 2007 2044 2011 2048
rect 2071 2044 2075 2048
rect 2119 2041 2123 2045
rect 1863 2035 1867 2039
rect 1135 2024 1139 2028
rect 1255 2027 1259 2031
rect 1327 2027 1331 2031
rect 1415 2027 1419 2031
rect 1503 2027 1507 2031
rect 1559 2027 1563 2031
rect 1571 2027 1575 2031
rect 1935 2027 1939 2031
rect 2023 2027 2027 2031
rect 2031 2027 2032 2031
rect 2032 2027 2035 2031
rect 247 2019 251 2023
rect 303 2019 307 2023
rect 367 2019 371 2023
rect 439 2019 443 2023
rect 511 2019 515 2023
rect 539 2019 543 2023
rect 547 2019 551 2023
rect 735 2019 739 2023
rect 791 2019 795 2023
rect 855 2019 859 2023
rect 911 2019 915 2023
rect 967 2019 971 2023
rect 1023 2019 1027 2023
rect 1063 2019 1067 2023
rect 2119 2024 2123 2028
rect 1071 2019 1072 2023
rect 1072 2019 1075 2023
rect 191 2012 195 2016
rect 231 2012 235 2016
rect 287 2012 291 2016
rect 351 2012 355 2016
rect 423 2012 427 2016
rect 495 2012 499 2016
rect 575 2012 579 2016
rect 647 2012 651 2016
rect 719 2012 723 2016
rect 783 2012 787 2016
rect 839 2012 843 2016
rect 895 2012 899 2016
rect 951 2012 955 2016
rect 1007 2012 1011 2016
rect 1047 2012 1051 2016
rect 1183 2016 1187 2020
rect 1239 2016 1243 2020
rect 1311 2016 1315 2020
rect 1399 2016 1403 2020
rect 1487 2016 1491 2020
rect 1583 2016 1587 2020
rect 1671 2016 1675 2020
rect 1759 2016 1763 2020
rect 1839 2016 1843 2020
rect 1919 2016 1923 2020
rect 2007 2016 2011 2020
rect 2071 2016 2075 2020
rect 111 2004 115 2008
rect 1095 2004 1099 2008
rect 1211 2007 1212 2011
rect 1212 2007 1215 2011
rect 1255 2007 1259 2011
rect 1327 2007 1331 2011
rect 1415 2007 1419 2011
rect 1503 2007 1507 2011
rect 1559 2007 1563 2011
rect 1831 2007 1835 2011
rect 1863 2007 1864 2011
rect 1864 2007 1867 2011
rect 1935 2007 1939 2011
rect 2023 2007 2027 2011
rect 2095 2007 2096 2011
rect 2096 2007 2099 2011
rect 215 1999 216 2003
rect 216 1999 219 2003
rect 247 1999 251 2003
rect 303 1999 307 2003
rect 367 1999 371 2003
rect 439 1999 443 2003
rect 511 1999 515 2003
rect 539 1999 543 2003
rect 735 1999 739 2003
rect 791 1999 795 2003
rect 855 1999 859 2003
rect 911 1999 915 2003
rect 967 1999 971 2003
rect 1023 1999 1027 2003
rect 1063 1999 1067 2003
rect 111 1987 115 1991
rect 191 1984 195 1988
rect 231 1984 235 1988
rect 287 1984 291 1988
rect 351 1984 355 1988
rect 423 1984 427 1988
rect 495 1984 499 1988
rect 575 1984 579 1988
rect 647 1984 651 1988
rect 719 1984 723 1988
rect 783 1984 787 1988
rect 839 1984 843 1988
rect 895 1984 899 1988
rect 951 1984 955 1988
rect 1007 1984 1011 1988
rect 1047 1984 1051 1988
rect 1095 1987 1099 1991
rect 1399 1987 1403 1991
rect 1479 1987 1483 1991
rect 1551 1987 1555 1991
rect 1571 1987 1572 1991
rect 1572 1987 1575 1991
rect 1695 1987 1699 1991
rect 1767 1987 1771 1991
rect 1807 1987 1811 1991
rect 1895 1987 1899 1991
rect 1967 1987 1971 1991
rect 1975 1987 1976 1991
rect 1976 1987 1979 1991
rect 2087 1987 2091 1991
rect 1303 1980 1307 1984
rect 1383 1980 1387 1984
rect 1463 1980 1467 1984
rect 1543 1980 1547 1984
rect 1615 1980 1619 1984
rect 1687 1980 1691 1984
rect 1751 1980 1755 1984
rect 1815 1980 1819 1984
rect 1879 1980 1883 1984
rect 1951 1980 1955 1984
rect 2023 1980 2027 1984
rect 2071 1980 2075 1984
rect 111 1969 115 1973
rect 191 1972 195 1976
rect 247 1972 251 1976
rect 311 1972 315 1976
rect 375 1972 379 1976
rect 447 1972 451 1976
rect 519 1972 523 1976
rect 591 1972 595 1976
rect 655 1972 659 1976
rect 719 1972 723 1976
rect 775 1972 779 1976
rect 823 1972 827 1976
rect 871 1972 875 1976
rect 919 1972 923 1976
rect 967 1972 971 1976
rect 1007 1972 1011 1976
rect 1047 1972 1051 1976
rect 1095 1969 1099 1973
rect 1135 1972 1139 1976
rect 2119 1972 2123 1976
rect 895 1963 899 1967
rect 1071 1963 1075 1967
rect 1327 1967 1328 1971
rect 1328 1967 1331 1971
rect 1399 1967 1403 1971
rect 1479 1967 1483 1971
rect 1551 1967 1555 1971
rect 1643 1967 1644 1971
rect 1644 1967 1647 1971
rect 1695 1967 1699 1971
rect 1767 1967 1771 1971
rect 1831 1967 1835 1971
rect 1895 1967 1899 1971
rect 1967 1967 1971 1971
rect 2079 1967 2083 1971
rect 2087 1967 2091 1971
rect 111 1952 115 1956
rect 263 1955 267 1959
rect 327 1955 331 1959
rect 335 1955 336 1959
rect 336 1955 339 1959
rect 463 1955 467 1959
rect 535 1955 539 1959
rect 547 1955 548 1959
rect 548 1955 551 1959
rect 607 1955 611 1959
rect 859 1955 863 1959
rect 1015 1955 1019 1959
rect 1055 1955 1059 1959
rect 1095 1952 1099 1956
rect 1135 1955 1139 1959
rect 1303 1952 1307 1956
rect 1383 1952 1387 1956
rect 1463 1952 1467 1956
rect 1543 1952 1547 1956
rect 1615 1952 1619 1956
rect 1687 1952 1691 1956
rect 1751 1952 1755 1956
rect 1815 1952 1819 1956
rect 1879 1952 1883 1956
rect 1951 1952 1955 1956
rect 2023 1952 2027 1956
rect 2071 1952 2075 1956
rect 2119 1955 2123 1959
rect 191 1944 195 1948
rect 247 1944 251 1948
rect 311 1944 315 1948
rect 375 1944 379 1948
rect 447 1944 451 1948
rect 519 1944 523 1948
rect 591 1944 595 1948
rect 655 1944 659 1948
rect 719 1944 723 1948
rect 775 1944 779 1948
rect 823 1944 827 1948
rect 871 1944 875 1948
rect 919 1944 923 1948
rect 967 1944 971 1948
rect 1007 1944 1011 1948
rect 1047 1944 1051 1948
rect 215 1935 216 1939
rect 216 1935 219 1939
rect 263 1935 267 1939
rect 327 1935 331 1939
rect 395 1935 399 1939
rect 463 1935 467 1939
rect 535 1935 539 1939
rect 859 1935 863 1939
rect 895 1935 896 1939
rect 896 1935 899 1939
rect 1015 1935 1019 1939
rect 1055 1935 1059 1939
rect 607 1923 611 1927
rect 1135 1933 1139 1937
rect 1159 1936 1163 1940
rect 1223 1936 1227 1940
rect 1303 1936 1307 1940
rect 1383 1936 1387 1940
rect 1463 1936 1467 1940
rect 1535 1936 1539 1940
rect 1615 1936 1619 1940
rect 1695 1936 1699 1940
rect 1783 1936 1787 1940
rect 1879 1936 1883 1940
rect 1983 1936 1987 1940
rect 2071 1936 2075 1940
rect 2119 1933 2123 1937
rect 2007 1927 2011 1931
rect 191 1915 195 1919
rect 247 1915 251 1919
rect 287 1915 291 1919
rect 335 1915 339 1919
rect 439 1915 443 1919
rect 503 1915 507 1919
rect 511 1915 515 1919
rect 631 1915 635 1919
rect 687 1915 691 1919
rect 743 1915 747 1919
rect 799 1915 803 1919
rect 855 1915 859 1919
rect 1135 1916 1139 1920
rect 1399 1919 1403 1923
rect 1447 1919 1451 1923
rect 1475 1919 1479 1923
rect 1807 1919 1808 1923
rect 1808 1919 1811 1923
rect 2095 1919 2096 1923
rect 2096 1919 2099 1923
rect 2119 1916 2123 1920
rect 135 1908 139 1912
rect 175 1908 179 1912
rect 231 1908 235 1912
rect 295 1908 299 1912
rect 367 1908 371 1912
rect 431 1908 435 1912
rect 495 1908 499 1912
rect 559 1908 563 1912
rect 615 1908 619 1912
rect 671 1908 675 1912
rect 727 1908 731 1912
rect 783 1908 787 1912
rect 847 1908 851 1912
rect 1159 1908 1163 1912
rect 1223 1908 1227 1912
rect 1303 1908 1307 1912
rect 1383 1908 1387 1912
rect 1463 1908 1467 1912
rect 1535 1908 1539 1912
rect 1615 1908 1619 1912
rect 1695 1908 1699 1912
rect 1783 1908 1787 1912
rect 1879 1908 1883 1912
rect 1983 1908 1987 1912
rect 2071 1908 2075 1912
rect 111 1900 115 1904
rect 1095 1900 1099 1904
rect 159 1895 160 1899
rect 160 1895 163 1899
rect 191 1895 195 1899
rect 247 1895 251 1899
rect 287 1895 291 1899
rect 395 1895 396 1899
rect 396 1895 399 1899
rect 439 1895 443 1899
rect 503 1895 507 1899
rect 623 1895 627 1899
rect 631 1895 635 1899
rect 687 1895 691 1899
rect 743 1895 747 1899
rect 799 1895 803 1899
rect 855 1895 859 1899
rect 1207 1899 1211 1903
rect 1327 1899 1328 1903
rect 1328 1899 1331 1903
rect 1399 1899 1403 1903
rect 1447 1899 1451 1903
rect 1735 1899 1739 1903
rect 2007 1899 2008 1903
rect 2008 1899 2011 1903
rect 2079 1899 2083 1903
rect 111 1883 115 1887
rect 135 1880 139 1884
rect 175 1880 179 1884
rect 231 1880 235 1884
rect 295 1880 299 1884
rect 367 1880 371 1884
rect 431 1880 435 1884
rect 495 1880 499 1884
rect 559 1880 563 1884
rect 615 1880 619 1884
rect 671 1880 675 1884
rect 727 1880 731 1884
rect 783 1880 787 1884
rect 847 1880 851 1884
rect 1095 1883 1099 1887
rect 1215 1875 1219 1879
rect 1279 1875 1283 1879
rect 1319 1875 1323 1879
rect 1407 1875 1411 1879
rect 1463 1875 1467 1879
rect 1475 1875 1476 1879
rect 1476 1875 1479 1879
rect 1575 1875 1579 1879
rect 1647 1875 1651 1879
rect 1671 1875 1675 1879
rect 1815 1875 1819 1879
rect 1911 1875 1915 1879
rect 2087 1875 2091 1879
rect 2095 1875 2096 1879
rect 2096 1875 2099 1879
rect 111 1861 115 1865
rect 135 1864 139 1868
rect 199 1864 203 1868
rect 271 1864 275 1868
rect 335 1864 339 1868
rect 399 1864 403 1868
rect 455 1864 459 1868
rect 503 1864 507 1868
rect 551 1864 555 1868
rect 599 1864 603 1868
rect 647 1864 651 1868
rect 695 1864 699 1868
rect 751 1864 755 1868
rect 1159 1868 1163 1872
rect 1199 1868 1203 1872
rect 1263 1868 1267 1872
rect 1327 1868 1331 1872
rect 1391 1868 1395 1872
rect 1447 1868 1451 1872
rect 1503 1868 1507 1872
rect 1559 1868 1563 1872
rect 1631 1868 1635 1872
rect 1711 1868 1715 1872
rect 1799 1868 1803 1872
rect 1895 1868 1899 1872
rect 1991 1868 1995 1872
rect 2071 1868 2075 1872
rect 1095 1861 1099 1865
rect 1135 1860 1139 1864
rect 2119 1860 2123 1864
rect 111 1844 115 1848
rect 295 1855 299 1859
rect 479 1855 483 1859
rect 1207 1855 1211 1859
rect 1215 1855 1219 1859
rect 1279 1855 1283 1859
rect 1399 1855 1403 1859
rect 1407 1855 1411 1859
rect 1463 1855 1467 1859
rect 1575 1855 1579 1859
rect 1647 1855 1651 1859
rect 1735 1855 1736 1859
rect 1736 1855 1739 1859
rect 1815 1855 1819 1859
rect 1911 1855 1915 1859
rect 2079 1855 2083 1859
rect 2087 1855 2091 1859
rect 207 1847 211 1851
rect 235 1847 239 1851
rect 511 1847 515 1851
rect 519 1847 523 1851
rect 1095 1844 1099 1848
rect 1135 1843 1139 1847
rect 135 1836 139 1840
rect 199 1836 203 1840
rect 271 1836 275 1840
rect 335 1836 339 1840
rect 399 1836 403 1840
rect 455 1836 459 1840
rect 503 1836 507 1840
rect 551 1836 555 1840
rect 599 1836 603 1840
rect 647 1836 651 1840
rect 695 1836 699 1840
rect 751 1836 755 1840
rect 1159 1840 1163 1844
rect 1199 1840 1203 1844
rect 1263 1840 1267 1844
rect 1327 1840 1331 1844
rect 1391 1840 1395 1844
rect 1447 1840 1451 1844
rect 1503 1840 1507 1844
rect 1559 1840 1563 1844
rect 1631 1840 1635 1844
rect 1711 1840 1715 1844
rect 1799 1840 1803 1844
rect 1895 1840 1899 1844
rect 1991 1840 1995 1844
rect 2071 1840 2075 1844
rect 2119 1843 2123 1847
rect 159 1827 160 1831
rect 160 1827 163 1831
rect 235 1827 239 1831
rect 295 1827 296 1831
rect 296 1827 299 1831
rect 439 1827 443 1831
rect 479 1827 480 1831
rect 480 1827 483 1831
rect 623 1819 627 1823
rect 1135 1825 1139 1829
rect 1159 1828 1163 1832
rect 1231 1828 1235 1832
rect 1303 1828 1307 1832
rect 1383 1828 1387 1832
rect 1463 1828 1467 1832
rect 1551 1828 1555 1832
rect 1647 1828 1651 1832
rect 1751 1828 1755 1832
rect 1855 1828 1859 1832
rect 1967 1828 1971 1832
rect 2071 1828 2075 1832
rect 2119 1825 2123 1829
rect 519 1807 523 1811
rect 1135 1808 1139 1812
rect 1247 1811 1251 1815
rect 1311 1811 1315 1815
rect 1319 1811 1323 1815
rect 1479 1811 1483 1815
rect 1559 1811 1563 1815
rect 1567 1811 1571 1815
rect 1671 1811 1672 1815
rect 1672 1811 1675 1815
rect 1951 1811 1955 1815
rect 1959 1811 1963 1815
rect 2095 1811 2096 1815
rect 2096 1811 2099 1815
rect 2119 1808 2123 1812
rect 207 1799 211 1803
rect 223 1799 227 1803
rect 375 1799 379 1803
rect 391 1799 395 1803
rect 543 1799 547 1803
rect 591 1799 595 1803
rect 639 1799 643 1803
rect 151 1792 155 1796
rect 215 1792 219 1796
rect 271 1792 275 1796
rect 327 1792 331 1796
rect 383 1792 387 1796
rect 431 1792 435 1796
rect 479 1792 483 1796
rect 527 1792 531 1796
rect 575 1792 579 1796
rect 623 1792 627 1796
rect 719 1799 723 1803
rect 1159 1800 1163 1804
rect 1231 1800 1235 1804
rect 1303 1800 1307 1804
rect 1383 1800 1387 1804
rect 1463 1800 1467 1804
rect 1551 1800 1555 1804
rect 1647 1800 1651 1804
rect 1751 1800 1755 1804
rect 1855 1800 1859 1804
rect 1967 1800 1971 1804
rect 2071 1800 2075 1804
rect 671 1792 675 1796
rect 727 1792 731 1796
rect 1215 1791 1219 1795
rect 1247 1791 1251 1795
rect 1311 1791 1315 1795
rect 1399 1791 1403 1795
rect 1479 1791 1483 1795
rect 1559 1791 1563 1795
rect 1715 1791 1719 1795
rect 1959 1791 1963 1795
rect 2031 1791 2035 1795
rect 2079 1791 2083 1795
rect 111 1784 115 1788
rect 223 1779 227 1783
rect 259 1779 263 1783
rect 391 1779 395 1783
rect 439 1779 443 1783
rect 1095 1784 1099 1788
rect 543 1779 547 1783
rect 591 1779 595 1783
rect 639 1779 643 1783
rect 719 1779 723 1783
rect 783 1779 787 1783
rect 111 1767 115 1771
rect 151 1764 155 1768
rect 215 1764 219 1768
rect 271 1764 275 1768
rect 327 1764 331 1768
rect 383 1764 387 1768
rect 431 1764 435 1768
rect 479 1764 483 1768
rect 527 1764 531 1768
rect 575 1764 579 1768
rect 623 1764 627 1768
rect 671 1764 675 1768
rect 727 1764 731 1768
rect 1095 1767 1099 1771
rect 1271 1771 1275 1775
rect 1335 1771 1339 1775
rect 1367 1771 1371 1775
rect 1471 1771 1475 1775
rect 1543 1771 1547 1775
rect 1567 1775 1571 1779
rect 1695 1771 1699 1775
rect 1703 1771 1707 1775
rect 1863 1771 1867 1775
rect 1943 1771 1947 1775
rect 1951 1771 1952 1775
rect 1952 1771 1955 1775
rect 2015 1771 2019 1775
rect 2095 1771 2096 1775
rect 2096 1771 2099 1775
rect 1191 1764 1195 1768
rect 1255 1764 1259 1768
rect 1319 1764 1323 1768
rect 1383 1764 1387 1768
rect 1455 1764 1459 1768
rect 1527 1764 1531 1768
rect 1607 1764 1611 1768
rect 1687 1764 1691 1768
rect 1767 1764 1771 1768
rect 1847 1764 1851 1768
rect 1927 1764 1931 1768
rect 2007 1764 2011 1768
rect 2071 1764 2075 1768
rect 111 1749 115 1753
rect 231 1752 235 1756
rect 295 1752 299 1756
rect 351 1752 355 1756
rect 415 1752 419 1756
rect 479 1752 483 1756
rect 543 1752 547 1756
rect 615 1752 619 1756
rect 687 1752 691 1756
rect 759 1752 763 1756
rect 831 1752 835 1756
rect 911 1752 915 1756
rect 991 1752 995 1756
rect 1135 1756 1139 1760
rect 2119 1756 2123 1760
rect 1095 1749 1099 1753
rect 1215 1751 1216 1755
rect 1216 1751 1219 1755
rect 1271 1751 1275 1755
rect 1335 1751 1339 1755
rect 1411 1751 1412 1755
rect 1412 1751 1415 1755
rect 1471 1751 1475 1755
rect 1543 1751 1547 1755
rect 1703 1751 1707 1755
rect 1715 1751 1716 1755
rect 1716 1751 1719 1755
rect 1783 1751 1787 1755
rect 1863 1751 1867 1755
rect 1943 1751 1947 1755
rect 2031 1751 2032 1755
rect 2032 1751 2035 1755
rect 2095 1751 2096 1755
rect 2096 1751 2099 1755
rect 111 1732 115 1736
rect 287 1735 291 1739
rect 307 1735 311 1739
rect 375 1735 376 1739
rect 376 1735 379 1739
rect 463 1735 467 1739
rect 663 1735 667 1739
rect 675 1735 679 1739
rect 927 1735 931 1739
rect 1003 1735 1007 1739
rect 1011 1735 1015 1739
rect 1135 1739 1139 1743
rect 1095 1732 1099 1736
rect 1191 1736 1195 1740
rect 1255 1736 1259 1740
rect 1319 1736 1323 1740
rect 1383 1736 1387 1740
rect 1455 1736 1459 1740
rect 1527 1736 1531 1740
rect 1607 1736 1611 1740
rect 1687 1736 1691 1740
rect 1767 1736 1771 1740
rect 1847 1736 1851 1740
rect 1927 1736 1931 1740
rect 2007 1736 2011 1740
rect 2071 1736 2075 1740
rect 2119 1739 2123 1743
rect 231 1724 235 1728
rect 295 1724 299 1728
rect 351 1724 355 1728
rect 415 1724 419 1728
rect 479 1724 483 1728
rect 543 1724 547 1728
rect 615 1724 619 1728
rect 687 1724 691 1728
rect 759 1724 763 1728
rect 831 1724 835 1728
rect 911 1724 915 1728
rect 991 1724 995 1728
rect 1135 1721 1139 1725
rect 1247 1724 1251 1728
rect 1295 1724 1299 1728
rect 1343 1724 1347 1728
rect 1399 1724 1403 1728
rect 1463 1724 1467 1728
rect 1527 1724 1531 1728
rect 1599 1724 1603 1728
rect 1671 1724 1675 1728
rect 1743 1724 1747 1728
rect 1807 1724 1811 1728
rect 1879 1724 1883 1728
rect 1951 1724 1955 1728
rect 2023 1724 2027 1728
rect 2071 1724 2075 1728
rect 2119 1721 2123 1725
rect 259 1715 260 1719
rect 260 1715 263 1719
rect 287 1715 291 1719
rect 463 1715 467 1719
rect 571 1715 572 1719
rect 572 1715 575 1719
rect 675 1715 679 1719
rect 783 1715 784 1719
rect 784 1715 787 1719
rect 799 1715 803 1719
rect 927 1715 931 1719
rect 1003 1715 1007 1719
rect 1135 1704 1139 1708
rect 1311 1707 1315 1711
rect 1359 1707 1363 1711
rect 1367 1707 1368 1711
rect 1368 1707 1371 1711
rect 1479 1707 1483 1711
rect 1535 1707 1539 1711
rect 1543 1707 1547 1711
rect 1687 1707 1691 1711
rect 1695 1707 1696 1711
rect 1696 1707 1699 1711
rect 1815 1707 1819 1711
rect 1895 1707 1899 1711
rect 1935 1707 1939 1711
rect 2015 1707 2019 1711
rect 2047 1707 2048 1711
rect 2048 1707 2051 1711
rect 2119 1704 2123 1708
rect 1247 1696 1251 1700
rect 207 1691 211 1695
rect 295 1691 299 1695
rect 307 1691 308 1695
rect 308 1691 311 1695
rect 315 1691 319 1695
rect 663 1691 664 1695
rect 664 1691 667 1695
rect 807 1691 811 1695
rect 863 1691 867 1695
rect 871 1691 875 1695
rect 999 1691 1003 1695
rect 1011 1691 1012 1695
rect 1012 1691 1015 1695
rect 1295 1696 1299 1700
rect 1343 1696 1347 1700
rect 1399 1696 1403 1700
rect 1463 1696 1467 1700
rect 1527 1696 1531 1700
rect 1599 1696 1603 1700
rect 1671 1696 1675 1700
rect 1743 1696 1747 1700
rect 1807 1696 1811 1700
rect 1879 1696 1883 1700
rect 1951 1696 1955 1700
rect 2023 1696 2027 1700
rect 2071 1696 2075 1700
rect 135 1684 139 1688
rect 199 1684 203 1688
rect 279 1684 283 1688
rect 367 1684 371 1688
rect 463 1684 467 1688
rect 551 1684 555 1688
rect 639 1684 643 1688
rect 719 1684 723 1688
rect 791 1684 795 1688
rect 855 1684 859 1688
rect 919 1684 923 1688
rect 983 1684 987 1688
rect 1047 1684 1051 1688
rect 1287 1687 1291 1691
rect 1311 1687 1315 1691
rect 1359 1687 1363 1691
rect 1411 1687 1415 1691
rect 1479 1687 1483 1691
rect 1535 1687 1539 1691
rect 1611 1687 1615 1691
rect 1687 1687 1691 1691
rect 1783 1691 1787 1695
rect 1815 1687 1819 1691
rect 1895 1687 1899 1691
rect 1987 1687 1991 1691
rect 2095 1687 2096 1691
rect 2096 1687 2099 1691
rect 111 1676 115 1680
rect 191 1671 195 1675
rect 207 1671 211 1675
rect 295 1671 299 1675
rect 571 1671 575 1675
rect 611 1671 615 1675
rect 799 1671 803 1675
rect 807 1671 811 1675
rect 863 1671 867 1675
rect 1095 1676 1099 1680
rect 999 1671 1003 1675
rect 1035 1671 1039 1675
rect 111 1659 115 1663
rect 135 1656 139 1660
rect 199 1656 203 1660
rect 279 1656 283 1660
rect 367 1656 371 1660
rect 463 1656 467 1660
rect 551 1656 555 1660
rect 639 1656 643 1660
rect 719 1656 723 1660
rect 791 1656 795 1660
rect 855 1656 859 1660
rect 919 1656 923 1660
rect 983 1656 987 1660
rect 1047 1656 1051 1660
rect 1095 1659 1099 1663
rect 1319 1663 1323 1667
rect 1359 1663 1363 1667
rect 1407 1663 1411 1667
rect 1463 1663 1467 1667
rect 1519 1663 1523 1667
rect 1543 1667 1547 1671
rect 1643 1663 1647 1667
rect 1651 1663 1655 1667
rect 1775 1663 1779 1667
rect 1847 1663 1851 1667
rect 1927 1663 1931 1667
rect 1935 1663 1936 1667
rect 1936 1663 1939 1667
rect 2011 1663 2015 1667
rect 2047 1663 2051 1667
rect 1263 1656 1267 1660
rect 1303 1656 1307 1660
rect 1343 1656 1347 1660
rect 1391 1656 1395 1660
rect 1447 1656 1451 1660
rect 1503 1656 1507 1660
rect 1567 1656 1571 1660
rect 1631 1656 1635 1660
rect 1695 1656 1699 1660
rect 1759 1656 1763 1660
rect 1831 1656 1835 1660
rect 1911 1656 1915 1660
rect 1999 1656 2003 1660
rect 2071 1656 2075 1660
rect 1135 1648 1139 1652
rect 2119 1648 2123 1652
rect 111 1637 115 1641
rect 135 1640 139 1644
rect 183 1640 187 1644
rect 263 1640 267 1644
rect 343 1640 347 1644
rect 423 1640 427 1644
rect 503 1640 507 1644
rect 583 1640 587 1644
rect 655 1640 659 1644
rect 727 1640 731 1644
rect 791 1640 795 1644
rect 847 1640 851 1644
rect 903 1640 907 1644
rect 959 1640 963 1644
rect 1007 1640 1011 1644
rect 1047 1640 1051 1644
rect 1287 1643 1288 1647
rect 1288 1643 1291 1647
rect 1319 1643 1323 1647
rect 1359 1643 1363 1647
rect 1407 1643 1411 1647
rect 1463 1643 1467 1647
rect 1519 1643 1523 1647
rect 1611 1643 1615 1647
rect 1643 1643 1647 1647
rect 1735 1643 1739 1647
rect 1775 1643 1779 1647
rect 1847 1643 1851 1647
rect 1927 1643 1931 1647
rect 1987 1643 1991 1647
rect 2095 1643 2096 1647
rect 2096 1643 2099 1647
rect 1095 1637 1099 1641
rect 315 1631 319 1635
rect 111 1620 115 1624
rect 159 1623 160 1627
rect 160 1623 163 1627
rect 171 1623 175 1627
rect 671 1623 675 1627
rect 803 1623 807 1627
rect 863 1623 867 1627
rect 871 1623 872 1627
rect 872 1623 875 1627
rect 931 1623 932 1627
rect 932 1623 935 1627
rect 939 1623 943 1627
rect 1115 1627 1119 1631
rect 1135 1631 1139 1635
rect 1263 1628 1267 1632
rect 1303 1628 1307 1632
rect 1343 1628 1347 1632
rect 1391 1628 1395 1632
rect 1447 1628 1451 1632
rect 1503 1628 1507 1632
rect 1567 1628 1571 1632
rect 1631 1628 1635 1632
rect 1695 1628 1699 1632
rect 1759 1628 1763 1632
rect 1831 1628 1835 1632
rect 1911 1628 1915 1632
rect 1999 1628 2003 1632
rect 2071 1628 2075 1632
rect 2119 1631 2123 1635
rect 1095 1620 1099 1624
rect 135 1612 139 1616
rect 183 1612 187 1616
rect 263 1612 267 1616
rect 343 1612 347 1616
rect 423 1612 427 1616
rect 503 1612 507 1616
rect 583 1612 587 1616
rect 655 1612 659 1616
rect 727 1612 731 1616
rect 779 1615 783 1619
rect 791 1612 795 1616
rect 847 1612 851 1616
rect 903 1612 907 1616
rect 959 1612 963 1616
rect 1007 1612 1011 1616
rect 1047 1612 1051 1616
rect 171 1603 175 1607
rect 191 1603 195 1607
rect 483 1603 487 1607
rect 611 1603 612 1607
rect 612 1603 615 1607
rect 671 1603 675 1607
rect 767 1603 771 1607
rect 803 1603 807 1607
rect 863 1603 867 1607
rect 939 1603 943 1607
rect 1035 1603 1036 1607
rect 1036 1603 1039 1607
rect 931 1595 935 1599
rect 1135 1601 1139 1605
rect 1159 1604 1163 1608
rect 1215 1604 1219 1608
rect 1303 1604 1307 1608
rect 1383 1604 1387 1608
rect 1463 1604 1467 1608
rect 1543 1604 1547 1608
rect 1623 1604 1627 1608
rect 1711 1604 1715 1608
rect 1799 1604 1803 1608
rect 1887 1604 1891 1608
rect 1983 1604 1987 1608
rect 2071 1604 2075 1608
rect 2119 1601 2123 1605
rect 1615 1595 1619 1599
rect 159 1583 160 1587
rect 160 1583 163 1587
rect 183 1583 187 1587
rect 591 1583 595 1587
rect 607 1583 611 1587
rect 707 1583 711 1587
rect 779 1583 783 1587
rect 135 1576 139 1580
rect 175 1576 179 1580
rect 231 1576 235 1580
rect 303 1576 307 1580
rect 375 1576 379 1580
rect 455 1576 459 1580
rect 527 1576 531 1580
rect 599 1576 603 1580
rect 671 1576 675 1580
rect 743 1576 747 1580
rect 815 1576 819 1580
rect 1135 1584 1139 1588
rect 1231 1587 1235 1591
rect 1319 1587 1323 1591
rect 1399 1587 1403 1591
rect 1651 1587 1652 1591
rect 1652 1587 1655 1591
rect 1775 1587 1779 1591
rect 1783 1587 1787 1591
rect 2011 1587 2012 1591
rect 2012 1587 2015 1591
rect 2119 1584 2123 1588
rect 887 1576 891 1580
rect 1159 1576 1163 1580
rect 1215 1576 1219 1580
rect 1303 1576 1307 1580
rect 1383 1576 1387 1580
rect 1463 1576 1467 1580
rect 1503 1579 1507 1583
rect 1543 1576 1547 1580
rect 1623 1576 1627 1580
rect 1711 1576 1715 1580
rect 1799 1576 1803 1580
rect 1887 1576 1891 1580
rect 1983 1576 1987 1580
rect 2071 1576 2075 1580
rect 111 1568 115 1572
rect 1095 1568 1099 1572
rect 183 1563 187 1567
rect 483 1563 484 1567
rect 484 1563 487 1567
rect 607 1563 611 1567
rect 707 1563 711 1567
rect 767 1563 768 1567
rect 768 1563 771 1567
rect 851 1563 855 1567
rect 1115 1567 1119 1571
rect 1231 1567 1235 1571
rect 1319 1567 1323 1571
rect 1399 1567 1403 1571
rect 1583 1567 1587 1571
rect 1615 1567 1619 1571
rect 1735 1567 1736 1571
rect 1736 1567 1739 1571
rect 1947 1567 1951 1571
rect 2095 1567 2096 1571
rect 2096 1567 2099 1571
rect 1775 1559 1779 1563
rect 111 1551 115 1555
rect 135 1548 139 1552
rect 175 1548 179 1552
rect 231 1548 235 1552
rect 303 1548 307 1552
rect 375 1548 379 1552
rect 455 1548 459 1552
rect 527 1548 531 1552
rect 599 1548 603 1552
rect 671 1548 675 1552
rect 743 1548 747 1552
rect 815 1548 819 1552
rect 887 1548 891 1552
rect 1095 1551 1099 1555
rect 1215 1547 1219 1551
rect 1255 1547 1259 1551
rect 1335 1547 1339 1551
rect 1415 1547 1419 1551
rect 1495 1547 1499 1551
rect 1503 1547 1504 1551
rect 1504 1547 1507 1551
rect 1663 1547 1667 1551
rect 1751 1547 1755 1551
rect 1783 1547 1787 1551
rect 1799 1547 1803 1551
rect 111 1533 115 1537
rect 135 1536 139 1540
rect 175 1536 179 1540
rect 231 1536 235 1540
rect 311 1536 315 1540
rect 391 1536 395 1540
rect 479 1536 483 1540
rect 567 1536 571 1540
rect 655 1536 659 1540
rect 743 1536 747 1540
rect 823 1536 827 1540
rect 911 1536 915 1540
rect 999 1536 1003 1540
rect 1159 1540 1163 1544
rect 1199 1540 1203 1544
rect 1247 1540 1251 1544
rect 1319 1540 1323 1544
rect 1399 1540 1403 1544
rect 1479 1540 1483 1544
rect 1559 1540 1563 1544
rect 1647 1540 1651 1544
rect 1735 1540 1739 1544
rect 1823 1540 1827 1544
rect 1911 1540 1915 1544
rect 1999 1540 2003 1544
rect 2071 1540 2075 1544
rect 1095 1533 1099 1537
rect 1135 1532 1139 1536
rect 2119 1532 2123 1536
rect 1183 1527 1184 1531
rect 1184 1527 1187 1531
rect 1215 1527 1219 1531
rect 1255 1527 1259 1531
rect 1335 1527 1339 1531
rect 1415 1527 1419 1531
rect 1495 1527 1499 1531
rect 1583 1527 1584 1531
rect 1584 1527 1587 1531
rect 1663 1527 1667 1531
rect 1751 1527 1755 1531
rect 2019 1527 2023 1531
rect 2039 1527 2043 1531
rect 111 1516 115 1520
rect 163 1519 164 1523
rect 164 1519 167 1523
rect 183 1519 187 1523
rect 591 1519 592 1523
rect 592 1519 595 1523
rect 927 1519 931 1523
rect 963 1519 967 1523
rect 971 1519 975 1523
rect 1095 1516 1099 1520
rect 1135 1515 1139 1519
rect 135 1508 139 1512
rect 175 1508 179 1512
rect 231 1508 235 1512
rect 311 1508 315 1512
rect 391 1508 395 1512
rect 479 1508 483 1512
rect 567 1508 571 1512
rect 655 1508 659 1512
rect 743 1508 747 1512
rect 823 1508 827 1512
rect 911 1508 915 1512
rect 999 1508 1003 1512
rect 1159 1512 1163 1516
rect 1199 1512 1203 1516
rect 1247 1512 1251 1516
rect 1319 1512 1323 1516
rect 1399 1512 1403 1516
rect 1479 1512 1483 1516
rect 1559 1512 1563 1516
rect 1647 1512 1651 1516
rect 1735 1512 1739 1516
rect 1823 1512 1827 1516
rect 1911 1512 1915 1516
rect 1999 1512 2003 1516
rect 2071 1512 2075 1516
rect 2119 1515 2123 1519
rect 183 1499 187 1503
rect 435 1499 439 1503
rect 707 1499 711 1503
rect 851 1499 852 1503
rect 852 1499 855 1503
rect 927 1499 931 1503
rect 963 1499 967 1503
rect 1135 1497 1139 1501
rect 1159 1500 1163 1504
rect 1199 1500 1203 1504
rect 1239 1500 1243 1504
rect 1303 1500 1307 1504
rect 1375 1500 1379 1504
rect 1455 1500 1459 1504
rect 1543 1500 1547 1504
rect 1623 1500 1627 1504
rect 1703 1500 1707 1504
rect 1775 1500 1779 1504
rect 1847 1500 1851 1504
rect 1919 1500 1923 1504
rect 1991 1500 1995 1504
rect 2063 1500 2067 1504
rect 2119 1497 2123 1501
rect 163 1487 167 1491
rect 1799 1491 1803 1495
rect 215 1479 219 1483
rect 291 1479 295 1483
rect 535 1479 539 1483
rect 615 1479 619 1483
rect 655 1479 659 1483
rect 783 1479 787 1483
rect 819 1479 823 1483
rect 827 1479 831 1483
rect 971 1479 972 1483
rect 972 1479 975 1483
rect 979 1479 983 1483
rect 1135 1480 1139 1484
rect 1215 1483 1219 1487
rect 1255 1483 1259 1487
rect 1319 1483 1323 1487
rect 1391 1483 1395 1487
rect 1471 1483 1475 1487
rect 1535 1483 1539 1487
rect 1947 1483 1948 1487
rect 1948 1483 1951 1487
rect 2079 1483 2083 1487
rect 2087 1483 2088 1487
rect 2088 1483 2091 1487
rect 2119 1480 2123 1484
rect 135 1472 139 1476
rect 199 1472 203 1476
rect 279 1472 283 1476
rect 359 1472 363 1476
rect 439 1472 443 1476
rect 519 1472 523 1476
rect 599 1472 603 1476
rect 679 1472 683 1476
rect 767 1472 771 1476
rect 855 1472 859 1476
rect 943 1472 947 1476
rect 1031 1472 1035 1476
rect 1159 1472 1163 1476
rect 1199 1472 1203 1476
rect 1239 1472 1243 1476
rect 1303 1472 1307 1476
rect 1375 1472 1379 1476
rect 1455 1472 1459 1476
rect 1543 1472 1547 1476
rect 1623 1472 1627 1476
rect 1703 1472 1707 1476
rect 1775 1472 1779 1476
rect 1847 1472 1851 1476
rect 1919 1472 1923 1476
rect 1991 1472 1995 1476
rect 111 1464 115 1468
rect 1095 1464 1099 1468
rect 159 1459 160 1463
rect 160 1459 163 1463
rect 215 1459 219 1463
rect 431 1459 435 1463
rect 447 1459 451 1463
rect 535 1459 539 1463
rect 615 1459 619 1463
rect 707 1459 708 1463
rect 708 1459 711 1463
rect 783 1459 787 1463
rect 819 1459 823 1463
rect 979 1459 983 1463
rect 1183 1463 1184 1467
rect 1184 1463 1187 1467
rect 1071 1459 1075 1463
rect 1215 1463 1219 1467
rect 1255 1463 1259 1467
rect 1319 1463 1323 1467
rect 1391 1463 1395 1467
rect 1471 1463 1475 1467
rect 1911 1463 1915 1467
rect 2039 1471 2043 1475
rect 2063 1472 2067 1476
rect 2019 1463 2020 1467
rect 2020 1463 2023 1467
rect 2079 1463 2083 1467
rect 111 1447 115 1451
rect 135 1444 139 1448
rect 199 1444 203 1448
rect 279 1444 283 1448
rect 359 1444 363 1448
rect 439 1444 443 1448
rect 519 1444 523 1448
rect 599 1444 603 1448
rect 679 1444 683 1448
rect 767 1444 771 1448
rect 855 1444 859 1448
rect 943 1444 947 1448
rect 1031 1444 1035 1448
rect 1095 1447 1099 1451
rect 1579 1447 1583 1451
rect 1343 1439 1347 1443
rect 1399 1439 1403 1443
rect 1447 1439 1451 1443
rect 1511 1439 1515 1443
rect 1535 1439 1539 1443
rect 1615 1439 1619 1443
rect 1687 1439 1691 1443
rect 1743 1439 1747 1443
rect 2079 1439 2083 1443
rect 2087 1439 2088 1443
rect 2088 1439 2091 1443
rect 111 1429 115 1433
rect 135 1432 139 1436
rect 191 1432 195 1436
rect 263 1432 267 1436
rect 335 1432 339 1436
rect 407 1432 411 1436
rect 479 1432 483 1436
rect 551 1432 555 1436
rect 631 1432 635 1436
rect 711 1432 715 1436
rect 799 1432 803 1436
rect 887 1432 891 1436
rect 975 1432 979 1436
rect 1047 1432 1051 1436
rect 1095 1429 1099 1433
rect 1279 1432 1283 1436
rect 1327 1432 1331 1436
rect 1383 1432 1387 1436
rect 1439 1432 1443 1436
rect 1495 1432 1499 1436
rect 1551 1432 1555 1436
rect 1607 1432 1611 1436
rect 1671 1432 1675 1436
rect 1735 1432 1739 1436
rect 1807 1432 1811 1436
rect 1887 1432 1891 1436
rect 1975 1432 1979 1436
rect 2063 1432 2067 1436
rect 1135 1424 1139 1428
rect 2119 1424 2123 1428
rect 111 1412 115 1416
rect 151 1415 155 1419
rect 279 1415 283 1419
rect 291 1415 292 1419
rect 292 1415 295 1419
rect 359 1415 360 1419
rect 360 1415 363 1419
rect 527 1415 531 1419
rect 135 1404 139 1408
rect 191 1404 195 1408
rect 263 1404 267 1408
rect 335 1404 339 1408
rect 407 1404 411 1408
rect 479 1404 483 1408
rect 551 1404 555 1408
rect 631 1404 635 1408
rect 655 1415 656 1419
rect 656 1415 659 1419
rect 827 1415 828 1419
rect 828 1415 831 1419
rect 835 1415 839 1419
rect 1023 1415 1027 1419
rect 1035 1415 1039 1419
rect 1343 1419 1347 1423
rect 1399 1419 1403 1423
rect 1447 1419 1451 1423
rect 1511 1419 1515 1423
rect 1579 1419 1580 1423
rect 1580 1419 1583 1423
rect 1615 1419 1619 1423
rect 1687 1419 1691 1423
rect 1911 1419 1912 1423
rect 1912 1419 1915 1423
rect 2015 1419 2019 1423
rect 2079 1419 2083 1423
rect 1095 1412 1099 1416
rect 159 1395 160 1399
rect 160 1395 163 1399
rect 203 1395 207 1399
rect 279 1395 283 1399
rect 447 1395 451 1399
rect 599 1395 603 1399
rect 711 1404 715 1408
rect 799 1404 803 1408
rect 887 1404 891 1408
rect 975 1404 979 1408
rect 1047 1404 1051 1408
rect 1135 1407 1139 1411
rect 1279 1404 1283 1408
rect 1327 1404 1331 1408
rect 1383 1404 1387 1408
rect 1439 1404 1443 1408
rect 1495 1404 1499 1408
rect 1551 1404 1555 1408
rect 1607 1404 1611 1408
rect 1671 1404 1675 1408
rect 1735 1404 1739 1408
rect 1807 1404 1811 1408
rect 1887 1404 1891 1408
rect 1975 1404 1979 1408
rect 2063 1404 2067 1408
rect 2119 1407 2123 1411
rect 835 1395 839 1399
rect 951 1395 955 1399
rect 1035 1395 1039 1399
rect 1071 1395 1072 1399
rect 1072 1395 1075 1399
rect 359 1387 363 1391
rect 1135 1385 1139 1389
rect 1335 1388 1339 1392
rect 1375 1388 1379 1392
rect 1415 1388 1419 1392
rect 1455 1388 1459 1392
rect 1495 1388 1499 1392
rect 1535 1388 1539 1392
rect 1583 1388 1587 1392
rect 1647 1388 1651 1392
rect 1719 1388 1723 1392
rect 1807 1388 1811 1392
rect 1895 1388 1899 1392
rect 1991 1388 1995 1392
rect 2071 1388 2075 1392
rect 2119 1385 2123 1389
rect 151 1375 155 1379
rect 251 1375 255 1379
rect 135 1368 139 1372
rect 175 1368 179 1372
rect 239 1368 243 1372
rect 303 1368 307 1372
rect 383 1375 387 1379
rect 455 1375 459 1379
rect 511 1375 515 1379
rect 527 1375 528 1379
rect 528 1375 531 1379
rect 663 1375 667 1379
rect 719 1375 723 1379
rect 731 1375 735 1379
rect 807 1375 808 1379
rect 808 1375 811 1379
rect 891 1375 895 1379
rect 1023 1375 1024 1379
rect 1024 1375 1027 1379
rect 359 1367 363 1371
rect 367 1368 371 1372
rect 439 1368 443 1372
rect 503 1368 507 1372
rect 575 1368 579 1372
rect 647 1368 651 1372
rect 711 1368 715 1372
rect 783 1368 787 1372
rect 855 1368 859 1372
rect 927 1368 931 1372
rect 999 1368 1003 1372
rect 1047 1368 1051 1372
rect 1135 1368 1139 1372
rect 1391 1371 1395 1375
rect 1423 1371 1427 1375
rect 1431 1371 1435 1375
rect 1483 1371 1484 1375
rect 1484 1371 1487 1375
rect 1503 1371 1507 1375
rect 1543 1371 1547 1375
rect 1663 1371 1667 1375
rect 1919 1379 1923 1383
rect 1743 1371 1744 1375
rect 1744 1371 1747 1375
rect 2087 1371 2091 1375
rect 2095 1371 2096 1375
rect 2096 1371 2099 1375
rect 2119 1368 2123 1372
rect 111 1360 115 1364
rect 1095 1360 1099 1364
rect 159 1355 160 1359
rect 160 1355 163 1359
rect 203 1355 204 1359
rect 204 1355 207 1359
rect 251 1355 255 1359
rect 375 1355 379 1359
rect 383 1355 387 1359
rect 455 1355 459 1359
rect 511 1355 515 1359
rect 599 1355 600 1359
rect 600 1355 603 1359
rect 663 1355 667 1359
rect 719 1355 723 1359
rect 891 1355 895 1359
rect 951 1355 952 1359
rect 952 1355 955 1359
rect 1335 1360 1339 1364
rect 1375 1360 1379 1364
rect 1415 1360 1419 1364
rect 1455 1360 1459 1364
rect 1495 1360 1499 1364
rect 1535 1360 1539 1364
rect 1583 1360 1587 1364
rect 1647 1360 1651 1364
rect 1719 1360 1723 1364
rect 1807 1360 1811 1364
rect 1895 1360 1899 1364
rect 1991 1360 1995 1364
rect 2071 1360 2075 1364
rect 1087 1355 1091 1359
rect 1391 1351 1395 1355
rect 1423 1351 1427 1355
rect 1503 1351 1507 1355
rect 1543 1351 1547 1355
rect 1591 1351 1595 1355
rect 1663 1351 1667 1355
rect 1919 1351 1920 1355
rect 1920 1351 1923 1355
rect 2015 1351 2016 1355
rect 2016 1351 2019 1355
rect 2087 1351 2091 1355
rect 111 1343 115 1347
rect 135 1340 139 1344
rect 175 1340 179 1344
rect 239 1340 243 1344
rect 303 1340 307 1344
rect 367 1340 371 1344
rect 439 1340 443 1344
rect 503 1340 507 1344
rect 575 1340 579 1344
rect 647 1340 651 1344
rect 711 1340 715 1344
rect 783 1340 787 1344
rect 855 1340 859 1344
rect 927 1340 931 1344
rect 999 1340 1003 1344
rect 1047 1340 1051 1344
rect 1095 1343 1099 1347
rect 1483 1343 1487 1347
rect 1087 1331 1091 1335
rect 1431 1331 1432 1335
rect 1432 1331 1435 1335
rect 1775 1331 1779 1335
rect 1847 1331 1851 1335
rect 1911 1331 1915 1335
rect 1975 1331 1979 1335
rect 2039 1331 2043 1335
rect 2047 1331 2048 1335
rect 2048 1331 2051 1335
rect 2095 1331 2096 1335
rect 2096 1331 2099 1335
rect 111 1317 115 1321
rect 135 1320 139 1324
rect 175 1320 179 1324
rect 215 1320 219 1324
rect 255 1320 259 1324
rect 319 1320 323 1324
rect 391 1320 395 1324
rect 463 1320 467 1324
rect 543 1320 547 1324
rect 623 1320 627 1324
rect 703 1320 707 1324
rect 783 1320 787 1324
rect 863 1320 867 1324
rect 943 1320 947 1324
rect 1023 1320 1027 1324
rect 1159 1324 1163 1328
rect 1223 1324 1227 1328
rect 1311 1324 1315 1328
rect 1407 1324 1411 1328
rect 1503 1324 1507 1328
rect 1599 1324 1603 1328
rect 1679 1324 1683 1328
rect 1759 1324 1763 1328
rect 1831 1324 1835 1328
rect 1895 1324 1899 1328
rect 1959 1324 1963 1328
rect 2023 1324 2027 1328
rect 2071 1324 2075 1328
rect 1095 1317 1099 1321
rect 1135 1316 1139 1320
rect 2119 1316 2123 1320
rect 111 1300 115 1304
rect 191 1303 195 1307
rect 231 1303 235 1307
rect 343 1311 347 1315
rect 1331 1311 1335 1315
rect 1591 1311 1595 1315
rect 1767 1311 1771 1315
rect 1775 1311 1779 1315
rect 1847 1311 1851 1315
rect 1911 1311 1915 1315
rect 1975 1311 1979 1315
rect 2039 1311 2043 1315
rect 2095 1311 2096 1315
rect 2096 1311 2099 1315
rect 279 1303 280 1307
rect 280 1303 283 1307
rect 359 1303 363 1307
rect 639 1303 643 1307
rect 719 1303 723 1307
rect 731 1303 732 1307
rect 732 1303 735 1307
rect 807 1303 808 1307
rect 808 1303 811 1307
rect 1095 1300 1099 1304
rect 1135 1299 1139 1303
rect 135 1292 139 1296
rect 175 1292 179 1296
rect 215 1292 219 1296
rect 255 1292 259 1296
rect 319 1292 323 1296
rect 391 1292 395 1296
rect 463 1292 467 1296
rect 543 1292 547 1296
rect 623 1292 627 1296
rect 703 1292 707 1296
rect 783 1292 787 1296
rect 863 1292 867 1296
rect 943 1292 947 1296
rect 1023 1292 1027 1296
rect 1159 1296 1163 1300
rect 1223 1296 1227 1300
rect 1311 1296 1315 1300
rect 1407 1296 1411 1300
rect 1503 1296 1507 1300
rect 1599 1296 1603 1300
rect 1679 1296 1683 1300
rect 1759 1296 1763 1300
rect 1831 1296 1835 1300
rect 1895 1296 1899 1300
rect 1959 1296 1963 1300
rect 2023 1296 2027 1300
rect 2071 1296 2075 1300
rect 2119 1299 2123 1303
rect 159 1283 160 1287
rect 160 1283 163 1287
rect 191 1283 195 1287
rect 231 1283 235 1287
rect 343 1283 344 1287
rect 344 1283 347 1287
rect 375 1275 379 1279
rect 551 1283 555 1287
rect 639 1283 643 1287
rect 719 1283 723 1287
rect 1071 1283 1075 1287
rect 1135 1281 1139 1285
rect 1175 1284 1179 1288
rect 1231 1284 1235 1288
rect 1303 1284 1307 1288
rect 1391 1284 1395 1288
rect 1479 1284 1483 1288
rect 1567 1284 1571 1288
rect 1655 1284 1659 1288
rect 1743 1284 1747 1288
rect 1831 1284 1835 1288
rect 1919 1284 1923 1288
rect 2007 1284 2011 1288
rect 2071 1284 2075 1288
rect 2119 1281 2123 1285
rect 191 1259 195 1263
rect 231 1259 235 1263
rect 279 1267 283 1271
rect 575 1267 579 1271
rect 1135 1264 1139 1268
rect 1199 1267 1200 1271
rect 1200 1267 1203 1271
rect 1411 1267 1415 1271
rect 1671 1267 1675 1271
rect 2047 1267 2051 1271
rect 135 1252 139 1256
rect 175 1252 179 1256
rect 215 1252 219 1256
rect 255 1252 259 1256
rect 111 1244 115 1248
rect 599 1259 603 1263
rect 703 1259 707 1263
rect 815 1259 819 1263
rect 1007 1259 1011 1263
rect 1015 1259 1019 1263
rect 2119 1264 2123 1268
rect 319 1252 323 1256
rect 399 1252 403 1256
rect 487 1252 491 1256
rect 583 1252 587 1256
rect 687 1252 691 1256
rect 799 1252 803 1256
rect 919 1252 923 1256
rect 1047 1252 1051 1256
rect 1175 1256 1179 1260
rect 1231 1256 1235 1260
rect 1303 1256 1307 1260
rect 1391 1256 1395 1260
rect 1479 1256 1483 1260
rect 1567 1256 1571 1260
rect 1655 1256 1659 1260
rect 1743 1256 1747 1260
rect 1831 1256 1835 1260
rect 1919 1256 1923 1260
rect 2007 1256 2011 1260
rect 2071 1256 2075 1260
rect 1095 1244 1099 1248
rect 1331 1247 1332 1251
rect 1332 1247 1335 1251
rect 1591 1247 1592 1251
rect 1592 1247 1595 1251
rect 1995 1247 1999 1251
rect 2095 1247 2096 1251
rect 2096 1247 2099 1251
rect 191 1239 195 1243
rect 231 1239 235 1243
rect 379 1239 383 1243
rect 551 1239 555 1243
rect 599 1239 603 1243
rect 703 1239 707 1243
rect 815 1239 819 1243
rect 1015 1239 1019 1243
rect 1071 1239 1072 1243
rect 1072 1239 1075 1243
rect 1767 1239 1771 1243
rect 111 1227 115 1231
rect 135 1224 139 1228
rect 175 1224 179 1228
rect 215 1224 219 1228
rect 255 1224 259 1228
rect 319 1224 323 1228
rect 399 1224 403 1228
rect 487 1224 491 1228
rect 583 1224 587 1228
rect 687 1224 691 1228
rect 799 1224 803 1228
rect 919 1224 923 1228
rect 1047 1224 1051 1228
rect 1095 1227 1099 1231
rect 1315 1231 1319 1235
rect 1343 1223 1347 1227
rect 1391 1223 1395 1227
rect 1411 1223 1415 1227
rect 1459 1231 1463 1235
rect 1671 1231 1675 1235
rect 1575 1223 1579 1227
rect 1687 1223 1691 1227
rect 1751 1223 1755 1227
rect 1807 1223 1811 1227
rect 1855 1223 1859 1227
rect 1919 1223 1923 1227
rect 2007 1223 2011 1227
rect 2087 1223 2091 1227
rect 1287 1216 1291 1220
rect 1327 1216 1331 1220
rect 1375 1216 1379 1220
rect 1431 1216 1435 1220
rect 1495 1216 1499 1220
rect 1559 1216 1563 1220
rect 1623 1216 1627 1220
rect 1679 1216 1683 1220
rect 1735 1216 1739 1220
rect 1791 1216 1795 1220
rect 1847 1216 1851 1220
rect 1903 1216 1907 1220
rect 1967 1216 1971 1220
rect 2031 1216 2035 1220
rect 2071 1216 2075 1220
rect 111 1205 115 1209
rect 271 1208 275 1212
rect 311 1208 315 1212
rect 351 1208 355 1212
rect 399 1208 403 1212
rect 447 1208 451 1212
rect 495 1208 499 1212
rect 551 1208 555 1212
rect 607 1208 611 1212
rect 671 1208 675 1212
rect 743 1208 747 1212
rect 815 1208 819 1212
rect 895 1208 899 1212
rect 983 1208 987 1212
rect 1095 1205 1099 1209
rect 1135 1208 1139 1212
rect 2119 1208 2123 1212
rect 111 1188 115 1192
rect 423 1199 427 1203
rect 1315 1203 1316 1207
rect 1316 1203 1319 1207
rect 1343 1203 1347 1207
rect 1391 1203 1395 1207
rect 1459 1203 1460 1207
rect 1460 1203 1463 1207
rect 1515 1203 1519 1207
rect 1575 1203 1579 1207
rect 1671 1203 1675 1207
rect 1687 1203 1691 1207
rect 1751 1203 1755 1207
rect 1807 1203 1811 1207
rect 1855 1203 1859 1207
rect 1919 1203 1923 1207
rect 1995 1203 1996 1207
rect 1996 1203 1999 1207
rect 2079 1203 2083 1207
rect 2087 1203 2091 1207
rect 327 1191 331 1195
rect 359 1191 363 1195
rect 463 1191 467 1195
rect 511 1191 515 1195
rect 567 1191 571 1195
rect 575 1191 576 1195
rect 576 1191 579 1195
rect 1007 1191 1008 1195
rect 1008 1191 1011 1195
rect 1095 1188 1099 1192
rect 1135 1191 1139 1195
rect 1287 1188 1291 1192
rect 1327 1188 1331 1192
rect 1375 1188 1379 1192
rect 1431 1188 1435 1192
rect 1495 1188 1499 1192
rect 1559 1188 1563 1192
rect 1623 1188 1627 1192
rect 1679 1188 1683 1192
rect 1735 1188 1739 1192
rect 1791 1188 1795 1192
rect 1847 1188 1851 1192
rect 1903 1188 1907 1192
rect 1967 1188 1971 1192
rect 2031 1188 2035 1192
rect 2071 1188 2075 1192
rect 2119 1191 2123 1195
rect 271 1180 275 1184
rect 311 1180 315 1184
rect 351 1180 355 1184
rect 399 1180 403 1184
rect 447 1180 451 1184
rect 495 1180 499 1184
rect 551 1180 555 1184
rect 607 1180 611 1184
rect 671 1180 675 1184
rect 743 1180 747 1184
rect 815 1180 819 1184
rect 895 1180 899 1184
rect 983 1180 987 1184
rect 327 1171 331 1175
rect 359 1171 363 1175
rect 379 1171 380 1175
rect 380 1171 383 1175
rect 423 1171 424 1175
rect 424 1171 427 1175
rect 463 1171 467 1175
rect 511 1171 515 1175
rect 971 1171 975 1175
rect 1135 1173 1139 1177
rect 1159 1176 1163 1180
rect 1207 1176 1211 1180
rect 1279 1176 1283 1180
rect 1351 1176 1355 1180
rect 1423 1176 1427 1180
rect 1487 1176 1491 1180
rect 1559 1176 1563 1180
rect 1631 1176 1635 1180
rect 1711 1176 1715 1180
rect 1799 1176 1803 1180
rect 1887 1176 1891 1180
rect 1983 1176 1987 1180
rect 2071 1176 2075 1180
rect 2119 1173 2123 1177
rect 699 1163 703 1167
rect 567 1155 571 1159
rect 455 1147 459 1151
rect 495 1147 499 1151
rect 543 1147 547 1151
rect 591 1147 595 1151
rect 631 1147 635 1151
rect 663 1155 667 1159
rect 1135 1156 1139 1160
rect 735 1147 739 1151
rect 791 1147 795 1151
rect 847 1147 851 1151
rect 903 1147 907 1151
rect 1023 1147 1027 1151
rect 1063 1147 1067 1151
rect 1371 1159 1375 1163
rect 1583 1159 1584 1163
rect 1584 1159 1587 1163
rect 2007 1159 2008 1163
rect 2008 1159 2011 1163
rect 2095 1159 2096 1163
rect 2096 1159 2099 1163
rect 2119 1156 2123 1160
rect 1159 1148 1163 1152
rect 1207 1148 1211 1152
rect 1279 1148 1283 1152
rect 1351 1148 1355 1152
rect 1423 1148 1427 1152
rect 1487 1148 1491 1152
rect 1559 1148 1563 1152
rect 1631 1148 1635 1152
rect 1711 1148 1715 1152
rect 1799 1148 1803 1152
rect 1887 1148 1891 1152
rect 1983 1148 1987 1152
rect 2071 1148 2075 1152
rect 399 1140 403 1144
rect 439 1140 443 1144
rect 479 1140 483 1144
rect 527 1140 531 1144
rect 575 1140 579 1144
rect 623 1140 627 1144
rect 671 1140 675 1144
rect 719 1140 723 1144
rect 775 1140 779 1144
rect 831 1140 835 1144
rect 887 1140 891 1144
rect 943 1140 947 1144
rect 1007 1140 1011 1144
rect 1047 1140 1051 1144
rect 1515 1139 1516 1143
rect 1516 1139 1519 1143
rect 111 1132 115 1136
rect 1095 1132 1099 1136
rect 427 1127 428 1131
rect 428 1127 431 1131
rect 455 1127 459 1131
rect 495 1127 499 1131
rect 543 1127 547 1131
rect 591 1127 595 1131
rect 631 1127 635 1131
rect 699 1127 700 1131
rect 700 1127 703 1131
rect 735 1127 739 1131
rect 791 1127 795 1131
rect 847 1127 851 1131
rect 903 1127 907 1131
rect 971 1127 972 1131
rect 972 1127 975 1131
rect 1055 1127 1059 1131
rect 1063 1127 1067 1131
rect 1687 1131 1691 1135
rect 2003 1139 2007 1143
rect 2079 1139 2083 1143
rect 1583 1123 1587 1127
rect 111 1115 115 1119
rect 399 1112 403 1116
rect 439 1112 443 1116
rect 479 1112 483 1116
rect 527 1112 531 1116
rect 575 1112 579 1116
rect 623 1112 627 1116
rect 671 1112 675 1116
rect 719 1112 723 1116
rect 775 1112 779 1116
rect 831 1112 835 1116
rect 887 1112 891 1116
rect 943 1112 947 1116
rect 1007 1112 1011 1116
rect 1047 1112 1051 1116
rect 1095 1115 1099 1119
rect 1287 1115 1291 1119
rect 1327 1115 1331 1119
rect 1371 1115 1372 1119
rect 1372 1115 1375 1119
rect 1479 1115 1483 1119
rect 1583 1115 1587 1119
rect 1671 1115 1675 1119
rect 1767 1115 1771 1119
rect 1871 1115 1875 1119
rect 1983 1115 1984 1119
rect 1984 1115 1987 1119
rect 2095 1115 2096 1119
rect 2096 1115 2099 1119
rect 1191 1108 1195 1112
rect 1271 1108 1275 1112
rect 1343 1108 1347 1112
rect 1415 1108 1419 1112
rect 1487 1108 1491 1112
rect 1567 1108 1571 1112
rect 1655 1108 1659 1112
rect 1751 1108 1755 1112
rect 1855 1108 1859 1112
rect 1959 1108 1963 1112
rect 2071 1108 2075 1112
rect 111 1097 115 1101
rect 159 1100 163 1104
rect 199 1100 203 1104
rect 255 1100 259 1104
rect 319 1100 323 1104
rect 399 1100 403 1104
rect 479 1100 483 1104
rect 559 1100 563 1104
rect 639 1100 643 1104
rect 711 1100 715 1104
rect 783 1100 787 1104
rect 855 1100 859 1104
rect 927 1100 931 1104
rect 999 1100 1003 1104
rect 1047 1100 1051 1104
rect 1095 1097 1099 1101
rect 1135 1100 1139 1104
rect 1287 1095 1291 1099
rect 1371 1095 1372 1099
rect 1372 1095 1375 1099
rect 1471 1095 1475 1099
rect 1495 1095 1499 1099
rect 1583 1095 1587 1099
rect 1671 1095 1675 1099
rect 1767 1095 1771 1099
rect 1871 1095 1875 1099
rect 2003 1099 2007 1103
rect 2119 1100 2123 1104
rect 2095 1095 2096 1099
rect 2096 1095 2099 1099
rect 111 1080 115 1084
rect 187 1083 188 1087
rect 188 1083 191 1087
rect 207 1083 211 1087
rect 663 1083 664 1087
rect 664 1083 667 1087
rect 1015 1083 1019 1087
rect 1023 1083 1024 1087
rect 1024 1083 1027 1087
rect 1087 1083 1091 1087
rect 1095 1080 1099 1084
rect 1135 1083 1139 1087
rect 1191 1080 1195 1084
rect 1271 1080 1275 1084
rect 1343 1080 1347 1084
rect 1415 1080 1419 1084
rect 1487 1080 1491 1084
rect 1567 1080 1571 1084
rect 1655 1080 1659 1084
rect 1751 1080 1755 1084
rect 1855 1080 1859 1084
rect 1959 1080 1963 1084
rect 2071 1080 2075 1084
rect 2119 1083 2123 1087
rect 159 1072 163 1076
rect 199 1072 203 1076
rect 255 1072 259 1076
rect 319 1072 323 1076
rect 399 1072 403 1076
rect 479 1072 483 1076
rect 559 1072 563 1076
rect 639 1072 643 1076
rect 711 1072 715 1076
rect 783 1072 787 1076
rect 855 1072 859 1076
rect 927 1072 931 1076
rect 999 1072 1003 1076
rect 1047 1072 1051 1076
rect 207 1063 211 1067
rect 883 1063 884 1067
rect 884 1063 887 1067
rect 1015 1063 1019 1067
rect 1055 1063 1059 1067
rect 1135 1065 1139 1069
rect 1159 1068 1163 1072
rect 1199 1068 1203 1072
rect 1247 1068 1251 1072
rect 1303 1068 1307 1072
rect 1351 1068 1355 1072
rect 1399 1068 1403 1072
rect 1455 1068 1459 1072
rect 1511 1068 1515 1072
rect 1583 1068 1587 1072
rect 1663 1068 1667 1072
rect 1759 1068 1763 1072
rect 1863 1068 1867 1072
rect 1967 1068 1971 1072
rect 2071 1068 2075 1072
rect 2119 1065 2123 1069
rect 167 1055 171 1059
rect 187 1047 191 1051
rect 427 1055 431 1059
rect 603 1055 607 1059
rect 1887 1059 1891 1063
rect 1135 1048 1139 1052
rect 1215 1051 1219 1055
rect 1223 1051 1224 1055
rect 1224 1051 1227 1055
rect 1319 1051 1323 1055
rect 1327 1051 1328 1055
rect 1328 1051 1331 1055
rect 1415 1051 1419 1055
rect 1427 1051 1428 1055
rect 1428 1051 1431 1055
rect 1479 1051 1480 1055
rect 1480 1051 1483 1055
rect 1599 1051 1603 1055
rect 1679 1051 1683 1055
rect 1991 1051 1992 1055
rect 1992 1051 1995 1055
rect 2047 1051 2051 1055
rect 2119 1048 2123 1052
rect 191 1039 195 1043
rect 231 1039 235 1043
rect 271 1039 275 1043
rect 399 1039 403 1043
rect 463 1039 467 1043
rect 547 1039 551 1043
rect 555 1039 559 1043
rect 611 1039 615 1043
rect 735 1039 739 1043
rect 1159 1040 1163 1044
rect 1199 1040 1203 1044
rect 1247 1040 1251 1044
rect 1303 1040 1307 1044
rect 1351 1040 1355 1044
rect 1399 1040 1403 1044
rect 1455 1040 1459 1044
rect 1471 1039 1475 1043
rect 135 1032 139 1036
rect 175 1032 179 1036
rect 215 1032 219 1036
rect 255 1032 259 1036
rect 319 1032 323 1036
rect 383 1032 387 1036
rect 447 1032 451 1036
rect 511 1032 515 1036
rect 575 1032 579 1036
rect 631 1032 635 1036
rect 687 1032 691 1036
rect 743 1032 747 1036
rect 799 1032 803 1036
rect 863 1032 867 1036
rect 1087 1031 1091 1035
rect 1215 1031 1219 1035
rect 1267 1031 1271 1035
rect 1319 1031 1323 1035
rect 1371 1031 1375 1035
rect 1415 1031 1419 1035
rect 1495 1031 1499 1035
rect 1511 1040 1515 1044
rect 1583 1040 1587 1044
rect 1663 1040 1667 1044
rect 1759 1040 1763 1044
rect 1863 1040 1867 1044
rect 1967 1040 1971 1044
rect 2071 1040 2075 1044
rect 1599 1031 1603 1035
rect 1887 1031 1888 1035
rect 1888 1031 1891 1035
rect 2047 1031 2051 1035
rect 2095 1031 2096 1035
rect 2096 1031 2099 1035
rect 111 1024 115 1028
rect 1095 1024 1099 1028
rect 160 1019 164 1023
rect 191 1019 195 1023
rect 231 1019 235 1023
rect 271 1019 275 1023
rect 291 1019 295 1023
rect 399 1019 403 1023
rect 463 1019 467 1023
rect 555 1019 559 1023
rect 603 1019 604 1023
rect 604 1019 607 1023
rect 735 1019 739 1023
rect 883 1019 887 1023
rect 111 1007 115 1011
rect 135 1004 139 1008
rect 175 1004 179 1008
rect 215 1004 219 1008
rect 255 1004 259 1008
rect 319 1004 323 1008
rect 383 1004 387 1008
rect 447 1004 451 1008
rect 511 1004 515 1008
rect 575 1004 579 1008
rect 631 1004 635 1008
rect 687 1004 691 1008
rect 743 1004 747 1008
rect 799 1004 803 1008
rect 863 1004 867 1008
rect 1095 1007 1099 1011
rect 1215 1007 1219 1011
rect 1223 1007 1224 1011
rect 1224 1007 1227 1011
rect 1311 1007 1315 1011
rect 1359 1007 1363 1011
rect 1399 1007 1403 1011
rect 1427 1007 1431 1011
rect 1591 1007 1595 1011
rect 1655 1007 1659 1011
rect 1679 1011 1683 1015
rect 1991 1015 1995 1019
rect 1159 1000 1163 1004
rect 1199 1000 1203 1004
rect 1239 1000 1243 1004
rect 1295 1000 1299 1004
rect 1351 1000 1355 1004
rect 1407 1000 1411 1004
rect 1463 1000 1467 1004
rect 1519 1000 1523 1004
rect 1575 1000 1579 1004
rect 1639 1000 1643 1004
rect 1895 1007 1899 1011
rect 1711 1000 1715 1004
rect 111 985 115 989
rect 135 988 139 992
rect 175 988 179 992
rect 223 988 227 992
rect 279 988 283 992
rect 343 988 347 992
rect 407 988 411 992
rect 471 988 475 992
rect 527 988 531 992
rect 583 988 587 992
rect 631 988 635 992
rect 687 988 691 992
rect 743 988 747 992
rect 799 988 803 992
rect 1135 992 1139 996
rect 1095 985 1099 989
rect 1207 987 1211 991
rect 1215 987 1219 991
rect 1267 987 1268 991
rect 1268 987 1271 991
rect 1311 987 1315 991
rect 1359 987 1363 991
rect 1483 987 1487 991
rect 1791 1000 1795 1004
rect 1879 1000 1883 1004
rect 1967 1000 1971 1004
rect 1591 987 1595 991
rect 1655 987 1659 991
rect 1779 987 1783 991
rect 1895 987 1899 991
rect 1983 987 1987 991
rect 2063 1000 2067 1004
rect 2119 992 2123 996
rect 111 968 115 972
rect 303 979 307 983
rect 183 971 187 975
rect 359 971 363 975
rect 419 971 423 975
rect 427 971 431 975
rect 539 971 543 975
rect 547 971 551 975
rect 607 971 608 975
rect 608 971 611 975
rect 1135 975 1139 979
rect 1095 968 1099 972
rect 1159 972 1163 976
rect 1199 972 1203 976
rect 1239 972 1243 976
rect 1295 972 1299 976
rect 1351 972 1355 976
rect 1407 972 1411 976
rect 1463 972 1467 976
rect 1519 972 1523 976
rect 1575 972 1579 976
rect 1639 972 1643 976
rect 1711 972 1715 976
rect 1791 972 1795 976
rect 1879 972 1883 976
rect 1967 972 1971 976
rect 2063 972 2067 976
rect 2119 975 2123 979
rect 135 960 139 964
rect 175 960 179 964
rect 223 960 227 964
rect 279 960 283 964
rect 343 960 347 964
rect 407 960 411 964
rect 471 960 475 964
rect 527 960 531 964
rect 583 960 587 964
rect 631 960 635 964
rect 687 960 691 964
rect 743 960 747 964
rect 799 960 803 964
rect 183 951 187 955
rect 291 951 295 955
rect 303 951 304 955
rect 304 951 307 955
rect 359 951 363 955
rect 419 951 423 955
rect 483 951 487 955
rect 539 951 543 955
rect 715 943 719 947
rect 1135 949 1139 953
rect 1159 952 1163 956
rect 1207 952 1211 956
rect 1287 952 1291 956
rect 1375 952 1379 956
rect 1455 952 1459 956
rect 1535 952 1539 956
rect 1615 952 1619 956
rect 1687 952 1691 956
rect 1751 952 1755 956
rect 1815 952 1819 956
rect 1879 952 1883 956
rect 1951 952 1955 956
rect 2023 952 2027 956
rect 2071 952 2075 956
rect 2119 949 2123 953
rect 1839 943 1843 947
rect 1135 932 1139 936
rect 1215 935 1219 939
rect 1391 935 1395 939
rect 1399 935 1400 939
rect 1400 935 1403 939
rect 1551 935 1555 939
rect 1607 935 1611 939
rect 1887 935 1891 939
rect 1967 935 1971 939
rect 2039 935 2043 939
rect 2047 935 2048 939
rect 2048 935 2051 939
rect 2095 935 2096 939
rect 2096 935 2099 939
rect 319 927 323 931
rect 367 927 371 931
rect 415 927 419 931
rect 427 927 428 931
rect 428 927 431 931
rect 523 927 527 931
rect 575 927 579 931
rect 639 927 643 931
rect 647 927 648 931
rect 648 927 651 931
rect 767 927 771 931
rect 831 927 835 931
rect 895 927 899 931
rect 959 927 963 931
rect 967 927 968 931
rect 968 927 971 931
rect 1063 927 1067 931
rect 2119 932 2123 936
rect 263 920 267 924
rect 303 920 307 924
rect 351 920 355 924
rect 399 920 403 924
rect 455 920 459 924
rect 511 920 515 924
rect 567 920 571 924
rect 623 920 627 924
rect 687 920 691 924
rect 751 920 755 924
rect 815 920 819 924
rect 879 920 883 924
rect 943 920 947 924
rect 1007 920 1011 924
rect 1047 920 1051 924
rect 1159 924 1163 928
rect 1207 924 1211 928
rect 1287 924 1291 928
rect 1375 924 1379 928
rect 1455 924 1459 928
rect 1535 924 1539 928
rect 1615 924 1619 928
rect 1687 924 1691 928
rect 1751 924 1755 928
rect 1815 924 1819 928
rect 1879 924 1883 928
rect 1951 924 1955 928
rect 2023 924 2027 928
rect 2071 924 2075 928
rect 111 912 115 916
rect 1095 912 1099 916
rect 1215 915 1219 919
rect 1223 915 1227 919
rect 1267 915 1271 919
rect 1391 915 1395 919
rect 1483 915 1484 919
rect 1484 915 1487 919
rect 1551 915 1555 919
rect 1779 915 1780 919
rect 1780 915 1783 919
rect 1839 915 1840 919
rect 1840 915 1843 919
rect 1887 915 1891 919
rect 1967 915 1971 919
rect 2039 915 2043 919
rect 291 907 292 911
rect 292 907 295 911
rect 319 907 323 911
rect 367 907 371 911
rect 415 907 419 911
rect 483 907 484 911
rect 484 907 487 911
rect 523 907 527 911
rect 575 907 579 911
rect 639 907 643 911
rect 715 907 716 911
rect 716 907 719 911
rect 767 907 771 911
rect 831 907 835 911
rect 895 907 899 911
rect 959 907 963 911
rect 1055 907 1059 911
rect 1063 907 1067 911
rect 111 895 115 899
rect 263 892 267 896
rect 303 892 307 896
rect 351 892 355 896
rect 399 892 403 896
rect 455 892 459 896
rect 511 892 515 896
rect 567 892 571 896
rect 623 892 627 896
rect 687 892 691 896
rect 751 892 755 896
rect 815 892 819 896
rect 879 892 883 896
rect 943 892 947 896
rect 1007 892 1011 896
rect 1047 892 1051 896
rect 1095 895 1099 899
rect 1335 895 1339 899
rect 1379 895 1383 899
rect 1387 895 1391 899
rect 1599 895 1603 899
rect 1607 895 1608 899
rect 1608 895 1611 899
rect 1759 895 1763 899
rect 1807 895 1811 899
rect 1903 895 1907 899
rect 1967 895 1971 899
rect 2039 895 2043 899
rect 2047 895 2048 899
rect 2048 895 2051 899
rect 2095 895 2096 899
rect 2096 895 2099 899
rect 1239 888 1243 892
rect 1319 888 1323 892
rect 1407 888 1411 892
rect 1495 888 1499 892
rect 1583 888 1587 892
rect 1663 888 1667 892
rect 1743 888 1747 892
rect 1815 888 1819 892
rect 1887 888 1891 892
rect 1951 888 1955 892
rect 2023 888 2027 892
rect 2071 888 2075 892
rect 111 873 115 877
rect 303 876 307 880
rect 351 876 355 880
rect 415 876 419 880
rect 479 876 483 880
rect 551 876 555 880
rect 623 876 627 880
rect 695 876 699 880
rect 767 876 771 880
rect 831 876 835 880
rect 887 876 891 880
rect 943 876 947 880
rect 1007 876 1011 880
rect 1047 876 1051 880
rect 1135 880 1139 884
rect 2119 880 2123 884
rect 1095 873 1099 877
rect 1267 875 1268 879
rect 1268 875 1271 879
rect 1335 875 1339 879
rect 1379 875 1383 879
rect 1483 875 1487 879
rect 1599 875 1603 879
rect 1735 875 1739 879
rect 1759 875 1763 879
rect 1895 875 1899 879
rect 1903 875 1907 879
rect 1967 875 1971 879
rect 2039 875 2043 879
rect 2095 875 2096 879
rect 2096 875 2099 879
rect 967 867 971 871
rect 111 856 115 860
rect 311 859 315 863
rect 303 848 307 852
rect 351 848 355 852
rect 567 859 571 863
rect 639 859 643 863
rect 647 859 648 863
rect 648 859 651 863
rect 731 859 735 863
rect 935 859 939 863
rect 1055 859 1059 863
rect 1135 863 1139 867
rect 1095 856 1099 860
rect 1239 860 1243 864
rect 1319 860 1323 864
rect 1407 860 1411 864
rect 1495 860 1499 864
rect 1583 860 1587 864
rect 1663 860 1667 864
rect 1743 860 1747 864
rect 1815 860 1819 864
rect 1887 860 1891 864
rect 1951 860 1955 864
rect 2023 860 2027 864
rect 2071 860 2075 864
rect 2119 863 2123 867
rect 415 848 419 852
rect 479 848 483 852
rect 551 848 555 852
rect 623 848 627 852
rect 695 848 699 852
rect 767 848 771 852
rect 831 848 835 852
rect 887 848 891 852
rect 943 848 947 852
rect 1007 848 1011 852
rect 1047 848 1051 852
rect 1135 845 1139 849
rect 1159 848 1163 852
rect 1247 848 1251 852
rect 1359 848 1363 852
rect 1455 848 1459 852
rect 1543 848 1547 852
rect 1631 848 1635 852
rect 1711 848 1715 852
rect 1783 848 1787 852
rect 1855 848 1859 852
rect 1935 848 1939 852
rect 2015 848 2019 852
rect 2071 848 2075 852
rect 2119 845 2123 849
rect 291 831 295 835
rect 507 839 508 843
rect 508 839 511 843
rect 567 839 571 843
rect 639 839 643 843
rect 731 839 735 843
rect 755 831 759 835
rect 1055 839 1059 843
rect 1063 839 1067 843
rect 304 819 308 823
rect 335 819 339 823
rect 583 819 587 823
rect 663 819 667 823
rect 671 819 672 823
rect 672 819 675 823
rect 815 819 819 823
rect 935 827 939 831
rect 1135 828 1139 832
rect 1263 831 1267 835
rect 1375 831 1379 835
rect 1387 831 1388 835
rect 1388 831 1391 835
rect 1463 831 1467 835
rect 1559 831 1563 835
rect 1807 831 1808 835
rect 1808 831 1811 835
rect 1819 831 1823 835
rect 2119 828 2123 832
rect 887 819 888 823
rect 888 819 891 823
rect 1071 819 1072 823
rect 1072 819 1075 823
rect 1159 820 1163 824
rect 1247 820 1251 824
rect 1359 820 1363 824
rect 1455 820 1459 824
rect 1543 820 1547 824
rect 1631 820 1635 824
rect 1711 820 1715 824
rect 1783 820 1787 824
rect 1855 820 1859 824
rect 1935 820 1939 824
rect 2015 820 2019 824
rect 2071 820 2075 824
rect 279 812 283 816
rect 343 812 347 816
rect 415 812 419 816
rect 487 812 491 816
rect 567 812 571 816
rect 647 812 651 816
rect 727 812 731 816
rect 799 812 803 816
rect 863 812 867 816
rect 927 812 931 816
rect 999 812 1003 816
rect 1047 812 1051 816
rect 1183 811 1184 815
rect 1184 811 1187 815
rect 1263 811 1267 815
rect 1375 811 1379 815
rect 1483 811 1484 815
rect 1484 811 1487 815
rect 1735 811 1736 815
rect 1736 811 1739 815
rect 1819 811 1823 815
rect 1911 811 1915 815
rect 111 804 115 808
rect 1095 804 1099 808
rect 335 799 339 803
rect 443 799 444 803
rect 444 799 447 803
rect 507 799 511 803
rect 583 799 587 803
rect 663 799 667 803
rect 755 799 756 803
rect 756 799 759 803
rect 815 799 819 803
rect 1015 799 1019 803
rect 1895 803 1899 807
rect 2095 811 2096 815
rect 2096 811 2099 815
rect 111 787 115 791
rect 279 784 283 788
rect 343 784 347 788
rect 415 784 419 788
rect 487 784 491 788
rect 567 784 571 788
rect 647 784 651 788
rect 727 784 731 788
rect 799 784 803 788
rect 863 784 867 788
rect 927 784 931 788
rect 999 784 1003 788
rect 1047 784 1051 788
rect 1095 787 1099 791
rect 1423 791 1427 795
rect 1463 791 1467 795
rect 1559 791 1563 795
rect 1567 791 1571 795
rect 1919 791 1923 795
rect 1979 791 1983 795
rect 1987 791 1991 795
rect 1159 784 1163 788
rect 1279 784 1283 788
rect 1407 784 1411 788
rect 1519 784 1523 788
rect 1623 784 1627 788
rect 1719 784 1723 788
rect 1815 784 1819 788
rect 1903 784 1907 788
rect 1999 784 2003 788
rect 2071 784 2075 788
rect 111 769 115 773
rect 215 772 219 776
rect 279 772 283 776
rect 351 772 355 776
rect 423 772 427 776
rect 495 772 499 776
rect 567 772 571 776
rect 639 772 643 776
rect 703 772 707 776
rect 759 772 763 776
rect 815 772 819 776
rect 863 772 867 776
rect 911 772 915 776
rect 959 772 963 776
rect 1007 772 1011 776
rect 1047 772 1051 776
rect 1135 776 1139 780
rect 2119 776 2123 780
rect 1095 769 1099 773
rect 1183 771 1184 775
rect 1184 771 1187 775
rect 1423 771 1427 775
rect 1567 771 1571 775
rect 1823 771 1827 775
rect 1911 771 1915 775
rect 1919 771 1923 775
rect 1979 771 1983 775
rect 2095 771 2096 775
rect 2096 771 2099 775
rect 111 752 115 756
rect 203 755 207 759
rect 583 755 587 759
rect 671 763 675 767
rect 887 763 891 767
rect 663 755 664 759
rect 664 755 667 759
rect 751 755 755 759
rect 879 755 883 759
rect 927 755 931 759
rect 1023 755 1027 759
rect 1063 755 1067 759
rect 1071 755 1072 759
rect 1072 755 1075 759
rect 1135 759 1139 763
rect 1095 752 1099 756
rect 1159 756 1163 760
rect 1279 756 1283 760
rect 1407 756 1411 760
rect 1519 756 1523 760
rect 1623 756 1627 760
rect 1719 756 1723 760
rect 1815 756 1819 760
rect 1903 756 1907 760
rect 1999 756 2003 760
rect 2071 756 2075 760
rect 2119 759 2123 763
rect 215 744 219 748
rect 279 744 283 748
rect 351 744 355 748
rect 423 744 427 748
rect 495 744 499 748
rect 567 744 571 748
rect 639 744 643 748
rect 703 744 707 748
rect 759 744 763 748
rect 815 744 819 748
rect 863 744 867 748
rect 911 744 915 748
rect 959 744 963 748
rect 1007 744 1011 748
rect 1047 744 1051 748
rect 443 735 447 739
rect 559 735 563 739
rect 583 735 587 739
rect 751 735 755 739
rect 823 735 827 739
rect 879 735 883 739
rect 927 735 931 739
rect 1015 735 1019 739
rect 1023 735 1027 739
rect 1063 735 1067 739
rect 1135 737 1139 741
rect 1335 740 1339 744
rect 1375 740 1379 744
rect 1415 740 1419 744
rect 1455 740 1459 744
rect 1503 740 1507 744
rect 1551 740 1555 744
rect 1599 740 1603 744
rect 1655 740 1659 744
rect 1711 740 1715 744
rect 1767 740 1771 744
rect 1831 740 1835 744
rect 1895 740 1899 744
rect 1959 740 1963 744
rect 2023 740 2027 744
rect 2071 740 2075 744
rect 2119 737 2123 741
rect 663 727 667 731
rect 1623 731 1627 735
rect 203 715 204 719
rect 204 715 207 719
rect 211 715 215 719
rect 419 715 420 719
rect 420 715 423 719
rect 427 715 431 719
rect 695 715 699 719
rect 727 715 731 719
rect 175 708 179 712
rect 239 708 243 712
rect 311 708 315 712
rect 391 708 395 712
rect 471 708 475 712
rect 543 708 547 712
rect 615 708 619 712
rect 679 708 683 712
rect 735 708 739 712
rect 111 700 115 704
rect 1135 720 1139 724
rect 1363 723 1364 727
rect 1364 723 1367 727
rect 1383 723 1387 727
rect 1423 723 1427 727
rect 1463 723 1467 727
rect 1679 723 1680 727
rect 1680 723 1683 727
rect 1759 723 1763 727
rect 1975 723 1979 727
rect 1987 723 1988 727
rect 1988 723 1991 727
rect 2047 723 2048 727
rect 2048 723 2051 727
rect 879 715 883 719
rect 943 715 947 719
rect 2119 720 2123 724
rect 799 708 803 712
rect 863 708 867 712
rect 927 708 931 712
rect 1335 712 1339 716
rect 1375 712 1379 716
rect 1415 712 1419 716
rect 1455 712 1459 716
rect 1503 712 1507 716
rect 1551 712 1555 716
rect 1599 712 1603 716
rect 1655 712 1659 716
rect 1711 712 1715 716
rect 1767 712 1771 716
rect 1831 712 1835 716
rect 1895 712 1899 716
rect 1959 712 1963 716
rect 2023 712 2027 716
rect 2071 712 2075 716
rect 1095 700 1099 704
rect 1383 703 1387 707
rect 1423 703 1427 707
rect 1463 703 1467 707
rect 1623 703 1624 707
rect 1624 703 1627 707
rect 1759 703 1763 707
rect 1823 703 1827 707
rect 1935 703 1939 707
rect 1975 703 1979 707
rect 2095 703 2096 707
rect 2096 703 2099 707
rect 211 695 215 699
rect 299 695 303 699
rect 427 695 431 699
rect 559 695 563 699
rect 695 695 699 699
rect 823 695 824 699
rect 824 695 827 699
rect 879 695 883 699
rect 943 695 947 699
rect 1363 691 1367 695
rect 1679 691 1683 695
rect 1947 691 1951 695
rect 111 683 115 687
rect 175 680 179 684
rect 239 680 243 684
rect 311 680 315 684
rect 391 680 395 684
rect 471 680 475 684
rect 543 680 547 684
rect 615 680 619 684
rect 679 680 683 684
rect 735 680 739 684
rect 799 680 803 684
rect 863 680 867 684
rect 927 680 931 684
rect 1095 683 1099 687
rect 1303 683 1307 687
rect 1351 683 1355 687
rect 1407 683 1411 687
rect 1463 683 1467 687
rect 1527 683 1531 687
rect 1671 683 1675 687
rect 1719 683 1723 687
rect 1839 683 1843 687
rect 1247 676 1251 680
rect 1287 676 1291 680
rect 1335 676 1339 680
rect 1391 676 1395 680
rect 1447 676 1451 680
rect 1511 676 1515 680
rect 1583 676 1587 680
rect 1655 676 1659 680
rect 1735 676 1739 680
rect 1823 676 1827 680
rect 1911 676 1915 680
rect 111 665 115 669
rect 135 668 139 672
rect 175 668 179 672
rect 215 668 219 672
rect 271 668 275 672
rect 335 668 339 672
rect 399 668 403 672
rect 463 668 467 672
rect 527 668 531 672
rect 591 668 595 672
rect 647 668 651 672
rect 703 668 707 672
rect 759 668 763 672
rect 823 668 827 672
rect 1095 665 1099 669
rect 1135 668 1139 672
rect 847 659 851 663
rect 1295 663 1299 667
rect 1303 663 1307 667
rect 1351 663 1355 667
rect 1407 663 1411 667
rect 1463 663 1467 667
rect 1527 663 1531 667
rect 1663 663 1667 667
rect 1671 663 1675 667
rect 1719 663 1723 667
rect 1839 663 1843 667
rect 1935 663 1936 667
rect 1936 663 1939 667
rect 2047 683 2051 687
rect 1999 676 2003 680
rect 2071 676 2075 680
rect 2119 668 2123 672
rect 2095 663 2096 667
rect 2096 663 2099 667
rect 111 648 115 652
rect 163 651 164 655
rect 164 651 167 655
rect 183 651 187 655
rect 223 651 227 655
rect 135 640 139 644
rect 175 640 179 644
rect 215 640 219 644
rect 271 640 275 644
rect 335 640 339 644
rect 399 640 403 644
rect 419 651 423 655
rect 551 651 552 655
rect 552 651 555 655
rect 727 651 728 655
rect 728 651 731 655
rect 751 651 755 655
rect 1095 648 1099 652
rect 1135 651 1139 655
rect 1247 648 1251 652
rect 1287 648 1291 652
rect 1335 648 1339 652
rect 1391 648 1395 652
rect 1447 648 1451 652
rect 1511 648 1515 652
rect 1583 648 1587 652
rect 1655 648 1659 652
rect 1735 648 1739 652
rect 1823 648 1827 652
rect 1911 648 1915 652
rect 1999 648 2003 652
rect 2071 648 2075 652
rect 2119 651 2123 655
rect 183 631 187 635
rect 223 631 227 635
rect 299 631 300 635
rect 300 631 303 635
rect 343 631 347 635
rect 463 640 467 644
rect 527 640 531 644
rect 591 640 595 644
rect 647 640 651 644
rect 703 640 707 644
rect 759 640 763 644
rect 823 640 827 644
rect 655 631 659 635
rect 751 631 755 635
rect 847 631 848 635
rect 848 631 851 635
rect 1135 633 1139 637
rect 1159 636 1163 640
rect 1199 636 1203 640
rect 1239 636 1243 640
rect 1279 636 1283 640
rect 1343 636 1347 640
rect 1415 636 1419 640
rect 1495 636 1499 640
rect 1583 636 1587 640
rect 1671 636 1675 640
rect 1759 636 1763 640
rect 1839 636 1843 640
rect 1919 636 1923 640
rect 2007 636 2011 640
rect 2071 636 2075 640
rect 2119 633 2123 637
rect 551 623 555 627
rect 1135 616 1139 620
rect 1183 619 1184 623
rect 1184 619 1187 623
rect 1207 619 1211 623
rect 1247 619 1251 623
rect 1287 619 1291 623
rect 1519 619 1520 623
rect 1520 619 1523 623
rect 1935 619 1939 623
rect 1947 619 1948 623
rect 1948 619 1951 623
rect 2047 619 2051 623
rect 2055 619 2059 623
rect 163 611 167 615
rect 2119 616 2123 620
rect 611 611 615 615
rect 1159 608 1163 612
rect 191 603 195 607
rect 231 603 235 607
rect 271 603 275 607
rect 367 603 371 607
rect 415 603 419 607
rect 447 603 451 607
rect 479 603 483 607
rect 495 603 499 607
rect 527 603 531 607
rect 687 603 691 607
rect 743 603 747 607
rect 1199 608 1203 612
rect 1239 608 1243 612
rect 1279 608 1283 612
rect 1343 608 1347 612
rect 1415 608 1419 612
rect 1495 608 1499 612
rect 1583 608 1587 612
rect 1671 608 1675 612
rect 1759 608 1763 612
rect 1839 608 1843 612
rect 1919 608 1923 612
rect 2007 608 2011 612
rect 2071 608 2075 612
rect 135 596 139 600
rect 175 596 179 600
rect 215 596 219 600
rect 255 596 259 600
rect 303 596 307 600
rect 351 596 355 600
rect 399 596 403 600
rect 439 596 443 600
rect 487 596 491 600
rect 535 596 539 600
rect 583 596 587 600
rect 631 596 635 600
rect 679 596 683 600
rect 727 596 731 600
rect 1207 599 1211 603
rect 1247 599 1251 603
rect 1287 599 1291 603
rect 111 588 115 592
rect 1095 588 1099 592
rect 1295 591 1299 595
rect 1663 591 1667 595
rect 1879 599 1883 603
rect 1935 599 1939 603
rect 2055 599 2059 603
rect 2095 599 2096 603
rect 2096 599 2099 603
rect 159 583 160 587
rect 160 583 163 587
rect 191 583 195 587
rect 231 583 235 587
rect 271 583 275 587
rect 343 583 347 587
rect 367 583 371 587
rect 415 583 419 587
rect 495 583 499 587
rect 527 583 531 587
rect 611 583 612 587
rect 612 583 615 587
rect 655 583 656 587
rect 656 583 659 587
rect 687 583 691 587
rect 743 583 747 587
rect 1519 583 1523 587
rect 111 571 115 575
rect 135 568 139 572
rect 175 568 179 572
rect 215 568 219 572
rect 255 568 259 572
rect 303 568 307 572
rect 351 568 355 572
rect 399 568 403 572
rect 439 568 443 572
rect 487 568 491 572
rect 535 568 539 572
rect 583 568 587 572
rect 631 568 635 572
rect 679 568 683 572
rect 727 568 731 572
rect 1095 571 1099 575
rect 1183 575 1184 579
rect 1184 575 1187 579
rect 1207 575 1211 579
rect 1247 575 1251 579
rect 1287 575 1291 579
rect 1327 575 1331 579
rect 1367 575 1371 579
rect 1671 575 1675 579
rect 1767 575 1771 579
rect 1939 575 1943 579
rect 1947 575 1951 579
rect 2047 575 2051 579
rect 1159 568 1163 572
rect 1199 568 1203 572
rect 1239 568 1243 572
rect 1279 568 1283 572
rect 1319 568 1323 572
rect 1359 568 1363 572
rect 1415 568 1419 572
rect 1487 568 1491 572
rect 1567 568 1571 572
rect 1655 568 1659 572
rect 1751 568 1755 572
rect 1855 568 1859 572
rect 1967 568 1971 572
rect 2071 568 2075 572
rect 1135 560 1139 564
rect 2119 560 2123 564
rect 111 549 115 553
rect 135 552 139 556
rect 175 552 179 556
rect 223 552 227 556
rect 279 552 283 556
rect 327 552 331 556
rect 375 552 379 556
rect 423 552 427 556
rect 463 552 467 556
rect 511 552 515 556
rect 559 552 563 556
rect 607 552 611 556
rect 655 552 659 556
rect 703 552 707 556
rect 751 552 755 556
rect 1207 555 1211 559
rect 1247 555 1251 559
rect 1287 555 1291 559
rect 1327 555 1331 559
rect 1367 555 1371 559
rect 1431 555 1435 559
rect 1535 555 1539 559
rect 1671 555 1675 559
rect 1767 555 1771 559
rect 1879 555 1880 559
rect 1880 555 1883 559
rect 1939 555 1943 559
rect 1095 549 1099 553
rect 1135 543 1139 547
rect 1159 540 1163 544
rect 111 532 115 536
rect 191 535 195 539
rect 239 535 243 539
rect 295 535 299 539
rect 319 535 323 539
rect 391 535 395 539
rect 439 535 443 539
rect 447 535 448 539
rect 448 535 451 539
rect 479 535 483 539
rect 499 535 503 539
rect 691 535 695 539
rect 1199 540 1203 544
rect 1239 540 1243 544
rect 1279 540 1283 544
rect 1319 540 1323 544
rect 1359 540 1363 544
rect 1415 540 1419 544
rect 1487 540 1491 544
rect 1567 540 1571 544
rect 1655 540 1659 544
rect 1751 540 1755 544
rect 1855 540 1859 544
rect 1967 540 1971 544
rect 2071 540 2075 544
rect 2119 543 2123 547
rect 1095 532 1099 536
rect 135 524 139 528
rect 175 524 179 528
rect 223 524 227 528
rect 279 524 283 528
rect 327 524 331 528
rect 375 524 379 528
rect 423 524 427 528
rect 463 524 467 528
rect 511 524 515 528
rect 559 524 563 528
rect 607 524 611 528
rect 655 524 659 528
rect 703 524 707 528
rect 751 524 755 528
rect 1135 521 1139 525
rect 1303 524 1307 528
rect 1343 524 1347 528
rect 1383 524 1387 528
rect 1423 524 1427 528
rect 1463 524 1467 528
rect 1503 524 1507 528
rect 1543 524 1547 528
rect 1591 524 1595 528
rect 1647 524 1651 528
rect 1703 524 1707 528
rect 1767 524 1771 528
rect 1839 524 1843 528
rect 1919 524 1923 528
rect 2007 524 2011 528
rect 2071 524 2075 528
rect 2119 521 2123 525
rect 159 515 160 519
rect 160 515 163 519
rect 191 515 195 519
rect 239 515 243 519
rect 295 515 299 519
rect 383 515 387 519
rect 391 515 395 519
rect 439 515 443 519
rect 499 515 503 519
rect 691 515 695 519
rect 583 507 587 511
rect 1135 504 1139 508
rect 1447 515 1451 519
rect 1351 507 1355 511
rect 1391 507 1395 511
rect 1479 507 1483 511
rect 1519 507 1523 511
rect 1303 496 1307 500
rect 1343 496 1347 500
rect 1383 496 1387 500
rect 1423 496 1427 500
rect 1463 496 1467 500
rect 1503 496 1507 500
rect 191 487 195 491
rect 247 487 251 491
rect 287 487 291 491
rect 319 487 320 491
rect 320 487 323 491
rect 439 487 443 491
rect 495 487 499 491
rect 551 487 555 491
rect 599 487 603 491
rect 655 487 659 491
rect 703 487 707 491
rect 751 487 755 491
rect 807 487 811 491
rect 855 487 859 491
rect 863 487 867 491
rect 1351 487 1355 491
rect 1391 487 1395 491
rect 1431 487 1435 491
rect 1447 487 1448 491
rect 1448 487 1451 491
rect 1479 487 1483 491
rect 1519 487 1523 491
rect 1555 507 1559 511
rect 1663 507 1667 511
rect 1719 507 1723 511
rect 1783 507 1787 511
rect 1847 507 1851 511
rect 1911 507 1915 511
rect 1947 507 1948 511
rect 1948 507 1951 511
rect 2079 507 2083 511
rect 2095 507 2096 511
rect 2096 507 2099 511
rect 2119 504 2123 508
rect 1543 496 1547 500
rect 1591 496 1595 500
rect 1647 496 1651 500
rect 1703 496 1707 500
rect 1767 496 1771 500
rect 1839 496 1843 500
rect 1919 496 1923 500
rect 2007 496 2011 500
rect 2071 496 2075 500
rect 135 480 139 484
rect 175 480 179 484
rect 231 480 235 484
rect 295 480 299 484
rect 359 480 363 484
rect 423 480 427 484
rect 479 480 483 484
rect 535 480 539 484
rect 591 480 595 484
rect 639 480 643 484
rect 687 480 691 484
rect 735 480 739 484
rect 791 480 795 484
rect 847 480 851 484
rect 1535 479 1539 483
rect 1663 487 1667 491
rect 1719 487 1723 491
rect 1783 487 1787 491
rect 1847 487 1851 491
rect 1999 487 2003 491
rect 2079 487 2083 491
rect 111 472 115 476
rect 183 467 187 471
rect 191 467 195 471
rect 247 467 251 471
rect 287 467 291 471
rect 383 467 384 471
rect 384 467 387 471
rect 439 467 443 471
rect 495 467 499 471
rect 583 471 587 475
rect 1095 472 1099 476
rect 599 467 603 471
rect 655 467 659 471
rect 703 467 707 471
rect 751 467 755 471
rect 807 467 811 471
rect 855 467 859 471
rect 1351 467 1355 471
rect 1391 467 1395 471
rect 1439 467 1443 471
rect 1487 467 1491 471
rect 1543 467 1547 471
rect 1555 467 1556 471
rect 1556 467 1559 471
rect 1663 467 1667 471
rect 1735 467 1739 471
rect 1823 467 1827 471
rect 1903 467 1907 471
rect 1911 467 1915 471
rect 2019 467 2020 471
rect 2020 467 2023 471
rect 2095 467 2096 471
rect 2096 467 2099 471
rect 1295 460 1299 464
rect 111 455 115 459
rect 1335 460 1339 464
rect 1375 460 1379 464
rect 1423 460 1427 464
rect 1471 460 1475 464
rect 1527 460 1531 464
rect 1583 460 1587 464
rect 1647 460 1651 464
rect 1719 460 1723 464
rect 1807 460 1811 464
rect 1895 460 1899 464
rect 1991 460 1995 464
rect 2071 460 2075 464
rect 135 452 139 456
rect 175 452 179 456
rect 231 452 235 456
rect 295 452 299 456
rect 359 452 363 456
rect 423 452 427 456
rect 479 452 483 456
rect 535 452 539 456
rect 591 452 595 456
rect 639 452 643 456
rect 687 452 691 456
rect 735 452 739 456
rect 791 452 795 456
rect 847 452 851 456
rect 1095 455 1099 459
rect 1135 452 1139 456
rect 2119 452 2123 456
rect 1343 447 1347 451
rect 1351 447 1355 451
rect 1391 447 1395 451
rect 1439 447 1443 451
rect 1487 447 1491 451
rect 1543 447 1547 451
rect 1611 447 1612 451
rect 1612 447 1615 451
rect 1663 447 1667 451
rect 1735 447 1739 451
rect 1823 447 1827 451
rect 1903 447 1907 451
rect 1999 447 2003 451
rect 2095 447 2096 451
rect 2096 447 2099 451
rect 111 433 115 437
rect 175 436 179 440
rect 215 436 219 440
rect 263 436 267 440
rect 327 436 331 440
rect 391 436 395 440
rect 463 436 467 440
rect 535 436 539 440
rect 607 436 611 440
rect 679 436 683 440
rect 743 436 747 440
rect 807 436 811 440
rect 871 436 875 440
rect 943 436 947 440
rect 1095 433 1099 437
rect 1135 435 1139 439
rect 1295 432 1299 436
rect 1335 432 1339 436
rect 1375 432 1379 436
rect 1423 432 1427 436
rect 1471 432 1475 436
rect 1527 432 1531 436
rect 1583 432 1587 436
rect 1647 432 1651 436
rect 1719 432 1723 436
rect 1807 432 1811 436
rect 1895 432 1899 436
rect 1991 432 1995 436
rect 2071 432 2075 436
rect 2119 435 2123 439
rect 863 427 867 431
rect 111 416 115 420
rect 199 419 200 423
rect 200 419 203 423
rect 223 419 227 423
rect 251 419 255 423
rect 351 419 352 423
rect 352 419 355 423
rect 551 419 555 423
rect 559 419 560 423
rect 560 419 563 423
rect 1095 416 1099 420
rect 1135 417 1139 421
rect 1159 420 1163 424
rect 1199 420 1203 424
rect 1255 420 1259 424
rect 1335 420 1339 424
rect 1415 420 1419 424
rect 1503 420 1507 424
rect 1591 420 1595 424
rect 1671 420 1675 424
rect 1751 420 1755 424
rect 1831 420 1835 424
rect 1911 420 1915 424
rect 1999 420 2003 424
rect 2071 420 2075 424
rect 2119 417 2123 421
rect 175 408 179 412
rect 215 408 219 412
rect 263 408 267 412
rect 327 408 331 412
rect 391 408 395 412
rect 463 408 467 412
rect 535 408 539 412
rect 607 408 611 412
rect 679 408 683 412
rect 743 408 747 412
rect 807 408 811 412
rect 871 408 875 412
rect 943 408 947 412
rect 1487 411 1491 415
rect 223 399 227 403
rect 251 399 255 403
rect 183 391 187 395
rect 431 399 435 403
rect 551 399 555 403
rect 915 399 919 403
rect 1135 400 1139 404
rect 1207 403 1211 407
rect 1855 411 1859 415
rect 1687 403 1691 407
rect 1707 403 1711 407
rect 2011 403 2015 407
rect 2019 403 2023 407
rect 2119 400 2123 404
rect 351 391 355 395
rect 1159 392 1163 396
rect 1199 392 1203 396
rect 1255 392 1259 396
rect 1335 392 1339 396
rect 1415 392 1419 396
rect 1503 392 1507 396
rect 1591 392 1595 396
rect 1671 392 1675 396
rect 1751 392 1755 396
rect 1831 392 1835 396
rect 1911 392 1915 396
rect 1999 392 2003 396
rect 2071 392 2075 396
rect 363 379 367 383
rect 1207 383 1211 387
rect 199 371 200 375
rect 200 371 203 375
rect 223 371 227 375
rect 503 371 507 375
rect 583 371 587 375
rect 727 371 731 375
rect 791 371 795 375
rect 855 371 859 375
rect 887 371 891 375
rect 967 371 971 375
rect 1023 371 1027 375
rect 1031 371 1032 375
rect 1032 371 1035 375
rect 1183 371 1187 375
rect 1343 375 1347 379
rect 1611 383 1615 387
rect 1707 383 1711 387
rect 1855 383 1856 387
rect 1856 383 1859 387
rect 1939 383 1940 387
rect 1940 383 1943 387
rect 2011 383 2015 387
rect 2095 383 2096 387
rect 2096 383 2099 387
rect 175 364 179 368
rect 215 364 219 368
rect 271 364 275 368
rect 335 364 339 368
rect 407 364 411 368
rect 487 364 491 368
rect 567 364 571 368
rect 639 364 643 368
rect 711 364 715 368
rect 775 364 779 368
rect 839 364 843 368
rect 895 364 899 368
rect 951 364 955 368
rect 1007 364 1011 368
rect 1047 364 1051 368
rect 111 356 115 360
rect 1095 356 1099 360
rect 1263 359 1267 363
rect 1327 359 1331 363
rect 1479 359 1483 363
rect 1487 359 1488 363
rect 1488 359 1491 363
rect 1663 359 1667 363
rect 1687 363 1691 367
rect 223 351 227 355
rect 363 351 364 355
rect 364 351 367 355
rect 431 351 432 355
rect 432 351 435 355
rect 503 351 507 355
rect 583 351 587 355
rect 667 351 668 355
rect 668 351 671 355
rect 727 351 731 355
rect 791 351 795 355
rect 855 351 859 355
rect 887 351 891 355
rect 967 351 971 355
rect 1023 351 1027 355
rect 1071 351 1072 355
rect 1072 351 1075 355
rect 1159 352 1163 356
rect 1247 352 1251 356
rect 1359 352 1363 356
rect 1463 352 1467 356
rect 1559 352 1563 356
rect 1647 352 1651 356
rect 1991 359 1995 363
rect 2047 359 2051 363
rect 2087 359 2091 363
rect 1727 352 1731 356
rect 1135 344 1139 348
rect 111 339 115 343
rect 175 336 179 340
rect 215 336 219 340
rect 271 336 275 340
rect 335 336 339 340
rect 407 336 411 340
rect 487 336 491 340
rect 567 336 571 340
rect 639 336 643 340
rect 711 336 715 340
rect 775 336 779 340
rect 839 336 843 340
rect 895 336 899 340
rect 951 336 955 340
rect 1007 336 1011 340
rect 1047 336 1051 340
rect 1095 339 1099 343
rect 1183 339 1184 343
rect 1184 339 1187 343
rect 1263 339 1267 343
rect 1327 339 1331 343
rect 1479 339 1483 343
rect 1799 352 1803 356
rect 1863 352 1867 356
rect 1919 352 1923 356
rect 1975 352 1979 356
rect 2031 352 2035 356
rect 2071 352 2075 356
rect 2119 344 2123 348
rect 1663 339 1667 343
rect 1911 339 1915 343
rect 1939 339 1943 343
rect 1991 339 1995 343
rect 2047 339 2051 343
rect 2087 339 2091 343
rect 1135 327 1139 331
rect 111 317 115 321
rect 383 320 387 324
rect 423 320 427 324
rect 463 320 467 324
rect 503 320 507 324
rect 543 320 547 324
rect 591 320 595 324
rect 639 320 643 324
rect 687 320 691 324
rect 735 320 739 324
rect 783 320 787 324
rect 831 320 835 324
rect 879 320 883 324
rect 927 320 931 324
rect 967 320 971 324
rect 1007 320 1011 324
rect 1047 320 1051 324
rect 1159 324 1163 328
rect 1247 324 1251 328
rect 1359 324 1363 328
rect 1463 324 1467 328
rect 1559 324 1563 328
rect 1647 324 1651 328
rect 1727 324 1731 328
rect 1799 324 1803 328
rect 1863 324 1867 328
rect 1919 324 1923 328
rect 1975 324 1979 328
rect 2031 324 2035 328
rect 2071 324 2075 328
rect 2119 327 2123 331
rect 1095 317 1099 321
rect 1031 311 1035 315
rect 111 300 115 304
rect 407 303 408 307
rect 408 303 411 307
rect 431 303 435 307
rect 471 303 475 307
rect 511 303 515 307
rect 551 303 555 307
rect 763 303 764 307
rect 764 303 767 307
rect 771 303 775 307
rect 975 303 979 307
rect 1015 303 1019 307
rect 1055 303 1059 307
rect 1095 300 1099 304
rect 1135 301 1139 305
rect 1351 304 1355 308
rect 1391 304 1395 308
rect 1431 304 1435 308
rect 1471 304 1475 308
rect 1511 304 1515 308
rect 1559 304 1563 308
rect 1615 304 1619 308
rect 1671 304 1675 308
rect 1735 304 1739 308
rect 1807 304 1811 308
rect 1887 304 1891 308
rect 1967 304 1971 308
rect 2047 304 2051 308
rect 2119 301 2123 305
rect 383 292 387 296
rect 423 292 427 296
rect 463 292 467 296
rect 503 292 507 296
rect 543 292 547 296
rect 591 292 595 296
rect 639 292 643 296
rect 687 292 691 296
rect 735 292 739 296
rect 783 292 787 296
rect 831 292 835 296
rect 879 292 883 296
rect 927 292 931 296
rect 967 292 971 296
rect 1007 292 1011 296
rect 1047 292 1051 296
rect 431 283 435 287
rect 471 283 475 287
rect 511 283 515 287
rect 551 283 555 287
rect 707 283 711 287
rect 771 283 775 287
rect 887 283 891 287
rect 975 283 979 287
rect 1015 283 1019 287
rect 1055 283 1059 287
rect 1071 283 1072 287
rect 1072 283 1075 287
rect 1135 284 1139 288
rect 1375 287 1376 291
rect 1376 287 1379 291
rect 1399 287 1403 291
rect 1439 287 1443 291
rect 1479 287 1483 291
rect 1519 287 1523 291
rect 1723 287 1727 291
rect 1983 287 1987 291
rect 2063 287 2067 291
rect 2095 287 2099 291
rect 2119 284 2123 288
rect 1351 276 1355 280
rect 1391 276 1395 280
rect 1431 276 1435 280
rect 1471 276 1475 280
rect 1511 276 1515 280
rect 1559 276 1563 280
rect 1615 276 1619 280
rect 1671 276 1675 280
rect 1735 276 1739 280
rect 1807 276 1811 280
rect 1887 276 1891 280
rect 1967 276 1971 280
rect 2047 276 2051 280
rect 407 263 411 267
rect 1399 267 1403 271
rect 1439 267 1443 271
rect 1479 267 1483 271
rect 1519 267 1523 271
rect 1723 267 1727 271
rect 343 255 347 259
rect 375 255 379 259
rect 431 255 435 259
rect 487 255 491 259
rect 551 255 555 259
rect 623 255 627 259
rect 699 255 703 259
rect 763 255 767 259
rect 287 248 291 252
rect 327 248 331 252
rect 367 248 371 252
rect 415 248 419 252
rect 471 248 475 252
rect 535 248 539 252
rect 607 248 611 252
rect 679 248 683 252
rect 743 248 747 252
rect 943 255 947 259
rect 1007 255 1011 259
rect 1063 255 1067 259
rect 1071 255 1072 259
rect 1072 255 1075 259
rect 1375 255 1379 259
rect 1571 259 1575 263
rect 1911 267 1912 271
rect 1912 267 1915 271
rect 1983 267 1987 271
rect 2063 267 2067 271
rect 807 248 811 252
rect 863 248 867 252
rect 927 248 931 252
rect 991 248 995 252
rect 1047 248 1051 252
rect 1319 247 1323 251
rect 1359 247 1363 251
rect 1399 247 1403 251
rect 1439 247 1443 251
rect 1479 247 1483 251
rect 1519 247 1523 251
rect 1615 247 1619 251
rect 1687 247 1691 251
rect 1775 247 1779 251
rect 1879 247 1883 251
rect 1999 247 2000 251
rect 2000 247 2003 251
rect 2095 247 2096 251
rect 2096 247 2099 251
rect 111 240 115 244
rect 1095 240 1099 244
rect 335 235 339 239
rect 343 235 347 239
rect 375 235 379 239
rect 431 235 435 239
rect 487 235 491 239
rect 551 235 555 239
rect 623 235 627 239
rect 707 235 708 239
rect 708 235 711 239
rect 779 235 783 239
rect 887 235 888 239
rect 888 235 891 239
rect 943 235 947 239
rect 1007 235 1011 239
rect 1063 235 1067 239
rect 1263 240 1267 244
rect 1303 240 1307 244
rect 1343 240 1347 244
rect 1383 240 1387 244
rect 1423 240 1427 244
rect 1463 240 1467 244
rect 1503 240 1507 244
rect 1543 240 1547 244
rect 1599 240 1603 244
rect 1671 240 1675 244
rect 1759 240 1763 244
rect 1863 240 1867 244
rect 1975 240 1979 244
rect 2071 240 2075 244
rect 1135 232 1139 236
rect 2119 232 2123 236
rect 111 223 115 227
rect 287 220 291 224
rect 327 220 331 224
rect 367 220 371 224
rect 415 220 419 224
rect 471 220 475 224
rect 535 220 539 224
rect 607 220 611 224
rect 679 220 683 224
rect 743 220 747 224
rect 807 220 811 224
rect 863 220 867 224
rect 927 220 931 224
rect 991 220 995 224
rect 1047 220 1051 224
rect 1095 223 1099 227
rect 1311 227 1315 231
rect 1319 227 1323 231
rect 1359 227 1363 231
rect 1399 227 1403 231
rect 1439 227 1443 231
rect 1479 227 1483 231
rect 1519 227 1523 231
rect 1571 227 1572 231
rect 1572 227 1575 231
rect 1615 227 1619 231
rect 1687 227 1691 231
rect 1775 227 1779 231
rect 1879 227 1883 231
rect 2063 227 2067 231
rect 1135 215 1139 219
rect 1263 212 1267 216
rect 1303 212 1307 216
rect 1343 212 1347 216
rect 1383 212 1387 216
rect 1423 212 1427 216
rect 1463 212 1467 216
rect 1503 212 1507 216
rect 1543 212 1547 216
rect 1599 212 1603 216
rect 1671 212 1675 216
rect 1759 212 1763 216
rect 1863 212 1867 216
rect 1975 212 1979 216
rect 2071 212 2075 216
rect 2119 215 2123 219
rect 1615 203 1619 207
rect 1999 203 2003 207
rect 111 193 115 197
rect 167 196 171 200
rect 207 196 211 200
rect 247 196 251 200
rect 295 196 299 200
rect 343 196 347 200
rect 399 196 403 200
rect 463 196 467 200
rect 527 196 531 200
rect 599 196 603 200
rect 671 196 675 200
rect 751 196 755 200
rect 831 196 835 200
rect 911 196 915 200
rect 991 196 995 200
rect 1047 196 1051 200
rect 1095 193 1099 197
rect 1135 193 1139 197
rect 1183 196 1187 200
rect 1231 196 1235 200
rect 1295 196 1299 200
rect 1359 196 1363 200
rect 1431 196 1435 200
rect 1511 196 1515 200
rect 1591 196 1595 200
rect 1663 196 1667 200
rect 1735 196 1739 200
rect 1807 196 1811 200
rect 1879 196 1883 200
rect 1951 196 1955 200
rect 2023 196 2027 200
rect 2071 196 2075 200
rect 2119 193 2123 197
rect 1975 187 1979 191
rect 111 176 115 180
rect 195 179 196 183
rect 196 179 199 183
rect 215 179 219 183
rect 255 179 259 183
rect 615 179 619 183
rect 679 179 683 183
rect 699 179 700 183
rect 700 179 703 183
rect 847 179 851 183
rect 927 179 931 183
rect 959 179 963 183
rect 1063 179 1067 183
rect 1071 179 1072 183
rect 1072 179 1075 183
rect 1095 176 1099 180
rect 1135 176 1139 180
rect 1211 179 1212 183
rect 1212 179 1215 183
rect 1219 179 1223 183
rect 1615 179 1616 183
rect 1616 179 1619 183
rect 2087 179 2091 183
rect 2095 179 2096 183
rect 2096 179 2099 183
rect 2119 176 2123 180
rect 167 168 171 172
rect 207 168 211 172
rect 247 168 251 172
rect 295 168 299 172
rect 343 168 347 172
rect 399 168 403 172
rect 463 168 467 172
rect 527 168 531 172
rect 599 168 603 172
rect 671 168 675 172
rect 751 168 755 172
rect 831 168 835 172
rect 911 168 915 172
rect 991 168 995 172
rect 1047 168 1051 172
rect 1183 168 1187 172
rect 1231 168 1235 172
rect 1295 168 1299 172
rect 1359 168 1363 172
rect 1431 168 1435 172
rect 1511 168 1515 172
rect 1591 168 1595 172
rect 1663 168 1667 172
rect 1735 168 1739 172
rect 1807 168 1811 172
rect 1879 168 1883 172
rect 1951 168 1955 172
rect 2023 168 2027 172
rect 2071 168 2075 172
rect 215 159 219 163
rect 255 159 259 163
rect 335 151 339 155
rect 555 159 556 163
rect 556 159 559 163
rect 615 159 619 163
rect 679 159 683 163
rect 779 159 780 163
rect 780 159 783 163
rect 847 159 851 163
rect 927 159 931 163
rect 1019 159 1020 163
rect 1020 159 1023 163
rect 1063 159 1067 163
rect 1219 159 1223 163
rect 1311 151 1315 155
rect 1599 151 1603 155
rect 2015 159 2019 163
rect 2063 159 2067 163
rect 2087 159 2091 163
rect 195 131 199 135
rect 191 123 195 127
rect 231 123 235 127
rect 271 123 275 127
rect 303 123 307 127
rect 351 123 355 127
rect 391 123 395 127
rect 431 123 435 127
rect 471 123 475 127
rect 511 123 515 127
rect 591 123 595 127
rect 631 123 635 127
rect 671 123 675 127
rect 711 123 715 127
rect 751 123 755 127
rect 791 123 795 127
rect 831 123 835 127
rect 887 123 891 127
rect 943 123 947 127
rect 959 123 960 127
rect 960 123 963 127
rect 1063 123 1067 127
rect 1175 123 1179 127
rect 1211 123 1215 127
rect 135 116 139 120
rect 175 116 179 120
rect 215 116 219 120
rect 255 116 259 120
rect 295 116 299 120
rect 335 116 339 120
rect 375 116 379 120
rect 415 116 419 120
rect 455 116 459 120
rect 495 116 499 120
rect 535 116 539 120
rect 575 116 579 120
rect 615 116 619 120
rect 655 116 659 120
rect 695 116 699 120
rect 735 116 739 120
rect 775 116 779 120
rect 815 116 819 120
rect 871 116 875 120
rect 935 116 939 120
rect 999 116 1003 120
rect 1047 116 1051 120
rect 1215 115 1219 119
rect 1255 115 1259 119
rect 1295 115 1299 119
rect 1335 115 1339 119
rect 1383 115 1387 119
rect 1447 115 1451 119
rect 1503 115 1507 119
rect 1631 115 1635 119
rect 1687 115 1691 119
rect 1735 115 1739 119
rect 1783 115 1787 119
rect 1823 115 1827 119
rect 1871 115 1875 119
rect 1919 115 1923 119
rect 1967 115 1971 119
rect 1975 115 1976 119
rect 1976 115 1979 119
rect 2047 115 2051 119
rect 2087 115 2091 119
rect 2095 115 2096 119
rect 2096 115 2099 119
rect 111 108 115 112
rect 1095 108 1099 112
rect 191 103 195 107
rect 231 103 235 107
rect 271 103 275 107
rect 303 103 307 107
rect 351 103 355 107
rect 391 103 395 107
rect 431 103 435 107
rect 471 103 475 107
rect 511 103 515 107
rect 555 103 559 107
rect 591 103 595 107
rect 631 103 635 107
rect 671 103 675 107
rect 711 103 715 107
rect 751 103 755 107
rect 791 103 795 107
rect 831 103 835 107
rect 887 103 891 107
rect 943 103 947 107
rect 1019 103 1023 107
rect 1063 103 1067 107
rect 1159 108 1163 112
rect 1199 108 1203 112
rect 1239 108 1243 112
rect 1279 108 1283 112
rect 1319 108 1323 112
rect 1367 108 1371 112
rect 1431 108 1435 112
rect 1495 108 1499 112
rect 1559 108 1563 112
rect 1615 108 1619 112
rect 1671 108 1675 112
rect 1719 108 1723 112
rect 1767 108 1771 112
rect 1807 108 1811 112
rect 1855 108 1859 112
rect 1903 108 1907 112
rect 1951 108 1955 112
rect 1991 108 1995 112
rect 2031 108 2035 112
rect 2071 108 2075 112
rect 1135 100 1139 104
rect 2119 100 2123 104
rect 111 91 115 95
rect 135 88 139 92
rect 175 88 179 92
rect 215 88 219 92
rect 255 88 259 92
rect 295 88 299 92
rect 335 88 339 92
rect 375 88 379 92
rect 415 88 419 92
rect 455 88 459 92
rect 495 88 499 92
rect 535 88 539 92
rect 575 88 579 92
rect 615 88 619 92
rect 655 88 659 92
rect 695 88 699 92
rect 735 88 739 92
rect 775 88 779 92
rect 815 88 819 92
rect 871 88 875 92
rect 935 88 939 92
rect 999 88 1003 92
rect 1047 88 1051 92
rect 1095 91 1099 95
rect 1175 95 1179 99
rect 1215 95 1219 99
rect 1255 95 1259 99
rect 1295 95 1299 99
rect 1335 95 1339 99
rect 1383 95 1387 99
rect 1447 95 1451 99
rect 1503 95 1507 99
rect 1599 95 1603 99
rect 1631 95 1635 99
rect 1687 95 1691 99
rect 1735 95 1739 99
rect 1783 95 1787 99
rect 1823 95 1827 99
rect 1871 95 1875 99
rect 1919 95 1923 99
rect 1967 95 1971 99
rect 2015 95 2016 99
rect 2016 95 2019 99
rect 2047 95 2051 99
rect 2087 95 2091 99
rect 1135 83 1139 87
rect 1159 80 1163 84
rect 1199 80 1203 84
rect 1239 80 1243 84
rect 1279 80 1283 84
rect 1319 80 1323 84
rect 1367 80 1371 84
rect 1431 80 1435 84
rect 1495 80 1499 84
rect 1559 80 1563 84
rect 1615 80 1619 84
rect 1671 80 1675 84
rect 1719 80 1723 84
rect 1767 80 1771 84
rect 1807 80 1811 84
rect 1855 80 1859 84
rect 1903 80 1907 84
rect 1951 80 1955 84
rect 1991 80 1995 84
rect 2031 80 2035 84
rect 2071 80 2075 84
rect 2119 83 2123 87
<< m3 >>
rect 1135 2214 1139 2215
rect 1135 2209 1139 2210
rect 1343 2214 1347 2215
rect 1343 2209 1347 2210
rect 1383 2214 1387 2215
rect 1383 2209 1387 2210
rect 1423 2214 1427 2215
rect 1423 2209 1427 2210
rect 1463 2214 1467 2215
rect 1463 2209 1467 2210
rect 1503 2214 1507 2215
rect 1503 2209 1507 2210
rect 1543 2214 1547 2215
rect 1543 2209 1547 2210
rect 1583 2214 1587 2215
rect 1583 2209 1587 2210
rect 1623 2214 1627 2215
rect 1663 2214 1667 2215
rect 1623 2209 1627 2210
rect 1646 2211 1652 2212
rect 1136 2189 1138 2209
rect 1344 2197 1346 2209
rect 1384 2197 1386 2209
rect 1398 2203 1404 2204
rect 1398 2199 1399 2203
rect 1403 2199 1404 2203
rect 1398 2198 1404 2199
rect 1342 2196 1348 2197
rect 1342 2192 1343 2196
rect 1347 2192 1348 2196
rect 1342 2191 1348 2192
rect 1382 2196 1388 2197
rect 1382 2192 1383 2196
rect 1387 2192 1388 2196
rect 1382 2191 1388 2192
rect 1134 2188 1140 2189
rect 1134 2184 1135 2188
rect 1139 2184 1140 2188
rect 1400 2184 1402 2198
rect 1424 2197 1426 2209
rect 1438 2203 1444 2204
rect 1438 2199 1439 2203
rect 1443 2199 1444 2203
rect 1438 2198 1444 2199
rect 1422 2196 1428 2197
rect 1422 2192 1423 2196
rect 1427 2192 1428 2196
rect 1422 2191 1428 2192
rect 1440 2184 1442 2198
rect 1464 2197 1466 2209
rect 1478 2203 1484 2204
rect 1478 2199 1479 2203
rect 1483 2199 1484 2203
rect 1478 2198 1484 2199
rect 1462 2196 1468 2197
rect 1462 2192 1463 2196
rect 1467 2192 1468 2196
rect 1462 2191 1468 2192
rect 1480 2184 1482 2198
rect 1504 2197 1506 2209
rect 1518 2203 1524 2204
rect 1518 2199 1519 2203
rect 1523 2199 1524 2203
rect 1518 2198 1524 2199
rect 1502 2196 1508 2197
rect 1502 2192 1503 2196
rect 1507 2192 1508 2196
rect 1502 2191 1508 2192
rect 1520 2184 1522 2198
rect 1544 2197 1546 2209
rect 1558 2203 1564 2204
rect 1558 2199 1559 2203
rect 1563 2199 1564 2203
rect 1558 2198 1564 2199
rect 1542 2196 1548 2197
rect 1542 2192 1543 2196
rect 1547 2192 1548 2196
rect 1542 2191 1548 2192
rect 1560 2184 1562 2198
rect 1584 2197 1586 2209
rect 1598 2203 1604 2204
rect 1598 2199 1599 2203
rect 1603 2199 1604 2203
rect 1598 2198 1604 2199
rect 1582 2196 1588 2197
rect 1582 2192 1583 2196
rect 1587 2192 1588 2196
rect 1582 2191 1588 2192
rect 1600 2184 1602 2198
rect 1624 2197 1626 2209
rect 1646 2207 1647 2211
rect 1651 2207 1652 2211
rect 1663 2209 1667 2210
rect 1703 2214 1707 2215
rect 1703 2209 1707 2210
rect 1743 2214 1747 2215
rect 1743 2209 1747 2210
rect 1783 2214 1787 2215
rect 1783 2209 1787 2210
rect 1823 2214 1827 2215
rect 1823 2209 1827 2210
rect 2119 2214 2123 2215
rect 2119 2209 2123 2210
rect 1646 2206 1652 2207
rect 1638 2203 1644 2204
rect 1638 2199 1639 2203
rect 1643 2199 1644 2203
rect 1638 2198 1644 2199
rect 1622 2196 1628 2197
rect 1622 2192 1623 2196
rect 1627 2192 1628 2196
rect 1622 2191 1628 2192
rect 1640 2184 1642 2198
rect 1134 2183 1140 2184
rect 1390 2183 1396 2184
rect 1390 2179 1391 2183
rect 1395 2179 1396 2183
rect 1390 2178 1396 2179
rect 1398 2183 1404 2184
rect 1398 2179 1399 2183
rect 1403 2179 1404 2183
rect 1398 2178 1404 2179
rect 1438 2183 1444 2184
rect 1438 2179 1439 2183
rect 1443 2179 1444 2183
rect 1438 2178 1444 2179
rect 1478 2183 1484 2184
rect 1478 2179 1479 2183
rect 1483 2179 1484 2183
rect 1478 2178 1484 2179
rect 1518 2183 1524 2184
rect 1518 2179 1519 2183
rect 1523 2179 1524 2183
rect 1518 2178 1524 2179
rect 1558 2183 1564 2184
rect 1558 2179 1559 2183
rect 1563 2179 1564 2183
rect 1558 2178 1564 2179
rect 1598 2183 1604 2184
rect 1598 2179 1599 2183
rect 1603 2179 1604 2183
rect 1598 2178 1604 2179
rect 1638 2183 1644 2184
rect 1638 2179 1639 2183
rect 1643 2179 1644 2183
rect 1638 2178 1644 2179
rect 1134 2171 1140 2172
rect 1134 2167 1135 2171
rect 1139 2167 1140 2171
rect 1134 2166 1140 2167
rect 1342 2168 1348 2169
rect 1136 2163 1138 2166
rect 1342 2164 1343 2168
rect 1347 2164 1348 2168
rect 1342 2163 1348 2164
rect 1382 2168 1388 2169
rect 1382 2164 1383 2168
rect 1387 2164 1388 2168
rect 1382 2163 1388 2164
rect 1135 2162 1139 2163
rect 1135 2157 1139 2158
rect 1287 2162 1291 2163
rect 1287 2157 1291 2158
rect 1327 2162 1331 2163
rect 1327 2157 1331 2158
rect 1343 2162 1347 2163
rect 1343 2157 1347 2158
rect 1367 2162 1371 2163
rect 1367 2157 1371 2158
rect 1383 2162 1387 2163
rect 1383 2157 1387 2158
rect 1136 2154 1138 2157
rect 1286 2156 1292 2157
rect 1134 2153 1140 2154
rect 1134 2149 1135 2153
rect 1139 2149 1140 2153
rect 1286 2152 1287 2156
rect 1291 2152 1292 2156
rect 1286 2151 1292 2152
rect 1326 2156 1332 2157
rect 1326 2152 1327 2156
rect 1331 2152 1332 2156
rect 1326 2151 1332 2152
rect 1366 2156 1372 2157
rect 1366 2152 1367 2156
rect 1371 2152 1372 2156
rect 1366 2151 1372 2152
rect 1134 2148 1140 2149
rect 1314 2139 1320 2140
rect 1134 2136 1140 2137
rect 1134 2132 1135 2136
rect 1139 2132 1140 2136
rect 1314 2135 1315 2139
rect 1319 2135 1320 2139
rect 1314 2134 1320 2135
rect 1334 2139 1340 2140
rect 1334 2135 1335 2139
rect 1339 2135 1340 2139
rect 1334 2134 1340 2135
rect 1374 2139 1380 2140
rect 1374 2135 1375 2139
rect 1379 2135 1380 2139
rect 1374 2134 1380 2135
rect 1134 2131 1140 2132
rect 1136 2107 1138 2131
rect 1286 2128 1292 2129
rect 1286 2124 1287 2128
rect 1291 2124 1292 2128
rect 1286 2123 1292 2124
rect 1288 2107 1290 2123
rect 1316 2117 1318 2134
rect 1326 2128 1332 2129
rect 1326 2124 1327 2128
rect 1331 2124 1332 2128
rect 1326 2123 1332 2124
rect 1315 2116 1319 2117
rect 1315 2111 1319 2112
rect 1328 2107 1330 2123
rect 1336 2120 1338 2134
rect 1366 2128 1372 2129
rect 1366 2124 1367 2128
rect 1371 2124 1372 2128
rect 1366 2123 1372 2124
rect 1334 2119 1340 2120
rect 1334 2115 1335 2119
rect 1339 2115 1340 2119
rect 1334 2114 1340 2115
rect 1368 2107 1370 2123
rect 1376 2120 1378 2134
rect 1374 2119 1380 2120
rect 1374 2115 1375 2119
rect 1379 2115 1380 2119
rect 1374 2114 1380 2115
rect 1392 2112 1394 2178
rect 1422 2168 1428 2169
rect 1422 2164 1423 2168
rect 1427 2164 1428 2168
rect 1422 2163 1428 2164
rect 1462 2168 1468 2169
rect 1462 2164 1463 2168
rect 1467 2164 1468 2168
rect 1462 2163 1468 2164
rect 1502 2168 1508 2169
rect 1502 2164 1503 2168
rect 1507 2164 1508 2168
rect 1502 2163 1508 2164
rect 1542 2168 1548 2169
rect 1542 2164 1543 2168
rect 1547 2164 1548 2168
rect 1542 2163 1548 2164
rect 1582 2168 1588 2169
rect 1582 2164 1583 2168
rect 1587 2164 1588 2168
rect 1582 2163 1588 2164
rect 1622 2168 1628 2169
rect 1622 2164 1623 2168
rect 1627 2164 1628 2168
rect 1622 2163 1628 2164
rect 1415 2162 1419 2163
rect 1415 2157 1419 2158
rect 1423 2162 1427 2163
rect 1423 2157 1427 2158
rect 1463 2162 1467 2163
rect 1463 2157 1467 2158
rect 1503 2162 1507 2163
rect 1503 2157 1507 2158
rect 1519 2162 1523 2163
rect 1519 2157 1523 2158
rect 1543 2162 1547 2163
rect 1543 2157 1547 2158
rect 1575 2162 1579 2163
rect 1575 2157 1579 2158
rect 1583 2162 1587 2163
rect 1583 2157 1587 2158
rect 1623 2162 1627 2163
rect 1623 2157 1627 2158
rect 1414 2156 1420 2157
rect 1414 2152 1415 2156
rect 1419 2152 1420 2156
rect 1414 2151 1420 2152
rect 1462 2156 1468 2157
rect 1462 2152 1463 2156
rect 1467 2152 1468 2156
rect 1462 2151 1468 2152
rect 1518 2156 1524 2157
rect 1518 2152 1519 2156
rect 1523 2152 1524 2156
rect 1518 2151 1524 2152
rect 1574 2156 1580 2157
rect 1574 2152 1575 2156
rect 1579 2152 1580 2156
rect 1574 2151 1580 2152
rect 1622 2156 1628 2157
rect 1622 2152 1623 2156
rect 1627 2152 1628 2156
rect 1622 2151 1628 2152
rect 1648 2140 1650 2206
rect 1664 2197 1666 2209
rect 1678 2203 1684 2204
rect 1678 2199 1679 2203
rect 1683 2199 1684 2203
rect 1678 2198 1684 2199
rect 1662 2196 1668 2197
rect 1662 2192 1663 2196
rect 1667 2192 1668 2196
rect 1662 2191 1668 2192
rect 1680 2184 1682 2198
rect 1704 2197 1706 2209
rect 1718 2203 1724 2204
rect 1718 2199 1719 2203
rect 1723 2199 1724 2203
rect 1718 2198 1724 2199
rect 1702 2196 1708 2197
rect 1702 2192 1703 2196
rect 1707 2192 1708 2196
rect 1702 2191 1708 2192
rect 1720 2184 1722 2198
rect 1744 2197 1746 2209
rect 1758 2203 1764 2204
rect 1758 2199 1759 2203
rect 1763 2199 1764 2203
rect 1758 2198 1764 2199
rect 1742 2196 1748 2197
rect 1742 2192 1743 2196
rect 1747 2192 1748 2196
rect 1742 2191 1748 2192
rect 1760 2184 1762 2198
rect 1784 2197 1786 2209
rect 1798 2203 1804 2204
rect 1798 2199 1799 2203
rect 1803 2199 1804 2203
rect 1798 2198 1804 2199
rect 1782 2196 1788 2197
rect 1782 2192 1783 2196
rect 1787 2192 1788 2196
rect 1782 2191 1788 2192
rect 1800 2184 1802 2198
rect 1824 2197 1826 2209
rect 1838 2203 1844 2204
rect 1838 2199 1839 2203
rect 1843 2199 1844 2203
rect 1838 2198 1844 2199
rect 1822 2196 1828 2197
rect 1822 2192 1823 2196
rect 1827 2192 1828 2196
rect 1822 2191 1828 2192
rect 1840 2184 1842 2198
rect 2120 2189 2122 2209
rect 2118 2188 2124 2189
rect 2118 2184 2119 2188
rect 2123 2184 2124 2188
rect 1678 2183 1684 2184
rect 1678 2179 1679 2183
rect 1683 2179 1684 2183
rect 1678 2178 1684 2179
rect 1718 2183 1724 2184
rect 1718 2179 1719 2183
rect 1723 2179 1724 2183
rect 1718 2178 1724 2179
rect 1758 2183 1764 2184
rect 1758 2179 1759 2183
rect 1763 2179 1764 2183
rect 1758 2178 1764 2179
rect 1798 2183 1804 2184
rect 1798 2179 1799 2183
rect 1803 2179 1804 2183
rect 1798 2178 1804 2179
rect 1838 2183 1844 2184
rect 2118 2183 2124 2184
rect 1838 2179 1839 2183
rect 1843 2179 1844 2183
rect 1838 2178 1844 2179
rect 2118 2171 2124 2172
rect 1662 2168 1668 2169
rect 1662 2164 1663 2168
rect 1667 2164 1668 2168
rect 1662 2163 1668 2164
rect 1702 2168 1708 2169
rect 1702 2164 1703 2168
rect 1707 2164 1708 2168
rect 1702 2163 1708 2164
rect 1742 2168 1748 2169
rect 1742 2164 1743 2168
rect 1747 2164 1748 2168
rect 1742 2163 1748 2164
rect 1782 2168 1788 2169
rect 1782 2164 1783 2168
rect 1787 2164 1788 2168
rect 1782 2163 1788 2164
rect 1822 2168 1828 2169
rect 1822 2164 1823 2168
rect 1827 2164 1828 2168
rect 2118 2167 2119 2171
rect 2123 2167 2124 2171
rect 2118 2166 2124 2167
rect 1822 2163 1828 2164
rect 2120 2163 2122 2166
rect 1663 2162 1667 2163
rect 1663 2157 1667 2158
rect 1671 2162 1675 2163
rect 1671 2157 1675 2158
rect 1703 2162 1707 2163
rect 1703 2157 1707 2158
rect 1719 2162 1723 2163
rect 1719 2157 1723 2158
rect 1743 2162 1747 2163
rect 1743 2157 1747 2158
rect 1775 2162 1779 2163
rect 1775 2157 1779 2158
rect 1783 2162 1787 2163
rect 1783 2157 1787 2158
rect 1823 2162 1827 2163
rect 1823 2157 1827 2158
rect 1831 2162 1835 2163
rect 1831 2157 1835 2158
rect 1887 2162 1891 2163
rect 1887 2157 1891 2158
rect 2119 2162 2123 2163
rect 2119 2157 2123 2158
rect 1670 2156 1676 2157
rect 1670 2152 1671 2156
rect 1675 2152 1676 2156
rect 1670 2151 1676 2152
rect 1718 2156 1724 2157
rect 1718 2152 1719 2156
rect 1723 2152 1724 2156
rect 1718 2151 1724 2152
rect 1774 2156 1780 2157
rect 1774 2152 1775 2156
rect 1779 2152 1780 2156
rect 1774 2151 1780 2152
rect 1830 2156 1836 2157
rect 1830 2152 1831 2156
rect 1835 2152 1836 2156
rect 1830 2151 1836 2152
rect 1886 2156 1892 2157
rect 1886 2152 1887 2156
rect 1891 2152 1892 2156
rect 2120 2154 2122 2157
rect 1886 2151 1892 2152
rect 2118 2153 2124 2154
rect 2118 2149 2119 2153
rect 2123 2149 2124 2153
rect 2118 2148 2124 2149
rect 1646 2139 1652 2140
rect 1646 2135 1647 2139
rect 1651 2135 1652 2139
rect 1646 2134 1652 2135
rect 1706 2139 1712 2140
rect 1706 2135 1707 2139
rect 1711 2135 1712 2139
rect 1706 2134 1712 2135
rect 1754 2139 1760 2140
rect 1754 2135 1755 2139
rect 1759 2135 1760 2139
rect 1754 2134 1760 2135
rect 1810 2139 1816 2140
rect 1810 2135 1811 2139
rect 1815 2135 1816 2139
rect 1810 2134 1816 2135
rect 2118 2136 2124 2137
rect 1414 2128 1420 2129
rect 1414 2124 1415 2128
rect 1419 2124 1420 2128
rect 1414 2123 1420 2124
rect 1462 2128 1468 2129
rect 1462 2124 1463 2128
rect 1467 2124 1468 2128
rect 1462 2123 1468 2124
rect 1518 2128 1524 2129
rect 1518 2124 1519 2128
rect 1523 2124 1524 2128
rect 1518 2123 1524 2124
rect 1574 2128 1580 2129
rect 1574 2124 1575 2128
rect 1579 2124 1580 2128
rect 1574 2123 1580 2124
rect 1622 2128 1628 2129
rect 1622 2124 1623 2128
rect 1627 2124 1628 2128
rect 1622 2123 1628 2124
rect 1670 2128 1676 2129
rect 1670 2124 1671 2128
rect 1675 2124 1676 2128
rect 1670 2123 1676 2124
rect 1390 2111 1396 2112
rect 1390 2107 1391 2111
rect 1395 2107 1396 2111
rect 1416 2107 1418 2123
rect 1464 2107 1466 2123
rect 1520 2107 1522 2123
rect 1576 2107 1578 2123
rect 1607 2116 1611 2117
rect 1607 2111 1611 2112
rect 1135 2106 1139 2107
rect 1135 2101 1139 2102
rect 1223 2106 1227 2107
rect 1223 2101 1227 2102
rect 1279 2106 1283 2107
rect 1279 2101 1283 2102
rect 1287 2106 1291 2107
rect 1287 2101 1291 2102
rect 1327 2106 1331 2107
rect 1327 2101 1331 2102
rect 1343 2106 1347 2107
rect 1343 2101 1347 2102
rect 1367 2106 1371 2107
rect 1390 2106 1396 2107
rect 1415 2106 1419 2107
rect 1367 2101 1371 2102
rect 1415 2101 1419 2102
rect 1423 2106 1427 2107
rect 1423 2101 1427 2102
rect 1463 2106 1467 2107
rect 1463 2101 1467 2102
rect 1503 2106 1507 2107
rect 1503 2101 1507 2102
rect 1519 2106 1523 2107
rect 1519 2101 1523 2102
rect 1575 2106 1579 2107
rect 1575 2101 1579 2102
rect 1583 2106 1587 2107
rect 1583 2101 1587 2102
rect 1136 2081 1138 2101
rect 1224 2089 1226 2101
rect 1280 2089 1282 2101
rect 1294 2095 1300 2096
rect 1294 2091 1295 2095
rect 1299 2091 1300 2095
rect 1294 2090 1300 2091
rect 1222 2088 1228 2089
rect 1222 2084 1223 2088
rect 1227 2084 1228 2088
rect 1222 2083 1228 2084
rect 1278 2088 1284 2089
rect 1278 2084 1279 2088
rect 1283 2084 1284 2088
rect 1278 2083 1284 2084
rect 1134 2080 1140 2081
rect 1134 2076 1135 2080
rect 1139 2076 1140 2080
rect 1296 2076 1298 2090
rect 1344 2089 1346 2101
rect 1350 2095 1356 2096
rect 1350 2091 1351 2095
rect 1355 2091 1356 2095
rect 1350 2090 1356 2091
rect 1342 2088 1348 2089
rect 1342 2084 1343 2088
rect 1347 2084 1348 2088
rect 1342 2083 1348 2084
rect 1352 2076 1354 2090
rect 1424 2089 1426 2101
rect 1438 2095 1444 2096
rect 1438 2091 1439 2095
rect 1443 2091 1444 2095
rect 1438 2090 1444 2091
rect 1422 2088 1428 2089
rect 1422 2084 1423 2088
rect 1427 2084 1428 2088
rect 1422 2083 1428 2084
rect 1440 2076 1442 2090
rect 1504 2089 1506 2101
rect 1518 2095 1524 2096
rect 1518 2091 1519 2095
rect 1523 2091 1524 2095
rect 1518 2090 1524 2091
rect 1502 2088 1508 2089
rect 1502 2084 1503 2088
rect 1507 2084 1508 2088
rect 1502 2083 1508 2084
rect 1520 2076 1522 2090
rect 1584 2089 1586 2101
rect 1608 2096 1610 2111
rect 1624 2107 1626 2123
rect 1672 2107 1674 2123
rect 1708 2120 1710 2134
rect 1718 2128 1724 2129
rect 1718 2124 1719 2128
rect 1723 2124 1724 2128
rect 1718 2123 1724 2124
rect 1706 2119 1712 2120
rect 1706 2115 1707 2119
rect 1711 2115 1712 2119
rect 1706 2114 1712 2115
rect 1690 2111 1696 2112
rect 1690 2107 1691 2111
rect 1695 2107 1696 2111
rect 1720 2107 1722 2123
rect 1756 2120 1758 2134
rect 1774 2128 1780 2129
rect 1774 2124 1775 2128
rect 1779 2124 1780 2128
rect 1774 2123 1780 2124
rect 1754 2119 1760 2120
rect 1754 2115 1755 2119
rect 1759 2115 1760 2119
rect 1754 2114 1760 2115
rect 1776 2107 1778 2123
rect 1812 2120 1814 2134
rect 2118 2132 2119 2136
rect 2123 2132 2124 2136
rect 2118 2131 2124 2132
rect 1830 2128 1836 2129
rect 1830 2124 1831 2128
rect 1835 2124 1836 2128
rect 1830 2123 1836 2124
rect 1886 2128 1892 2129
rect 1886 2124 1887 2128
rect 1891 2124 1892 2128
rect 1886 2123 1892 2124
rect 1810 2119 1816 2120
rect 1810 2115 1811 2119
rect 1815 2115 1816 2119
rect 1810 2114 1816 2115
rect 1832 2107 1834 2123
rect 1888 2107 1890 2123
rect 2120 2107 2122 2131
rect 1623 2106 1627 2107
rect 1623 2101 1627 2102
rect 1663 2106 1667 2107
rect 1663 2101 1667 2102
rect 1671 2106 1675 2107
rect 1690 2106 1696 2107
rect 1719 2106 1723 2107
rect 1671 2101 1675 2102
rect 1598 2095 1604 2096
rect 1598 2091 1599 2095
rect 1603 2091 1604 2095
rect 1598 2090 1604 2091
rect 1606 2095 1612 2096
rect 1606 2091 1607 2095
rect 1611 2091 1612 2095
rect 1606 2090 1612 2091
rect 1582 2088 1588 2089
rect 1582 2084 1583 2088
rect 1587 2084 1588 2088
rect 1582 2083 1588 2084
rect 1600 2076 1602 2090
rect 1664 2089 1666 2101
rect 1662 2088 1668 2089
rect 1662 2084 1663 2088
rect 1667 2084 1668 2088
rect 1662 2083 1668 2084
rect 1692 2076 1694 2106
rect 1719 2101 1723 2102
rect 1743 2106 1747 2107
rect 1743 2101 1747 2102
rect 1775 2106 1779 2107
rect 1775 2101 1779 2102
rect 1831 2106 1835 2107
rect 1831 2101 1835 2102
rect 1887 2106 1891 2107
rect 1887 2101 1891 2102
rect 1919 2106 1923 2107
rect 1919 2101 1923 2102
rect 2007 2106 2011 2107
rect 2007 2101 2011 2102
rect 2071 2106 2075 2107
rect 2071 2101 2075 2102
rect 2119 2106 2123 2107
rect 2119 2101 2123 2102
rect 1744 2089 1746 2101
rect 1758 2095 1764 2096
rect 1758 2091 1759 2095
rect 1763 2091 1764 2095
rect 1758 2090 1764 2091
rect 1742 2088 1748 2089
rect 1742 2084 1743 2088
rect 1747 2084 1748 2088
rect 1742 2083 1748 2084
rect 1760 2076 1762 2090
rect 1832 2089 1834 2101
rect 1846 2095 1852 2096
rect 1846 2091 1847 2095
rect 1851 2091 1852 2095
rect 1846 2090 1852 2091
rect 1830 2088 1836 2089
rect 1830 2084 1831 2088
rect 1835 2084 1836 2088
rect 1830 2083 1836 2084
rect 1848 2076 1850 2090
rect 1920 2089 1922 2101
rect 1934 2095 1940 2096
rect 1934 2091 1935 2095
rect 1939 2091 1940 2095
rect 1934 2090 1940 2091
rect 1918 2088 1924 2089
rect 1918 2084 1919 2088
rect 1923 2084 1924 2088
rect 1918 2083 1924 2084
rect 1936 2076 1938 2090
rect 2008 2089 2010 2101
rect 2022 2095 2028 2096
rect 2022 2091 2023 2095
rect 2027 2091 2028 2095
rect 2022 2090 2028 2091
rect 2030 2095 2036 2096
rect 2030 2091 2031 2095
rect 2035 2091 2036 2095
rect 2030 2090 2036 2091
rect 2006 2088 2012 2089
rect 2006 2084 2007 2088
rect 2011 2084 2012 2088
rect 2006 2083 2012 2084
rect 2024 2076 2026 2090
rect 1134 2075 1140 2076
rect 1210 2075 1216 2076
rect 1210 2071 1211 2075
rect 1215 2071 1216 2075
rect 1210 2070 1216 2071
rect 1294 2075 1300 2076
rect 1294 2071 1295 2075
rect 1299 2071 1300 2075
rect 1294 2070 1300 2071
rect 1350 2075 1356 2076
rect 1350 2071 1351 2075
rect 1355 2071 1356 2075
rect 1350 2070 1356 2071
rect 1438 2075 1444 2076
rect 1438 2071 1439 2075
rect 1443 2071 1444 2075
rect 1438 2070 1444 2071
rect 1518 2075 1524 2076
rect 1518 2071 1519 2075
rect 1523 2071 1524 2075
rect 1518 2070 1524 2071
rect 1598 2075 1604 2076
rect 1598 2071 1599 2075
rect 1603 2071 1604 2075
rect 1598 2070 1604 2071
rect 1690 2075 1696 2076
rect 1690 2071 1691 2075
rect 1695 2071 1696 2075
rect 1690 2070 1696 2071
rect 1758 2075 1764 2076
rect 1758 2071 1759 2075
rect 1763 2071 1764 2075
rect 1758 2070 1764 2071
rect 1846 2075 1852 2076
rect 1846 2071 1847 2075
rect 1851 2071 1852 2075
rect 1846 2070 1852 2071
rect 1934 2075 1940 2076
rect 1934 2071 1935 2075
rect 1939 2071 1940 2075
rect 1934 2070 1940 2071
rect 2022 2075 2028 2076
rect 2022 2071 2023 2075
rect 2027 2071 2028 2075
rect 2022 2070 2028 2071
rect 1134 2063 1140 2064
rect 1134 2059 1135 2063
rect 1139 2059 1140 2063
rect 1134 2058 1140 2059
rect 1136 2055 1138 2058
rect 1135 2054 1139 2055
rect 1135 2049 1139 2050
rect 1183 2054 1187 2055
rect 1183 2049 1187 2050
rect 1136 2046 1138 2049
rect 1182 2048 1188 2049
rect 1134 2045 1140 2046
rect 1134 2041 1135 2045
rect 1139 2041 1140 2045
rect 1182 2044 1183 2048
rect 1187 2044 1188 2048
rect 1182 2043 1188 2044
rect 1134 2040 1140 2041
rect 111 2034 115 2035
rect 111 2029 115 2030
rect 191 2034 195 2035
rect 191 2029 195 2030
rect 231 2034 235 2035
rect 231 2029 235 2030
rect 287 2034 291 2035
rect 287 2029 291 2030
rect 351 2034 355 2035
rect 351 2029 355 2030
rect 423 2034 427 2035
rect 423 2029 427 2030
rect 495 2034 499 2035
rect 495 2029 499 2030
rect 575 2034 579 2035
rect 575 2029 579 2030
rect 647 2034 651 2035
rect 647 2029 651 2030
rect 719 2034 723 2035
rect 719 2029 723 2030
rect 783 2034 787 2035
rect 783 2029 787 2030
rect 839 2034 843 2035
rect 839 2029 843 2030
rect 895 2034 899 2035
rect 895 2029 899 2030
rect 951 2034 955 2035
rect 951 2029 955 2030
rect 1007 2034 1011 2035
rect 1007 2029 1011 2030
rect 1047 2034 1051 2035
rect 1047 2029 1051 2030
rect 1095 2034 1099 2035
rect 1095 2029 1099 2030
rect 112 2009 114 2029
rect 192 2017 194 2029
rect 232 2017 234 2029
rect 246 2023 252 2024
rect 246 2019 247 2023
rect 251 2019 252 2023
rect 246 2018 252 2019
rect 190 2016 196 2017
rect 190 2012 191 2016
rect 195 2012 196 2016
rect 190 2011 196 2012
rect 230 2016 236 2017
rect 230 2012 231 2016
rect 235 2012 236 2016
rect 230 2011 236 2012
rect 110 2008 116 2009
rect 110 2004 111 2008
rect 115 2004 116 2008
rect 248 2004 250 2018
rect 288 2017 290 2029
rect 302 2023 308 2024
rect 302 2019 303 2023
rect 307 2019 308 2023
rect 302 2018 308 2019
rect 286 2016 292 2017
rect 286 2012 287 2016
rect 291 2012 292 2016
rect 286 2011 292 2012
rect 304 2004 306 2018
rect 352 2017 354 2029
rect 366 2023 372 2024
rect 366 2019 367 2023
rect 371 2019 372 2023
rect 366 2018 372 2019
rect 350 2016 356 2017
rect 350 2012 351 2016
rect 355 2012 356 2016
rect 350 2011 356 2012
rect 368 2004 370 2018
rect 424 2017 426 2029
rect 438 2023 444 2024
rect 438 2019 439 2023
rect 443 2019 444 2023
rect 438 2018 444 2019
rect 422 2016 428 2017
rect 422 2012 423 2016
rect 427 2012 428 2016
rect 422 2011 428 2012
rect 440 2004 442 2018
rect 496 2017 498 2029
rect 510 2023 516 2024
rect 510 2019 511 2023
rect 515 2019 516 2023
rect 510 2018 516 2019
rect 538 2023 544 2024
rect 538 2019 539 2023
rect 543 2019 544 2023
rect 538 2018 544 2019
rect 546 2023 552 2024
rect 546 2019 547 2023
rect 551 2019 552 2023
rect 546 2018 552 2019
rect 494 2016 500 2017
rect 494 2012 495 2016
rect 499 2012 500 2016
rect 494 2011 500 2012
rect 512 2004 514 2018
rect 540 2004 542 2018
rect 110 2003 116 2004
rect 214 2003 220 2004
rect 214 1999 215 2003
rect 219 1999 220 2003
rect 214 1998 220 1999
rect 246 2003 252 2004
rect 246 1999 247 2003
rect 251 1999 252 2003
rect 246 1998 252 1999
rect 302 2003 308 2004
rect 302 1999 303 2003
rect 307 1999 308 2003
rect 302 1998 308 1999
rect 366 2003 372 2004
rect 366 1999 367 2003
rect 371 1999 372 2003
rect 366 1998 372 1999
rect 438 2003 444 2004
rect 438 1999 439 2003
rect 443 1999 444 2003
rect 438 1998 444 1999
rect 510 2003 516 2004
rect 510 1999 511 2003
rect 515 1999 516 2003
rect 510 1998 516 1999
rect 538 2003 544 2004
rect 538 1999 539 2003
rect 543 1999 544 2003
rect 538 1998 544 1999
rect 110 1991 116 1992
rect 110 1987 111 1991
rect 115 1987 116 1991
rect 110 1986 116 1987
rect 190 1988 196 1989
rect 112 1983 114 1986
rect 190 1984 191 1988
rect 195 1984 196 1988
rect 190 1983 196 1984
rect 111 1982 115 1983
rect 111 1977 115 1978
rect 191 1982 195 1983
rect 191 1977 195 1978
rect 112 1974 114 1977
rect 190 1976 196 1977
rect 110 1973 116 1974
rect 110 1969 111 1973
rect 115 1969 116 1973
rect 190 1972 191 1976
rect 195 1972 196 1976
rect 190 1971 196 1972
rect 110 1968 116 1969
rect 110 1956 116 1957
rect 110 1952 111 1956
rect 115 1952 116 1956
rect 110 1951 116 1952
rect 112 1931 114 1951
rect 190 1948 196 1949
rect 190 1944 191 1948
rect 195 1944 196 1948
rect 190 1943 196 1944
rect 192 1931 194 1943
rect 216 1940 218 1998
rect 230 1988 236 1989
rect 230 1984 231 1988
rect 235 1984 236 1988
rect 230 1983 236 1984
rect 286 1988 292 1989
rect 286 1984 287 1988
rect 291 1984 292 1988
rect 286 1983 292 1984
rect 350 1988 356 1989
rect 350 1984 351 1988
rect 355 1984 356 1988
rect 350 1983 356 1984
rect 422 1988 428 1989
rect 422 1984 423 1988
rect 427 1984 428 1988
rect 422 1983 428 1984
rect 494 1988 500 1989
rect 494 1984 495 1988
rect 499 1984 500 1988
rect 494 1983 500 1984
rect 231 1982 235 1983
rect 231 1977 235 1978
rect 247 1982 251 1983
rect 247 1977 251 1978
rect 287 1982 291 1983
rect 287 1977 291 1978
rect 311 1982 315 1983
rect 311 1977 315 1978
rect 351 1982 355 1983
rect 351 1977 355 1978
rect 375 1982 379 1983
rect 375 1977 379 1978
rect 423 1982 427 1983
rect 423 1977 427 1978
rect 447 1982 451 1983
rect 447 1977 451 1978
rect 495 1982 499 1983
rect 495 1977 499 1978
rect 519 1982 523 1983
rect 519 1977 523 1978
rect 246 1976 252 1977
rect 246 1972 247 1976
rect 251 1972 252 1976
rect 246 1971 252 1972
rect 310 1976 316 1977
rect 310 1972 311 1976
rect 315 1972 316 1976
rect 310 1971 316 1972
rect 374 1976 380 1977
rect 374 1972 375 1976
rect 379 1972 380 1976
rect 374 1971 380 1972
rect 446 1976 452 1977
rect 446 1972 447 1976
rect 451 1972 452 1976
rect 446 1971 452 1972
rect 518 1976 524 1977
rect 518 1972 519 1976
rect 523 1972 524 1976
rect 518 1971 524 1972
rect 548 1960 550 2018
rect 576 2017 578 2029
rect 648 2017 650 2029
rect 720 2017 722 2029
rect 734 2023 740 2024
rect 734 2019 735 2023
rect 739 2019 740 2023
rect 734 2018 740 2019
rect 574 2016 580 2017
rect 574 2012 575 2016
rect 579 2012 580 2016
rect 574 2011 580 2012
rect 646 2016 652 2017
rect 646 2012 647 2016
rect 651 2012 652 2016
rect 646 2011 652 2012
rect 718 2016 724 2017
rect 718 2012 719 2016
rect 723 2012 724 2016
rect 718 2011 724 2012
rect 736 2004 738 2018
rect 784 2017 786 2029
rect 790 2023 796 2024
rect 790 2019 791 2023
rect 795 2019 796 2023
rect 790 2018 796 2019
rect 782 2016 788 2017
rect 782 2012 783 2016
rect 787 2012 788 2016
rect 782 2011 788 2012
rect 792 2004 794 2018
rect 840 2017 842 2029
rect 854 2023 860 2024
rect 854 2019 855 2023
rect 859 2019 860 2023
rect 854 2018 860 2019
rect 838 2016 844 2017
rect 838 2012 839 2016
rect 843 2012 844 2016
rect 838 2011 844 2012
rect 856 2004 858 2018
rect 896 2017 898 2029
rect 910 2023 916 2024
rect 910 2019 911 2023
rect 915 2019 916 2023
rect 910 2018 916 2019
rect 894 2016 900 2017
rect 894 2012 895 2016
rect 899 2012 900 2016
rect 894 2011 900 2012
rect 912 2004 914 2018
rect 952 2017 954 2029
rect 966 2023 972 2024
rect 966 2019 967 2023
rect 971 2019 972 2023
rect 966 2018 972 2019
rect 950 2016 956 2017
rect 950 2012 951 2016
rect 955 2012 956 2016
rect 950 2011 956 2012
rect 968 2004 970 2018
rect 1008 2017 1010 2029
rect 1022 2023 1028 2024
rect 1022 2019 1023 2023
rect 1027 2019 1028 2023
rect 1022 2018 1028 2019
rect 1006 2016 1012 2017
rect 1006 2012 1007 2016
rect 1011 2012 1012 2016
rect 1006 2011 1012 2012
rect 1024 2004 1026 2018
rect 1048 2017 1050 2029
rect 1062 2023 1068 2024
rect 1062 2019 1063 2023
rect 1067 2019 1068 2023
rect 1062 2018 1068 2019
rect 1070 2023 1076 2024
rect 1070 2019 1071 2023
rect 1075 2019 1076 2023
rect 1070 2018 1076 2019
rect 1046 2016 1052 2017
rect 1046 2012 1047 2016
rect 1051 2012 1052 2016
rect 1046 2011 1052 2012
rect 1064 2004 1066 2018
rect 734 2003 740 2004
rect 734 1999 735 2003
rect 739 1999 740 2003
rect 734 1998 740 1999
rect 790 2003 796 2004
rect 790 1999 791 2003
rect 795 1999 796 2003
rect 790 1998 796 1999
rect 854 2003 860 2004
rect 854 1999 855 2003
rect 859 1999 860 2003
rect 854 1998 860 1999
rect 910 2003 916 2004
rect 910 1999 911 2003
rect 915 1999 916 2003
rect 910 1998 916 1999
rect 966 2003 972 2004
rect 966 1999 967 2003
rect 971 1999 972 2003
rect 966 1998 972 1999
rect 1022 2003 1028 2004
rect 1022 1999 1023 2003
rect 1027 1999 1028 2003
rect 1022 1998 1028 1999
rect 1062 2003 1068 2004
rect 1062 1999 1063 2003
rect 1067 1999 1068 2003
rect 1062 1998 1068 1999
rect 574 1988 580 1989
rect 574 1984 575 1988
rect 579 1984 580 1988
rect 574 1983 580 1984
rect 646 1988 652 1989
rect 646 1984 647 1988
rect 651 1984 652 1988
rect 646 1983 652 1984
rect 718 1988 724 1989
rect 718 1984 719 1988
rect 723 1984 724 1988
rect 718 1983 724 1984
rect 782 1988 788 1989
rect 782 1984 783 1988
rect 787 1984 788 1988
rect 782 1983 788 1984
rect 838 1988 844 1989
rect 838 1984 839 1988
rect 843 1984 844 1988
rect 838 1983 844 1984
rect 894 1988 900 1989
rect 894 1984 895 1988
rect 899 1984 900 1988
rect 894 1983 900 1984
rect 950 1988 956 1989
rect 950 1984 951 1988
rect 955 1984 956 1988
rect 950 1983 956 1984
rect 1006 1988 1012 1989
rect 1006 1984 1007 1988
rect 1011 1984 1012 1988
rect 1006 1983 1012 1984
rect 1046 1988 1052 1989
rect 1046 1984 1047 1988
rect 1051 1984 1052 1988
rect 1046 1983 1052 1984
rect 575 1982 579 1983
rect 575 1977 579 1978
rect 591 1982 595 1983
rect 591 1977 595 1978
rect 647 1982 651 1983
rect 647 1977 651 1978
rect 655 1982 659 1983
rect 655 1977 659 1978
rect 719 1982 723 1983
rect 719 1977 723 1978
rect 775 1982 779 1983
rect 775 1977 779 1978
rect 783 1982 787 1983
rect 783 1977 787 1978
rect 823 1982 827 1983
rect 823 1977 827 1978
rect 839 1982 843 1983
rect 839 1977 843 1978
rect 871 1982 875 1983
rect 871 1977 875 1978
rect 895 1982 899 1983
rect 895 1977 899 1978
rect 919 1982 923 1983
rect 919 1977 923 1978
rect 951 1982 955 1983
rect 951 1977 955 1978
rect 967 1982 971 1983
rect 967 1977 971 1978
rect 1007 1982 1011 1983
rect 1007 1977 1011 1978
rect 1047 1982 1051 1983
rect 1047 1977 1051 1978
rect 590 1976 596 1977
rect 590 1972 591 1976
rect 595 1972 596 1976
rect 590 1971 596 1972
rect 654 1976 660 1977
rect 654 1972 655 1976
rect 659 1972 660 1976
rect 654 1971 660 1972
rect 718 1976 724 1977
rect 718 1972 719 1976
rect 723 1972 724 1976
rect 718 1971 724 1972
rect 774 1976 780 1977
rect 774 1972 775 1976
rect 779 1972 780 1976
rect 774 1971 780 1972
rect 822 1976 828 1977
rect 822 1972 823 1976
rect 827 1972 828 1976
rect 822 1971 828 1972
rect 870 1976 876 1977
rect 870 1972 871 1976
rect 875 1972 876 1976
rect 870 1971 876 1972
rect 918 1976 924 1977
rect 918 1972 919 1976
rect 923 1972 924 1976
rect 918 1971 924 1972
rect 966 1976 972 1977
rect 966 1972 967 1976
rect 971 1972 972 1976
rect 966 1971 972 1972
rect 1006 1976 1012 1977
rect 1006 1972 1007 1976
rect 1011 1972 1012 1976
rect 1006 1971 1012 1972
rect 1046 1976 1052 1977
rect 1046 1972 1047 1976
rect 1051 1972 1052 1976
rect 1046 1971 1052 1972
rect 1072 1968 1074 2018
rect 1096 2009 1098 2029
rect 1134 2028 1140 2029
rect 1134 2024 1135 2028
rect 1139 2024 1140 2028
rect 1134 2023 1140 2024
rect 1094 2008 1100 2009
rect 1094 2004 1095 2008
rect 1099 2004 1100 2008
rect 1094 2003 1100 2004
rect 1136 2003 1138 2023
rect 1182 2020 1188 2021
rect 1182 2016 1183 2020
rect 1187 2016 1188 2020
rect 1182 2015 1188 2016
rect 1184 2003 1186 2015
rect 1212 2012 1214 2070
rect 1222 2060 1228 2061
rect 1222 2056 1223 2060
rect 1227 2056 1228 2060
rect 1222 2055 1228 2056
rect 1278 2060 1284 2061
rect 1278 2056 1279 2060
rect 1283 2056 1284 2060
rect 1278 2055 1284 2056
rect 1342 2060 1348 2061
rect 1342 2056 1343 2060
rect 1347 2056 1348 2060
rect 1342 2055 1348 2056
rect 1422 2060 1428 2061
rect 1422 2056 1423 2060
rect 1427 2056 1428 2060
rect 1422 2055 1428 2056
rect 1502 2060 1508 2061
rect 1502 2056 1503 2060
rect 1507 2056 1508 2060
rect 1502 2055 1508 2056
rect 1582 2060 1588 2061
rect 1582 2056 1583 2060
rect 1587 2056 1588 2060
rect 1582 2055 1588 2056
rect 1662 2060 1668 2061
rect 1662 2056 1663 2060
rect 1667 2056 1668 2060
rect 1662 2055 1668 2056
rect 1742 2060 1748 2061
rect 1742 2056 1743 2060
rect 1747 2056 1748 2060
rect 1742 2055 1748 2056
rect 1830 2060 1836 2061
rect 1830 2056 1831 2060
rect 1835 2056 1836 2060
rect 1830 2055 1836 2056
rect 1918 2060 1924 2061
rect 1918 2056 1919 2060
rect 1923 2056 1924 2060
rect 1918 2055 1924 2056
rect 2006 2060 2012 2061
rect 2006 2056 2007 2060
rect 2011 2056 2012 2060
rect 2006 2055 2012 2056
rect 1223 2054 1227 2055
rect 1223 2049 1227 2050
rect 1239 2054 1243 2055
rect 1239 2049 1243 2050
rect 1279 2054 1283 2055
rect 1279 2049 1283 2050
rect 1311 2054 1315 2055
rect 1311 2049 1315 2050
rect 1343 2054 1347 2055
rect 1343 2049 1347 2050
rect 1399 2054 1403 2055
rect 1399 2049 1403 2050
rect 1423 2054 1427 2055
rect 1423 2049 1427 2050
rect 1487 2054 1491 2055
rect 1487 2049 1491 2050
rect 1503 2054 1507 2055
rect 1503 2049 1507 2050
rect 1583 2054 1587 2055
rect 1583 2049 1587 2050
rect 1663 2054 1667 2055
rect 1663 2049 1667 2050
rect 1671 2054 1675 2055
rect 1671 2049 1675 2050
rect 1743 2054 1747 2055
rect 1743 2049 1747 2050
rect 1759 2054 1763 2055
rect 1759 2049 1763 2050
rect 1831 2054 1835 2055
rect 1831 2049 1835 2050
rect 1839 2054 1843 2055
rect 1839 2049 1843 2050
rect 1919 2054 1923 2055
rect 1919 2049 1923 2050
rect 2007 2054 2011 2055
rect 2007 2049 2011 2050
rect 1238 2048 1244 2049
rect 1238 2044 1239 2048
rect 1243 2044 1244 2048
rect 1238 2043 1244 2044
rect 1310 2048 1316 2049
rect 1310 2044 1311 2048
rect 1315 2044 1316 2048
rect 1310 2043 1316 2044
rect 1398 2048 1404 2049
rect 1398 2044 1399 2048
rect 1403 2044 1404 2048
rect 1398 2043 1404 2044
rect 1486 2048 1492 2049
rect 1486 2044 1487 2048
rect 1491 2044 1492 2048
rect 1486 2043 1492 2044
rect 1582 2048 1588 2049
rect 1582 2044 1583 2048
rect 1587 2044 1588 2048
rect 1582 2043 1588 2044
rect 1670 2048 1676 2049
rect 1670 2044 1671 2048
rect 1675 2044 1676 2048
rect 1670 2043 1676 2044
rect 1758 2048 1764 2049
rect 1758 2044 1759 2048
rect 1763 2044 1764 2048
rect 1758 2043 1764 2044
rect 1838 2048 1844 2049
rect 1838 2044 1839 2048
rect 1843 2044 1844 2048
rect 1838 2043 1844 2044
rect 1918 2048 1924 2049
rect 1918 2044 1919 2048
rect 1923 2044 1924 2048
rect 1918 2043 1924 2044
rect 2006 2048 2012 2049
rect 2006 2044 2007 2048
rect 2011 2044 2012 2048
rect 2006 2043 2012 2044
rect 1862 2039 1868 2040
rect 1862 2035 1863 2039
rect 1867 2035 1868 2039
rect 1862 2034 1868 2035
rect 1254 2031 1260 2032
rect 1254 2027 1255 2031
rect 1259 2027 1260 2031
rect 1254 2026 1260 2027
rect 1326 2031 1332 2032
rect 1326 2027 1327 2031
rect 1331 2027 1332 2031
rect 1326 2026 1332 2027
rect 1414 2031 1420 2032
rect 1414 2027 1415 2031
rect 1419 2027 1420 2031
rect 1414 2026 1420 2027
rect 1502 2031 1508 2032
rect 1502 2027 1503 2031
rect 1507 2027 1508 2031
rect 1502 2026 1508 2027
rect 1558 2031 1564 2032
rect 1558 2027 1559 2031
rect 1563 2027 1564 2031
rect 1558 2026 1564 2027
rect 1570 2031 1576 2032
rect 1570 2027 1571 2031
rect 1575 2027 1576 2031
rect 1570 2026 1576 2027
rect 1238 2020 1244 2021
rect 1238 2016 1239 2020
rect 1243 2016 1244 2020
rect 1238 2015 1244 2016
rect 1210 2011 1216 2012
rect 1210 2007 1211 2011
rect 1215 2007 1216 2011
rect 1210 2006 1216 2007
rect 1240 2003 1242 2015
rect 1256 2012 1258 2026
rect 1310 2020 1316 2021
rect 1310 2016 1311 2020
rect 1315 2016 1316 2020
rect 1310 2015 1316 2016
rect 1254 2011 1260 2012
rect 1254 2007 1255 2011
rect 1259 2007 1260 2011
rect 1254 2006 1260 2007
rect 1312 2003 1314 2015
rect 1328 2012 1330 2026
rect 1398 2020 1404 2021
rect 1398 2016 1399 2020
rect 1403 2016 1404 2020
rect 1398 2015 1404 2016
rect 1326 2011 1332 2012
rect 1326 2007 1327 2011
rect 1331 2007 1332 2011
rect 1326 2006 1332 2007
rect 1400 2003 1402 2015
rect 1416 2012 1418 2026
rect 1486 2020 1492 2021
rect 1486 2016 1487 2020
rect 1491 2016 1492 2020
rect 1486 2015 1492 2016
rect 1414 2011 1420 2012
rect 1414 2007 1415 2011
rect 1419 2007 1420 2011
rect 1414 2006 1420 2007
rect 1488 2003 1490 2015
rect 1504 2012 1506 2026
rect 1560 2012 1562 2026
rect 1502 2011 1508 2012
rect 1502 2007 1503 2011
rect 1507 2007 1508 2011
rect 1502 2006 1508 2007
rect 1558 2011 1564 2012
rect 1558 2007 1559 2011
rect 1563 2007 1564 2011
rect 1558 2006 1564 2007
rect 1135 2002 1139 2003
rect 1135 1997 1139 1998
rect 1183 2002 1187 2003
rect 1183 1997 1187 1998
rect 1239 2002 1243 2003
rect 1239 1997 1243 1998
rect 1303 2002 1307 2003
rect 1303 1997 1307 1998
rect 1311 2002 1315 2003
rect 1311 1997 1315 1998
rect 1383 2002 1387 2003
rect 1383 1997 1387 1998
rect 1399 2002 1403 2003
rect 1399 1997 1403 1998
rect 1463 2002 1467 2003
rect 1463 1997 1467 1998
rect 1487 2002 1491 2003
rect 1487 1997 1491 1998
rect 1543 2002 1547 2003
rect 1543 1997 1547 1998
rect 1094 1991 1100 1992
rect 1094 1987 1095 1991
rect 1099 1987 1100 1991
rect 1094 1986 1100 1987
rect 1096 1983 1098 1986
rect 1095 1982 1099 1983
rect 1095 1977 1099 1978
rect 1136 1977 1138 1997
rect 1304 1985 1306 1997
rect 1384 1985 1386 1997
rect 1398 1991 1404 1992
rect 1398 1987 1399 1991
rect 1403 1987 1404 1991
rect 1398 1986 1404 1987
rect 1302 1984 1308 1985
rect 1302 1980 1303 1984
rect 1307 1980 1308 1984
rect 1302 1979 1308 1980
rect 1382 1984 1388 1985
rect 1382 1980 1383 1984
rect 1387 1980 1388 1984
rect 1382 1979 1388 1980
rect 1096 1974 1098 1977
rect 1134 1976 1140 1977
rect 1094 1973 1100 1974
rect 1094 1969 1095 1973
rect 1099 1969 1100 1973
rect 1134 1972 1135 1976
rect 1139 1972 1140 1976
rect 1400 1972 1402 1986
rect 1464 1985 1466 1997
rect 1478 1991 1484 1992
rect 1478 1987 1479 1991
rect 1483 1987 1484 1991
rect 1478 1986 1484 1987
rect 1462 1984 1468 1985
rect 1462 1980 1463 1984
rect 1467 1980 1468 1984
rect 1462 1979 1468 1980
rect 1480 1972 1482 1986
rect 1544 1985 1546 1997
rect 1572 1992 1574 2026
rect 1582 2020 1588 2021
rect 1582 2016 1583 2020
rect 1587 2016 1588 2020
rect 1582 2015 1588 2016
rect 1670 2020 1676 2021
rect 1670 2016 1671 2020
rect 1675 2016 1676 2020
rect 1670 2015 1676 2016
rect 1758 2020 1764 2021
rect 1758 2016 1759 2020
rect 1763 2016 1764 2020
rect 1758 2015 1764 2016
rect 1838 2020 1844 2021
rect 1838 2016 1839 2020
rect 1843 2016 1844 2020
rect 1838 2015 1844 2016
rect 1584 2003 1586 2015
rect 1672 2003 1674 2015
rect 1760 2003 1762 2015
rect 1830 2011 1836 2012
rect 1830 2007 1831 2011
rect 1835 2007 1836 2011
rect 1830 2006 1836 2007
rect 1583 2002 1587 2003
rect 1583 1997 1587 1998
rect 1615 2002 1619 2003
rect 1615 1997 1619 1998
rect 1671 2002 1675 2003
rect 1671 1997 1675 1998
rect 1687 2002 1691 2003
rect 1687 1997 1691 1998
rect 1751 2002 1755 2003
rect 1751 1997 1755 1998
rect 1759 2002 1763 2003
rect 1759 1997 1763 1998
rect 1815 2002 1819 2003
rect 1815 1997 1819 1998
rect 1550 1991 1556 1992
rect 1550 1987 1551 1991
rect 1555 1987 1556 1991
rect 1550 1986 1556 1987
rect 1570 1991 1576 1992
rect 1570 1987 1571 1991
rect 1575 1987 1576 1991
rect 1570 1986 1576 1987
rect 1542 1984 1548 1985
rect 1542 1980 1543 1984
rect 1547 1980 1548 1984
rect 1542 1979 1548 1980
rect 1552 1972 1554 1986
rect 1616 1985 1618 1997
rect 1688 1985 1690 1997
rect 1694 1991 1700 1992
rect 1694 1987 1695 1991
rect 1699 1987 1700 1991
rect 1694 1986 1700 1987
rect 1614 1984 1620 1985
rect 1614 1980 1615 1984
rect 1619 1980 1620 1984
rect 1686 1984 1692 1985
rect 1614 1979 1620 1980
rect 1643 1980 1647 1981
rect 1686 1980 1687 1984
rect 1691 1980 1692 1984
rect 1686 1979 1692 1980
rect 1643 1975 1647 1976
rect 1644 1972 1646 1975
rect 1696 1972 1698 1986
rect 1752 1985 1754 1997
rect 1766 1991 1772 1992
rect 1766 1987 1767 1991
rect 1771 1987 1772 1991
rect 1766 1986 1772 1987
rect 1806 1991 1812 1992
rect 1806 1987 1807 1991
rect 1811 1987 1812 1991
rect 1806 1986 1812 1987
rect 1750 1984 1756 1985
rect 1750 1980 1751 1984
rect 1755 1980 1756 1984
rect 1750 1979 1756 1980
rect 1768 1972 1770 1986
rect 1134 1971 1140 1972
rect 1326 1971 1332 1972
rect 1094 1968 1100 1969
rect 894 1967 900 1968
rect 894 1963 895 1967
rect 899 1963 900 1967
rect 894 1962 900 1963
rect 1070 1967 1076 1968
rect 1070 1963 1071 1967
rect 1075 1963 1076 1967
rect 1326 1967 1327 1971
rect 1331 1967 1332 1971
rect 1326 1966 1332 1967
rect 1398 1971 1404 1972
rect 1398 1967 1399 1971
rect 1403 1967 1404 1971
rect 1398 1966 1404 1967
rect 1478 1971 1484 1972
rect 1478 1967 1479 1971
rect 1483 1967 1484 1971
rect 1478 1966 1484 1967
rect 1550 1971 1556 1972
rect 1550 1967 1551 1971
rect 1555 1967 1556 1971
rect 1550 1966 1556 1967
rect 1642 1971 1648 1972
rect 1642 1967 1643 1971
rect 1647 1967 1648 1971
rect 1642 1966 1648 1967
rect 1694 1971 1700 1972
rect 1694 1967 1695 1971
rect 1699 1967 1700 1971
rect 1694 1966 1700 1967
rect 1766 1971 1772 1972
rect 1766 1967 1767 1971
rect 1771 1967 1772 1971
rect 1766 1966 1772 1967
rect 1070 1962 1076 1963
rect 262 1959 268 1960
rect 262 1955 263 1959
rect 267 1955 268 1959
rect 262 1954 268 1955
rect 326 1959 332 1960
rect 326 1955 327 1959
rect 331 1955 332 1959
rect 326 1954 332 1955
rect 334 1959 340 1960
rect 334 1955 335 1959
rect 339 1955 340 1959
rect 334 1954 340 1955
rect 462 1959 468 1960
rect 462 1955 463 1959
rect 467 1955 468 1959
rect 462 1954 468 1955
rect 534 1959 540 1960
rect 534 1955 535 1959
rect 539 1955 540 1959
rect 534 1954 540 1955
rect 546 1959 552 1960
rect 546 1955 547 1959
rect 551 1955 552 1959
rect 546 1954 552 1955
rect 606 1959 612 1960
rect 606 1955 607 1959
rect 611 1955 612 1959
rect 606 1954 612 1955
rect 858 1959 864 1960
rect 858 1955 859 1959
rect 863 1955 864 1959
rect 858 1954 864 1955
rect 246 1948 252 1949
rect 246 1944 247 1948
rect 251 1944 252 1948
rect 246 1943 252 1944
rect 214 1939 220 1940
rect 214 1935 215 1939
rect 219 1935 220 1939
rect 214 1934 220 1935
rect 248 1931 250 1943
rect 264 1940 266 1954
rect 310 1948 316 1949
rect 310 1944 311 1948
rect 315 1944 316 1948
rect 310 1943 316 1944
rect 262 1939 268 1940
rect 262 1935 263 1939
rect 267 1935 268 1939
rect 262 1934 268 1935
rect 312 1931 314 1943
rect 328 1940 330 1954
rect 326 1939 332 1940
rect 326 1935 327 1939
rect 331 1935 332 1939
rect 326 1934 332 1935
rect 111 1930 115 1931
rect 111 1925 115 1926
rect 135 1930 139 1931
rect 135 1925 139 1926
rect 175 1930 179 1931
rect 175 1925 179 1926
rect 191 1930 195 1931
rect 191 1925 195 1926
rect 231 1930 235 1931
rect 231 1925 235 1926
rect 247 1930 251 1931
rect 247 1925 251 1926
rect 295 1930 299 1931
rect 295 1925 299 1926
rect 311 1930 315 1931
rect 311 1925 315 1926
rect 112 1905 114 1925
rect 136 1913 138 1925
rect 176 1913 178 1925
rect 190 1919 196 1920
rect 190 1915 191 1919
rect 195 1915 196 1919
rect 190 1914 196 1915
rect 134 1912 140 1913
rect 134 1908 135 1912
rect 139 1908 140 1912
rect 134 1907 140 1908
rect 174 1912 180 1913
rect 174 1908 175 1912
rect 179 1908 180 1912
rect 174 1907 180 1908
rect 110 1904 116 1905
rect 110 1900 111 1904
rect 115 1900 116 1904
rect 192 1900 194 1914
rect 232 1913 234 1925
rect 246 1919 252 1920
rect 246 1915 247 1919
rect 251 1915 252 1919
rect 246 1914 252 1915
rect 286 1919 292 1920
rect 286 1915 287 1919
rect 291 1915 292 1919
rect 286 1914 292 1915
rect 230 1912 236 1913
rect 230 1908 231 1912
rect 235 1908 236 1912
rect 230 1907 236 1908
rect 248 1900 250 1914
rect 288 1900 290 1914
rect 296 1913 298 1925
rect 336 1920 338 1954
rect 374 1948 380 1949
rect 374 1944 375 1948
rect 379 1944 380 1948
rect 374 1943 380 1944
rect 446 1948 452 1949
rect 446 1944 447 1948
rect 451 1944 452 1948
rect 446 1943 452 1944
rect 376 1931 378 1943
rect 394 1939 400 1940
rect 394 1935 395 1939
rect 399 1935 400 1939
rect 394 1934 400 1935
rect 367 1930 371 1931
rect 367 1925 371 1926
rect 375 1930 379 1931
rect 375 1925 379 1926
rect 334 1919 340 1920
rect 334 1915 335 1919
rect 339 1915 340 1919
rect 334 1914 340 1915
rect 368 1913 370 1925
rect 294 1912 300 1913
rect 294 1908 295 1912
rect 299 1908 300 1912
rect 294 1907 300 1908
rect 366 1912 372 1913
rect 366 1908 367 1912
rect 371 1908 372 1912
rect 366 1907 372 1908
rect 396 1900 398 1934
rect 448 1931 450 1943
rect 464 1940 466 1954
rect 518 1948 524 1949
rect 518 1944 519 1948
rect 523 1944 524 1948
rect 518 1943 524 1944
rect 462 1939 468 1940
rect 462 1935 463 1939
rect 467 1935 468 1939
rect 462 1934 468 1935
rect 520 1931 522 1943
rect 536 1940 538 1954
rect 590 1948 596 1949
rect 590 1944 591 1948
rect 595 1944 596 1948
rect 590 1943 596 1944
rect 534 1939 540 1940
rect 534 1935 535 1939
rect 539 1935 540 1939
rect 534 1934 540 1935
rect 592 1931 594 1943
rect 431 1930 435 1931
rect 431 1925 435 1926
rect 447 1930 451 1931
rect 447 1925 451 1926
rect 495 1930 499 1931
rect 495 1925 499 1926
rect 519 1930 523 1931
rect 519 1925 523 1926
rect 559 1930 563 1931
rect 559 1925 563 1926
rect 591 1930 595 1931
rect 608 1928 610 1954
rect 654 1948 660 1949
rect 654 1944 655 1948
rect 659 1944 660 1948
rect 654 1943 660 1944
rect 718 1948 724 1949
rect 718 1944 719 1948
rect 723 1944 724 1948
rect 718 1943 724 1944
rect 774 1948 780 1949
rect 774 1944 775 1948
rect 779 1944 780 1948
rect 774 1943 780 1944
rect 822 1948 828 1949
rect 822 1944 823 1948
rect 827 1944 828 1948
rect 822 1943 828 1944
rect 656 1931 658 1943
rect 720 1931 722 1943
rect 776 1931 778 1943
rect 824 1931 826 1943
rect 860 1940 862 1954
rect 870 1948 876 1949
rect 870 1944 871 1948
rect 875 1944 876 1948
rect 870 1943 876 1944
rect 858 1939 864 1940
rect 858 1935 859 1939
rect 863 1935 864 1939
rect 858 1934 864 1935
rect 872 1931 874 1943
rect 896 1940 898 1962
rect 1014 1959 1020 1960
rect 1014 1955 1015 1959
rect 1019 1955 1020 1959
rect 1014 1954 1020 1955
rect 1054 1959 1060 1960
rect 1054 1955 1055 1959
rect 1059 1955 1060 1959
rect 1134 1959 1140 1960
rect 1054 1954 1060 1955
rect 1094 1956 1100 1957
rect 918 1948 924 1949
rect 918 1944 919 1948
rect 923 1944 924 1948
rect 918 1943 924 1944
rect 966 1948 972 1949
rect 966 1944 967 1948
rect 971 1944 972 1948
rect 966 1943 972 1944
rect 1006 1948 1012 1949
rect 1006 1944 1007 1948
rect 1011 1944 1012 1948
rect 1006 1943 1012 1944
rect 894 1939 900 1940
rect 894 1935 895 1939
rect 899 1935 900 1939
rect 894 1934 900 1935
rect 920 1931 922 1943
rect 968 1931 970 1943
rect 1008 1931 1010 1943
rect 1016 1940 1018 1954
rect 1046 1948 1052 1949
rect 1046 1944 1047 1948
rect 1051 1944 1052 1948
rect 1046 1943 1052 1944
rect 1014 1939 1020 1940
rect 1014 1935 1015 1939
rect 1019 1935 1020 1939
rect 1014 1934 1020 1935
rect 1048 1931 1050 1943
rect 1056 1940 1058 1954
rect 1094 1952 1095 1956
rect 1099 1952 1100 1956
rect 1134 1955 1135 1959
rect 1139 1955 1140 1959
rect 1134 1954 1140 1955
rect 1302 1956 1308 1957
rect 1094 1951 1100 1952
rect 1054 1939 1060 1940
rect 1054 1935 1055 1939
rect 1059 1935 1060 1939
rect 1054 1934 1060 1935
rect 1096 1931 1098 1951
rect 1136 1947 1138 1954
rect 1302 1952 1303 1956
rect 1307 1952 1308 1956
rect 1302 1951 1308 1952
rect 1304 1947 1306 1951
rect 1135 1946 1139 1947
rect 1135 1941 1139 1942
rect 1159 1946 1163 1947
rect 1159 1941 1163 1942
rect 1223 1946 1227 1947
rect 1223 1941 1227 1942
rect 1303 1946 1307 1947
rect 1303 1941 1307 1942
rect 1136 1938 1138 1941
rect 1158 1940 1164 1941
rect 1134 1937 1140 1938
rect 1134 1933 1135 1937
rect 1139 1933 1140 1937
rect 1158 1936 1159 1940
rect 1163 1936 1164 1940
rect 1158 1935 1164 1936
rect 1222 1940 1228 1941
rect 1222 1936 1223 1940
rect 1227 1936 1228 1940
rect 1222 1935 1228 1936
rect 1302 1940 1308 1941
rect 1302 1936 1303 1940
rect 1307 1936 1308 1940
rect 1302 1935 1308 1936
rect 1134 1932 1140 1933
rect 615 1930 619 1931
rect 591 1925 595 1926
rect 606 1927 612 1928
rect 432 1913 434 1925
rect 438 1919 444 1920
rect 438 1915 439 1919
rect 443 1915 444 1919
rect 438 1914 444 1915
rect 430 1912 436 1913
rect 430 1908 431 1912
rect 435 1908 436 1912
rect 430 1907 436 1908
rect 440 1900 442 1914
rect 496 1913 498 1925
rect 502 1919 508 1920
rect 502 1915 503 1919
rect 507 1915 508 1919
rect 502 1914 508 1915
rect 510 1919 516 1920
rect 510 1915 511 1919
rect 515 1915 516 1919
rect 510 1914 516 1915
rect 494 1912 500 1913
rect 494 1908 495 1912
rect 499 1908 500 1912
rect 494 1907 500 1908
rect 504 1900 506 1914
rect 110 1899 116 1900
rect 158 1899 164 1900
rect 158 1895 159 1899
rect 163 1895 164 1899
rect 158 1894 164 1895
rect 190 1899 196 1900
rect 190 1895 191 1899
rect 195 1895 196 1899
rect 190 1894 196 1895
rect 246 1899 252 1900
rect 246 1895 247 1899
rect 251 1895 252 1899
rect 246 1894 252 1895
rect 286 1899 292 1900
rect 286 1895 287 1899
rect 291 1895 292 1899
rect 286 1894 292 1895
rect 394 1899 400 1900
rect 394 1895 395 1899
rect 399 1895 400 1899
rect 394 1894 400 1895
rect 438 1899 444 1900
rect 438 1895 439 1899
rect 443 1895 444 1899
rect 438 1894 444 1895
rect 502 1899 508 1900
rect 502 1895 503 1899
rect 507 1895 508 1899
rect 502 1894 508 1895
rect 110 1887 116 1888
rect 110 1883 111 1887
rect 115 1883 116 1887
rect 110 1882 116 1883
rect 134 1884 140 1885
rect 112 1875 114 1882
rect 134 1880 135 1884
rect 139 1880 140 1884
rect 134 1879 140 1880
rect 136 1875 138 1879
rect 111 1874 115 1875
rect 111 1869 115 1870
rect 135 1874 139 1875
rect 135 1869 139 1870
rect 112 1866 114 1869
rect 134 1868 140 1869
rect 110 1865 116 1866
rect 110 1861 111 1865
rect 115 1861 116 1865
rect 134 1864 135 1868
rect 139 1864 140 1868
rect 134 1863 140 1864
rect 110 1860 116 1861
rect 110 1848 116 1849
rect 110 1844 111 1848
rect 115 1844 116 1848
rect 110 1843 116 1844
rect 112 1815 114 1843
rect 134 1840 140 1841
rect 134 1836 135 1840
rect 139 1836 140 1840
rect 134 1835 140 1836
rect 136 1815 138 1835
rect 160 1832 162 1894
rect 174 1884 180 1885
rect 174 1880 175 1884
rect 179 1880 180 1884
rect 174 1879 180 1880
rect 230 1884 236 1885
rect 230 1880 231 1884
rect 235 1880 236 1884
rect 230 1879 236 1880
rect 294 1884 300 1885
rect 294 1880 295 1884
rect 299 1880 300 1884
rect 294 1879 300 1880
rect 366 1884 372 1885
rect 366 1880 367 1884
rect 371 1880 372 1884
rect 366 1879 372 1880
rect 430 1884 436 1885
rect 430 1880 431 1884
rect 435 1880 436 1884
rect 430 1879 436 1880
rect 494 1884 500 1885
rect 494 1880 495 1884
rect 499 1880 500 1884
rect 494 1879 500 1880
rect 176 1875 178 1879
rect 232 1875 234 1879
rect 296 1875 298 1879
rect 368 1875 370 1879
rect 432 1875 434 1879
rect 496 1875 498 1879
rect 175 1874 179 1875
rect 175 1869 179 1870
rect 199 1874 203 1875
rect 199 1869 203 1870
rect 231 1874 235 1875
rect 231 1869 235 1870
rect 271 1874 275 1875
rect 271 1869 275 1870
rect 295 1874 299 1875
rect 295 1869 299 1870
rect 335 1874 339 1875
rect 335 1869 339 1870
rect 367 1874 371 1875
rect 367 1869 371 1870
rect 399 1874 403 1875
rect 399 1869 403 1870
rect 431 1874 435 1875
rect 431 1869 435 1870
rect 455 1874 459 1875
rect 455 1869 459 1870
rect 495 1874 499 1875
rect 495 1869 499 1870
rect 503 1874 507 1875
rect 503 1869 507 1870
rect 198 1868 204 1869
rect 198 1864 199 1868
rect 203 1864 204 1868
rect 198 1863 204 1864
rect 270 1868 276 1869
rect 270 1864 271 1868
rect 275 1864 276 1868
rect 270 1863 276 1864
rect 334 1868 340 1869
rect 334 1864 335 1868
rect 339 1864 340 1868
rect 334 1863 340 1864
rect 398 1868 404 1869
rect 398 1864 399 1868
rect 403 1864 404 1868
rect 398 1863 404 1864
rect 454 1868 460 1869
rect 454 1864 455 1868
rect 459 1864 460 1868
rect 454 1863 460 1864
rect 502 1868 508 1869
rect 502 1864 503 1868
rect 507 1864 508 1868
rect 502 1863 508 1864
rect 294 1859 300 1860
rect 294 1855 295 1859
rect 299 1855 300 1859
rect 294 1854 300 1855
rect 478 1859 484 1860
rect 478 1855 479 1859
rect 483 1855 484 1859
rect 478 1854 484 1855
rect 206 1851 212 1852
rect 206 1847 207 1851
rect 211 1847 212 1851
rect 206 1846 212 1847
rect 234 1851 240 1852
rect 234 1847 235 1851
rect 239 1847 240 1851
rect 234 1846 240 1847
rect 198 1840 204 1841
rect 198 1836 199 1840
rect 203 1836 204 1840
rect 198 1835 204 1836
rect 158 1831 164 1832
rect 158 1827 159 1831
rect 163 1827 164 1831
rect 158 1826 164 1827
rect 200 1815 202 1835
rect 111 1814 115 1815
rect 111 1809 115 1810
rect 135 1814 139 1815
rect 135 1809 139 1810
rect 151 1814 155 1815
rect 151 1809 155 1810
rect 199 1814 203 1815
rect 199 1809 203 1810
rect 112 1789 114 1809
rect 152 1797 154 1809
rect 208 1804 210 1846
rect 236 1832 238 1846
rect 270 1840 276 1841
rect 270 1836 271 1840
rect 275 1836 276 1840
rect 270 1835 276 1836
rect 234 1831 240 1832
rect 234 1827 235 1831
rect 239 1827 240 1831
rect 234 1826 240 1827
rect 272 1815 274 1835
rect 296 1832 298 1854
rect 334 1840 340 1841
rect 334 1836 335 1840
rect 339 1836 340 1840
rect 334 1835 340 1836
rect 398 1840 404 1841
rect 398 1836 399 1840
rect 403 1836 404 1840
rect 398 1835 404 1836
rect 454 1840 460 1841
rect 454 1836 455 1840
rect 459 1836 460 1840
rect 454 1835 460 1836
rect 294 1831 300 1832
rect 294 1827 295 1831
rect 299 1827 300 1831
rect 294 1826 300 1827
rect 336 1815 338 1835
rect 400 1815 402 1835
rect 438 1831 444 1832
rect 438 1827 439 1831
rect 443 1827 444 1831
rect 438 1826 444 1827
rect 215 1814 219 1815
rect 215 1809 219 1810
rect 271 1814 275 1815
rect 271 1809 275 1810
rect 327 1814 331 1815
rect 327 1809 331 1810
rect 335 1814 339 1815
rect 335 1809 339 1810
rect 383 1814 387 1815
rect 383 1809 387 1810
rect 399 1814 403 1815
rect 399 1809 403 1810
rect 431 1814 435 1815
rect 431 1809 435 1810
rect 206 1803 212 1804
rect 206 1799 207 1803
rect 211 1799 212 1803
rect 206 1798 212 1799
rect 216 1797 218 1809
rect 222 1803 228 1804
rect 222 1799 223 1803
rect 227 1799 228 1803
rect 222 1798 228 1799
rect 150 1796 156 1797
rect 150 1792 151 1796
rect 155 1792 156 1796
rect 150 1791 156 1792
rect 214 1796 220 1797
rect 214 1792 215 1796
rect 219 1792 220 1796
rect 214 1791 220 1792
rect 110 1788 116 1789
rect 110 1784 111 1788
rect 115 1784 116 1788
rect 224 1784 226 1798
rect 272 1797 274 1809
rect 328 1797 330 1809
rect 374 1803 380 1804
rect 374 1799 375 1803
rect 379 1799 380 1803
rect 374 1798 380 1799
rect 270 1796 276 1797
rect 270 1792 271 1796
rect 275 1792 276 1796
rect 270 1791 276 1792
rect 326 1796 332 1797
rect 326 1792 327 1796
rect 331 1792 332 1796
rect 326 1791 332 1792
rect 110 1783 116 1784
rect 222 1783 228 1784
rect 222 1779 223 1783
rect 227 1779 228 1783
rect 222 1778 228 1779
rect 258 1783 264 1784
rect 258 1779 259 1783
rect 263 1779 264 1783
rect 258 1778 264 1779
rect 110 1771 116 1772
rect 110 1767 111 1771
rect 115 1767 116 1771
rect 110 1766 116 1767
rect 150 1768 156 1769
rect 112 1763 114 1766
rect 150 1764 151 1768
rect 155 1764 156 1768
rect 150 1763 156 1764
rect 214 1768 220 1769
rect 214 1764 215 1768
rect 219 1764 220 1768
rect 214 1763 220 1764
rect 111 1762 115 1763
rect 111 1757 115 1758
rect 151 1762 155 1763
rect 151 1757 155 1758
rect 215 1762 219 1763
rect 215 1757 219 1758
rect 231 1762 235 1763
rect 231 1757 235 1758
rect 112 1754 114 1757
rect 230 1756 236 1757
rect 110 1753 116 1754
rect 110 1749 111 1753
rect 115 1749 116 1753
rect 230 1752 231 1756
rect 235 1752 236 1756
rect 230 1751 236 1752
rect 110 1748 116 1749
rect 110 1736 116 1737
rect 110 1732 111 1736
rect 115 1732 116 1736
rect 110 1731 116 1732
rect 112 1707 114 1731
rect 230 1728 236 1729
rect 230 1724 231 1728
rect 235 1724 236 1728
rect 230 1723 236 1724
rect 232 1707 234 1723
rect 260 1720 262 1778
rect 270 1768 276 1769
rect 270 1764 271 1768
rect 275 1764 276 1768
rect 270 1763 276 1764
rect 326 1768 332 1769
rect 326 1764 327 1768
rect 331 1764 332 1768
rect 326 1763 332 1764
rect 271 1762 275 1763
rect 271 1757 275 1758
rect 295 1762 299 1763
rect 295 1757 299 1758
rect 327 1762 331 1763
rect 327 1757 331 1758
rect 351 1762 355 1763
rect 351 1757 355 1758
rect 294 1756 300 1757
rect 294 1752 295 1756
rect 299 1752 300 1756
rect 294 1751 300 1752
rect 350 1756 356 1757
rect 350 1752 351 1756
rect 355 1752 356 1756
rect 350 1751 356 1752
rect 376 1740 378 1798
rect 384 1797 386 1809
rect 390 1803 396 1804
rect 390 1799 391 1803
rect 395 1799 396 1803
rect 390 1798 396 1799
rect 382 1796 388 1797
rect 382 1792 383 1796
rect 387 1792 388 1796
rect 382 1791 388 1792
rect 392 1784 394 1798
rect 432 1797 434 1809
rect 430 1796 436 1797
rect 430 1792 431 1796
rect 435 1792 436 1796
rect 430 1791 436 1792
rect 440 1784 442 1826
rect 456 1815 458 1835
rect 480 1832 482 1854
rect 512 1852 514 1914
rect 560 1913 562 1925
rect 606 1923 607 1927
rect 611 1923 612 1927
rect 615 1925 619 1926
rect 655 1930 659 1931
rect 655 1925 659 1926
rect 671 1930 675 1931
rect 671 1925 675 1926
rect 719 1930 723 1931
rect 719 1925 723 1926
rect 727 1930 731 1931
rect 727 1925 731 1926
rect 775 1930 779 1931
rect 775 1925 779 1926
rect 783 1930 787 1931
rect 783 1925 787 1926
rect 823 1930 827 1931
rect 823 1925 827 1926
rect 847 1930 851 1931
rect 847 1925 851 1926
rect 871 1930 875 1931
rect 871 1925 875 1926
rect 919 1930 923 1931
rect 919 1925 923 1926
rect 967 1930 971 1931
rect 967 1925 971 1926
rect 1007 1930 1011 1931
rect 1007 1925 1011 1926
rect 1047 1930 1051 1931
rect 1047 1925 1051 1926
rect 1095 1930 1099 1931
rect 1095 1925 1099 1926
rect 606 1922 612 1923
rect 616 1913 618 1925
rect 630 1919 636 1920
rect 630 1915 631 1919
rect 635 1915 636 1919
rect 630 1914 636 1915
rect 558 1912 564 1913
rect 558 1908 559 1912
rect 563 1908 564 1912
rect 558 1907 564 1908
rect 614 1912 620 1913
rect 614 1908 615 1912
rect 619 1908 620 1912
rect 614 1907 620 1908
rect 632 1900 634 1914
rect 672 1913 674 1925
rect 686 1919 692 1920
rect 686 1915 687 1919
rect 691 1915 692 1919
rect 686 1914 692 1915
rect 670 1912 676 1913
rect 670 1908 671 1912
rect 675 1908 676 1912
rect 670 1907 676 1908
rect 688 1900 690 1914
rect 728 1913 730 1925
rect 742 1919 748 1920
rect 742 1915 743 1919
rect 747 1915 748 1919
rect 742 1914 748 1915
rect 726 1912 732 1913
rect 726 1908 727 1912
rect 731 1908 732 1912
rect 726 1907 732 1908
rect 744 1900 746 1914
rect 784 1913 786 1925
rect 798 1919 804 1920
rect 798 1915 799 1919
rect 803 1915 804 1919
rect 798 1914 804 1915
rect 782 1912 788 1913
rect 782 1908 783 1912
rect 787 1908 788 1912
rect 782 1907 788 1908
rect 800 1900 802 1914
rect 848 1913 850 1925
rect 854 1919 860 1920
rect 854 1915 855 1919
rect 859 1915 860 1919
rect 854 1914 860 1915
rect 846 1912 852 1913
rect 846 1908 847 1912
rect 851 1908 852 1912
rect 846 1907 852 1908
rect 856 1900 858 1914
rect 1096 1905 1098 1925
rect 1134 1920 1140 1921
rect 1134 1916 1135 1920
rect 1139 1916 1140 1920
rect 1134 1915 1140 1916
rect 1094 1904 1100 1905
rect 1094 1900 1095 1904
rect 1099 1900 1100 1904
rect 622 1899 628 1900
rect 622 1895 623 1899
rect 627 1895 628 1899
rect 622 1894 628 1895
rect 630 1899 636 1900
rect 630 1895 631 1899
rect 635 1895 636 1899
rect 630 1894 636 1895
rect 686 1899 692 1900
rect 686 1895 687 1899
rect 691 1895 692 1899
rect 686 1894 692 1895
rect 742 1899 748 1900
rect 742 1895 743 1899
rect 747 1895 748 1899
rect 742 1894 748 1895
rect 798 1899 804 1900
rect 798 1895 799 1899
rect 803 1895 804 1899
rect 798 1894 804 1895
rect 854 1899 860 1900
rect 1094 1899 1100 1900
rect 854 1895 855 1899
rect 859 1895 860 1899
rect 854 1894 860 1895
rect 558 1884 564 1885
rect 558 1880 559 1884
rect 563 1880 564 1884
rect 558 1879 564 1880
rect 614 1884 620 1885
rect 614 1880 615 1884
rect 619 1880 620 1884
rect 614 1879 620 1880
rect 560 1875 562 1879
rect 616 1875 618 1879
rect 551 1874 555 1875
rect 551 1869 555 1870
rect 559 1874 563 1875
rect 559 1869 563 1870
rect 599 1874 603 1875
rect 599 1869 603 1870
rect 615 1874 619 1875
rect 615 1869 619 1870
rect 550 1868 556 1869
rect 550 1864 551 1868
rect 555 1864 556 1868
rect 550 1863 556 1864
rect 598 1868 604 1869
rect 598 1864 599 1868
rect 603 1864 604 1868
rect 598 1863 604 1864
rect 510 1851 516 1852
rect 510 1847 511 1851
rect 515 1847 516 1851
rect 510 1846 516 1847
rect 518 1851 524 1852
rect 518 1847 519 1851
rect 523 1847 524 1851
rect 518 1846 524 1847
rect 502 1840 508 1841
rect 502 1836 503 1840
rect 507 1836 508 1840
rect 502 1835 508 1836
rect 478 1831 484 1832
rect 478 1827 479 1831
rect 483 1827 484 1831
rect 478 1826 484 1827
rect 504 1815 506 1835
rect 455 1814 459 1815
rect 455 1809 459 1810
rect 479 1814 483 1815
rect 479 1809 483 1810
rect 503 1814 507 1815
rect 520 1812 522 1846
rect 550 1840 556 1841
rect 550 1836 551 1840
rect 555 1836 556 1840
rect 550 1835 556 1836
rect 598 1840 604 1841
rect 598 1836 599 1840
rect 603 1836 604 1840
rect 598 1835 604 1836
rect 552 1815 554 1835
rect 600 1815 602 1835
rect 624 1824 626 1894
rect 1136 1891 1138 1915
rect 1158 1912 1164 1913
rect 1158 1908 1159 1912
rect 1163 1908 1164 1912
rect 1158 1907 1164 1908
rect 1222 1912 1228 1913
rect 1222 1908 1223 1912
rect 1227 1908 1228 1912
rect 1222 1907 1228 1908
rect 1302 1912 1308 1913
rect 1302 1908 1303 1912
rect 1307 1908 1308 1912
rect 1302 1907 1308 1908
rect 1160 1891 1162 1907
rect 1206 1903 1212 1904
rect 1206 1899 1207 1903
rect 1211 1899 1212 1903
rect 1206 1898 1212 1899
rect 1135 1890 1139 1891
rect 1094 1887 1100 1888
rect 670 1884 676 1885
rect 670 1880 671 1884
rect 675 1880 676 1884
rect 670 1879 676 1880
rect 726 1884 732 1885
rect 726 1880 727 1884
rect 731 1880 732 1884
rect 726 1879 732 1880
rect 782 1884 788 1885
rect 782 1880 783 1884
rect 787 1880 788 1884
rect 782 1879 788 1880
rect 846 1884 852 1885
rect 846 1880 847 1884
rect 851 1880 852 1884
rect 1094 1883 1095 1887
rect 1099 1883 1100 1887
rect 1135 1885 1139 1886
rect 1159 1890 1163 1891
rect 1159 1885 1163 1886
rect 1199 1890 1203 1891
rect 1199 1885 1203 1886
rect 1094 1882 1100 1883
rect 846 1879 852 1880
rect 672 1875 674 1879
rect 728 1875 730 1879
rect 784 1875 786 1879
rect 848 1875 850 1879
rect 1096 1875 1098 1882
rect 647 1874 651 1875
rect 647 1869 651 1870
rect 671 1874 675 1875
rect 671 1869 675 1870
rect 695 1874 699 1875
rect 695 1869 699 1870
rect 727 1874 731 1875
rect 727 1869 731 1870
rect 751 1874 755 1875
rect 751 1869 755 1870
rect 783 1874 787 1875
rect 783 1869 787 1870
rect 847 1874 851 1875
rect 847 1869 851 1870
rect 1095 1874 1099 1875
rect 1095 1869 1099 1870
rect 646 1868 652 1869
rect 646 1864 647 1868
rect 651 1864 652 1868
rect 646 1863 652 1864
rect 694 1868 700 1869
rect 694 1864 695 1868
rect 699 1864 700 1868
rect 694 1863 700 1864
rect 750 1868 756 1869
rect 750 1864 751 1868
rect 755 1864 756 1868
rect 1096 1866 1098 1869
rect 750 1863 756 1864
rect 1094 1865 1100 1866
rect 1136 1865 1138 1885
rect 1160 1873 1162 1885
rect 1200 1873 1202 1885
rect 1158 1872 1164 1873
rect 1158 1868 1159 1872
rect 1163 1868 1164 1872
rect 1158 1867 1164 1868
rect 1198 1872 1204 1873
rect 1198 1868 1199 1872
rect 1203 1868 1204 1872
rect 1198 1867 1204 1868
rect 1094 1861 1095 1865
rect 1099 1861 1100 1865
rect 1094 1860 1100 1861
rect 1134 1864 1140 1865
rect 1134 1860 1135 1864
rect 1139 1860 1140 1864
rect 1208 1860 1210 1898
rect 1224 1891 1226 1907
rect 1304 1891 1306 1907
rect 1328 1904 1330 1966
rect 1382 1956 1388 1957
rect 1382 1952 1383 1956
rect 1387 1952 1388 1956
rect 1382 1951 1388 1952
rect 1462 1956 1468 1957
rect 1462 1952 1463 1956
rect 1467 1952 1468 1956
rect 1462 1951 1468 1952
rect 1542 1956 1548 1957
rect 1542 1952 1543 1956
rect 1547 1952 1548 1956
rect 1542 1951 1548 1952
rect 1614 1956 1620 1957
rect 1614 1952 1615 1956
rect 1619 1952 1620 1956
rect 1614 1951 1620 1952
rect 1686 1956 1692 1957
rect 1686 1952 1687 1956
rect 1691 1952 1692 1956
rect 1686 1951 1692 1952
rect 1750 1956 1756 1957
rect 1750 1952 1751 1956
rect 1755 1952 1756 1956
rect 1750 1951 1756 1952
rect 1384 1947 1386 1951
rect 1464 1947 1466 1951
rect 1544 1947 1546 1951
rect 1616 1947 1618 1951
rect 1688 1947 1690 1951
rect 1752 1947 1754 1951
rect 1383 1946 1387 1947
rect 1383 1941 1387 1942
rect 1463 1946 1467 1947
rect 1463 1941 1467 1942
rect 1535 1946 1539 1947
rect 1535 1941 1539 1942
rect 1543 1946 1547 1947
rect 1543 1941 1547 1942
rect 1615 1946 1619 1947
rect 1615 1941 1619 1942
rect 1687 1946 1691 1947
rect 1687 1941 1691 1942
rect 1695 1946 1699 1947
rect 1695 1941 1699 1942
rect 1751 1946 1755 1947
rect 1751 1941 1755 1942
rect 1783 1946 1787 1947
rect 1783 1941 1787 1942
rect 1382 1940 1388 1941
rect 1382 1936 1383 1940
rect 1387 1936 1388 1940
rect 1382 1935 1388 1936
rect 1462 1940 1468 1941
rect 1462 1936 1463 1940
rect 1467 1936 1468 1940
rect 1462 1935 1468 1936
rect 1534 1940 1540 1941
rect 1534 1936 1535 1940
rect 1539 1936 1540 1940
rect 1534 1935 1540 1936
rect 1614 1940 1620 1941
rect 1614 1936 1615 1940
rect 1619 1936 1620 1940
rect 1614 1935 1620 1936
rect 1694 1940 1700 1941
rect 1694 1936 1695 1940
rect 1699 1936 1700 1940
rect 1694 1935 1700 1936
rect 1782 1940 1788 1941
rect 1782 1936 1783 1940
rect 1787 1936 1788 1940
rect 1782 1935 1788 1936
rect 1808 1924 1810 1986
rect 1816 1985 1818 1997
rect 1814 1984 1820 1985
rect 1814 1980 1815 1984
rect 1819 1980 1820 1984
rect 1814 1979 1820 1980
rect 1832 1972 1834 2006
rect 1840 2003 1842 2015
rect 1864 2012 1866 2034
rect 2032 2032 2034 2090
rect 2072 2089 2074 2101
rect 2070 2088 2076 2089
rect 2070 2084 2071 2088
rect 2075 2084 2076 2088
rect 2070 2083 2076 2084
rect 2120 2081 2122 2101
rect 2118 2080 2124 2081
rect 2118 2076 2119 2080
rect 2123 2076 2124 2080
rect 2094 2075 2100 2076
rect 2118 2075 2124 2076
rect 2094 2071 2095 2075
rect 2099 2071 2100 2075
rect 2094 2070 2100 2071
rect 2070 2060 2076 2061
rect 2070 2056 2071 2060
rect 2075 2056 2076 2060
rect 2070 2055 2076 2056
rect 2071 2054 2075 2055
rect 2071 2049 2075 2050
rect 2070 2048 2076 2049
rect 2070 2044 2071 2048
rect 2075 2044 2076 2048
rect 2070 2043 2076 2044
rect 1934 2031 1940 2032
rect 1934 2027 1935 2031
rect 1939 2027 1940 2031
rect 1934 2026 1940 2027
rect 2022 2031 2028 2032
rect 2022 2027 2023 2031
rect 2027 2027 2028 2031
rect 2022 2026 2028 2027
rect 2030 2031 2036 2032
rect 2030 2027 2031 2031
rect 2035 2027 2036 2031
rect 2030 2026 2036 2027
rect 1918 2020 1924 2021
rect 1918 2016 1919 2020
rect 1923 2016 1924 2020
rect 1918 2015 1924 2016
rect 1862 2011 1868 2012
rect 1862 2007 1863 2011
rect 1867 2007 1868 2011
rect 1862 2006 1868 2007
rect 1920 2003 1922 2015
rect 1936 2012 1938 2026
rect 2006 2020 2012 2021
rect 2006 2016 2007 2020
rect 2011 2016 2012 2020
rect 2006 2015 2012 2016
rect 1934 2011 1940 2012
rect 1934 2007 1935 2011
rect 1939 2007 1940 2011
rect 1934 2006 1940 2007
rect 2008 2003 2010 2015
rect 2024 2012 2026 2026
rect 2070 2020 2076 2021
rect 2070 2016 2071 2020
rect 2075 2016 2076 2020
rect 2070 2015 2076 2016
rect 2022 2011 2028 2012
rect 2022 2007 2023 2011
rect 2027 2007 2028 2011
rect 2022 2006 2028 2007
rect 2072 2003 2074 2015
rect 2096 2012 2098 2070
rect 2118 2063 2124 2064
rect 2118 2059 2119 2063
rect 2123 2059 2124 2063
rect 2118 2058 2124 2059
rect 2120 2055 2122 2058
rect 2119 2054 2123 2055
rect 2119 2049 2123 2050
rect 2120 2046 2122 2049
rect 2118 2045 2124 2046
rect 2118 2041 2119 2045
rect 2123 2041 2124 2045
rect 2118 2040 2124 2041
rect 2118 2028 2124 2029
rect 2118 2024 2119 2028
rect 2123 2024 2124 2028
rect 2118 2023 2124 2024
rect 2094 2011 2100 2012
rect 2094 2007 2095 2011
rect 2099 2007 2100 2011
rect 2094 2006 2100 2007
rect 2120 2003 2122 2023
rect 1839 2002 1843 2003
rect 1839 1997 1843 1998
rect 1879 2002 1883 2003
rect 1879 1997 1883 1998
rect 1919 2002 1923 2003
rect 1919 1997 1923 1998
rect 1951 2002 1955 2003
rect 1951 1997 1955 1998
rect 2007 2002 2011 2003
rect 2007 1997 2011 1998
rect 2023 2002 2027 2003
rect 2023 1997 2027 1998
rect 2071 2002 2075 2003
rect 2071 1997 2075 1998
rect 2119 2002 2123 2003
rect 2119 1997 2123 1998
rect 1880 1985 1882 1997
rect 1894 1991 1900 1992
rect 1894 1987 1895 1991
rect 1899 1987 1900 1991
rect 1894 1986 1900 1987
rect 1878 1984 1884 1985
rect 1878 1980 1879 1984
rect 1883 1980 1884 1984
rect 1878 1979 1884 1980
rect 1896 1972 1898 1986
rect 1952 1985 1954 1997
rect 1966 1991 1972 1992
rect 1966 1987 1967 1991
rect 1971 1987 1972 1991
rect 1966 1986 1972 1987
rect 1974 1991 1980 1992
rect 1974 1987 1975 1991
rect 1979 1987 1980 1991
rect 1974 1986 1980 1987
rect 1950 1984 1956 1985
rect 1950 1980 1951 1984
rect 1955 1980 1956 1984
rect 1950 1979 1956 1980
rect 1968 1972 1970 1986
rect 1976 1981 1978 1986
rect 2024 1985 2026 1997
rect 2072 1985 2074 1997
rect 2086 1991 2092 1992
rect 2086 1987 2087 1991
rect 2091 1987 2092 1991
rect 2086 1986 2092 1987
rect 2022 1984 2028 1985
rect 1975 1980 1979 1981
rect 2022 1980 2023 1984
rect 2027 1980 2028 1984
rect 2022 1979 2028 1980
rect 2070 1984 2076 1985
rect 2070 1980 2071 1984
rect 2075 1980 2076 1984
rect 2070 1979 2076 1980
rect 1975 1975 1979 1976
rect 2088 1972 2090 1986
rect 2120 1977 2122 1997
rect 2118 1976 2124 1977
rect 2118 1972 2119 1976
rect 2123 1972 2124 1976
rect 1830 1971 1836 1972
rect 1830 1967 1831 1971
rect 1835 1967 1836 1971
rect 1830 1966 1836 1967
rect 1894 1971 1900 1972
rect 1894 1967 1895 1971
rect 1899 1967 1900 1971
rect 1894 1966 1900 1967
rect 1966 1971 1972 1972
rect 1966 1967 1967 1971
rect 1971 1967 1972 1971
rect 1966 1966 1972 1967
rect 2078 1971 2084 1972
rect 2078 1967 2079 1971
rect 2083 1967 2084 1971
rect 2078 1966 2084 1967
rect 2086 1971 2092 1972
rect 2118 1971 2124 1972
rect 2086 1967 2087 1971
rect 2091 1967 2092 1971
rect 2086 1966 2092 1967
rect 1814 1956 1820 1957
rect 1814 1952 1815 1956
rect 1819 1952 1820 1956
rect 1814 1951 1820 1952
rect 1878 1956 1884 1957
rect 1878 1952 1879 1956
rect 1883 1952 1884 1956
rect 1878 1951 1884 1952
rect 1950 1956 1956 1957
rect 1950 1952 1951 1956
rect 1955 1952 1956 1956
rect 1950 1951 1956 1952
rect 2022 1956 2028 1957
rect 2022 1952 2023 1956
rect 2027 1952 2028 1956
rect 2022 1951 2028 1952
rect 2070 1956 2076 1957
rect 2070 1952 2071 1956
rect 2075 1952 2076 1956
rect 2070 1951 2076 1952
rect 1816 1947 1818 1951
rect 1880 1947 1882 1951
rect 1952 1947 1954 1951
rect 2024 1947 2026 1951
rect 2072 1947 2074 1951
rect 1815 1946 1819 1947
rect 1815 1941 1819 1942
rect 1879 1946 1883 1947
rect 1879 1941 1883 1942
rect 1951 1946 1955 1947
rect 1951 1941 1955 1942
rect 1983 1946 1987 1947
rect 1983 1941 1987 1942
rect 2023 1946 2027 1947
rect 2023 1941 2027 1942
rect 2071 1946 2075 1947
rect 2071 1941 2075 1942
rect 1878 1940 1884 1941
rect 1878 1936 1879 1940
rect 1883 1936 1884 1940
rect 1878 1935 1884 1936
rect 1982 1940 1988 1941
rect 1982 1936 1983 1940
rect 1987 1936 1988 1940
rect 1982 1935 1988 1936
rect 2070 1940 2076 1941
rect 2070 1936 2071 1940
rect 2075 1936 2076 1940
rect 2070 1935 2076 1936
rect 2006 1931 2012 1932
rect 2006 1927 2007 1931
rect 2011 1927 2012 1931
rect 2006 1926 2012 1927
rect 1398 1923 1404 1924
rect 1398 1919 1399 1923
rect 1403 1919 1404 1923
rect 1398 1918 1404 1919
rect 1446 1923 1452 1924
rect 1446 1919 1447 1923
rect 1451 1919 1452 1923
rect 1446 1918 1452 1919
rect 1474 1923 1480 1924
rect 1474 1919 1475 1923
rect 1479 1919 1480 1923
rect 1474 1918 1480 1919
rect 1806 1923 1812 1924
rect 1806 1919 1807 1923
rect 1811 1919 1812 1923
rect 1806 1918 1812 1919
rect 1382 1912 1388 1913
rect 1382 1908 1383 1912
rect 1387 1908 1388 1912
rect 1382 1907 1388 1908
rect 1326 1903 1332 1904
rect 1326 1899 1327 1903
rect 1331 1899 1332 1903
rect 1326 1898 1332 1899
rect 1384 1891 1386 1907
rect 1400 1904 1402 1918
rect 1448 1904 1450 1918
rect 1462 1912 1468 1913
rect 1462 1908 1463 1912
rect 1467 1908 1468 1912
rect 1462 1907 1468 1908
rect 1398 1903 1404 1904
rect 1398 1899 1399 1903
rect 1403 1899 1404 1903
rect 1398 1898 1404 1899
rect 1446 1903 1452 1904
rect 1446 1899 1447 1903
rect 1451 1899 1452 1903
rect 1446 1898 1452 1899
rect 1464 1891 1466 1907
rect 1223 1890 1227 1891
rect 1223 1885 1227 1886
rect 1263 1890 1267 1891
rect 1263 1885 1267 1886
rect 1303 1890 1307 1891
rect 1303 1885 1307 1886
rect 1327 1890 1331 1891
rect 1327 1885 1331 1886
rect 1383 1890 1387 1891
rect 1383 1885 1387 1886
rect 1391 1890 1395 1891
rect 1391 1885 1395 1886
rect 1447 1890 1451 1891
rect 1447 1885 1451 1886
rect 1463 1890 1467 1891
rect 1463 1885 1467 1886
rect 1214 1879 1220 1880
rect 1214 1875 1215 1879
rect 1219 1875 1220 1879
rect 1214 1874 1220 1875
rect 1216 1860 1218 1874
rect 1264 1873 1266 1885
rect 1278 1879 1284 1880
rect 1278 1875 1279 1879
rect 1283 1875 1284 1879
rect 1278 1874 1284 1875
rect 1318 1879 1324 1880
rect 1318 1875 1319 1879
rect 1323 1875 1324 1879
rect 1318 1874 1324 1875
rect 1262 1872 1268 1873
rect 1262 1868 1263 1872
rect 1267 1868 1268 1872
rect 1262 1867 1268 1868
rect 1280 1860 1282 1874
rect 1134 1859 1140 1860
rect 1206 1859 1212 1860
rect 1206 1855 1207 1859
rect 1211 1855 1212 1859
rect 1206 1854 1212 1855
rect 1214 1859 1220 1860
rect 1214 1855 1215 1859
rect 1219 1855 1220 1859
rect 1214 1854 1220 1855
rect 1278 1859 1284 1860
rect 1278 1855 1279 1859
rect 1283 1855 1284 1859
rect 1278 1854 1284 1855
rect 1094 1848 1100 1849
rect 1094 1844 1095 1848
rect 1099 1844 1100 1848
rect 1094 1843 1100 1844
rect 1134 1847 1140 1848
rect 1134 1843 1135 1847
rect 1139 1843 1140 1847
rect 646 1840 652 1841
rect 646 1836 647 1840
rect 651 1836 652 1840
rect 646 1835 652 1836
rect 694 1840 700 1841
rect 694 1836 695 1840
rect 699 1836 700 1840
rect 694 1835 700 1836
rect 750 1840 756 1841
rect 750 1836 751 1840
rect 755 1836 756 1840
rect 750 1835 756 1836
rect 622 1823 628 1824
rect 622 1819 623 1823
rect 627 1819 628 1823
rect 622 1818 628 1819
rect 648 1815 650 1835
rect 696 1815 698 1835
rect 752 1815 754 1835
rect 1096 1815 1098 1843
rect 1134 1842 1140 1843
rect 1158 1844 1164 1845
rect 1136 1839 1138 1842
rect 1158 1840 1159 1844
rect 1163 1840 1164 1844
rect 1158 1839 1164 1840
rect 1198 1844 1204 1845
rect 1198 1840 1199 1844
rect 1203 1840 1204 1844
rect 1198 1839 1204 1840
rect 1262 1844 1268 1845
rect 1262 1840 1263 1844
rect 1267 1840 1268 1844
rect 1262 1839 1268 1840
rect 1135 1838 1139 1839
rect 1135 1833 1139 1834
rect 1159 1838 1163 1839
rect 1159 1833 1163 1834
rect 1199 1838 1203 1839
rect 1199 1833 1203 1834
rect 1231 1838 1235 1839
rect 1231 1833 1235 1834
rect 1263 1838 1267 1839
rect 1263 1833 1267 1834
rect 1303 1838 1307 1839
rect 1303 1833 1307 1834
rect 1136 1830 1138 1833
rect 1158 1832 1164 1833
rect 1134 1829 1140 1830
rect 1134 1825 1135 1829
rect 1139 1825 1140 1829
rect 1158 1828 1159 1832
rect 1163 1828 1164 1832
rect 1158 1827 1164 1828
rect 1230 1832 1236 1833
rect 1230 1828 1231 1832
rect 1235 1828 1236 1832
rect 1230 1827 1236 1828
rect 1302 1832 1308 1833
rect 1302 1828 1303 1832
rect 1307 1828 1308 1832
rect 1302 1827 1308 1828
rect 1134 1824 1140 1825
rect 1320 1816 1322 1874
rect 1328 1873 1330 1885
rect 1392 1873 1394 1885
rect 1406 1879 1412 1880
rect 1406 1875 1407 1879
rect 1411 1875 1412 1879
rect 1406 1874 1412 1875
rect 1326 1872 1332 1873
rect 1326 1868 1327 1872
rect 1331 1868 1332 1872
rect 1326 1867 1332 1868
rect 1390 1872 1396 1873
rect 1390 1868 1391 1872
rect 1395 1868 1396 1872
rect 1390 1867 1396 1868
rect 1408 1860 1410 1874
rect 1448 1873 1450 1885
rect 1476 1880 1478 1918
rect 1534 1912 1540 1913
rect 1534 1908 1535 1912
rect 1539 1908 1540 1912
rect 1534 1907 1540 1908
rect 1614 1912 1620 1913
rect 1614 1908 1615 1912
rect 1619 1908 1620 1912
rect 1614 1907 1620 1908
rect 1694 1912 1700 1913
rect 1694 1908 1695 1912
rect 1699 1908 1700 1912
rect 1694 1907 1700 1908
rect 1782 1912 1788 1913
rect 1782 1908 1783 1912
rect 1787 1908 1788 1912
rect 1782 1907 1788 1908
rect 1878 1912 1884 1913
rect 1878 1908 1879 1912
rect 1883 1908 1884 1912
rect 1878 1907 1884 1908
rect 1982 1912 1988 1913
rect 1982 1908 1983 1912
rect 1987 1908 1988 1912
rect 1982 1907 1988 1908
rect 1536 1891 1538 1907
rect 1616 1891 1618 1907
rect 1696 1891 1698 1907
rect 1734 1903 1740 1904
rect 1734 1899 1735 1903
rect 1739 1899 1740 1903
rect 1734 1898 1740 1899
rect 1503 1890 1507 1891
rect 1503 1885 1507 1886
rect 1535 1890 1539 1891
rect 1535 1885 1539 1886
rect 1559 1890 1563 1891
rect 1559 1885 1563 1886
rect 1615 1890 1619 1891
rect 1615 1885 1619 1886
rect 1631 1890 1635 1891
rect 1631 1885 1635 1886
rect 1695 1890 1699 1891
rect 1695 1885 1699 1886
rect 1711 1890 1715 1891
rect 1711 1885 1715 1886
rect 1462 1879 1468 1880
rect 1462 1875 1463 1879
rect 1467 1875 1468 1879
rect 1462 1874 1468 1875
rect 1474 1879 1480 1880
rect 1474 1875 1475 1879
rect 1479 1875 1480 1879
rect 1474 1874 1480 1875
rect 1446 1872 1452 1873
rect 1446 1868 1447 1872
rect 1451 1868 1452 1872
rect 1446 1867 1452 1868
rect 1464 1860 1466 1874
rect 1504 1873 1506 1885
rect 1560 1873 1562 1885
rect 1574 1879 1580 1880
rect 1574 1875 1575 1879
rect 1579 1875 1580 1879
rect 1574 1874 1580 1875
rect 1502 1872 1508 1873
rect 1502 1868 1503 1872
rect 1507 1868 1508 1872
rect 1502 1867 1508 1868
rect 1558 1872 1564 1873
rect 1558 1868 1559 1872
rect 1563 1868 1564 1872
rect 1558 1867 1564 1868
rect 1576 1860 1578 1874
rect 1632 1873 1634 1885
rect 1646 1879 1652 1880
rect 1646 1875 1647 1879
rect 1651 1875 1652 1879
rect 1646 1874 1652 1875
rect 1670 1879 1676 1880
rect 1670 1875 1671 1879
rect 1675 1875 1676 1879
rect 1670 1874 1676 1875
rect 1630 1872 1636 1873
rect 1630 1868 1631 1872
rect 1635 1868 1636 1872
rect 1630 1867 1636 1868
rect 1648 1860 1650 1874
rect 1398 1859 1404 1860
rect 1398 1855 1399 1859
rect 1403 1855 1404 1859
rect 1398 1854 1404 1855
rect 1406 1859 1412 1860
rect 1406 1855 1407 1859
rect 1411 1855 1412 1859
rect 1406 1854 1412 1855
rect 1462 1859 1468 1860
rect 1462 1855 1463 1859
rect 1467 1855 1468 1859
rect 1462 1854 1468 1855
rect 1574 1859 1580 1860
rect 1574 1855 1575 1859
rect 1579 1855 1580 1859
rect 1574 1854 1580 1855
rect 1646 1859 1652 1860
rect 1646 1855 1647 1859
rect 1651 1855 1652 1859
rect 1646 1854 1652 1855
rect 1326 1844 1332 1845
rect 1326 1840 1327 1844
rect 1331 1840 1332 1844
rect 1326 1839 1332 1840
rect 1390 1844 1396 1845
rect 1390 1840 1391 1844
rect 1395 1840 1396 1844
rect 1390 1839 1396 1840
rect 1327 1838 1331 1839
rect 1327 1833 1331 1834
rect 1383 1838 1387 1839
rect 1383 1833 1387 1834
rect 1391 1838 1395 1839
rect 1391 1833 1395 1834
rect 1382 1832 1388 1833
rect 1382 1828 1383 1832
rect 1387 1828 1388 1832
rect 1382 1827 1388 1828
rect 1246 1815 1252 1816
rect 527 1814 531 1815
rect 503 1809 507 1810
rect 518 1811 524 1812
rect 480 1797 482 1809
rect 518 1807 519 1811
rect 523 1807 524 1811
rect 527 1809 531 1810
rect 551 1814 555 1815
rect 551 1809 555 1810
rect 575 1814 579 1815
rect 575 1809 579 1810
rect 599 1814 603 1815
rect 599 1809 603 1810
rect 623 1814 627 1815
rect 623 1809 627 1810
rect 647 1814 651 1815
rect 647 1809 651 1810
rect 671 1814 675 1815
rect 671 1809 675 1810
rect 695 1814 699 1815
rect 695 1809 699 1810
rect 727 1814 731 1815
rect 727 1809 731 1810
rect 751 1814 755 1815
rect 751 1809 755 1810
rect 1095 1814 1099 1815
rect 1095 1809 1099 1810
rect 1134 1812 1140 1813
rect 518 1806 524 1807
rect 528 1797 530 1809
rect 542 1803 548 1804
rect 542 1799 543 1803
rect 547 1799 548 1803
rect 542 1798 548 1799
rect 478 1796 484 1797
rect 478 1792 479 1796
rect 483 1792 484 1796
rect 478 1791 484 1792
rect 526 1796 532 1797
rect 526 1792 527 1796
rect 531 1792 532 1796
rect 526 1791 532 1792
rect 544 1784 546 1798
rect 576 1797 578 1809
rect 590 1803 596 1804
rect 590 1799 591 1803
rect 595 1799 596 1803
rect 590 1798 596 1799
rect 574 1796 580 1797
rect 574 1792 575 1796
rect 579 1792 580 1796
rect 574 1791 580 1792
rect 592 1784 594 1798
rect 624 1797 626 1809
rect 638 1803 644 1804
rect 638 1799 639 1803
rect 643 1799 644 1803
rect 638 1798 644 1799
rect 622 1796 628 1797
rect 622 1792 623 1796
rect 627 1792 628 1796
rect 622 1791 628 1792
rect 640 1784 642 1798
rect 672 1797 674 1809
rect 718 1803 724 1804
rect 718 1799 719 1803
rect 723 1799 724 1803
rect 718 1798 724 1799
rect 670 1796 676 1797
rect 670 1792 671 1796
rect 675 1792 676 1796
rect 670 1791 676 1792
rect 720 1784 722 1798
rect 728 1797 730 1809
rect 726 1796 732 1797
rect 726 1792 727 1796
rect 731 1792 732 1796
rect 726 1791 732 1792
rect 1096 1789 1098 1809
rect 1134 1808 1135 1812
rect 1139 1808 1140 1812
rect 1246 1811 1247 1815
rect 1251 1811 1252 1815
rect 1246 1810 1252 1811
rect 1310 1815 1316 1816
rect 1310 1811 1311 1815
rect 1315 1811 1316 1815
rect 1310 1810 1316 1811
rect 1318 1815 1324 1816
rect 1318 1811 1319 1815
rect 1323 1811 1324 1815
rect 1318 1810 1324 1811
rect 1134 1807 1140 1808
rect 1094 1788 1100 1789
rect 1094 1784 1095 1788
rect 1099 1784 1100 1788
rect 1136 1787 1138 1807
rect 1158 1804 1164 1805
rect 1158 1800 1159 1804
rect 1163 1800 1164 1804
rect 1158 1799 1164 1800
rect 1230 1804 1236 1805
rect 1230 1800 1231 1804
rect 1235 1800 1236 1804
rect 1230 1799 1236 1800
rect 1160 1787 1162 1799
rect 1214 1795 1220 1796
rect 1214 1791 1215 1795
rect 1219 1791 1220 1795
rect 1214 1790 1220 1791
rect 390 1783 396 1784
rect 390 1779 391 1783
rect 395 1779 396 1783
rect 390 1778 396 1779
rect 438 1783 444 1784
rect 438 1779 439 1783
rect 443 1779 444 1783
rect 438 1778 444 1779
rect 542 1783 548 1784
rect 542 1779 543 1783
rect 547 1779 548 1783
rect 542 1778 548 1779
rect 590 1783 596 1784
rect 590 1779 591 1783
rect 595 1779 596 1783
rect 590 1778 596 1779
rect 638 1783 644 1784
rect 638 1779 639 1783
rect 643 1779 644 1783
rect 638 1778 644 1779
rect 718 1783 724 1784
rect 718 1779 719 1783
rect 723 1779 724 1783
rect 718 1778 724 1779
rect 782 1783 788 1784
rect 1094 1783 1100 1784
rect 1135 1786 1139 1787
rect 782 1779 783 1783
rect 787 1779 788 1783
rect 1135 1781 1139 1782
rect 1159 1786 1163 1787
rect 1159 1781 1163 1782
rect 1191 1786 1195 1787
rect 1191 1781 1195 1782
rect 782 1778 788 1779
rect 382 1768 388 1769
rect 382 1764 383 1768
rect 387 1764 388 1768
rect 382 1763 388 1764
rect 430 1768 436 1769
rect 430 1764 431 1768
rect 435 1764 436 1768
rect 430 1763 436 1764
rect 478 1768 484 1769
rect 478 1764 479 1768
rect 483 1764 484 1768
rect 478 1763 484 1764
rect 526 1768 532 1769
rect 526 1764 527 1768
rect 531 1764 532 1768
rect 526 1763 532 1764
rect 574 1768 580 1769
rect 574 1764 575 1768
rect 579 1764 580 1768
rect 574 1763 580 1764
rect 622 1768 628 1769
rect 622 1764 623 1768
rect 627 1764 628 1768
rect 622 1763 628 1764
rect 670 1768 676 1769
rect 670 1764 671 1768
rect 675 1764 676 1768
rect 670 1763 676 1764
rect 726 1768 732 1769
rect 726 1764 727 1768
rect 731 1764 732 1768
rect 726 1763 732 1764
rect 383 1762 387 1763
rect 383 1757 387 1758
rect 415 1762 419 1763
rect 415 1757 419 1758
rect 431 1762 435 1763
rect 431 1757 435 1758
rect 479 1762 483 1763
rect 479 1757 483 1758
rect 527 1762 531 1763
rect 527 1757 531 1758
rect 543 1762 547 1763
rect 543 1757 547 1758
rect 575 1762 579 1763
rect 575 1757 579 1758
rect 615 1762 619 1763
rect 615 1757 619 1758
rect 623 1762 627 1763
rect 623 1757 627 1758
rect 671 1762 675 1763
rect 671 1757 675 1758
rect 687 1762 691 1763
rect 687 1757 691 1758
rect 727 1762 731 1763
rect 727 1757 731 1758
rect 759 1762 763 1763
rect 759 1757 763 1758
rect 414 1756 420 1757
rect 414 1752 415 1756
rect 419 1752 420 1756
rect 414 1751 420 1752
rect 478 1756 484 1757
rect 478 1752 479 1756
rect 483 1752 484 1756
rect 478 1751 484 1752
rect 542 1756 548 1757
rect 542 1752 543 1756
rect 547 1752 548 1756
rect 542 1751 548 1752
rect 614 1756 620 1757
rect 614 1752 615 1756
rect 619 1752 620 1756
rect 614 1751 620 1752
rect 686 1756 692 1757
rect 686 1752 687 1756
rect 691 1752 692 1756
rect 686 1751 692 1752
rect 758 1756 764 1757
rect 758 1752 759 1756
rect 763 1752 764 1756
rect 758 1751 764 1752
rect 286 1739 292 1740
rect 286 1735 287 1739
rect 291 1735 292 1739
rect 286 1734 292 1735
rect 306 1739 312 1740
rect 306 1735 307 1739
rect 311 1735 312 1739
rect 306 1734 312 1735
rect 374 1739 380 1740
rect 374 1735 375 1739
rect 379 1735 380 1739
rect 374 1734 380 1735
rect 462 1739 468 1740
rect 462 1735 463 1739
rect 467 1735 468 1739
rect 462 1734 468 1735
rect 662 1739 668 1740
rect 662 1735 663 1739
rect 667 1735 668 1739
rect 662 1734 668 1735
rect 674 1739 680 1740
rect 674 1735 675 1739
rect 679 1735 680 1739
rect 674 1734 680 1735
rect 288 1720 290 1734
rect 294 1728 300 1729
rect 294 1724 295 1728
rect 299 1724 300 1728
rect 294 1723 300 1724
rect 258 1719 264 1720
rect 258 1715 259 1719
rect 263 1715 264 1719
rect 258 1714 264 1715
rect 286 1719 292 1720
rect 286 1715 287 1719
rect 291 1715 292 1719
rect 286 1714 292 1715
rect 296 1707 298 1723
rect 111 1706 115 1707
rect 111 1701 115 1702
rect 135 1706 139 1707
rect 135 1701 139 1702
rect 199 1706 203 1707
rect 199 1701 203 1702
rect 231 1706 235 1707
rect 231 1701 235 1702
rect 279 1706 283 1707
rect 279 1701 283 1702
rect 295 1706 299 1707
rect 295 1701 299 1702
rect 112 1681 114 1701
rect 136 1689 138 1701
rect 200 1689 202 1701
rect 206 1695 212 1696
rect 206 1691 207 1695
rect 211 1691 212 1695
rect 206 1690 212 1691
rect 134 1688 140 1689
rect 134 1684 135 1688
rect 139 1684 140 1688
rect 134 1683 140 1684
rect 198 1688 204 1689
rect 198 1684 199 1688
rect 203 1684 204 1688
rect 198 1683 204 1684
rect 110 1680 116 1681
rect 110 1676 111 1680
rect 115 1676 116 1680
rect 208 1676 210 1690
rect 280 1689 282 1701
rect 308 1696 310 1734
rect 350 1728 356 1729
rect 350 1724 351 1728
rect 355 1724 356 1728
rect 350 1723 356 1724
rect 414 1728 420 1729
rect 414 1724 415 1728
rect 419 1724 420 1728
rect 414 1723 420 1724
rect 352 1707 354 1723
rect 416 1707 418 1723
rect 464 1720 466 1734
rect 478 1728 484 1729
rect 478 1724 479 1728
rect 483 1724 484 1728
rect 478 1723 484 1724
rect 542 1728 548 1729
rect 542 1724 543 1728
rect 547 1724 548 1728
rect 542 1723 548 1724
rect 614 1728 620 1729
rect 614 1724 615 1728
rect 619 1724 620 1728
rect 614 1723 620 1724
rect 462 1719 468 1720
rect 462 1715 463 1719
rect 467 1715 468 1719
rect 462 1714 468 1715
rect 480 1707 482 1723
rect 544 1707 546 1723
rect 570 1719 576 1720
rect 570 1715 571 1719
rect 575 1715 576 1719
rect 570 1714 576 1715
rect 351 1706 355 1707
rect 351 1701 355 1702
rect 367 1706 371 1707
rect 367 1701 371 1702
rect 415 1706 419 1707
rect 415 1701 419 1702
rect 463 1706 467 1707
rect 463 1701 467 1702
rect 479 1706 483 1707
rect 479 1701 483 1702
rect 543 1706 547 1707
rect 543 1701 547 1702
rect 551 1706 555 1707
rect 551 1701 555 1702
rect 294 1695 300 1696
rect 294 1691 295 1695
rect 299 1691 300 1695
rect 294 1690 300 1691
rect 306 1695 312 1696
rect 306 1691 307 1695
rect 311 1691 312 1695
rect 306 1690 312 1691
rect 314 1695 320 1696
rect 314 1691 315 1695
rect 319 1691 320 1695
rect 314 1690 320 1691
rect 278 1688 284 1689
rect 278 1684 279 1688
rect 283 1684 284 1688
rect 278 1683 284 1684
rect 296 1676 298 1690
rect 110 1675 116 1676
rect 190 1675 196 1676
rect 190 1671 191 1675
rect 195 1671 196 1675
rect 190 1670 196 1671
rect 206 1675 212 1676
rect 206 1671 207 1675
rect 211 1671 212 1675
rect 206 1670 212 1671
rect 294 1675 300 1676
rect 294 1671 295 1675
rect 299 1671 300 1675
rect 294 1670 300 1671
rect 110 1663 116 1664
rect 110 1659 111 1663
rect 115 1659 116 1663
rect 110 1658 116 1659
rect 134 1660 140 1661
rect 112 1651 114 1658
rect 134 1656 135 1660
rect 139 1656 140 1660
rect 134 1655 140 1656
rect 136 1651 138 1655
rect 111 1650 115 1651
rect 111 1645 115 1646
rect 135 1650 139 1651
rect 135 1645 139 1646
rect 183 1650 187 1651
rect 183 1645 187 1646
rect 112 1642 114 1645
rect 134 1644 140 1645
rect 110 1641 116 1642
rect 110 1637 111 1641
rect 115 1637 116 1641
rect 134 1640 135 1644
rect 139 1640 140 1644
rect 134 1639 140 1640
rect 182 1644 188 1645
rect 182 1640 183 1644
rect 187 1640 188 1644
rect 182 1639 188 1640
rect 110 1636 116 1637
rect 158 1627 164 1628
rect 110 1624 116 1625
rect 110 1620 111 1624
rect 115 1620 116 1624
rect 158 1623 159 1627
rect 163 1623 164 1627
rect 158 1622 164 1623
rect 170 1627 176 1628
rect 170 1623 171 1627
rect 175 1623 176 1627
rect 170 1622 176 1623
rect 110 1619 116 1620
rect 112 1599 114 1619
rect 134 1616 140 1617
rect 134 1612 135 1616
rect 139 1612 140 1616
rect 134 1611 140 1612
rect 136 1599 138 1611
rect 111 1598 115 1599
rect 111 1593 115 1594
rect 135 1598 139 1599
rect 135 1593 139 1594
rect 112 1573 114 1593
rect 136 1581 138 1593
rect 160 1588 162 1622
rect 172 1608 174 1622
rect 182 1616 188 1617
rect 182 1612 183 1616
rect 187 1612 188 1616
rect 182 1611 188 1612
rect 170 1607 176 1608
rect 170 1603 171 1607
rect 175 1603 176 1607
rect 170 1602 176 1603
rect 184 1599 186 1611
rect 192 1608 194 1670
rect 198 1660 204 1661
rect 198 1656 199 1660
rect 203 1656 204 1660
rect 198 1655 204 1656
rect 278 1660 284 1661
rect 278 1656 279 1660
rect 283 1656 284 1660
rect 278 1655 284 1656
rect 200 1651 202 1655
rect 280 1651 282 1655
rect 199 1650 203 1651
rect 199 1645 203 1646
rect 263 1650 267 1651
rect 263 1645 267 1646
rect 279 1650 283 1651
rect 279 1645 283 1646
rect 262 1644 268 1645
rect 262 1640 263 1644
rect 267 1640 268 1644
rect 262 1639 268 1640
rect 316 1636 318 1690
rect 368 1689 370 1701
rect 464 1689 466 1701
rect 552 1689 554 1701
rect 366 1688 372 1689
rect 366 1684 367 1688
rect 371 1684 372 1688
rect 366 1683 372 1684
rect 462 1688 468 1689
rect 462 1684 463 1688
rect 467 1684 468 1688
rect 462 1683 468 1684
rect 550 1688 556 1689
rect 550 1684 551 1688
rect 555 1684 556 1688
rect 550 1683 556 1684
rect 572 1676 574 1714
rect 616 1707 618 1723
rect 615 1706 619 1707
rect 615 1701 619 1702
rect 639 1706 643 1707
rect 639 1701 643 1702
rect 640 1689 642 1701
rect 664 1696 666 1734
rect 676 1720 678 1734
rect 686 1728 692 1729
rect 686 1724 687 1728
rect 691 1724 692 1728
rect 686 1723 692 1724
rect 758 1728 764 1729
rect 758 1724 759 1728
rect 763 1724 764 1728
rect 758 1723 764 1724
rect 674 1719 680 1720
rect 674 1715 675 1719
rect 679 1715 680 1719
rect 674 1714 680 1715
rect 688 1707 690 1723
rect 760 1707 762 1723
rect 784 1720 786 1778
rect 1094 1771 1100 1772
rect 1094 1767 1095 1771
rect 1099 1767 1100 1771
rect 1094 1766 1100 1767
rect 1096 1763 1098 1766
rect 831 1762 835 1763
rect 831 1757 835 1758
rect 911 1762 915 1763
rect 911 1757 915 1758
rect 991 1762 995 1763
rect 991 1757 995 1758
rect 1095 1762 1099 1763
rect 1136 1761 1138 1781
rect 1192 1769 1194 1781
rect 1190 1768 1196 1769
rect 1190 1764 1191 1768
rect 1195 1764 1196 1768
rect 1190 1763 1196 1764
rect 1095 1757 1099 1758
rect 1134 1760 1140 1761
rect 830 1756 836 1757
rect 830 1752 831 1756
rect 835 1752 836 1756
rect 830 1751 836 1752
rect 910 1756 916 1757
rect 910 1752 911 1756
rect 915 1752 916 1756
rect 910 1751 916 1752
rect 990 1756 996 1757
rect 990 1752 991 1756
rect 995 1752 996 1756
rect 1096 1754 1098 1757
rect 1134 1756 1135 1760
rect 1139 1756 1140 1760
rect 1216 1756 1218 1790
rect 1232 1787 1234 1799
rect 1248 1796 1250 1810
rect 1302 1804 1308 1805
rect 1302 1800 1303 1804
rect 1307 1800 1308 1804
rect 1302 1799 1308 1800
rect 1246 1795 1252 1796
rect 1246 1791 1247 1795
rect 1251 1791 1252 1795
rect 1246 1790 1252 1791
rect 1304 1787 1306 1799
rect 1312 1796 1314 1810
rect 1382 1804 1388 1805
rect 1382 1800 1383 1804
rect 1387 1800 1388 1804
rect 1382 1799 1388 1800
rect 1310 1795 1316 1796
rect 1310 1791 1311 1795
rect 1315 1791 1316 1795
rect 1310 1790 1316 1791
rect 1384 1787 1386 1799
rect 1400 1796 1402 1854
rect 1446 1844 1452 1845
rect 1446 1840 1447 1844
rect 1451 1840 1452 1844
rect 1446 1839 1452 1840
rect 1502 1844 1508 1845
rect 1502 1840 1503 1844
rect 1507 1840 1508 1844
rect 1502 1839 1508 1840
rect 1558 1844 1564 1845
rect 1558 1840 1559 1844
rect 1563 1840 1564 1844
rect 1558 1839 1564 1840
rect 1630 1844 1636 1845
rect 1630 1840 1631 1844
rect 1635 1840 1636 1844
rect 1630 1839 1636 1840
rect 1447 1838 1451 1839
rect 1447 1833 1451 1834
rect 1463 1838 1467 1839
rect 1463 1833 1467 1834
rect 1503 1838 1507 1839
rect 1503 1833 1507 1834
rect 1551 1838 1555 1839
rect 1551 1833 1555 1834
rect 1559 1838 1563 1839
rect 1559 1833 1563 1834
rect 1631 1838 1635 1839
rect 1631 1833 1635 1834
rect 1647 1838 1651 1839
rect 1647 1833 1651 1834
rect 1462 1832 1468 1833
rect 1462 1828 1463 1832
rect 1467 1828 1468 1832
rect 1462 1827 1468 1828
rect 1550 1832 1556 1833
rect 1550 1828 1551 1832
rect 1555 1828 1556 1832
rect 1550 1827 1556 1828
rect 1646 1832 1652 1833
rect 1646 1828 1647 1832
rect 1651 1828 1652 1832
rect 1646 1827 1652 1828
rect 1672 1816 1674 1874
rect 1712 1873 1714 1885
rect 1710 1872 1716 1873
rect 1710 1868 1711 1872
rect 1715 1868 1716 1872
rect 1710 1867 1716 1868
rect 1736 1860 1738 1898
rect 1784 1891 1786 1907
rect 1880 1891 1882 1907
rect 1984 1891 1986 1907
rect 2008 1904 2010 1926
rect 2070 1912 2076 1913
rect 2070 1908 2071 1912
rect 2075 1908 2076 1912
rect 2070 1907 2076 1908
rect 2006 1903 2012 1904
rect 2006 1899 2007 1903
rect 2011 1899 2012 1903
rect 2006 1898 2012 1899
rect 2072 1891 2074 1907
rect 2080 1904 2082 1966
rect 2118 1959 2124 1960
rect 2118 1955 2119 1959
rect 2123 1955 2124 1959
rect 2118 1954 2124 1955
rect 2120 1947 2122 1954
rect 2119 1946 2123 1947
rect 2119 1941 2123 1942
rect 2120 1938 2122 1941
rect 2118 1937 2124 1938
rect 2118 1933 2119 1937
rect 2123 1933 2124 1937
rect 2118 1932 2124 1933
rect 2094 1923 2100 1924
rect 2094 1919 2095 1923
rect 2099 1919 2100 1923
rect 2094 1918 2100 1919
rect 2118 1920 2124 1921
rect 2078 1903 2084 1904
rect 2078 1899 2079 1903
rect 2083 1899 2084 1903
rect 2078 1898 2084 1899
rect 1783 1890 1787 1891
rect 1783 1885 1787 1886
rect 1799 1890 1803 1891
rect 1799 1885 1803 1886
rect 1879 1890 1883 1891
rect 1879 1885 1883 1886
rect 1895 1890 1899 1891
rect 1895 1885 1899 1886
rect 1983 1890 1987 1891
rect 1983 1885 1987 1886
rect 1991 1890 1995 1891
rect 1991 1885 1995 1886
rect 2071 1890 2075 1891
rect 2071 1885 2075 1886
rect 1800 1873 1802 1885
rect 1814 1879 1820 1880
rect 1814 1875 1815 1879
rect 1819 1875 1820 1879
rect 1814 1874 1820 1875
rect 1798 1872 1804 1873
rect 1798 1868 1799 1872
rect 1803 1868 1804 1872
rect 1798 1867 1804 1868
rect 1816 1860 1818 1874
rect 1896 1873 1898 1885
rect 1910 1879 1916 1880
rect 1910 1875 1911 1879
rect 1915 1875 1916 1879
rect 1910 1874 1916 1875
rect 1894 1872 1900 1873
rect 1894 1868 1895 1872
rect 1899 1868 1900 1872
rect 1894 1867 1900 1868
rect 1912 1860 1914 1874
rect 1992 1873 1994 1885
rect 2072 1873 2074 1885
rect 2096 1880 2098 1918
rect 2118 1916 2119 1920
rect 2123 1916 2124 1920
rect 2118 1915 2124 1916
rect 2120 1891 2122 1915
rect 2119 1890 2123 1891
rect 2119 1885 2123 1886
rect 2086 1879 2092 1880
rect 2086 1875 2087 1879
rect 2091 1875 2092 1879
rect 2086 1874 2092 1875
rect 2094 1879 2100 1880
rect 2094 1875 2095 1879
rect 2099 1875 2100 1879
rect 2094 1874 2100 1875
rect 1990 1872 1996 1873
rect 1990 1868 1991 1872
rect 1995 1868 1996 1872
rect 1990 1867 1996 1868
rect 2070 1872 2076 1873
rect 2070 1868 2071 1872
rect 2075 1868 2076 1872
rect 2070 1867 2076 1868
rect 2088 1860 2090 1874
rect 2120 1865 2122 1885
rect 2118 1864 2124 1865
rect 2118 1860 2119 1864
rect 2123 1860 2124 1864
rect 1734 1859 1740 1860
rect 1734 1855 1735 1859
rect 1739 1855 1740 1859
rect 1734 1854 1740 1855
rect 1814 1859 1820 1860
rect 1814 1855 1815 1859
rect 1819 1855 1820 1859
rect 1814 1854 1820 1855
rect 1910 1859 1916 1860
rect 1910 1855 1911 1859
rect 1915 1855 1916 1859
rect 1910 1854 1916 1855
rect 2078 1859 2084 1860
rect 2078 1855 2079 1859
rect 2083 1855 2084 1859
rect 2078 1854 2084 1855
rect 2086 1859 2092 1860
rect 2118 1859 2124 1860
rect 2086 1855 2087 1859
rect 2091 1855 2092 1859
rect 2086 1854 2092 1855
rect 1710 1844 1716 1845
rect 1710 1840 1711 1844
rect 1715 1840 1716 1844
rect 1710 1839 1716 1840
rect 1798 1844 1804 1845
rect 1798 1840 1799 1844
rect 1803 1840 1804 1844
rect 1798 1839 1804 1840
rect 1894 1844 1900 1845
rect 1894 1840 1895 1844
rect 1899 1840 1900 1844
rect 1894 1839 1900 1840
rect 1990 1844 1996 1845
rect 1990 1840 1991 1844
rect 1995 1840 1996 1844
rect 1990 1839 1996 1840
rect 2070 1844 2076 1845
rect 2070 1840 2071 1844
rect 2075 1840 2076 1844
rect 2070 1839 2076 1840
rect 1711 1838 1715 1839
rect 1711 1833 1715 1834
rect 1751 1838 1755 1839
rect 1751 1833 1755 1834
rect 1799 1838 1803 1839
rect 1799 1833 1803 1834
rect 1855 1838 1859 1839
rect 1855 1833 1859 1834
rect 1895 1838 1899 1839
rect 1895 1833 1899 1834
rect 1967 1838 1971 1839
rect 1967 1833 1971 1834
rect 1991 1838 1995 1839
rect 1991 1833 1995 1834
rect 2071 1838 2075 1839
rect 2071 1833 2075 1834
rect 1750 1832 1756 1833
rect 1750 1828 1751 1832
rect 1755 1828 1756 1832
rect 1750 1827 1756 1828
rect 1854 1832 1860 1833
rect 1854 1828 1855 1832
rect 1859 1828 1860 1832
rect 1854 1827 1860 1828
rect 1966 1832 1972 1833
rect 1966 1828 1967 1832
rect 1971 1828 1972 1832
rect 1966 1827 1972 1828
rect 2070 1832 2076 1833
rect 2070 1828 2071 1832
rect 2075 1828 2076 1832
rect 2070 1827 2076 1828
rect 1478 1815 1484 1816
rect 1478 1811 1479 1815
rect 1483 1811 1484 1815
rect 1478 1810 1484 1811
rect 1558 1815 1564 1816
rect 1558 1811 1559 1815
rect 1563 1811 1564 1815
rect 1558 1810 1564 1811
rect 1566 1815 1572 1816
rect 1566 1811 1567 1815
rect 1571 1811 1572 1815
rect 1566 1810 1572 1811
rect 1670 1815 1676 1816
rect 1670 1811 1671 1815
rect 1675 1811 1676 1815
rect 1670 1810 1676 1811
rect 1950 1815 1956 1816
rect 1950 1811 1951 1815
rect 1955 1811 1956 1815
rect 1950 1810 1956 1811
rect 1958 1815 1964 1816
rect 1958 1811 1959 1815
rect 1963 1811 1964 1815
rect 1958 1810 1964 1811
rect 1462 1804 1468 1805
rect 1462 1800 1463 1804
rect 1467 1800 1468 1804
rect 1462 1799 1468 1800
rect 1398 1795 1404 1796
rect 1398 1791 1399 1795
rect 1403 1791 1404 1795
rect 1398 1790 1404 1791
rect 1464 1787 1466 1799
rect 1480 1796 1482 1810
rect 1550 1804 1556 1805
rect 1550 1800 1551 1804
rect 1555 1800 1556 1804
rect 1550 1799 1556 1800
rect 1478 1795 1484 1796
rect 1478 1791 1479 1795
rect 1483 1791 1484 1795
rect 1478 1790 1484 1791
rect 1552 1787 1554 1799
rect 1560 1796 1562 1810
rect 1558 1795 1564 1796
rect 1558 1791 1559 1795
rect 1563 1791 1564 1795
rect 1558 1790 1564 1791
rect 1231 1786 1235 1787
rect 1231 1781 1235 1782
rect 1255 1786 1259 1787
rect 1255 1781 1259 1782
rect 1303 1786 1307 1787
rect 1303 1781 1307 1782
rect 1319 1786 1323 1787
rect 1319 1781 1323 1782
rect 1383 1786 1387 1787
rect 1383 1781 1387 1782
rect 1455 1786 1459 1787
rect 1455 1781 1459 1782
rect 1463 1786 1467 1787
rect 1463 1781 1467 1782
rect 1527 1786 1531 1787
rect 1527 1781 1531 1782
rect 1551 1786 1555 1787
rect 1551 1781 1555 1782
rect 1256 1769 1258 1781
rect 1270 1775 1276 1776
rect 1270 1771 1271 1775
rect 1275 1771 1276 1775
rect 1270 1770 1276 1771
rect 1254 1768 1260 1769
rect 1254 1764 1255 1768
rect 1259 1764 1260 1768
rect 1254 1763 1260 1764
rect 1272 1756 1274 1770
rect 1320 1769 1322 1781
rect 1334 1775 1340 1776
rect 1334 1771 1335 1775
rect 1339 1771 1340 1775
rect 1334 1770 1340 1771
rect 1366 1775 1372 1776
rect 1366 1771 1367 1775
rect 1371 1771 1372 1775
rect 1366 1770 1372 1771
rect 1318 1768 1324 1769
rect 1318 1764 1319 1768
rect 1323 1764 1324 1768
rect 1318 1763 1324 1764
rect 1336 1756 1338 1770
rect 1134 1755 1140 1756
rect 1214 1755 1220 1756
rect 990 1751 996 1752
rect 1094 1753 1100 1754
rect 1094 1749 1095 1753
rect 1099 1749 1100 1753
rect 1214 1751 1215 1755
rect 1219 1751 1220 1755
rect 1214 1750 1220 1751
rect 1270 1755 1276 1756
rect 1270 1751 1271 1755
rect 1275 1751 1276 1755
rect 1270 1750 1276 1751
rect 1334 1755 1340 1756
rect 1334 1751 1335 1755
rect 1339 1751 1340 1755
rect 1334 1750 1340 1751
rect 1094 1748 1100 1749
rect 1134 1743 1140 1744
rect 926 1739 932 1740
rect 926 1735 927 1739
rect 931 1735 932 1739
rect 926 1734 932 1735
rect 1002 1739 1008 1740
rect 1002 1735 1003 1739
rect 1007 1735 1008 1739
rect 1002 1734 1008 1735
rect 1010 1739 1016 1740
rect 1010 1735 1011 1739
rect 1015 1735 1016 1739
rect 1134 1739 1135 1743
rect 1139 1739 1140 1743
rect 1134 1738 1140 1739
rect 1190 1740 1196 1741
rect 1010 1734 1016 1735
rect 1094 1736 1100 1737
rect 830 1728 836 1729
rect 830 1724 831 1728
rect 835 1724 836 1728
rect 830 1723 836 1724
rect 910 1728 916 1729
rect 910 1724 911 1728
rect 915 1724 916 1728
rect 910 1723 916 1724
rect 782 1719 788 1720
rect 782 1715 783 1719
rect 787 1715 788 1719
rect 782 1714 788 1715
rect 798 1719 804 1720
rect 798 1715 799 1719
rect 803 1715 804 1719
rect 798 1714 804 1715
rect 687 1706 691 1707
rect 687 1701 691 1702
rect 719 1706 723 1707
rect 719 1701 723 1702
rect 759 1706 763 1707
rect 759 1701 763 1702
rect 791 1706 795 1707
rect 791 1701 795 1702
rect 662 1695 668 1696
rect 662 1691 663 1695
rect 667 1691 668 1695
rect 662 1690 668 1691
rect 720 1689 722 1701
rect 792 1689 794 1701
rect 638 1688 644 1689
rect 638 1684 639 1688
rect 643 1684 644 1688
rect 638 1683 644 1684
rect 718 1688 724 1689
rect 718 1684 719 1688
rect 723 1684 724 1688
rect 718 1683 724 1684
rect 790 1688 796 1689
rect 790 1684 791 1688
rect 795 1684 796 1688
rect 790 1683 796 1684
rect 800 1676 802 1714
rect 832 1707 834 1723
rect 912 1707 914 1723
rect 928 1720 930 1734
rect 990 1728 996 1729
rect 990 1724 991 1728
rect 995 1724 996 1728
rect 990 1723 996 1724
rect 926 1719 932 1720
rect 926 1715 927 1719
rect 931 1715 932 1719
rect 926 1714 932 1715
rect 992 1707 994 1723
rect 1004 1720 1006 1734
rect 1002 1719 1008 1720
rect 1002 1715 1003 1719
rect 1007 1715 1008 1719
rect 1002 1714 1008 1715
rect 831 1706 835 1707
rect 831 1701 835 1702
rect 855 1706 859 1707
rect 855 1701 859 1702
rect 911 1706 915 1707
rect 911 1701 915 1702
rect 919 1706 923 1707
rect 919 1701 923 1702
rect 983 1706 987 1707
rect 983 1701 987 1702
rect 991 1706 995 1707
rect 991 1701 995 1702
rect 806 1695 812 1696
rect 806 1691 807 1695
rect 811 1691 812 1695
rect 806 1690 812 1691
rect 808 1676 810 1690
rect 856 1689 858 1701
rect 862 1695 868 1696
rect 862 1691 863 1695
rect 867 1691 868 1695
rect 862 1690 868 1691
rect 870 1695 876 1696
rect 870 1691 871 1695
rect 875 1691 876 1695
rect 870 1690 876 1691
rect 854 1688 860 1689
rect 854 1684 855 1688
rect 859 1684 860 1688
rect 854 1683 860 1684
rect 864 1676 866 1690
rect 570 1675 576 1676
rect 570 1671 571 1675
rect 575 1671 576 1675
rect 570 1670 576 1671
rect 610 1675 616 1676
rect 610 1671 611 1675
rect 615 1671 616 1675
rect 610 1670 616 1671
rect 798 1675 804 1676
rect 798 1671 799 1675
rect 803 1671 804 1675
rect 798 1670 804 1671
rect 806 1675 812 1676
rect 806 1671 807 1675
rect 811 1671 812 1675
rect 806 1670 812 1671
rect 862 1675 868 1676
rect 862 1671 863 1675
rect 867 1671 868 1675
rect 862 1670 868 1671
rect 366 1660 372 1661
rect 366 1656 367 1660
rect 371 1656 372 1660
rect 366 1655 372 1656
rect 462 1660 468 1661
rect 462 1656 463 1660
rect 467 1656 468 1660
rect 462 1655 468 1656
rect 550 1660 556 1661
rect 550 1656 551 1660
rect 555 1656 556 1660
rect 550 1655 556 1656
rect 368 1651 370 1655
rect 464 1651 466 1655
rect 552 1651 554 1655
rect 343 1650 347 1651
rect 343 1645 347 1646
rect 367 1650 371 1651
rect 367 1645 371 1646
rect 423 1650 427 1651
rect 423 1645 427 1646
rect 463 1650 467 1651
rect 463 1645 467 1646
rect 503 1650 507 1651
rect 503 1645 507 1646
rect 551 1650 555 1651
rect 551 1645 555 1646
rect 583 1650 587 1651
rect 583 1645 587 1646
rect 342 1644 348 1645
rect 342 1640 343 1644
rect 347 1640 348 1644
rect 342 1639 348 1640
rect 422 1644 428 1645
rect 422 1640 423 1644
rect 427 1640 428 1644
rect 422 1639 428 1640
rect 502 1644 508 1645
rect 502 1640 503 1644
rect 507 1640 508 1644
rect 502 1639 508 1640
rect 582 1644 588 1645
rect 582 1640 583 1644
rect 587 1640 588 1644
rect 582 1639 588 1640
rect 314 1635 320 1636
rect 314 1631 315 1635
rect 319 1631 320 1635
rect 314 1630 320 1631
rect 262 1616 268 1617
rect 262 1612 263 1616
rect 267 1612 268 1616
rect 262 1611 268 1612
rect 342 1616 348 1617
rect 342 1612 343 1616
rect 347 1612 348 1616
rect 342 1611 348 1612
rect 422 1616 428 1617
rect 422 1612 423 1616
rect 427 1612 428 1616
rect 422 1611 428 1612
rect 502 1616 508 1617
rect 502 1612 503 1616
rect 507 1612 508 1616
rect 502 1611 508 1612
rect 582 1616 588 1617
rect 582 1612 583 1616
rect 587 1612 588 1616
rect 582 1611 588 1612
rect 190 1607 196 1608
rect 190 1603 191 1607
rect 195 1603 196 1607
rect 190 1602 196 1603
rect 264 1599 266 1611
rect 344 1599 346 1611
rect 424 1599 426 1611
rect 482 1607 488 1608
rect 482 1603 483 1607
rect 487 1603 488 1607
rect 482 1602 488 1603
rect 175 1598 179 1599
rect 175 1593 179 1594
rect 183 1598 187 1599
rect 183 1593 187 1594
rect 231 1598 235 1599
rect 231 1593 235 1594
rect 263 1598 267 1599
rect 263 1593 267 1594
rect 303 1598 307 1599
rect 303 1593 307 1594
rect 343 1598 347 1599
rect 343 1593 347 1594
rect 375 1598 379 1599
rect 375 1593 379 1594
rect 423 1598 427 1599
rect 423 1593 427 1594
rect 455 1598 459 1599
rect 455 1593 459 1594
rect 158 1587 164 1588
rect 158 1583 159 1587
rect 163 1583 164 1587
rect 158 1582 164 1583
rect 176 1581 178 1593
rect 182 1587 188 1588
rect 182 1583 183 1587
rect 187 1583 188 1587
rect 182 1582 188 1583
rect 134 1580 140 1581
rect 134 1576 135 1580
rect 139 1576 140 1580
rect 134 1575 140 1576
rect 174 1580 180 1581
rect 174 1576 175 1580
rect 179 1576 180 1580
rect 174 1575 180 1576
rect 110 1572 116 1573
rect 110 1568 111 1572
rect 115 1568 116 1572
rect 184 1568 186 1582
rect 232 1581 234 1593
rect 304 1581 306 1593
rect 376 1581 378 1593
rect 456 1581 458 1593
rect 230 1580 236 1581
rect 230 1576 231 1580
rect 235 1576 236 1580
rect 230 1575 236 1576
rect 302 1580 308 1581
rect 302 1576 303 1580
rect 307 1576 308 1580
rect 302 1575 308 1576
rect 374 1580 380 1581
rect 374 1576 375 1580
rect 379 1576 380 1580
rect 374 1575 380 1576
rect 454 1580 460 1581
rect 454 1576 455 1580
rect 459 1576 460 1580
rect 454 1575 460 1576
rect 484 1568 486 1602
rect 504 1599 506 1611
rect 584 1599 586 1611
rect 612 1608 614 1670
rect 638 1660 644 1661
rect 638 1656 639 1660
rect 643 1656 644 1660
rect 638 1655 644 1656
rect 718 1660 724 1661
rect 718 1656 719 1660
rect 723 1656 724 1660
rect 718 1655 724 1656
rect 790 1660 796 1661
rect 790 1656 791 1660
rect 795 1656 796 1660
rect 790 1655 796 1656
rect 854 1660 860 1661
rect 854 1656 855 1660
rect 859 1656 860 1660
rect 854 1655 860 1656
rect 640 1651 642 1655
rect 720 1651 722 1655
rect 792 1651 794 1655
rect 856 1651 858 1655
rect 639 1650 643 1651
rect 639 1645 643 1646
rect 655 1650 659 1651
rect 655 1645 659 1646
rect 719 1650 723 1651
rect 719 1645 723 1646
rect 727 1650 731 1651
rect 727 1645 731 1646
rect 791 1650 795 1651
rect 791 1645 795 1646
rect 847 1650 851 1651
rect 847 1645 851 1646
rect 855 1650 859 1651
rect 855 1645 859 1646
rect 654 1644 660 1645
rect 654 1640 655 1644
rect 659 1640 660 1644
rect 654 1639 660 1640
rect 726 1644 732 1645
rect 726 1640 727 1644
rect 731 1640 732 1644
rect 726 1639 732 1640
rect 790 1644 796 1645
rect 790 1640 791 1644
rect 795 1640 796 1644
rect 790 1639 796 1640
rect 846 1644 852 1645
rect 846 1640 847 1644
rect 851 1640 852 1644
rect 846 1639 852 1640
rect 872 1628 874 1690
rect 920 1689 922 1701
rect 984 1689 986 1701
rect 1012 1696 1014 1734
rect 1094 1732 1095 1736
rect 1099 1732 1100 1736
rect 1136 1735 1138 1738
rect 1190 1736 1191 1740
rect 1195 1736 1196 1740
rect 1190 1735 1196 1736
rect 1254 1740 1260 1741
rect 1254 1736 1255 1740
rect 1259 1736 1260 1740
rect 1254 1735 1260 1736
rect 1318 1740 1324 1741
rect 1318 1736 1319 1740
rect 1323 1736 1324 1740
rect 1318 1735 1324 1736
rect 1094 1731 1100 1732
rect 1135 1734 1139 1735
rect 1096 1707 1098 1731
rect 1135 1729 1139 1730
rect 1191 1734 1195 1735
rect 1191 1729 1195 1730
rect 1247 1734 1251 1735
rect 1247 1729 1251 1730
rect 1255 1734 1259 1735
rect 1255 1729 1259 1730
rect 1295 1734 1299 1735
rect 1295 1729 1299 1730
rect 1319 1734 1323 1735
rect 1319 1729 1323 1730
rect 1343 1734 1347 1735
rect 1343 1729 1347 1730
rect 1136 1726 1138 1729
rect 1246 1728 1252 1729
rect 1134 1725 1140 1726
rect 1134 1721 1135 1725
rect 1139 1721 1140 1725
rect 1246 1724 1247 1728
rect 1251 1724 1252 1728
rect 1246 1723 1252 1724
rect 1294 1728 1300 1729
rect 1294 1724 1295 1728
rect 1299 1724 1300 1728
rect 1294 1723 1300 1724
rect 1342 1728 1348 1729
rect 1342 1724 1343 1728
rect 1347 1724 1348 1728
rect 1342 1723 1348 1724
rect 1134 1720 1140 1721
rect 1368 1712 1370 1770
rect 1384 1769 1386 1781
rect 1456 1769 1458 1781
rect 1470 1775 1476 1776
rect 1470 1771 1471 1775
rect 1475 1771 1476 1775
rect 1470 1770 1476 1771
rect 1382 1768 1388 1769
rect 1382 1764 1383 1768
rect 1387 1764 1388 1768
rect 1382 1763 1388 1764
rect 1454 1768 1460 1769
rect 1454 1764 1455 1768
rect 1459 1764 1460 1768
rect 1454 1763 1460 1764
rect 1472 1756 1474 1770
rect 1528 1769 1530 1781
rect 1568 1780 1570 1810
rect 1646 1804 1652 1805
rect 1646 1800 1647 1804
rect 1651 1800 1652 1804
rect 1646 1799 1652 1800
rect 1750 1804 1756 1805
rect 1750 1800 1751 1804
rect 1755 1800 1756 1804
rect 1750 1799 1756 1800
rect 1854 1804 1860 1805
rect 1854 1800 1855 1804
rect 1859 1800 1860 1804
rect 1854 1799 1860 1800
rect 1648 1787 1650 1799
rect 1714 1795 1720 1796
rect 1714 1791 1715 1795
rect 1719 1791 1720 1795
rect 1714 1790 1720 1791
rect 1607 1786 1611 1787
rect 1607 1781 1611 1782
rect 1647 1786 1651 1787
rect 1647 1781 1651 1782
rect 1687 1786 1691 1787
rect 1687 1781 1691 1782
rect 1566 1779 1572 1780
rect 1542 1775 1548 1776
rect 1542 1771 1543 1775
rect 1547 1771 1548 1775
rect 1566 1775 1567 1779
rect 1571 1775 1572 1779
rect 1566 1774 1572 1775
rect 1542 1770 1548 1771
rect 1526 1768 1532 1769
rect 1526 1764 1527 1768
rect 1531 1764 1532 1768
rect 1526 1763 1532 1764
rect 1544 1756 1546 1770
rect 1608 1769 1610 1781
rect 1688 1769 1690 1781
rect 1694 1775 1700 1776
rect 1694 1771 1695 1775
rect 1699 1771 1700 1775
rect 1694 1770 1700 1771
rect 1702 1775 1708 1776
rect 1702 1771 1703 1775
rect 1707 1771 1708 1775
rect 1702 1770 1708 1771
rect 1606 1768 1612 1769
rect 1606 1764 1607 1768
rect 1611 1764 1612 1768
rect 1606 1763 1612 1764
rect 1686 1768 1692 1769
rect 1686 1764 1687 1768
rect 1691 1764 1692 1768
rect 1686 1763 1692 1764
rect 1410 1755 1416 1756
rect 1410 1751 1411 1755
rect 1415 1751 1416 1755
rect 1410 1750 1416 1751
rect 1470 1755 1476 1756
rect 1470 1751 1471 1755
rect 1475 1751 1476 1755
rect 1470 1750 1476 1751
rect 1542 1755 1548 1756
rect 1542 1751 1543 1755
rect 1547 1751 1548 1755
rect 1542 1750 1548 1751
rect 1382 1740 1388 1741
rect 1382 1736 1383 1740
rect 1387 1736 1388 1740
rect 1382 1735 1388 1736
rect 1383 1734 1387 1735
rect 1383 1729 1387 1730
rect 1399 1734 1403 1735
rect 1399 1729 1403 1730
rect 1398 1728 1404 1729
rect 1398 1724 1399 1728
rect 1403 1724 1404 1728
rect 1398 1723 1404 1724
rect 1310 1711 1316 1712
rect 1134 1708 1140 1709
rect 1047 1706 1051 1707
rect 1047 1701 1051 1702
rect 1095 1706 1099 1707
rect 1134 1704 1135 1708
rect 1139 1704 1140 1708
rect 1310 1707 1311 1711
rect 1315 1707 1316 1711
rect 1310 1706 1316 1707
rect 1358 1711 1364 1712
rect 1358 1707 1359 1711
rect 1363 1707 1364 1711
rect 1358 1706 1364 1707
rect 1366 1711 1372 1712
rect 1366 1707 1367 1711
rect 1371 1707 1372 1711
rect 1366 1706 1372 1707
rect 1134 1703 1140 1704
rect 1095 1701 1099 1702
rect 998 1695 1004 1696
rect 998 1691 999 1695
rect 1003 1691 1004 1695
rect 998 1690 1004 1691
rect 1010 1695 1016 1696
rect 1010 1691 1011 1695
rect 1015 1691 1016 1695
rect 1010 1690 1016 1691
rect 918 1688 924 1689
rect 918 1684 919 1688
rect 923 1684 924 1688
rect 918 1683 924 1684
rect 982 1688 988 1689
rect 982 1684 983 1688
rect 987 1684 988 1688
rect 982 1683 988 1684
rect 1000 1676 1002 1690
rect 1048 1689 1050 1701
rect 1046 1688 1052 1689
rect 1046 1684 1047 1688
rect 1051 1684 1052 1688
rect 1046 1683 1052 1684
rect 1096 1681 1098 1701
rect 1094 1680 1100 1681
rect 1094 1676 1095 1680
rect 1099 1676 1100 1680
rect 1136 1679 1138 1703
rect 1246 1700 1252 1701
rect 1246 1696 1247 1700
rect 1251 1696 1252 1700
rect 1246 1695 1252 1696
rect 1294 1700 1300 1701
rect 1294 1696 1295 1700
rect 1299 1696 1300 1700
rect 1294 1695 1300 1696
rect 1248 1679 1250 1695
rect 1286 1691 1292 1692
rect 1286 1687 1287 1691
rect 1291 1687 1292 1691
rect 1286 1686 1292 1687
rect 998 1675 1004 1676
rect 998 1671 999 1675
rect 1003 1671 1004 1675
rect 998 1670 1004 1671
rect 1034 1675 1040 1676
rect 1094 1675 1100 1676
rect 1135 1678 1139 1679
rect 1034 1671 1035 1675
rect 1039 1671 1040 1675
rect 1135 1673 1139 1674
rect 1247 1678 1251 1679
rect 1247 1673 1251 1674
rect 1263 1678 1267 1679
rect 1263 1673 1267 1674
rect 1034 1670 1040 1671
rect 918 1660 924 1661
rect 918 1656 919 1660
rect 923 1656 924 1660
rect 918 1655 924 1656
rect 982 1660 988 1661
rect 982 1656 983 1660
rect 987 1656 988 1660
rect 982 1655 988 1656
rect 920 1651 922 1655
rect 984 1651 986 1655
rect 903 1650 907 1651
rect 903 1645 907 1646
rect 919 1650 923 1651
rect 919 1645 923 1646
rect 959 1650 963 1651
rect 959 1645 963 1646
rect 983 1650 987 1651
rect 983 1645 987 1646
rect 1007 1650 1011 1651
rect 1007 1645 1011 1646
rect 902 1644 908 1645
rect 902 1640 903 1644
rect 907 1640 908 1644
rect 902 1639 908 1640
rect 958 1644 964 1645
rect 958 1640 959 1644
rect 963 1640 964 1644
rect 958 1639 964 1640
rect 1006 1644 1012 1645
rect 1006 1640 1007 1644
rect 1011 1640 1012 1644
rect 1006 1639 1012 1640
rect 670 1627 676 1628
rect 670 1623 671 1627
rect 675 1623 676 1627
rect 670 1622 676 1623
rect 802 1627 808 1628
rect 802 1623 803 1627
rect 807 1623 808 1627
rect 802 1622 808 1623
rect 862 1627 868 1628
rect 862 1623 863 1627
rect 867 1623 868 1627
rect 862 1622 868 1623
rect 870 1627 876 1628
rect 870 1623 871 1627
rect 875 1623 876 1627
rect 870 1622 876 1623
rect 930 1627 936 1628
rect 930 1623 931 1627
rect 935 1623 936 1627
rect 930 1622 936 1623
rect 938 1627 944 1628
rect 938 1623 939 1627
rect 943 1623 944 1627
rect 938 1622 944 1623
rect 654 1616 660 1617
rect 654 1612 655 1616
rect 659 1612 660 1616
rect 654 1611 660 1612
rect 610 1607 616 1608
rect 610 1603 611 1607
rect 615 1603 616 1607
rect 610 1602 616 1603
rect 656 1599 658 1611
rect 672 1608 674 1622
rect 778 1619 784 1620
rect 726 1616 732 1617
rect 726 1612 727 1616
rect 731 1612 732 1616
rect 778 1615 779 1619
rect 783 1615 784 1619
rect 778 1614 784 1615
rect 790 1616 796 1617
rect 726 1611 732 1612
rect 670 1607 676 1608
rect 670 1603 671 1607
rect 675 1603 676 1607
rect 670 1602 676 1603
rect 728 1599 730 1611
rect 766 1607 772 1608
rect 766 1603 767 1607
rect 771 1603 772 1607
rect 766 1602 772 1603
rect 503 1598 507 1599
rect 503 1593 507 1594
rect 527 1598 531 1599
rect 527 1593 531 1594
rect 583 1598 587 1599
rect 583 1593 587 1594
rect 599 1598 603 1599
rect 599 1593 603 1594
rect 655 1598 659 1599
rect 655 1593 659 1594
rect 671 1598 675 1599
rect 671 1593 675 1594
rect 727 1598 731 1599
rect 727 1593 731 1594
rect 743 1598 747 1599
rect 743 1593 747 1594
rect 528 1581 530 1593
rect 590 1587 596 1588
rect 590 1583 591 1587
rect 595 1583 596 1587
rect 590 1582 596 1583
rect 526 1580 532 1581
rect 526 1576 527 1580
rect 531 1576 532 1580
rect 526 1575 532 1576
rect 110 1567 116 1568
rect 182 1567 188 1568
rect 182 1563 183 1567
rect 187 1563 188 1567
rect 182 1562 188 1563
rect 482 1567 488 1568
rect 482 1563 483 1567
rect 487 1563 488 1567
rect 482 1562 488 1563
rect 110 1555 116 1556
rect 110 1551 111 1555
rect 115 1551 116 1555
rect 110 1550 116 1551
rect 134 1552 140 1553
rect 112 1547 114 1550
rect 134 1548 135 1552
rect 139 1548 140 1552
rect 134 1547 140 1548
rect 174 1552 180 1553
rect 174 1548 175 1552
rect 179 1548 180 1552
rect 174 1547 180 1548
rect 230 1552 236 1553
rect 230 1548 231 1552
rect 235 1548 236 1552
rect 230 1547 236 1548
rect 302 1552 308 1553
rect 302 1548 303 1552
rect 307 1548 308 1552
rect 302 1547 308 1548
rect 374 1552 380 1553
rect 374 1548 375 1552
rect 379 1548 380 1552
rect 374 1547 380 1548
rect 454 1552 460 1553
rect 454 1548 455 1552
rect 459 1548 460 1552
rect 454 1547 460 1548
rect 526 1552 532 1553
rect 526 1548 527 1552
rect 531 1548 532 1552
rect 526 1547 532 1548
rect 111 1546 115 1547
rect 111 1541 115 1542
rect 135 1546 139 1547
rect 135 1541 139 1542
rect 175 1546 179 1547
rect 175 1541 179 1542
rect 231 1546 235 1547
rect 231 1541 235 1542
rect 303 1546 307 1547
rect 303 1541 307 1542
rect 311 1546 315 1547
rect 311 1541 315 1542
rect 375 1546 379 1547
rect 375 1541 379 1542
rect 391 1546 395 1547
rect 391 1541 395 1542
rect 455 1546 459 1547
rect 455 1541 459 1542
rect 479 1546 483 1547
rect 479 1541 483 1542
rect 527 1546 531 1547
rect 527 1541 531 1542
rect 567 1546 571 1547
rect 567 1541 571 1542
rect 112 1538 114 1541
rect 134 1540 140 1541
rect 110 1537 116 1538
rect 110 1533 111 1537
rect 115 1533 116 1537
rect 134 1536 135 1540
rect 139 1536 140 1540
rect 134 1535 140 1536
rect 174 1540 180 1541
rect 174 1536 175 1540
rect 179 1536 180 1540
rect 174 1535 180 1536
rect 230 1540 236 1541
rect 230 1536 231 1540
rect 235 1536 236 1540
rect 230 1535 236 1536
rect 310 1540 316 1541
rect 310 1536 311 1540
rect 315 1536 316 1540
rect 310 1535 316 1536
rect 390 1540 396 1541
rect 390 1536 391 1540
rect 395 1536 396 1540
rect 390 1535 396 1536
rect 478 1540 484 1541
rect 478 1536 479 1540
rect 483 1536 484 1540
rect 478 1535 484 1536
rect 566 1540 572 1541
rect 566 1536 567 1540
rect 571 1536 572 1540
rect 566 1535 572 1536
rect 110 1532 116 1533
rect 592 1524 594 1582
rect 600 1581 602 1593
rect 606 1587 612 1588
rect 606 1583 607 1587
rect 611 1583 612 1587
rect 606 1582 612 1583
rect 598 1580 604 1581
rect 598 1576 599 1580
rect 603 1576 604 1580
rect 598 1575 604 1576
rect 608 1568 610 1582
rect 672 1581 674 1593
rect 706 1587 712 1588
rect 706 1583 707 1587
rect 711 1583 712 1587
rect 706 1582 712 1583
rect 670 1580 676 1581
rect 670 1576 671 1580
rect 675 1576 676 1580
rect 670 1575 676 1576
rect 708 1568 710 1582
rect 744 1581 746 1593
rect 742 1580 748 1581
rect 742 1576 743 1580
rect 747 1576 748 1580
rect 742 1575 748 1576
rect 768 1568 770 1602
rect 780 1588 782 1614
rect 790 1612 791 1616
rect 795 1612 796 1616
rect 790 1611 796 1612
rect 792 1599 794 1611
rect 804 1608 806 1622
rect 846 1616 852 1617
rect 846 1612 847 1616
rect 851 1612 852 1616
rect 846 1611 852 1612
rect 802 1607 808 1608
rect 802 1603 803 1607
rect 807 1603 808 1607
rect 802 1602 808 1603
rect 848 1599 850 1611
rect 864 1608 866 1622
rect 902 1616 908 1617
rect 902 1612 903 1616
rect 907 1612 908 1616
rect 902 1611 908 1612
rect 862 1607 868 1608
rect 862 1603 863 1607
rect 867 1603 868 1607
rect 862 1602 868 1603
rect 904 1599 906 1611
rect 932 1600 934 1622
rect 940 1608 942 1622
rect 958 1616 964 1617
rect 958 1612 959 1616
rect 963 1612 964 1616
rect 958 1611 964 1612
rect 1006 1616 1012 1617
rect 1006 1612 1007 1616
rect 1011 1612 1012 1616
rect 1006 1611 1012 1612
rect 938 1607 944 1608
rect 938 1603 939 1607
rect 943 1603 944 1607
rect 938 1602 944 1603
rect 930 1599 936 1600
rect 960 1599 962 1611
rect 1008 1599 1010 1611
rect 1036 1608 1038 1670
rect 1094 1663 1100 1664
rect 1046 1660 1052 1661
rect 1046 1656 1047 1660
rect 1051 1656 1052 1660
rect 1094 1659 1095 1663
rect 1099 1659 1100 1663
rect 1094 1658 1100 1659
rect 1046 1655 1052 1656
rect 1048 1651 1050 1655
rect 1096 1651 1098 1658
rect 1136 1653 1138 1673
rect 1264 1661 1266 1673
rect 1262 1660 1268 1661
rect 1262 1656 1263 1660
rect 1267 1656 1268 1660
rect 1262 1655 1268 1656
rect 1134 1652 1140 1653
rect 1047 1650 1051 1651
rect 1047 1645 1051 1646
rect 1095 1650 1099 1651
rect 1134 1648 1135 1652
rect 1139 1648 1140 1652
rect 1288 1648 1290 1686
rect 1296 1679 1298 1695
rect 1312 1692 1314 1706
rect 1342 1700 1348 1701
rect 1342 1696 1343 1700
rect 1347 1696 1348 1700
rect 1342 1695 1348 1696
rect 1310 1691 1316 1692
rect 1310 1687 1311 1691
rect 1315 1687 1316 1691
rect 1310 1686 1316 1687
rect 1344 1679 1346 1695
rect 1360 1692 1362 1706
rect 1398 1700 1404 1701
rect 1398 1696 1399 1700
rect 1403 1696 1404 1700
rect 1398 1695 1404 1696
rect 1358 1691 1364 1692
rect 1358 1687 1359 1691
rect 1363 1687 1364 1691
rect 1358 1686 1364 1687
rect 1400 1679 1402 1695
rect 1412 1692 1414 1750
rect 1454 1740 1460 1741
rect 1454 1736 1455 1740
rect 1459 1736 1460 1740
rect 1454 1735 1460 1736
rect 1526 1740 1532 1741
rect 1526 1736 1527 1740
rect 1531 1736 1532 1740
rect 1526 1735 1532 1736
rect 1606 1740 1612 1741
rect 1606 1736 1607 1740
rect 1611 1736 1612 1740
rect 1606 1735 1612 1736
rect 1686 1740 1692 1741
rect 1686 1736 1687 1740
rect 1691 1736 1692 1740
rect 1686 1735 1692 1736
rect 1455 1734 1459 1735
rect 1455 1729 1459 1730
rect 1463 1734 1467 1735
rect 1463 1729 1467 1730
rect 1527 1734 1531 1735
rect 1527 1729 1531 1730
rect 1599 1734 1603 1735
rect 1599 1729 1603 1730
rect 1607 1734 1611 1735
rect 1607 1729 1611 1730
rect 1671 1734 1675 1735
rect 1671 1729 1675 1730
rect 1687 1734 1691 1735
rect 1687 1729 1691 1730
rect 1462 1728 1468 1729
rect 1462 1724 1463 1728
rect 1467 1724 1468 1728
rect 1462 1723 1468 1724
rect 1526 1728 1532 1729
rect 1526 1724 1527 1728
rect 1531 1724 1532 1728
rect 1526 1723 1532 1724
rect 1598 1728 1604 1729
rect 1598 1724 1599 1728
rect 1603 1724 1604 1728
rect 1598 1723 1604 1724
rect 1670 1728 1676 1729
rect 1670 1724 1671 1728
rect 1675 1724 1676 1728
rect 1670 1723 1676 1724
rect 1696 1712 1698 1770
rect 1704 1756 1706 1770
rect 1716 1756 1718 1790
rect 1752 1787 1754 1799
rect 1856 1787 1858 1799
rect 1751 1786 1755 1787
rect 1751 1781 1755 1782
rect 1767 1786 1771 1787
rect 1767 1781 1771 1782
rect 1847 1786 1851 1787
rect 1847 1781 1851 1782
rect 1855 1786 1859 1787
rect 1855 1781 1859 1782
rect 1927 1786 1931 1787
rect 1927 1781 1931 1782
rect 1768 1769 1770 1781
rect 1848 1769 1850 1781
rect 1862 1775 1868 1776
rect 1862 1771 1863 1775
rect 1867 1771 1868 1775
rect 1862 1770 1868 1771
rect 1766 1768 1772 1769
rect 1766 1764 1767 1768
rect 1771 1764 1772 1768
rect 1766 1763 1772 1764
rect 1846 1768 1852 1769
rect 1846 1764 1847 1768
rect 1851 1764 1852 1768
rect 1846 1763 1852 1764
rect 1864 1756 1866 1770
rect 1928 1769 1930 1781
rect 1952 1776 1954 1810
rect 1960 1796 1962 1810
rect 1966 1804 1972 1805
rect 1966 1800 1967 1804
rect 1971 1800 1972 1804
rect 1966 1799 1972 1800
rect 2070 1804 2076 1805
rect 2070 1800 2071 1804
rect 2075 1800 2076 1804
rect 2070 1799 2076 1800
rect 1958 1795 1964 1796
rect 1958 1791 1959 1795
rect 1963 1791 1964 1795
rect 1958 1790 1964 1791
rect 1968 1787 1970 1799
rect 2030 1795 2036 1796
rect 2030 1791 2031 1795
rect 2035 1791 2036 1795
rect 2030 1790 2036 1791
rect 1967 1786 1971 1787
rect 1967 1781 1971 1782
rect 2007 1786 2011 1787
rect 2007 1781 2011 1782
rect 1942 1775 1948 1776
rect 1942 1771 1943 1775
rect 1947 1771 1948 1775
rect 1942 1770 1948 1771
rect 1950 1775 1956 1776
rect 1950 1771 1951 1775
rect 1955 1771 1956 1775
rect 1950 1770 1956 1771
rect 1926 1768 1932 1769
rect 1926 1764 1927 1768
rect 1931 1764 1932 1768
rect 1926 1763 1932 1764
rect 1944 1756 1946 1770
rect 2008 1769 2010 1781
rect 2014 1775 2020 1776
rect 2014 1771 2015 1775
rect 2019 1771 2020 1775
rect 2014 1770 2020 1771
rect 2006 1768 2012 1769
rect 2006 1764 2007 1768
rect 2011 1764 2012 1768
rect 2006 1763 2012 1764
rect 1702 1755 1708 1756
rect 1702 1751 1703 1755
rect 1707 1751 1708 1755
rect 1702 1750 1708 1751
rect 1714 1755 1720 1756
rect 1714 1751 1715 1755
rect 1719 1751 1720 1755
rect 1714 1750 1720 1751
rect 1782 1755 1788 1756
rect 1782 1751 1783 1755
rect 1787 1751 1788 1755
rect 1782 1750 1788 1751
rect 1862 1755 1868 1756
rect 1862 1751 1863 1755
rect 1867 1751 1868 1755
rect 1862 1750 1868 1751
rect 1942 1755 1948 1756
rect 1942 1751 1943 1755
rect 1947 1751 1948 1755
rect 1942 1750 1948 1751
rect 1766 1740 1772 1741
rect 1766 1736 1767 1740
rect 1771 1736 1772 1740
rect 1766 1735 1772 1736
rect 1743 1734 1747 1735
rect 1743 1729 1747 1730
rect 1767 1734 1771 1735
rect 1767 1729 1771 1730
rect 1742 1728 1748 1729
rect 1742 1724 1743 1728
rect 1747 1724 1748 1728
rect 1742 1723 1748 1724
rect 1478 1711 1484 1712
rect 1478 1707 1479 1711
rect 1483 1707 1484 1711
rect 1478 1706 1484 1707
rect 1534 1711 1540 1712
rect 1534 1707 1535 1711
rect 1539 1707 1540 1711
rect 1534 1706 1540 1707
rect 1542 1711 1548 1712
rect 1542 1707 1543 1711
rect 1547 1707 1548 1711
rect 1542 1706 1548 1707
rect 1686 1711 1692 1712
rect 1686 1707 1687 1711
rect 1691 1707 1692 1711
rect 1686 1706 1692 1707
rect 1694 1711 1700 1712
rect 1694 1707 1695 1711
rect 1699 1707 1700 1711
rect 1694 1706 1700 1707
rect 1462 1700 1468 1701
rect 1462 1696 1463 1700
rect 1467 1696 1468 1700
rect 1462 1695 1468 1696
rect 1410 1691 1416 1692
rect 1410 1687 1411 1691
rect 1415 1687 1416 1691
rect 1410 1686 1416 1687
rect 1464 1679 1466 1695
rect 1480 1692 1482 1706
rect 1526 1700 1532 1701
rect 1526 1696 1527 1700
rect 1531 1696 1532 1700
rect 1526 1695 1532 1696
rect 1478 1691 1484 1692
rect 1478 1687 1479 1691
rect 1483 1687 1484 1691
rect 1478 1686 1484 1687
rect 1528 1679 1530 1695
rect 1536 1692 1538 1706
rect 1534 1691 1540 1692
rect 1534 1687 1535 1691
rect 1539 1687 1540 1691
rect 1534 1686 1540 1687
rect 1295 1678 1299 1679
rect 1295 1673 1299 1674
rect 1303 1678 1307 1679
rect 1303 1673 1307 1674
rect 1343 1678 1347 1679
rect 1343 1673 1347 1674
rect 1391 1678 1395 1679
rect 1391 1673 1395 1674
rect 1399 1678 1403 1679
rect 1399 1673 1403 1674
rect 1447 1678 1451 1679
rect 1447 1673 1451 1674
rect 1463 1678 1467 1679
rect 1463 1673 1467 1674
rect 1503 1678 1507 1679
rect 1503 1673 1507 1674
rect 1527 1678 1531 1679
rect 1527 1673 1531 1674
rect 1304 1661 1306 1673
rect 1318 1667 1324 1668
rect 1318 1663 1319 1667
rect 1323 1663 1324 1667
rect 1318 1662 1324 1663
rect 1302 1660 1308 1661
rect 1302 1656 1303 1660
rect 1307 1656 1308 1660
rect 1302 1655 1308 1656
rect 1320 1648 1322 1662
rect 1344 1661 1346 1673
rect 1358 1667 1364 1668
rect 1358 1663 1359 1667
rect 1363 1663 1364 1667
rect 1358 1662 1364 1663
rect 1342 1660 1348 1661
rect 1342 1656 1343 1660
rect 1347 1656 1348 1660
rect 1342 1655 1348 1656
rect 1360 1648 1362 1662
rect 1392 1661 1394 1673
rect 1406 1667 1412 1668
rect 1406 1663 1407 1667
rect 1411 1663 1412 1667
rect 1406 1662 1412 1663
rect 1390 1660 1396 1661
rect 1390 1656 1391 1660
rect 1395 1656 1396 1660
rect 1390 1655 1396 1656
rect 1408 1648 1410 1662
rect 1448 1661 1450 1673
rect 1462 1667 1468 1668
rect 1462 1663 1463 1667
rect 1467 1663 1468 1667
rect 1462 1662 1468 1663
rect 1446 1660 1452 1661
rect 1446 1656 1447 1660
rect 1451 1656 1452 1660
rect 1446 1655 1452 1656
rect 1464 1648 1466 1662
rect 1504 1661 1506 1673
rect 1544 1672 1546 1706
rect 1598 1700 1604 1701
rect 1598 1696 1599 1700
rect 1603 1696 1604 1700
rect 1598 1695 1604 1696
rect 1670 1700 1676 1701
rect 1670 1696 1671 1700
rect 1675 1696 1676 1700
rect 1670 1695 1676 1696
rect 1600 1679 1602 1695
rect 1610 1691 1616 1692
rect 1610 1687 1611 1691
rect 1615 1687 1616 1691
rect 1610 1686 1616 1687
rect 1567 1678 1571 1679
rect 1567 1673 1571 1674
rect 1599 1678 1603 1679
rect 1599 1673 1603 1674
rect 1542 1671 1548 1672
rect 1518 1667 1524 1668
rect 1518 1663 1519 1667
rect 1523 1663 1524 1667
rect 1542 1667 1543 1671
rect 1547 1667 1548 1671
rect 1542 1666 1548 1667
rect 1518 1662 1524 1663
rect 1502 1660 1508 1661
rect 1502 1656 1503 1660
rect 1507 1656 1508 1660
rect 1502 1655 1508 1656
rect 1520 1648 1522 1662
rect 1568 1661 1570 1673
rect 1566 1660 1572 1661
rect 1566 1656 1567 1660
rect 1571 1656 1572 1660
rect 1566 1655 1572 1656
rect 1612 1648 1614 1686
rect 1672 1679 1674 1695
rect 1688 1692 1690 1706
rect 1742 1700 1748 1701
rect 1742 1696 1743 1700
rect 1747 1696 1748 1700
rect 1784 1696 1786 1750
rect 1846 1740 1852 1741
rect 1846 1736 1847 1740
rect 1851 1736 1852 1740
rect 1846 1735 1852 1736
rect 1926 1740 1932 1741
rect 1926 1736 1927 1740
rect 1931 1736 1932 1740
rect 1926 1735 1932 1736
rect 2006 1740 2012 1741
rect 2006 1736 2007 1740
rect 2011 1736 2012 1740
rect 2006 1735 2012 1736
rect 1807 1734 1811 1735
rect 1807 1729 1811 1730
rect 1847 1734 1851 1735
rect 1847 1729 1851 1730
rect 1879 1734 1883 1735
rect 1879 1729 1883 1730
rect 1927 1734 1931 1735
rect 1927 1729 1931 1730
rect 1951 1734 1955 1735
rect 1951 1729 1955 1730
rect 2007 1734 2011 1735
rect 2007 1729 2011 1730
rect 1806 1728 1812 1729
rect 1806 1724 1807 1728
rect 1811 1724 1812 1728
rect 1806 1723 1812 1724
rect 1878 1728 1884 1729
rect 1878 1724 1879 1728
rect 1883 1724 1884 1728
rect 1878 1723 1884 1724
rect 1950 1728 1956 1729
rect 1950 1724 1951 1728
rect 1955 1724 1956 1728
rect 1950 1723 1956 1724
rect 2016 1712 2018 1770
rect 2032 1756 2034 1790
rect 2072 1787 2074 1799
rect 2080 1796 2082 1854
rect 2118 1847 2124 1848
rect 2118 1843 2119 1847
rect 2123 1843 2124 1847
rect 2118 1842 2124 1843
rect 2120 1839 2122 1842
rect 2119 1838 2123 1839
rect 2119 1833 2123 1834
rect 2120 1830 2122 1833
rect 2118 1829 2124 1830
rect 2118 1825 2119 1829
rect 2123 1825 2124 1829
rect 2118 1824 2124 1825
rect 2094 1815 2100 1816
rect 2094 1811 2095 1815
rect 2099 1811 2100 1815
rect 2094 1810 2100 1811
rect 2118 1812 2124 1813
rect 2078 1795 2084 1796
rect 2078 1791 2079 1795
rect 2083 1791 2084 1795
rect 2078 1790 2084 1791
rect 2071 1786 2075 1787
rect 2071 1781 2075 1782
rect 2072 1769 2074 1781
rect 2096 1776 2098 1810
rect 2118 1808 2119 1812
rect 2123 1808 2124 1812
rect 2118 1807 2124 1808
rect 2120 1787 2122 1807
rect 2119 1786 2123 1787
rect 2119 1781 2123 1782
rect 2094 1775 2100 1776
rect 2094 1771 2095 1775
rect 2099 1771 2100 1775
rect 2094 1770 2100 1771
rect 2070 1768 2076 1769
rect 2070 1764 2071 1768
rect 2075 1764 2076 1768
rect 2070 1763 2076 1764
rect 2120 1761 2122 1781
rect 2118 1760 2124 1761
rect 2118 1756 2119 1760
rect 2123 1756 2124 1760
rect 2030 1755 2036 1756
rect 2030 1751 2031 1755
rect 2035 1751 2036 1755
rect 2030 1750 2036 1751
rect 2094 1755 2100 1756
rect 2118 1755 2124 1756
rect 2094 1751 2095 1755
rect 2099 1751 2100 1755
rect 2094 1750 2100 1751
rect 2070 1740 2076 1741
rect 2070 1736 2071 1740
rect 2075 1736 2076 1740
rect 2070 1735 2076 1736
rect 2023 1734 2027 1735
rect 2023 1729 2027 1730
rect 2071 1734 2075 1735
rect 2071 1729 2075 1730
rect 2022 1728 2028 1729
rect 2022 1724 2023 1728
rect 2027 1724 2028 1728
rect 2022 1723 2028 1724
rect 2070 1728 2076 1729
rect 2070 1724 2071 1728
rect 2075 1724 2076 1728
rect 2070 1723 2076 1724
rect 1814 1711 1820 1712
rect 1814 1707 1815 1711
rect 1819 1707 1820 1711
rect 1814 1706 1820 1707
rect 1894 1711 1900 1712
rect 1894 1707 1895 1711
rect 1899 1707 1900 1711
rect 1894 1706 1900 1707
rect 1934 1711 1940 1712
rect 1934 1707 1935 1711
rect 1939 1707 1940 1711
rect 1934 1706 1940 1707
rect 2014 1711 2020 1712
rect 2014 1707 2015 1711
rect 2019 1707 2020 1711
rect 2014 1706 2020 1707
rect 2046 1711 2052 1712
rect 2046 1707 2047 1711
rect 2051 1707 2052 1711
rect 2046 1706 2052 1707
rect 1806 1700 1812 1701
rect 1806 1696 1807 1700
rect 1811 1696 1812 1700
rect 1742 1695 1748 1696
rect 1782 1695 1788 1696
rect 1806 1695 1812 1696
rect 1686 1691 1692 1692
rect 1686 1687 1687 1691
rect 1691 1687 1692 1691
rect 1686 1686 1692 1687
rect 1744 1679 1746 1695
rect 1782 1691 1783 1695
rect 1787 1691 1788 1695
rect 1782 1690 1788 1691
rect 1808 1679 1810 1695
rect 1816 1692 1818 1706
rect 1878 1700 1884 1701
rect 1878 1696 1879 1700
rect 1883 1696 1884 1700
rect 1878 1695 1884 1696
rect 1814 1691 1820 1692
rect 1814 1687 1815 1691
rect 1819 1687 1820 1691
rect 1814 1686 1820 1687
rect 1880 1679 1882 1695
rect 1896 1692 1898 1706
rect 1894 1691 1900 1692
rect 1894 1687 1895 1691
rect 1899 1687 1900 1691
rect 1894 1686 1900 1687
rect 1631 1678 1635 1679
rect 1631 1673 1635 1674
rect 1671 1678 1675 1679
rect 1671 1673 1675 1674
rect 1695 1678 1699 1679
rect 1695 1673 1699 1674
rect 1743 1678 1747 1679
rect 1743 1673 1747 1674
rect 1759 1678 1763 1679
rect 1759 1673 1763 1674
rect 1807 1678 1811 1679
rect 1807 1673 1811 1674
rect 1831 1678 1835 1679
rect 1831 1673 1835 1674
rect 1879 1678 1883 1679
rect 1879 1673 1883 1674
rect 1911 1678 1915 1679
rect 1911 1673 1915 1674
rect 1632 1661 1634 1673
rect 1642 1667 1648 1668
rect 1642 1663 1643 1667
rect 1647 1663 1648 1667
rect 1642 1662 1648 1663
rect 1650 1667 1656 1668
rect 1650 1663 1651 1667
rect 1655 1663 1656 1667
rect 1650 1662 1656 1663
rect 1630 1660 1636 1661
rect 1630 1656 1631 1660
rect 1635 1656 1636 1660
rect 1630 1655 1636 1656
rect 1644 1648 1646 1662
rect 1134 1647 1140 1648
rect 1286 1647 1292 1648
rect 1095 1645 1099 1646
rect 1046 1644 1052 1645
rect 1046 1640 1047 1644
rect 1051 1640 1052 1644
rect 1096 1642 1098 1645
rect 1286 1643 1287 1647
rect 1291 1643 1292 1647
rect 1286 1642 1292 1643
rect 1318 1647 1324 1648
rect 1318 1643 1319 1647
rect 1323 1643 1324 1647
rect 1318 1642 1324 1643
rect 1358 1647 1364 1648
rect 1358 1643 1359 1647
rect 1363 1643 1364 1647
rect 1358 1642 1364 1643
rect 1406 1647 1412 1648
rect 1406 1643 1407 1647
rect 1411 1643 1412 1647
rect 1406 1642 1412 1643
rect 1462 1647 1468 1648
rect 1462 1643 1463 1647
rect 1467 1643 1468 1647
rect 1462 1642 1468 1643
rect 1518 1647 1524 1648
rect 1518 1643 1519 1647
rect 1523 1643 1524 1647
rect 1518 1642 1524 1643
rect 1610 1647 1616 1648
rect 1610 1643 1611 1647
rect 1615 1643 1616 1647
rect 1610 1642 1616 1643
rect 1642 1647 1648 1648
rect 1642 1643 1643 1647
rect 1647 1643 1648 1647
rect 1642 1642 1648 1643
rect 1046 1639 1052 1640
rect 1094 1641 1100 1642
rect 1094 1637 1095 1641
rect 1099 1637 1100 1641
rect 1094 1636 1100 1637
rect 1134 1635 1140 1636
rect 1114 1631 1120 1632
rect 1114 1627 1115 1631
rect 1119 1627 1120 1631
rect 1134 1631 1135 1635
rect 1139 1631 1140 1635
rect 1134 1630 1140 1631
rect 1262 1632 1268 1633
rect 1114 1626 1120 1627
rect 1094 1624 1100 1625
rect 1094 1620 1095 1624
rect 1099 1620 1100 1624
rect 1094 1619 1100 1620
rect 1046 1616 1052 1617
rect 1046 1612 1047 1616
rect 1051 1612 1052 1616
rect 1046 1611 1052 1612
rect 1034 1607 1040 1608
rect 1034 1603 1035 1607
rect 1039 1603 1040 1607
rect 1034 1602 1040 1603
rect 1048 1599 1050 1611
rect 1096 1599 1098 1619
rect 791 1598 795 1599
rect 791 1593 795 1594
rect 815 1598 819 1599
rect 815 1593 819 1594
rect 847 1598 851 1599
rect 847 1593 851 1594
rect 887 1598 891 1599
rect 887 1593 891 1594
rect 903 1598 907 1599
rect 930 1595 931 1599
rect 935 1595 936 1599
rect 930 1594 936 1595
rect 959 1598 963 1599
rect 903 1593 907 1594
rect 959 1593 963 1594
rect 1007 1598 1011 1599
rect 1007 1593 1011 1594
rect 1047 1598 1051 1599
rect 1047 1593 1051 1594
rect 1095 1598 1099 1599
rect 1095 1593 1099 1594
rect 778 1587 784 1588
rect 778 1583 779 1587
rect 783 1583 784 1587
rect 778 1582 784 1583
rect 816 1581 818 1593
rect 888 1581 890 1593
rect 814 1580 820 1581
rect 814 1576 815 1580
rect 819 1576 820 1580
rect 814 1575 820 1576
rect 886 1580 892 1581
rect 886 1576 887 1580
rect 891 1576 892 1580
rect 886 1575 892 1576
rect 1096 1573 1098 1593
rect 1094 1572 1100 1573
rect 1116 1572 1118 1626
rect 1136 1615 1138 1630
rect 1262 1628 1263 1632
rect 1267 1628 1268 1632
rect 1262 1627 1268 1628
rect 1302 1632 1308 1633
rect 1302 1628 1303 1632
rect 1307 1628 1308 1632
rect 1302 1627 1308 1628
rect 1342 1632 1348 1633
rect 1342 1628 1343 1632
rect 1347 1628 1348 1632
rect 1342 1627 1348 1628
rect 1390 1632 1396 1633
rect 1390 1628 1391 1632
rect 1395 1628 1396 1632
rect 1390 1627 1396 1628
rect 1446 1632 1452 1633
rect 1446 1628 1447 1632
rect 1451 1628 1452 1632
rect 1446 1627 1452 1628
rect 1502 1632 1508 1633
rect 1502 1628 1503 1632
rect 1507 1628 1508 1632
rect 1502 1627 1508 1628
rect 1566 1632 1572 1633
rect 1566 1628 1567 1632
rect 1571 1628 1572 1632
rect 1566 1627 1572 1628
rect 1630 1632 1636 1633
rect 1630 1628 1631 1632
rect 1635 1628 1636 1632
rect 1630 1627 1636 1628
rect 1264 1615 1266 1627
rect 1304 1615 1306 1627
rect 1344 1615 1346 1627
rect 1392 1615 1394 1627
rect 1448 1615 1450 1627
rect 1504 1615 1506 1627
rect 1568 1615 1570 1627
rect 1632 1615 1634 1627
rect 1135 1614 1139 1615
rect 1135 1609 1139 1610
rect 1159 1614 1163 1615
rect 1159 1609 1163 1610
rect 1215 1614 1219 1615
rect 1215 1609 1219 1610
rect 1263 1614 1267 1615
rect 1263 1609 1267 1610
rect 1303 1614 1307 1615
rect 1303 1609 1307 1610
rect 1343 1614 1347 1615
rect 1343 1609 1347 1610
rect 1383 1614 1387 1615
rect 1383 1609 1387 1610
rect 1391 1614 1395 1615
rect 1391 1609 1395 1610
rect 1447 1614 1451 1615
rect 1447 1609 1451 1610
rect 1463 1614 1467 1615
rect 1463 1609 1467 1610
rect 1503 1614 1507 1615
rect 1503 1609 1507 1610
rect 1543 1614 1547 1615
rect 1543 1609 1547 1610
rect 1567 1614 1571 1615
rect 1567 1609 1571 1610
rect 1623 1614 1627 1615
rect 1623 1609 1627 1610
rect 1631 1614 1635 1615
rect 1631 1609 1635 1610
rect 1136 1606 1138 1609
rect 1158 1608 1164 1609
rect 1134 1605 1140 1606
rect 1134 1601 1135 1605
rect 1139 1601 1140 1605
rect 1158 1604 1159 1608
rect 1163 1604 1164 1608
rect 1158 1603 1164 1604
rect 1214 1608 1220 1609
rect 1214 1604 1215 1608
rect 1219 1604 1220 1608
rect 1214 1603 1220 1604
rect 1302 1608 1308 1609
rect 1302 1604 1303 1608
rect 1307 1604 1308 1608
rect 1302 1603 1308 1604
rect 1382 1608 1388 1609
rect 1382 1604 1383 1608
rect 1387 1604 1388 1608
rect 1382 1603 1388 1604
rect 1462 1608 1468 1609
rect 1462 1604 1463 1608
rect 1467 1604 1468 1608
rect 1462 1603 1468 1604
rect 1542 1608 1548 1609
rect 1542 1604 1543 1608
rect 1547 1604 1548 1608
rect 1542 1603 1548 1604
rect 1622 1608 1628 1609
rect 1622 1604 1623 1608
rect 1627 1604 1628 1608
rect 1622 1603 1628 1604
rect 1134 1600 1140 1601
rect 1614 1599 1620 1600
rect 1614 1595 1615 1599
rect 1619 1595 1620 1599
rect 1614 1594 1620 1595
rect 1230 1591 1236 1592
rect 1134 1588 1140 1589
rect 1134 1584 1135 1588
rect 1139 1584 1140 1588
rect 1230 1587 1231 1591
rect 1235 1587 1236 1591
rect 1230 1586 1236 1587
rect 1318 1591 1324 1592
rect 1318 1587 1319 1591
rect 1323 1587 1324 1591
rect 1318 1586 1324 1587
rect 1398 1591 1404 1592
rect 1398 1587 1399 1591
rect 1403 1587 1404 1591
rect 1398 1586 1404 1587
rect 1134 1583 1140 1584
rect 1094 1568 1095 1572
rect 1099 1568 1100 1572
rect 606 1567 612 1568
rect 606 1563 607 1567
rect 611 1563 612 1567
rect 606 1562 612 1563
rect 706 1567 712 1568
rect 706 1563 707 1567
rect 711 1563 712 1567
rect 706 1562 712 1563
rect 766 1567 772 1568
rect 766 1563 767 1567
rect 771 1563 772 1567
rect 766 1562 772 1563
rect 850 1567 856 1568
rect 1094 1567 1100 1568
rect 1114 1571 1120 1572
rect 1114 1567 1115 1571
rect 1119 1567 1120 1571
rect 850 1563 851 1567
rect 855 1563 856 1567
rect 1114 1566 1120 1567
rect 1136 1563 1138 1583
rect 1158 1580 1164 1581
rect 1158 1576 1159 1580
rect 1163 1576 1164 1580
rect 1158 1575 1164 1576
rect 1214 1580 1220 1581
rect 1214 1576 1215 1580
rect 1219 1576 1220 1580
rect 1214 1575 1220 1576
rect 1160 1563 1162 1575
rect 1216 1563 1218 1575
rect 1232 1572 1234 1586
rect 1302 1580 1308 1581
rect 1302 1576 1303 1580
rect 1307 1576 1308 1580
rect 1302 1575 1308 1576
rect 1230 1571 1236 1572
rect 1230 1567 1231 1571
rect 1235 1567 1236 1571
rect 1230 1566 1236 1567
rect 1304 1563 1306 1575
rect 1320 1572 1322 1586
rect 1382 1580 1388 1581
rect 1382 1576 1383 1580
rect 1387 1576 1388 1580
rect 1382 1575 1388 1576
rect 1318 1571 1324 1572
rect 1318 1567 1319 1571
rect 1323 1567 1324 1571
rect 1318 1566 1324 1567
rect 1384 1563 1386 1575
rect 1400 1572 1402 1586
rect 1502 1583 1508 1584
rect 1462 1580 1468 1581
rect 1462 1576 1463 1580
rect 1467 1576 1468 1580
rect 1502 1579 1503 1583
rect 1507 1579 1508 1583
rect 1502 1578 1508 1579
rect 1542 1580 1548 1581
rect 1462 1575 1468 1576
rect 1398 1571 1404 1572
rect 1398 1567 1399 1571
rect 1403 1567 1404 1571
rect 1398 1566 1404 1567
rect 1464 1563 1466 1575
rect 850 1562 856 1563
rect 1135 1562 1139 1563
rect 598 1552 604 1553
rect 598 1548 599 1552
rect 603 1548 604 1552
rect 598 1547 604 1548
rect 670 1552 676 1553
rect 670 1548 671 1552
rect 675 1548 676 1552
rect 670 1547 676 1548
rect 742 1552 748 1553
rect 742 1548 743 1552
rect 747 1548 748 1552
rect 742 1547 748 1548
rect 814 1552 820 1553
rect 814 1548 815 1552
rect 819 1548 820 1552
rect 814 1547 820 1548
rect 599 1546 603 1547
rect 599 1541 603 1542
rect 655 1546 659 1547
rect 655 1541 659 1542
rect 671 1546 675 1547
rect 671 1541 675 1542
rect 743 1546 747 1547
rect 743 1541 747 1542
rect 815 1546 819 1547
rect 815 1541 819 1542
rect 823 1546 827 1547
rect 823 1541 827 1542
rect 654 1540 660 1541
rect 654 1536 655 1540
rect 659 1536 660 1540
rect 654 1535 660 1536
rect 742 1540 748 1541
rect 742 1536 743 1540
rect 747 1536 748 1540
rect 742 1535 748 1536
rect 822 1540 828 1541
rect 822 1536 823 1540
rect 827 1536 828 1540
rect 822 1535 828 1536
rect 162 1523 168 1524
rect 110 1520 116 1521
rect 110 1516 111 1520
rect 115 1516 116 1520
rect 162 1519 163 1523
rect 167 1519 168 1523
rect 162 1518 168 1519
rect 182 1523 188 1524
rect 182 1519 183 1523
rect 187 1519 188 1523
rect 182 1518 188 1519
rect 590 1523 596 1524
rect 590 1519 591 1523
rect 595 1519 596 1523
rect 590 1518 596 1519
rect 110 1515 116 1516
rect 112 1495 114 1515
rect 134 1512 140 1513
rect 134 1508 135 1512
rect 139 1508 140 1512
rect 134 1507 140 1508
rect 136 1495 138 1507
rect 111 1494 115 1495
rect 111 1489 115 1490
rect 135 1494 139 1495
rect 164 1492 166 1518
rect 174 1512 180 1513
rect 174 1508 175 1512
rect 179 1508 180 1512
rect 174 1507 180 1508
rect 176 1495 178 1507
rect 184 1504 186 1518
rect 230 1512 236 1513
rect 230 1508 231 1512
rect 235 1508 236 1512
rect 230 1507 236 1508
rect 310 1512 316 1513
rect 310 1508 311 1512
rect 315 1508 316 1512
rect 310 1507 316 1508
rect 390 1512 396 1513
rect 390 1508 391 1512
rect 395 1508 396 1512
rect 390 1507 396 1508
rect 478 1512 484 1513
rect 478 1508 479 1512
rect 483 1508 484 1512
rect 478 1507 484 1508
rect 566 1512 572 1513
rect 566 1508 567 1512
rect 571 1508 572 1512
rect 566 1507 572 1508
rect 654 1512 660 1513
rect 654 1508 655 1512
rect 659 1508 660 1512
rect 654 1507 660 1508
rect 742 1512 748 1513
rect 742 1508 743 1512
rect 747 1508 748 1512
rect 742 1507 748 1508
rect 822 1512 828 1513
rect 822 1508 823 1512
rect 827 1508 828 1512
rect 822 1507 828 1508
rect 182 1503 188 1504
rect 182 1499 183 1503
rect 187 1499 188 1503
rect 182 1498 188 1499
rect 232 1495 234 1507
rect 312 1495 314 1507
rect 392 1495 394 1507
rect 434 1503 440 1504
rect 434 1499 435 1503
rect 439 1499 440 1503
rect 432 1498 440 1499
rect 432 1497 438 1498
rect 175 1494 179 1495
rect 135 1489 139 1490
rect 162 1491 168 1492
rect 112 1469 114 1489
rect 136 1477 138 1489
rect 162 1487 163 1491
rect 167 1487 168 1491
rect 175 1489 179 1490
rect 199 1494 203 1495
rect 199 1489 203 1490
rect 231 1494 235 1495
rect 231 1489 235 1490
rect 279 1494 283 1495
rect 279 1489 283 1490
rect 311 1494 315 1495
rect 311 1489 315 1490
rect 359 1494 363 1495
rect 359 1489 363 1490
rect 391 1494 395 1495
rect 391 1489 395 1490
rect 162 1486 168 1487
rect 200 1477 202 1489
rect 214 1483 220 1484
rect 214 1479 215 1483
rect 219 1479 220 1483
rect 214 1478 220 1479
rect 134 1476 140 1477
rect 134 1472 135 1476
rect 139 1472 140 1476
rect 134 1471 140 1472
rect 198 1476 204 1477
rect 198 1472 199 1476
rect 203 1472 204 1476
rect 198 1471 204 1472
rect 110 1468 116 1469
rect 110 1464 111 1468
rect 115 1464 116 1468
rect 216 1464 218 1478
rect 280 1477 282 1489
rect 290 1483 296 1484
rect 290 1479 291 1483
rect 295 1479 296 1483
rect 290 1478 296 1479
rect 278 1476 284 1477
rect 278 1472 279 1476
rect 283 1472 284 1476
rect 278 1471 284 1472
rect 110 1463 116 1464
rect 158 1463 164 1464
rect 158 1459 159 1463
rect 163 1459 164 1463
rect 158 1458 164 1459
rect 214 1463 220 1464
rect 214 1459 215 1463
rect 219 1459 220 1463
rect 214 1458 220 1459
rect 110 1451 116 1452
rect 110 1447 111 1451
rect 115 1447 116 1451
rect 110 1446 116 1447
rect 134 1448 140 1449
rect 112 1443 114 1446
rect 134 1444 135 1448
rect 139 1444 140 1448
rect 134 1443 140 1444
rect 111 1442 115 1443
rect 111 1437 115 1438
rect 135 1442 139 1443
rect 135 1437 139 1438
rect 112 1434 114 1437
rect 134 1436 140 1437
rect 110 1433 116 1434
rect 110 1429 111 1433
rect 115 1429 116 1433
rect 134 1432 135 1436
rect 139 1432 140 1436
rect 134 1431 140 1432
rect 110 1428 116 1429
rect 150 1419 156 1420
rect 110 1416 116 1417
rect 110 1412 111 1416
rect 115 1412 116 1416
rect 150 1415 151 1419
rect 155 1415 156 1419
rect 150 1414 156 1415
rect 110 1411 116 1412
rect 112 1391 114 1411
rect 134 1408 140 1409
rect 134 1404 135 1408
rect 139 1404 140 1408
rect 134 1403 140 1404
rect 136 1391 138 1403
rect 111 1390 115 1391
rect 111 1385 115 1386
rect 135 1390 139 1391
rect 135 1385 139 1386
rect 112 1365 114 1385
rect 136 1373 138 1385
rect 152 1380 154 1414
rect 160 1400 162 1458
rect 198 1448 204 1449
rect 198 1444 199 1448
rect 203 1444 204 1448
rect 198 1443 204 1444
rect 278 1448 284 1449
rect 278 1444 279 1448
rect 283 1444 284 1448
rect 278 1443 284 1444
rect 191 1442 195 1443
rect 191 1437 195 1438
rect 199 1442 203 1443
rect 199 1437 203 1438
rect 263 1442 267 1443
rect 263 1437 267 1438
rect 279 1442 283 1443
rect 279 1437 283 1438
rect 190 1436 196 1437
rect 190 1432 191 1436
rect 195 1432 196 1436
rect 190 1431 196 1432
rect 262 1436 268 1437
rect 262 1432 263 1436
rect 267 1432 268 1436
rect 262 1431 268 1432
rect 292 1420 294 1478
rect 360 1477 362 1489
rect 358 1476 364 1477
rect 358 1472 359 1476
rect 363 1472 364 1476
rect 358 1471 364 1472
rect 432 1464 434 1497
rect 480 1495 482 1507
rect 568 1495 570 1507
rect 656 1495 658 1507
rect 706 1503 712 1504
rect 706 1499 707 1503
rect 711 1499 712 1503
rect 706 1498 712 1499
rect 439 1494 443 1495
rect 439 1489 443 1490
rect 479 1494 483 1495
rect 479 1489 483 1490
rect 519 1494 523 1495
rect 519 1489 523 1490
rect 567 1494 571 1495
rect 567 1489 571 1490
rect 599 1494 603 1495
rect 599 1489 603 1490
rect 655 1494 659 1495
rect 655 1489 659 1490
rect 679 1494 683 1495
rect 679 1489 683 1490
rect 440 1477 442 1489
rect 520 1477 522 1489
rect 534 1483 540 1484
rect 534 1479 535 1483
rect 539 1479 540 1483
rect 534 1478 540 1479
rect 438 1476 444 1477
rect 438 1472 439 1476
rect 443 1472 444 1476
rect 438 1471 444 1472
rect 518 1476 524 1477
rect 518 1472 519 1476
rect 523 1472 524 1476
rect 518 1471 524 1472
rect 536 1464 538 1478
rect 600 1477 602 1489
rect 614 1483 620 1484
rect 614 1479 615 1483
rect 619 1479 620 1483
rect 614 1478 620 1479
rect 654 1483 660 1484
rect 654 1479 655 1483
rect 659 1479 660 1483
rect 654 1478 660 1479
rect 598 1476 604 1477
rect 598 1472 599 1476
rect 603 1472 604 1476
rect 598 1471 604 1472
rect 616 1464 618 1478
rect 430 1463 436 1464
rect 430 1459 431 1463
rect 435 1459 436 1463
rect 430 1458 436 1459
rect 446 1463 452 1464
rect 446 1459 447 1463
rect 451 1459 452 1463
rect 446 1458 452 1459
rect 534 1463 540 1464
rect 534 1459 535 1463
rect 539 1459 540 1463
rect 534 1458 540 1459
rect 614 1463 620 1464
rect 614 1459 615 1463
rect 619 1459 620 1463
rect 614 1458 620 1459
rect 358 1448 364 1449
rect 358 1444 359 1448
rect 363 1444 364 1448
rect 358 1443 364 1444
rect 438 1448 444 1449
rect 438 1444 439 1448
rect 443 1444 444 1448
rect 438 1443 444 1444
rect 335 1442 339 1443
rect 335 1437 339 1438
rect 359 1442 363 1443
rect 359 1437 363 1438
rect 407 1442 411 1443
rect 407 1437 411 1438
rect 439 1442 443 1443
rect 439 1437 443 1438
rect 334 1436 340 1437
rect 334 1432 335 1436
rect 339 1432 340 1436
rect 334 1431 340 1432
rect 406 1436 412 1437
rect 406 1432 407 1436
rect 411 1432 412 1436
rect 406 1431 412 1432
rect 278 1419 284 1420
rect 278 1415 279 1419
rect 283 1415 284 1419
rect 278 1414 284 1415
rect 290 1419 296 1420
rect 290 1415 291 1419
rect 295 1415 296 1419
rect 290 1414 296 1415
rect 358 1419 364 1420
rect 358 1415 359 1419
rect 363 1415 364 1419
rect 358 1414 364 1415
rect 190 1408 196 1409
rect 190 1404 191 1408
rect 195 1404 196 1408
rect 190 1403 196 1404
rect 262 1408 268 1409
rect 262 1404 263 1408
rect 267 1404 268 1408
rect 262 1403 268 1404
rect 158 1399 164 1400
rect 158 1395 159 1399
rect 163 1395 164 1399
rect 158 1394 164 1395
rect 192 1391 194 1403
rect 202 1399 208 1400
rect 202 1395 203 1399
rect 207 1395 208 1399
rect 202 1394 208 1395
rect 175 1390 179 1391
rect 175 1385 179 1386
rect 191 1390 195 1391
rect 191 1385 195 1386
rect 150 1379 156 1380
rect 150 1375 151 1379
rect 155 1375 156 1379
rect 150 1374 156 1375
rect 176 1373 178 1385
rect 134 1372 140 1373
rect 134 1368 135 1372
rect 139 1368 140 1372
rect 134 1367 140 1368
rect 174 1372 180 1373
rect 174 1368 175 1372
rect 179 1368 180 1372
rect 174 1367 180 1368
rect 110 1364 116 1365
rect 110 1360 111 1364
rect 115 1360 116 1364
rect 204 1360 206 1394
rect 264 1391 266 1403
rect 280 1400 282 1414
rect 334 1408 340 1409
rect 334 1404 335 1408
rect 339 1404 340 1408
rect 334 1403 340 1404
rect 278 1399 284 1400
rect 278 1395 279 1399
rect 283 1395 284 1399
rect 278 1394 284 1395
rect 336 1391 338 1403
rect 360 1392 362 1414
rect 406 1408 412 1409
rect 406 1404 407 1408
rect 411 1404 412 1408
rect 406 1403 412 1404
rect 358 1391 364 1392
rect 408 1391 410 1403
rect 448 1400 450 1458
rect 518 1448 524 1449
rect 518 1444 519 1448
rect 523 1444 524 1448
rect 518 1443 524 1444
rect 598 1448 604 1449
rect 598 1444 599 1448
rect 603 1444 604 1448
rect 598 1443 604 1444
rect 479 1442 483 1443
rect 479 1437 483 1438
rect 519 1442 523 1443
rect 519 1437 523 1438
rect 551 1442 555 1443
rect 551 1437 555 1438
rect 599 1442 603 1443
rect 599 1437 603 1438
rect 631 1442 635 1443
rect 631 1437 635 1438
rect 478 1436 484 1437
rect 478 1432 479 1436
rect 483 1432 484 1436
rect 478 1431 484 1432
rect 550 1436 556 1437
rect 550 1432 551 1436
rect 555 1432 556 1436
rect 550 1431 556 1432
rect 630 1436 636 1437
rect 630 1432 631 1436
rect 635 1432 636 1436
rect 630 1431 636 1432
rect 656 1420 658 1478
rect 680 1477 682 1489
rect 678 1476 684 1477
rect 678 1472 679 1476
rect 683 1472 684 1476
rect 678 1471 684 1472
rect 708 1464 710 1498
rect 744 1495 746 1507
rect 824 1495 826 1507
rect 852 1504 854 1562
rect 1135 1557 1139 1558
rect 1159 1562 1163 1563
rect 1159 1557 1163 1558
rect 1199 1562 1203 1563
rect 1199 1557 1203 1558
rect 1215 1562 1219 1563
rect 1215 1557 1219 1558
rect 1247 1562 1251 1563
rect 1247 1557 1251 1558
rect 1303 1562 1307 1563
rect 1303 1557 1307 1558
rect 1319 1562 1323 1563
rect 1319 1557 1323 1558
rect 1383 1562 1387 1563
rect 1383 1557 1387 1558
rect 1399 1562 1403 1563
rect 1399 1557 1403 1558
rect 1463 1562 1467 1563
rect 1463 1557 1467 1558
rect 1479 1562 1483 1563
rect 1479 1557 1483 1558
rect 1094 1555 1100 1556
rect 886 1552 892 1553
rect 886 1548 887 1552
rect 891 1548 892 1552
rect 1094 1551 1095 1555
rect 1099 1551 1100 1555
rect 1094 1550 1100 1551
rect 886 1547 892 1548
rect 1096 1547 1098 1550
rect 887 1546 891 1547
rect 887 1541 891 1542
rect 911 1546 915 1547
rect 911 1541 915 1542
rect 999 1546 1003 1547
rect 999 1541 1003 1542
rect 1095 1546 1099 1547
rect 1095 1541 1099 1542
rect 910 1540 916 1541
rect 910 1536 911 1540
rect 915 1536 916 1540
rect 910 1535 916 1536
rect 998 1540 1004 1541
rect 998 1536 999 1540
rect 1003 1536 1004 1540
rect 1096 1538 1098 1541
rect 998 1535 1004 1536
rect 1094 1537 1100 1538
rect 1136 1537 1138 1557
rect 1160 1545 1162 1557
rect 1200 1545 1202 1557
rect 1214 1551 1220 1552
rect 1214 1547 1215 1551
rect 1219 1547 1220 1551
rect 1214 1546 1220 1547
rect 1158 1544 1164 1545
rect 1158 1540 1159 1544
rect 1163 1540 1164 1544
rect 1158 1539 1164 1540
rect 1198 1544 1204 1545
rect 1198 1540 1199 1544
rect 1203 1540 1204 1544
rect 1198 1539 1204 1540
rect 1094 1533 1095 1537
rect 1099 1533 1100 1537
rect 1094 1532 1100 1533
rect 1134 1536 1140 1537
rect 1134 1532 1135 1536
rect 1139 1532 1140 1536
rect 1216 1532 1218 1546
rect 1248 1545 1250 1557
rect 1254 1551 1260 1552
rect 1254 1547 1255 1551
rect 1259 1547 1260 1551
rect 1254 1546 1260 1547
rect 1246 1544 1252 1545
rect 1246 1540 1247 1544
rect 1251 1540 1252 1544
rect 1246 1539 1252 1540
rect 1256 1532 1258 1546
rect 1320 1545 1322 1557
rect 1334 1551 1340 1552
rect 1334 1547 1335 1551
rect 1339 1547 1340 1551
rect 1334 1546 1340 1547
rect 1318 1544 1324 1545
rect 1318 1540 1319 1544
rect 1323 1540 1324 1544
rect 1318 1539 1324 1540
rect 1336 1532 1338 1546
rect 1400 1545 1402 1557
rect 1414 1551 1420 1552
rect 1414 1547 1415 1551
rect 1419 1547 1420 1551
rect 1414 1546 1420 1547
rect 1398 1544 1404 1545
rect 1398 1540 1399 1544
rect 1403 1540 1404 1544
rect 1398 1539 1404 1540
rect 1416 1532 1418 1546
rect 1480 1545 1482 1557
rect 1504 1552 1506 1578
rect 1542 1576 1543 1580
rect 1547 1576 1548 1580
rect 1542 1575 1548 1576
rect 1544 1563 1546 1575
rect 1616 1572 1618 1594
rect 1652 1592 1654 1662
rect 1696 1661 1698 1673
rect 1760 1661 1762 1673
rect 1774 1667 1780 1668
rect 1774 1663 1775 1667
rect 1779 1663 1780 1667
rect 1774 1662 1780 1663
rect 1694 1660 1700 1661
rect 1694 1656 1695 1660
rect 1699 1656 1700 1660
rect 1694 1655 1700 1656
rect 1758 1660 1764 1661
rect 1758 1656 1759 1660
rect 1763 1656 1764 1660
rect 1758 1655 1764 1656
rect 1776 1648 1778 1662
rect 1832 1661 1834 1673
rect 1846 1667 1852 1668
rect 1846 1663 1847 1667
rect 1851 1663 1852 1667
rect 1846 1662 1852 1663
rect 1830 1660 1836 1661
rect 1830 1656 1831 1660
rect 1835 1656 1836 1660
rect 1830 1655 1836 1656
rect 1848 1648 1850 1662
rect 1912 1661 1914 1673
rect 1936 1668 1938 1706
rect 1950 1700 1956 1701
rect 1950 1696 1951 1700
rect 1955 1696 1956 1700
rect 1950 1695 1956 1696
rect 2022 1700 2028 1701
rect 2022 1696 2023 1700
rect 2027 1696 2028 1700
rect 2022 1695 2028 1696
rect 1952 1679 1954 1695
rect 1986 1691 1992 1692
rect 1986 1687 1987 1691
rect 1991 1687 1992 1691
rect 1986 1686 1992 1687
rect 1951 1678 1955 1679
rect 1951 1673 1955 1674
rect 1926 1667 1932 1668
rect 1926 1663 1927 1667
rect 1931 1663 1932 1667
rect 1926 1662 1932 1663
rect 1934 1667 1940 1668
rect 1934 1663 1935 1667
rect 1939 1663 1940 1667
rect 1934 1662 1940 1663
rect 1910 1660 1916 1661
rect 1910 1656 1911 1660
rect 1915 1656 1916 1660
rect 1910 1655 1916 1656
rect 1928 1648 1930 1662
rect 1988 1648 1990 1686
rect 2024 1679 2026 1695
rect 1999 1678 2003 1679
rect 1999 1673 2003 1674
rect 2023 1678 2027 1679
rect 2023 1673 2027 1674
rect 2000 1661 2002 1673
rect 2048 1668 2050 1706
rect 2070 1700 2076 1701
rect 2070 1696 2071 1700
rect 2075 1696 2076 1700
rect 2070 1695 2076 1696
rect 2072 1679 2074 1695
rect 2096 1692 2098 1750
rect 2118 1743 2124 1744
rect 2118 1739 2119 1743
rect 2123 1739 2124 1743
rect 2118 1738 2124 1739
rect 2120 1735 2122 1738
rect 2119 1734 2123 1735
rect 2119 1729 2123 1730
rect 2120 1726 2122 1729
rect 2118 1725 2124 1726
rect 2118 1721 2119 1725
rect 2123 1721 2124 1725
rect 2118 1720 2124 1721
rect 2118 1708 2124 1709
rect 2118 1704 2119 1708
rect 2123 1704 2124 1708
rect 2118 1703 2124 1704
rect 2094 1691 2100 1692
rect 2094 1687 2095 1691
rect 2099 1687 2100 1691
rect 2094 1686 2100 1687
rect 2120 1679 2122 1703
rect 2071 1678 2075 1679
rect 2071 1673 2075 1674
rect 2119 1678 2123 1679
rect 2119 1673 2123 1674
rect 2010 1667 2016 1668
rect 2010 1663 2011 1667
rect 2015 1663 2016 1667
rect 2010 1662 2016 1663
rect 2046 1667 2052 1668
rect 2046 1663 2047 1667
rect 2051 1663 2052 1667
rect 2046 1662 2052 1663
rect 1998 1660 2004 1661
rect 1998 1656 1999 1660
rect 2003 1656 2004 1660
rect 1998 1655 2004 1656
rect 1734 1647 1740 1648
rect 1734 1643 1735 1647
rect 1739 1643 1740 1647
rect 1734 1642 1740 1643
rect 1774 1647 1780 1648
rect 1774 1643 1775 1647
rect 1779 1643 1780 1647
rect 1774 1642 1780 1643
rect 1846 1647 1852 1648
rect 1846 1643 1847 1647
rect 1851 1643 1852 1647
rect 1846 1642 1852 1643
rect 1926 1647 1932 1648
rect 1926 1643 1927 1647
rect 1931 1643 1932 1647
rect 1926 1642 1932 1643
rect 1986 1647 1992 1648
rect 1986 1643 1987 1647
rect 1991 1643 1992 1647
rect 1986 1642 1992 1643
rect 1694 1632 1700 1633
rect 1694 1628 1695 1632
rect 1699 1628 1700 1632
rect 1694 1627 1700 1628
rect 1696 1615 1698 1627
rect 1695 1614 1699 1615
rect 1695 1609 1699 1610
rect 1711 1614 1715 1615
rect 1711 1609 1715 1610
rect 1710 1608 1716 1609
rect 1710 1604 1711 1608
rect 1715 1604 1716 1608
rect 1710 1603 1716 1604
rect 1650 1591 1656 1592
rect 1650 1587 1651 1591
rect 1655 1587 1656 1591
rect 1650 1586 1656 1587
rect 1622 1580 1628 1581
rect 1622 1576 1623 1580
rect 1627 1576 1628 1580
rect 1622 1575 1628 1576
rect 1710 1580 1716 1581
rect 1710 1576 1711 1580
rect 1715 1576 1716 1580
rect 1710 1575 1716 1576
rect 1582 1571 1588 1572
rect 1582 1567 1583 1571
rect 1587 1567 1588 1571
rect 1582 1566 1588 1567
rect 1614 1571 1620 1572
rect 1614 1567 1615 1571
rect 1619 1567 1620 1571
rect 1614 1566 1620 1567
rect 1543 1562 1547 1563
rect 1543 1557 1547 1558
rect 1559 1562 1563 1563
rect 1559 1557 1563 1558
rect 1494 1551 1500 1552
rect 1494 1547 1495 1551
rect 1499 1547 1500 1551
rect 1494 1546 1500 1547
rect 1502 1551 1508 1552
rect 1502 1547 1503 1551
rect 1507 1547 1508 1551
rect 1502 1546 1508 1547
rect 1478 1544 1484 1545
rect 1478 1540 1479 1544
rect 1483 1540 1484 1544
rect 1478 1539 1484 1540
rect 1496 1532 1498 1546
rect 1560 1545 1562 1557
rect 1558 1544 1564 1545
rect 1558 1540 1559 1544
rect 1563 1540 1564 1544
rect 1558 1539 1564 1540
rect 1584 1532 1586 1566
rect 1624 1563 1626 1575
rect 1712 1563 1714 1575
rect 1736 1572 1738 1642
rect 1758 1632 1764 1633
rect 1758 1628 1759 1632
rect 1763 1628 1764 1632
rect 1758 1627 1764 1628
rect 1830 1632 1836 1633
rect 1830 1628 1831 1632
rect 1835 1628 1836 1632
rect 1830 1627 1836 1628
rect 1910 1632 1916 1633
rect 1910 1628 1911 1632
rect 1915 1628 1916 1632
rect 1910 1627 1916 1628
rect 1998 1632 2004 1633
rect 1998 1628 1999 1632
rect 2003 1628 2004 1632
rect 1998 1627 2004 1628
rect 1760 1615 1762 1627
rect 1832 1615 1834 1627
rect 1912 1615 1914 1627
rect 2000 1615 2002 1627
rect 1759 1614 1763 1615
rect 1759 1609 1763 1610
rect 1799 1614 1803 1615
rect 1799 1609 1803 1610
rect 1831 1614 1835 1615
rect 1831 1609 1835 1610
rect 1887 1614 1891 1615
rect 1887 1609 1891 1610
rect 1911 1614 1915 1615
rect 1911 1609 1915 1610
rect 1983 1614 1987 1615
rect 1983 1609 1987 1610
rect 1999 1614 2003 1615
rect 1999 1609 2003 1610
rect 1798 1608 1804 1609
rect 1798 1604 1799 1608
rect 1803 1604 1804 1608
rect 1798 1603 1804 1604
rect 1886 1608 1892 1609
rect 1886 1604 1887 1608
rect 1891 1604 1892 1608
rect 1886 1603 1892 1604
rect 1982 1608 1988 1609
rect 1982 1604 1983 1608
rect 1987 1604 1988 1608
rect 1982 1603 1988 1604
rect 2012 1592 2014 1662
rect 2072 1661 2074 1673
rect 2070 1660 2076 1661
rect 2070 1656 2071 1660
rect 2075 1656 2076 1660
rect 2070 1655 2076 1656
rect 2120 1653 2122 1673
rect 2118 1652 2124 1653
rect 2118 1648 2119 1652
rect 2123 1648 2124 1652
rect 2094 1647 2100 1648
rect 2118 1647 2124 1648
rect 2094 1643 2095 1647
rect 2099 1643 2100 1647
rect 2094 1642 2100 1643
rect 2070 1632 2076 1633
rect 2070 1628 2071 1632
rect 2075 1628 2076 1632
rect 2070 1627 2076 1628
rect 2072 1615 2074 1627
rect 2071 1614 2075 1615
rect 2071 1609 2075 1610
rect 2070 1608 2076 1609
rect 2070 1604 2071 1608
rect 2075 1604 2076 1608
rect 2070 1603 2076 1604
rect 1774 1591 1780 1592
rect 1774 1587 1775 1591
rect 1779 1587 1780 1591
rect 1774 1586 1780 1587
rect 1782 1591 1788 1592
rect 1782 1587 1783 1591
rect 1787 1587 1788 1591
rect 1782 1586 1788 1587
rect 2010 1591 2016 1592
rect 2010 1587 2011 1591
rect 2015 1587 2016 1591
rect 2010 1586 2016 1587
rect 1734 1571 1740 1572
rect 1734 1567 1735 1571
rect 1739 1567 1740 1571
rect 1734 1566 1740 1567
rect 1776 1564 1778 1586
rect 1774 1563 1780 1564
rect 1623 1562 1627 1563
rect 1623 1557 1627 1558
rect 1647 1562 1651 1563
rect 1647 1557 1651 1558
rect 1711 1562 1715 1563
rect 1711 1557 1715 1558
rect 1735 1562 1739 1563
rect 1774 1559 1775 1563
rect 1779 1559 1780 1563
rect 1774 1558 1780 1559
rect 1735 1557 1739 1558
rect 1648 1545 1650 1557
rect 1662 1551 1668 1552
rect 1662 1547 1663 1551
rect 1667 1547 1668 1551
rect 1662 1546 1668 1547
rect 1646 1544 1652 1545
rect 1646 1540 1647 1544
rect 1651 1540 1652 1544
rect 1646 1539 1652 1540
rect 1664 1532 1666 1546
rect 1736 1545 1738 1557
rect 1784 1552 1786 1586
rect 1798 1580 1804 1581
rect 1798 1576 1799 1580
rect 1803 1576 1804 1580
rect 1798 1575 1804 1576
rect 1886 1580 1892 1581
rect 1886 1576 1887 1580
rect 1891 1576 1892 1580
rect 1886 1575 1892 1576
rect 1982 1580 1988 1581
rect 1982 1576 1983 1580
rect 1987 1576 1988 1580
rect 1982 1575 1988 1576
rect 2070 1580 2076 1581
rect 2070 1576 2071 1580
rect 2075 1576 2076 1580
rect 2070 1575 2076 1576
rect 1800 1563 1802 1575
rect 1888 1563 1890 1575
rect 1946 1571 1952 1572
rect 1946 1567 1947 1571
rect 1951 1567 1952 1571
rect 1946 1566 1952 1567
rect 1799 1562 1803 1563
rect 1799 1557 1803 1558
rect 1823 1562 1827 1563
rect 1823 1557 1827 1558
rect 1887 1562 1891 1563
rect 1887 1557 1891 1558
rect 1911 1562 1915 1563
rect 1911 1557 1915 1558
rect 1750 1551 1756 1552
rect 1750 1547 1751 1551
rect 1755 1547 1756 1551
rect 1750 1546 1756 1547
rect 1782 1551 1788 1552
rect 1782 1547 1783 1551
rect 1787 1547 1788 1551
rect 1782 1546 1788 1547
rect 1798 1551 1804 1552
rect 1798 1547 1799 1551
rect 1803 1547 1804 1551
rect 1798 1546 1804 1547
rect 1734 1544 1740 1545
rect 1734 1540 1735 1544
rect 1739 1540 1740 1544
rect 1734 1539 1740 1540
rect 1752 1532 1754 1546
rect 1134 1531 1140 1532
rect 1182 1531 1188 1532
rect 1182 1527 1183 1531
rect 1187 1527 1188 1531
rect 1182 1526 1188 1527
rect 1214 1531 1220 1532
rect 1214 1527 1215 1531
rect 1219 1527 1220 1531
rect 1214 1526 1220 1527
rect 1254 1531 1260 1532
rect 1254 1527 1255 1531
rect 1259 1527 1260 1531
rect 1254 1526 1260 1527
rect 1334 1531 1340 1532
rect 1334 1527 1335 1531
rect 1339 1527 1340 1531
rect 1334 1526 1340 1527
rect 1414 1531 1420 1532
rect 1414 1527 1415 1531
rect 1419 1527 1420 1531
rect 1414 1526 1420 1527
rect 1494 1531 1500 1532
rect 1494 1527 1495 1531
rect 1499 1527 1500 1531
rect 1494 1526 1500 1527
rect 1582 1531 1588 1532
rect 1582 1527 1583 1531
rect 1587 1527 1588 1531
rect 1582 1526 1588 1527
rect 1662 1531 1668 1532
rect 1662 1527 1663 1531
rect 1667 1527 1668 1531
rect 1662 1526 1668 1527
rect 1750 1531 1756 1532
rect 1750 1527 1751 1531
rect 1755 1527 1756 1531
rect 1750 1526 1756 1527
rect 926 1523 932 1524
rect 926 1519 927 1523
rect 931 1519 932 1523
rect 926 1518 932 1519
rect 962 1523 968 1524
rect 962 1519 963 1523
rect 967 1519 968 1523
rect 962 1518 968 1519
rect 970 1523 976 1524
rect 970 1519 971 1523
rect 975 1519 976 1523
rect 970 1518 976 1519
rect 1094 1520 1100 1521
rect 910 1512 916 1513
rect 910 1508 911 1512
rect 915 1508 916 1512
rect 910 1507 916 1508
rect 850 1503 856 1504
rect 850 1499 851 1503
rect 855 1499 856 1503
rect 850 1498 856 1499
rect 912 1495 914 1507
rect 928 1504 930 1518
rect 964 1504 966 1518
rect 926 1503 932 1504
rect 926 1499 927 1503
rect 931 1499 932 1503
rect 926 1498 932 1499
rect 962 1503 968 1504
rect 962 1499 963 1503
rect 967 1499 968 1503
rect 962 1498 968 1499
rect 743 1494 747 1495
rect 743 1489 747 1490
rect 767 1494 771 1495
rect 767 1489 771 1490
rect 823 1494 827 1495
rect 823 1489 827 1490
rect 855 1494 859 1495
rect 855 1489 859 1490
rect 911 1494 915 1495
rect 911 1489 915 1490
rect 943 1494 947 1495
rect 943 1489 947 1490
rect 768 1477 770 1489
rect 782 1483 788 1484
rect 782 1479 783 1483
rect 787 1479 788 1483
rect 782 1478 788 1479
rect 818 1483 824 1484
rect 818 1479 819 1483
rect 823 1479 824 1483
rect 818 1478 824 1479
rect 826 1483 832 1484
rect 826 1479 827 1483
rect 831 1479 832 1483
rect 826 1478 832 1479
rect 766 1476 772 1477
rect 766 1472 767 1476
rect 771 1472 772 1476
rect 766 1471 772 1472
rect 784 1464 786 1478
rect 820 1464 822 1478
rect 706 1463 712 1464
rect 706 1459 707 1463
rect 711 1459 712 1463
rect 706 1458 712 1459
rect 782 1463 788 1464
rect 782 1459 783 1463
rect 787 1459 788 1463
rect 782 1458 788 1459
rect 818 1463 824 1464
rect 818 1459 819 1463
rect 823 1459 824 1463
rect 818 1458 824 1459
rect 678 1448 684 1449
rect 678 1444 679 1448
rect 683 1444 684 1448
rect 678 1443 684 1444
rect 766 1448 772 1449
rect 766 1444 767 1448
rect 771 1444 772 1448
rect 766 1443 772 1444
rect 679 1442 683 1443
rect 679 1437 683 1438
rect 711 1442 715 1443
rect 711 1437 715 1438
rect 767 1442 771 1443
rect 767 1437 771 1438
rect 799 1442 803 1443
rect 799 1437 803 1438
rect 710 1436 716 1437
rect 710 1432 711 1436
rect 715 1432 716 1436
rect 710 1431 716 1432
rect 798 1436 804 1437
rect 798 1432 799 1436
rect 803 1432 804 1436
rect 798 1431 804 1432
rect 828 1420 830 1478
rect 856 1477 858 1489
rect 944 1477 946 1489
rect 972 1484 974 1518
rect 1094 1516 1095 1520
rect 1099 1516 1100 1520
rect 1094 1515 1100 1516
rect 1134 1519 1140 1520
rect 1134 1515 1135 1519
rect 1139 1515 1140 1519
rect 998 1512 1004 1513
rect 998 1508 999 1512
rect 1003 1508 1004 1512
rect 998 1507 1004 1508
rect 1000 1495 1002 1507
rect 1096 1495 1098 1515
rect 1134 1514 1140 1515
rect 1158 1516 1164 1517
rect 1136 1511 1138 1514
rect 1158 1512 1159 1516
rect 1163 1512 1164 1516
rect 1158 1511 1164 1512
rect 1135 1510 1139 1511
rect 1135 1505 1139 1506
rect 1159 1510 1163 1511
rect 1159 1505 1163 1506
rect 1136 1502 1138 1505
rect 1158 1504 1164 1505
rect 1134 1501 1140 1502
rect 1134 1497 1135 1501
rect 1139 1497 1140 1501
rect 1158 1500 1159 1504
rect 1163 1500 1164 1504
rect 1158 1499 1164 1500
rect 1134 1496 1140 1497
rect 999 1494 1003 1495
rect 999 1489 1003 1490
rect 1031 1494 1035 1495
rect 1031 1489 1035 1490
rect 1095 1494 1099 1495
rect 1095 1489 1099 1490
rect 970 1483 976 1484
rect 970 1479 971 1483
rect 975 1479 976 1483
rect 970 1478 976 1479
rect 978 1483 984 1484
rect 978 1479 979 1483
rect 983 1479 984 1483
rect 978 1478 984 1479
rect 854 1476 860 1477
rect 854 1472 855 1476
rect 859 1472 860 1476
rect 854 1471 860 1472
rect 942 1476 948 1477
rect 942 1472 943 1476
rect 947 1472 948 1476
rect 942 1471 948 1472
rect 980 1464 982 1478
rect 1032 1477 1034 1489
rect 1030 1476 1036 1477
rect 1030 1472 1031 1476
rect 1035 1472 1036 1476
rect 1030 1471 1036 1472
rect 1096 1469 1098 1489
rect 1134 1484 1140 1485
rect 1134 1480 1135 1484
rect 1139 1480 1140 1484
rect 1134 1479 1140 1480
rect 1094 1468 1100 1469
rect 1094 1464 1095 1468
rect 1099 1464 1100 1468
rect 978 1463 984 1464
rect 978 1459 979 1463
rect 983 1459 984 1463
rect 978 1458 984 1459
rect 1070 1463 1076 1464
rect 1094 1463 1100 1464
rect 1070 1459 1071 1463
rect 1075 1459 1076 1463
rect 1070 1458 1076 1459
rect 854 1448 860 1449
rect 854 1444 855 1448
rect 859 1444 860 1448
rect 854 1443 860 1444
rect 942 1448 948 1449
rect 942 1444 943 1448
rect 947 1444 948 1448
rect 942 1443 948 1444
rect 1030 1448 1036 1449
rect 1030 1444 1031 1448
rect 1035 1444 1036 1448
rect 1030 1443 1036 1444
rect 855 1442 859 1443
rect 855 1437 859 1438
rect 887 1442 891 1443
rect 887 1437 891 1438
rect 943 1442 947 1443
rect 943 1437 947 1438
rect 975 1442 979 1443
rect 975 1437 979 1438
rect 1031 1442 1035 1443
rect 1031 1437 1035 1438
rect 1047 1442 1051 1443
rect 1047 1437 1051 1438
rect 886 1436 892 1437
rect 886 1432 887 1436
rect 891 1432 892 1436
rect 886 1431 892 1432
rect 974 1436 980 1437
rect 974 1432 975 1436
rect 979 1432 980 1436
rect 974 1431 980 1432
rect 1046 1436 1052 1437
rect 1046 1432 1047 1436
rect 1051 1432 1052 1436
rect 1046 1431 1052 1432
rect 526 1419 532 1420
rect 526 1415 527 1419
rect 531 1415 532 1419
rect 526 1414 532 1415
rect 654 1419 660 1420
rect 654 1415 655 1419
rect 659 1415 660 1419
rect 654 1414 660 1415
rect 826 1419 832 1420
rect 826 1415 827 1419
rect 831 1415 832 1419
rect 826 1414 832 1415
rect 834 1419 840 1420
rect 834 1415 835 1419
rect 839 1415 840 1419
rect 834 1414 840 1415
rect 1022 1419 1028 1420
rect 1022 1415 1023 1419
rect 1027 1415 1028 1419
rect 1022 1414 1028 1415
rect 1034 1419 1040 1420
rect 1034 1415 1035 1419
rect 1039 1415 1040 1419
rect 1034 1414 1040 1415
rect 478 1408 484 1409
rect 478 1404 479 1408
rect 483 1404 484 1408
rect 478 1403 484 1404
rect 446 1399 452 1400
rect 446 1395 447 1399
rect 451 1395 452 1399
rect 446 1394 452 1395
rect 480 1391 482 1403
rect 239 1390 243 1391
rect 239 1385 243 1386
rect 263 1390 267 1391
rect 263 1385 267 1386
rect 303 1390 307 1391
rect 303 1385 307 1386
rect 335 1390 339 1391
rect 358 1387 359 1391
rect 363 1387 364 1391
rect 358 1386 364 1387
rect 367 1390 371 1391
rect 335 1385 339 1386
rect 367 1385 371 1386
rect 407 1390 411 1391
rect 407 1385 411 1386
rect 439 1390 443 1391
rect 439 1385 443 1386
rect 479 1390 483 1391
rect 479 1385 483 1386
rect 503 1390 507 1391
rect 503 1385 507 1386
rect 240 1373 242 1385
rect 250 1379 256 1380
rect 250 1375 251 1379
rect 255 1375 256 1379
rect 250 1374 256 1375
rect 238 1372 244 1373
rect 238 1368 239 1372
rect 243 1368 244 1372
rect 238 1367 244 1368
rect 252 1360 254 1374
rect 304 1373 306 1385
rect 368 1373 370 1385
rect 382 1379 388 1380
rect 382 1375 383 1379
rect 387 1375 388 1379
rect 382 1374 388 1375
rect 302 1372 308 1373
rect 366 1372 372 1373
rect 302 1368 303 1372
rect 307 1368 308 1372
rect 302 1367 308 1368
rect 358 1371 364 1372
rect 358 1367 359 1371
rect 363 1367 364 1371
rect 366 1368 367 1372
rect 371 1368 372 1372
rect 366 1367 372 1368
rect 358 1366 364 1367
rect 110 1359 116 1360
rect 158 1359 164 1360
rect 158 1355 159 1359
rect 163 1355 164 1359
rect 158 1354 164 1355
rect 202 1359 208 1360
rect 202 1355 203 1359
rect 207 1355 208 1359
rect 202 1354 208 1355
rect 250 1359 256 1360
rect 250 1355 251 1359
rect 255 1355 256 1359
rect 250 1354 256 1355
rect 110 1347 116 1348
rect 110 1343 111 1347
rect 115 1343 116 1347
rect 110 1342 116 1343
rect 134 1344 140 1345
rect 112 1331 114 1342
rect 134 1340 135 1344
rect 139 1340 140 1344
rect 134 1339 140 1340
rect 136 1331 138 1339
rect 111 1330 115 1331
rect 111 1325 115 1326
rect 135 1330 139 1331
rect 135 1325 139 1326
rect 112 1322 114 1325
rect 134 1324 140 1325
rect 110 1321 116 1322
rect 110 1317 111 1321
rect 115 1317 116 1321
rect 134 1320 135 1324
rect 139 1320 140 1324
rect 134 1319 140 1320
rect 110 1316 116 1317
rect 110 1304 116 1305
rect 110 1300 111 1304
rect 115 1300 116 1304
rect 110 1299 116 1300
rect 112 1275 114 1299
rect 134 1296 140 1297
rect 134 1292 135 1296
rect 139 1292 140 1296
rect 134 1291 140 1292
rect 136 1275 138 1291
rect 160 1288 162 1354
rect 174 1344 180 1345
rect 174 1340 175 1344
rect 179 1340 180 1344
rect 174 1339 180 1340
rect 238 1344 244 1345
rect 238 1340 239 1344
rect 243 1340 244 1344
rect 238 1339 244 1340
rect 302 1344 308 1345
rect 302 1340 303 1344
rect 307 1340 308 1344
rect 302 1339 308 1340
rect 176 1331 178 1339
rect 240 1331 242 1339
rect 304 1331 306 1339
rect 175 1330 179 1331
rect 175 1325 179 1326
rect 215 1330 219 1331
rect 215 1325 219 1326
rect 239 1330 243 1331
rect 239 1325 243 1326
rect 255 1330 259 1331
rect 255 1325 259 1326
rect 303 1330 307 1331
rect 303 1325 307 1326
rect 319 1330 323 1331
rect 319 1325 323 1326
rect 174 1324 180 1325
rect 174 1320 175 1324
rect 179 1320 180 1324
rect 174 1319 180 1320
rect 214 1324 220 1325
rect 214 1320 215 1324
rect 219 1320 220 1324
rect 214 1319 220 1320
rect 254 1324 260 1325
rect 254 1320 255 1324
rect 259 1320 260 1324
rect 254 1319 260 1320
rect 318 1324 324 1325
rect 318 1320 319 1324
rect 323 1320 324 1324
rect 318 1319 324 1320
rect 342 1315 348 1316
rect 342 1311 343 1315
rect 347 1311 348 1315
rect 342 1310 348 1311
rect 190 1307 196 1308
rect 190 1303 191 1307
rect 195 1303 196 1307
rect 190 1302 196 1303
rect 230 1307 236 1308
rect 230 1303 231 1307
rect 235 1303 236 1307
rect 230 1302 236 1303
rect 278 1307 284 1308
rect 278 1303 279 1307
rect 283 1303 284 1307
rect 278 1302 284 1303
rect 174 1296 180 1297
rect 174 1292 175 1296
rect 179 1292 180 1296
rect 174 1291 180 1292
rect 158 1287 164 1288
rect 158 1283 159 1287
rect 163 1283 164 1287
rect 158 1282 164 1283
rect 176 1275 178 1291
rect 192 1288 194 1302
rect 214 1296 220 1297
rect 214 1292 215 1296
rect 219 1292 220 1296
rect 214 1291 220 1292
rect 190 1287 196 1288
rect 190 1283 191 1287
rect 195 1283 196 1287
rect 190 1282 196 1283
rect 216 1275 218 1291
rect 232 1288 234 1302
rect 254 1296 260 1297
rect 254 1292 255 1296
rect 259 1292 260 1296
rect 254 1291 260 1292
rect 230 1287 236 1288
rect 230 1283 231 1287
rect 235 1283 236 1287
rect 230 1282 236 1283
rect 256 1275 258 1291
rect 111 1274 115 1275
rect 111 1269 115 1270
rect 135 1274 139 1275
rect 135 1269 139 1270
rect 175 1274 179 1275
rect 175 1269 179 1270
rect 215 1274 219 1275
rect 215 1269 219 1270
rect 255 1274 259 1275
rect 280 1272 282 1302
rect 318 1296 324 1297
rect 318 1292 319 1296
rect 323 1292 324 1296
rect 318 1291 324 1292
rect 320 1275 322 1291
rect 344 1288 346 1310
rect 360 1308 362 1366
rect 384 1360 386 1374
rect 440 1373 442 1385
rect 454 1379 460 1380
rect 454 1375 455 1379
rect 459 1375 460 1379
rect 454 1374 460 1375
rect 438 1372 444 1373
rect 438 1368 439 1372
rect 443 1368 444 1372
rect 438 1367 444 1368
rect 456 1360 458 1374
rect 504 1373 506 1385
rect 528 1380 530 1414
rect 550 1408 556 1409
rect 550 1404 551 1408
rect 555 1404 556 1408
rect 550 1403 556 1404
rect 630 1408 636 1409
rect 630 1404 631 1408
rect 635 1404 636 1408
rect 630 1403 636 1404
rect 710 1408 716 1409
rect 710 1404 711 1408
rect 715 1404 716 1408
rect 710 1403 716 1404
rect 798 1408 804 1409
rect 798 1404 799 1408
rect 803 1404 804 1408
rect 798 1403 804 1404
rect 552 1391 554 1403
rect 598 1399 604 1400
rect 598 1395 599 1399
rect 603 1395 604 1399
rect 598 1394 604 1395
rect 551 1390 555 1391
rect 551 1385 555 1386
rect 575 1390 579 1391
rect 575 1385 579 1386
rect 510 1379 516 1380
rect 510 1375 511 1379
rect 515 1375 516 1379
rect 510 1374 516 1375
rect 526 1379 532 1380
rect 526 1375 527 1379
rect 531 1375 532 1379
rect 526 1374 532 1375
rect 502 1372 508 1373
rect 502 1368 503 1372
rect 507 1368 508 1372
rect 502 1367 508 1368
rect 512 1360 514 1374
rect 576 1373 578 1385
rect 574 1372 580 1373
rect 574 1368 575 1372
rect 579 1368 580 1372
rect 574 1367 580 1368
rect 600 1360 602 1394
rect 632 1391 634 1403
rect 712 1391 714 1403
rect 800 1391 802 1403
rect 836 1400 838 1414
rect 886 1408 892 1409
rect 886 1404 887 1408
rect 891 1404 892 1408
rect 886 1403 892 1404
rect 974 1408 980 1409
rect 974 1404 975 1408
rect 979 1404 980 1408
rect 974 1403 980 1404
rect 834 1399 840 1400
rect 834 1395 835 1399
rect 839 1395 840 1399
rect 834 1394 840 1395
rect 888 1391 890 1403
rect 950 1399 956 1400
rect 950 1395 951 1399
rect 955 1395 956 1399
rect 950 1394 956 1395
rect 631 1390 635 1391
rect 631 1385 635 1386
rect 647 1390 651 1391
rect 647 1385 651 1386
rect 711 1390 715 1391
rect 711 1385 715 1386
rect 783 1390 787 1391
rect 783 1385 787 1386
rect 799 1390 803 1391
rect 799 1385 803 1386
rect 855 1390 859 1391
rect 855 1385 859 1386
rect 887 1390 891 1391
rect 887 1385 891 1386
rect 927 1390 931 1391
rect 927 1385 931 1386
rect 648 1373 650 1385
rect 662 1379 668 1380
rect 662 1375 663 1379
rect 667 1375 668 1379
rect 662 1374 668 1375
rect 646 1372 652 1373
rect 646 1368 647 1372
rect 651 1368 652 1372
rect 646 1367 652 1368
rect 664 1360 666 1374
rect 712 1373 714 1385
rect 718 1379 724 1380
rect 718 1375 719 1379
rect 723 1375 724 1379
rect 718 1374 724 1375
rect 730 1379 736 1380
rect 730 1375 731 1379
rect 735 1375 736 1379
rect 730 1374 736 1375
rect 710 1372 716 1373
rect 710 1368 711 1372
rect 715 1368 716 1372
rect 710 1367 716 1368
rect 720 1360 722 1374
rect 374 1359 380 1360
rect 374 1355 375 1359
rect 379 1355 380 1359
rect 374 1354 380 1355
rect 382 1359 388 1360
rect 382 1355 383 1359
rect 387 1355 388 1359
rect 382 1354 388 1355
rect 454 1359 460 1360
rect 454 1355 455 1359
rect 459 1355 460 1359
rect 454 1354 460 1355
rect 510 1359 516 1360
rect 510 1355 511 1359
rect 515 1355 516 1359
rect 510 1354 516 1355
rect 598 1359 604 1360
rect 598 1355 599 1359
rect 603 1355 604 1359
rect 598 1354 604 1355
rect 662 1359 668 1360
rect 662 1355 663 1359
rect 667 1355 668 1359
rect 662 1354 668 1355
rect 718 1359 724 1360
rect 718 1355 719 1359
rect 723 1355 724 1359
rect 718 1354 724 1355
rect 366 1344 372 1345
rect 366 1340 367 1344
rect 371 1340 372 1344
rect 366 1339 372 1340
rect 368 1331 370 1339
rect 367 1330 371 1331
rect 367 1325 371 1326
rect 358 1307 364 1308
rect 358 1303 359 1307
rect 363 1303 364 1307
rect 358 1302 364 1303
rect 342 1287 348 1288
rect 342 1283 343 1287
rect 347 1283 348 1287
rect 342 1282 348 1283
rect 376 1280 378 1354
rect 438 1344 444 1345
rect 438 1340 439 1344
rect 443 1340 444 1344
rect 438 1339 444 1340
rect 502 1344 508 1345
rect 502 1340 503 1344
rect 507 1340 508 1344
rect 502 1339 508 1340
rect 574 1344 580 1345
rect 574 1340 575 1344
rect 579 1340 580 1344
rect 574 1339 580 1340
rect 646 1344 652 1345
rect 646 1340 647 1344
rect 651 1340 652 1344
rect 646 1339 652 1340
rect 710 1344 716 1345
rect 710 1340 711 1344
rect 715 1340 716 1344
rect 710 1339 716 1340
rect 440 1331 442 1339
rect 504 1331 506 1339
rect 576 1331 578 1339
rect 648 1331 650 1339
rect 712 1331 714 1339
rect 391 1330 395 1331
rect 391 1325 395 1326
rect 439 1330 443 1331
rect 439 1325 443 1326
rect 463 1330 467 1331
rect 463 1325 467 1326
rect 503 1330 507 1331
rect 503 1325 507 1326
rect 543 1330 547 1331
rect 543 1325 547 1326
rect 575 1330 579 1331
rect 575 1325 579 1326
rect 623 1330 627 1331
rect 623 1325 627 1326
rect 647 1330 651 1331
rect 647 1325 651 1326
rect 703 1330 707 1331
rect 703 1325 707 1326
rect 711 1330 715 1331
rect 711 1325 715 1326
rect 390 1324 396 1325
rect 390 1320 391 1324
rect 395 1320 396 1324
rect 390 1319 396 1320
rect 462 1324 468 1325
rect 462 1320 463 1324
rect 467 1320 468 1324
rect 462 1319 468 1320
rect 542 1324 548 1325
rect 542 1320 543 1324
rect 547 1320 548 1324
rect 542 1319 548 1320
rect 622 1324 628 1325
rect 622 1320 623 1324
rect 627 1320 628 1324
rect 622 1319 628 1320
rect 702 1324 708 1325
rect 702 1320 703 1324
rect 707 1320 708 1324
rect 702 1319 708 1320
rect 732 1308 734 1374
rect 784 1373 786 1385
rect 806 1379 812 1380
rect 806 1375 807 1379
rect 811 1375 812 1379
rect 806 1374 812 1375
rect 782 1372 788 1373
rect 782 1368 783 1372
rect 787 1368 788 1372
rect 782 1367 788 1368
rect 782 1344 788 1345
rect 782 1340 783 1344
rect 787 1340 788 1344
rect 782 1339 788 1340
rect 784 1331 786 1339
rect 783 1330 787 1331
rect 783 1325 787 1326
rect 782 1324 788 1325
rect 782 1320 783 1324
rect 787 1320 788 1324
rect 782 1319 788 1320
rect 808 1308 810 1374
rect 856 1373 858 1385
rect 890 1379 896 1380
rect 890 1375 891 1379
rect 895 1375 896 1379
rect 890 1374 896 1375
rect 854 1372 860 1373
rect 854 1368 855 1372
rect 859 1368 860 1372
rect 854 1367 860 1368
rect 892 1360 894 1374
rect 928 1373 930 1385
rect 926 1372 932 1373
rect 926 1368 927 1372
rect 931 1368 932 1372
rect 926 1367 932 1368
rect 952 1360 954 1394
rect 976 1391 978 1403
rect 975 1390 979 1391
rect 975 1385 979 1386
rect 999 1390 1003 1391
rect 999 1385 1003 1386
rect 1000 1373 1002 1385
rect 1024 1380 1026 1414
rect 1036 1400 1038 1414
rect 1046 1408 1052 1409
rect 1046 1404 1047 1408
rect 1051 1404 1052 1408
rect 1046 1403 1052 1404
rect 1034 1399 1040 1400
rect 1034 1395 1035 1399
rect 1039 1395 1040 1399
rect 1034 1394 1040 1395
rect 1048 1391 1050 1403
rect 1072 1400 1074 1458
rect 1136 1455 1138 1479
rect 1158 1476 1164 1477
rect 1158 1472 1159 1476
rect 1163 1472 1164 1476
rect 1158 1471 1164 1472
rect 1160 1455 1162 1471
rect 1184 1468 1186 1526
rect 1198 1516 1204 1517
rect 1198 1512 1199 1516
rect 1203 1512 1204 1516
rect 1198 1511 1204 1512
rect 1246 1516 1252 1517
rect 1246 1512 1247 1516
rect 1251 1512 1252 1516
rect 1246 1511 1252 1512
rect 1318 1516 1324 1517
rect 1318 1512 1319 1516
rect 1323 1512 1324 1516
rect 1318 1511 1324 1512
rect 1398 1516 1404 1517
rect 1398 1512 1399 1516
rect 1403 1512 1404 1516
rect 1398 1511 1404 1512
rect 1478 1516 1484 1517
rect 1478 1512 1479 1516
rect 1483 1512 1484 1516
rect 1478 1511 1484 1512
rect 1558 1516 1564 1517
rect 1558 1512 1559 1516
rect 1563 1512 1564 1516
rect 1558 1511 1564 1512
rect 1646 1516 1652 1517
rect 1646 1512 1647 1516
rect 1651 1512 1652 1516
rect 1646 1511 1652 1512
rect 1734 1516 1740 1517
rect 1734 1512 1735 1516
rect 1739 1512 1740 1516
rect 1734 1511 1740 1512
rect 1199 1510 1203 1511
rect 1199 1505 1203 1506
rect 1239 1510 1243 1511
rect 1239 1505 1243 1506
rect 1247 1510 1251 1511
rect 1247 1505 1251 1506
rect 1303 1510 1307 1511
rect 1303 1505 1307 1506
rect 1319 1510 1323 1511
rect 1319 1505 1323 1506
rect 1375 1510 1379 1511
rect 1375 1505 1379 1506
rect 1399 1510 1403 1511
rect 1399 1505 1403 1506
rect 1455 1510 1459 1511
rect 1455 1505 1459 1506
rect 1479 1510 1483 1511
rect 1479 1505 1483 1506
rect 1543 1510 1547 1511
rect 1543 1505 1547 1506
rect 1559 1510 1563 1511
rect 1559 1505 1563 1506
rect 1623 1510 1627 1511
rect 1623 1505 1627 1506
rect 1647 1510 1651 1511
rect 1647 1505 1651 1506
rect 1703 1510 1707 1511
rect 1703 1505 1707 1506
rect 1735 1510 1739 1511
rect 1735 1505 1739 1506
rect 1775 1510 1779 1511
rect 1775 1505 1779 1506
rect 1198 1504 1204 1505
rect 1198 1500 1199 1504
rect 1203 1500 1204 1504
rect 1198 1499 1204 1500
rect 1238 1504 1244 1505
rect 1238 1500 1239 1504
rect 1243 1500 1244 1504
rect 1238 1499 1244 1500
rect 1302 1504 1308 1505
rect 1302 1500 1303 1504
rect 1307 1500 1308 1504
rect 1302 1499 1308 1500
rect 1374 1504 1380 1505
rect 1374 1500 1375 1504
rect 1379 1500 1380 1504
rect 1374 1499 1380 1500
rect 1454 1504 1460 1505
rect 1454 1500 1455 1504
rect 1459 1500 1460 1504
rect 1454 1499 1460 1500
rect 1542 1504 1548 1505
rect 1542 1500 1543 1504
rect 1547 1500 1548 1504
rect 1542 1499 1548 1500
rect 1622 1504 1628 1505
rect 1622 1500 1623 1504
rect 1627 1500 1628 1504
rect 1622 1499 1628 1500
rect 1702 1504 1708 1505
rect 1702 1500 1703 1504
rect 1707 1500 1708 1504
rect 1702 1499 1708 1500
rect 1774 1504 1780 1505
rect 1774 1500 1775 1504
rect 1779 1500 1780 1504
rect 1774 1499 1780 1500
rect 1800 1496 1802 1546
rect 1824 1545 1826 1557
rect 1912 1545 1914 1557
rect 1822 1544 1828 1545
rect 1822 1540 1823 1544
rect 1827 1540 1828 1544
rect 1822 1539 1828 1540
rect 1910 1544 1916 1545
rect 1910 1540 1911 1544
rect 1915 1540 1916 1544
rect 1910 1539 1916 1540
rect 1822 1516 1828 1517
rect 1822 1512 1823 1516
rect 1827 1512 1828 1516
rect 1822 1511 1828 1512
rect 1910 1516 1916 1517
rect 1910 1512 1911 1516
rect 1915 1512 1916 1516
rect 1910 1511 1916 1512
rect 1823 1510 1827 1511
rect 1823 1505 1827 1506
rect 1847 1510 1851 1511
rect 1847 1505 1851 1506
rect 1911 1510 1915 1511
rect 1911 1505 1915 1506
rect 1919 1510 1923 1511
rect 1919 1505 1923 1506
rect 1846 1504 1852 1505
rect 1846 1500 1847 1504
rect 1851 1500 1852 1504
rect 1846 1499 1852 1500
rect 1918 1504 1924 1505
rect 1918 1500 1919 1504
rect 1923 1500 1924 1504
rect 1918 1499 1924 1500
rect 1798 1495 1804 1496
rect 1798 1491 1799 1495
rect 1803 1491 1804 1495
rect 1798 1490 1804 1491
rect 1948 1488 1950 1566
rect 1984 1563 1986 1575
rect 2072 1563 2074 1575
rect 2096 1572 2098 1642
rect 2118 1635 2124 1636
rect 2118 1631 2119 1635
rect 2123 1631 2124 1635
rect 2118 1630 2124 1631
rect 2120 1615 2122 1630
rect 2119 1614 2123 1615
rect 2119 1609 2123 1610
rect 2120 1606 2122 1609
rect 2118 1605 2124 1606
rect 2118 1601 2119 1605
rect 2123 1601 2124 1605
rect 2118 1600 2124 1601
rect 2118 1588 2124 1589
rect 2118 1584 2119 1588
rect 2123 1584 2124 1588
rect 2118 1583 2124 1584
rect 2094 1571 2100 1572
rect 2094 1567 2095 1571
rect 2099 1567 2100 1571
rect 2094 1566 2100 1567
rect 2120 1563 2122 1583
rect 1983 1562 1987 1563
rect 1983 1557 1987 1558
rect 1999 1562 2003 1563
rect 1999 1557 2003 1558
rect 2071 1562 2075 1563
rect 2071 1557 2075 1558
rect 2119 1562 2123 1563
rect 2119 1557 2123 1558
rect 2000 1545 2002 1557
rect 2072 1545 2074 1557
rect 1998 1544 2004 1545
rect 1998 1540 1999 1544
rect 2003 1540 2004 1544
rect 1998 1539 2004 1540
rect 2070 1544 2076 1545
rect 2070 1540 2071 1544
rect 2075 1540 2076 1544
rect 2070 1539 2076 1540
rect 2120 1537 2122 1557
rect 2118 1536 2124 1537
rect 2118 1532 2119 1536
rect 2123 1532 2124 1536
rect 2018 1531 2024 1532
rect 2018 1527 2019 1531
rect 2023 1527 2024 1531
rect 2018 1526 2024 1527
rect 2038 1531 2044 1532
rect 2118 1531 2124 1532
rect 2038 1527 2039 1531
rect 2043 1527 2044 1531
rect 2038 1526 2044 1527
rect 1998 1516 2004 1517
rect 1998 1512 1999 1516
rect 2003 1512 2004 1516
rect 1998 1511 2004 1512
rect 1991 1510 1995 1511
rect 1991 1505 1995 1506
rect 1999 1510 2003 1511
rect 1999 1505 2003 1506
rect 1990 1504 1996 1505
rect 1990 1500 1991 1504
rect 1995 1500 1996 1504
rect 1990 1499 1996 1500
rect 1214 1487 1220 1488
rect 1214 1483 1215 1487
rect 1219 1483 1220 1487
rect 1214 1482 1220 1483
rect 1254 1487 1260 1488
rect 1254 1483 1255 1487
rect 1259 1483 1260 1487
rect 1254 1482 1260 1483
rect 1318 1487 1324 1488
rect 1318 1483 1319 1487
rect 1323 1483 1324 1487
rect 1318 1482 1324 1483
rect 1390 1487 1396 1488
rect 1390 1483 1391 1487
rect 1395 1483 1396 1487
rect 1390 1482 1396 1483
rect 1470 1487 1476 1488
rect 1470 1483 1471 1487
rect 1475 1483 1476 1487
rect 1470 1482 1476 1483
rect 1534 1487 1540 1488
rect 1534 1483 1535 1487
rect 1539 1483 1540 1487
rect 1534 1482 1540 1483
rect 1946 1487 1952 1488
rect 1946 1483 1947 1487
rect 1951 1483 1952 1487
rect 1946 1482 1952 1483
rect 1198 1476 1204 1477
rect 1198 1472 1199 1476
rect 1203 1472 1204 1476
rect 1198 1471 1204 1472
rect 1182 1467 1188 1468
rect 1182 1463 1183 1467
rect 1187 1463 1188 1467
rect 1182 1462 1188 1463
rect 1200 1455 1202 1471
rect 1216 1468 1218 1482
rect 1238 1476 1244 1477
rect 1238 1472 1239 1476
rect 1243 1472 1244 1476
rect 1238 1471 1244 1472
rect 1214 1467 1220 1468
rect 1214 1463 1215 1467
rect 1219 1463 1220 1467
rect 1214 1462 1220 1463
rect 1240 1455 1242 1471
rect 1256 1468 1258 1482
rect 1302 1476 1308 1477
rect 1302 1472 1303 1476
rect 1307 1472 1308 1476
rect 1302 1471 1308 1472
rect 1254 1467 1260 1468
rect 1254 1463 1255 1467
rect 1259 1463 1260 1467
rect 1254 1462 1260 1463
rect 1304 1455 1306 1471
rect 1320 1468 1322 1482
rect 1374 1476 1380 1477
rect 1374 1472 1375 1476
rect 1379 1472 1380 1476
rect 1374 1471 1380 1472
rect 1318 1467 1324 1468
rect 1318 1463 1319 1467
rect 1323 1463 1324 1467
rect 1318 1462 1324 1463
rect 1376 1455 1378 1471
rect 1392 1468 1394 1482
rect 1454 1476 1460 1477
rect 1454 1472 1455 1476
rect 1459 1472 1460 1476
rect 1454 1471 1460 1472
rect 1390 1467 1396 1468
rect 1390 1463 1391 1467
rect 1395 1463 1396 1467
rect 1390 1462 1396 1463
rect 1456 1455 1458 1471
rect 1472 1468 1474 1482
rect 1470 1467 1476 1468
rect 1470 1463 1471 1467
rect 1475 1463 1476 1467
rect 1470 1462 1476 1463
rect 1135 1454 1139 1455
rect 1094 1451 1100 1452
rect 1094 1447 1095 1451
rect 1099 1447 1100 1451
rect 1135 1449 1139 1450
rect 1159 1454 1163 1455
rect 1159 1449 1163 1450
rect 1199 1454 1203 1455
rect 1199 1449 1203 1450
rect 1239 1454 1243 1455
rect 1239 1449 1243 1450
rect 1279 1454 1283 1455
rect 1279 1449 1283 1450
rect 1303 1454 1307 1455
rect 1303 1449 1307 1450
rect 1327 1454 1331 1455
rect 1327 1449 1331 1450
rect 1375 1454 1379 1455
rect 1375 1449 1379 1450
rect 1383 1454 1387 1455
rect 1383 1449 1387 1450
rect 1439 1454 1443 1455
rect 1439 1449 1443 1450
rect 1455 1454 1459 1455
rect 1455 1449 1459 1450
rect 1495 1454 1499 1455
rect 1495 1449 1499 1450
rect 1094 1446 1100 1447
rect 1096 1443 1098 1446
rect 1095 1442 1099 1443
rect 1095 1437 1099 1438
rect 1096 1434 1098 1437
rect 1094 1433 1100 1434
rect 1094 1429 1095 1433
rect 1099 1429 1100 1433
rect 1136 1429 1138 1449
rect 1280 1437 1282 1449
rect 1328 1437 1330 1449
rect 1342 1443 1348 1444
rect 1342 1439 1343 1443
rect 1347 1439 1348 1443
rect 1342 1438 1348 1439
rect 1278 1436 1284 1437
rect 1278 1432 1279 1436
rect 1283 1432 1284 1436
rect 1278 1431 1284 1432
rect 1326 1436 1332 1437
rect 1326 1432 1327 1436
rect 1331 1432 1332 1436
rect 1326 1431 1332 1432
rect 1094 1428 1100 1429
rect 1134 1428 1140 1429
rect 1134 1424 1135 1428
rect 1139 1424 1140 1428
rect 1344 1424 1346 1438
rect 1384 1437 1386 1449
rect 1398 1443 1404 1444
rect 1398 1439 1399 1443
rect 1403 1439 1404 1443
rect 1398 1438 1404 1439
rect 1382 1436 1388 1437
rect 1382 1432 1383 1436
rect 1387 1432 1388 1436
rect 1382 1431 1388 1432
rect 1400 1424 1402 1438
rect 1440 1437 1442 1449
rect 1446 1443 1452 1444
rect 1446 1439 1447 1443
rect 1451 1439 1452 1443
rect 1446 1438 1452 1439
rect 1438 1436 1444 1437
rect 1438 1432 1439 1436
rect 1443 1432 1444 1436
rect 1438 1431 1444 1432
rect 1448 1424 1450 1438
rect 1496 1437 1498 1449
rect 1536 1444 1538 1482
rect 1542 1476 1548 1477
rect 1542 1472 1543 1476
rect 1547 1472 1548 1476
rect 1542 1471 1548 1472
rect 1622 1476 1628 1477
rect 1622 1472 1623 1476
rect 1627 1472 1628 1476
rect 1622 1471 1628 1472
rect 1702 1476 1708 1477
rect 1702 1472 1703 1476
rect 1707 1472 1708 1476
rect 1702 1471 1708 1472
rect 1774 1476 1780 1477
rect 1774 1472 1775 1476
rect 1779 1472 1780 1476
rect 1774 1471 1780 1472
rect 1846 1476 1852 1477
rect 1846 1472 1847 1476
rect 1851 1472 1852 1476
rect 1846 1471 1852 1472
rect 1918 1476 1924 1477
rect 1918 1472 1919 1476
rect 1923 1472 1924 1476
rect 1918 1471 1924 1472
rect 1990 1476 1996 1477
rect 1990 1472 1991 1476
rect 1995 1472 1996 1476
rect 1990 1471 1996 1472
rect 1544 1455 1546 1471
rect 1624 1455 1626 1471
rect 1704 1455 1706 1471
rect 1776 1455 1778 1471
rect 1848 1455 1850 1471
rect 1910 1467 1916 1468
rect 1910 1463 1911 1467
rect 1915 1463 1916 1467
rect 1910 1462 1916 1463
rect 1543 1454 1547 1455
rect 1543 1449 1547 1450
rect 1551 1454 1555 1455
rect 1607 1454 1611 1455
rect 1551 1449 1555 1450
rect 1578 1451 1584 1452
rect 1510 1443 1516 1444
rect 1510 1439 1511 1443
rect 1515 1439 1516 1443
rect 1510 1438 1516 1439
rect 1534 1443 1540 1444
rect 1534 1439 1535 1443
rect 1539 1439 1540 1443
rect 1534 1438 1540 1439
rect 1494 1436 1500 1437
rect 1494 1432 1495 1436
rect 1499 1432 1500 1436
rect 1494 1431 1500 1432
rect 1512 1424 1514 1438
rect 1552 1437 1554 1449
rect 1578 1447 1579 1451
rect 1583 1447 1584 1451
rect 1607 1449 1611 1450
rect 1623 1454 1627 1455
rect 1623 1449 1627 1450
rect 1671 1454 1675 1455
rect 1671 1449 1675 1450
rect 1703 1454 1707 1455
rect 1703 1449 1707 1450
rect 1735 1454 1739 1455
rect 1735 1449 1739 1450
rect 1775 1454 1779 1455
rect 1775 1449 1779 1450
rect 1807 1454 1811 1455
rect 1807 1449 1811 1450
rect 1847 1454 1851 1455
rect 1847 1449 1851 1450
rect 1887 1454 1891 1455
rect 1887 1449 1891 1450
rect 1578 1446 1584 1447
rect 1550 1436 1556 1437
rect 1550 1432 1551 1436
rect 1555 1432 1556 1436
rect 1550 1431 1556 1432
rect 1580 1424 1582 1446
rect 1608 1437 1610 1449
rect 1614 1443 1620 1444
rect 1614 1439 1615 1443
rect 1619 1439 1620 1443
rect 1614 1438 1620 1439
rect 1606 1436 1612 1437
rect 1606 1432 1607 1436
rect 1611 1432 1612 1436
rect 1606 1431 1612 1432
rect 1616 1424 1618 1438
rect 1672 1437 1674 1449
rect 1686 1443 1692 1444
rect 1686 1439 1687 1443
rect 1691 1439 1692 1443
rect 1686 1438 1692 1439
rect 1670 1436 1676 1437
rect 1670 1432 1671 1436
rect 1675 1432 1676 1436
rect 1670 1431 1676 1432
rect 1688 1424 1690 1438
rect 1736 1437 1738 1449
rect 1742 1443 1748 1444
rect 1742 1439 1743 1443
rect 1747 1439 1748 1443
rect 1742 1438 1748 1439
rect 1734 1436 1740 1437
rect 1734 1432 1735 1436
rect 1739 1432 1740 1436
rect 1734 1431 1740 1432
rect 1134 1423 1140 1424
rect 1342 1423 1348 1424
rect 1342 1419 1343 1423
rect 1347 1419 1348 1423
rect 1342 1418 1348 1419
rect 1398 1423 1404 1424
rect 1398 1419 1399 1423
rect 1403 1419 1404 1423
rect 1398 1418 1404 1419
rect 1446 1423 1452 1424
rect 1446 1419 1447 1423
rect 1451 1419 1452 1423
rect 1446 1418 1452 1419
rect 1510 1423 1516 1424
rect 1510 1419 1511 1423
rect 1515 1419 1516 1423
rect 1510 1418 1516 1419
rect 1578 1423 1584 1424
rect 1578 1419 1579 1423
rect 1583 1419 1584 1423
rect 1578 1418 1584 1419
rect 1614 1423 1620 1424
rect 1614 1419 1615 1423
rect 1619 1419 1620 1423
rect 1614 1418 1620 1419
rect 1686 1423 1692 1424
rect 1686 1419 1687 1423
rect 1691 1419 1692 1423
rect 1686 1418 1692 1419
rect 1094 1416 1100 1417
rect 1094 1412 1095 1416
rect 1099 1412 1100 1416
rect 1094 1411 1100 1412
rect 1134 1411 1140 1412
rect 1070 1399 1076 1400
rect 1070 1395 1071 1399
rect 1075 1395 1076 1399
rect 1070 1394 1076 1395
rect 1096 1391 1098 1411
rect 1134 1407 1135 1411
rect 1139 1407 1140 1411
rect 1134 1406 1140 1407
rect 1278 1408 1284 1409
rect 1136 1399 1138 1406
rect 1278 1404 1279 1408
rect 1283 1404 1284 1408
rect 1278 1403 1284 1404
rect 1326 1408 1332 1409
rect 1326 1404 1327 1408
rect 1331 1404 1332 1408
rect 1326 1403 1332 1404
rect 1382 1408 1388 1409
rect 1382 1404 1383 1408
rect 1387 1404 1388 1408
rect 1382 1403 1388 1404
rect 1438 1408 1444 1409
rect 1438 1404 1439 1408
rect 1443 1404 1444 1408
rect 1438 1403 1444 1404
rect 1494 1408 1500 1409
rect 1494 1404 1495 1408
rect 1499 1404 1500 1408
rect 1494 1403 1500 1404
rect 1550 1408 1556 1409
rect 1550 1404 1551 1408
rect 1555 1404 1556 1408
rect 1550 1403 1556 1404
rect 1606 1408 1612 1409
rect 1606 1404 1607 1408
rect 1611 1404 1612 1408
rect 1606 1403 1612 1404
rect 1670 1408 1676 1409
rect 1670 1404 1671 1408
rect 1675 1404 1676 1408
rect 1670 1403 1676 1404
rect 1734 1408 1740 1409
rect 1734 1404 1735 1408
rect 1739 1404 1740 1408
rect 1734 1403 1740 1404
rect 1280 1399 1282 1403
rect 1328 1399 1330 1403
rect 1384 1399 1386 1403
rect 1440 1399 1442 1403
rect 1496 1399 1498 1403
rect 1552 1399 1554 1403
rect 1608 1399 1610 1403
rect 1672 1399 1674 1403
rect 1736 1399 1738 1403
rect 1135 1398 1139 1399
rect 1135 1393 1139 1394
rect 1279 1398 1283 1399
rect 1279 1393 1283 1394
rect 1327 1398 1331 1399
rect 1327 1393 1331 1394
rect 1335 1398 1339 1399
rect 1335 1393 1339 1394
rect 1375 1398 1379 1399
rect 1375 1393 1379 1394
rect 1383 1398 1387 1399
rect 1383 1393 1387 1394
rect 1415 1398 1419 1399
rect 1415 1393 1419 1394
rect 1439 1398 1443 1399
rect 1439 1393 1443 1394
rect 1455 1398 1459 1399
rect 1455 1393 1459 1394
rect 1495 1398 1499 1399
rect 1495 1393 1499 1394
rect 1535 1398 1539 1399
rect 1535 1393 1539 1394
rect 1551 1398 1555 1399
rect 1551 1393 1555 1394
rect 1583 1398 1587 1399
rect 1583 1393 1587 1394
rect 1607 1398 1611 1399
rect 1607 1393 1611 1394
rect 1647 1398 1651 1399
rect 1647 1393 1651 1394
rect 1671 1398 1675 1399
rect 1671 1393 1675 1394
rect 1719 1398 1723 1399
rect 1719 1393 1723 1394
rect 1735 1398 1739 1399
rect 1735 1393 1739 1394
rect 1047 1390 1051 1391
rect 1047 1385 1051 1386
rect 1095 1390 1099 1391
rect 1136 1390 1138 1393
rect 1334 1392 1340 1393
rect 1095 1385 1099 1386
rect 1134 1389 1140 1390
rect 1134 1385 1135 1389
rect 1139 1385 1140 1389
rect 1334 1388 1335 1392
rect 1339 1388 1340 1392
rect 1334 1387 1340 1388
rect 1374 1392 1380 1393
rect 1374 1388 1375 1392
rect 1379 1388 1380 1392
rect 1374 1387 1380 1388
rect 1414 1392 1420 1393
rect 1414 1388 1415 1392
rect 1419 1388 1420 1392
rect 1414 1387 1420 1388
rect 1454 1392 1460 1393
rect 1454 1388 1455 1392
rect 1459 1388 1460 1392
rect 1454 1387 1460 1388
rect 1494 1392 1500 1393
rect 1494 1388 1495 1392
rect 1499 1388 1500 1392
rect 1494 1387 1500 1388
rect 1534 1392 1540 1393
rect 1534 1388 1535 1392
rect 1539 1388 1540 1392
rect 1534 1387 1540 1388
rect 1582 1392 1588 1393
rect 1582 1388 1583 1392
rect 1587 1388 1588 1392
rect 1582 1387 1588 1388
rect 1646 1392 1652 1393
rect 1646 1388 1647 1392
rect 1651 1388 1652 1392
rect 1646 1387 1652 1388
rect 1718 1392 1724 1393
rect 1718 1388 1719 1392
rect 1723 1388 1724 1392
rect 1718 1387 1724 1388
rect 1022 1379 1028 1380
rect 1022 1375 1023 1379
rect 1027 1375 1028 1379
rect 1022 1374 1028 1375
rect 1048 1373 1050 1385
rect 998 1372 1004 1373
rect 998 1368 999 1372
rect 1003 1368 1004 1372
rect 998 1367 1004 1368
rect 1046 1372 1052 1373
rect 1046 1368 1047 1372
rect 1051 1368 1052 1372
rect 1046 1367 1052 1368
rect 1096 1365 1098 1385
rect 1134 1384 1140 1385
rect 1744 1376 1746 1438
rect 1808 1437 1810 1449
rect 1888 1437 1890 1449
rect 1806 1436 1812 1437
rect 1806 1432 1807 1436
rect 1811 1432 1812 1436
rect 1806 1431 1812 1432
rect 1886 1436 1892 1437
rect 1886 1432 1887 1436
rect 1891 1432 1892 1436
rect 1886 1431 1892 1432
rect 1912 1424 1914 1462
rect 1920 1455 1922 1471
rect 1992 1455 1994 1471
rect 2020 1468 2022 1526
rect 2040 1476 2042 1526
rect 2118 1519 2124 1520
rect 2070 1516 2076 1517
rect 2070 1512 2071 1516
rect 2075 1512 2076 1516
rect 2118 1515 2119 1519
rect 2123 1515 2124 1519
rect 2118 1514 2124 1515
rect 2070 1511 2076 1512
rect 2120 1511 2122 1514
rect 2063 1510 2067 1511
rect 2063 1505 2067 1506
rect 2071 1510 2075 1511
rect 2071 1505 2075 1506
rect 2119 1510 2123 1511
rect 2119 1505 2123 1506
rect 2062 1504 2068 1505
rect 2062 1500 2063 1504
rect 2067 1500 2068 1504
rect 2120 1502 2122 1505
rect 2062 1499 2068 1500
rect 2118 1501 2124 1502
rect 2118 1497 2119 1501
rect 2123 1497 2124 1501
rect 2118 1496 2124 1497
rect 2078 1487 2084 1488
rect 2078 1483 2079 1487
rect 2083 1483 2084 1487
rect 2078 1482 2084 1483
rect 2086 1487 2092 1488
rect 2086 1483 2087 1487
rect 2091 1483 2092 1487
rect 2086 1482 2092 1483
rect 2118 1484 2124 1485
rect 2062 1476 2068 1477
rect 2038 1475 2044 1476
rect 2038 1471 2039 1475
rect 2043 1471 2044 1475
rect 2062 1472 2063 1476
rect 2067 1472 2068 1476
rect 2062 1471 2068 1472
rect 2038 1470 2044 1471
rect 2018 1467 2024 1468
rect 2018 1463 2019 1467
rect 2023 1463 2024 1467
rect 2018 1462 2024 1463
rect 2064 1455 2066 1471
rect 2080 1468 2082 1482
rect 2078 1467 2084 1468
rect 2078 1463 2079 1467
rect 2083 1463 2084 1467
rect 2078 1462 2084 1463
rect 1919 1454 1923 1455
rect 1919 1449 1923 1450
rect 1975 1454 1979 1455
rect 1975 1449 1979 1450
rect 1991 1454 1995 1455
rect 1991 1449 1995 1450
rect 2063 1454 2067 1455
rect 2063 1449 2067 1450
rect 1976 1437 1978 1449
rect 2064 1437 2066 1449
rect 2088 1444 2090 1482
rect 2118 1480 2119 1484
rect 2123 1480 2124 1484
rect 2118 1479 2124 1480
rect 2120 1455 2122 1479
rect 2119 1454 2123 1455
rect 2119 1449 2123 1450
rect 2078 1443 2084 1444
rect 2078 1439 2079 1443
rect 2083 1439 2084 1443
rect 2078 1438 2084 1439
rect 2086 1443 2092 1444
rect 2086 1439 2087 1443
rect 2091 1439 2092 1443
rect 2086 1438 2092 1439
rect 1974 1436 1980 1437
rect 1974 1432 1975 1436
rect 1979 1432 1980 1436
rect 1974 1431 1980 1432
rect 2062 1436 2068 1437
rect 2062 1432 2063 1436
rect 2067 1432 2068 1436
rect 2062 1431 2068 1432
rect 2080 1424 2082 1438
rect 2120 1429 2122 1449
rect 2118 1428 2124 1429
rect 2118 1424 2119 1428
rect 2123 1424 2124 1428
rect 1910 1423 1916 1424
rect 1910 1419 1911 1423
rect 1915 1419 1916 1423
rect 1910 1418 1916 1419
rect 2014 1423 2020 1424
rect 2014 1419 2015 1423
rect 2019 1419 2020 1423
rect 2014 1418 2020 1419
rect 2078 1423 2084 1424
rect 2118 1423 2124 1424
rect 2078 1419 2079 1423
rect 2083 1419 2084 1423
rect 2078 1418 2084 1419
rect 1806 1408 1812 1409
rect 1806 1404 1807 1408
rect 1811 1404 1812 1408
rect 1806 1403 1812 1404
rect 1886 1408 1892 1409
rect 1886 1404 1887 1408
rect 1891 1404 1892 1408
rect 1886 1403 1892 1404
rect 1974 1408 1980 1409
rect 1974 1404 1975 1408
rect 1979 1404 1980 1408
rect 1974 1403 1980 1404
rect 1808 1399 1810 1403
rect 1888 1399 1890 1403
rect 1976 1399 1978 1403
rect 1807 1398 1811 1399
rect 1807 1393 1811 1394
rect 1887 1398 1891 1399
rect 1887 1393 1891 1394
rect 1895 1398 1899 1399
rect 1895 1393 1899 1394
rect 1975 1398 1979 1399
rect 1975 1393 1979 1394
rect 1991 1398 1995 1399
rect 1991 1393 1995 1394
rect 1806 1392 1812 1393
rect 1806 1388 1807 1392
rect 1811 1388 1812 1392
rect 1806 1387 1812 1388
rect 1894 1392 1900 1393
rect 1894 1388 1895 1392
rect 1899 1388 1900 1392
rect 1894 1387 1900 1388
rect 1990 1392 1996 1393
rect 1990 1388 1991 1392
rect 1995 1388 1996 1392
rect 1990 1387 1996 1388
rect 1918 1383 1924 1384
rect 1918 1379 1919 1383
rect 1923 1379 1924 1383
rect 1918 1378 1924 1379
rect 1390 1375 1396 1376
rect 1134 1372 1140 1373
rect 1134 1368 1135 1372
rect 1139 1368 1140 1372
rect 1390 1371 1391 1375
rect 1395 1371 1396 1375
rect 1390 1370 1396 1371
rect 1422 1375 1428 1376
rect 1422 1371 1423 1375
rect 1427 1371 1428 1375
rect 1422 1370 1428 1371
rect 1430 1375 1436 1376
rect 1430 1371 1431 1375
rect 1435 1371 1436 1375
rect 1430 1370 1436 1371
rect 1482 1375 1488 1376
rect 1482 1371 1483 1375
rect 1487 1371 1488 1375
rect 1482 1370 1488 1371
rect 1502 1375 1508 1376
rect 1502 1371 1503 1375
rect 1507 1371 1508 1375
rect 1502 1370 1508 1371
rect 1542 1375 1548 1376
rect 1542 1371 1543 1375
rect 1547 1371 1548 1375
rect 1542 1370 1548 1371
rect 1662 1375 1668 1376
rect 1662 1371 1663 1375
rect 1667 1371 1668 1375
rect 1662 1370 1668 1371
rect 1742 1375 1748 1376
rect 1742 1371 1743 1375
rect 1747 1371 1748 1375
rect 1742 1370 1748 1371
rect 1134 1367 1140 1368
rect 1094 1364 1100 1365
rect 1094 1360 1095 1364
rect 1099 1360 1100 1364
rect 890 1359 896 1360
rect 890 1355 891 1359
rect 895 1355 896 1359
rect 890 1354 896 1355
rect 950 1359 956 1360
rect 950 1355 951 1359
rect 955 1355 956 1359
rect 950 1354 956 1355
rect 1086 1359 1092 1360
rect 1094 1359 1100 1360
rect 1086 1355 1087 1359
rect 1091 1355 1092 1359
rect 1086 1354 1092 1355
rect 854 1344 860 1345
rect 854 1340 855 1344
rect 859 1340 860 1344
rect 854 1339 860 1340
rect 926 1344 932 1345
rect 926 1340 927 1344
rect 931 1340 932 1344
rect 926 1339 932 1340
rect 998 1344 1004 1345
rect 998 1340 999 1344
rect 1003 1340 1004 1344
rect 998 1339 1004 1340
rect 1046 1344 1052 1345
rect 1046 1340 1047 1344
rect 1051 1340 1052 1344
rect 1046 1339 1052 1340
rect 856 1331 858 1339
rect 928 1331 930 1339
rect 1000 1331 1002 1339
rect 1048 1331 1050 1339
rect 1088 1336 1090 1354
rect 1094 1347 1100 1348
rect 1136 1347 1138 1367
rect 1334 1364 1340 1365
rect 1334 1360 1335 1364
rect 1339 1360 1340 1364
rect 1334 1359 1340 1360
rect 1374 1364 1380 1365
rect 1374 1360 1375 1364
rect 1379 1360 1380 1364
rect 1374 1359 1380 1360
rect 1336 1347 1338 1359
rect 1376 1347 1378 1359
rect 1392 1356 1394 1370
rect 1414 1364 1420 1365
rect 1414 1360 1415 1364
rect 1419 1360 1420 1364
rect 1414 1359 1420 1360
rect 1390 1355 1396 1356
rect 1390 1351 1391 1355
rect 1395 1351 1396 1355
rect 1390 1350 1396 1351
rect 1416 1347 1418 1359
rect 1424 1356 1426 1370
rect 1422 1355 1428 1356
rect 1422 1351 1423 1355
rect 1427 1351 1428 1355
rect 1422 1350 1428 1351
rect 1094 1343 1095 1347
rect 1099 1343 1100 1347
rect 1094 1342 1100 1343
rect 1135 1346 1139 1347
rect 1086 1335 1092 1336
rect 1086 1331 1087 1335
rect 1091 1331 1092 1335
rect 1096 1331 1098 1342
rect 1135 1341 1139 1342
rect 1159 1346 1163 1347
rect 1159 1341 1163 1342
rect 1223 1346 1227 1347
rect 1223 1341 1227 1342
rect 1311 1346 1315 1347
rect 1311 1341 1315 1342
rect 1335 1346 1339 1347
rect 1335 1341 1339 1342
rect 1375 1346 1379 1347
rect 1375 1341 1379 1342
rect 1407 1346 1411 1347
rect 1407 1341 1411 1342
rect 1415 1346 1419 1347
rect 1415 1341 1419 1342
rect 855 1330 859 1331
rect 855 1325 859 1326
rect 863 1330 867 1331
rect 863 1325 867 1326
rect 927 1330 931 1331
rect 927 1325 931 1326
rect 943 1330 947 1331
rect 943 1325 947 1326
rect 999 1330 1003 1331
rect 999 1325 1003 1326
rect 1023 1330 1027 1331
rect 1023 1325 1027 1326
rect 1047 1330 1051 1331
rect 1086 1330 1092 1331
rect 1095 1330 1099 1331
rect 1047 1325 1051 1326
rect 1095 1325 1099 1326
rect 862 1324 868 1325
rect 862 1320 863 1324
rect 867 1320 868 1324
rect 862 1319 868 1320
rect 942 1324 948 1325
rect 942 1320 943 1324
rect 947 1320 948 1324
rect 942 1319 948 1320
rect 1022 1324 1028 1325
rect 1022 1320 1023 1324
rect 1027 1320 1028 1324
rect 1096 1322 1098 1325
rect 1022 1319 1028 1320
rect 1094 1321 1100 1322
rect 1136 1321 1138 1341
rect 1160 1329 1162 1341
rect 1224 1329 1226 1341
rect 1312 1329 1314 1341
rect 1408 1329 1410 1341
rect 1432 1336 1434 1370
rect 1454 1364 1460 1365
rect 1454 1360 1455 1364
rect 1459 1360 1460 1364
rect 1454 1359 1460 1360
rect 1456 1347 1458 1359
rect 1484 1348 1486 1370
rect 1494 1364 1500 1365
rect 1494 1360 1495 1364
rect 1499 1360 1500 1364
rect 1494 1359 1500 1360
rect 1482 1347 1488 1348
rect 1496 1347 1498 1359
rect 1504 1356 1506 1370
rect 1534 1364 1540 1365
rect 1534 1360 1535 1364
rect 1539 1360 1540 1364
rect 1534 1359 1540 1360
rect 1502 1355 1508 1356
rect 1502 1351 1503 1355
rect 1507 1351 1508 1355
rect 1502 1350 1508 1351
rect 1536 1347 1538 1359
rect 1544 1356 1546 1370
rect 1582 1364 1588 1365
rect 1582 1360 1583 1364
rect 1587 1360 1588 1364
rect 1582 1359 1588 1360
rect 1646 1364 1652 1365
rect 1646 1360 1647 1364
rect 1651 1360 1652 1364
rect 1646 1359 1652 1360
rect 1542 1355 1548 1356
rect 1542 1351 1543 1355
rect 1547 1351 1548 1355
rect 1542 1350 1548 1351
rect 1584 1347 1586 1359
rect 1590 1355 1596 1356
rect 1590 1351 1591 1355
rect 1595 1351 1596 1355
rect 1590 1350 1596 1351
rect 1455 1346 1459 1347
rect 1482 1343 1483 1347
rect 1487 1343 1488 1347
rect 1482 1342 1488 1343
rect 1495 1346 1499 1347
rect 1455 1341 1459 1342
rect 1495 1341 1499 1342
rect 1503 1346 1507 1347
rect 1503 1341 1507 1342
rect 1535 1346 1539 1347
rect 1535 1341 1539 1342
rect 1583 1346 1587 1347
rect 1583 1341 1587 1342
rect 1430 1335 1436 1336
rect 1430 1331 1431 1335
rect 1435 1331 1436 1335
rect 1430 1330 1436 1331
rect 1504 1329 1506 1341
rect 1158 1328 1164 1329
rect 1158 1324 1159 1328
rect 1163 1324 1164 1328
rect 1158 1323 1164 1324
rect 1222 1328 1228 1329
rect 1222 1324 1223 1328
rect 1227 1324 1228 1328
rect 1222 1323 1228 1324
rect 1310 1328 1316 1329
rect 1310 1324 1311 1328
rect 1315 1324 1316 1328
rect 1310 1323 1316 1324
rect 1406 1328 1412 1329
rect 1406 1324 1407 1328
rect 1411 1324 1412 1328
rect 1406 1323 1412 1324
rect 1502 1328 1508 1329
rect 1502 1324 1503 1328
rect 1507 1324 1508 1328
rect 1502 1323 1508 1324
rect 1094 1317 1095 1321
rect 1099 1317 1100 1321
rect 1094 1316 1100 1317
rect 1134 1320 1140 1321
rect 1134 1316 1135 1320
rect 1139 1316 1140 1320
rect 1592 1316 1594 1350
rect 1648 1347 1650 1359
rect 1664 1356 1666 1370
rect 1718 1364 1724 1365
rect 1718 1360 1719 1364
rect 1723 1360 1724 1364
rect 1718 1359 1724 1360
rect 1806 1364 1812 1365
rect 1806 1360 1807 1364
rect 1811 1360 1812 1364
rect 1806 1359 1812 1360
rect 1894 1364 1900 1365
rect 1894 1360 1895 1364
rect 1899 1360 1900 1364
rect 1894 1359 1900 1360
rect 1662 1355 1668 1356
rect 1662 1351 1663 1355
rect 1667 1351 1668 1355
rect 1662 1350 1668 1351
rect 1720 1347 1722 1359
rect 1808 1347 1810 1359
rect 1896 1347 1898 1359
rect 1920 1356 1922 1378
rect 1990 1364 1996 1365
rect 1990 1360 1991 1364
rect 1995 1360 1996 1364
rect 1990 1359 1996 1360
rect 1918 1355 1924 1356
rect 1918 1351 1919 1355
rect 1923 1351 1924 1355
rect 1918 1350 1924 1351
rect 1992 1347 1994 1359
rect 2016 1356 2018 1418
rect 2118 1411 2124 1412
rect 2062 1408 2068 1409
rect 2062 1404 2063 1408
rect 2067 1404 2068 1408
rect 2118 1407 2119 1411
rect 2123 1407 2124 1411
rect 2118 1406 2124 1407
rect 2062 1403 2068 1404
rect 2064 1399 2066 1403
rect 2120 1399 2122 1406
rect 2063 1398 2067 1399
rect 2063 1393 2067 1394
rect 2071 1398 2075 1399
rect 2071 1393 2075 1394
rect 2119 1398 2123 1399
rect 2119 1393 2123 1394
rect 2070 1392 2076 1393
rect 2070 1388 2071 1392
rect 2075 1388 2076 1392
rect 2120 1390 2122 1393
rect 2070 1387 2076 1388
rect 2118 1389 2124 1390
rect 2118 1385 2119 1389
rect 2123 1385 2124 1389
rect 2118 1384 2124 1385
rect 2086 1375 2092 1376
rect 2086 1371 2087 1375
rect 2091 1371 2092 1375
rect 2086 1370 2092 1371
rect 2094 1375 2100 1376
rect 2094 1371 2095 1375
rect 2099 1371 2100 1375
rect 2094 1370 2100 1371
rect 2118 1372 2124 1373
rect 2070 1364 2076 1365
rect 2070 1360 2071 1364
rect 2075 1360 2076 1364
rect 2070 1359 2076 1360
rect 2014 1355 2020 1356
rect 2014 1351 2015 1355
rect 2019 1351 2020 1355
rect 2014 1350 2020 1351
rect 2072 1347 2074 1359
rect 2088 1356 2090 1370
rect 2086 1355 2092 1356
rect 2086 1351 2087 1355
rect 2091 1351 2092 1355
rect 2086 1350 2092 1351
rect 1599 1346 1603 1347
rect 1599 1341 1603 1342
rect 1647 1346 1651 1347
rect 1647 1341 1651 1342
rect 1679 1346 1683 1347
rect 1679 1341 1683 1342
rect 1719 1346 1723 1347
rect 1719 1341 1723 1342
rect 1759 1346 1763 1347
rect 1759 1341 1763 1342
rect 1807 1346 1811 1347
rect 1807 1341 1811 1342
rect 1831 1346 1835 1347
rect 1831 1341 1835 1342
rect 1895 1346 1899 1347
rect 1895 1341 1899 1342
rect 1959 1346 1963 1347
rect 1959 1341 1963 1342
rect 1991 1346 1995 1347
rect 1991 1341 1995 1342
rect 2023 1346 2027 1347
rect 2023 1341 2027 1342
rect 2071 1346 2075 1347
rect 2071 1341 2075 1342
rect 1600 1329 1602 1341
rect 1680 1329 1682 1341
rect 1760 1329 1762 1341
rect 1774 1335 1780 1336
rect 1774 1331 1775 1335
rect 1779 1331 1780 1335
rect 1774 1330 1780 1331
rect 1598 1328 1604 1329
rect 1598 1324 1599 1328
rect 1603 1324 1604 1328
rect 1598 1323 1604 1324
rect 1678 1328 1684 1329
rect 1678 1324 1679 1328
rect 1683 1324 1684 1328
rect 1678 1323 1684 1324
rect 1758 1328 1764 1329
rect 1758 1324 1759 1328
rect 1763 1324 1764 1328
rect 1758 1323 1764 1324
rect 1776 1316 1778 1330
rect 1832 1329 1834 1341
rect 1846 1335 1852 1336
rect 1846 1331 1847 1335
rect 1851 1331 1852 1335
rect 1846 1330 1852 1331
rect 1830 1328 1836 1329
rect 1830 1324 1831 1328
rect 1835 1324 1836 1328
rect 1830 1323 1836 1324
rect 1848 1316 1850 1330
rect 1896 1329 1898 1341
rect 1910 1335 1916 1336
rect 1910 1331 1911 1335
rect 1915 1331 1916 1335
rect 1910 1330 1916 1331
rect 1894 1328 1900 1329
rect 1894 1324 1895 1328
rect 1899 1324 1900 1328
rect 1894 1323 1900 1324
rect 1912 1316 1914 1330
rect 1960 1329 1962 1341
rect 1974 1335 1980 1336
rect 1974 1331 1975 1335
rect 1979 1331 1980 1335
rect 1974 1330 1980 1331
rect 1958 1328 1964 1329
rect 1958 1324 1959 1328
rect 1963 1324 1964 1328
rect 1958 1323 1964 1324
rect 1976 1316 1978 1330
rect 2024 1329 2026 1341
rect 2038 1335 2044 1336
rect 2038 1331 2039 1335
rect 2043 1331 2044 1335
rect 2038 1330 2044 1331
rect 2046 1335 2052 1336
rect 2046 1331 2047 1335
rect 2051 1331 2052 1335
rect 2046 1330 2052 1331
rect 2022 1328 2028 1329
rect 2022 1324 2023 1328
rect 2027 1324 2028 1328
rect 2022 1323 2028 1324
rect 2040 1316 2042 1330
rect 1134 1315 1140 1316
rect 1330 1315 1336 1316
rect 1330 1311 1331 1315
rect 1335 1311 1336 1315
rect 1330 1310 1336 1311
rect 1590 1315 1596 1316
rect 1590 1311 1591 1315
rect 1595 1311 1596 1315
rect 1590 1310 1596 1311
rect 1766 1315 1772 1316
rect 1766 1311 1767 1315
rect 1771 1311 1772 1315
rect 1766 1310 1772 1311
rect 1774 1315 1780 1316
rect 1774 1311 1775 1315
rect 1779 1311 1780 1315
rect 1774 1310 1780 1311
rect 1846 1315 1852 1316
rect 1846 1311 1847 1315
rect 1851 1311 1852 1315
rect 1846 1310 1852 1311
rect 1910 1315 1916 1316
rect 1910 1311 1911 1315
rect 1915 1311 1916 1315
rect 1910 1310 1916 1311
rect 1974 1315 1980 1316
rect 1974 1311 1975 1315
rect 1979 1311 1980 1315
rect 1974 1310 1980 1311
rect 2038 1315 2044 1316
rect 2038 1311 2039 1315
rect 2043 1311 2044 1315
rect 2038 1310 2044 1311
rect 638 1307 644 1308
rect 638 1303 639 1307
rect 643 1303 644 1307
rect 638 1302 644 1303
rect 718 1307 724 1308
rect 718 1303 719 1307
rect 723 1303 724 1307
rect 718 1302 724 1303
rect 730 1307 736 1308
rect 730 1303 731 1307
rect 735 1303 736 1307
rect 730 1302 736 1303
rect 806 1307 812 1308
rect 806 1303 807 1307
rect 811 1303 812 1307
rect 806 1302 812 1303
rect 1094 1304 1100 1305
rect 390 1296 396 1297
rect 390 1292 391 1296
rect 395 1292 396 1296
rect 390 1291 396 1292
rect 462 1296 468 1297
rect 462 1292 463 1296
rect 467 1292 468 1296
rect 462 1291 468 1292
rect 542 1296 548 1297
rect 542 1292 543 1296
rect 547 1292 548 1296
rect 542 1291 548 1292
rect 622 1296 628 1297
rect 622 1292 623 1296
rect 627 1292 628 1296
rect 622 1291 628 1292
rect 374 1279 380 1280
rect 374 1275 375 1279
rect 379 1275 380 1279
rect 392 1275 394 1291
rect 464 1275 466 1291
rect 544 1275 546 1291
rect 550 1287 556 1288
rect 550 1283 551 1287
rect 555 1283 556 1287
rect 550 1282 556 1283
rect 319 1274 323 1275
rect 374 1274 380 1275
rect 391 1274 395 1275
rect 255 1269 259 1270
rect 278 1271 284 1272
rect 112 1249 114 1269
rect 136 1257 138 1269
rect 176 1257 178 1269
rect 190 1263 196 1264
rect 190 1259 191 1263
rect 195 1259 196 1263
rect 190 1258 196 1259
rect 134 1256 140 1257
rect 134 1252 135 1256
rect 139 1252 140 1256
rect 134 1251 140 1252
rect 174 1256 180 1257
rect 174 1252 175 1256
rect 179 1252 180 1256
rect 174 1251 180 1252
rect 110 1248 116 1249
rect 110 1244 111 1248
rect 115 1244 116 1248
rect 192 1244 194 1258
rect 216 1257 218 1269
rect 230 1263 236 1264
rect 230 1259 231 1263
rect 235 1259 236 1263
rect 230 1258 236 1259
rect 214 1256 220 1257
rect 214 1252 215 1256
rect 219 1252 220 1256
rect 214 1251 220 1252
rect 232 1244 234 1258
rect 256 1257 258 1269
rect 278 1267 279 1271
rect 283 1267 284 1271
rect 319 1269 323 1270
rect 391 1269 395 1270
rect 399 1274 403 1275
rect 399 1269 403 1270
rect 463 1274 467 1275
rect 463 1269 467 1270
rect 487 1274 491 1275
rect 487 1269 491 1270
rect 543 1274 547 1275
rect 543 1269 547 1270
rect 278 1266 284 1267
rect 320 1257 322 1269
rect 400 1257 402 1269
rect 488 1257 490 1269
rect 254 1256 260 1257
rect 254 1252 255 1256
rect 259 1252 260 1256
rect 254 1251 260 1252
rect 318 1256 324 1257
rect 318 1252 319 1256
rect 323 1252 324 1256
rect 318 1251 324 1252
rect 398 1256 404 1257
rect 398 1252 399 1256
rect 403 1252 404 1256
rect 398 1251 404 1252
rect 486 1256 492 1257
rect 486 1252 487 1256
rect 491 1252 492 1256
rect 486 1251 492 1252
rect 552 1244 554 1282
rect 624 1275 626 1291
rect 640 1288 642 1302
rect 702 1296 708 1297
rect 702 1292 703 1296
rect 707 1292 708 1296
rect 702 1291 708 1292
rect 638 1287 644 1288
rect 638 1283 639 1287
rect 643 1283 644 1287
rect 638 1282 644 1283
rect 704 1275 706 1291
rect 720 1288 722 1302
rect 1094 1300 1095 1304
rect 1099 1300 1100 1304
rect 1094 1299 1100 1300
rect 1134 1303 1140 1304
rect 1134 1299 1135 1303
rect 1139 1299 1140 1303
rect 782 1296 788 1297
rect 782 1292 783 1296
rect 787 1292 788 1296
rect 782 1291 788 1292
rect 862 1296 868 1297
rect 862 1292 863 1296
rect 867 1292 868 1296
rect 862 1291 868 1292
rect 942 1296 948 1297
rect 942 1292 943 1296
rect 947 1292 948 1296
rect 942 1291 948 1292
rect 1022 1296 1028 1297
rect 1022 1292 1023 1296
rect 1027 1292 1028 1296
rect 1022 1291 1028 1292
rect 718 1287 724 1288
rect 718 1283 719 1287
rect 723 1283 724 1287
rect 718 1282 724 1283
rect 784 1275 786 1291
rect 864 1275 866 1291
rect 944 1275 946 1291
rect 1024 1275 1026 1291
rect 1070 1287 1076 1288
rect 1070 1283 1071 1287
rect 1075 1283 1076 1287
rect 1070 1282 1076 1283
rect 583 1274 587 1275
rect 574 1271 580 1272
rect 574 1267 575 1271
rect 579 1267 580 1271
rect 583 1269 587 1270
rect 623 1274 627 1275
rect 623 1269 627 1270
rect 687 1274 691 1275
rect 687 1269 691 1270
rect 703 1274 707 1275
rect 703 1269 707 1270
rect 783 1274 787 1275
rect 783 1269 787 1270
rect 799 1274 803 1275
rect 799 1269 803 1270
rect 863 1274 867 1275
rect 863 1269 867 1270
rect 919 1274 923 1275
rect 919 1269 923 1270
rect 943 1274 947 1275
rect 943 1269 947 1270
rect 1023 1274 1027 1275
rect 1023 1269 1027 1270
rect 1047 1274 1051 1275
rect 1047 1269 1051 1270
rect 574 1266 580 1267
rect 110 1243 116 1244
rect 190 1243 196 1244
rect 190 1239 191 1243
rect 195 1239 196 1243
rect 190 1238 196 1239
rect 230 1243 236 1244
rect 230 1239 231 1243
rect 235 1239 236 1243
rect 230 1238 236 1239
rect 378 1243 384 1244
rect 378 1239 379 1243
rect 383 1239 384 1243
rect 378 1238 384 1239
rect 550 1243 556 1244
rect 550 1239 551 1243
rect 555 1239 556 1243
rect 550 1238 556 1239
rect 110 1231 116 1232
rect 110 1227 111 1231
rect 115 1227 116 1231
rect 110 1226 116 1227
rect 134 1228 140 1229
rect 112 1219 114 1226
rect 134 1224 135 1228
rect 139 1224 140 1228
rect 134 1223 140 1224
rect 174 1228 180 1229
rect 174 1224 175 1228
rect 179 1224 180 1228
rect 174 1223 180 1224
rect 214 1228 220 1229
rect 214 1224 215 1228
rect 219 1224 220 1228
rect 214 1223 220 1224
rect 254 1228 260 1229
rect 254 1224 255 1228
rect 259 1224 260 1228
rect 254 1223 260 1224
rect 318 1228 324 1229
rect 318 1224 319 1228
rect 323 1224 324 1228
rect 318 1223 324 1224
rect 136 1219 138 1223
rect 176 1219 178 1223
rect 216 1219 218 1223
rect 256 1219 258 1223
rect 320 1219 322 1223
rect 111 1218 115 1219
rect 111 1213 115 1214
rect 135 1218 139 1219
rect 135 1213 139 1214
rect 175 1218 179 1219
rect 175 1213 179 1214
rect 215 1218 219 1219
rect 215 1213 219 1214
rect 255 1218 259 1219
rect 255 1213 259 1214
rect 271 1218 275 1219
rect 271 1213 275 1214
rect 311 1218 315 1219
rect 311 1213 315 1214
rect 319 1218 323 1219
rect 319 1213 323 1214
rect 351 1218 355 1219
rect 351 1213 355 1214
rect 112 1210 114 1213
rect 270 1212 276 1213
rect 110 1209 116 1210
rect 110 1205 111 1209
rect 115 1205 116 1209
rect 270 1208 271 1212
rect 275 1208 276 1212
rect 270 1207 276 1208
rect 310 1212 316 1213
rect 310 1208 311 1212
rect 315 1208 316 1212
rect 310 1207 316 1208
rect 350 1212 356 1213
rect 350 1208 351 1212
rect 355 1208 356 1212
rect 350 1207 356 1208
rect 110 1204 116 1205
rect 326 1195 332 1196
rect 110 1192 116 1193
rect 110 1188 111 1192
rect 115 1188 116 1192
rect 326 1191 327 1195
rect 331 1191 332 1195
rect 326 1190 332 1191
rect 358 1195 364 1196
rect 358 1191 359 1195
rect 363 1191 364 1195
rect 358 1190 364 1191
rect 110 1187 116 1188
rect 112 1163 114 1187
rect 270 1184 276 1185
rect 270 1180 271 1184
rect 275 1180 276 1184
rect 270 1179 276 1180
rect 310 1184 316 1185
rect 310 1180 311 1184
rect 315 1180 316 1184
rect 310 1179 316 1180
rect 272 1163 274 1179
rect 312 1163 314 1179
rect 328 1176 330 1190
rect 350 1184 356 1185
rect 350 1180 351 1184
rect 355 1180 356 1184
rect 350 1179 356 1180
rect 326 1175 332 1176
rect 326 1171 327 1175
rect 331 1171 332 1175
rect 326 1170 332 1171
rect 352 1163 354 1179
rect 360 1176 362 1190
rect 380 1176 382 1238
rect 398 1228 404 1229
rect 398 1224 399 1228
rect 403 1224 404 1228
rect 398 1223 404 1224
rect 486 1228 492 1229
rect 486 1224 487 1228
rect 491 1224 492 1228
rect 486 1223 492 1224
rect 400 1219 402 1223
rect 488 1219 490 1223
rect 399 1218 403 1219
rect 399 1213 403 1214
rect 447 1218 451 1219
rect 447 1213 451 1214
rect 487 1218 491 1219
rect 487 1213 491 1214
rect 495 1218 499 1219
rect 495 1213 499 1214
rect 551 1218 555 1219
rect 551 1213 555 1214
rect 398 1212 404 1213
rect 398 1208 399 1212
rect 403 1208 404 1212
rect 398 1207 404 1208
rect 446 1212 452 1213
rect 446 1208 447 1212
rect 451 1208 452 1212
rect 446 1207 452 1208
rect 494 1212 500 1213
rect 494 1208 495 1212
rect 499 1208 500 1212
rect 494 1207 500 1208
rect 550 1212 556 1213
rect 550 1208 551 1212
rect 555 1208 556 1212
rect 550 1207 556 1208
rect 422 1203 428 1204
rect 422 1199 423 1203
rect 427 1199 428 1203
rect 422 1198 428 1199
rect 398 1184 404 1185
rect 398 1180 399 1184
rect 403 1180 404 1184
rect 398 1179 404 1180
rect 358 1175 364 1176
rect 358 1171 359 1175
rect 363 1171 364 1175
rect 358 1170 364 1171
rect 378 1175 384 1176
rect 378 1171 379 1175
rect 383 1171 384 1175
rect 378 1170 384 1171
rect 400 1163 402 1179
rect 424 1176 426 1198
rect 576 1196 578 1266
rect 584 1257 586 1269
rect 598 1263 604 1264
rect 598 1259 599 1263
rect 603 1259 604 1263
rect 598 1258 604 1259
rect 582 1256 588 1257
rect 582 1252 583 1256
rect 587 1252 588 1256
rect 582 1251 588 1252
rect 600 1244 602 1258
rect 688 1257 690 1269
rect 702 1263 708 1264
rect 702 1259 703 1263
rect 707 1259 708 1263
rect 702 1258 708 1259
rect 686 1256 692 1257
rect 686 1252 687 1256
rect 691 1252 692 1256
rect 686 1251 692 1252
rect 704 1244 706 1258
rect 800 1257 802 1269
rect 814 1263 820 1264
rect 814 1259 815 1263
rect 819 1259 820 1263
rect 814 1258 820 1259
rect 798 1256 804 1257
rect 798 1252 799 1256
rect 803 1252 804 1256
rect 798 1251 804 1252
rect 816 1244 818 1258
rect 920 1257 922 1269
rect 1006 1263 1012 1264
rect 1006 1259 1007 1263
rect 1011 1259 1012 1263
rect 1006 1258 1012 1259
rect 1014 1263 1020 1264
rect 1014 1259 1015 1263
rect 1019 1259 1020 1263
rect 1014 1258 1020 1259
rect 918 1256 924 1257
rect 918 1252 919 1256
rect 923 1252 924 1256
rect 918 1251 924 1252
rect 598 1243 604 1244
rect 598 1239 599 1243
rect 603 1239 604 1243
rect 598 1238 604 1239
rect 702 1243 708 1244
rect 702 1239 703 1243
rect 707 1239 708 1243
rect 702 1238 708 1239
rect 814 1243 820 1244
rect 814 1239 815 1243
rect 819 1239 820 1243
rect 814 1238 820 1239
rect 582 1228 588 1229
rect 582 1224 583 1228
rect 587 1224 588 1228
rect 582 1223 588 1224
rect 686 1228 692 1229
rect 686 1224 687 1228
rect 691 1224 692 1228
rect 686 1223 692 1224
rect 798 1228 804 1229
rect 798 1224 799 1228
rect 803 1224 804 1228
rect 798 1223 804 1224
rect 918 1228 924 1229
rect 918 1224 919 1228
rect 923 1224 924 1228
rect 918 1223 924 1224
rect 584 1219 586 1223
rect 688 1219 690 1223
rect 800 1219 802 1223
rect 920 1219 922 1223
rect 583 1218 587 1219
rect 583 1213 587 1214
rect 607 1218 611 1219
rect 607 1213 611 1214
rect 671 1218 675 1219
rect 671 1213 675 1214
rect 687 1218 691 1219
rect 687 1213 691 1214
rect 743 1218 747 1219
rect 743 1213 747 1214
rect 799 1218 803 1219
rect 799 1213 803 1214
rect 815 1218 819 1219
rect 815 1213 819 1214
rect 895 1218 899 1219
rect 895 1213 899 1214
rect 919 1218 923 1219
rect 919 1213 923 1214
rect 983 1218 987 1219
rect 983 1213 987 1214
rect 606 1212 612 1213
rect 606 1208 607 1212
rect 611 1208 612 1212
rect 606 1207 612 1208
rect 670 1212 676 1213
rect 670 1208 671 1212
rect 675 1208 676 1212
rect 670 1207 676 1208
rect 742 1212 748 1213
rect 742 1208 743 1212
rect 747 1208 748 1212
rect 742 1207 748 1208
rect 814 1212 820 1213
rect 814 1208 815 1212
rect 819 1208 820 1212
rect 814 1207 820 1208
rect 894 1212 900 1213
rect 894 1208 895 1212
rect 899 1208 900 1212
rect 894 1207 900 1208
rect 982 1212 988 1213
rect 982 1208 983 1212
rect 987 1208 988 1212
rect 982 1207 988 1208
rect 1008 1196 1010 1258
rect 1016 1244 1018 1258
rect 1048 1257 1050 1269
rect 1046 1256 1052 1257
rect 1046 1252 1047 1256
rect 1051 1252 1052 1256
rect 1046 1251 1052 1252
rect 1072 1244 1074 1282
rect 1096 1275 1098 1299
rect 1134 1298 1140 1299
rect 1158 1300 1164 1301
rect 1136 1295 1138 1298
rect 1158 1296 1159 1300
rect 1163 1296 1164 1300
rect 1158 1295 1164 1296
rect 1222 1300 1228 1301
rect 1222 1296 1223 1300
rect 1227 1296 1228 1300
rect 1222 1295 1228 1296
rect 1310 1300 1316 1301
rect 1310 1296 1311 1300
rect 1315 1296 1316 1300
rect 1310 1295 1316 1296
rect 1135 1294 1139 1295
rect 1135 1289 1139 1290
rect 1159 1294 1163 1295
rect 1159 1289 1163 1290
rect 1175 1294 1179 1295
rect 1175 1289 1179 1290
rect 1223 1294 1227 1295
rect 1223 1289 1227 1290
rect 1231 1294 1235 1295
rect 1231 1289 1235 1290
rect 1303 1294 1307 1295
rect 1303 1289 1307 1290
rect 1311 1294 1315 1295
rect 1311 1289 1315 1290
rect 1136 1286 1138 1289
rect 1174 1288 1180 1289
rect 1134 1285 1140 1286
rect 1134 1281 1135 1285
rect 1139 1281 1140 1285
rect 1174 1284 1175 1288
rect 1179 1284 1180 1288
rect 1174 1283 1180 1284
rect 1230 1288 1236 1289
rect 1230 1284 1231 1288
rect 1235 1284 1236 1288
rect 1230 1283 1236 1284
rect 1302 1288 1308 1289
rect 1302 1284 1303 1288
rect 1307 1284 1308 1288
rect 1302 1283 1308 1284
rect 1134 1280 1140 1281
rect 1095 1274 1099 1275
rect 1095 1269 1099 1270
rect 1198 1271 1204 1272
rect 1096 1249 1098 1269
rect 1134 1268 1140 1269
rect 1134 1264 1135 1268
rect 1139 1264 1140 1268
rect 1198 1267 1199 1271
rect 1203 1267 1204 1271
rect 1198 1266 1204 1267
rect 1134 1263 1140 1264
rect 1094 1248 1100 1249
rect 1094 1244 1095 1248
rect 1099 1244 1100 1248
rect 1014 1243 1020 1244
rect 1014 1239 1015 1243
rect 1019 1239 1020 1243
rect 1014 1238 1020 1239
rect 1070 1243 1076 1244
rect 1094 1243 1100 1244
rect 1070 1239 1071 1243
rect 1075 1239 1076 1243
rect 1136 1239 1138 1263
rect 1200 1261 1202 1266
rect 1174 1260 1180 1261
rect 1174 1256 1175 1260
rect 1179 1256 1180 1260
rect 1174 1255 1180 1256
rect 1199 1260 1203 1261
rect 1199 1255 1203 1256
rect 1230 1260 1236 1261
rect 1230 1256 1231 1260
rect 1235 1256 1236 1260
rect 1230 1255 1236 1256
rect 1302 1260 1308 1261
rect 1302 1256 1303 1260
rect 1307 1256 1308 1260
rect 1302 1255 1308 1256
rect 1176 1239 1178 1255
rect 1232 1239 1234 1255
rect 1304 1239 1306 1255
rect 1332 1252 1334 1310
rect 1406 1300 1412 1301
rect 1406 1296 1407 1300
rect 1411 1296 1412 1300
rect 1406 1295 1412 1296
rect 1502 1300 1508 1301
rect 1502 1296 1503 1300
rect 1507 1296 1508 1300
rect 1502 1295 1508 1296
rect 1598 1300 1604 1301
rect 1598 1296 1599 1300
rect 1603 1296 1604 1300
rect 1598 1295 1604 1296
rect 1678 1300 1684 1301
rect 1678 1296 1679 1300
rect 1683 1296 1684 1300
rect 1678 1295 1684 1296
rect 1758 1300 1764 1301
rect 1758 1296 1759 1300
rect 1763 1296 1764 1300
rect 1758 1295 1764 1296
rect 1391 1294 1395 1295
rect 1391 1289 1395 1290
rect 1407 1294 1411 1295
rect 1407 1289 1411 1290
rect 1479 1294 1483 1295
rect 1479 1289 1483 1290
rect 1503 1294 1507 1295
rect 1503 1289 1507 1290
rect 1567 1294 1571 1295
rect 1567 1289 1571 1290
rect 1599 1294 1603 1295
rect 1599 1289 1603 1290
rect 1655 1294 1659 1295
rect 1655 1289 1659 1290
rect 1679 1294 1683 1295
rect 1679 1289 1683 1290
rect 1743 1294 1747 1295
rect 1743 1289 1747 1290
rect 1759 1294 1763 1295
rect 1759 1289 1763 1290
rect 1390 1288 1396 1289
rect 1390 1284 1391 1288
rect 1395 1284 1396 1288
rect 1390 1283 1396 1284
rect 1478 1288 1484 1289
rect 1478 1284 1479 1288
rect 1483 1284 1484 1288
rect 1478 1283 1484 1284
rect 1566 1288 1572 1289
rect 1566 1284 1567 1288
rect 1571 1284 1572 1288
rect 1566 1283 1572 1284
rect 1654 1288 1660 1289
rect 1654 1284 1655 1288
rect 1659 1284 1660 1288
rect 1654 1283 1660 1284
rect 1742 1288 1748 1289
rect 1742 1284 1743 1288
rect 1747 1284 1748 1288
rect 1742 1283 1748 1284
rect 1410 1271 1416 1272
rect 1410 1267 1411 1271
rect 1415 1267 1416 1271
rect 1410 1266 1416 1267
rect 1670 1271 1676 1272
rect 1670 1267 1671 1271
rect 1675 1267 1676 1271
rect 1670 1266 1676 1267
rect 1390 1260 1396 1261
rect 1390 1256 1391 1260
rect 1395 1256 1396 1260
rect 1390 1255 1396 1256
rect 1330 1251 1336 1252
rect 1330 1247 1331 1251
rect 1335 1247 1336 1251
rect 1330 1246 1336 1247
rect 1392 1239 1394 1255
rect 1070 1238 1076 1239
rect 1135 1238 1139 1239
rect 1135 1233 1139 1234
rect 1175 1238 1179 1239
rect 1175 1233 1179 1234
rect 1231 1238 1235 1239
rect 1231 1233 1235 1234
rect 1287 1238 1291 1239
rect 1287 1233 1291 1234
rect 1303 1238 1307 1239
rect 1327 1238 1331 1239
rect 1303 1233 1307 1234
rect 1314 1235 1320 1236
rect 1094 1231 1100 1232
rect 1046 1228 1052 1229
rect 1046 1224 1047 1228
rect 1051 1224 1052 1228
rect 1094 1227 1095 1231
rect 1099 1227 1100 1231
rect 1094 1226 1100 1227
rect 1046 1223 1052 1224
rect 1048 1219 1050 1223
rect 1096 1219 1098 1226
rect 1047 1218 1051 1219
rect 1047 1213 1051 1214
rect 1095 1218 1099 1219
rect 1095 1213 1099 1214
rect 1136 1213 1138 1233
rect 1288 1221 1290 1233
rect 1314 1231 1315 1235
rect 1319 1231 1320 1235
rect 1327 1233 1331 1234
rect 1375 1238 1379 1239
rect 1375 1233 1379 1234
rect 1391 1238 1395 1239
rect 1391 1233 1395 1234
rect 1314 1230 1320 1231
rect 1286 1220 1292 1221
rect 1286 1216 1287 1220
rect 1291 1216 1292 1220
rect 1286 1215 1292 1216
rect 1096 1210 1098 1213
rect 1134 1212 1140 1213
rect 1094 1209 1100 1210
rect 1094 1205 1095 1209
rect 1099 1205 1100 1209
rect 1134 1208 1135 1212
rect 1139 1208 1140 1212
rect 1316 1208 1318 1230
rect 1328 1221 1330 1233
rect 1342 1227 1348 1228
rect 1342 1223 1343 1227
rect 1347 1223 1348 1227
rect 1342 1222 1348 1223
rect 1326 1220 1332 1221
rect 1326 1216 1327 1220
rect 1331 1216 1332 1220
rect 1326 1215 1332 1216
rect 1344 1208 1346 1222
rect 1376 1221 1378 1233
rect 1412 1228 1414 1266
rect 1478 1260 1484 1261
rect 1478 1256 1479 1260
rect 1483 1256 1484 1260
rect 1478 1255 1484 1256
rect 1566 1260 1572 1261
rect 1566 1256 1567 1260
rect 1571 1256 1572 1260
rect 1566 1255 1572 1256
rect 1591 1260 1595 1261
rect 1591 1255 1595 1256
rect 1654 1260 1660 1261
rect 1654 1256 1655 1260
rect 1659 1256 1660 1260
rect 1654 1255 1660 1256
rect 1480 1239 1482 1255
rect 1568 1239 1570 1255
rect 1592 1252 1594 1255
rect 1590 1251 1596 1252
rect 1590 1247 1591 1251
rect 1595 1247 1596 1251
rect 1590 1246 1596 1247
rect 1656 1239 1658 1255
rect 1431 1238 1435 1239
rect 1479 1238 1483 1239
rect 1431 1233 1435 1234
rect 1458 1235 1464 1236
rect 1390 1227 1396 1228
rect 1390 1223 1391 1227
rect 1395 1223 1396 1227
rect 1390 1222 1396 1223
rect 1410 1227 1416 1228
rect 1410 1223 1411 1227
rect 1415 1223 1416 1227
rect 1410 1222 1416 1223
rect 1374 1220 1380 1221
rect 1374 1216 1375 1220
rect 1379 1216 1380 1220
rect 1374 1215 1380 1216
rect 1392 1208 1394 1222
rect 1432 1221 1434 1233
rect 1458 1231 1459 1235
rect 1463 1231 1464 1235
rect 1479 1233 1483 1234
rect 1495 1238 1499 1239
rect 1495 1233 1499 1234
rect 1559 1238 1563 1239
rect 1559 1233 1563 1234
rect 1567 1238 1571 1239
rect 1567 1233 1571 1234
rect 1623 1238 1627 1239
rect 1623 1233 1627 1234
rect 1655 1238 1659 1239
rect 1672 1236 1674 1266
rect 1742 1260 1748 1261
rect 1742 1256 1743 1260
rect 1747 1256 1748 1260
rect 1742 1255 1748 1256
rect 1744 1239 1746 1255
rect 1768 1244 1770 1310
rect 1830 1300 1836 1301
rect 1830 1296 1831 1300
rect 1835 1296 1836 1300
rect 1830 1295 1836 1296
rect 1894 1300 1900 1301
rect 1894 1296 1895 1300
rect 1899 1296 1900 1300
rect 1894 1295 1900 1296
rect 1958 1300 1964 1301
rect 1958 1296 1959 1300
rect 1963 1296 1964 1300
rect 1958 1295 1964 1296
rect 2022 1300 2028 1301
rect 2022 1296 2023 1300
rect 2027 1296 2028 1300
rect 2022 1295 2028 1296
rect 1831 1294 1835 1295
rect 1831 1289 1835 1290
rect 1895 1294 1899 1295
rect 1895 1289 1899 1290
rect 1919 1294 1923 1295
rect 1919 1289 1923 1290
rect 1959 1294 1963 1295
rect 1959 1289 1963 1290
rect 2007 1294 2011 1295
rect 2007 1289 2011 1290
rect 2023 1294 2027 1295
rect 2023 1289 2027 1290
rect 1830 1288 1836 1289
rect 1830 1284 1831 1288
rect 1835 1284 1836 1288
rect 1830 1283 1836 1284
rect 1918 1288 1924 1289
rect 1918 1284 1919 1288
rect 1923 1284 1924 1288
rect 1918 1283 1924 1284
rect 2006 1288 2012 1289
rect 2006 1284 2007 1288
rect 2011 1284 2012 1288
rect 2006 1283 2012 1284
rect 2048 1272 2050 1330
rect 2072 1329 2074 1341
rect 2096 1336 2098 1370
rect 2118 1368 2119 1372
rect 2123 1368 2124 1372
rect 2118 1367 2124 1368
rect 2120 1347 2122 1367
rect 2119 1346 2123 1347
rect 2119 1341 2123 1342
rect 2094 1335 2100 1336
rect 2094 1331 2095 1335
rect 2099 1331 2100 1335
rect 2094 1330 2100 1331
rect 2070 1328 2076 1329
rect 2070 1324 2071 1328
rect 2075 1324 2076 1328
rect 2070 1323 2076 1324
rect 2120 1321 2122 1341
rect 2118 1320 2124 1321
rect 2118 1316 2119 1320
rect 2123 1316 2124 1320
rect 2094 1315 2100 1316
rect 2118 1315 2124 1316
rect 2094 1311 2095 1315
rect 2099 1311 2100 1315
rect 2094 1310 2100 1311
rect 2070 1300 2076 1301
rect 2070 1296 2071 1300
rect 2075 1296 2076 1300
rect 2070 1295 2076 1296
rect 2071 1294 2075 1295
rect 2071 1289 2075 1290
rect 2070 1288 2076 1289
rect 2070 1284 2071 1288
rect 2075 1284 2076 1288
rect 2070 1283 2076 1284
rect 2046 1271 2052 1272
rect 2046 1267 2047 1271
rect 2051 1267 2052 1271
rect 2046 1266 2052 1267
rect 1830 1260 1836 1261
rect 1830 1256 1831 1260
rect 1835 1256 1836 1260
rect 1830 1255 1836 1256
rect 1918 1260 1924 1261
rect 1918 1256 1919 1260
rect 1923 1256 1924 1260
rect 1918 1255 1924 1256
rect 2006 1260 2012 1261
rect 2006 1256 2007 1260
rect 2011 1256 2012 1260
rect 2006 1255 2012 1256
rect 2070 1260 2076 1261
rect 2070 1256 2071 1260
rect 2075 1256 2076 1260
rect 2070 1255 2076 1256
rect 1766 1243 1772 1244
rect 1766 1239 1767 1243
rect 1771 1239 1772 1243
rect 1832 1239 1834 1255
rect 1920 1239 1922 1255
rect 1994 1251 2000 1252
rect 1994 1247 1995 1251
rect 1999 1247 2000 1251
rect 1994 1246 2000 1247
rect 1679 1238 1683 1239
rect 1655 1233 1659 1234
rect 1670 1235 1676 1236
rect 1458 1230 1464 1231
rect 1430 1220 1436 1221
rect 1430 1216 1431 1220
rect 1435 1216 1436 1220
rect 1430 1215 1436 1216
rect 1460 1208 1462 1230
rect 1496 1221 1498 1233
rect 1560 1221 1562 1233
rect 1574 1227 1580 1228
rect 1574 1223 1575 1227
rect 1579 1223 1580 1227
rect 1574 1222 1580 1223
rect 1494 1220 1500 1221
rect 1494 1216 1495 1220
rect 1499 1216 1500 1220
rect 1494 1215 1500 1216
rect 1558 1220 1564 1221
rect 1558 1216 1559 1220
rect 1563 1216 1564 1220
rect 1558 1215 1564 1216
rect 1576 1208 1578 1222
rect 1624 1221 1626 1233
rect 1670 1231 1671 1235
rect 1675 1231 1676 1235
rect 1679 1233 1683 1234
rect 1735 1238 1739 1239
rect 1735 1233 1739 1234
rect 1743 1238 1747 1239
rect 1766 1238 1772 1239
rect 1791 1238 1795 1239
rect 1743 1233 1747 1234
rect 1791 1233 1795 1234
rect 1831 1238 1835 1239
rect 1831 1233 1835 1234
rect 1847 1238 1851 1239
rect 1847 1233 1851 1234
rect 1903 1238 1907 1239
rect 1903 1233 1907 1234
rect 1919 1238 1923 1239
rect 1919 1233 1923 1234
rect 1967 1238 1971 1239
rect 1967 1233 1971 1234
rect 1670 1230 1676 1231
rect 1680 1221 1682 1233
rect 1686 1227 1692 1228
rect 1686 1223 1687 1227
rect 1691 1223 1692 1227
rect 1686 1222 1692 1223
rect 1622 1220 1628 1221
rect 1622 1216 1623 1220
rect 1627 1216 1628 1220
rect 1622 1215 1628 1216
rect 1678 1220 1684 1221
rect 1678 1216 1679 1220
rect 1683 1216 1684 1220
rect 1678 1215 1684 1216
rect 1688 1208 1690 1222
rect 1736 1221 1738 1233
rect 1750 1227 1756 1228
rect 1750 1223 1751 1227
rect 1755 1223 1756 1227
rect 1750 1222 1756 1223
rect 1734 1220 1740 1221
rect 1734 1216 1735 1220
rect 1739 1216 1740 1220
rect 1734 1215 1740 1216
rect 1752 1208 1754 1222
rect 1792 1221 1794 1233
rect 1806 1227 1812 1228
rect 1806 1223 1807 1227
rect 1811 1223 1812 1227
rect 1806 1222 1812 1223
rect 1790 1220 1796 1221
rect 1790 1216 1791 1220
rect 1795 1216 1796 1220
rect 1790 1215 1796 1216
rect 1808 1208 1810 1222
rect 1848 1221 1850 1233
rect 1854 1227 1860 1228
rect 1854 1223 1855 1227
rect 1859 1223 1860 1227
rect 1854 1222 1860 1223
rect 1846 1220 1852 1221
rect 1846 1216 1847 1220
rect 1851 1216 1852 1220
rect 1846 1215 1852 1216
rect 1856 1208 1858 1222
rect 1904 1221 1906 1233
rect 1918 1227 1924 1228
rect 1918 1223 1919 1227
rect 1923 1223 1924 1227
rect 1918 1222 1924 1223
rect 1902 1220 1908 1221
rect 1902 1216 1903 1220
rect 1907 1216 1908 1220
rect 1902 1215 1908 1216
rect 1920 1208 1922 1222
rect 1968 1221 1970 1233
rect 1966 1220 1972 1221
rect 1966 1216 1967 1220
rect 1971 1216 1972 1220
rect 1966 1215 1972 1216
rect 1996 1208 1998 1246
rect 2008 1239 2010 1255
rect 2072 1239 2074 1255
rect 2096 1252 2098 1310
rect 2118 1303 2124 1304
rect 2118 1299 2119 1303
rect 2123 1299 2124 1303
rect 2118 1298 2124 1299
rect 2120 1295 2122 1298
rect 2119 1294 2123 1295
rect 2119 1289 2123 1290
rect 2120 1286 2122 1289
rect 2118 1285 2124 1286
rect 2118 1281 2119 1285
rect 2123 1281 2124 1285
rect 2118 1280 2124 1281
rect 2118 1268 2124 1269
rect 2118 1264 2119 1268
rect 2123 1264 2124 1268
rect 2118 1263 2124 1264
rect 2094 1251 2100 1252
rect 2094 1247 2095 1251
rect 2099 1247 2100 1251
rect 2094 1246 2100 1247
rect 2120 1239 2122 1263
rect 2007 1238 2011 1239
rect 2007 1233 2011 1234
rect 2031 1238 2035 1239
rect 2031 1233 2035 1234
rect 2071 1238 2075 1239
rect 2071 1233 2075 1234
rect 2119 1238 2123 1239
rect 2119 1233 2123 1234
rect 2006 1227 2012 1228
rect 2006 1223 2007 1227
rect 2011 1223 2012 1227
rect 2006 1222 2012 1223
rect 1134 1207 1140 1208
rect 1314 1207 1320 1208
rect 1094 1204 1100 1205
rect 1314 1203 1315 1207
rect 1319 1203 1320 1207
rect 1314 1202 1320 1203
rect 1342 1207 1348 1208
rect 1342 1203 1343 1207
rect 1347 1203 1348 1207
rect 1342 1202 1348 1203
rect 1390 1207 1396 1208
rect 1390 1203 1391 1207
rect 1395 1203 1396 1207
rect 1390 1202 1396 1203
rect 1458 1207 1464 1208
rect 1458 1203 1459 1207
rect 1463 1203 1464 1207
rect 1458 1202 1464 1203
rect 1514 1207 1520 1208
rect 1514 1203 1515 1207
rect 1519 1203 1520 1207
rect 1514 1202 1520 1203
rect 1574 1207 1580 1208
rect 1574 1203 1575 1207
rect 1579 1203 1580 1207
rect 1574 1202 1580 1203
rect 1670 1207 1676 1208
rect 1670 1203 1671 1207
rect 1675 1203 1676 1207
rect 1670 1202 1676 1203
rect 1686 1207 1692 1208
rect 1686 1203 1687 1207
rect 1691 1203 1692 1207
rect 1686 1202 1692 1203
rect 1750 1207 1756 1208
rect 1750 1203 1751 1207
rect 1755 1203 1756 1207
rect 1750 1202 1756 1203
rect 1806 1207 1812 1208
rect 1806 1203 1807 1207
rect 1811 1203 1812 1207
rect 1806 1202 1812 1203
rect 1854 1207 1860 1208
rect 1854 1203 1855 1207
rect 1859 1203 1860 1207
rect 1854 1202 1860 1203
rect 1918 1207 1924 1208
rect 1918 1203 1919 1207
rect 1923 1203 1924 1207
rect 1918 1202 1924 1203
rect 1994 1207 2000 1208
rect 1994 1203 1995 1207
rect 1999 1203 2000 1207
rect 1994 1202 2000 1203
rect 462 1195 468 1196
rect 462 1191 463 1195
rect 467 1191 468 1195
rect 462 1190 468 1191
rect 510 1195 516 1196
rect 510 1191 511 1195
rect 515 1191 516 1195
rect 510 1190 516 1191
rect 566 1195 572 1196
rect 566 1191 567 1195
rect 571 1191 572 1195
rect 566 1190 572 1191
rect 574 1195 580 1196
rect 574 1191 575 1195
rect 579 1191 580 1195
rect 574 1190 580 1191
rect 1006 1195 1012 1196
rect 1006 1191 1007 1195
rect 1011 1191 1012 1195
rect 1134 1195 1140 1196
rect 1006 1190 1012 1191
rect 1094 1192 1100 1193
rect 446 1184 452 1185
rect 446 1180 447 1184
rect 451 1180 452 1184
rect 446 1179 452 1180
rect 422 1175 428 1176
rect 422 1171 423 1175
rect 427 1171 428 1175
rect 422 1170 428 1171
rect 448 1163 450 1179
rect 464 1176 466 1190
rect 494 1184 500 1185
rect 494 1180 495 1184
rect 499 1180 500 1184
rect 494 1179 500 1180
rect 462 1175 468 1176
rect 462 1171 463 1175
rect 467 1171 468 1175
rect 462 1170 468 1171
rect 496 1163 498 1179
rect 512 1176 514 1190
rect 550 1184 556 1185
rect 550 1180 551 1184
rect 555 1180 556 1184
rect 550 1179 556 1180
rect 510 1175 516 1176
rect 510 1171 511 1175
rect 515 1171 516 1175
rect 510 1170 516 1171
rect 552 1163 554 1179
rect 111 1162 115 1163
rect 111 1157 115 1158
rect 271 1162 275 1163
rect 271 1157 275 1158
rect 311 1162 315 1163
rect 311 1157 315 1158
rect 351 1162 355 1163
rect 351 1157 355 1158
rect 399 1162 403 1163
rect 399 1157 403 1158
rect 439 1162 443 1163
rect 439 1157 443 1158
rect 447 1162 451 1163
rect 447 1157 451 1158
rect 479 1162 483 1163
rect 479 1157 483 1158
rect 495 1162 499 1163
rect 495 1157 499 1158
rect 527 1162 531 1163
rect 527 1157 531 1158
rect 551 1162 555 1163
rect 568 1160 570 1190
rect 1094 1188 1095 1192
rect 1099 1188 1100 1192
rect 1134 1191 1135 1195
rect 1139 1191 1140 1195
rect 1134 1190 1140 1191
rect 1286 1192 1292 1193
rect 1094 1187 1100 1188
rect 1136 1187 1138 1190
rect 1286 1188 1287 1192
rect 1291 1188 1292 1192
rect 1286 1187 1292 1188
rect 1326 1192 1332 1193
rect 1326 1188 1327 1192
rect 1331 1188 1332 1192
rect 1326 1187 1332 1188
rect 1374 1192 1380 1193
rect 1374 1188 1375 1192
rect 1379 1188 1380 1192
rect 1374 1187 1380 1188
rect 1430 1192 1436 1193
rect 1430 1188 1431 1192
rect 1435 1188 1436 1192
rect 1430 1187 1436 1188
rect 1494 1192 1500 1193
rect 1494 1188 1495 1192
rect 1499 1188 1500 1192
rect 1494 1187 1500 1188
rect 606 1184 612 1185
rect 606 1180 607 1184
rect 611 1180 612 1184
rect 606 1179 612 1180
rect 670 1184 676 1185
rect 670 1180 671 1184
rect 675 1180 676 1184
rect 670 1179 676 1180
rect 742 1184 748 1185
rect 742 1180 743 1184
rect 747 1180 748 1184
rect 742 1179 748 1180
rect 814 1184 820 1185
rect 814 1180 815 1184
rect 819 1180 820 1184
rect 814 1179 820 1180
rect 894 1184 900 1185
rect 894 1180 895 1184
rect 899 1180 900 1184
rect 894 1179 900 1180
rect 982 1184 988 1185
rect 982 1180 983 1184
rect 987 1180 988 1184
rect 982 1179 988 1180
rect 608 1163 610 1179
rect 672 1163 674 1179
rect 698 1167 704 1168
rect 698 1163 699 1167
rect 703 1163 704 1167
rect 744 1163 746 1179
rect 816 1163 818 1179
rect 896 1163 898 1179
rect 970 1175 976 1176
rect 970 1171 971 1175
rect 975 1171 976 1175
rect 970 1170 976 1171
rect 575 1162 579 1163
rect 551 1157 555 1158
rect 566 1159 572 1160
rect 112 1137 114 1157
rect 400 1145 402 1157
rect 440 1145 442 1157
rect 454 1151 460 1152
rect 454 1147 455 1151
rect 459 1147 460 1151
rect 454 1146 460 1147
rect 398 1144 404 1145
rect 398 1140 399 1144
rect 403 1140 404 1144
rect 398 1139 404 1140
rect 438 1144 444 1145
rect 438 1140 439 1144
rect 443 1140 444 1144
rect 438 1139 444 1140
rect 110 1136 116 1137
rect 110 1132 111 1136
rect 115 1132 116 1136
rect 456 1132 458 1146
rect 480 1145 482 1157
rect 494 1151 500 1152
rect 494 1147 495 1151
rect 499 1147 500 1151
rect 494 1146 500 1147
rect 478 1144 484 1145
rect 478 1140 479 1144
rect 483 1140 484 1144
rect 478 1139 484 1140
rect 496 1132 498 1146
rect 528 1145 530 1157
rect 566 1155 567 1159
rect 571 1155 572 1159
rect 575 1157 579 1158
rect 607 1162 611 1163
rect 607 1157 611 1158
rect 623 1162 627 1163
rect 671 1162 675 1163
rect 698 1162 704 1163
rect 719 1162 723 1163
rect 623 1157 627 1158
rect 662 1159 668 1160
rect 566 1154 572 1155
rect 542 1151 548 1152
rect 542 1147 543 1151
rect 547 1147 548 1151
rect 542 1146 548 1147
rect 526 1144 532 1145
rect 526 1140 527 1144
rect 531 1140 532 1144
rect 526 1139 532 1140
rect 544 1132 546 1146
rect 576 1145 578 1157
rect 590 1151 596 1152
rect 590 1147 591 1151
rect 595 1147 596 1151
rect 590 1146 596 1147
rect 574 1144 580 1145
rect 574 1140 575 1144
rect 579 1140 580 1144
rect 574 1139 580 1140
rect 592 1132 594 1146
rect 624 1145 626 1157
rect 662 1155 663 1159
rect 667 1155 668 1159
rect 671 1157 675 1158
rect 662 1154 668 1155
rect 630 1151 636 1152
rect 630 1147 631 1151
rect 635 1147 636 1151
rect 630 1146 636 1147
rect 622 1144 628 1145
rect 622 1140 623 1144
rect 627 1140 628 1144
rect 622 1139 628 1140
rect 632 1132 634 1146
rect 110 1131 116 1132
rect 426 1131 432 1132
rect 426 1127 427 1131
rect 431 1127 432 1131
rect 426 1126 432 1127
rect 454 1131 460 1132
rect 454 1127 455 1131
rect 459 1127 460 1131
rect 454 1126 460 1127
rect 494 1131 500 1132
rect 494 1127 495 1131
rect 499 1127 500 1131
rect 494 1126 500 1127
rect 542 1131 548 1132
rect 542 1127 543 1131
rect 547 1127 548 1131
rect 542 1126 548 1127
rect 590 1131 596 1132
rect 590 1127 591 1131
rect 595 1127 596 1131
rect 590 1126 596 1127
rect 630 1131 636 1132
rect 630 1127 631 1131
rect 635 1127 636 1131
rect 630 1126 636 1127
rect 110 1119 116 1120
rect 110 1115 111 1119
rect 115 1115 116 1119
rect 110 1114 116 1115
rect 398 1116 404 1117
rect 112 1111 114 1114
rect 398 1112 399 1116
rect 403 1112 404 1116
rect 398 1111 404 1112
rect 111 1110 115 1111
rect 111 1105 115 1106
rect 159 1110 163 1111
rect 159 1105 163 1106
rect 199 1110 203 1111
rect 199 1105 203 1106
rect 255 1110 259 1111
rect 255 1105 259 1106
rect 319 1110 323 1111
rect 319 1105 323 1106
rect 399 1110 403 1111
rect 399 1105 403 1106
rect 112 1102 114 1105
rect 158 1104 164 1105
rect 110 1101 116 1102
rect 110 1097 111 1101
rect 115 1097 116 1101
rect 158 1100 159 1104
rect 163 1100 164 1104
rect 158 1099 164 1100
rect 198 1104 204 1105
rect 198 1100 199 1104
rect 203 1100 204 1104
rect 198 1099 204 1100
rect 254 1104 260 1105
rect 254 1100 255 1104
rect 259 1100 260 1104
rect 254 1099 260 1100
rect 318 1104 324 1105
rect 318 1100 319 1104
rect 323 1100 324 1104
rect 318 1099 324 1100
rect 398 1104 404 1105
rect 398 1100 399 1104
rect 403 1100 404 1104
rect 398 1099 404 1100
rect 110 1096 116 1097
rect 186 1087 192 1088
rect 110 1084 116 1085
rect 110 1080 111 1084
rect 115 1080 116 1084
rect 186 1083 187 1087
rect 191 1083 192 1087
rect 186 1082 192 1083
rect 206 1087 212 1088
rect 206 1083 207 1087
rect 211 1083 212 1087
rect 206 1082 212 1083
rect 110 1079 116 1080
rect 112 1055 114 1079
rect 158 1076 164 1077
rect 158 1072 159 1076
rect 163 1072 164 1076
rect 158 1071 164 1072
rect 160 1055 162 1071
rect 166 1059 172 1060
rect 166 1055 167 1059
rect 171 1055 172 1059
rect 111 1054 115 1055
rect 111 1049 115 1050
rect 135 1054 139 1055
rect 135 1049 139 1050
rect 159 1054 163 1055
rect 166 1054 172 1055
rect 175 1054 179 1055
rect 159 1049 163 1050
rect 112 1029 114 1049
rect 136 1037 138 1049
rect 134 1036 140 1037
rect 134 1032 135 1036
rect 139 1032 140 1036
rect 134 1031 140 1032
rect 110 1028 116 1029
rect 110 1024 111 1028
rect 115 1024 116 1028
rect 110 1023 116 1024
rect 159 1023 165 1024
rect 159 1019 160 1023
rect 164 1022 165 1023
rect 168 1022 170 1054
rect 188 1052 190 1082
rect 198 1076 204 1077
rect 198 1072 199 1076
rect 203 1072 204 1076
rect 198 1071 204 1072
rect 200 1055 202 1071
rect 208 1068 210 1082
rect 254 1076 260 1077
rect 254 1072 255 1076
rect 259 1072 260 1076
rect 254 1071 260 1072
rect 318 1076 324 1077
rect 318 1072 319 1076
rect 323 1072 324 1076
rect 318 1071 324 1072
rect 398 1076 404 1077
rect 398 1072 399 1076
rect 403 1072 404 1076
rect 398 1071 404 1072
rect 206 1067 212 1068
rect 206 1063 207 1067
rect 211 1063 212 1067
rect 206 1062 212 1063
rect 256 1055 258 1071
rect 320 1055 322 1071
rect 400 1055 402 1071
rect 428 1060 430 1126
rect 438 1116 444 1117
rect 438 1112 439 1116
rect 443 1112 444 1116
rect 438 1111 444 1112
rect 478 1116 484 1117
rect 478 1112 479 1116
rect 483 1112 484 1116
rect 478 1111 484 1112
rect 526 1116 532 1117
rect 526 1112 527 1116
rect 531 1112 532 1116
rect 526 1111 532 1112
rect 574 1116 580 1117
rect 574 1112 575 1116
rect 579 1112 580 1116
rect 574 1111 580 1112
rect 622 1116 628 1117
rect 622 1112 623 1116
rect 627 1112 628 1116
rect 622 1111 628 1112
rect 439 1110 443 1111
rect 439 1105 443 1106
rect 479 1110 483 1111
rect 479 1105 483 1106
rect 527 1110 531 1111
rect 527 1105 531 1106
rect 559 1110 563 1111
rect 559 1105 563 1106
rect 575 1110 579 1111
rect 575 1105 579 1106
rect 623 1110 627 1111
rect 623 1105 627 1106
rect 639 1110 643 1111
rect 639 1105 643 1106
rect 478 1104 484 1105
rect 478 1100 479 1104
rect 483 1100 484 1104
rect 478 1099 484 1100
rect 558 1104 564 1105
rect 558 1100 559 1104
rect 563 1100 564 1104
rect 558 1099 564 1100
rect 638 1104 644 1105
rect 638 1100 639 1104
rect 643 1100 644 1104
rect 638 1099 644 1100
rect 664 1088 666 1154
rect 672 1145 674 1157
rect 670 1144 676 1145
rect 670 1140 671 1144
rect 675 1140 676 1144
rect 670 1139 676 1140
rect 700 1132 702 1162
rect 719 1157 723 1158
rect 743 1162 747 1163
rect 743 1157 747 1158
rect 775 1162 779 1163
rect 775 1157 779 1158
rect 815 1162 819 1163
rect 815 1157 819 1158
rect 831 1162 835 1163
rect 831 1157 835 1158
rect 887 1162 891 1163
rect 887 1157 891 1158
rect 895 1162 899 1163
rect 895 1157 899 1158
rect 943 1162 947 1163
rect 943 1157 947 1158
rect 720 1145 722 1157
rect 734 1151 740 1152
rect 734 1147 735 1151
rect 739 1147 740 1151
rect 734 1146 740 1147
rect 718 1144 724 1145
rect 718 1140 719 1144
rect 723 1140 724 1144
rect 718 1139 724 1140
rect 736 1132 738 1146
rect 776 1145 778 1157
rect 790 1151 796 1152
rect 790 1147 791 1151
rect 795 1147 796 1151
rect 790 1146 796 1147
rect 774 1144 780 1145
rect 774 1140 775 1144
rect 779 1140 780 1144
rect 774 1139 780 1140
rect 792 1132 794 1146
rect 832 1145 834 1157
rect 846 1151 852 1152
rect 846 1147 847 1151
rect 851 1147 852 1151
rect 846 1146 852 1147
rect 830 1144 836 1145
rect 830 1140 831 1144
rect 835 1140 836 1144
rect 830 1139 836 1140
rect 848 1132 850 1146
rect 888 1145 890 1157
rect 902 1151 908 1152
rect 902 1147 903 1151
rect 907 1147 908 1151
rect 902 1146 908 1147
rect 886 1144 892 1145
rect 886 1140 887 1144
rect 891 1140 892 1144
rect 886 1139 892 1140
rect 904 1132 906 1146
rect 944 1145 946 1157
rect 942 1144 948 1145
rect 942 1140 943 1144
rect 947 1140 948 1144
rect 942 1139 948 1140
rect 972 1132 974 1170
rect 984 1163 986 1179
rect 1096 1163 1098 1187
rect 1135 1186 1139 1187
rect 1135 1181 1139 1182
rect 1159 1186 1163 1187
rect 1159 1181 1163 1182
rect 1207 1186 1211 1187
rect 1207 1181 1211 1182
rect 1279 1186 1283 1187
rect 1279 1181 1283 1182
rect 1287 1186 1291 1187
rect 1287 1181 1291 1182
rect 1327 1186 1331 1187
rect 1327 1181 1331 1182
rect 1351 1186 1355 1187
rect 1351 1181 1355 1182
rect 1375 1186 1379 1187
rect 1375 1181 1379 1182
rect 1423 1186 1427 1187
rect 1423 1181 1427 1182
rect 1431 1186 1435 1187
rect 1431 1181 1435 1182
rect 1487 1186 1491 1187
rect 1487 1181 1491 1182
rect 1495 1186 1499 1187
rect 1495 1181 1499 1182
rect 1136 1178 1138 1181
rect 1158 1180 1164 1181
rect 1134 1177 1140 1178
rect 1134 1173 1135 1177
rect 1139 1173 1140 1177
rect 1158 1176 1159 1180
rect 1163 1176 1164 1180
rect 1158 1175 1164 1176
rect 1206 1180 1212 1181
rect 1206 1176 1207 1180
rect 1211 1176 1212 1180
rect 1206 1175 1212 1176
rect 1278 1180 1284 1181
rect 1278 1176 1279 1180
rect 1283 1176 1284 1180
rect 1278 1175 1284 1176
rect 1350 1180 1356 1181
rect 1350 1176 1351 1180
rect 1355 1176 1356 1180
rect 1350 1175 1356 1176
rect 1422 1180 1428 1181
rect 1422 1176 1423 1180
rect 1427 1176 1428 1180
rect 1422 1175 1428 1176
rect 1486 1180 1492 1181
rect 1486 1176 1487 1180
rect 1491 1176 1492 1180
rect 1486 1175 1492 1176
rect 1134 1172 1140 1173
rect 1370 1163 1376 1164
rect 983 1162 987 1163
rect 983 1157 987 1158
rect 1007 1162 1011 1163
rect 1007 1157 1011 1158
rect 1047 1162 1051 1163
rect 1047 1157 1051 1158
rect 1095 1162 1099 1163
rect 1095 1157 1099 1158
rect 1134 1160 1140 1161
rect 1008 1145 1010 1157
rect 1022 1151 1028 1152
rect 1022 1147 1023 1151
rect 1027 1147 1028 1151
rect 1022 1146 1028 1147
rect 1006 1144 1012 1145
rect 1006 1140 1007 1144
rect 1011 1140 1012 1144
rect 1006 1139 1012 1140
rect 698 1131 704 1132
rect 698 1127 699 1131
rect 703 1127 704 1131
rect 698 1126 704 1127
rect 734 1131 740 1132
rect 734 1127 735 1131
rect 739 1127 740 1131
rect 734 1126 740 1127
rect 790 1131 796 1132
rect 790 1127 791 1131
rect 795 1127 796 1131
rect 790 1126 796 1127
rect 846 1131 852 1132
rect 846 1127 847 1131
rect 851 1127 852 1131
rect 846 1126 852 1127
rect 902 1131 908 1132
rect 902 1127 903 1131
rect 907 1127 908 1131
rect 902 1126 908 1127
rect 970 1131 976 1132
rect 970 1127 971 1131
rect 975 1127 976 1131
rect 970 1126 976 1127
rect 670 1116 676 1117
rect 670 1112 671 1116
rect 675 1112 676 1116
rect 670 1111 676 1112
rect 718 1116 724 1117
rect 718 1112 719 1116
rect 723 1112 724 1116
rect 718 1111 724 1112
rect 774 1116 780 1117
rect 774 1112 775 1116
rect 779 1112 780 1116
rect 774 1111 780 1112
rect 830 1116 836 1117
rect 830 1112 831 1116
rect 835 1112 836 1116
rect 830 1111 836 1112
rect 886 1116 892 1117
rect 886 1112 887 1116
rect 891 1112 892 1116
rect 886 1111 892 1112
rect 942 1116 948 1117
rect 942 1112 943 1116
rect 947 1112 948 1116
rect 942 1111 948 1112
rect 1006 1116 1012 1117
rect 1006 1112 1007 1116
rect 1011 1112 1012 1116
rect 1006 1111 1012 1112
rect 671 1110 675 1111
rect 671 1105 675 1106
rect 711 1110 715 1111
rect 711 1105 715 1106
rect 719 1110 723 1111
rect 719 1105 723 1106
rect 775 1110 779 1111
rect 775 1105 779 1106
rect 783 1110 787 1111
rect 783 1105 787 1106
rect 831 1110 835 1111
rect 831 1105 835 1106
rect 855 1110 859 1111
rect 855 1105 859 1106
rect 887 1110 891 1111
rect 887 1105 891 1106
rect 927 1110 931 1111
rect 927 1105 931 1106
rect 943 1110 947 1111
rect 943 1105 947 1106
rect 999 1110 1003 1111
rect 999 1105 1003 1106
rect 1007 1110 1011 1111
rect 1007 1105 1011 1106
rect 710 1104 716 1105
rect 710 1100 711 1104
rect 715 1100 716 1104
rect 710 1099 716 1100
rect 782 1104 788 1105
rect 782 1100 783 1104
rect 787 1100 788 1104
rect 782 1099 788 1100
rect 854 1104 860 1105
rect 854 1100 855 1104
rect 859 1100 860 1104
rect 854 1099 860 1100
rect 926 1104 932 1105
rect 926 1100 927 1104
rect 931 1100 932 1104
rect 926 1099 932 1100
rect 998 1104 1004 1105
rect 998 1100 999 1104
rect 1003 1100 1004 1104
rect 998 1099 1004 1100
rect 1024 1088 1026 1146
rect 1048 1145 1050 1157
rect 1062 1151 1068 1152
rect 1062 1147 1063 1151
rect 1067 1147 1068 1151
rect 1062 1146 1068 1147
rect 1046 1144 1052 1145
rect 1046 1140 1047 1144
rect 1051 1140 1052 1144
rect 1046 1139 1052 1140
rect 1064 1132 1066 1146
rect 1096 1137 1098 1157
rect 1134 1156 1135 1160
rect 1139 1156 1140 1160
rect 1370 1159 1371 1163
rect 1375 1159 1376 1163
rect 1370 1158 1376 1159
rect 1134 1155 1140 1156
rect 1094 1136 1100 1137
rect 1094 1132 1095 1136
rect 1099 1132 1100 1136
rect 1054 1131 1060 1132
rect 1054 1127 1055 1131
rect 1059 1127 1060 1131
rect 1054 1126 1060 1127
rect 1062 1131 1068 1132
rect 1094 1131 1100 1132
rect 1136 1131 1138 1155
rect 1158 1152 1164 1153
rect 1158 1148 1159 1152
rect 1163 1148 1164 1152
rect 1158 1147 1164 1148
rect 1206 1152 1212 1153
rect 1206 1148 1207 1152
rect 1211 1148 1212 1152
rect 1206 1147 1212 1148
rect 1278 1152 1284 1153
rect 1278 1148 1279 1152
rect 1283 1148 1284 1152
rect 1278 1147 1284 1148
rect 1350 1152 1356 1153
rect 1350 1148 1351 1152
rect 1355 1148 1356 1152
rect 1350 1147 1356 1148
rect 1160 1131 1162 1147
rect 1208 1131 1210 1147
rect 1280 1131 1282 1147
rect 1352 1131 1354 1147
rect 1062 1127 1063 1131
rect 1067 1127 1068 1131
rect 1062 1126 1068 1127
rect 1135 1130 1139 1131
rect 1046 1116 1052 1117
rect 1046 1112 1047 1116
rect 1051 1112 1052 1116
rect 1046 1111 1052 1112
rect 1047 1110 1051 1111
rect 1047 1105 1051 1106
rect 1046 1104 1052 1105
rect 1046 1100 1047 1104
rect 1051 1100 1052 1104
rect 1046 1099 1052 1100
rect 662 1087 668 1088
rect 662 1083 663 1087
rect 667 1083 668 1087
rect 662 1082 668 1083
rect 1014 1087 1020 1088
rect 1014 1083 1015 1087
rect 1019 1083 1020 1087
rect 1014 1082 1020 1083
rect 1022 1087 1028 1088
rect 1022 1083 1023 1087
rect 1027 1083 1028 1087
rect 1022 1082 1028 1083
rect 478 1076 484 1077
rect 478 1072 479 1076
rect 483 1072 484 1076
rect 478 1071 484 1072
rect 558 1076 564 1077
rect 558 1072 559 1076
rect 563 1072 564 1076
rect 558 1071 564 1072
rect 638 1076 644 1077
rect 638 1072 639 1076
rect 643 1072 644 1076
rect 638 1071 644 1072
rect 710 1076 716 1077
rect 710 1072 711 1076
rect 715 1072 716 1076
rect 710 1071 716 1072
rect 782 1076 788 1077
rect 782 1072 783 1076
rect 787 1072 788 1076
rect 782 1071 788 1072
rect 854 1076 860 1077
rect 854 1072 855 1076
rect 859 1072 860 1076
rect 854 1071 860 1072
rect 926 1076 932 1077
rect 926 1072 927 1076
rect 931 1072 932 1076
rect 926 1071 932 1072
rect 998 1076 1004 1077
rect 998 1072 999 1076
rect 1003 1072 1004 1076
rect 998 1071 1004 1072
rect 426 1059 432 1060
rect 426 1055 427 1059
rect 431 1055 432 1059
rect 480 1055 482 1071
rect 560 1055 562 1071
rect 602 1059 608 1060
rect 602 1055 603 1059
rect 607 1055 608 1059
rect 640 1055 642 1071
rect 712 1055 714 1071
rect 784 1055 786 1071
rect 856 1055 858 1071
rect 882 1067 888 1068
rect 882 1063 883 1067
rect 887 1063 888 1067
rect 882 1062 888 1063
rect 199 1054 203 1055
rect 175 1049 179 1050
rect 186 1051 192 1052
rect 176 1037 178 1049
rect 186 1047 187 1051
rect 191 1047 192 1051
rect 199 1049 203 1050
rect 215 1054 219 1055
rect 215 1049 219 1050
rect 255 1054 259 1055
rect 255 1049 259 1050
rect 319 1054 323 1055
rect 319 1049 323 1050
rect 383 1054 387 1055
rect 383 1049 387 1050
rect 399 1054 403 1055
rect 426 1054 432 1055
rect 447 1054 451 1055
rect 399 1049 403 1050
rect 447 1049 451 1050
rect 479 1054 483 1055
rect 479 1049 483 1050
rect 511 1054 515 1055
rect 511 1049 515 1050
rect 559 1054 563 1055
rect 559 1049 563 1050
rect 575 1054 579 1055
rect 602 1054 608 1055
rect 631 1054 635 1055
rect 575 1049 579 1050
rect 186 1046 192 1047
rect 190 1043 196 1044
rect 190 1039 191 1043
rect 195 1039 196 1043
rect 190 1038 196 1039
rect 174 1036 180 1037
rect 174 1032 175 1036
rect 179 1032 180 1036
rect 174 1031 180 1032
rect 192 1024 194 1038
rect 216 1037 218 1049
rect 230 1043 236 1044
rect 230 1039 231 1043
rect 235 1039 236 1043
rect 230 1038 236 1039
rect 214 1036 220 1037
rect 214 1032 215 1036
rect 219 1032 220 1036
rect 214 1031 220 1032
rect 232 1024 234 1038
rect 256 1037 258 1049
rect 270 1043 276 1044
rect 270 1039 271 1043
rect 275 1039 276 1043
rect 270 1038 276 1039
rect 254 1036 260 1037
rect 254 1032 255 1036
rect 259 1032 260 1036
rect 254 1031 260 1032
rect 272 1024 274 1038
rect 320 1037 322 1049
rect 384 1037 386 1049
rect 398 1043 404 1044
rect 398 1039 399 1043
rect 403 1039 404 1043
rect 398 1038 404 1039
rect 318 1036 324 1037
rect 318 1032 319 1036
rect 323 1032 324 1036
rect 318 1031 324 1032
rect 382 1036 388 1037
rect 382 1032 383 1036
rect 387 1032 388 1036
rect 382 1031 388 1032
rect 400 1024 402 1038
rect 448 1037 450 1049
rect 462 1043 468 1044
rect 462 1039 463 1043
rect 467 1039 468 1043
rect 462 1038 468 1039
rect 446 1036 452 1037
rect 446 1032 447 1036
rect 451 1032 452 1036
rect 446 1031 452 1032
rect 464 1024 466 1038
rect 512 1037 514 1049
rect 546 1043 552 1044
rect 546 1039 547 1043
rect 551 1039 552 1043
rect 546 1038 552 1039
rect 554 1043 560 1044
rect 554 1039 555 1043
rect 559 1039 560 1043
rect 554 1038 560 1039
rect 510 1036 516 1037
rect 510 1032 511 1036
rect 515 1032 516 1036
rect 510 1031 516 1032
rect 164 1020 170 1022
rect 190 1023 196 1024
rect 164 1019 165 1020
rect 159 1018 165 1019
rect 190 1019 191 1023
rect 195 1019 196 1023
rect 190 1018 196 1019
rect 230 1023 236 1024
rect 230 1019 231 1023
rect 235 1019 236 1023
rect 230 1018 236 1019
rect 270 1023 276 1024
rect 270 1019 271 1023
rect 275 1019 276 1023
rect 270 1018 276 1019
rect 290 1023 296 1024
rect 290 1019 291 1023
rect 295 1019 296 1023
rect 290 1018 296 1019
rect 398 1023 404 1024
rect 398 1019 399 1023
rect 403 1019 404 1023
rect 398 1018 404 1019
rect 462 1023 468 1024
rect 462 1019 463 1023
rect 467 1019 468 1023
rect 462 1018 468 1019
rect 110 1011 116 1012
rect 110 1007 111 1011
rect 115 1007 116 1011
rect 110 1006 116 1007
rect 134 1008 140 1009
rect 112 999 114 1006
rect 134 1004 135 1008
rect 139 1004 140 1008
rect 134 1003 140 1004
rect 174 1008 180 1009
rect 174 1004 175 1008
rect 179 1004 180 1008
rect 174 1003 180 1004
rect 214 1008 220 1009
rect 214 1004 215 1008
rect 219 1004 220 1008
rect 214 1003 220 1004
rect 254 1008 260 1009
rect 254 1004 255 1008
rect 259 1004 260 1008
rect 254 1003 260 1004
rect 136 999 138 1003
rect 176 999 178 1003
rect 216 999 218 1003
rect 256 999 258 1003
rect 111 998 115 999
rect 111 993 115 994
rect 135 998 139 999
rect 135 993 139 994
rect 175 998 179 999
rect 175 993 179 994
rect 215 998 219 999
rect 215 993 219 994
rect 223 998 227 999
rect 223 993 227 994
rect 255 998 259 999
rect 255 993 259 994
rect 279 998 283 999
rect 279 993 283 994
rect 112 990 114 993
rect 134 992 140 993
rect 110 989 116 990
rect 110 985 111 989
rect 115 985 116 989
rect 134 988 135 992
rect 139 988 140 992
rect 134 987 140 988
rect 174 992 180 993
rect 174 988 175 992
rect 179 988 180 992
rect 174 987 180 988
rect 222 992 228 993
rect 222 988 223 992
rect 227 988 228 992
rect 222 987 228 988
rect 278 992 284 993
rect 278 988 279 992
rect 283 988 284 992
rect 278 987 284 988
rect 110 984 116 985
rect 182 975 188 976
rect 110 972 116 973
rect 110 968 111 972
rect 115 968 116 972
rect 182 971 183 975
rect 187 971 188 975
rect 182 970 188 971
rect 110 967 116 968
rect 112 943 114 967
rect 134 964 140 965
rect 134 960 135 964
rect 139 960 140 964
rect 134 959 140 960
rect 174 964 180 965
rect 174 960 175 964
rect 179 960 180 964
rect 174 959 180 960
rect 136 943 138 959
rect 176 943 178 959
rect 184 956 186 970
rect 222 964 228 965
rect 222 960 223 964
rect 227 960 228 964
rect 222 959 228 960
rect 278 964 284 965
rect 278 960 279 964
rect 283 960 284 964
rect 278 959 284 960
rect 182 955 188 956
rect 182 951 183 955
rect 187 951 188 955
rect 182 950 188 951
rect 224 943 226 959
rect 280 943 282 959
rect 292 956 294 1018
rect 318 1008 324 1009
rect 318 1004 319 1008
rect 323 1004 324 1008
rect 318 1003 324 1004
rect 382 1008 388 1009
rect 382 1004 383 1008
rect 387 1004 388 1008
rect 382 1003 388 1004
rect 446 1008 452 1009
rect 446 1004 447 1008
rect 451 1004 452 1008
rect 446 1003 452 1004
rect 510 1008 516 1009
rect 510 1004 511 1008
rect 515 1004 516 1008
rect 510 1003 516 1004
rect 320 999 322 1003
rect 384 999 386 1003
rect 448 999 450 1003
rect 512 999 514 1003
rect 319 998 323 999
rect 319 993 323 994
rect 343 998 347 999
rect 343 993 347 994
rect 383 998 387 999
rect 383 993 387 994
rect 407 998 411 999
rect 407 993 411 994
rect 447 998 451 999
rect 447 993 451 994
rect 471 998 475 999
rect 471 993 475 994
rect 511 998 515 999
rect 511 993 515 994
rect 527 998 531 999
rect 527 993 531 994
rect 342 992 348 993
rect 342 988 343 992
rect 347 988 348 992
rect 342 987 348 988
rect 406 992 412 993
rect 406 988 407 992
rect 411 988 412 992
rect 406 987 412 988
rect 470 992 476 993
rect 470 988 471 992
rect 475 988 476 992
rect 470 987 476 988
rect 526 992 532 993
rect 526 988 527 992
rect 531 988 532 992
rect 526 987 532 988
rect 302 983 308 984
rect 302 979 303 983
rect 307 979 308 983
rect 302 978 308 979
rect 304 956 306 978
rect 548 976 550 1038
rect 556 1024 558 1038
rect 576 1037 578 1049
rect 574 1036 580 1037
rect 574 1032 575 1036
rect 579 1032 580 1036
rect 574 1031 580 1032
rect 604 1024 606 1054
rect 631 1049 635 1050
rect 639 1054 643 1055
rect 639 1049 643 1050
rect 687 1054 691 1055
rect 687 1049 691 1050
rect 711 1054 715 1055
rect 711 1049 715 1050
rect 743 1054 747 1055
rect 743 1049 747 1050
rect 783 1054 787 1055
rect 783 1049 787 1050
rect 799 1054 803 1055
rect 799 1049 803 1050
rect 855 1054 859 1055
rect 855 1049 859 1050
rect 863 1054 867 1055
rect 863 1049 867 1050
rect 610 1043 616 1044
rect 610 1039 611 1043
rect 615 1039 616 1043
rect 610 1038 616 1039
rect 554 1023 560 1024
rect 554 1019 555 1023
rect 559 1019 560 1023
rect 554 1018 560 1019
rect 602 1023 608 1024
rect 602 1019 603 1023
rect 607 1019 608 1023
rect 602 1018 608 1019
rect 574 1008 580 1009
rect 574 1004 575 1008
rect 579 1004 580 1008
rect 574 1003 580 1004
rect 576 999 578 1003
rect 575 998 579 999
rect 575 993 579 994
rect 583 998 587 999
rect 583 993 587 994
rect 582 992 588 993
rect 582 988 583 992
rect 587 988 588 992
rect 582 987 588 988
rect 612 987 614 1038
rect 632 1037 634 1049
rect 688 1037 690 1049
rect 734 1043 740 1044
rect 734 1039 735 1043
rect 739 1039 740 1043
rect 734 1038 740 1039
rect 630 1036 636 1037
rect 630 1032 631 1036
rect 635 1032 636 1036
rect 630 1031 636 1032
rect 686 1036 692 1037
rect 686 1032 687 1036
rect 691 1032 692 1036
rect 686 1031 692 1032
rect 736 1024 738 1038
rect 744 1037 746 1049
rect 800 1037 802 1049
rect 864 1037 866 1049
rect 742 1036 748 1037
rect 742 1032 743 1036
rect 747 1032 748 1036
rect 742 1031 748 1032
rect 798 1036 804 1037
rect 798 1032 799 1036
rect 803 1032 804 1036
rect 798 1031 804 1032
rect 862 1036 868 1037
rect 862 1032 863 1036
rect 867 1032 868 1036
rect 862 1031 868 1032
rect 884 1024 886 1062
rect 928 1055 930 1071
rect 1000 1055 1002 1071
rect 1016 1068 1018 1082
rect 1046 1076 1052 1077
rect 1046 1072 1047 1076
rect 1051 1072 1052 1076
rect 1046 1071 1052 1072
rect 1014 1067 1020 1068
rect 1014 1063 1015 1067
rect 1019 1063 1020 1067
rect 1014 1062 1020 1063
rect 1048 1055 1050 1071
rect 1056 1068 1058 1126
rect 1135 1125 1139 1126
rect 1159 1130 1163 1131
rect 1159 1125 1163 1126
rect 1191 1130 1195 1131
rect 1191 1125 1195 1126
rect 1207 1130 1211 1131
rect 1207 1125 1211 1126
rect 1271 1130 1275 1131
rect 1271 1125 1275 1126
rect 1279 1130 1283 1131
rect 1279 1125 1283 1126
rect 1343 1130 1347 1131
rect 1343 1125 1347 1126
rect 1351 1130 1355 1131
rect 1351 1125 1355 1126
rect 1094 1119 1100 1120
rect 1094 1115 1095 1119
rect 1099 1115 1100 1119
rect 1094 1114 1100 1115
rect 1096 1111 1098 1114
rect 1095 1110 1099 1111
rect 1095 1105 1099 1106
rect 1136 1105 1138 1125
rect 1192 1113 1194 1125
rect 1272 1113 1274 1125
rect 1286 1119 1292 1120
rect 1286 1115 1287 1119
rect 1291 1115 1292 1119
rect 1286 1114 1292 1115
rect 1326 1119 1332 1120
rect 1326 1115 1327 1119
rect 1331 1115 1332 1119
rect 1326 1114 1332 1115
rect 1190 1112 1196 1113
rect 1190 1108 1191 1112
rect 1195 1108 1196 1112
rect 1190 1107 1196 1108
rect 1270 1112 1276 1113
rect 1270 1108 1271 1112
rect 1275 1108 1276 1112
rect 1270 1107 1276 1108
rect 1096 1102 1098 1105
rect 1134 1104 1140 1105
rect 1094 1101 1100 1102
rect 1094 1097 1095 1101
rect 1099 1097 1100 1101
rect 1134 1100 1135 1104
rect 1139 1100 1140 1104
rect 1288 1100 1290 1114
rect 1134 1099 1140 1100
rect 1286 1099 1292 1100
rect 1094 1096 1100 1097
rect 1286 1095 1287 1099
rect 1291 1095 1292 1099
rect 1286 1094 1292 1095
rect 1086 1087 1092 1088
rect 1086 1083 1087 1087
rect 1091 1083 1092 1087
rect 1134 1087 1140 1088
rect 1086 1082 1092 1083
rect 1094 1084 1100 1085
rect 1054 1067 1060 1068
rect 1054 1063 1055 1067
rect 1059 1063 1060 1067
rect 1054 1062 1060 1063
rect 927 1054 931 1055
rect 927 1049 931 1050
rect 999 1054 1003 1055
rect 999 1049 1003 1050
rect 1047 1054 1051 1055
rect 1047 1049 1051 1050
rect 1088 1036 1090 1082
rect 1094 1080 1095 1084
rect 1099 1080 1100 1084
rect 1134 1083 1135 1087
rect 1139 1083 1140 1087
rect 1134 1082 1140 1083
rect 1190 1084 1196 1085
rect 1094 1079 1100 1080
rect 1136 1079 1138 1082
rect 1190 1080 1191 1084
rect 1195 1080 1196 1084
rect 1190 1079 1196 1080
rect 1270 1084 1276 1085
rect 1270 1080 1271 1084
rect 1275 1080 1276 1084
rect 1270 1079 1276 1080
rect 1096 1055 1098 1079
rect 1135 1078 1139 1079
rect 1135 1073 1139 1074
rect 1159 1078 1163 1079
rect 1159 1073 1163 1074
rect 1191 1078 1195 1079
rect 1191 1073 1195 1074
rect 1199 1078 1203 1079
rect 1199 1073 1203 1074
rect 1247 1078 1251 1079
rect 1247 1073 1251 1074
rect 1271 1078 1275 1079
rect 1271 1073 1275 1074
rect 1303 1078 1307 1079
rect 1303 1073 1307 1074
rect 1136 1070 1138 1073
rect 1158 1072 1164 1073
rect 1134 1069 1140 1070
rect 1134 1065 1135 1069
rect 1139 1065 1140 1069
rect 1158 1068 1159 1072
rect 1163 1068 1164 1072
rect 1158 1067 1164 1068
rect 1198 1072 1204 1073
rect 1198 1068 1199 1072
rect 1203 1068 1204 1072
rect 1198 1067 1204 1068
rect 1246 1072 1252 1073
rect 1246 1068 1247 1072
rect 1251 1068 1252 1072
rect 1246 1067 1252 1068
rect 1302 1072 1308 1073
rect 1302 1068 1303 1072
rect 1307 1068 1308 1072
rect 1302 1067 1308 1068
rect 1134 1064 1140 1065
rect 1328 1056 1330 1114
rect 1344 1113 1346 1125
rect 1372 1120 1374 1158
rect 1422 1152 1428 1153
rect 1422 1148 1423 1152
rect 1427 1148 1428 1152
rect 1422 1147 1428 1148
rect 1486 1152 1492 1153
rect 1486 1148 1487 1152
rect 1491 1148 1492 1152
rect 1486 1147 1492 1148
rect 1424 1131 1426 1147
rect 1488 1131 1490 1147
rect 1516 1144 1518 1202
rect 1558 1192 1564 1193
rect 1558 1188 1559 1192
rect 1563 1188 1564 1192
rect 1558 1187 1564 1188
rect 1622 1192 1628 1193
rect 1622 1188 1623 1192
rect 1627 1188 1628 1192
rect 1622 1187 1628 1188
rect 1559 1186 1563 1187
rect 1559 1181 1563 1182
rect 1623 1186 1627 1187
rect 1623 1181 1627 1182
rect 1631 1186 1635 1187
rect 1631 1181 1635 1182
rect 1558 1180 1564 1181
rect 1558 1176 1559 1180
rect 1563 1176 1564 1180
rect 1558 1175 1564 1176
rect 1630 1180 1636 1181
rect 1630 1176 1631 1180
rect 1635 1176 1636 1180
rect 1630 1175 1636 1176
rect 1582 1163 1588 1164
rect 1582 1159 1583 1163
rect 1587 1159 1588 1163
rect 1582 1158 1588 1159
rect 1558 1152 1564 1153
rect 1558 1148 1559 1152
rect 1563 1148 1564 1152
rect 1558 1147 1564 1148
rect 1514 1143 1520 1144
rect 1514 1139 1515 1143
rect 1519 1139 1520 1143
rect 1514 1138 1520 1139
rect 1560 1131 1562 1147
rect 1415 1130 1419 1131
rect 1415 1125 1419 1126
rect 1423 1130 1427 1131
rect 1423 1125 1427 1126
rect 1487 1130 1491 1131
rect 1487 1125 1491 1126
rect 1559 1130 1563 1131
rect 1559 1125 1563 1126
rect 1567 1130 1571 1131
rect 1584 1128 1586 1158
rect 1672 1153 1674 1202
rect 1678 1192 1684 1193
rect 1678 1188 1679 1192
rect 1683 1188 1684 1192
rect 1678 1187 1684 1188
rect 1734 1192 1740 1193
rect 1734 1188 1735 1192
rect 1739 1188 1740 1192
rect 1734 1187 1740 1188
rect 1790 1192 1796 1193
rect 1790 1188 1791 1192
rect 1795 1188 1796 1192
rect 1790 1187 1796 1188
rect 1846 1192 1852 1193
rect 1846 1188 1847 1192
rect 1851 1188 1852 1192
rect 1846 1187 1852 1188
rect 1902 1192 1908 1193
rect 1902 1188 1903 1192
rect 1907 1188 1908 1192
rect 1902 1187 1908 1188
rect 1966 1192 1972 1193
rect 1966 1188 1967 1192
rect 1971 1188 1972 1192
rect 1966 1187 1972 1188
rect 1679 1186 1683 1187
rect 1679 1181 1683 1182
rect 1711 1186 1715 1187
rect 1711 1181 1715 1182
rect 1735 1186 1739 1187
rect 1735 1181 1739 1182
rect 1791 1186 1795 1187
rect 1791 1181 1795 1182
rect 1799 1186 1803 1187
rect 1799 1181 1803 1182
rect 1847 1186 1851 1187
rect 1847 1181 1851 1182
rect 1887 1186 1891 1187
rect 1887 1181 1891 1182
rect 1903 1186 1907 1187
rect 1903 1181 1907 1182
rect 1967 1186 1971 1187
rect 1967 1181 1971 1182
rect 1983 1186 1987 1187
rect 1983 1181 1987 1182
rect 1710 1180 1716 1181
rect 1710 1176 1711 1180
rect 1715 1176 1716 1180
rect 1710 1175 1716 1176
rect 1798 1180 1804 1181
rect 1798 1176 1799 1180
rect 1803 1176 1804 1180
rect 1798 1175 1804 1176
rect 1886 1180 1892 1181
rect 1886 1176 1887 1180
rect 1891 1176 1892 1180
rect 1886 1175 1892 1176
rect 1982 1180 1988 1181
rect 1982 1176 1983 1180
rect 1987 1176 1988 1180
rect 1982 1175 1988 1176
rect 2008 1164 2010 1222
rect 2032 1221 2034 1233
rect 2072 1221 2074 1233
rect 2086 1227 2092 1228
rect 2086 1223 2087 1227
rect 2091 1223 2092 1227
rect 2086 1222 2092 1223
rect 2030 1220 2036 1221
rect 2030 1216 2031 1220
rect 2035 1216 2036 1220
rect 2030 1215 2036 1216
rect 2070 1220 2076 1221
rect 2070 1216 2071 1220
rect 2075 1216 2076 1220
rect 2070 1215 2076 1216
rect 2088 1208 2090 1222
rect 2120 1213 2122 1233
rect 2118 1212 2124 1213
rect 2118 1208 2119 1212
rect 2123 1208 2124 1212
rect 2078 1207 2084 1208
rect 2078 1203 2079 1207
rect 2083 1203 2084 1207
rect 2078 1202 2084 1203
rect 2086 1207 2092 1208
rect 2118 1207 2124 1208
rect 2086 1203 2087 1207
rect 2091 1203 2092 1207
rect 2086 1202 2092 1203
rect 2030 1192 2036 1193
rect 2030 1188 2031 1192
rect 2035 1188 2036 1192
rect 2030 1187 2036 1188
rect 2070 1192 2076 1193
rect 2070 1188 2071 1192
rect 2075 1188 2076 1192
rect 2070 1187 2076 1188
rect 2031 1186 2035 1187
rect 2031 1181 2035 1182
rect 2071 1186 2075 1187
rect 2071 1181 2075 1182
rect 2070 1180 2076 1181
rect 2070 1176 2071 1180
rect 2075 1176 2076 1180
rect 2070 1175 2076 1176
rect 2006 1163 2012 1164
rect 2006 1159 2007 1163
rect 2011 1159 2012 1163
rect 2006 1158 2012 1159
rect 1630 1152 1636 1153
rect 1630 1148 1631 1152
rect 1635 1148 1636 1152
rect 1672 1151 1690 1153
rect 1630 1147 1636 1148
rect 1632 1131 1634 1147
rect 1688 1136 1690 1151
rect 1710 1152 1716 1153
rect 1710 1148 1711 1152
rect 1715 1148 1716 1152
rect 1710 1147 1716 1148
rect 1798 1152 1804 1153
rect 1798 1148 1799 1152
rect 1803 1148 1804 1152
rect 1798 1147 1804 1148
rect 1886 1152 1892 1153
rect 1886 1148 1887 1152
rect 1891 1148 1892 1152
rect 1886 1147 1892 1148
rect 1982 1152 1988 1153
rect 1982 1148 1983 1152
rect 1987 1148 1988 1152
rect 1982 1147 1988 1148
rect 2070 1152 2076 1153
rect 2070 1148 2071 1152
rect 2075 1148 2076 1152
rect 2070 1147 2076 1148
rect 1686 1135 1692 1136
rect 1686 1131 1687 1135
rect 1691 1131 1692 1135
rect 1712 1131 1714 1147
rect 1800 1131 1802 1147
rect 1888 1131 1890 1147
rect 1984 1131 1986 1147
rect 2002 1143 2008 1144
rect 2002 1139 2003 1143
rect 2007 1139 2008 1143
rect 2002 1138 2008 1139
rect 1631 1130 1635 1131
rect 1567 1125 1571 1126
rect 1582 1127 1588 1128
rect 1370 1119 1376 1120
rect 1370 1115 1371 1119
rect 1375 1115 1376 1119
rect 1370 1114 1376 1115
rect 1416 1113 1418 1125
rect 1478 1119 1484 1120
rect 1478 1115 1479 1119
rect 1483 1115 1484 1119
rect 1478 1114 1484 1115
rect 1342 1112 1348 1113
rect 1342 1108 1343 1112
rect 1347 1108 1348 1112
rect 1342 1107 1348 1108
rect 1414 1112 1420 1113
rect 1414 1108 1415 1112
rect 1419 1108 1420 1112
rect 1414 1107 1420 1108
rect 1370 1099 1376 1100
rect 1370 1095 1371 1099
rect 1375 1095 1376 1099
rect 1370 1094 1376 1095
rect 1470 1099 1476 1100
rect 1470 1095 1471 1099
rect 1475 1095 1476 1099
rect 1470 1094 1476 1095
rect 1342 1084 1348 1085
rect 1342 1080 1343 1084
rect 1347 1080 1348 1084
rect 1342 1079 1348 1080
rect 1343 1078 1347 1079
rect 1343 1073 1347 1074
rect 1351 1078 1355 1079
rect 1351 1073 1355 1074
rect 1350 1072 1356 1073
rect 1350 1068 1351 1072
rect 1355 1068 1356 1072
rect 1350 1067 1356 1068
rect 1214 1055 1220 1056
rect 1095 1054 1099 1055
rect 1095 1049 1099 1050
rect 1134 1052 1140 1053
rect 1086 1035 1092 1036
rect 1086 1031 1087 1035
rect 1091 1031 1092 1035
rect 1086 1030 1092 1031
rect 1096 1029 1098 1049
rect 1134 1048 1135 1052
rect 1139 1048 1140 1052
rect 1214 1051 1215 1055
rect 1219 1051 1220 1055
rect 1214 1050 1220 1051
rect 1222 1055 1228 1056
rect 1222 1051 1223 1055
rect 1227 1051 1228 1055
rect 1222 1050 1228 1051
rect 1318 1055 1324 1056
rect 1318 1051 1319 1055
rect 1323 1051 1324 1055
rect 1318 1050 1324 1051
rect 1326 1055 1332 1056
rect 1326 1051 1327 1055
rect 1331 1051 1332 1055
rect 1326 1050 1332 1051
rect 1134 1047 1140 1048
rect 1094 1028 1100 1029
rect 1094 1024 1095 1028
rect 1099 1024 1100 1028
rect 734 1023 740 1024
rect 734 1019 735 1023
rect 739 1019 740 1023
rect 734 1018 740 1019
rect 882 1023 888 1024
rect 1094 1023 1100 1024
rect 1136 1023 1138 1047
rect 1158 1044 1164 1045
rect 1158 1040 1159 1044
rect 1163 1040 1164 1044
rect 1158 1039 1164 1040
rect 1198 1044 1204 1045
rect 1198 1040 1199 1044
rect 1203 1040 1204 1044
rect 1198 1039 1204 1040
rect 1160 1023 1162 1039
rect 1200 1023 1202 1039
rect 1216 1036 1218 1050
rect 1214 1035 1220 1036
rect 1214 1031 1215 1035
rect 1219 1031 1220 1035
rect 1214 1030 1220 1031
rect 882 1019 883 1023
rect 887 1019 888 1023
rect 882 1018 888 1019
rect 1135 1022 1139 1023
rect 1135 1017 1139 1018
rect 1159 1022 1163 1023
rect 1159 1017 1163 1018
rect 1199 1022 1203 1023
rect 1199 1017 1203 1018
rect 1094 1011 1100 1012
rect 630 1008 636 1009
rect 630 1004 631 1008
rect 635 1004 636 1008
rect 630 1003 636 1004
rect 686 1008 692 1009
rect 686 1004 687 1008
rect 691 1004 692 1008
rect 686 1003 692 1004
rect 742 1008 748 1009
rect 742 1004 743 1008
rect 747 1004 748 1008
rect 742 1003 748 1004
rect 798 1008 804 1009
rect 798 1004 799 1008
rect 803 1004 804 1008
rect 798 1003 804 1004
rect 862 1008 868 1009
rect 862 1004 863 1008
rect 867 1004 868 1008
rect 1094 1007 1095 1011
rect 1099 1007 1100 1011
rect 1094 1006 1100 1007
rect 862 1003 868 1004
rect 632 999 634 1003
rect 688 999 690 1003
rect 744 999 746 1003
rect 800 999 802 1003
rect 864 999 866 1003
rect 1096 999 1098 1006
rect 631 998 635 999
rect 631 993 635 994
rect 687 998 691 999
rect 687 993 691 994
rect 743 998 747 999
rect 743 993 747 994
rect 799 998 803 999
rect 799 993 803 994
rect 863 998 867 999
rect 863 993 867 994
rect 1095 998 1099 999
rect 1136 997 1138 1017
rect 1160 1005 1162 1017
rect 1200 1005 1202 1017
rect 1224 1012 1226 1050
rect 1246 1044 1252 1045
rect 1246 1040 1247 1044
rect 1251 1040 1252 1044
rect 1246 1039 1252 1040
rect 1302 1044 1308 1045
rect 1302 1040 1303 1044
rect 1307 1040 1308 1044
rect 1302 1039 1308 1040
rect 1248 1023 1250 1039
rect 1266 1035 1272 1036
rect 1266 1031 1267 1035
rect 1271 1031 1272 1035
rect 1266 1030 1272 1031
rect 1239 1022 1243 1023
rect 1239 1017 1243 1018
rect 1247 1022 1251 1023
rect 1247 1017 1251 1018
rect 1214 1011 1220 1012
rect 1214 1007 1215 1011
rect 1219 1007 1220 1011
rect 1214 1006 1220 1007
rect 1222 1011 1228 1012
rect 1222 1007 1223 1011
rect 1227 1007 1228 1011
rect 1222 1006 1228 1007
rect 1158 1004 1164 1005
rect 1158 1000 1159 1004
rect 1163 1000 1164 1004
rect 1158 999 1164 1000
rect 1198 1004 1204 1005
rect 1198 1000 1199 1004
rect 1203 1000 1204 1004
rect 1198 999 1204 1000
rect 1095 993 1099 994
rect 1134 996 1140 997
rect 630 992 636 993
rect 630 988 631 992
rect 635 988 636 992
rect 630 987 636 988
rect 686 992 692 993
rect 686 988 687 992
rect 691 988 692 992
rect 686 987 692 988
rect 742 992 748 993
rect 742 988 743 992
rect 747 988 748 992
rect 742 987 748 988
rect 798 992 804 993
rect 798 988 799 992
rect 803 988 804 992
rect 1096 990 1098 993
rect 1134 992 1135 996
rect 1139 992 1140 996
rect 1216 992 1218 1006
rect 1240 1005 1242 1017
rect 1238 1004 1244 1005
rect 1238 1000 1239 1004
rect 1243 1000 1244 1004
rect 1238 999 1244 1000
rect 1268 992 1270 1030
rect 1304 1023 1306 1039
rect 1320 1036 1322 1050
rect 1350 1044 1356 1045
rect 1350 1040 1351 1044
rect 1355 1040 1356 1044
rect 1350 1039 1356 1040
rect 1318 1035 1324 1036
rect 1318 1031 1319 1035
rect 1323 1031 1324 1035
rect 1318 1030 1324 1031
rect 1352 1023 1354 1039
rect 1372 1036 1374 1094
rect 1414 1084 1420 1085
rect 1414 1080 1415 1084
rect 1419 1080 1420 1084
rect 1414 1079 1420 1080
rect 1399 1078 1403 1079
rect 1399 1073 1403 1074
rect 1415 1078 1419 1079
rect 1415 1073 1419 1074
rect 1455 1078 1459 1079
rect 1455 1073 1459 1074
rect 1398 1072 1404 1073
rect 1398 1068 1399 1072
rect 1403 1068 1404 1072
rect 1398 1067 1404 1068
rect 1454 1072 1460 1073
rect 1454 1068 1455 1072
rect 1459 1068 1460 1072
rect 1454 1067 1460 1068
rect 1414 1055 1420 1056
rect 1414 1051 1415 1055
rect 1419 1051 1420 1055
rect 1414 1050 1420 1051
rect 1426 1055 1432 1056
rect 1426 1051 1427 1055
rect 1431 1051 1432 1055
rect 1426 1050 1432 1051
rect 1398 1044 1404 1045
rect 1398 1040 1399 1044
rect 1403 1040 1404 1044
rect 1398 1039 1404 1040
rect 1370 1035 1376 1036
rect 1370 1031 1371 1035
rect 1375 1031 1376 1035
rect 1370 1030 1376 1031
rect 1400 1023 1402 1039
rect 1416 1036 1418 1050
rect 1414 1035 1420 1036
rect 1414 1031 1415 1035
rect 1419 1031 1420 1035
rect 1414 1030 1420 1031
rect 1295 1022 1299 1023
rect 1295 1017 1299 1018
rect 1303 1022 1307 1023
rect 1303 1017 1307 1018
rect 1351 1022 1355 1023
rect 1351 1017 1355 1018
rect 1399 1022 1403 1023
rect 1399 1017 1403 1018
rect 1407 1022 1411 1023
rect 1407 1017 1411 1018
rect 1296 1005 1298 1017
rect 1310 1011 1316 1012
rect 1310 1007 1311 1011
rect 1315 1007 1316 1011
rect 1310 1006 1316 1007
rect 1294 1004 1300 1005
rect 1294 1000 1295 1004
rect 1299 1000 1300 1004
rect 1294 999 1300 1000
rect 1312 992 1314 1006
rect 1352 1005 1354 1017
rect 1358 1011 1364 1012
rect 1358 1007 1359 1011
rect 1363 1007 1364 1011
rect 1358 1006 1364 1007
rect 1398 1011 1404 1012
rect 1398 1007 1399 1011
rect 1403 1007 1404 1011
rect 1398 1006 1404 1007
rect 1350 1004 1356 1005
rect 1350 1000 1351 1004
rect 1355 1000 1356 1004
rect 1350 999 1356 1000
rect 1360 992 1362 1006
rect 1134 991 1140 992
rect 1206 991 1212 992
rect 798 987 804 988
rect 1094 989 1100 990
rect 608 985 614 987
rect 1094 985 1095 989
rect 1099 985 1100 989
rect 1206 987 1207 991
rect 1211 987 1212 991
rect 1206 986 1212 987
rect 1214 991 1220 992
rect 1214 987 1215 991
rect 1219 987 1220 991
rect 1214 986 1220 987
rect 1266 991 1272 992
rect 1266 987 1267 991
rect 1271 987 1272 991
rect 1266 986 1272 987
rect 1310 991 1316 992
rect 1310 987 1311 991
rect 1315 987 1316 991
rect 1310 986 1316 987
rect 1358 991 1364 992
rect 1358 987 1359 991
rect 1363 987 1364 991
rect 1358 986 1364 987
rect 608 976 610 985
rect 1094 984 1100 985
rect 1134 979 1140 980
rect 358 975 364 976
rect 358 971 359 975
rect 363 971 364 975
rect 358 970 364 971
rect 418 975 424 976
rect 418 971 419 975
rect 423 971 424 975
rect 418 970 424 971
rect 426 975 432 976
rect 426 971 427 975
rect 431 971 432 975
rect 426 970 432 971
rect 538 975 544 976
rect 538 971 539 975
rect 543 971 544 975
rect 538 970 544 971
rect 546 975 552 976
rect 546 971 547 975
rect 551 971 552 975
rect 546 970 552 971
rect 606 975 612 976
rect 606 971 607 975
rect 611 971 612 975
rect 1134 975 1135 979
rect 1139 975 1140 979
rect 1134 974 1140 975
rect 1158 976 1164 977
rect 606 970 612 971
rect 1094 972 1100 973
rect 342 964 348 965
rect 342 960 343 964
rect 347 960 348 964
rect 342 959 348 960
rect 290 955 296 956
rect 290 951 291 955
rect 295 951 296 955
rect 290 950 296 951
rect 302 955 308 956
rect 302 951 303 955
rect 307 951 308 955
rect 302 950 308 951
rect 344 943 346 959
rect 360 956 362 970
rect 406 964 412 965
rect 406 960 407 964
rect 411 960 412 964
rect 406 959 412 960
rect 358 955 364 956
rect 358 951 359 955
rect 363 951 364 955
rect 358 950 364 951
rect 408 943 410 959
rect 420 956 422 970
rect 418 955 424 956
rect 418 951 419 955
rect 423 951 424 955
rect 418 950 424 951
rect 111 942 115 943
rect 111 937 115 938
rect 135 942 139 943
rect 135 937 139 938
rect 175 942 179 943
rect 175 937 179 938
rect 223 942 227 943
rect 223 937 227 938
rect 263 942 267 943
rect 263 937 267 938
rect 279 942 283 943
rect 279 937 283 938
rect 303 942 307 943
rect 303 937 307 938
rect 343 942 347 943
rect 343 937 347 938
rect 351 942 355 943
rect 351 937 355 938
rect 399 942 403 943
rect 399 937 403 938
rect 407 942 411 943
rect 407 937 411 938
rect 112 917 114 937
rect 264 925 266 937
rect 304 925 306 937
rect 318 931 324 932
rect 318 927 319 931
rect 323 927 324 931
rect 318 926 324 927
rect 262 924 268 925
rect 262 920 263 924
rect 267 920 268 924
rect 262 919 268 920
rect 302 924 308 925
rect 302 920 303 924
rect 307 920 308 924
rect 302 919 308 920
rect 110 916 116 917
rect 110 912 111 916
rect 115 912 116 916
rect 320 912 322 926
rect 352 925 354 937
rect 366 931 372 932
rect 366 927 367 931
rect 371 927 372 931
rect 366 926 372 927
rect 350 924 356 925
rect 350 920 351 924
rect 355 920 356 924
rect 350 919 356 920
rect 368 912 370 926
rect 400 925 402 937
rect 428 932 430 970
rect 470 964 476 965
rect 470 960 471 964
rect 475 960 476 964
rect 470 959 476 960
rect 526 964 532 965
rect 526 960 527 964
rect 531 960 532 964
rect 526 959 532 960
rect 472 943 474 959
rect 482 955 488 956
rect 482 951 483 955
rect 487 951 488 955
rect 482 950 488 951
rect 455 942 459 943
rect 455 937 459 938
rect 471 942 475 943
rect 471 937 475 938
rect 414 931 420 932
rect 414 927 415 931
rect 419 927 420 931
rect 414 926 420 927
rect 426 931 432 932
rect 426 927 427 931
rect 431 927 432 931
rect 426 926 432 927
rect 398 924 404 925
rect 398 920 399 924
rect 403 920 404 924
rect 398 919 404 920
rect 416 912 418 926
rect 456 925 458 937
rect 454 924 460 925
rect 454 920 455 924
rect 459 920 460 924
rect 454 919 460 920
rect 484 912 486 950
rect 528 943 530 959
rect 540 956 542 970
rect 1094 968 1095 972
rect 1099 968 1100 972
rect 1094 967 1100 968
rect 582 964 588 965
rect 582 960 583 964
rect 587 960 588 964
rect 582 959 588 960
rect 630 964 636 965
rect 630 960 631 964
rect 635 960 636 964
rect 630 959 636 960
rect 686 964 692 965
rect 686 960 687 964
rect 691 960 692 964
rect 686 959 692 960
rect 742 964 748 965
rect 742 960 743 964
rect 747 960 748 964
rect 742 959 748 960
rect 798 964 804 965
rect 798 960 799 964
rect 803 960 804 964
rect 798 959 804 960
rect 538 955 544 956
rect 538 951 539 955
rect 543 951 544 955
rect 538 950 544 951
rect 584 943 586 959
rect 632 943 634 959
rect 688 943 690 959
rect 714 947 720 948
rect 714 943 715 947
rect 719 943 720 947
rect 744 943 746 959
rect 800 943 802 959
rect 1096 943 1098 967
rect 1136 963 1138 974
rect 1158 972 1159 976
rect 1163 972 1164 976
rect 1158 971 1164 972
rect 1198 976 1204 977
rect 1198 972 1199 976
rect 1203 972 1204 976
rect 1198 971 1204 972
rect 1208 971 1210 986
rect 1238 976 1244 977
rect 1238 972 1239 976
rect 1243 972 1244 976
rect 1238 971 1244 972
rect 1294 976 1300 977
rect 1294 972 1295 976
rect 1299 972 1300 976
rect 1294 971 1300 972
rect 1350 976 1356 977
rect 1350 972 1351 976
rect 1355 972 1356 976
rect 1350 971 1356 972
rect 1160 963 1162 971
rect 1200 963 1202 971
rect 1208 969 1226 971
rect 1135 962 1139 963
rect 1135 957 1139 958
rect 1159 962 1163 963
rect 1159 957 1163 958
rect 1199 962 1203 963
rect 1199 957 1203 958
rect 1207 962 1211 963
rect 1207 957 1211 958
rect 1136 954 1138 957
rect 1158 956 1164 957
rect 1134 953 1140 954
rect 1134 949 1135 953
rect 1139 949 1140 953
rect 1158 952 1159 956
rect 1163 952 1164 956
rect 1158 951 1164 952
rect 1206 956 1212 957
rect 1206 952 1207 956
rect 1211 952 1212 956
rect 1206 951 1212 952
rect 1134 948 1140 949
rect 511 942 515 943
rect 511 937 515 938
rect 527 942 531 943
rect 527 937 531 938
rect 567 942 571 943
rect 567 937 571 938
rect 583 942 587 943
rect 583 937 587 938
rect 623 942 627 943
rect 623 937 627 938
rect 631 942 635 943
rect 631 937 635 938
rect 687 942 691 943
rect 714 942 720 943
rect 743 942 747 943
rect 687 937 691 938
rect 512 925 514 937
rect 522 931 528 932
rect 522 927 523 931
rect 527 927 528 931
rect 522 926 528 927
rect 510 924 516 925
rect 510 920 511 924
rect 515 920 516 924
rect 510 919 516 920
rect 524 912 526 926
rect 568 925 570 937
rect 574 931 580 932
rect 574 927 575 931
rect 579 927 580 931
rect 574 926 580 927
rect 566 924 572 925
rect 566 920 567 924
rect 571 920 572 924
rect 566 919 572 920
rect 576 912 578 926
rect 624 925 626 937
rect 638 931 644 932
rect 638 927 639 931
rect 643 927 644 931
rect 638 926 644 927
rect 646 931 652 932
rect 646 927 647 931
rect 651 927 652 931
rect 646 926 652 927
rect 622 924 628 925
rect 622 920 623 924
rect 627 920 628 924
rect 622 919 628 920
rect 640 912 642 926
rect 110 911 116 912
rect 290 911 296 912
rect 290 907 291 911
rect 295 907 296 911
rect 290 906 296 907
rect 318 911 324 912
rect 318 907 319 911
rect 323 907 324 911
rect 318 906 324 907
rect 366 911 372 912
rect 366 907 367 911
rect 371 907 372 911
rect 366 906 372 907
rect 414 911 420 912
rect 414 907 415 911
rect 419 907 420 911
rect 414 906 420 907
rect 482 911 488 912
rect 482 907 483 911
rect 487 907 488 911
rect 482 906 488 907
rect 522 911 528 912
rect 522 907 523 911
rect 527 907 528 911
rect 522 906 528 907
rect 574 911 580 912
rect 574 907 575 911
rect 579 907 580 911
rect 574 906 580 907
rect 638 911 644 912
rect 638 907 639 911
rect 643 907 644 911
rect 638 906 644 907
rect 110 899 116 900
rect 110 895 111 899
rect 115 895 116 899
rect 110 894 116 895
rect 262 896 268 897
rect 112 887 114 894
rect 262 892 263 896
rect 267 892 268 896
rect 262 891 268 892
rect 264 887 266 891
rect 111 886 115 887
rect 111 881 115 882
rect 263 886 267 887
rect 263 881 267 882
rect 112 878 114 881
rect 110 877 116 878
rect 110 873 111 877
rect 115 873 116 877
rect 110 872 116 873
rect 110 860 116 861
rect 110 856 111 860
rect 115 856 116 860
rect 110 855 116 856
rect 112 835 114 855
rect 292 836 294 906
rect 302 896 308 897
rect 302 892 303 896
rect 307 892 308 896
rect 302 891 308 892
rect 350 896 356 897
rect 350 892 351 896
rect 355 892 356 896
rect 350 891 356 892
rect 398 896 404 897
rect 398 892 399 896
rect 403 892 404 896
rect 398 891 404 892
rect 454 896 460 897
rect 454 892 455 896
rect 459 892 460 896
rect 454 891 460 892
rect 510 896 516 897
rect 510 892 511 896
rect 515 892 516 896
rect 510 891 516 892
rect 566 896 572 897
rect 566 892 567 896
rect 571 892 572 896
rect 566 891 572 892
rect 622 896 628 897
rect 622 892 623 896
rect 627 892 628 896
rect 622 891 628 892
rect 304 887 306 891
rect 352 887 354 891
rect 400 887 402 891
rect 456 887 458 891
rect 512 887 514 891
rect 568 887 570 891
rect 624 887 626 891
rect 303 886 307 887
rect 303 881 307 882
rect 351 886 355 887
rect 351 881 355 882
rect 399 886 403 887
rect 399 881 403 882
rect 415 886 419 887
rect 415 881 419 882
rect 455 886 459 887
rect 455 881 459 882
rect 479 886 483 887
rect 479 881 483 882
rect 511 886 515 887
rect 511 881 515 882
rect 551 886 555 887
rect 551 881 555 882
rect 567 886 571 887
rect 567 881 571 882
rect 623 886 627 887
rect 623 881 627 882
rect 302 880 308 881
rect 302 876 303 880
rect 307 876 308 880
rect 302 875 308 876
rect 350 880 356 881
rect 350 876 351 880
rect 355 876 356 880
rect 350 875 356 876
rect 414 880 420 881
rect 414 876 415 880
rect 419 876 420 880
rect 414 875 420 876
rect 478 880 484 881
rect 478 876 479 880
rect 483 876 484 880
rect 478 875 484 876
rect 550 880 556 881
rect 550 876 551 880
rect 555 876 556 880
rect 550 875 556 876
rect 622 880 628 881
rect 622 876 623 880
rect 627 876 628 880
rect 622 875 628 876
rect 648 864 650 926
rect 688 925 690 937
rect 686 924 692 925
rect 686 920 687 924
rect 691 920 692 924
rect 686 919 692 920
rect 716 912 718 942
rect 743 937 747 938
rect 751 942 755 943
rect 751 937 755 938
rect 799 942 803 943
rect 799 937 803 938
rect 815 942 819 943
rect 815 937 819 938
rect 879 942 883 943
rect 879 937 883 938
rect 943 942 947 943
rect 943 937 947 938
rect 1007 942 1011 943
rect 1007 937 1011 938
rect 1047 942 1051 943
rect 1047 937 1051 938
rect 1095 942 1099 943
rect 1095 937 1099 938
rect 1214 939 1220 940
rect 752 925 754 937
rect 766 931 772 932
rect 766 927 767 931
rect 771 927 772 931
rect 766 926 772 927
rect 750 924 756 925
rect 750 920 751 924
rect 755 920 756 924
rect 750 919 756 920
rect 768 912 770 926
rect 816 925 818 937
rect 830 931 836 932
rect 830 927 831 931
rect 835 927 836 931
rect 830 926 836 927
rect 814 924 820 925
rect 814 920 815 924
rect 819 920 820 924
rect 814 919 820 920
rect 832 912 834 926
rect 880 925 882 937
rect 894 931 900 932
rect 894 927 895 931
rect 899 927 900 931
rect 894 926 900 927
rect 878 924 884 925
rect 878 920 879 924
rect 883 920 884 924
rect 878 919 884 920
rect 896 912 898 926
rect 944 925 946 937
rect 958 931 964 932
rect 958 927 959 931
rect 963 927 964 931
rect 958 926 964 927
rect 966 931 972 932
rect 966 927 967 931
rect 971 927 972 931
rect 966 926 972 927
rect 942 924 948 925
rect 942 920 943 924
rect 947 920 948 924
rect 942 919 948 920
rect 960 912 962 926
rect 714 911 720 912
rect 714 907 715 911
rect 719 907 720 911
rect 714 906 720 907
rect 766 911 772 912
rect 766 907 767 911
rect 771 907 772 911
rect 766 906 772 907
rect 830 911 836 912
rect 830 907 831 911
rect 835 907 836 911
rect 830 906 836 907
rect 894 911 900 912
rect 894 907 895 911
rect 899 907 900 911
rect 894 906 900 907
rect 958 911 964 912
rect 958 907 959 911
rect 963 907 964 911
rect 958 906 964 907
rect 686 896 692 897
rect 686 892 687 896
rect 691 892 692 896
rect 686 891 692 892
rect 750 896 756 897
rect 750 892 751 896
rect 755 892 756 896
rect 750 891 756 892
rect 814 896 820 897
rect 814 892 815 896
rect 819 892 820 896
rect 814 891 820 892
rect 878 896 884 897
rect 878 892 879 896
rect 883 892 884 896
rect 878 891 884 892
rect 942 896 948 897
rect 942 892 943 896
rect 947 892 948 896
rect 942 891 948 892
rect 688 887 690 891
rect 752 887 754 891
rect 816 887 818 891
rect 880 887 882 891
rect 944 887 946 891
rect 687 886 691 887
rect 687 881 691 882
rect 695 886 699 887
rect 695 881 699 882
rect 751 886 755 887
rect 751 881 755 882
rect 767 886 771 887
rect 767 881 771 882
rect 815 886 819 887
rect 815 881 819 882
rect 831 886 835 887
rect 831 881 835 882
rect 879 886 883 887
rect 879 881 883 882
rect 887 886 891 887
rect 887 881 891 882
rect 943 886 947 887
rect 943 881 947 882
rect 694 880 700 881
rect 694 876 695 880
rect 699 876 700 880
rect 694 875 700 876
rect 766 880 772 881
rect 766 876 767 880
rect 771 876 772 880
rect 766 875 772 876
rect 830 880 836 881
rect 830 876 831 880
rect 835 876 836 880
rect 830 875 836 876
rect 886 880 892 881
rect 886 876 887 880
rect 891 876 892 880
rect 886 875 892 876
rect 942 880 948 881
rect 942 876 943 880
rect 947 876 948 880
rect 942 875 948 876
rect 968 872 970 926
rect 1008 925 1010 937
rect 1048 925 1050 937
rect 1062 931 1068 932
rect 1062 927 1063 931
rect 1067 927 1068 931
rect 1062 926 1068 927
rect 1006 924 1012 925
rect 1006 920 1007 924
rect 1011 920 1012 924
rect 1006 919 1012 920
rect 1046 924 1052 925
rect 1046 920 1047 924
rect 1051 920 1052 924
rect 1046 919 1052 920
rect 1064 912 1066 926
rect 1096 917 1098 937
rect 1134 936 1140 937
rect 1134 932 1135 936
rect 1139 932 1140 936
rect 1214 935 1215 939
rect 1219 935 1220 939
rect 1214 934 1220 935
rect 1134 931 1140 932
rect 1094 916 1100 917
rect 1094 912 1095 916
rect 1099 912 1100 916
rect 1054 911 1060 912
rect 1054 907 1055 911
rect 1059 907 1060 911
rect 1054 906 1060 907
rect 1062 911 1068 912
rect 1094 911 1100 912
rect 1136 911 1138 931
rect 1158 928 1164 929
rect 1158 924 1159 928
rect 1163 924 1164 928
rect 1158 923 1164 924
rect 1206 928 1212 929
rect 1206 924 1207 928
rect 1211 924 1212 928
rect 1206 923 1212 924
rect 1160 911 1162 923
rect 1208 911 1210 923
rect 1216 920 1218 934
rect 1224 920 1226 969
rect 1240 963 1242 971
rect 1296 963 1298 971
rect 1352 963 1354 971
rect 1239 962 1243 963
rect 1239 957 1243 958
rect 1287 962 1291 963
rect 1287 957 1291 958
rect 1295 962 1299 963
rect 1295 957 1299 958
rect 1351 962 1355 963
rect 1351 957 1355 958
rect 1375 962 1379 963
rect 1375 957 1379 958
rect 1286 956 1292 957
rect 1286 952 1287 956
rect 1291 952 1292 956
rect 1286 951 1292 952
rect 1374 956 1380 957
rect 1374 952 1375 956
rect 1379 952 1380 956
rect 1374 951 1380 952
rect 1400 940 1402 1006
rect 1408 1005 1410 1017
rect 1428 1012 1430 1050
rect 1454 1044 1460 1045
rect 1472 1044 1474 1094
rect 1480 1056 1482 1114
rect 1488 1113 1490 1125
rect 1568 1113 1570 1125
rect 1582 1123 1583 1127
rect 1587 1123 1588 1127
rect 1631 1125 1635 1126
rect 1655 1130 1659 1131
rect 1686 1130 1692 1131
rect 1711 1130 1715 1131
rect 1655 1125 1659 1126
rect 1711 1125 1715 1126
rect 1751 1130 1755 1131
rect 1751 1125 1755 1126
rect 1799 1130 1803 1131
rect 1799 1125 1803 1126
rect 1855 1130 1859 1131
rect 1855 1125 1859 1126
rect 1887 1130 1891 1131
rect 1887 1125 1891 1126
rect 1959 1130 1963 1131
rect 1959 1125 1963 1126
rect 1983 1130 1987 1131
rect 1983 1125 1987 1126
rect 1582 1122 1588 1123
rect 1582 1119 1588 1120
rect 1582 1115 1583 1119
rect 1587 1115 1588 1119
rect 1582 1114 1588 1115
rect 1486 1112 1492 1113
rect 1486 1108 1487 1112
rect 1491 1108 1492 1112
rect 1486 1107 1492 1108
rect 1566 1112 1572 1113
rect 1566 1108 1567 1112
rect 1571 1108 1572 1112
rect 1566 1107 1572 1108
rect 1584 1100 1586 1114
rect 1656 1113 1658 1125
rect 1670 1119 1676 1120
rect 1670 1115 1671 1119
rect 1675 1115 1676 1119
rect 1670 1114 1676 1115
rect 1654 1112 1660 1113
rect 1654 1108 1655 1112
rect 1659 1108 1660 1112
rect 1654 1107 1660 1108
rect 1672 1100 1674 1114
rect 1752 1113 1754 1125
rect 1766 1119 1772 1120
rect 1766 1115 1767 1119
rect 1771 1115 1772 1119
rect 1766 1114 1772 1115
rect 1750 1112 1756 1113
rect 1750 1108 1751 1112
rect 1755 1108 1756 1112
rect 1750 1107 1756 1108
rect 1768 1100 1770 1114
rect 1856 1113 1858 1125
rect 1870 1119 1876 1120
rect 1870 1115 1871 1119
rect 1875 1115 1876 1119
rect 1870 1114 1876 1115
rect 1854 1112 1860 1113
rect 1854 1108 1855 1112
rect 1859 1108 1860 1112
rect 1854 1107 1860 1108
rect 1872 1100 1874 1114
rect 1960 1113 1962 1125
rect 1982 1119 1988 1120
rect 1982 1115 1983 1119
rect 1987 1115 1988 1119
rect 1982 1114 1988 1115
rect 1958 1112 1964 1113
rect 1958 1108 1959 1112
rect 1963 1108 1964 1112
rect 1958 1107 1964 1108
rect 1494 1099 1500 1100
rect 1494 1095 1495 1099
rect 1499 1095 1500 1099
rect 1494 1094 1500 1095
rect 1582 1099 1588 1100
rect 1582 1095 1583 1099
rect 1587 1095 1588 1099
rect 1582 1094 1588 1095
rect 1670 1099 1676 1100
rect 1670 1095 1671 1099
rect 1675 1095 1676 1099
rect 1670 1094 1676 1095
rect 1766 1099 1772 1100
rect 1766 1095 1767 1099
rect 1771 1095 1772 1099
rect 1766 1094 1772 1095
rect 1870 1099 1876 1100
rect 1870 1095 1871 1099
rect 1875 1095 1876 1099
rect 1870 1094 1876 1095
rect 1486 1084 1492 1085
rect 1486 1080 1487 1084
rect 1491 1080 1492 1084
rect 1486 1079 1492 1080
rect 1487 1078 1491 1079
rect 1487 1073 1491 1074
rect 1478 1055 1484 1056
rect 1478 1051 1479 1055
rect 1483 1051 1484 1055
rect 1478 1050 1484 1051
rect 1454 1040 1455 1044
rect 1459 1040 1460 1044
rect 1454 1039 1460 1040
rect 1470 1043 1476 1044
rect 1470 1039 1471 1043
rect 1475 1039 1476 1043
rect 1456 1023 1458 1039
rect 1470 1038 1476 1039
rect 1496 1036 1498 1094
rect 1566 1084 1572 1085
rect 1566 1080 1567 1084
rect 1571 1080 1572 1084
rect 1566 1079 1572 1080
rect 1654 1084 1660 1085
rect 1654 1080 1655 1084
rect 1659 1080 1660 1084
rect 1654 1079 1660 1080
rect 1750 1084 1756 1085
rect 1750 1080 1751 1084
rect 1755 1080 1756 1084
rect 1750 1079 1756 1080
rect 1854 1084 1860 1085
rect 1854 1080 1855 1084
rect 1859 1080 1860 1084
rect 1854 1079 1860 1080
rect 1958 1084 1964 1085
rect 1958 1080 1959 1084
rect 1963 1080 1964 1084
rect 1958 1079 1964 1080
rect 1511 1078 1515 1079
rect 1511 1073 1515 1074
rect 1567 1078 1571 1079
rect 1567 1073 1571 1074
rect 1583 1078 1587 1079
rect 1583 1073 1587 1074
rect 1655 1078 1659 1079
rect 1655 1073 1659 1074
rect 1663 1078 1667 1079
rect 1663 1073 1667 1074
rect 1751 1078 1755 1079
rect 1751 1073 1755 1074
rect 1759 1078 1763 1079
rect 1759 1073 1763 1074
rect 1855 1078 1859 1079
rect 1855 1073 1859 1074
rect 1863 1078 1867 1079
rect 1863 1073 1867 1074
rect 1959 1078 1963 1079
rect 1959 1073 1963 1074
rect 1967 1078 1971 1079
rect 1967 1073 1971 1074
rect 1510 1072 1516 1073
rect 1510 1068 1511 1072
rect 1515 1068 1516 1072
rect 1510 1067 1516 1068
rect 1582 1072 1588 1073
rect 1582 1068 1583 1072
rect 1587 1068 1588 1072
rect 1582 1067 1588 1068
rect 1662 1072 1668 1073
rect 1662 1068 1663 1072
rect 1667 1068 1668 1072
rect 1662 1067 1668 1068
rect 1758 1072 1764 1073
rect 1758 1068 1759 1072
rect 1763 1068 1764 1072
rect 1758 1067 1764 1068
rect 1862 1072 1868 1073
rect 1862 1068 1863 1072
rect 1867 1068 1868 1072
rect 1862 1067 1868 1068
rect 1966 1072 1972 1073
rect 1966 1068 1967 1072
rect 1971 1068 1972 1072
rect 1966 1067 1972 1068
rect 1886 1063 1892 1064
rect 1886 1059 1887 1063
rect 1891 1059 1892 1063
rect 1886 1058 1892 1059
rect 1598 1055 1604 1056
rect 1598 1051 1599 1055
rect 1603 1051 1604 1055
rect 1598 1050 1604 1051
rect 1678 1055 1684 1056
rect 1678 1051 1679 1055
rect 1683 1051 1684 1055
rect 1678 1050 1684 1051
rect 1510 1044 1516 1045
rect 1510 1040 1511 1044
rect 1515 1040 1516 1044
rect 1510 1039 1516 1040
rect 1582 1044 1588 1045
rect 1582 1040 1583 1044
rect 1587 1040 1588 1044
rect 1582 1039 1588 1040
rect 1494 1035 1500 1036
rect 1494 1031 1495 1035
rect 1499 1031 1500 1035
rect 1494 1030 1500 1031
rect 1512 1023 1514 1039
rect 1584 1023 1586 1039
rect 1600 1036 1602 1050
rect 1662 1044 1668 1045
rect 1662 1040 1663 1044
rect 1667 1040 1668 1044
rect 1662 1039 1668 1040
rect 1598 1035 1604 1036
rect 1598 1031 1599 1035
rect 1603 1031 1604 1035
rect 1598 1030 1604 1031
rect 1664 1023 1666 1039
rect 1455 1022 1459 1023
rect 1455 1017 1459 1018
rect 1463 1022 1467 1023
rect 1463 1017 1467 1018
rect 1511 1022 1515 1023
rect 1511 1017 1515 1018
rect 1519 1022 1523 1023
rect 1519 1017 1523 1018
rect 1575 1022 1579 1023
rect 1575 1017 1579 1018
rect 1583 1022 1587 1023
rect 1583 1017 1587 1018
rect 1639 1022 1643 1023
rect 1639 1017 1643 1018
rect 1663 1022 1667 1023
rect 1663 1017 1667 1018
rect 1426 1011 1432 1012
rect 1426 1007 1427 1011
rect 1431 1007 1432 1011
rect 1426 1006 1432 1007
rect 1464 1005 1466 1017
rect 1520 1005 1522 1017
rect 1576 1005 1578 1017
rect 1590 1011 1596 1012
rect 1590 1007 1591 1011
rect 1595 1007 1596 1011
rect 1590 1006 1596 1007
rect 1406 1004 1412 1005
rect 1406 1000 1407 1004
rect 1411 1000 1412 1004
rect 1406 999 1412 1000
rect 1462 1004 1468 1005
rect 1462 1000 1463 1004
rect 1467 1000 1468 1004
rect 1462 999 1468 1000
rect 1518 1004 1524 1005
rect 1518 1000 1519 1004
rect 1523 1000 1524 1004
rect 1518 999 1524 1000
rect 1574 1004 1580 1005
rect 1574 1000 1575 1004
rect 1579 1000 1580 1004
rect 1574 999 1580 1000
rect 1592 992 1594 1006
rect 1640 1005 1642 1017
rect 1680 1016 1682 1050
rect 1758 1044 1764 1045
rect 1758 1040 1759 1044
rect 1763 1040 1764 1044
rect 1758 1039 1764 1040
rect 1862 1044 1868 1045
rect 1862 1040 1863 1044
rect 1867 1040 1868 1044
rect 1862 1039 1868 1040
rect 1760 1023 1762 1039
rect 1864 1023 1866 1039
rect 1888 1036 1890 1058
rect 1966 1044 1972 1045
rect 1966 1040 1967 1044
rect 1971 1040 1972 1044
rect 1966 1039 1972 1040
rect 1886 1035 1892 1036
rect 1886 1031 1887 1035
rect 1891 1031 1892 1035
rect 1886 1030 1892 1031
rect 1968 1023 1970 1039
rect 1711 1022 1715 1023
rect 1711 1017 1715 1018
rect 1759 1022 1763 1023
rect 1759 1017 1763 1018
rect 1791 1022 1795 1023
rect 1791 1017 1795 1018
rect 1863 1022 1867 1023
rect 1863 1017 1867 1018
rect 1879 1022 1883 1023
rect 1879 1017 1883 1018
rect 1967 1022 1971 1023
rect 1967 1017 1971 1018
rect 1678 1015 1684 1016
rect 1654 1011 1660 1012
rect 1654 1007 1655 1011
rect 1659 1007 1660 1011
rect 1678 1011 1679 1015
rect 1683 1011 1684 1015
rect 1678 1010 1684 1011
rect 1654 1006 1660 1007
rect 1638 1004 1644 1005
rect 1638 1000 1639 1004
rect 1643 1000 1644 1004
rect 1638 999 1644 1000
rect 1656 992 1658 1006
rect 1712 1005 1714 1017
rect 1792 1005 1794 1017
rect 1880 1005 1882 1017
rect 1894 1011 1900 1012
rect 1894 1007 1895 1011
rect 1899 1007 1900 1011
rect 1894 1006 1900 1007
rect 1710 1004 1716 1005
rect 1710 1000 1711 1004
rect 1715 1000 1716 1004
rect 1710 999 1716 1000
rect 1790 1004 1796 1005
rect 1790 1000 1791 1004
rect 1795 1000 1796 1004
rect 1790 999 1796 1000
rect 1878 1004 1884 1005
rect 1878 1000 1879 1004
rect 1883 1000 1884 1004
rect 1878 999 1884 1000
rect 1896 992 1898 1006
rect 1968 1005 1970 1017
rect 1966 1004 1972 1005
rect 1966 1000 1967 1004
rect 1971 1000 1972 1004
rect 1966 999 1972 1000
rect 1984 992 1986 1114
rect 2004 1104 2006 1138
rect 2072 1131 2074 1147
rect 2080 1144 2082 1202
rect 2118 1195 2124 1196
rect 2118 1191 2119 1195
rect 2123 1191 2124 1195
rect 2118 1190 2124 1191
rect 2120 1187 2122 1190
rect 2119 1186 2123 1187
rect 2119 1181 2123 1182
rect 2120 1178 2122 1181
rect 2118 1177 2124 1178
rect 2118 1173 2119 1177
rect 2123 1173 2124 1177
rect 2118 1172 2124 1173
rect 2094 1163 2100 1164
rect 2094 1159 2095 1163
rect 2099 1159 2100 1163
rect 2094 1158 2100 1159
rect 2118 1160 2124 1161
rect 2078 1143 2084 1144
rect 2078 1139 2079 1143
rect 2083 1139 2084 1143
rect 2078 1138 2084 1139
rect 2071 1130 2075 1131
rect 2071 1125 2075 1126
rect 2072 1113 2074 1125
rect 2096 1120 2098 1158
rect 2118 1156 2119 1160
rect 2123 1156 2124 1160
rect 2118 1155 2124 1156
rect 2120 1131 2122 1155
rect 2119 1130 2123 1131
rect 2119 1125 2123 1126
rect 2094 1119 2100 1120
rect 2094 1115 2095 1119
rect 2099 1115 2100 1119
rect 2094 1114 2100 1115
rect 2070 1112 2076 1113
rect 2070 1108 2071 1112
rect 2075 1108 2076 1112
rect 2070 1107 2076 1108
rect 2120 1105 2122 1125
rect 2118 1104 2124 1105
rect 2002 1103 2008 1104
rect 2002 1099 2003 1103
rect 2007 1099 2008 1103
rect 2118 1100 2119 1104
rect 2123 1100 2124 1104
rect 2002 1098 2008 1099
rect 2094 1099 2100 1100
rect 2118 1099 2124 1100
rect 2094 1095 2095 1099
rect 2099 1095 2100 1099
rect 2094 1094 2100 1095
rect 2070 1084 2076 1085
rect 2070 1080 2071 1084
rect 2075 1080 2076 1084
rect 2070 1079 2076 1080
rect 2071 1078 2075 1079
rect 2071 1073 2075 1074
rect 2070 1072 2076 1073
rect 2070 1068 2071 1072
rect 2075 1068 2076 1072
rect 2070 1067 2076 1068
rect 1990 1055 1996 1056
rect 1990 1051 1991 1055
rect 1995 1051 1996 1055
rect 1990 1050 1996 1051
rect 2046 1055 2052 1056
rect 2046 1051 2047 1055
rect 2051 1051 2052 1055
rect 2046 1050 2052 1051
rect 1992 1020 1994 1050
rect 2048 1036 2050 1050
rect 2070 1044 2076 1045
rect 2070 1040 2071 1044
rect 2075 1040 2076 1044
rect 2070 1039 2076 1040
rect 2046 1035 2052 1036
rect 2046 1031 2047 1035
rect 2051 1031 2052 1035
rect 2046 1030 2052 1031
rect 2072 1023 2074 1039
rect 2096 1036 2098 1094
rect 2118 1087 2124 1088
rect 2118 1083 2119 1087
rect 2123 1083 2124 1087
rect 2118 1082 2124 1083
rect 2120 1079 2122 1082
rect 2119 1078 2123 1079
rect 2119 1073 2123 1074
rect 2120 1070 2122 1073
rect 2118 1069 2124 1070
rect 2118 1065 2119 1069
rect 2123 1065 2124 1069
rect 2118 1064 2124 1065
rect 2118 1052 2124 1053
rect 2118 1048 2119 1052
rect 2123 1048 2124 1052
rect 2118 1047 2124 1048
rect 2094 1035 2100 1036
rect 2094 1031 2095 1035
rect 2099 1031 2100 1035
rect 2094 1030 2100 1031
rect 2120 1023 2122 1047
rect 2063 1022 2067 1023
rect 1990 1019 1996 1020
rect 1990 1015 1991 1019
rect 1995 1015 1996 1019
rect 2063 1017 2067 1018
rect 2071 1022 2075 1023
rect 2071 1017 2075 1018
rect 2119 1022 2123 1023
rect 2119 1017 2123 1018
rect 1990 1014 1996 1015
rect 2064 1005 2066 1017
rect 2062 1004 2068 1005
rect 2062 1000 2063 1004
rect 2067 1000 2068 1004
rect 2062 999 2068 1000
rect 2120 997 2122 1017
rect 2118 996 2124 997
rect 2118 992 2119 996
rect 2123 992 2124 996
rect 1482 991 1488 992
rect 1482 987 1483 991
rect 1487 987 1488 991
rect 1482 986 1488 987
rect 1590 991 1596 992
rect 1590 987 1591 991
rect 1595 987 1596 991
rect 1590 986 1596 987
rect 1654 991 1660 992
rect 1654 987 1655 991
rect 1659 987 1660 991
rect 1654 986 1660 987
rect 1778 991 1784 992
rect 1778 987 1779 991
rect 1783 987 1784 991
rect 1778 986 1784 987
rect 1894 991 1900 992
rect 1894 987 1895 991
rect 1899 987 1900 991
rect 1894 986 1900 987
rect 1982 991 1988 992
rect 2118 991 2124 992
rect 1982 987 1983 991
rect 1987 987 1988 991
rect 1982 986 1988 987
rect 1406 976 1412 977
rect 1406 972 1407 976
rect 1411 972 1412 976
rect 1406 971 1412 972
rect 1462 976 1468 977
rect 1462 972 1463 976
rect 1467 972 1468 976
rect 1462 971 1468 972
rect 1408 963 1410 971
rect 1464 963 1466 971
rect 1407 962 1411 963
rect 1407 957 1411 958
rect 1455 962 1459 963
rect 1455 957 1459 958
rect 1463 962 1467 963
rect 1463 957 1467 958
rect 1454 956 1460 957
rect 1454 952 1455 956
rect 1459 952 1460 956
rect 1454 951 1460 952
rect 1390 939 1396 940
rect 1390 935 1391 939
rect 1395 935 1396 939
rect 1390 934 1396 935
rect 1398 939 1404 940
rect 1398 935 1399 939
rect 1403 935 1404 939
rect 1398 934 1404 935
rect 1286 928 1292 929
rect 1286 924 1287 928
rect 1291 924 1292 928
rect 1286 923 1292 924
rect 1374 928 1380 929
rect 1374 924 1375 928
rect 1379 924 1380 928
rect 1374 923 1380 924
rect 1214 919 1220 920
rect 1214 915 1215 919
rect 1219 915 1220 919
rect 1214 914 1220 915
rect 1222 919 1228 920
rect 1222 915 1223 919
rect 1227 915 1228 919
rect 1222 914 1228 915
rect 1266 919 1272 920
rect 1266 915 1267 919
rect 1271 915 1272 919
rect 1266 914 1272 915
rect 1062 907 1063 911
rect 1067 907 1068 911
rect 1062 906 1068 907
rect 1135 910 1139 911
rect 1006 896 1012 897
rect 1006 892 1007 896
rect 1011 892 1012 896
rect 1006 891 1012 892
rect 1046 896 1052 897
rect 1046 892 1047 896
rect 1051 892 1052 896
rect 1046 891 1052 892
rect 1008 887 1010 891
rect 1048 887 1050 891
rect 1007 886 1011 887
rect 1007 881 1011 882
rect 1047 886 1051 887
rect 1047 881 1051 882
rect 1006 880 1012 881
rect 1006 876 1007 880
rect 1011 876 1012 880
rect 1006 875 1012 876
rect 1046 880 1052 881
rect 1046 876 1047 880
rect 1051 876 1052 880
rect 1046 875 1052 876
rect 1056 875 1058 906
rect 1135 905 1139 906
rect 1159 910 1163 911
rect 1159 905 1163 906
rect 1207 910 1211 911
rect 1207 905 1211 906
rect 1239 910 1243 911
rect 1239 905 1243 906
rect 1094 899 1100 900
rect 1094 895 1095 899
rect 1099 895 1100 899
rect 1094 894 1100 895
rect 1096 887 1098 894
rect 1095 886 1099 887
rect 1136 885 1138 905
rect 1240 893 1242 905
rect 1238 892 1244 893
rect 1238 888 1239 892
rect 1243 888 1244 892
rect 1238 887 1244 888
rect 1095 881 1099 882
rect 1134 884 1140 885
rect 1096 878 1098 881
rect 1134 880 1135 884
rect 1139 880 1140 884
rect 1268 880 1270 914
rect 1288 911 1290 923
rect 1376 911 1378 923
rect 1392 920 1394 934
rect 1454 928 1460 929
rect 1454 924 1455 928
rect 1459 924 1460 928
rect 1454 923 1460 924
rect 1390 919 1396 920
rect 1390 915 1391 919
rect 1395 915 1396 919
rect 1390 914 1396 915
rect 1456 911 1458 923
rect 1484 920 1486 986
rect 1518 976 1524 977
rect 1518 972 1519 976
rect 1523 972 1524 976
rect 1518 971 1524 972
rect 1574 976 1580 977
rect 1574 972 1575 976
rect 1579 972 1580 976
rect 1574 971 1580 972
rect 1638 976 1644 977
rect 1638 972 1639 976
rect 1643 972 1644 976
rect 1638 971 1644 972
rect 1710 976 1716 977
rect 1710 972 1711 976
rect 1715 972 1716 976
rect 1710 971 1716 972
rect 1520 963 1522 971
rect 1576 963 1578 971
rect 1640 963 1642 971
rect 1712 963 1714 971
rect 1519 962 1523 963
rect 1519 957 1523 958
rect 1535 962 1539 963
rect 1535 957 1539 958
rect 1575 962 1579 963
rect 1575 957 1579 958
rect 1615 962 1619 963
rect 1615 957 1619 958
rect 1639 962 1643 963
rect 1639 957 1643 958
rect 1687 962 1691 963
rect 1687 957 1691 958
rect 1711 962 1715 963
rect 1711 957 1715 958
rect 1751 962 1755 963
rect 1751 957 1755 958
rect 1534 956 1540 957
rect 1534 952 1535 956
rect 1539 952 1540 956
rect 1534 951 1540 952
rect 1614 956 1620 957
rect 1614 952 1615 956
rect 1619 952 1620 956
rect 1614 951 1620 952
rect 1686 956 1692 957
rect 1686 952 1687 956
rect 1691 952 1692 956
rect 1686 951 1692 952
rect 1750 956 1756 957
rect 1750 952 1751 956
rect 1755 952 1756 956
rect 1750 951 1756 952
rect 1550 939 1556 940
rect 1550 935 1551 939
rect 1555 935 1556 939
rect 1550 934 1556 935
rect 1606 939 1612 940
rect 1606 935 1607 939
rect 1611 935 1612 939
rect 1606 934 1612 935
rect 1534 928 1540 929
rect 1534 924 1535 928
rect 1539 924 1540 928
rect 1534 923 1540 924
rect 1482 919 1488 920
rect 1482 915 1483 919
rect 1487 915 1488 919
rect 1482 914 1488 915
rect 1536 911 1538 923
rect 1552 920 1554 934
rect 1550 919 1556 920
rect 1550 915 1551 919
rect 1555 915 1556 919
rect 1550 914 1556 915
rect 1287 910 1291 911
rect 1287 905 1291 906
rect 1319 910 1323 911
rect 1319 905 1323 906
rect 1375 910 1379 911
rect 1375 905 1379 906
rect 1407 910 1411 911
rect 1407 905 1411 906
rect 1455 910 1459 911
rect 1455 905 1459 906
rect 1495 910 1499 911
rect 1495 905 1499 906
rect 1535 910 1539 911
rect 1535 905 1539 906
rect 1583 910 1587 911
rect 1583 905 1587 906
rect 1320 893 1322 905
rect 1334 899 1340 900
rect 1334 895 1335 899
rect 1339 895 1340 899
rect 1334 894 1340 895
rect 1378 899 1384 900
rect 1378 895 1379 899
rect 1383 895 1384 899
rect 1378 894 1384 895
rect 1386 899 1392 900
rect 1386 895 1387 899
rect 1391 895 1392 899
rect 1386 894 1392 895
rect 1318 892 1324 893
rect 1318 888 1319 892
rect 1323 888 1324 892
rect 1318 887 1324 888
rect 1336 880 1338 894
rect 1380 880 1382 894
rect 1134 879 1140 880
rect 1266 879 1272 880
rect 1094 877 1100 878
rect 1056 873 1066 875
rect 966 871 972 872
rect 966 867 967 871
rect 971 867 972 871
rect 966 866 972 867
rect 310 863 316 864
rect 310 859 311 863
rect 315 859 316 863
rect 310 858 316 859
rect 566 863 572 864
rect 566 859 567 863
rect 571 859 572 863
rect 566 858 572 859
rect 638 863 644 864
rect 638 859 639 863
rect 643 859 644 863
rect 638 858 644 859
rect 646 863 652 864
rect 646 859 647 863
rect 651 859 652 863
rect 646 858 652 859
rect 730 863 736 864
rect 730 859 731 863
rect 735 859 736 863
rect 730 858 736 859
rect 934 863 940 864
rect 934 859 935 863
rect 939 859 940 863
rect 934 858 940 859
rect 1054 863 1060 864
rect 1054 859 1055 863
rect 1059 859 1060 863
rect 1054 858 1060 859
rect 302 852 308 853
rect 302 848 303 852
rect 307 848 308 852
rect 302 847 308 848
rect 290 835 296 836
rect 304 835 306 847
rect 111 834 115 835
rect 111 829 115 830
rect 279 834 283 835
rect 290 831 291 835
rect 295 831 296 835
rect 290 830 296 831
rect 303 834 307 835
rect 279 829 283 830
rect 303 829 307 830
rect 112 809 114 829
rect 280 817 282 829
rect 303 823 309 824
rect 303 819 304 823
rect 308 822 309 823
rect 312 822 314 858
rect 350 852 356 853
rect 350 848 351 852
rect 355 848 356 852
rect 350 847 356 848
rect 414 852 420 853
rect 414 848 415 852
rect 419 848 420 852
rect 414 847 420 848
rect 478 852 484 853
rect 478 848 479 852
rect 483 848 484 852
rect 478 847 484 848
rect 550 852 556 853
rect 550 848 551 852
rect 555 848 556 852
rect 550 847 556 848
rect 352 835 354 847
rect 416 835 418 847
rect 480 835 482 847
rect 506 843 512 844
rect 506 839 507 843
rect 511 839 512 843
rect 506 838 512 839
rect 343 834 347 835
rect 343 829 347 830
rect 351 834 355 835
rect 351 829 355 830
rect 415 834 419 835
rect 415 829 419 830
rect 479 834 483 835
rect 479 829 483 830
rect 487 834 491 835
rect 487 829 491 830
rect 308 820 314 822
rect 334 823 340 824
rect 308 819 309 820
rect 303 818 309 819
rect 334 819 335 823
rect 339 819 340 823
rect 334 818 340 819
rect 278 816 284 817
rect 278 812 279 816
rect 283 812 284 816
rect 278 811 284 812
rect 110 808 116 809
rect 110 804 111 808
rect 115 804 116 808
rect 336 804 338 818
rect 344 817 346 829
rect 416 817 418 829
rect 488 817 490 829
rect 342 816 348 817
rect 342 812 343 816
rect 347 812 348 816
rect 342 811 348 812
rect 414 816 420 817
rect 414 812 415 816
rect 419 812 420 816
rect 414 811 420 812
rect 486 816 492 817
rect 486 812 487 816
rect 491 812 492 816
rect 486 811 492 812
rect 508 804 510 838
rect 552 835 554 847
rect 568 844 570 858
rect 622 852 628 853
rect 622 848 623 852
rect 627 848 628 852
rect 622 847 628 848
rect 566 843 572 844
rect 566 839 567 843
rect 571 839 572 843
rect 566 838 572 839
rect 624 835 626 847
rect 640 844 642 858
rect 694 852 700 853
rect 694 848 695 852
rect 699 848 700 852
rect 694 847 700 848
rect 638 843 644 844
rect 638 839 639 843
rect 643 839 644 843
rect 638 838 644 839
rect 696 835 698 847
rect 732 844 734 858
rect 766 852 772 853
rect 766 848 767 852
rect 771 848 772 852
rect 766 847 772 848
rect 830 852 836 853
rect 830 848 831 852
rect 835 848 836 852
rect 830 847 836 848
rect 886 852 892 853
rect 886 848 887 852
rect 891 848 892 852
rect 886 847 892 848
rect 730 843 736 844
rect 730 839 731 843
rect 735 839 736 843
rect 730 838 736 839
rect 754 835 760 836
rect 768 835 770 847
rect 832 835 834 847
rect 888 835 890 847
rect 551 834 555 835
rect 551 829 555 830
rect 567 834 571 835
rect 567 829 571 830
rect 623 834 627 835
rect 623 829 627 830
rect 647 834 651 835
rect 647 829 651 830
rect 695 834 699 835
rect 695 829 699 830
rect 727 834 731 835
rect 754 831 755 835
rect 759 831 760 835
rect 754 830 760 831
rect 767 834 771 835
rect 727 829 731 830
rect 568 817 570 829
rect 582 823 588 824
rect 582 819 583 823
rect 587 819 588 823
rect 582 818 588 819
rect 566 816 572 817
rect 566 812 567 816
rect 571 812 572 816
rect 566 811 572 812
rect 584 804 586 818
rect 648 817 650 829
rect 662 823 668 824
rect 662 819 663 823
rect 667 819 668 823
rect 662 818 668 819
rect 670 823 676 824
rect 670 819 671 823
rect 675 819 676 823
rect 670 818 676 819
rect 646 816 652 817
rect 646 812 647 816
rect 651 812 652 816
rect 646 811 652 812
rect 664 804 666 818
rect 110 803 116 804
rect 334 803 340 804
rect 334 799 335 803
rect 339 799 340 803
rect 334 798 340 799
rect 442 803 448 804
rect 442 799 443 803
rect 447 799 448 803
rect 442 798 448 799
rect 506 803 512 804
rect 506 799 507 803
rect 511 799 512 803
rect 506 798 512 799
rect 582 803 588 804
rect 582 799 583 803
rect 587 799 588 803
rect 582 798 588 799
rect 662 803 668 804
rect 662 799 663 803
rect 667 799 668 803
rect 662 798 668 799
rect 110 791 116 792
rect 110 787 111 791
rect 115 787 116 791
rect 110 786 116 787
rect 278 788 284 789
rect 112 783 114 786
rect 278 784 279 788
rect 283 784 284 788
rect 278 783 284 784
rect 342 788 348 789
rect 342 784 343 788
rect 347 784 348 788
rect 342 783 348 784
rect 414 788 420 789
rect 414 784 415 788
rect 419 784 420 788
rect 414 783 420 784
rect 111 782 115 783
rect 111 777 115 778
rect 215 782 219 783
rect 215 777 219 778
rect 279 782 283 783
rect 279 777 283 778
rect 343 782 347 783
rect 343 777 347 778
rect 351 782 355 783
rect 351 777 355 778
rect 415 782 419 783
rect 415 777 419 778
rect 423 782 427 783
rect 423 777 427 778
rect 112 774 114 777
rect 214 776 220 777
rect 110 773 116 774
rect 110 769 111 773
rect 115 769 116 773
rect 214 772 215 776
rect 219 772 220 776
rect 214 771 220 772
rect 278 776 284 777
rect 278 772 279 776
rect 283 772 284 776
rect 278 771 284 772
rect 350 776 356 777
rect 350 772 351 776
rect 355 772 356 776
rect 350 771 356 772
rect 422 776 428 777
rect 422 772 423 776
rect 427 772 428 776
rect 422 771 428 772
rect 110 768 116 769
rect 202 759 208 760
rect 110 756 116 757
rect 110 752 111 756
rect 115 752 116 756
rect 202 755 203 759
rect 207 755 208 759
rect 202 754 208 755
rect 110 751 116 752
rect 112 731 114 751
rect 111 730 115 731
rect 111 725 115 726
rect 175 730 179 731
rect 175 725 179 726
rect 112 705 114 725
rect 176 713 178 725
rect 204 720 206 754
rect 214 748 220 749
rect 214 744 215 748
rect 219 744 220 748
rect 214 743 220 744
rect 278 748 284 749
rect 278 744 279 748
rect 283 744 284 748
rect 278 743 284 744
rect 350 748 356 749
rect 350 744 351 748
rect 355 744 356 748
rect 350 743 356 744
rect 422 748 428 749
rect 422 744 423 748
rect 427 744 428 748
rect 422 743 428 744
rect 216 731 218 743
rect 280 731 282 743
rect 352 731 354 743
rect 424 731 426 743
rect 444 740 446 798
rect 486 788 492 789
rect 486 784 487 788
rect 491 784 492 788
rect 486 783 492 784
rect 566 788 572 789
rect 566 784 567 788
rect 571 784 572 788
rect 566 783 572 784
rect 646 788 652 789
rect 646 784 647 788
rect 651 784 652 788
rect 646 783 652 784
rect 487 782 491 783
rect 487 777 491 778
rect 495 782 499 783
rect 495 777 499 778
rect 567 782 571 783
rect 567 777 571 778
rect 639 782 643 783
rect 639 777 643 778
rect 647 782 651 783
rect 647 777 651 778
rect 494 776 500 777
rect 494 772 495 776
rect 499 772 500 776
rect 494 771 500 772
rect 566 776 572 777
rect 566 772 567 776
rect 571 772 572 776
rect 566 771 572 772
rect 638 776 644 777
rect 638 772 639 776
rect 643 772 644 776
rect 638 771 644 772
rect 672 768 674 818
rect 728 817 730 829
rect 726 816 732 817
rect 726 812 727 816
rect 731 812 732 816
rect 726 811 732 812
rect 756 804 758 830
rect 767 829 771 830
rect 799 834 803 835
rect 799 829 803 830
rect 831 834 835 835
rect 831 829 835 830
rect 863 834 867 835
rect 863 829 867 830
rect 887 834 891 835
rect 887 829 891 830
rect 927 834 931 835
rect 936 832 938 858
rect 942 852 948 853
rect 942 848 943 852
rect 947 848 948 852
rect 942 847 948 848
rect 1006 852 1012 853
rect 1006 848 1007 852
rect 1011 848 1012 852
rect 1006 847 1012 848
rect 1046 852 1052 853
rect 1046 848 1047 852
rect 1051 848 1052 852
rect 1046 847 1052 848
rect 944 835 946 847
rect 1008 835 1010 847
rect 1048 835 1050 847
rect 1056 844 1058 858
rect 1064 844 1066 873
rect 1094 873 1095 877
rect 1099 873 1100 877
rect 1266 875 1267 879
rect 1271 875 1272 879
rect 1266 874 1272 875
rect 1334 879 1340 880
rect 1334 875 1335 879
rect 1339 875 1340 879
rect 1334 874 1340 875
rect 1378 879 1384 880
rect 1378 875 1379 879
rect 1383 875 1384 879
rect 1378 874 1384 875
rect 1094 872 1100 873
rect 1134 867 1140 868
rect 1134 863 1135 867
rect 1139 863 1140 867
rect 1134 862 1140 863
rect 1238 864 1244 865
rect 1094 860 1100 861
rect 1094 856 1095 860
rect 1099 856 1100 860
rect 1136 859 1138 862
rect 1238 860 1239 864
rect 1243 860 1244 864
rect 1238 859 1244 860
rect 1318 864 1324 865
rect 1318 860 1319 864
rect 1323 860 1324 864
rect 1318 859 1324 860
rect 1094 855 1100 856
rect 1135 858 1139 859
rect 1054 843 1060 844
rect 1054 839 1055 843
rect 1059 839 1060 843
rect 1054 838 1060 839
rect 1062 843 1068 844
rect 1062 839 1063 843
rect 1067 839 1068 843
rect 1062 838 1068 839
rect 1096 835 1098 855
rect 1135 853 1139 854
rect 1159 858 1163 859
rect 1159 853 1163 854
rect 1239 858 1243 859
rect 1239 853 1243 854
rect 1247 858 1251 859
rect 1247 853 1251 854
rect 1319 858 1323 859
rect 1319 853 1323 854
rect 1359 858 1363 859
rect 1359 853 1363 854
rect 1136 850 1138 853
rect 1158 852 1164 853
rect 1134 849 1140 850
rect 1134 845 1135 849
rect 1139 845 1140 849
rect 1158 848 1159 852
rect 1163 848 1164 852
rect 1158 847 1164 848
rect 1246 852 1252 853
rect 1246 848 1247 852
rect 1251 848 1252 852
rect 1246 847 1252 848
rect 1358 852 1364 853
rect 1358 848 1359 852
rect 1363 848 1364 852
rect 1358 847 1364 848
rect 1134 844 1140 845
rect 1388 836 1390 894
rect 1408 893 1410 905
rect 1496 893 1498 905
rect 1584 893 1586 905
rect 1608 900 1610 934
rect 1614 928 1620 929
rect 1614 924 1615 928
rect 1619 924 1620 928
rect 1614 923 1620 924
rect 1686 928 1692 929
rect 1686 924 1687 928
rect 1691 924 1692 928
rect 1686 923 1692 924
rect 1750 928 1756 929
rect 1750 924 1751 928
rect 1755 924 1756 928
rect 1750 923 1756 924
rect 1616 911 1618 923
rect 1688 911 1690 923
rect 1752 911 1754 923
rect 1780 920 1782 986
rect 2118 979 2124 980
rect 1790 976 1796 977
rect 1790 972 1791 976
rect 1795 972 1796 976
rect 1790 971 1796 972
rect 1878 976 1884 977
rect 1878 972 1879 976
rect 1883 972 1884 976
rect 1878 971 1884 972
rect 1966 976 1972 977
rect 1966 972 1967 976
rect 1971 972 1972 976
rect 1966 971 1972 972
rect 2062 976 2068 977
rect 2062 972 2063 976
rect 2067 972 2068 976
rect 2118 975 2119 979
rect 2123 975 2124 979
rect 2118 974 2124 975
rect 2062 971 2068 972
rect 1792 963 1794 971
rect 1880 963 1882 971
rect 1968 963 1970 971
rect 2064 963 2066 971
rect 2120 963 2122 974
rect 1791 962 1795 963
rect 1791 957 1795 958
rect 1815 962 1819 963
rect 1815 957 1819 958
rect 1879 962 1883 963
rect 1879 957 1883 958
rect 1951 962 1955 963
rect 1951 957 1955 958
rect 1967 962 1971 963
rect 1967 957 1971 958
rect 2023 962 2027 963
rect 2023 957 2027 958
rect 2063 962 2067 963
rect 2063 957 2067 958
rect 2071 962 2075 963
rect 2071 957 2075 958
rect 2119 962 2123 963
rect 2119 957 2123 958
rect 1814 956 1820 957
rect 1814 952 1815 956
rect 1819 952 1820 956
rect 1814 951 1820 952
rect 1878 956 1884 957
rect 1878 952 1879 956
rect 1883 952 1884 956
rect 1878 951 1884 952
rect 1950 956 1956 957
rect 1950 952 1951 956
rect 1955 952 1956 956
rect 1950 951 1956 952
rect 2022 956 2028 957
rect 2022 952 2023 956
rect 2027 952 2028 956
rect 2022 951 2028 952
rect 2070 956 2076 957
rect 2070 952 2071 956
rect 2075 952 2076 956
rect 2120 954 2122 957
rect 2070 951 2076 952
rect 2118 953 2124 954
rect 2118 949 2119 953
rect 2123 949 2124 953
rect 2118 948 2124 949
rect 1838 947 1844 948
rect 1838 943 1839 947
rect 1843 943 1844 947
rect 1838 942 1844 943
rect 1814 928 1820 929
rect 1814 924 1815 928
rect 1819 924 1820 928
rect 1814 923 1820 924
rect 1778 919 1784 920
rect 1778 915 1779 919
rect 1783 915 1784 919
rect 1778 914 1784 915
rect 1816 911 1818 923
rect 1840 920 1842 942
rect 1886 939 1892 940
rect 1886 935 1887 939
rect 1891 935 1892 939
rect 1886 934 1892 935
rect 1966 939 1972 940
rect 1966 935 1967 939
rect 1971 935 1972 939
rect 1966 934 1972 935
rect 2038 939 2044 940
rect 2038 935 2039 939
rect 2043 935 2044 939
rect 2038 934 2044 935
rect 2046 939 2052 940
rect 2046 935 2047 939
rect 2051 935 2052 939
rect 2046 934 2052 935
rect 2094 939 2100 940
rect 2094 935 2095 939
rect 2099 935 2100 939
rect 2094 934 2100 935
rect 2118 936 2124 937
rect 1878 928 1884 929
rect 1878 924 1879 928
rect 1883 924 1884 928
rect 1878 923 1884 924
rect 1838 919 1844 920
rect 1838 915 1839 919
rect 1843 915 1844 919
rect 1838 914 1844 915
rect 1880 911 1882 923
rect 1888 920 1890 934
rect 1950 928 1956 929
rect 1950 924 1951 928
rect 1955 924 1956 928
rect 1950 923 1956 924
rect 1886 919 1892 920
rect 1886 915 1887 919
rect 1891 915 1892 919
rect 1886 914 1892 915
rect 1952 911 1954 923
rect 1968 920 1970 934
rect 2022 928 2028 929
rect 2022 924 2023 928
rect 2027 924 2028 928
rect 2022 923 2028 924
rect 1966 919 1972 920
rect 1966 915 1967 919
rect 1971 915 1972 919
rect 1966 914 1972 915
rect 2024 911 2026 923
rect 2040 920 2042 934
rect 2038 919 2044 920
rect 2038 915 2039 919
rect 2043 915 2044 919
rect 2038 914 2044 915
rect 1615 910 1619 911
rect 1615 905 1619 906
rect 1663 910 1667 911
rect 1663 905 1667 906
rect 1687 910 1691 911
rect 1687 905 1691 906
rect 1743 910 1747 911
rect 1743 905 1747 906
rect 1751 910 1755 911
rect 1751 905 1755 906
rect 1815 910 1819 911
rect 1815 905 1819 906
rect 1879 910 1883 911
rect 1879 905 1883 906
rect 1887 910 1891 911
rect 1887 905 1891 906
rect 1951 910 1955 911
rect 1951 905 1955 906
rect 2023 910 2027 911
rect 2023 905 2027 906
rect 1598 899 1604 900
rect 1598 895 1599 899
rect 1603 895 1604 899
rect 1598 894 1604 895
rect 1606 899 1612 900
rect 1606 895 1607 899
rect 1611 895 1612 899
rect 1606 894 1612 895
rect 1406 892 1412 893
rect 1406 888 1407 892
rect 1411 888 1412 892
rect 1406 887 1412 888
rect 1494 892 1500 893
rect 1494 888 1495 892
rect 1499 888 1500 892
rect 1494 887 1500 888
rect 1582 892 1588 893
rect 1582 888 1583 892
rect 1587 888 1588 892
rect 1582 887 1588 888
rect 1600 880 1602 894
rect 1664 893 1666 905
rect 1744 893 1746 905
rect 1758 899 1764 900
rect 1758 895 1759 899
rect 1763 895 1764 899
rect 1758 894 1764 895
rect 1806 899 1812 900
rect 1806 895 1807 899
rect 1811 895 1812 899
rect 1806 894 1812 895
rect 1662 892 1668 893
rect 1662 888 1663 892
rect 1667 888 1668 892
rect 1662 887 1668 888
rect 1742 892 1748 893
rect 1742 888 1743 892
rect 1747 888 1748 892
rect 1742 887 1748 888
rect 1760 880 1762 894
rect 1482 879 1488 880
rect 1482 875 1483 879
rect 1487 875 1488 879
rect 1482 874 1488 875
rect 1598 879 1604 880
rect 1598 875 1599 879
rect 1603 875 1604 879
rect 1598 874 1604 875
rect 1734 879 1740 880
rect 1734 875 1735 879
rect 1739 875 1740 879
rect 1734 874 1740 875
rect 1758 879 1764 880
rect 1758 875 1759 879
rect 1763 875 1764 879
rect 1758 874 1764 875
rect 1406 864 1412 865
rect 1406 860 1407 864
rect 1411 860 1412 864
rect 1406 859 1412 860
rect 1407 858 1411 859
rect 1407 853 1411 854
rect 1455 858 1459 859
rect 1455 853 1459 854
rect 1454 852 1460 853
rect 1454 848 1455 852
rect 1459 848 1460 852
rect 1454 847 1460 848
rect 1262 835 1268 836
rect 943 834 947 835
rect 927 829 931 830
rect 934 831 940 832
rect 800 817 802 829
rect 814 823 820 824
rect 814 819 815 823
rect 819 819 820 823
rect 814 818 820 819
rect 798 816 804 817
rect 798 812 799 816
rect 803 812 804 816
rect 798 811 804 812
rect 816 804 818 818
rect 864 817 866 829
rect 886 823 892 824
rect 886 819 887 823
rect 891 819 892 823
rect 886 818 892 819
rect 862 816 868 817
rect 862 812 863 816
rect 867 812 868 816
rect 862 811 868 812
rect 754 803 760 804
rect 754 799 755 803
rect 759 799 760 803
rect 754 798 760 799
rect 814 803 820 804
rect 814 799 815 803
rect 819 799 820 803
rect 814 798 820 799
rect 726 788 732 789
rect 726 784 727 788
rect 731 784 732 788
rect 726 783 732 784
rect 798 788 804 789
rect 798 784 799 788
rect 803 784 804 788
rect 798 783 804 784
rect 862 788 868 789
rect 862 784 863 788
rect 867 784 868 788
rect 862 783 868 784
rect 703 782 707 783
rect 703 777 707 778
rect 727 782 731 783
rect 727 777 731 778
rect 759 782 763 783
rect 759 777 763 778
rect 799 782 803 783
rect 799 777 803 778
rect 815 782 819 783
rect 815 777 819 778
rect 863 782 867 783
rect 863 777 867 778
rect 702 776 708 777
rect 702 772 703 776
rect 707 772 708 776
rect 702 771 708 772
rect 758 776 764 777
rect 758 772 759 776
rect 763 772 764 776
rect 758 771 764 772
rect 814 776 820 777
rect 814 772 815 776
rect 819 772 820 776
rect 814 771 820 772
rect 862 776 868 777
rect 862 772 863 776
rect 867 772 868 776
rect 862 771 868 772
rect 888 768 890 818
rect 928 817 930 829
rect 934 827 935 831
rect 939 827 940 831
rect 943 829 947 830
rect 999 834 1003 835
rect 999 829 1003 830
rect 1007 834 1011 835
rect 1007 829 1011 830
rect 1047 834 1051 835
rect 1047 829 1051 830
rect 1095 834 1099 835
rect 1095 829 1099 830
rect 1134 832 1140 833
rect 934 826 940 827
rect 1000 817 1002 829
rect 1048 817 1050 829
rect 1070 823 1076 824
rect 1070 819 1071 823
rect 1075 819 1076 823
rect 1070 818 1076 819
rect 926 816 932 817
rect 926 812 927 816
rect 931 812 932 816
rect 926 811 932 812
rect 998 816 1004 817
rect 998 812 999 816
rect 1003 812 1004 816
rect 998 811 1004 812
rect 1046 816 1052 817
rect 1046 812 1047 816
rect 1051 812 1052 816
rect 1046 811 1052 812
rect 1014 803 1020 804
rect 1014 799 1015 803
rect 1019 799 1020 803
rect 1014 798 1020 799
rect 926 788 932 789
rect 926 784 927 788
rect 931 784 932 788
rect 926 783 932 784
rect 998 788 1004 789
rect 998 784 999 788
rect 1003 784 1004 788
rect 998 783 1004 784
rect 911 782 915 783
rect 911 777 915 778
rect 927 782 931 783
rect 927 777 931 778
rect 959 782 963 783
rect 959 777 963 778
rect 999 782 1003 783
rect 999 777 1003 778
rect 1007 782 1011 783
rect 1007 777 1011 778
rect 910 776 916 777
rect 910 772 911 776
rect 915 772 916 776
rect 910 771 916 772
rect 958 776 964 777
rect 958 772 959 776
rect 963 772 964 776
rect 958 771 964 772
rect 1006 776 1012 777
rect 1006 772 1007 776
rect 1011 772 1012 776
rect 1006 771 1012 772
rect 670 767 676 768
rect 670 763 671 767
rect 675 763 676 767
rect 670 762 676 763
rect 886 767 892 768
rect 886 763 887 767
rect 891 763 892 767
rect 886 762 892 763
rect 582 759 588 760
rect 582 755 583 759
rect 587 755 588 759
rect 582 754 588 755
rect 662 759 668 760
rect 662 755 663 759
rect 667 755 668 759
rect 662 754 668 755
rect 750 759 756 760
rect 750 755 751 759
rect 755 755 756 759
rect 750 754 756 755
rect 878 759 884 760
rect 878 755 879 759
rect 883 755 884 759
rect 878 754 884 755
rect 926 759 932 760
rect 926 755 927 759
rect 931 755 932 759
rect 926 754 932 755
rect 494 748 500 749
rect 494 744 495 748
rect 499 744 500 748
rect 494 743 500 744
rect 566 748 572 749
rect 566 744 567 748
rect 571 744 572 748
rect 566 743 572 744
rect 442 739 448 740
rect 442 735 443 739
rect 447 735 448 739
rect 442 734 448 735
rect 496 731 498 743
rect 558 739 564 740
rect 558 735 559 739
rect 563 735 564 739
rect 558 734 564 735
rect 215 730 219 731
rect 215 725 219 726
rect 239 730 243 731
rect 239 725 243 726
rect 279 730 283 731
rect 279 725 283 726
rect 311 730 315 731
rect 311 725 315 726
rect 351 730 355 731
rect 351 725 355 726
rect 391 730 395 731
rect 391 725 395 726
rect 423 730 427 731
rect 423 725 427 726
rect 471 730 475 731
rect 471 725 475 726
rect 495 730 499 731
rect 495 725 499 726
rect 543 730 547 731
rect 543 725 547 726
rect 202 719 208 720
rect 202 715 203 719
rect 207 715 208 719
rect 202 714 208 715
rect 210 719 216 720
rect 210 715 211 719
rect 215 715 216 719
rect 210 714 216 715
rect 174 712 180 713
rect 174 708 175 712
rect 179 708 180 712
rect 174 707 180 708
rect 110 704 116 705
rect 110 700 111 704
rect 115 700 116 704
rect 212 700 214 714
rect 240 713 242 725
rect 312 713 314 725
rect 392 713 394 725
rect 418 719 424 720
rect 418 715 419 719
rect 423 715 424 719
rect 418 714 424 715
rect 426 719 432 720
rect 426 715 427 719
rect 431 715 432 719
rect 426 714 432 715
rect 238 712 244 713
rect 238 708 239 712
rect 243 708 244 712
rect 238 707 244 708
rect 310 712 316 713
rect 310 708 311 712
rect 315 708 316 712
rect 310 707 316 708
rect 390 712 396 713
rect 390 708 391 712
rect 395 708 396 712
rect 390 707 396 708
rect 110 699 116 700
rect 210 699 216 700
rect 210 695 211 699
rect 215 695 216 699
rect 210 694 216 695
rect 298 699 304 700
rect 298 695 299 699
rect 303 695 304 699
rect 298 694 304 695
rect 110 687 116 688
rect 110 683 111 687
rect 115 683 116 687
rect 110 682 116 683
rect 174 684 180 685
rect 112 679 114 682
rect 174 680 175 684
rect 179 680 180 684
rect 174 679 180 680
rect 238 684 244 685
rect 238 680 239 684
rect 243 680 244 684
rect 238 679 244 680
rect 111 678 115 679
rect 111 673 115 674
rect 135 678 139 679
rect 135 673 139 674
rect 175 678 179 679
rect 175 673 179 674
rect 215 678 219 679
rect 215 673 219 674
rect 239 678 243 679
rect 239 673 243 674
rect 271 678 275 679
rect 271 673 275 674
rect 112 670 114 673
rect 134 672 140 673
rect 110 669 116 670
rect 110 665 111 669
rect 115 665 116 669
rect 134 668 135 672
rect 139 668 140 672
rect 134 667 140 668
rect 174 672 180 673
rect 174 668 175 672
rect 179 668 180 672
rect 174 667 180 668
rect 214 672 220 673
rect 214 668 215 672
rect 219 668 220 672
rect 214 667 220 668
rect 270 672 276 673
rect 270 668 271 672
rect 275 668 276 672
rect 270 667 276 668
rect 110 664 116 665
rect 162 655 168 656
rect 110 652 116 653
rect 110 648 111 652
rect 115 648 116 652
rect 162 651 163 655
rect 167 651 168 655
rect 162 650 168 651
rect 182 655 188 656
rect 182 651 183 655
rect 187 651 188 655
rect 182 650 188 651
rect 222 655 228 656
rect 222 651 223 655
rect 227 651 228 655
rect 222 650 228 651
rect 110 647 116 648
rect 112 619 114 647
rect 134 644 140 645
rect 134 640 135 644
rect 139 640 140 644
rect 134 639 140 640
rect 136 619 138 639
rect 111 618 115 619
rect 111 613 115 614
rect 135 618 139 619
rect 164 616 166 650
rect 174 644 180 645
rect 174 640 175 644
rect 179 640 180 644
rect 174 639 180 640
rect 176 619 178 639
rect 184 636 186 650
rect 214 644 220 645
rect 214 640 215 644
rect 219 640 220 644
rect 214 639 220 640
rect 182 635 188 636
rect 182 631 183 635
rect 187 631 188 635
rect 182 630 188 631
rect 216 619 218 639
rect 224 636 226 650
rect 270 644 276 645
rect 270 640 271 644
rect 275 640 276 644
rect 270 639 276 640
rect 222 635 228 636
rect 222 631 223 635
rect 227 631 228 635
rect 222 630 228 631
rect 272 619 274 639
rect 300 636 302 694
rect 310 684 316 685
rect 310 680 311 684
rect 315 680 316 684
rect 310 679 316 680
rect 390 684 396 685
rect 390 680 391 684
rect 395 680 396 684
rect 390 679 396 680
rect 311 678 315 679
rect 311 673 315 674
rect 335 678 339 679
rect 335 673 339 674
rect 391 678 395 679
rect 391 673 395 674
rect 399 678 403 679
rect 399 673 403 674
rect 334 672 340 673
rect 334 668 335 672
rect 339 668 340 672
rect 334 667 340 668
rect 398 672 404 673
rect 398 668 399 672
rect 403 668 404 672
rect 398 667 404 668
rect 420 656 422 714
rect 428 700 430 714
rect 472 713 474 725
rect 544 713 546 725
rect 470 712 476 713
rect 470 708 471 712
rect 475 708 476 712
rect 470 707 476 708
rect 542 712 548 713
rect 542 708 543 712
rect 547 708 548 712
rect 542 707 548 708
rect 560 700 562 734
rect 568 731 570 743
rect 584 740 586 754
rect 638 748 644 749
rect 638 744 639 748
rect 643 744 644 748
rect 638 743 644 744
rect 582 739 588 740
rect 582 735 583 739
rect 587 735 588 739
rect 582 734 588 735
rect 640 731 642 743
rect 664 732 666 754
rect 702 748 708 749
rect 702 744 703 748
rect 707 744 708 748
rect 702 743 708 744
rect 662 731 668 732
rect 704 731 706 743
rect 752 740 754 754
rect 758 748 764 749
rect 758 744 759 748
rect 763 744 764 748
rect 758 743 764 744
rect 814 748 820 749
rect 814 744 815 748
rect 819 744 820 748
rect 814 743 820 744
rect 862 748 868 749
rect 862 744 863 748
rect 867 744 868 748
rect 862 743 868 744
rect 750 739 756 740
rect 750 735 751 739
rect 755 735 756 739
rect 750 734 756 735
rect 760 731 762 743
rect 816 731 818 743
rect 822 739 828 740
rect 822 735 823 739
rect 827 735 828 739
rect 822 734 828 735
rect 567 730 571 731
rect 567 725 571 726
rect 615 730 619 731
rect 615 725 619 726
rect 639 730 643 731
rect 662 727 663 731
rect 667 727 668 731
rect 662 726 668 727
rect 679 730 683 731
rect 639 725 643 726
rect 679 725 683 726
rect 703 730 707 731
rect 703 725 707 726
rect 735 730 739 731
rect 735 725 739 726
rect 759 730 763 731
rect 759 725 763 726
rect 799 730 803 731
rect 799 725 803 726
rect 815 730 819 731
rect 815 725 819 726
rect 616 713 618 725
rect 680 713 682 725
rect 694 719 700 720
rect 694 715 695 719
rect 699 715 700 719
rect 694 714 700 715
rect 726 719 732 720
rect 726 715 727 719
rect 731 715 732 719
rect 726 714 732 715
rect 614 712 620 713
rect 614 708 615 712
rect 619 708 620 712
rect 614 707 620 708
rect 678 712 684 713
rect 678 708 679 712
rect 683 708 684 712
rect 678 707 684 708
rect 696 700 698 714
rect 426 699 432 700
rect 426 695 427 699
rect 431 695 432 699
rect 426 694 432 695
rect 558 699 564 700
rect 558 695 559 699
rect 563 695 564 699
rect 558 694 564 695
rect 694 699 700 700
rect 694 695 695 699
rect 699 695 700 699
rect 694 694 700 695
rect 470 684 476 685
rect 470 680 471 684
rect 475 680 476 684
rect 470 679 476 680
rect 542 684 548 685
rect 542 680 543 684
rect 547 680 548 684
rect 542 679 548 680
rect 614 684 620 685
rect 614 680 615 684
rect 619 680 620 684
rect 614 679 620 680
rect 678 684 684 685
rect 678 680 679 684
rect 683 680 684 684
rect 678 679 684 680
rect 463 678 467 679
rect 463 673 467 674
rect 471 678 475 679
rect 471 673 475 674
rect 527 678 531 679
rect 527 673 531 674
rect 543 678 547 679
rect 543 673 547 674
rect 591 678 595 679
rect 591 673 595 674
rect 615 678 619 679
rect 615 673 619 674
rect 647 678 651 679
rect 647 673 651 674
rect 679 678 683 679
rect 679 673 683 674
rect 703 678 707 679
rect 703 673 707 674
rect 462 672 468 673
rect 462 668 463 672
rect 467 668 468 672
rect 462 667 468 668
rect 526 672 532 673
rect 526 668 527 672
rect 531 668 532 672
rect 526 667 532 668
rect 590 672 596 673
rect 590 668 591 672
rect 595 668 596 672
rect 590 667 596 668
rect 646 672 652 673
rect 646 668 647 672
rect 651 668 652 672
rect 646 667 652 668
rect 702 672 708 673
rect 702 668 703 672
rect 707 668 708 672
rect 702 667 708 668
rect 728 656 730 714
rect 736 713 738 725
rect 800 713 802 725
rect 734 712 740 713
rect 734 708 735 712
rect 739 708 740 712
rect 734 707 740 708
rect 798 712 804 713
rect 798 708 799 712
rect 803 708 804 712
rect 798 707 804 708
rect 824 700 826 734
rect 864 731 866 743
rect 880 740 882 754
rect 910 748 916 749
rect 910 744 911 748
rect 915 744 916 748
rect 910 743 916 744
rect 878 739 884 740
rect 878 735 879 739
rect 883 735 884 739
rect 878 734 884 735
rect 912 731 914 743
rect 928 740 930 754
rect 958 748 964 749
rect 958 744 959 748
rect 963 744 964 748
rect 958 743 964 744
rect 1006 748 1012 749
rect 1006 744 1007 748
rect 1011 744 1012 748
rect 1006 743 1012 744
rect 926 739 932 740
rect 926 735 927 739
rect 931 735 932 739
rect 926 734 932 735
rect 960 731 962 743
rect 1008 731 1010 743
rect 1016 740 1018 798
rect 1046 788 1052 789
rect 1046 784 1047 788
rect 1051 784 1052 788
rect 1046 783 1052 784
rect 1047 782 1051 783
rect 1047 777 1051 778
rect 1046 776 1052 777
rect 1046 772 1047 776
rect 1051 772 1052 776
rect 1046 771 1052 772
rect 1072 760 1074 818
rect 1096 809 1098 829
rect 1134 828 1135 832
rect 1139 828 1140 832
rect 1262 831 1263 835
rect 1267 831 1268 835
rect 1262 830 1268 831
rect 1374 835 1380 836
rect 1374 831 1375 835
rect 1379 831 1380 835
rect 1374 830 1380 831
rect 1386 835 1392 836
rect 1386 831 1387 835
rect 1391 831 1392 835
rect 1386 830 1392 831
rect 1462 835 1468 836
rect 1462 831 1463 835
rect 1467 831 1468 835
rect 1462 830 1468 831
rect 1134 827 1140 828
rect 1094 808 1100 809
rect 1094 804 1095 808
rect 1099 804 1100 808
rect 1136 807 1138 827
rect 1158 824 1164 825
rect 1158 820 1159 824
rect 1163 820 1164 824
rect 1158 819 1164 820
rect 1246 824 1252 825
rect 1246 820 1247 824
rect 1251 820 1252 824
rect 1246 819 1252 820
rect 1160 807 1162 819
rect 1182 815 1188 816
rect 1182 811 1183 815
rect 1187 811 1188 815
rect 1182 810 1188 811
rect 1094 803 1100 804
rect 1135 806 1139 807
rect 1135 801 1139 802
rect 1159 806 1163 807
rect 1159 801 1163 802
rect 1094 791 1100 792
rect 1094 787 1095 791
rect 1099 787 1100 791
rect 1094 786 1100 787
rect 1096 783 1098 786
rect 1095 782 1099 783
rect 1136 781 1138 801
rect 1160 789 1162 801
rect 1158 788 1164 789
rect 1158 784 1159 788
rect 1163 784 1164 788
rect 1158 783 1164 784
rect 1095 777 1099 778
rect 1134 780 1140 781
rect 1096 774 1098 777
rect 1134 776 1135 780
rect 1139 776 1140 780
rect 1184 776 1186 810
rect 1248 807 1250 819
rect 1264 816 1266 830
rect 1358 824 1364 825
rect 1358 820 1359 824
rect 1363 820 1364 824
rect 1358 819 1364 820
rect 1262 815 1268 816
rect 1262 811 1263 815
rect 1267 811 1268 815
rect 1262 810 1268 811
rect 1360 807 1362 819
rect 1376 816 1378 830
rect 1454 824 1460 825
rect 1454 820 1455 824
rect 1459 820 1460 824
rect 1454 819 1460 820
rect 1374 815 1380 816
rect 1374 811 1375 815
rect 1379 811 1380 815
rect 1374 810 1380 811
rect 1456 807 1458 819
rect 1247 806 1251 807
rect 1247 801 1251 802
rect 1279 806 1283 807
rect 1279 801 1283 802
rect 1359 806 1363 807
rect 1359 801 1363 802
rect 1407 806 1411 807
rect 1407 801 1411 802
rect 1455 806 1459 807
rect 1455 801 1459 802
rect 1280 789 1282 801
rect 1408 789 1410 801
rect 1464 796 1466 830
rect 1484 816 1486 874
rect 1494 864 1500 865
rect 1494 860 1495 864
rect 1499 860 1500 864
rect 1494 859 1500 860
rect 1582 864 1588 865
rect 1582 860 1583 864
rect 1587 860 1588 864
rect 1582 859 1588 860
rect 1662 864 1668 865
rect 1662 860 1663 864
rect 1667 860 1668 864
rect 1662 859 1668 860
rect 1495 858 1499 859
rect 1495 853 1499 854
rect 1543 858 1547 859
rect 1543 853 1547 854
rect 1583 858 1587 859
rect 1583 853 1587 854
rect 1631 858 1635 859
rect 1631 853 1635 854
rect 1663 858 1667 859
rect 1663 853 1667 854
rect 1711 858 1715 859
rect 1711 853 1715 854
rect 1542 852 1548 853
rect 1542 848 1543 852
rect 1547 848 1548 852
rect 1542 847 1548 848
rect 1630 852 1636 853
rect 1630 848 1631 852
rect 1635 848 1636 852
rect 1630 847 1636 848
rect 1710 852 1716 853
rect 1710 848 1711 852
rect 1715 848 1716 852
rect 1710 847 1716 848
rect 1558 835 1564 836
rect 1558 831 1559 835
rect 1563 831 1564 835
rect 1558 830 1564 831
rect 1542 824 1548 825
rect 1542 820 1543 824
rect 1547 820 1548 824
rect 1542 819 1548 820
rect 1482 815 1488 816
rect 1482 811 1483 815
rect 1487 811 1488 815
rect 1482 810 1488 811
rect 1544 807 1546 819
rect 1519 806 1523 807
rect 1519 801 1523 802
rect 1543 806 1547 807
rect 1543 801 1547 802
rect 1422 795 1428 796
rect 1422 791 1423 795
rect 1427 791 1428 795
rect 1422 790 1428 791
rect 1462 795 1468 796
rect 1462 791 1463 795
rect 1467 791 1468 795
rect 1462 790 1468 791
rect 1278 788 1284 789
rect 1278 784 1279 788
rect 1283 784 1284 788
rect 1278 783 1284 784
rect 1406 788 1412 789
rect 1406 784 1407 788
rect 1411 784 1412 788
rect 1406 783 1412 784
rect 1424 776 1426 790
rect 1520 789 1522 801
rect 1560 796 1562 830
rect 1630 824 1636 825
rect 1630 820 1631 824
rect 1635 820 1636 824
rect 1630 819 1636 820
rect 1710 824 1716 825
rect 1710 820 1711 824
rect 1715 820 1716 824
rect 1710 819 1716 820
rect 1632 807 1634 819
rect 1712 807 1714 819
rect 1736 816 1738 874
rect 1742 864 1748 865
rect 1742 860 1743 864
rect 1747 860 1748 864
rect 1742 859 1748 860
rect 1743 858 1747 859
rect 1743 853 1747 854
rect 1783 858 1787 859
rect 1783 853 1787 854
rect 1782 852 1788 853
rect 1782 848 1783 852
rect 1787 848 1788 852
rect 1782 847 1788 848
rect 1808 836 1810 894
rect 1816 893 1818 905
rect 1888 893 1890 905
rect 1902 899 1908 900
rect 1902 895 1903 899
rect 1907 895 1908 899
rect 1902 894 1908 895
rect 1814 892 1820 893
rect 1814 888 1815 892
rect 1819 888 1820 892
rect 1814 887 1820 888
rect 1886 892 1892 893
rect 1886 888 1887 892
rect 1891 888 1892 892
rect 1886 887 1892 888
rect 1904 880 1906 894
rect 1952 893 1954 905
rect 1966 899 1972 900
rect 1966 895 1967 899
rect 1971 895 1972 899
rect 1966 894 1972 895
rect 1950 892 1956 893
rect 1950 888 1951 892
rect 1955 888 1956 892
rect 1950 887 1956 888
rect 1968 880 1970 894
rect 2024 893 2026 905
rect 2048 900 2050 934
rect 2070 928 2076 929
rect 2070 924 2071 928
rect 2075 924 2076 928
rect 2070 923 2076 924
rect 2072 911 2074 923
rect 2071 910 2075 911
rect 2071 905 2075 906
rect 2038 899 2044 900
rect 2038 895 2039 899
rect 2043 895 2044 899
rect 2038 894 2044 895
rect 2046 899 2052 900
rect 2046 895 2047 899
rect 2051 895 2052 899
rect 2046 894 2052 895
rect 2022 892 2028 893
rect 2022 888 2023 892
rect 2027 888 2028 892
rect 2022 887 2028 888
rect 2040 880 2042 894
rect 2072 893 2074 905
rect 2096 900 2098 934
rect 2118 932 2119 936
rect 2123 932 2124 936
rect 2118 931 2124 932
rect 2120 911 2122 931
rect 2119 910 2123 911
rect 2119 905 2123 906
rect 2094 899 2100 900
rect 2094 895 2095 899
rect 2099 895 2100 899
rect 2094 894 2100 895
rect 2070 892 2076 893
rect 2070 888 2071 892
rect 2075 888 2076 892
rect 2070 887 2076 888
rect 2120 885 2122 905
rect 2118 884 2124 885
rect 2118 880 2119 884
rect 2123 880 2124 884
rect 1894 879 1900 880
rect 1894 875 1895 879
rect 1899 875 1900 879
rect 1894 874 1900 875
rect 1902 879 1908 880
rect 1902 875 1903 879
rect 1907 875 1908 879
rect 1902 874 1908 875
rect 1966 879 1972 880
rect 1966 875 1967 879
rect 1971 875 1972 879
rect 1966 874 1972 875
rect 2038 879 2044 880
rect 2038 875 2039 879
rect 2043 875 2044 879
rect 2038 874 2044 875
rect 2094 879 2100 880
rect 2118 879 2124 880
rect 2094 875 2095 879
rect 2099 875 2100 879
rect 2094 874 2100 875
rect 1814 864 1820 865
rect 1814 860 1815 864
rect 1819 860 1820 864
rect 1814 859 1820 860
rect 1886 864 1892 865
rect 1886 860 1887 864
rect 1891 860 1892 864
rect 1886 859 1892 860
rect 1815 858 1819 859
rect 1815 853 1819 854
rect 1855 858 1859 859
rect 1855 853 1859 854
rect 1887 858 1891 859
rect 1887 853 1891 854
rect 1854 852 1860 853
rect 1854 848 1855 852
rect 1859 848 1860 852
rect 1854 847 1860 848
rect 1806 835 1812 836
rect 1806 831 1807 835
rect 1811 831 1812 835
rect 1806 830 1812 831
rect 1818 835 1824 836
rect 1818 831 1819 835
rect 1823 831 1824 835
rect 1818 830 1824 831
rect 1782 824 1788 825
rect 1782 820 1783 824
rect 1787 820 1788 824
rect 1782 819 1788 820
rect 1734 815 1740 816
rect 1734 811 1735 815
rect 1739 811 1740 815
rect 1734 810 1740 811
rect 1784 807 1786 819
rect 1820 816 1822 830
rect 1854 824 1860 825
rect 1854 820 1855 824
rect 1859 820 1860 824
rect 1854 819 1860 820
rect 1818 815 1824 816
rect 1818 811 1819 815
rect 1823 811 1824 815
rect 1818 810 1824 811
rect 1856 807 1858 819
rect 1896 808 1898 874
rect 1950 864 1956 865
rect 1950 860 1951 864
rect 1955 860 1956 864
rect 1950 859 1956 860
rect 2022 864 2028 865
rect 2022 860 2023 864
rect 2027 860 2028 864
rect 2022 859 2028 860
rect 2070 864 2076 865
rect 2070 860 2071 864
rect 2075 860 2076 864
rect 2070 859 2076 860
rect 1935 858 1939 859
rect 1935 853 1939 854
rect 1951 858 1955 859
rect 1951 853 1955 854
rect 2015 858 2019 859
rect 2015 853 2019 854
rect 2023 858 2027 859
rect 2023 853 2027 854
rect 2071 858 2075 859
rect 2071 853 2075 854
rect 1934 852 1940 853
rect 1934 848 1935 852
rect 1939 848 1940 852
rect 1934 847 1940 848
rect 2014 852 2020 853
rect 2014 848 2015 852
rect 2019 848 2020 852
rect 2014 847 2020 848
rect 2070 852 2076 853
rect 2070 848 2071 852
rect 2075 848 2076 852
rect 2070 847 2076 848
rect 1934 824 1940 825
rect 1934 820 1935 824
rect 1939 820 1940 824
rect 1934 819 1940 820
rect 2014 824 2020 825
rect 2014 820 2015 824
rect 2019 820 2020 824
rect 2014 819 2020 820
rect 2070 824 2076 825
rect 2070 820 2071 824
rect 2075 820 2076 824
rect 2070 819 2076 820
rect 1910 815 1916 816
rect 1910 811 1911 815
rect 1915 811 1916 815
rect 1910 810 1916 811
rect 1894 807 1900 808
rect 1623 806 1627 807
rect 1623 801 1627 802
rect 1631 806 1635 807
rect 1631 801 1635 802
rect 1711 806 1715 807
rect 1711 801 1715 802
rect 1719 806 1723 807
rect 1719 801 1723 802
rect 1783 806 1787 807
rect 1783 801 1787 802
rect 1815 806 1819 807
rect 1815 801 1819 802
rect 1855 806 1859 807
rect 1894 803 1895 807
rect 1899 803 1900 807
rect 1894 802 1900 803
rect 1903 806 1907 807
rect 1855 801 1859 802
rect 1903 801 1907 802
rect 1558 795 1564 796
rect 1558 791 1559 795
rect 1563 791 1564 795
rect 1558 790 1564 791
rect 1566 795 1572 796
rect 1566 791 1567 795
rect 1571 791 1572 795
rect 1566 790 1572 791
rect 1518 788 1524 789
rect 1518 784 1519 788
rect 1523 784 1524 788
rect 1518 783 1524 784
rect 1568 776 1570 790
rect 1624 789 1626 801
rect 1720 789 1722 801
rect 1816 789 1818 801
rect 1904 789 1906 801
rect 1622 788 1628 789
rect 1622 784 1623 788
rect 1627 784 1628 788
rect 1622 783 1628 784
rect 1718 788 1724 789
rect 1718 784 1719 788
rect 1723 784 1724 788
rect 1718 783 1724 784
rect 1814 788 1820 789
rect 1814 784 1815 788
rect 1819 784 1820 788
rect 1814 783 1820 784
rect 1902 788 1908 789
rect 1902 784 1903 788
rect 1907 784 1908 788
rect 1902 783 1908 784
rect 1912 776 1914 810
rect 1936 807 1938 819
rect 2016 807 2018 819
rect 2072 807 2074 819
rect 2096 816 2098 874
rect 2118 867 2124 868
rect 2118 863 2119 867
rect 2123 863 2124 867
rect 2118 862 2124 863
rect 2120 859 2122 862
rect 2119 858 2123 859
rect 2119 853 2123 854
rect 2120 850 2122 853
rect 2118 849 2124 850
rect 2118 845 2119 849
rect 2123 845 2124 849
rect 2118 844 2124 845
rect 2118 832 2124 833
rect 2118 828 2119 832
rect 2123 828 2124 832
rect 2118 827 2124 828
rect 2094 815 2100 816
rect 2094 811 2095 815
rect 2099 811 2100 815
rect 2094 810 2100 811
rect 2120 807 2122 827
rect 1935 806 1939 807
rect 1935 801 1939 802
rect 1999 806 2003 807
rect 1999 801 2003 802
rect 2015 806 2019 807
rect 2015 801 2019 802
rect 2071 806 2075 807
rect 2071 801 2075 802
rect 2119 806 2123 807
rect 2119 801 2123 802
rect 1918 795 1924 796
rect 1918 791 1919 795
rect 1923 791 1924 795
rect 1918 790 1924 791
rect 1978 795 1984 796
rect 1978 791 1979 795
rect 1983 791 1984 795
rect 1978 790 1984 791
rect 1986 795 1992 796
rect 1986 791 1987 795
rect 1991 791 1992 795
rect 1986 790 1992 791
rect 1920 776 1922 790
rect 1980 776 1982 790
rect 1134 775 1140 776
rect 1182 775 1188 776
rect 1094 773 1100 774
rect 1094 769 1095 773
rect 1099 769 1100 773
rect 1182 771 1183 775
rect 1187 771 1188 775
rect 1182 770 1188 771
rect 1422 775 1428 776
rect 1422 771 1423 775
rect 1427 771 1428 775
rect 1422 770 1428 771
rect 1566 775 1572 776
rect 1566 771 1567 775
rect 1571 771 1572 775
rect 1566 770 1572 771
rect 1822 775 1828 776
rect 1822 771 1823 775
rect 1827 771 1828 775
rect 1822 770 1828 771
rect 1910 775 1916 776
rect 1910 771 1911 775
rect 1915 771 1916 775
rect 1910 770 1916 771
rect 1918 775 1924 776
rect 1918 771 1919 775
rect 1923 771 1924 775
rect 1918 770 1924 771
rect 1978 775 1984 776
rect 1978 771 1979 775
rect 1983 771 1984 775
rect 1978 770 1984 771
rect 1094 768 1100 769
rect 1134 763 1140 764
rect 1022 759 1028 760
rect 1022 755 1023 759
rect 1027 755 1028 759
rect 1022 754 1028 755
rect 1062 759 1068 760
rect 1062 755 1063 759
rect 1067 755 1068 759
rect 1062 754 1068 755
rect 1070 759 1076 760
rect 1070 755 1071 759
rect 1075 755 1076 759
rect 1134 759 1135 763
rect 1139 759 1140 763
rect 1134 758 1140 759
rect 1158 760 1164 761
rect 1070 754 1076 755
rect 1094 756 1100 757
rect 1024 740 1026 754
rect 1046 748 1052 749
rect 1046 744 1047 748
rect 1051 744 1052 748
rect 1046 743 1052 744
rect 1014 739 1020 740
rect 1014 735 1015 739
rect 1019 735 1020 739
rect 1014 734 1020 735
rect 1022 739 1028 740
rect 1022 735 1023 739
rect 1027 735 1028 739
rect 1022 734 1028 735
rect 1048 731 1050 743
rect 1064 740 1066 754
rect 1094 752 1095 756
rect 1099 752 1100 756
rect 1094 751 1100 752
rect 1136 751 1138 758
rect 1158 756 1159 760
rect 1163 756 1164 760
rect 1158 755 1164 756
rect 1278 760 1284 761
rect 1278 756 1279 760
rect 1283 756 1284 760
rect 1278 755 1284 756
rect 1406 760 1412 761
rect 1406 756 1407 760
rect 1411 756 1412 760
rect 1406 755 1412 756
rect 1518 760 1524 761
rect 1518 756 1519 760
rect 1523 756 1524 760
rect 1518 755 1524 756
rect 1622 760 1628 761
rect 1622 756 1623 760
rect 1627 756 1628 760
rect 1622 755 1628 756
rect 1718 760 1724 761
rect 1718 756 1719 760
rect 1723 756 1724 760
rect 1718 755 1724 756
rect 1814 760 1820 761
rect 1814 756 1815 760
rect 1819 756 1820 760
rect 1814 755 1820 756
rect 1160 751 1162 755
rect 1280 751 1282 755
rect 1408 751 1410 755
rect 1520 751 1522 755
rect 1624 751 1626 755
rect 1720 751 1722 755
rect 1816 751 1818 755
rect 1062 739 1068 740
rect 1062 735 1063 739
rect 1067 735 1068 739
rect 1062 734 1068 735
rect 1096 731 1098 751
rect 1135 750 1139 751
rect 1135 745 1139 746
rect 1159 750 1163 751
rect 1159 745 1163 746
rect 1279 750 1283 751
rect 1279 745 1283 746
rect 1335 750 1339 751
rect 1335 745 1339 746
rect 1375 750 1379 751
rect 1375 745 1379 746
rect 1407 750 1411 751
rect 1407 745 1411 746
rect 1415 750 1419 751
rect 1415 745 1419 746
rect 1455 750 1459 751
rect 1455 745 1459 746
rect 1503 750 1507 751
rect 1503 745 1507 746
rect 1519 750 1523 751
rect 1519 745 1523 746
rect 1551 750 1555 751
rect 1551 745 1555 746
rect 1599 750 1603 751
rect 1599 745 1603 746
rect 1623 750 1627 751
rect 1623 745 1627 746
rect 1655 750 1659 751
rect 1655 745 1659 746
rect 1711 750 1715 751
rect 1711 745 1715 746
rect 1719 750 1723 751
rect 1719 745 1723 746
rect 1767 750 1771 751
rect 1767 745 1771 746
rect 1815 750 1819 751
rect 1815 745 1819 746
rect 1136 742 1138 745
rect 1334 744 1340 745
rect 1134 741 1140 742
rect 1134 737 1135 741
rect 1139 737 1140 741
rect 1334 740 1335 744
rect 1339 740 1340 744
rect 1334 739 1340 740
rect 1374 744 1380 745
rect 1374 740 1375 744
rect 1379 740 1380 744
rect 1374 739 1380 740
rect 1414 744 1420 745
rect 1414 740 1415 744
rect 1419 740 1420 744
rect 1414 739 1420 740
rect 1454 744 1460 745
rect 1454 740 1455 744
rect 1459 740 1460 744
rect 1454 739 1460 740
rect 1502 744 1508 745
rect 1502 740 1503 744
rect 1507 740 1508 744
rect 1502 739 1508 740
rect 1550 744 1556 745
rect 1550 740 1551 744
rect 1555 740 1556 744
rect 1550 739 1556 740
rect 1598 744 1604 745
rect 1598 740 1599 744
rect 1603 740 1604 744
rect 1598 739 1604 740
rect 1654 744 1660 745
rect 1654 740 1655 744
rect 1659 740 1660 744
rect 1654 739 1660 740
rect 1710 744 1716 745
rect 1710 740 1711 744
rect 1715 740 1716 744
rect 1710 739 1716 740
rect 1766 744 1772 745
rect 1766 740 1767 744
rect 1771 740 1772 744
rect 1766 739 1772 740
rect 1134 736 1140 737
rect 1622 735 1628 736
rect 1622 731 1623 735
rect 1627 731 1628 735
rect 863 730 867 731
rect 863 725 867 726
rect 911 730 915 731
rect 911 725 915 726
rect 927 730 931 731
rect 927 725 931 726
rect 959 730 963 731
rect 959 725 963 726
rect 1007 730 1011 731
rect 1007 725 1011 726
rect 1047 730 1051 731
rect 1047 725 1051 726
rect 1095 730 1099 731
rect 1622 730 1628 731
rect 1095 725 1099 726
rect 1362 727 1368 728
rect 864 713 866 725
rect 878 719 884 720
rect 878 715 879 719
rect 883 715 884 719
rect 878 714 884 715
rect 862 712 868 713
rect 862 708 863 712
rect 867 708 868 712
rect 862 707 868 708
rect 880 700 882 714
rect 928 713 930 725
rect 942 719 948 720
rect 942 715 943 719
rect 947 715 948 719
rect 942 714 948 715
rect 926 712 932 713
rect 926 708 927 712
rect 931 708 932 712
rect 926 707 932 708
rect 944 700 946 714
rect 1096 705 1098 725
rect 1134 724 1140 725
rect 1134 720 1135 724
rect 1139 720 1140 724
rect 1362 723 1363 727
rect 1367 723 1368 727
rect 1362 722 1368 723
rect 1382 727 1388 728
rect 1382 723 1383 727
rect 1387 723 1388 727
rect 1382 722 1388 723
rect 1422 727 1428 728
rect 1422 723 1423 727
rect 1427 723 1428 727
rect 1422 722 1428 723
rect 1462 727 1468 728
rect 1462 723 1463 727
rect 1467 723 1468 727
rect 1462 722 1468 723
rect 1134 719 1140 720
rect 1094 704 1100 705
rect 1094 700 1095 704
rect 1099 700 1100 704
rect 822 699 828 700
rect 822 695 823 699
rect 827 695 828 699
rect 822 694 828 695
rect 878 699 884 700
rect 878 695 879 699
rect 883 695 884 699
rect 878 694 884 695
rect 942 699 948 700
rect 1094 699 1100 700
rect 1136 699 1138 719
rect 1334 716 1340 717
rect 1334 712 1335 716
rect 1339 712 1340 716
rect 1334 711 1340 712
rect 1336 699 1338 711
rect 942 695 943 699
rect 947 695 948 699
rect 942 694 948 695
rect 1135 698 1139 699
rect 1135 693 1139 694
rect 1247 698 1251 699
rect 1247 693 1251 694
rect 1287 698 1291 699
rect 1287 693 1291 694
rect 1335 698 1339 699
rect 1364 696 1366 722
rect 1374 716 1380 717
rect 1374 712 1375 716
rect 1379 712 1380 716
rect 1374 711 1380 712
rect 1376 699 1378 711
rect 1384 708 1386 722
rect 1414 716 1420 717
rect 1414 712 1415 716
rect 1419 712 1420 716
rect 1414 711 1420 712
rect 1382 707 1388 708
rect 1382 703 1383 707
rect 1387 703 1388 707
rect 1382 702 1388 703
rect 1416 699 1418 711
rect 1424 708 1426 722
rect 1454 716 1460 717
rect 1454 712 1455 716
rect 1459 712 1460 716
rect 1454 711 1460 712
rect 1422 707 1428 708
rect 1422 703 1423 707
rect 1427 703 1428 707
rect 1422 702 1428 703
rect 1456 699 1458 711
rect 1464 708 1466 722
rect 1502 716 1508 717
rect 1502 712 1503 716
rect 1507 712 1508 716
rect 1502 711 1508 712
rect 1550 716 1556 717
rect 1550 712 1551 716
rect 1555 712 1556 716
rect 1550 711 1556 712
rect 1598 716 1604 717
rect 1598 712 1599 716
rect 1603 712 1604 716
rect 1598 711 1604 712
rect 1462 707 1468 708
rect 1462 703 1463 707
rect 1467 703 1468 707
rect 1462 702 1468 703
rect 1504 699 1506 711
rect 1552 699 1554 711
rect 1600 699 1602 711
rect 1624 708 1626 730
rect 1678 727 1684 728
rect 1678 723 1679 727
rect 1683 723 1684 727
rect 1678 722 1684 723
rect 1758 727 1764 728
rect 1758 723 1759 727
rect 1763 723 1764 727
rect 1758 722 1764 723
rect 1654 716 1660 717
rect 1654 712 1655 716
rect 1659 712 1660 716
rect 1654 711 1660 712
rect 1622 707 1628 708
rect 1622 703 1623 707
rect 1627 703 1628 707
rect 1622 702 1628 703
rect 1656 699 1658 711
rect 1375 698 1379 699
rect 1335 693 1339 694
rect 1362 695 1368 696
rect 1094 687 1100 688
rect 734 684 740 685
rect 734 680 735 684
rect 739 680 740 684
rect 734 679 740 680
rect 798 684 804 685
rect 798 680 799 684
rect 803 680 804 684
rect 798 679 804 680
rect 862 684 868 685
rect 862 680 863 684
rect 867 680 868 684
rect 862 679 868 680
rect 926 684 932 685
rect 926 680 927 684
rect 931 680 932 684
rect 1094 683 1095 687
rect 1099 683 1100 687
rect 1094 682 1100 683
rect 926 679 932 680
rect 1096 679 1098 682
rect 735 678 739 679
rect 735 673 739 674
rect 759 678 763 679
rect 759 673 763 674
rect 799 678 803 679
rect 799 673 803 674
rect 823 678 827 679
rect 823 673 827 674
rect 863 678 867 679
rect 863 673 867 674
rect 927 678 931 679
rect 927 673 931 674
rect 1095 678 1099 679
rect 1095 673 1099 674
rect 1136 673 1138 693
rect 1248 681 1250 693
rect 1288 681 1290 693
rect 1302 687 1308 688
rect 1302 683 1303 687
rect 1307 683 1308 687
rect 1302 682 1308 683
rect 1246 680 1252 681
rect 1246 676 1247 680
rect 1251 676 1252 680
rect 1246 675 1252 676
rect 1286 680 1292 681
rect 1286 676 1287 680
rect 1291 676 1292 680
rect 1286 675 1292 676
rect 758 672 764 673
rect 758 668 759 672
rect 763 668 764 672
rect 758 667 764 668
rect 822 672 828 673
rect 822 668 823 672
rect 827 668 828 672
rect 1096 670 1098 673
rect 1134 672 1140 673
rect 822 667 828 668
rect 1094 669 1100 670
rect 1094 665 1095 669
rect 1099 665 1100 669
rect 1134 668 1135 672
rect 1139 668 1140 672
rect 1304 668 1306 682
rect 1336 681 1338 693
rect 1362 691 1363 695
rect 1367 691 1368 695
rect 1375 693 1379 694
rect 1391 698 1395 699
rect 1391 693 1395 694
rect 1415 698 1419 699
rect 1415 693 1419 694
rect 1447 698 1451 699
rect 1447 693 1451 694
rect 1455 698 1459 699
rect 1455 693 1459 694
rect 1503 698 1507 699
rect 1503 693 1507 694
rect 1511 698 1515 699
rect 1511 693 1515 694
rect 1551 698 1555 699
rect 1551 693 1555 694
rect 1583 698 1587 699
rect 1583 693 1587 694
rect 1599 698 1603 699
rect 1599 693 1603 694
rect 1655 698 1659 699
rect 1680 696 1682 722
rect 1710 716 1716 717
rect 1710 712 1711 716
rect 1715 712 1716 716
rect 1710 711 1716 712
rect 1712 699 1714 711
rect 1760 708 1762 722
rect 1766 716 1772 717
rect 1766 712 1767 716
rect 1771 712 1772 716
rect 1766 711 1772 712
rect 1758 707 1764 708
rect 1758 703 1759 707
rect 1763 703 1764 707
rect 1758 702 1764 703
rect 1768 699 1770 711
rect 1824 708 1826 770
rect 1902 760 1908 761
rect 1902 756 1903 760
rect 1907 756 1908 760
rect 1902 755 1908 756
rect 1904 751 1906 755
rect 1831 750 1835 751
rect 1831 745 1835 746
rect 1895 750 1899 751
rect 1895 745 1899 746
rect 1903 750 1907 751
rect 1903 745 1907 746
rect 1959 750 1963 751
rect 1959 745 1963 746
rect 1830 744 1836 745
rect 1830 740 1831 744
rect 1835 740 1836 744
rect 1830 739 1836 740
rect 1894 744 1900 745
rect 1894 740 1895 744
rect 1899 740 1900 744
rect 1894 739 1900 740
rect 1958 744 1964 745
rect 1958 740 1959 744
rect 1963 740 1964 744
rect 1958 739 1964 740
rect 1988 728 1990 790
rect 2000 789 2002 801
rect 2072 789 2074 801
rect 1998 788 2004 789
rect 1998 784 1999 788
rect 2003 784 2004 788
rect 1998 783 2004 784
rect 2070 788 2076 789
rect 2070 784 2071 788
rect 2075 784 2076 788
rect 2070 783 2076 784
rect 2120 781 2122 801
rect 2118 780 2124 781
rect 2118 776 2119 780
rect 2123 776 2124 780
rect 2094 775 2100 776
rect 2118 775 2124 776
rect 2094 771 2095 775
rect 2099 771 2100 775
rect 2094 770 2100 771
rect 1998 760 2004 761
rect 1998 756 1999 760
rect 2003 756 2004 760
rect 1998 755 2004 756
rect 2070 760 2076 761
rect 2070 756 2071 760
rect 2075 756 2076 760
rect 2070 755 2076 756
rect 2000 751 2002 755
rect 2072 751 2074 755
rect 1999 750 2003 751
rect 1999 745 2003 746
rect 2023 750 2027 751
rect 2023 745 2027 746
rect 2071 750 2075 751
rect 2071 745 2075 746
rect 2022 744 2028 745
rect 2022 740 2023 744
rect 2027 740 2028 744
rect 2022 739 2028 740
rect 2070 744 2076 745
rect 2070 740 2071 744
rect 2075 740 2076 744
rect 2070 739 2076 740
rect 1974 727 1980 728
rect 1974 723 1975 727
rect 1979 723 1980 727
rect 1974 722 1980 723
rect 1986 727 1992 728
rect 1986 723 1987 727
rect 1991 723 1992 727
rect 1986 722 1992 723
rect 2046 727 2052 728
rect 2046 723 2047 727
rect 2051 723 2052 727
rect 2046 722 2052 723
rect 1830 716 1836 717
rect 1830 712 1831 716
rect 1835 712 1836 716
rect 1830 711 1836 712
rect 1894 716 1900 717
rect 1894 712 1895 716
rect 1899 712 1900 716
rect 1894 711 1900 712
rect 1958 716 1964 717
rect 1958 712 1959 716
rect 1963 712 1964 716
rect 1958 711 1964 712
rect 1822 707 1828 708
rect 1822 703 1823 707
rect 1827 703 1828 707
rect 1822 702 1828 703
rect 1832 699 1834 711
rect 1896 699 1898 711
rect 1934 707 1940 708
rect 1934 703 1935 707
rect 1939 703 1940 707
rect 1934 702 1940 703
rect 1711 698 1715 699
rect 1655 693 1659 694
rect 1678 695 1684 696
rect 1362 690 1368 691
rect 1350 687 1356 688
rect 1350 683 1351 687
rect 1355 683 1356 687
rect 1350 682 1356 683
rect 1334 680 1340 681
rect 1334 676 1335 680
rect 1339 676 1340 680
rect 1334 675 1340 676
rect 1352 668 1354 682
rect 1392 681 1394 693
rect 1406 687 1412 688
rect 1406 683 1407 687
rect 1411 683 1412 687
rect 1406 682 1412 683
rect 1390 680 1396 681
rect 1390 676 1391 680
rect 1395 676 1396 680
rect 1390 675 1396 676
rect 1408 668 1410 682
rect 1448 681 1450 693
rect 1462 687 1468 688
rect 1462 683 1463 687
rect 1467 683 1468 687
rect 1462 682 1468 683
rect 1446 680 1452 681
rect 1446 676 1447 680
rect 1451 676 1452 680
rect 1446 675 1452 676
rect 1464 668 1466 682
rect 1512 681 1514 693
rect 1526 687 1532 688
rect 1526 683 1527 687
rect 1531 683 1532 687
rect 1526 682 1532 683
rect 1510 680 1516 681
rect 1510 676 1511 680
rect 1515 676 1516 680
rect 1510 675 1516 676
rect 1528 668 1530 682
rect 1584 681 1586 693
rect 1656 681 1658 693
rect 1678 691 1679 695
rect 1683 691 1684 695
rect 1711 693 1715 694
rect 1735 698 1739 699
rect 1735 693 1739 694
rect 1767 698 1771 699
rect 1767 693 1771 694
rect 1823 698 1827 699
rect 1823 693 1827 694
rect 1831 698 1835 699
rect 1831 693 1835 694
rect 1895 698 1899 699
rect 1895 693 1899 694
rect 1911 698 1915 699
rect 1911 693 1915 694
rect 1678 690 1684 691
rect 1670 687 1676 688
rect 1670 683 1671 687
rect 1675 683 1676 687
rect 1670 682 1676 683
rect 1718 687 1724 688
rect 1718 683 1719 687
rect 1723 683 1724 687
rect 1718 682 1724 683
rect 1582 680 1588 681
rect 1582 676 1583 680
rect 1587 676 1588 680
rect 1582 675 1588 676
rect 1654 680 1660 681
rect 1654 676 1655 680
rect 1659 676 1660 680
rect 1654 675 1660 676
rect 1672 668 1674 682
rect 1720 668 1722 682
rect 1736 681 1738 693
rect 1824 681 1826 693
rect 1838 687 1844 688
rect 1838 683 1839 687
rect 1843 683 1844 687
rect 1838 682 1844 683
rect 1734 680 1740 681
rect 1734 676 1735 680
rect 1739 676 1740 680
rect 1734 675 1740 676
rect 1822 680 1828 681
rect 1822 676 1823 680
rect 1827 676 1828 680
rect 1822 675 1828 676
rect 1840 668 1842 682
rect 1912 681 1914 693
rect 1910 680 1916 681
rect 1910 676 1911 680
rect 1915 676 1916 680
rect 1910 675 1916 676
rect 1936 668 1938 702
rect 1960 699 1962 711
rect 1976 708 1978 722
rect 2022 716 2028 717
rect 2022 712 2023 716
rect 2027 712 2028 716
rect 2022 711 2028 712
rect 1974 707 1980 708
rect 1974 703 1975 707
rect 1979 703 1980 707
rect 1974 702 1980 703
rect 2024 699 2026 711
rect 1959 698 1963 699
rect 1946 695 1952 696
rect 1946 691 1947 695
rect 1951 691 1952 695
rect 1959 693 1963 694
rect 1999 698 2003 699
rect 1999 693 2003 694
rect 2023 698 2027 699
rect 2023 693 2027 694
rect 1946 690 1952 691
rect 1134 667 1140 668
rect 1294 667 1300 668
rect 1094 664 1100 665
rect 846 663 852 664
rect 846 659 847 663
rect 851 659 852 663
rect 1294 663 1295 667
rect 1299 663 1300 667
rect 1294 662 1300 663
rect 1302 667 1308 668
rect 1302 663 1303 667
rect 1307 663 1308 667
rect 1302 662 1308 663
rect 1350 667 1356 668
rect 1350 663 1351 667
rect 1355 663 1356 667
rect 1350 662 1356 663
rect 1406 667 1412 668
rect 1406 663 1407 667
rect 1411 663 1412 667
rect 1406 662 1412 663
rect 1462 667 1468 668
rect 1462 663 1463 667
rect 1467 663 1468 667
rect 1462 662 1468 663
rect 1526 667 1532 668
rect 1526 663 1527 667
rect 1531 663 1532 667
rect 1526 662 1532 663
rect 1662 667 1668 668
rect 1662 663 1663 667
rect 1667 663 1668 667
rect 1662 662 1668 663
rect 1670 667 1676 668
rect 1670 663 1671 667
rect 1675 663 1676 667
rect 1670 662 1676 663
rect 1718 667 1724 668
rect 1718 663 1719 667
rect 1723 663 1724 667
rect 1718 662 1724 663
rect 1838 667 1844 668
rect 1838 663 1839 667
rect 1843 663 1844 667
rect 1838 662 1844 663
rect 1934 667 1940 668
rect 1934 663 1935 667
rect 1939 663 1940 667
rect 1934 662 1940 663
rect 846 658 852 659
rect 418 655 424 656
rect 418 651 419 655
rect 423 651 424 655
rect 418 650 424 651
rect 550 655 556 656
rect 550 651 551 655
rect 555 651 556 655
rect 550 650 556 651
rect 726 655 732 656
rect 726 651 727 655
rect 731 651 732 655
rect 726 650 732 651
rect 750 655 756 656
rect 750 651 751 655
rect 755 651 756 655
rect 750 650 756 651
rect 334 644 340 645
rect 334 640 335 644
rect 339 640 340 644
rect 334 639 340 640
rect 398 644 404 645
rect 398 640 399 644
rect 403 640 404 644
rect 398 639 404 640
rect 462 644 468 645
rect 462 640 463 644
rect 467 640 468 644
rect 462 639 468 640
rect 526 644 532 645
rect 526 640 527 644
rect 531 640 532 644
rect 526 639 532 640
rect 298 635 304 636
rect 298 631 299 635
rect 303 631 304 635
rect 298 630 304 631
rect 336 619 338 639
rect 342 635 348 636
rect 342 631 343 635
rect 347 631 348 635
rect 342 630 348 631
rect 175 618 179 619
rect 135 613 139 614
rect 162 615 168 616
rect 112 593 114 613
rect 136 601 138 613
rect 162 611 163 615
rect 167 611 168 615
rect 175 613 179 614
rect 215 618 219 619
rect 215 613 219 614
rect 255 618 259 619
rect 255 613 259 614
rect 271 618 275 619
rect 271 613 275 614
rect 303 618 307 619
rect 303 613 307 614
rect 335 618 339 619
rect 335 613 339 614
rect 162 610 168 611
rect 176 601 178 613
rect 190 607 196 608
rect 190 603 191 607
rect 195 603 196 607
rect 190 602 196 603
rect 134 600 140 601
rect 134 596 135 600
rect 139 596 140 600
rect 134 595 140 596
rect 174 600 180 601
rect 174 596 175 600
rect 179 596 180 600
rect 174 595 180 596
rect 110 592 116 593
rect 110 588 111 592
rect 115 588 116 592
rect 192 588 194 602
rect 216 601 218 613
rect 230 607 236 608
rect 230 603 231 607
rect 235 603 236 607
rect 230 602 236 603
rect 214 600 220 601
rect 214 596 215 600
rect 219 596 220 600
rect 214 595 220 596
rect 232 588 234 602
rect 256 601 258 613
rect 270 607 276 608
rect 270 603 271 607
rect 275 603 276 607
rect 270 602 276 603
rect 254 600 260 601
rect 254 596 255 600
rect 259 596 260 600
rect 254 595 260 596
rect 272 588 274 602
rect 304 601 306 613
rect 302 600 308 601
rect 302 596 303 600
rect 307 596 308 600
rect 302 595 308 596
rect 344 588 346 630
rect 400 619 402 639
rect 464 619 466 639
rect 528 619 530 639
rect 552 628 554 650
rect 590 644 596 645
rect 590 640 591 644
rect 595 640 596 644
rect 590 639 596 640
rect 646 644 652 645
rect 646 640 647 644
rect 651 640 652 644
rect 646 639 652 640
rect 702 644 708 645
rect 702 640 703 644
rect 707 640 708 644
rect 702 639 708 640
rect 550 627 556 628
rect 550 623 551 627
rect 555 623 556 627
rect 550 622 556 623
rect 592 619 594 639
rect 648 619 650 639
rect 654 635 660 636
rect 654 631 655 635
rect 659 631 660 635
rect 654 630 660 631
rect 351 618 355 619
rect 351 613 355 614
rect 399 618 403 619
rect 399 613 403 614
rect 439 618 443 619
rect 439 613 443 614
rect 463 618 467 619
rect 463 613 467 614
rect 487 618 491 619
rect 487 613 491 614
rect 527 618 531 619
rect 527 613 531 614
rect 535 618 539 619
rect 535 613 539 614
rect 583 618 587 619
rect 583 613 587 614
rect 591 618 595 619
rect 631 618 635 619
rect 591 613 595 614
rect 610 615 616 616
rect 352 601 354 613
rect 366 607 372 608
rect 366 603 367 607
rect 371 603 372 607
rect 366 602 372 603
rect 350 600 356 601
rect 350 596 351 600
rect 355 596 356 600
rect 350 595 356 596
rect 368 588 370 602
rect 400 601 402 613
rect 414 607 420 608
rect 414 603 415 607
rect 419 603 420 607
rect 414 602 420 603
rect 398 600 404 601
rect 398 596 399 600
rect 403 596 404 600
rect 398 595 404 596
rect 416 588 418 602
rect 440 601 442 613
rect 446 607 452 608
rect 446 603 447 607
rect 451 603 452 607
rect 446 602 452 603
rect 478 607 484 608
rect 478 603 479 607
rect 483 603 484 607
rect 478 602 484 603
rect 438 600 444 601
rect 438 596 439 600
rect 443 596 444 600
rect 438 595 444 596
rect 110 587 116 588
rect 158 587 164 588
rect 158 583 159 587
rect 163 583 164 587
rect 158 582 164 583
rect 190 587 196 588
rect 190 583 191 587
rect 195 583 196 587
rect 190 582 196 583
rect 230 587 236 588
rect 230 583 231 587
rect 235 583 236 587
rect 230 582 236 583
rect 270 587 276 588
rect 270 583 271 587
rect 275 583 276 587
rect 270 582 276 583
rect 342 587 348 588
rect 342 583 343 587
rect 347 583 348 587
rect 342 582 348 583
rect 366 587 372 588
rect 366 583 367 587
rect 371 583 372 587
rect 366 582 372 583
rect 414 587 420 588
rect 414 583 415 587
rect 419 583 420 587
rect 414 582 420 583
rect 110 575 116 576
rect 110 571 111 575
rect 115 571 116 575
rect 110 570 116 571
rect 134 572 140 573
rect 112 563 114 570
rect 134 568 135 572
rect 139 568 140 572
rect 134 567 140 568
rect 136 563 138 567
rect 111 562 115 563
rect 111 557 115 558
rect 135 562 139 563
rect 135 557 139 558
rect 112 554 114 557
rect 134 556 140 557
rect 110 553 116 554
rect 110 549 111 553
rect 115 549 116 553
rect 134 552 135 556
rect 139 552 140 556
rect 134 551 140 552
rect 110 548 116 549
rect 110 536 116 537
rect 110 532 111 536
rect 115 532 116 536
rect 110 531 116 532
rect 112 503 114 531
rect 134 528 140 529
rect 134 524 135 528
rect 139 524 140 528
rect 134 523 140 524
rect 136 503 138 523
rect 160 520 162 582
rect 174 572 180 573
rect 174 568 175 572
rect 179 568 180 572
rect 174 567 180 568
rect 214 572 220 573
rect 214 568 215 572
rect 219 568 220 572
rect 214 567 220 568
rect 254 572 260 573
rect 254 568 255 572
rect 259 568 260 572
rect 254 567 260 568
rect 302 572 308 573
rect 302 568 303 572
rect 307 568 308 572
rect 302 567 308 568
rect 350 572 356 573
rect 350 568 351 572
rect 355 568 356 572
rect 350 567 356 568
rect 398 572 404 573
rect 398 568 399 572
rect 403 568 404 572
rect 398 567 404 568
rect 438 572 444 573
rect 438 568 439 572
rect 443 568 444 572
rect 438 567 444 568
rect 176 563 178 567
rect 216 563 218 567
rect 256 563 258 567
rect 304 563 306 567
rect 352 563 354 567
rect 400 563 402 567
rect 440 563 442 567
rect 175 562 179 563
rect 175 557 179 558
rect 215 562 219 563
rect 215 557 219 558
rect 223 562 227 563
rect 223 557 227 558
rect 255 562 259 563
rect 255 557 259 558
rect 279 562 283 563
rect 279 557 283 558
rect 303 562 307 563
rect 303 557 307 558
rect 327 562 331 563
rect 327 557 331 558
rect 351 562 355 563
rect 351 557 355 558
rect 375 562 379 563
rect 375 557 379 558
rect 399 562 403 563
rect 399 557 403 558
rect 423 562 427 563
rect 423 557 427 558
rect 439 562 443 563
rect 439 557 443 558
rect 174 556 180 557
rect 174 552 175 556
rect 179 552 180 556
rect 174 551 180 552
rect 222 556 228 557
rect 222 552 223 556
rect 227 552 228 556
rect 222 551 228 552
rect 278 556 284 557
rect 278 552 279 556
rect 283 552 284 556
rect 278 551 284 552
rect 326 556 332 557
rect 326 552 327 556
rect 331 552 332 556
rect 326 551 332 552
rect 374 556 380 557
rect 374 552 375 556
rect 379 552 380 556
rect 374 551 380 552
rect 422 556 428 557
rect 422 552 423 556
rect 427 552 428 556
rect 422 551 428 552
rect 448 540 450 602
rect 463 562 467 563
rect 463 557 467 558
rect 462 556 468 557
rect 462 552 463 556
rect 467 552 468 556
rect 462 551 468 552
rect 480 540 482 602
rect 488 601 490 613
rect 494 607 500 608
rect 494 603 495 607
rect 499 603 500 607
rect 494 602 500 603
rect 526 607 532 608
rect 526 603 527 607
rect 531 603 532 607
rect 526 602 532 603
rect 486 600 492 601
rect 486 596 487 600
rect 491 596 492 600
rect 486 595 492 596
rect 496 588 498 602
rect 528 588 530 602
rect 536 601 538 613
rect 584 601 586 613
rect 610 611 611 615
rect 615 611 616 615
rect 631 613 635 614
rect 647 618 651 619
rect 647 613 651 614
rect 610 610 616 611
rect 534 600 540 601
rect 534 596 535 600
rect 539 596 540 600
rect 534 595 540 596
rect 582 600 588 601
rect 582 596 583 600
rect 587 596 588 600
rect 582 595 588 596
rect 612 588 614 610
rect 632 601 634 613
rect 630 600 636 601
rect 630 596 631 600
rect 635 596 636 600
rect 630 595 636 596
rect 656 588 658 630
rect 704 619 706 639
rect 752 636 754 650
rect 758 644 764 645
rect 758 640 759 644
rect 763 640 764 644
rect 758 639 764 640
rect 822 644 828 645
rect 822 640 823 644
rect 827 640 828 644
rect 822 639 828 640
rect 750 635 756 636
rect 750 631 751 635
rect 755 631 756 635
rect 750 630 756 631
rect 760 619 762 639
rect 824 619 826 639
rect 848 636 850 658
rect 1134 655 1140 656
rect 1094 652 1100 653
rect 1094 648 1095 652
rect 1099 648 1100 652
rect 1134 651 1135 655
rect 1139 651 1140 655
rect 1134 650 1140 651
rect 1246 652 1252 653
rect 1094 647 1100 648
rect 1136 647 1138 650
rect 1246 648 1247 652
rect 1251 648 1252 652
rect 1246 647 1252 648
rect 1286 652 1292 653
rect 1286 648 1287 652
rect 1291 648 1292 652
rect 1286 647 1292 648
rect 846 635 852 636
rect 846 631 847 635
rect 851 631 852 635
rect 846 630 852 631
rect 1096 619 1098 647
rect 1135 646 1139 647
rect 1135 641 1139 642
rect 1159 646 1163 647
rect 1159 641 1163 642
rect 1199 646 1203 647
rect 1199 641 1203 642
rect 1239 646 1243 647
rect 1239 641 1243 642
rect 1247 646 1251 647
rect 1247 641 1251 642
rect 1279 646 1283 647
rect 1279 641 1283 642
rect 1287 646 1291 647
rect 1287 641 1291 642
rect 1136 638 1138 641
rect 1158 640 1164 641
rect 1134 637 1140 638
rect 1134 633 1135 637
rect 1139 633 1140 637
rect 1158 636 1159 640
rect 1163 636 1164 640
rect 1158 635 1164 636
rect 1198 640 1204 641
rect 1198 636 1199 640
rect 1203 636 1204 640
rect 1198 635 1204 636
rect 1238 640 1244 641
rect 1238 636 1239 640
rect 1243 636 1244 640
rect 1238 635 1244 636
rect 1278 640 1284 641
rect 1278 636 1279 640
rect 1283 636 1284 640
rect 1278 635 1284 636
rect 1134 632 1140 633
rect 1182 623 1188 624
rect 1134 620 1140 621
rect 679 618 683 619
rect 679 613 683 614
rect 703 618 707 619
rect 703 613 707 614
rect 727 618 731 619
rect 727 613 731 614
rect 759 618 763 619
rect 759 613 763 614
rect 823 618 827 619
rect 823 613 827 614
rect 1095 618 1099 619
rect 1134 616 1135 620
rect 1139 616 1140 620
rect 1182 619 1183 623
rect 1187 619 1188 623
rect 1182 618 1188 619
rect 1206 623 1212 624
rect 1206 619 1207 623
rect 1211 619 1212 623
rect 1206 618 1212 619
rect 1246 623 1252 624
rect 1246 619 1247 623
rect 1251 619 1252 623
rect 1246 618 1252 619
rect 1286 623 1292 624
rect 1286 619 1287 623
rect 1291 619 1292 623
rect 1286 618 1292 619
rect 1134 615 1140 616
rect 1095 613 1099 614
rect 680 601 682 613
rect 686 607 692 608
rect 686 603 687 607
rect 691 603 692 607
rect 686 602 692 603
rect 678 600 684 601
rect 678 596 679 600
rect 683 596 684 600
rect 678 595 684 596
rect 688 588 690 602
rect 728 601 730 613
rect 742 607 748 608
rect 742 603 743 607
rect 747 603 748 607
rect 742 602 748 603
rect 726 600 732 601
rect 726 596 727 600
rect 731 596 732 600
rect 726 595 732 596
rect 744 588 746 602
rect 1096 593 1098 613
rect 1094 592 1100 593
rect 1094 588 1095 592
rect 1099 588 1100 592
rect 1136 591 1138 615
rect 1158 612 1164 613
rect 1158 608 1159 612
rect 1163 608 1164 612
rect 1158 607 1164 608
rect 1160 591 1162 607
rect 494 587 500 588
rect 494 583 495 587
rect 499 583 500 587
rect 494 582 500 583
rect 526 587 532 588
rect 526 583 527 587
rect 531 583 532 587
rect 526 582 532 583
rect 610 587 616 588
rect 610 583 611 587
rect 615 583 616 587
rect 610 582 616 583
rect 654 587 660 588
rect 654 583 655 587
rect 659 583 660 587
rect 654 582 660 583
rect 686 587 692 588
rect 686 583 687 587
rect 691 583 692 587
rect 686 582 692 583
rect 742 587 748 588
rect 1094 587 1100 588
rect 1135 590 1139 591
rect 742 583 743 587
rect 747 583 748 587
rect 1135 585 1139 586
rect 1159 590 1163 591
rect 1159 585 1163 586
rect 742 582 748 583
rect 1094 575 1100 576
rect 486 572 492 573
rect 486 568 487 572
rect 491 568 492 572
rect 486 567 492 568
rect 534 572 540 573
rect 534 568 535 572
rect 539 568 540 572
rect 534 567 540 568
rect 582 572 588 573
rect 582 568 583 572
rect 587 568 588 572
rect 582 567 588 568
rect 630 572 636 573
rect 630 568 631 572
rect 635 568 636 572
rect 630 567 636 568
rect 678 572 684 573
rect 678 568 679 572
rect 683 568 684 572
rect 678 567 684 568
rect 726 572 732 573
rect 726 568 727 572
rect 731 568 732 572
rect 1094 571 1095 575
rect 1099 571 1100 575
rect 1094 570 1100 571
rect 726 567 732 568
rect 488 563 490 567
rect 536 563 538 567
rect 584 563 586 567
rect 632 563 634 567
rect 680 563 682 567
rect 728 563 730 567
rect 1096 563 1098 570
rect 1136 565 1138 585
rect 1160 573 1162 585
rect 1184 580 1186 618
rect 1198 612 1204 613
rect 1198 608 1199 612
rect 1203 608 1204 612
rect 1198 607 1204 608
rect 1200 591 1202 607
rect 1208 604 1210 618
rect 1238 612 1244 613
rect 1238 608 1239 612
rect 1243 608 1244 612
rect 1238 607 1244 608
rect 1206 603 1212 604
rect 1206 599 1207 603
rect 1211 599 1212 603
rect 1206 598 1212 599
rect 1240 591 1242 607
rect 1248 604 1250 618
rect 1278 612 1284 613
rect 1278 608 1279 612
rect 1283 608 1284 612
rect 1278 607 1284 608
rect 1246 603 1252 604
rect 1246 599 1247 603
rect 1251 599 1252 603
rect 1246 598 1252 599
rect 1280 591 1282 607
rect 1288 604 1290 618
rect 1286 603 1292 604
rect 1286 599 1287 603
rect 1291 599 1292 603
rect 1286 598 1292 599
rect 1296 596 1298 662
rect 1334 652 1340 653
rect 1334 648 1335 652
rect 1339 648 1340 652
rect 1334 647 1340 648
rect 1390 652 1396 653
rect 1390 648 1391 652
rect 1395 648 1396 652
rect 1390 647 1396 648
rect 1446 652 1452 653
rect 1446 648 1447 652
rect 1451 648 1452 652
rect 1446 647 1452 648
rect 1510 652 1516 653
rect 1510 648 1511 652
rect 1515 648 1516 652
rect 1510 647 1516 648
rect 1582 652 1588 653
rect 1582 648 1583 652
rect 1587 648 1588 652
rect 1582 647 1588 648
rect 1654 652 1660 653
rect 1654 648 1655 652
rect 1659 648 1660 652
rect 1654 647 1660 648
rect 1335 646 1339 647
rect 1335 641 1339 642
rect 1343 646 1347 647
rect 1343 641 1347 642
rect 1391 646 1395 647
rect 1391 641 1395 642
rect 1415 646 1419 647
rect 1415 641 1419 642
rect 1447 646 1451 647
rect 1447 641 1451 642
rect 1495 646 1499 647
rect 1495 641 1499 642
rect 1511 646 1515 647
rect 1511 641 1515 642
rect 1583 646 1587 647
rect 1583 641 1587 642
rect 1655 646 1659 647
rect 1655 641 1659 642
rect 1342 640 1348 641
rect 1342 636 1343 640
rect 1347 636 1348 640
rect 1342 635 1348 636
rect 1414 640 1420 641
rect 1414 636 1415 640
rect 1419 636 1420 640
rect 1414 635 1420 636
rect 1494 640 1500 641
rect 1494 636 1495 640
rect 1499 636 1500 640
rect 1494 635 1500 636
rect 1582 640 1588 641
rect 1582 636 1583 640
rect 1587 636 1588 640
rect 1582 635 1588 636
rect 1518 623 1524 624
rect 1518 619 1519 623
rect 1523 619 1524 623
rect 1518 618 1524 619
rect 1342 612 1348 613
rect 1342 608 1343 612
rect 1347 608 1348 612
rect 1342 607 1348 608
rect 1414 612 1420 613
rect 1414 608 1415 612
rect 1419 608 1420 612
rect 1414 607 1420 608
rect 1494 612 1500 613
rect 1494 608 1495 612
rect 1499 608 1500 612
rect 1494 607 1500 608
rect 1294 595 1300 596
rect 1294 591 1295 595
rect 1299 591 1300 595
rect 1344 591 1346 607
rect 1416 591 1418 607
rect 1496 591 1498 607
rect 1199 590 1203 591
rect 1199 585 1203 586
rect 1239 590 1243 591
rect 1239 585 1243 586
rect 1279 590 1283 591
rect 1294 590 1300 591
rect 1319 590 1323 591
rect 1279 585 1283 586
rect 1319 585 1323 586
rect 1343 590 1347 591
rect 1343 585 1347 586
rect 1359 590 1363 591
rect 1359 585 1363 586
rect 1415 590 1419 591
rect 1415 585 1419 586
rect 1487 590 1491 591
rect 1487 585 1491 586
rect 1495 590 1499 591
rect 1520 588 1522 618
rect 1582 612 1588 613
rect 1582 608 1583 612
rect 1587 608 1588 612
rect 1582 607 1588 608
rect 1584 591 1586 607
rect 1664 596 1666 662
rect 1734 652 1740 653
rect 1734 648 1735 652
rect 1739 648 1740 652
rect 1734 647 1740 648
rect 1822 652 1828 653
rect 1822 648 1823 652
rect 1827 648 1828 652
rect 1822 647 1828 648
rect 1910 652 1916 653
rect 1910 648 1911 652
rect 1915 648 1916 652
rect 1910 647 1916 648
rect 1671 646 1675 647
rect 1671 641 1675 642
rect 1735 646 1739 647
rect 1735 641 1739 642
rect 1759 646 1763 647
rect 1759 641 1763 642
rect 1823 646 1827 647
rect 1823 641 1827 642
rect 1839 646 1843 647
rect 1839 641 1843 642
rect 1911 646 1915 647
rect 1911 641 1915 642
rect 1919 646 1923 647
rect 1919 641 1923 642
rect 1670 640 1676 641
rect 1670 636 1671 640
rect 1675 636 1676 640
rect 1670 635 1676 636
rect 1758 640 1764 641
rect 1758 636 1759 640
rect 1763 636 1764 640
rect 1758 635 1764 636
rect 1838 640 1844 641
rect 1838 636 1839 640
rect 1843 636 1844 640
rect 1838 635 1844 636
rect 1918 640 1924 641
rect 1918 636 1919 640
rect 1923 636 1924 640
rect 1918 635 1924 636
rect 1948 624 1950 690
rect 2000 681 2002 693
rect 2048 688 2050 722
rect 2070 716 2076 717
rect 2070 712 2071 716
rect 2075 712 2076 716
rect 2070 711 2076 712
rect 2072 699 2074 711
rect 2096 708 2098 770
rect 2118 763 2124 764
rect 2118 759 2119 763
rect 2123 759 2124 763
rect 2118 758 2124 759
rect 2120 751 2122 758
rect 2119 750 2123 751
rect 2119 745 2123 746
rect 2120 742 2122 745
rect 2118 741 2124 742
rect 2118 737 2119 741
rect 2123 737 2124 741
rect 2118 736 2124 737
rect 2118 724 2124 725
rect 2118 720 2119 724
rect 2123 720 2124 724
rect 2118 719 2124 720
rect 2094 707 2100 708
rect 2094 703 2095 707
rect 2099 703 2100 707
rect 2094 702 2100 703
rect 2120 699 2122 719
rect 2071 698 2075 699
rect 2071 693 2075 694
rect 2119 698 2123 699
rect 2119 693 2123 694
rect 2046 687 2052 688
rect 2046 683 2047 687
rect 2051 683 2052 687
rect 2046 682 2052 683
rect 2072 681 2074 693
rect 1998 680 2004 681
rect 1998 676 1999 680
rect 2003 676 2004 680
rect 1998 675 2004 676
rect 2070 680 2076 681
rect 2070 676 2071 680
rect 2075 676 2076 680
rect 2070 675 2076 676
rect 2120 673 2122 693
rect 2118 672 2124 673
rect 2118 668 2119 672
rect 2123 668 2124 672
rect 2094 667 2100 668
rect 2118 667 2124 668
rect 2094 663 2095 667
rect 2099 663 2100 667
rect 2094 662 2100 663
rect 1998 652 2004 653
rect 1998 648 1999 652
rect 2003 648 2004 652
rect 1998 647 2004 648
rect 2070 652 2076 653
rect 2070 648 2071 652
rect 2075 648 2076 652
rect 2070 647 2076 648
rect 1999 646 2003 647
rect 1999 641 2003 642
rect 2007 646 2011 647
rect 2007 641 2011 642
rect 2071 646 2075 647
rect 2071 641 2075 642
rect 2006 640 2012 641
rect 2006 636 2007 640
rect 2011 636 2012 640
rect 2006 635 2012 636
rect 2070 640 2076 641
rect 2070 636 2071 640
rect 2075 636 2076 640
rect 2070 635 2076 636
rect 1934 623 1940 624
rect 1934 619 1935 623
rect 1939 619 1940 623
rect 1934 618 1940 619
rect 1946 623 1952 624
rect 1946 619 1947 623
rect 1951 619 1952 623
rect 1946 618 1952 619
rect 2046 623 2052 624
rect 2046 619 2047 623
rect 2051 619 2052 623
rect 2046 618 2052 619
rect 2054 623 2060 624
rect 2054 619 2055 623
rect 2059 619 2060 623
rect 2054 618 2060 619
rect 1670 612 1676 613
rect 1670 608 1671 612
rect 1675 608 1676 612
rect 1670 607 1676 608
rect 1758 612 1764 613
rect 1758 608 1759 612
rect 1763 608 1764 612
rect 1758 607 1764 608
rect 1838 612 1844 613
rect 1838 608 1839 612
rect 1843 608 1844 612
rect 1838 607 1844 608
rect 1918 612 1924 613
rect 1918 608 1919 612
rect 1923 608 1924 612
rect 1918 607 1924 608
rect 1662 595 1668 596
rect 1662 591 1663 595
rect 1667 591 1668 595
rect 1672 591 1674 607
rect 1760 591 1762 607
rect 1840 591 1842 607
rect 1878 603 1884 604
rect 1878 599 1879 603
rect 1883 599 1884 603
rect 1878 598 1884 599
rect 1567 590 1571 591
rect 1495 585 1499 586
rect 1518 587 1524 588
rect 1182 579 1188 580
rect 1182 575 1183 579
rect 1187 575 1188 579
rect 1182 574 1188 575
rect 1200 573 1202 585
rect 1206 579 1212 580
rect 1206 575 1207 579
rect 1211 575 1212 579
rect 1206 574 1212 575
rect 1158 572 1164 573
rect 1158 568 1159 572
rect 1163 568 1164 572
rect 1158 567 1164 568
rect 1198 572 1204 573
rect 1198 568 1199 572
rect 1203 568 1204 572
rect 1198 567 1204 568
rect 1134 564 1140 565
rect 487 562 491 563
rect 487 557 491 558
rect 511 562 515 563
rect 511 557 515 558
rect 535 562 539 563
rect 535 557 539 558
rect 559 562 563 563
rect 559 557 563 558
rect 583 562 587 563
rect 583 557 587 558
rect 607 562 611 563
rect 607 557 611 558
rect 631 562 635 563
rect 631 557 635 558
rect 655 562 659 563
rect 655 557 659 558
rect 679 562 683 563
rect 679 557 683 558
rect 703 562 707 563
rect 703 557 707 558
rect 727 562 731 563
rect 727 557 731 558
rect 751 562 755 563
rect 751 557 755 558
rect 1095 562 1099 563
rect 1134 560 1135 564
rect 1139 560 1140 564
rect 1208 560 1210 574
rect 1240 573 1242 585
rect 1246 579 1252 580
rect 1246 575 1247 579
rect 1251 575 1252 579
rect 1246 574 1252 575
rect 1238 572 1244 573
rect 1238 568 1239 572
rect 1243 568 1244 572
rect 1238 567 1244 568
rect 1248 560 1250 574
rect 1280 573 1282 585
rect 1286 579 1292 580
rect 1286 575 1287 579
rect 1291 575 1292 579
rect 1286 574 1292 575
rect 1278 572 1284 573
rect 1278 568 1279 572
rect 1283 568 1284 572
rect 1278 567 1284 568
rect 1288 560 1290 574
rect 1320 573 1322 585
rect 1326 579 1332 580
rect 1326 575 1327 579
rect 1331 575 1332 579
rect 1326 574 1332 575
rect 1318 572 1324 573
rect 1318 568 1319 572
rect 1323 568 1324 572
rect 1318 567 1324 568
rect 1328 560 1330 574
rect 1360 573 1362 585
rect 1366 579 1372 580
rect 1366 575 1367 579
rect 1371 575 1372 579
rect 1366 574 1372 575
rect 1358 572 1364 573
rect 1358 568 1359 572
rect 1363 568 1364 572
rect 1358 567 1364 568
rect 1368 560 1370 574
rect 1416 573 1418 585
rect 1488 573 1490 585
rect 1518 583 1519 587
rect 1523 583 1524 587
rect 1567 585 1571 586
rect 1583 590 1587 591
rect 1583 585 1587 586
rect 1655 590 1659 591
rect 1662 590 1668 591
rect 1671 590 1675 591
rect 1655 585 1659 586
rect 1671 585 1675 586
rect 1751 590 1755 591
rect 1751 585 1755 586
rect 1759 590 1763 591
rect 1759 585 1763 586
rect 1839 590 1843 591
rect 1839 585 1843 586
rect 1855 590 1859 591
rect 1855 585 1859 586
rect 1518 582 1524 583
rect 1568 573 1570 585
rect 1656 573 1658 585
rect 1670 579 1676 580
rect 1670 575 1671 579
rect 1675 575 1676 579
rect 1670 574 1676 575
rect 1414 572 1420 573
rect 1414 568 1415 572
rect 1419 568 1420 572
rect 1414 567 1420 568
rect 1486 572 1492 573
rect 1486 568 1487 572
rect 1491 568 1492 572
rect 1486 567 1492 568
rect 1566 572 1572 573
rect 1566 568 1567 572
rect 1571 568 1572 572
rect 1566 567 1572 568
rect 1654 572 1660 573
rect 1654 568 1655 572
rect 1659 568 1660 572
rect 1654 567 1660 568
rect 1672 560 1674 574
rect 1752 573 1754 585
rect 1766 579 1772 580
rect 1766 575 1767 579
rect 1771 575 1772 579
rect 1766 574 1772 575
rect 1750 572 1756 573
rect 1750 568 1751 572
rect 1755 568 1756 572
rect 1750 567 1756 568
rect 1768 560 1770 574
rect 1856 573 1858 585
rect 1854 572 1860 573
rect 1854 568 1855 572
rect 1859 568 1860 572
rect 1854 567 1860 568
rect 1880 560 1882 598
rect 1920 591 1922 607
rect 1936 604 1938 618
rect 2006 612 2012 613
rect 2006 608 2007 612
rect 2011 608 2012 612
rect 2006 607 2012 608
rect 1934 603 1940 604
rect 1934 599 1935 603
rect 1939 599 1940 603
rect 1934 598 1940 599
rect 2008 591 2010 607
rect 1919 590 1923 591
rect 1919 585 1923 586
rect 1967 590 1971 591
rect 1967 585 1971 586
rect 2007 590 2011 591
rect 2007 585 2011 586
rect 1938 579 1944 580
rect 1938 575 1939 579
rect 1943 575 1944 579
rect 1938 574 1944 575
rect 1946 579 1952 580
rect 1946 575 1947 579
rect 1951 575 1952 579
rect 1946 574 1952 575
rect 1940 560 1942 574
rect 1134 559 1140 560
rect 1206 559 1212 560
rect 1095 557 1099 558
rect 510 556 516 557
rect 510 552 511 556
rect 515 552 516 556
rect 510 551 516 552
rect 558 556 564 557
rect 558 552 559 556
rect 563 552 564 556
rect 558 551 564 552
rect 606 556 612 557
rect 606 552 607 556
rect 611 552 612 556
rect 606 551 612 552
rect 654 556 660 557
rect 654 552 655 556
rect 659 552 660 556
rect 654 551 660 552
rect 702 556 708 557
rect 702 552 703 556
rect 707 552 708 556
rect 702 551 708 552
rect 750 556 756 557
rect 750 552 751 556
rect 755 552 756 556
rect 1096 554 1098 557
rect 1206 555 1207 559
rect 1211 555 1212 559
rect 1206 554 1212 555
rect 1246 559 1252 560
rect 1246 555 1247 559
rect 1251 555 1252 559
rect 1246 554 1252 555
rect 1286 559 1292 560
rect 1286 555 1287 559
rect 1291 555 1292 559
rect 1286 554 1292 555
rect 1326 559 1332 560
rect 1326 555 1327 559
rect 1331 555 1332 559
rect 1326 554 1332 555
rect 1366 559 1372 560
rect 1366 555 1367 559
rect 1371 555 1372 559
rect 1366 554 1372 555
rect 1430 559 1436 560
rect 1430 555 1431 559
rect 1435 555 1436 559
rect 1430 554 1436 555
rect 1534 559 1540 560
rect 1534 555 1535 559
rect 1539 555 1540 559
rect 1534 554 1540 555
rect 1670 559 1676 560
rect 1670 555 1671 559
rect 1675 555 1676 559
rect 1670 554 1676 555
rect 1766 559 1772 560
rect 1766 555 1767 559
rect 1771 555 1772 559
rect 1766 554 1772 555
rect 1878 559 1884 560
rect 1878 555 1879 559
rect 1883 555 1884 559
rect 1878 554 1884 555
rect 1938 559 1944 560
rect 1938 555 1939 559
rect 1943 555 1944 559
rect 1938 554 1944 555
rect 750 551 756 552
rect 1094 553 1100 554
rect 1094 549 1095 553
rect 1099 549 1100 553
rect 1094 548 1100 549
rect 1134 547 1140 548
rect 1134 543 1135 547
rect 1139 543 1140 547
rect 1134 542 1140 543
rect 1158 544 1164 545
rect 190 539 196 540
rect 190 535 191 539
rect 195 535 196 539
rect 190 534 196 535
rect 238 539 244 540
rect 238 535 239 539
rect 243 535 244 539
rect 238 534 244 535
rect 294 539 300 540
rect 294 535 295 539
rect 299 535 300 539
rect 294 534 300 535
rect 318 539 324 540
rect 318 535 319 539
rect 323 535 324 539
rect 318 534 324 535
rect 390 539 396 540
rect 390 535 391 539
rect 395 535 396 539
rect 390 534 396 535
rect 438 539 444 540
rect 438 535 439 539
rect 443 535 444 539
rect 438 534 444 535
rect 446 539 452 540
rect 446 535 447 539
rect 451 535 452 539
rect 446 534 452 535
rect 478 539 484 540
rect 478 535 479 539
rect 483 535 484 539
rect 478 534 484 535
rect 498 539 504 540
rect 498 535 499 539
rect 503 535 504 539
rect 498 534 504 535
rect 690 539 696 540
rect 690 535 691 539
rect 695 535 696 539
rect 690 534 696 535
rect 1094 536 1100 537
rect 174 528 180 529
rect 174 524 175 528
rect 179 524 180 528
rect 174 523 180 524
rect 158 519 164 520
rect 158 515 159 519
rect 163 515 164 519
rect 158 514 164 515
rect 176 503 178 523
rect 192 520 194 534
rect 222 528 228 529
rect 222 524 223 528
rect 227 524 228 528
rect 222 523 228 524
rect 190 519 196 520
rect 190 515 191 519
rect 195 515 196 519
rect 190 514 196 515
rect 224 503 226 523
rect 240 520 242 534
rect 278 528 284 529
rect 278 524 279 528
rect 283 524 284 528
rect 278 523 284 524
rect 238 519 244 520
rect 238 515 239 519
rect 243 515 244 519
rect 238 514 244 515
rect 280 503 282 523
rect 296 520 298 534
rect 294 519 300 520
rect 294 515 295 519
rect 299 515 300 519
rect 294 514 300 515
rect 111 502 115 503
rect 111 497 115 498
rect 135 502 139 503
rect 135 497 139 498
rect 175 502 179 503
rect 175 497 179 498
rect 223 502 227 503
rect 223 497 227 498
rect 231 502 235 503
rect 231 497 235 498
rect 279 502 283 503
rect 279 497 283 498
rect 295 502 299 503
rect 295 497 299 498
rect 112 477 114 497
rect 136 485 138 497
rect 176 485 178 497
rect 190 491 196 492
rect 190 487 191 491
rect 195 487 196 491
rect 190 486 196 487
rect 134 484 140 485
rect 134 480 135 484
rect 139 480 140 484
rect 134 479 140 480
rect 174 484 180 485
rect 174 480 175 484
rect 179 480 180 484
rect 174 479 180 480
rect 110 476 116 477
rect 110 472 111 476
rect 115 472 116 476
rect 192 472 194 486
rect 232 485 234 497
rect 246 491 252 492
rect 246 487 247 491
rect 251 487 252 491
rect 246 486 252 487
rect 286 491 292 492
rect 286 487 287 491
rect 291 487 292 491
rect 286 486 292 487
rect 230 484 236 485
rect 230 480 231 484
rect 235 480 236 484
rect 230 479 236 480
rect 248 472 250 486
rect 288 472 290 486
rect 296 485 298 497
rect 320 492 322 534
rect 326 528 332 529
rect 326 524 327 528
rect 331 524 332 528
rect 326 523 332 524
rect 374 528 380 529
rect 374 524 375 528
rect 379 524 380 528
rect 374 523 380 524
rect 328 503 330 523
rect 376 503 378 523
rect 392 520 394 534
rect 422 528 428 529
rect 422 524 423 528
rect 427 524 428 528
rect 422 523 428 524
rect 382 519 388 520
rect 382 515 383 519
rect 387 515 388 519
rect 382 514 388 515
rect 390 519 396 520
rect 390 515 391 519
rect 395 515 396 519
rect 390 514 396 515
rect 327 502 331 503
rect 327 497 331 498
rect 359 502 363 503
rect 359 497 363 498
rect 375 502 379 503
rect 375 497 379 498
rect 318 491 324 492
rect 318 487 319 491
rect 323 487 324 491
rect 318 486 324 487
rect 360 485 362 497
rect 294 484 300 485
rect 294 480 295 484
rect 299 480 300 484
rect 294 479 300 480
rect 358 484 364 485
rect 358 480 359 484
rect 363 480 364 484
rect 358 479 364 480
rect 384 472 386 514
rect 424 503 426 523
rect 440 520 442 534
rect 462 528 468 529
rect 462 524 463 528
rect 467 524 468 528
rect 462 523 468 524
rect 438 519 444 520
rect 438 515 439 519
rect 443 515 444 519
rect 438 514 444 515
rect 464 503 466 523
rect 500 520 502 534
rect 510 528 516 529
rect 510 524 511 528
rect 515 524 516 528
rect 510 523 516 524
rect 558 528 564 529
rect 558 524 559 528
rect 563 524 564 528
rect 558 523 564 524
rect 606 528 612 529
rect 606 524 607 528
rect 611 524 612 528
rect 606 523 612 524
rect 654 528 660 529
rect 654 524 655 528
rect 659 524 660 528
rect 654 523 660 524
rect 498 519 504 520
rect 498 515 499 519
rect 503 515 504 519
rect 498 514 504 515
rect 512 503 514 523
rect 560 503 562 523
rect 582 511 588 512
rect 582 507 583 511
rect 587 507 588 511
rect 582 506 588 507
rect 423 502 427 503
rect 423 497 427 498
rect 463 502 467 503
rect 463 497 467 498
rect 479 502 483 503
rect 479 497 483 498
rect 511 502 515 503
rect 511 497 515 498
rect 535 502 539 503
rect 535 497 539 498
rect 559 502 563 503
rect 559 497 563 498
rect 424 485 426 497
rect 438 491 444 492
rect 438 487 439 491
rect 443 487 444 491
rect 438 486 444 487
rect 422 484 428 485
rect 422 480 423 484
rect 427 480 428 484
rect 422 479 428 480
rect 440 472 442 486
rect 480 485 482 497
rect 494 491 500 492
rect 494 487 495 491
rect 499 487 500 491
rect 494 486 500 487
rect 478 484 484 485
rect 478 480 479 484
rect 483 480 484 484
rect 478 479 484 480
rect 496 472 498 486
rect 536 485 538 497
rect 550 491 556 492
rect 550 487 551 491
rect 555 487 556 491
rect 550 486 556 487
rect 534 484 540 485
rect 534 480 535 484
rect 539 480 540 484
rect 534 479 540 480
rect 110 471 116 472
rect 182 471 188 472
rect 182 467 183 471
rect 187 467 188 471
rect 182 466 188 467
rect 190 471 196 472
rect 190 467 191 471
rect 195 467 196 471
rect 190 466 196 467
rect 246 471 252 472
rect 246 467 247 471
rect 251 467 252 471
rect 246 466 252 467
rect 286 471 292 472
rect 286 467 287 471
rect 291 467 292 471
rect 286 466 292 467
rect 382 471 388 472
rect 382 467 383 471
rect 387 467 388 471
rect 382 466 388 467
rect 438 471 444 472
rect 438 467 439 471
rect 443 467 444 471
rect 438 466 444 467
rect 494 471 500 472
rect 494 467 495 471
rect 499 467 500 471
rect 494 466 500 467
rect 110 459 116 460
rect 110 455 111 459
rect 115 455 116 459
rect 110 454 116 455
rect 134 456 140 457
rect 112 447 114 454
rect 134 452 135 456
rect 139 452 140 456
rect 134 451 140 452
rect 174 456 180 457
rect 174 452 175 456
rect 179 452 180 456
rect 174 451 180 452
rect 136 447 138 451
rect 176 447 178 451
rect 111 446 115 447
rect 111 441 115 442
rect 135 446 139 447
rect 135 441 139 442
rect 175 446 179 447
rect 175 441 179 442
rect 112 438 114 441
rect 174 440 180 441
rect 110 437 116 438
rect 110 433 111 437
rect 115 433 116 437
rect 174 436 175 440
rect 179 436 180 440
rect 174 435 180 436
rect 110 432 116 433
rect 110 420 116 421
rect 110 416 111 420
rect 115 416 116 420
rect 110 415 116 416
rect 112 387 114 415
rect 174 412 180 413
rect 174 408 175 412
rect 179 408 180 412
rect 174 407 180 408
rect 176 387 178 407
rect 184 396 186 466
rect 230 456 236 457
rect 230 452 231 456
rect 235 452 236 456
rect 230 451 236 452
rect 294 456 300 457
rect 294 452 295 456
rect 299 452 300 456
rect 294 451 300 452
rect 358 456 364 457
rect 358 452 359 456
rect 363 452 364 456
rect 358 451 364 452
rect 422 456 428 457
rect 422 452 423 456
rect 427 452 428 456
rect 422 451 428 452
rect 478 456 484 457
rect 478 452 479 456
rect 483 452 484 456
rect 478 451 484 452
rect 534 456 540 457
rect 534 452 535 456
rect 539 452 540 456
rect 534 451 540 452
rect 232 447 234 451
rect 296 447 298 451
rect 360 447 362 451
rect 424 447 426 451
rect 480 447 482 451
rect 536 447 538 451
rect 215 446 219 447
rect 215 441 219 442
rect 231 446 235 447
rect 231 441 235 442
rect 263 446 267 447
rect 263 441 267 442
rect 295 446 299 447
rect 295 441 299 442
rect 327 446 331 447
rect 327 441 331 442
rect 359 446 363 447
rect 359 441 363 442
rect 391 446 395 447
rect 391 441 395 442
rect 423 446 427 447
rect 423 441 427 442
rect 463 446 467 447
rect 463 441 467 442
rect 479 446 483 447
rect 479 441 483 442
rect 535 446 539 447
rect 535 441 539 442
rect 214 440 220 441
rect 214 436 215 440
rect 219 436 220 440
rect 214 435 220 436
rect 262 440 268 441
rect 262 436 263 440
rect 267 436 268 440
rect 262 435 268 436
rect 326 440 332 441
rect 326 436 327 440
rect 331 436 332 440
rect 326 435 332 436
rect 390 440 396 441
rect 390 436 391 440
rect 395 436 396 440
rect 390 435 396 436
rect 462 440 468 441
rect 462 436 463 440
rect 467 436 468 440
rect 462 435 468 436
rect 534 440 540 441
rect 534 436 535 440
rect 539 436 540 440
rect 534 435 540 436
rect 552 435 554 486
rect 584 476 586 506
rect 608 503 610 523
rect 656 503 658 523
rect 692 520 694 534
rect 1094 532 1095 536
rect 1099 532 1100 536
rect 1136 535 1138 542
rect 1158 540 1159 544
rect 1163 540 1164 544
rect 1158 539 1164 540
rect 1198 544 1204 545
rect 1198 540 1199 544
rect 1203 540 1204 544
rect 1198 539 1204 540
rect 1238 544 1244 545
rect 1238 540 1239 544
rect 1243 540 1244 544
rect 1238 539 1244 540
rect 1278 544 1284 545
rect 1278 540 1279 544
rect 1283 540 1284 544
rect 1278 539 1284 540
rect 1318 544 1324 545
rect 1318 540 1319 544
rect 1323 540 1324 544
rect 1318 539 1324 540
rect 1358 544 1364 545
rect 1358 540 1359 544
rect 1363 540 1364 544
rect 1358 539 1364 540
rect 1414 544 1420 545
rect 1414 540 1415 544
rect 1419 540 1420 544
rect 1414 539 1420 540
rect 1160 535 1162 539
rect 1200 535 1202 539
rect 1240 535 1242 539
rect 1280 535 1282 539
rect 1320 535 1322 539
rect 1360 535 1362 539
rect 1416 535 1418 539
rect 1094 531 1100 532
rect 1135 534 1139 535
rect 702 528 708 529
rect 702 524 703 528
rect 707 524 708 528
rect 702 523 708 524
rect 750 528 756 529
rect 750 524 751 528
rect 755 524 756 528
rect 750 523 756 524
rect 690 519 696 520
rect 690 515 691 519
rect 695 515 696 519
rect 690 514 696 515
rect 704 503 706 523
rect 752 503 754 523
rect 1096 503 1098 531
rect 1135 529 1139 530
rect 1159 534 1163 535
rect 1159 529 1163 530
rect 1199 534 1203 535
rect 1199 529 1203 530
rect 1239 534 1243 535
rect 1239 529 1243 530
rect 1279 534 1283 535
rect 1279 529 1283 530
rect 1303 534 1307 535
rect 1303 529 1307 530
rect 1319 534 1323 535
rect 1319 529 1323 530
rect 1343 534 1347 535
rect 1343 529 1347 530
rect 1359 534 1363 535
rect 1359 529 1363 530
rect 1383 534 1387 535
rect 1383 529 1387 530
rect 1415 534 1419 535
rect 1415 529 1419 530
rect 1423 534 1427 535
rect 1423 529 1427 530
rect 1136 526 1138 529
rect 1302 528 1308 529
rect 1134 525 1140 526
rect 1134 521 1135 525
rect 1139 521 1140 525
rect 1302 524 1303 528
rect 1307 524 1308 528
rect 1302 523 1308 524
rect 1342 528 1348 529
rect 1342 524 1343 528
rect 1347 524 1348 528
rect 1342 523 1348 524
rect 1382 528 1388 529
rect 1382 524 1383 528
rect 1387 524 1388 528
rect 1382 523 1388 524
rect 1422 528 1428 529
rect 1422 524 1423 528
rect 1427 524 1428 528
rect 1422 523 1428 524
rect 1134 520 1140 521
rect 1350 511 1356 512
rect 1134 508 1140 509
rect 1134 504 1135 508
rect 1139 504 1140 508
rect 1350 507 1351 511
rect 1355 507 1356 511
rect 1350 506 1356 507
rect 1390 511 1396 512
rect 1390 507 1391 511
rect 1395 507 1396 511
rect 1390 506 1396 507
rect 1134 503 1140 504
rect 591 502 595 503
rect 591 497 595 498
rect 607 502 611 503
rect 607 497 611 498
rect 639 502 643 503
rect 639 497 643 498
rect 655 502 659 503
rect 655 497 659 498
rect 687 502 691 503
rect 687 497 691 498
rect 703 502 707 503
rect 703 497 707 498
rect 735 502 739 503
rect 735 497 739 498
rect 751 502 755 503
rect 751 497 755 498
rect 791 502 795 503
rect 791 497 795 498
rect 847 502 851 503
rect 847 497 851 498
rect 1095 502 1099 503
rect 1095 497 1099 498
rect 592 485 594 497
rect 598 491 604 492
rect 598 487 599 491
rect 603 487 604 491
rect 598 486 604 487
rect 590 484 596 485
rect 590 480 591 484
rect 595 480 596 484
rect 590 479 596 480
rect 582 475 588 476
rect 582 471 583 475
rect 587 471 588 475
rect 600 472 602 486
rect 640 485 642 497
rect 654 491 660 492
rect 654 487 655 491
rect 659 487 660 491
rect 654 486 660 487
rect 638 484 644 485
rect 638 480 639 484
rect 643 480 644 484
rect 638 479 644 480
rect 656 472 658 486
rect 688 485 690 497
rect 702 491 708 492
rect 702 487 703 491
rect 707 487 708 491
rect 702 486 708 487
rect 686 484 692 485
rect 686 480 687 484
rect 691 480 692 484
rect 686 479 692 480
rect 704 472 706 486
rect 736 485 738 497
rect 750 491 756 492
rect 750 487 751 491
rect 755 487 756 491
rect 750 486 756 487
rect 734 484 740 485
rect 734 480 735 484
rect 739 480 740 484
rect 734 479 740 480
rect 752 472 754 486
rect 792 485 794 497
rect 806 491 812 492
rect 806 487 807 491
rect 811 487 812 491
rect 806 486 812 487
rect 790 484 796 485
rect 790 480 791 484
rect 795 480 796 484
rect 790 479 796 480
rect 808 472 810 486
rect 848 485 850 497
rect 854 491 860 492
rect 854 487 855 491
rect 859 487 860 491
rect 854 486 860 487
rect 862 491 868 492
rect 862 487 863 491
rect 867 487 868 491
rect 862 486 868 487
rect 846 484 852 485
rect 846 480 847 484
rect 851 480 852 484
rect 846 479 852 480
rect 856 472 858 486
rect 582 470 588 471
rect 598 471 604 472
rect 598 467 599 471
rect 603 467 604 471
rect 598 466 604 467
rect 654 471 660 472
rect 654 467 655 471
rect 659 467 660 471
rect 654 466 660 467
rect 702 471 708 472
rect 702 467 703 471
rect 707 467 708 471
rect 702 466 708 467
rect 750 471 756 472
rect 750 467 751 471
rect 755 467 756 471
rect 750 466 756 467
rect 806 471 812 472
rect 806 467 807 471
rect 811 467 812 471
rect 806 466 812 467
rect 854 471 860 472
rect 854 467 855 471
rect 859 467 860 471
rect 854 466 860 467
rect 590 456 596 457
rect 590 452 591 456
rect 595 452 596 456
rect 590 451 596 452
rect 638 456 644 457
rect 638 452 639 456
rect 643 452 644 456
rect 638 451 644 452
rect 686 456 692 457
rect 686 452 687 456
rect 691 452 692 456
rect 686 451 692 452
rect 734 456 740 457
rect 734 452 735 456
rect 739 452 740 456
rect 734 451 740 452
rect 790 456 796 457
rect 790 452 791 456
rect 795 452 796 456
rect 790 451 796 452
rect 846 456 852 457
rect 846 452 847 456
rect 851 452 852 456
rect 846 451 852 452
rect 592 447 594 451
rect 640 447 642 451
rect 688 447 690 451
rect 736 447 738 451
rect 792 447 794 451
rect 848 447 850 451
rect 591 446 595 447
rect 591 441 595 442
rect 607 446 611 447
rect 607 441 611 442
rect 639 446 643 447
rect 639 441 643 442
rect 679 446 683 447
rect 679 441 683 442
rect 687 446 691 447
rect 687 441 691 442
rect 735 446 739 447
rect 735 441 739 442
rect 743 446 747 447
rect 743 441 747 442
rect 791 446 795 447
rect 791 441 795 442
rect 807 446 811 447
rect 807 441 811 442
rect 847 446 851 447
rect 847 441 851 442
rect 606 440 612 441
rect 606 436 607 440
rect 611 436 612 440
rect 606 435 612 436
rect 678 440 684 441
rect 678 436 679 440
rect 683 436 684 440
rect 678 435 684 436
rect 742 440 748 441
rect 742 436 743 440
rect 747 436 748 440
rect 742 435 748 436
rect 806 440 812 441
rect 806 436 807 440
rect 811 436 812 440
rect 806 435 812 436
rect 552 433 562 435
rect 560 424 562 433
rect 864 432 866 486
rect 1096 477 1098 497
rect 1136 483 1138 503
rect 1302 500 1308 501
rect 1302 496 1303 500
rect 1307 496 1308 500
rect 1302 495 1308 496
rect 1342 500 1348 501
rect 1342 496 1343 500
rect 1347 496 1348 500
rect 1342 495 1348 496
rect 1304 483 1306 495
rect 1344 483 1346 495
rect 1352 492 1354 506
rect 1382 500 1388 501
rect 1382 496 1383 500
rect 1387 496 1388 500
rect 1382 495 1388 496
rect 1350 491 1356 492
rect 1350 487 1351 491
rect 1355 487 1356 491
rect 1350 486 1356 487
rect 1384 483 1386 495
rect 1392 492 1394 506
rect 1422 500 1428 501
rect 1422 496 1423 500
rect 1427 496 1428 500
rect 1422 495 1428 496
rect 1390 491 1396 492
rect 1390 487 1391 491
rect 1395 487 1396 491
rect 1390 486 1396 487
rect 1424 483 1426 495
rect 1432 492 1434 554
rect 1486 544 1492 545
rect 1486 540 1487 544
rect 1491 540 1492 544
rect 1486 539 1492 540
rect 1488 535 1490 539
rect 1463 534 1467 535
rect 1463 529 1467 530
rect 1487 534 1491 535
rect 1487 529 1491 530
rect 1503 534 1507 535
rect 1503 529 1507 530
rect 1462 528 1468 529
rect 1462 524 1463 528
rect 1467 524 1468 528
rect 1462 523 1468 524
rect 1502 528 1508 529
rect 1502 524 1503 528
rect 1507 524 1508 528
rect 1502 523 1508 524
rect 1446 519 1452 520
rect 1446 515 1447 519
rect 1451 515 1452 519
rect 1446 514 1452 515
rect 1448 492 1450 514
rect 1478 511 1484 512
rect 1478 507 1479 511
rect 1483 507 1484 511
rect 1478 506 1484 507
rect 1518 511 1524 512
rect 1518 507 1519 511
rect 1523 507 1524 511
rect 1518 506 1524 507
rect 1462 500 1468 501
rect 1462 496 1463 500
rect 1467 496 1468 500
rect 1462 495 1468 496
rect 1430 491 1436 492
rect 1430 487 1431 491
rect 1435 487 1436 491
rect 1430 486 1436 487
rect 1446 491 1452 492
rect 1446 487 1447 491
rect 1451 487 1452 491
rect 1446 486 1452 487
rect 1464 483 1466 495
rect 1480 492 1482 506
rect 1502 500 1508 501
rect 1502 496 1503 500
rect 1507 496 1508 500
rect 1502 495 1508 496
rect 1478 491 1484 492
rect 1478 487 1479 491
rect 1483 487 1484 491
rect 1478 486 1484 487
rect 1504 483 1506 495
rect 1520 492 1522 506
rect 1518 491 1524 492
rect 1518 487 1519 491
rect 1523 487 1524 491
rect 1518 486 1524 487
rect 1536 484 1538 554
rect 1566 544 1572 545
rect 1566 540 1567 544
rect 1571 540 1572 544
rect 1566 539 1572 540
rect 1654 544 1660 545
rect 1654 540 1655 544
rect 1659 540 1660 544
rect 1654 539 1660 540
rect 1750 544 1756 545
rect 1750 540 1751 544
rect 1755 540 1756 544
rect 1750 539 1756 540
rect 1854 544 1860 545
rect 1854 540 1855 544
rect 1859 540 1860 544
rect 1854 539 1860 540
rect 1568 535 1570 539
rect 1656 535 1658 539
rect 1752 535 1754 539
rect 1856 535 1858 539
rect 1543 534 1547 535
rect 1543 529 1547 530
rect 1567 534 1571 535
rect 1567 529 1571 530
rect 1591 534 1595 535
rect 1591 529 1595 530
rect 1647 534 1651 535
rect 1647 529 1651 530
rect 1655 534 1659 535
rect 1655 529 1659 530
rect 1703 534 1707 535
rect 1703 529 1707 530
rect 1751 534 1755 535
rect 1751 529 1755 530
rect 1767 534 1771 535
rect 1767 529 1771 530
rect 1839 534 1843 535
rect 1839 529 1843 530
rect 1855 534 1859 535
rect 1855 529 1859 530
rect 1919 534 1923 535
rect 1919 529 1923 530
rect 1542 528 1548 529
rect 1542 524 1543 528
rect 1547 524 1548 528
rect 1542 523 1548 524
rect 1590 528 1596 529
rect 1590 524 1591 528
rect 1595 524 1596 528
rect 1590 523 1596 524
rect 1646 528 1652 529
rect 1646 524 1647 528
rect 1651 524 1652 528
rect 1646 523 1652 524
rect 1702 528 1708 529
rect 1702 524 1703 528
rect 1707 524 1708 528
rect 1702 523 1708 524
rect 1766 528 1772 529
rect 1766 524 1767 528
rect 1771 524 1772 528
rect 1766 523 1772 524
rect 1838 528 1844 529
rect 1838 524 1839 528
rect 1843 524 1844 528
rect 1838 523 1844 524
rect 1918 528 1924 529
rect 1918 524 1919 528
rect 1923 524 1924 528
rect 1918 523 1924 524
rect 1948 512 1950 574
rect 1968 573 1970 585
rect 2048 580 2050 618
rect 2056 604 2058 618
rect 2070 612 2076 613
rect 2070 608 2071 612
rect 2075 608 2076 612
rect 2070 607 2076 608
rect 2054 603 2060 604
rect 2054 599 2055 603
rect 2059 599 2060 603
rect 2054 598 2060 599
rect 2072 591 2074 607
rect 2096 604 2098 662
rect 2118 655 2124 656
rect 2118 651 2119 655
rect 2123 651 2124 655
rect 2118 650 2124 651
rect 2120 647 2122 650
rect 2119 646 2123 647
rect 2119 641 2123 642
rect 2120 638 2122 641
rect 2118 637 2124 638
rect 2118 633 2119 637
rect 2123 633 2124 637
rect 2118 632 2124 633
rect 2118 620 2124 621
rect 2118 616 2119 620
rect 2123 616 2124 620
rect 2118 615 2124 616
rect 2094 603 2100 604
rect 2094 599 2095 603
rect 2099 599 2100 603
rect 2094 598 2100 599
rect 2120 591 2122 615
rect 2071 590 2075 591
rect 2071 585 2075 586
rect 2119 590 2123 591
rect 2119 585 2123 586
rect 2046 579 2052 580
rect 2046 575 2047 579
rect 2051 575 2052 579
rect 2046 574 2052 575
rect 2072 573 2074 585
rect 1966 572 1972 573
rect 1966 568 1967 572
rect 1971 568 1972 572
rect 1966 567 1972 568
rect 2070 572 2076 573
rect 2070 568 2071 572
rect 2075 568 2076 572
rect 2070 567 2076 568
rect 2120 565 2122 585
rect 2118 564 2124 565
rect 2118 560 2119 564
rect 2123 560 2124 564
rect 2118 559 2124 560
rect 2118 547 2124 548
rect 1966 544 1972 545
rect 1966 540 1967 544
rect 1971 540 1972 544
rect 1966 539 1972 540
rect 2070 544 2076 545
rect 2070 540 2071 544
rect 2075 540 2076 544
rect 2118 543 2119 547
rect 2123 543 2124 547
rect 2118 542 2124 543
rect 2070 539 2076 540
rect 1968 535 1970 539
rect 2072 535 2074 539
rect 2120 535 2122 542
rect 1967 534 1971 535
rect 1967 529 1971 530
rect 2007 534 2011 535
rect 2007 529 2011 530
rect 2071 534 2075 535
rect 2071 529 2075 530
rect 2119 534 2123 535
rect 2119 529 2123 530
rect 2006 528 2012 529
rect 2006 524 2007 528
rect 2011 524 2012 528
rect 2006 523 2012 524
rect 2070 528 2076 529
rect 2070 524 2071 528
rect 2075 524 2076 528
rect 2120 526 2122 529
rect 2070 523 2076 524
rect 2118 525 2124 526
rect 2118 521 2119 525
rect 2123 521 2124 525
rect 2118 520 2124 521
rect 1554 511 1560 512
rect 1554 507 1555 511
rect 1559 507 1560 511
rect 1554 506 1560 507
rect 1662 511 1668 512
rect 1662 507 1663 511
rect 1667 507 1668 511
rect 1662 506 1668 507
rect 1718 511 1724 512
rect 1718 507 1719 511
rect 1723 507 1724 511
rect 1718 506 1724 507
rect 1782 511 1788 512
rect 1782 507 1783 511
rect 1787 507 1788 511
rect 1782 506 1788 507
rect 1846 511 1852 512
rect 1846 507 1847 511
rect 1851 507 1852 511
rect 1846 506 1852 507
rect 1910 511 1916 512
rect 1910 507 1911 511
rect 1915 507 1916 511
rect 1910 506 1916 507
rect 1946 511 1952 512
rect 1946 507 1947 511
rect 1951 507 1952 511
rect 1946 506 1952 507
rect 2078 511 2084 512
rect 2078 507 2079 511
rect 2083 507 2084 511
rect 2078 506 2084 507
rect 2094 511 2100 512
rect 2094 507 2095 511
rect 2099 507 2100 511
rect 2094 506 2100 507
rect 2118 508 2124 509
rect 1542 500 1548 501
rect 1542 496 1543 500
rect 1547 496 1548 500
rect 1542 495 1548 496
rect 1534 483 1540 484
rect 1544 483 1546 495
rect 1135 482 1139 483
rect 1135 477 1139 478
rect 1295 482 1299 483
rect 1295 477 1299 478
rect 1303 482 1307 483
rect 1303 477 1307 478
rect 1335 482 1339 483
rect 1335 477 1339 478
rect 1343 482 1347 483
rect 1343 477 1347 478
rect 1375 482 1379 483
rect 1375 477 1379 478
rect 1383 482 1387 483
rect 1383 477 1387 478
rect 1423 482 1427 483
rect 1423 477 1427 478
rect 1463 482 1467 483
rect 1463 477 1467 478
rect 1471 482 1475 483
rect 1471 477 1475 478
rect 1503 482 1507 483
rect 1503 477 1507 478
rect 1527 482 1531 483
rect 1534 479 1535 483
rect 1539 479 1540 483
rect 1534 478 1540 479
rect 1543 482 1547 483
rect 1527 477 1531 478
rect 1543 477 1547 478
rect 1094 476 1100 477
rect 1094 472 1095 476
rect 1099 472 1100 476
rect 1094 471 1100 472
rect 1094 459 1100 460
rect 1094 455 1095 459
rect 1099 455 1100 459
rect 1136 457 1138 477
rect 1296 465 1298 477
rect 1336 465 1338 477
rect 1350 471 1356 472
rect 1350 467 1351 471
rect 1355 467 1356 471
rect 1350 466 1356 467
rect 1294 464 1300 465
rect 1294 460 1295 464
rect 1299 460 1300 464
rect 1294 459 1300 460
rect 1334 464 1340 465
rect 1334 460 1335 464
rect 1339 460 1340 464
rect 1334 459 1340 460
rect 1094 454 1100 455
rect 1134 456 1140 457
rect 1096 447 1098 454
rect 1134 452 1135 456
rect 1139 452 1140 456
rect 1352 452 1354 466
rect 1376 465 1378 477
rect 1390 471 1396 472
rect 1390 467 1391 471
rect 1395 467 1396 471
rect 1390 466 1396 467
rect 1374 464 1380 465
rect 1374 460 1375 464
rect 1379 460 1380 464
rect 1374 459 1380 460
rect 1392 452 1394 466
rect 1424 465 1426 477
rect 1438 471 1444 472
rect 1438 467 1439 471
rect 1443 467 1444 471
rect 1438 466 1444 467
rect 1422 464 1428 465
rect 1422 460 1423 464
rect 1427 460 1428 464
rect 1422 459 1428 460
rect 1440 452 1442 466
rect 1472 465 1474 477
rect 1486 471 1492 472
rect 1486 467 1487 471
rect 1491 467 1492 471
rect 1486 466 1492 467
rect 1470 464 1476 465
rect 1470 460 1471 464
rect 1475 460 1476 464
rect 1470 459 1476 460
rect 1488 452 1490 466
rect 1528 465 1530 477
rect 1556 472 1558 506
rect 1590 500 1596 501
rect 1590 496 1591 500
rect 1595 496 1596 500
rect 1590 495 1596 496
rect 1646 500 1652 501
rect 1646 496 1647 500
rect 1651 496 1652 500
rect 1646 495 1652 496
rect 1592 483 1594 495
rect 1648 483 1650 495
rect 1664 492 1666 506
rect 1702 500 1708 501
rect 1702 496 1703 500
rect 1707 496 1708 500
rect 1702 495 1708 496
rect 1662 491 1668 492
rect 1662 487 1663 491
rect 1667 487 1668 491
rect 1662 486 1668 487
rect 1704 483 1706 495
rect 1720 492 1722 506
rect 1766 500 1772 501
rect 1766 496 1767 500
rect 1771 496 1772 500
rect 1766 495 1772 496
rect 1718 491 1724 492
rect 1718 487 1719 491
rect 1723 487 1724 491
rect 1718 486 1724 487
rect 1768 483 1770 495
rect 1784 492 1786 506
rect 1838 500 1844 501
rect 1838 496 1839 500
rect 1843 496 1844 500
rect 1838 495 1844 496
rect 1782 491 1788 492
rect 1782 487 1783 491
rect 1787 487 1788 491
rect 1782 486 1788 487
rect 1840 483 1842 495
rect 1848 492 1850 506
rect 1846 491 1852 492
rect 1846 487 1847 491
rect 1851 487 1852 491
rect 1846 486 1852 487
rect 1583 482 1587 483
rect 1583 477 1587 478
rect 1591 482 1595 483
rect 1591 477 1595 478
rect 1647 482 1651 483
rect 1647 477 1651 478
rect 1703 482 1707 483
rect 1703 477 1707 478
rect 1719 482 1723 483
rect 1719 477 1723 478
rect 1767 482 1771 483
rect 1767 477 1771 478
rect 1807 482 1811 483
rect 1807 477 1811 478
rect 1839 482 1843 483
rect 1839 477 1843 478
rect 1895 482 1899 483
rect 1895 477 1899 478
rect 1542 471 1548 472
rect 1542 467 1543 471
rect 1547 467 1548 471
rect 1542 466 1548 467
rect 1554 471 1560 472
rect 1554 467 1555 471
rect 1559 467 1560 471
rect 1554 466 1560 467
rect 1526 464 1532 465
rect 1526 460 1527 464
rect 1531 460 1532 464
rect 1526 459 1532 460
rect 1544 452 1546 466
rect 1584 465 1586 477
rect 1648 465 1650 477
rect 1662 471 1668 472
rect 1662 467 1663 471
rect 1667 467 1668 471
rect 1662 466 1668 467
rect 1582 464 1588 465
rect 1582 460 1583 464
rect 1587 460 1588 464
rect 1582 459 1588 460
rect 1646 464 1652 465
rect 1646 460 1647 464
rect 1651 460 1652 464
rect 1646 459 1652 460
rect 1664 452 1666 466
rect 1720 465 1722 477
rect 1734 471 1740 472
rect 1734 467 1735 471
rect 1739 467 1740 471
rect 1734 466 1740 467
rect 1718 464 1724 465
rect 1718 460 1719 464
rect 1723 460 1724 464
rect 1718 459 1724 460
rect 1736 452 1738 466
rect 1808 465 1810 477
rect 1822 471 1828 472
rect 1822 467 1823 471
rect 1827 467 1828 471
rect 1822 466 1828 467
rect 1806 464 1812 465
rect 1806 460 1807 464
rect 1811 460 1812 464
rect 1806 459 1812 460
rect 1824 452 1826 466
rect 1896 465 1898 477
rect 1912 472 1914 506
rect 1918 500 1924 501
rect 1918 496 1919 500
rect 1923 496 1924 500
rect 1918 495 1924 496
rect 2006 500 2012 501
rect 2006 496 2007 500
rect 2011 496 2012 500
rect 2006 495 2012 496
rect 2070 500 2076 501
rect 2070 496 2071 500
rect 2075 496 2076 500
rect 2070 495 2076 496
rect 1920 483 1922 495
rect 1998 491 2004 492
rect 1998 487 1999 491
rect 2003 487 2004 491
rect 1998 486 2004 487
rect 1919 482 1923 483
rect 1919 477 1923 478
rect 1991 482 1995 483
rect 1991 477 1995 478
rect 1902 471 1908 472
rect 1902 467 1903 471
rect 1907 467 1908 471
rect 1902 466 1908 467
rect 1910 471 1916 472
rect 1910 467 1911 471
rect 1915 467 1916 471
rect 1910 466 1916 467
rect 1894 464 1900 465
rect 1894 460 1895 464
rect 1899 460 1900 464
rect 1894 459 1900 460
rect 1904 452 1906 466
rect 1992 465 1994 477
rect 1990 464 1996 465
rect 1990 460 1991 464
rect 1995 460 1996 464
rect 1990 459 1996 460
rect 2000 452 2002 486
rect 2008 483 2010 495
rect 2072 483 2074 495
rect 2080 492 2082 506
rect 2078 491 2084 492
rect 2078 487 2079 491
rect 2083 487 2084 491
rect 2078 486 2084 487
rect 2007 482 2011 483
rect 2007 477 2011 478
rect 2071 482 2075 483
rect 2071 477 2075 478
rect 2018 471 2024 472
rect 2018 467 2019 471
rect 2023 467 2024 471
rect 2018 466 2024 467
rect 1134 451 1140 452
rect 1342 451 1348 452
rect 1342 447 1343 451
rect 1347 447 1348 451
rect 871 446 875 447
rect 871 441 875 442
rect 943 446 947 447
rect 943 441 947 442
rect 1095 446 1099 447
rect 1342 446 1348 447
rect 1350 451 1356 452
rect 1350 447 1351 451
rect 1355 447 1356 451
rect 1350 446 1356 447
rect 1390 451 1396 452
rect 1390 447 1391 451
rect 1395 447 1396 451
rect 1390 446 1396 447
rect 1438 451 1444 452
rect 1438 447 1439 451
rect 1443 447 1444 451
rect 1438 446 1444 447
rect 1486 451 1492 452
rect 1486 447 1487 451
rect 1491 447 1492 451
rect 1486 446 1492 447
rect 1542 451 1548 452
rect 1542 447 1543 451
rect 1547 447 1548 451
rect 1542 446 1548 447
rect 1610 451 1616 452
rect 1610 447 1611 451
rect 1615 447 1616 451
rect 1610 446 1616 447
rect 1662 451 1668 452
rect 1662 447 1663 451
rect 1667 447 1668 451
rect 1662 446 1668 447
rect 1734 451 1740 452
rect 1734 447 1735 451
rect 1739 447 1740 451
rect 1734 446 1740 447
rect 1822 451 1828 452
rect 1822 447 1823 451
rect 1827 447 1828 451
rect 1822 446 1828 447
rect 1902 451 1908 452
rect 1902 447 1903 451
rect 1907 447 1908 451
rect 1902 446 1908 447
rect 1998 451 2004 452
rect 1998 447 1999 451
rect 2003 447 2004 451
rect 1998 446 2004 447
rect 1095 441 1099 442
rect 870 440 876 441
rect 870 436 871 440
rect 875 436 876 440
rect 870 435 876 436
rect 942 440 948 441
rect 942 436 943 440
rect 947 436 948 440
rect 1096 438 1098 441
rect 1134 439 1140 440
rect 942 435 948 436
rect 1094 437 1100 438
rect 1094 433 1095 437
rect 1099 433 1100 437
rect 1134 435 1135 439
rect 1139 435 1140 439
rect 1134 434 1140 435
rect 1294 436 1300 437
rect 1094 432 1100 433
rect 862 431 868 432
rect 1136 431 1138 434
rect 1294 432 1295 436
rect 1299 432 1300 436
rect 1294 431 1300 432
rect 1334 436 1340 437
rect 1334 432 1335 436
rect 1339 432 1340 436
rect 1334 431 1340 432
rect 862 427 863 431
rect 867 427 868 431
rect 862 426 868 427
rect 1135 430 1139 431
rect 1135 425 1139 426
rect 1159 430 1163 431
rect 1159 425 1163 426
rect 1199 430 1203 431
rect 1199 425 1203 426
rect 1255 430 1259 431
rect 1255 425 1259 426
rect 1295 430 1299 431
rect 1295 425 1299 426
rect 1335 430 1339 431
rect 1335 425 1339 426
rect 198 423 204 424
rect 198 419 199 423
rect 203 419 204 423
rect 198 418 204 419
rect 222 423 228 424
rect 222 419 223 423
rect 227 419 228 423
rect 222 418 228 419
rect 250 423 256 424
rect 250 419 251 423
rect 255 419 256 423
rect 250 418 256 419
rect 350 423 356 424
rect 350 419 351 423
rect 355 419 356 423
rect 350 418 356 419
rect 550 423 556 424
rect 550 419 551 423
rect 555 419 556 423
rect 550 418 556 419
rect 558 423 564 424
rect 558 419 559 423
rect 563 419 564 423
rect 1136 422 1138 425
rect 1158 424 1164 425
rect 1134 421 1140 422
rect 558 418 564 419
rect 1094 420 1100 421
rect 182 395 188 396
rect 182 391 183 395
rect 187 391 188 395
rect 182 390 188 391
rect 111 386 115 387
rect 111 381 115 382
rect 175 386 179 387
rect 175 381 179 382
rect 112 361 114 381
rect 176 369 178 381
rect 200 376 202 418
rect 214 412 220 413
rect 214 408 215 412
rect 219 408 220 412
rect 214 407 220 408
rect 216 387 218 407
rect 224 404 226 418
rect 252 404 254 418
rect 262 412 268 413
rect 262 408 263 412
rect 267 408 268 412
rect 262 407 268 408
rect 326 412 332 413
rect 326 408 327 412
rect 331 408 332 412
rect 326 407 332 408
rect 222 403 228 404
rect 222 399 223 403
rect 227 399 228 403
rect 222 398 228 399
rect 250 403 256 404
rect 250 399 251 403
rect 255 399 256 403
rect 250 398 256 399
rect 264 387 266 407
rect 328 387 330 407
rect 352 396 354 418
rect 390 412 396 413
rect 390 408 391 412
rect 395 408 396 412
rect 390 407 396 408
rect 462 412 468 413
rect 462 408 463 412
rect 467 408 468 412
rect 462 407 468 408
rect 534 412 540 413
rect 534 408 535 412
rect 539 408 540 412
rect 534 407 540 408
rect 350 395 356 396
rect 350 391 351 395
rect 355 391 356 395
rect 350 390 356 391
rect 392 387 394 407
rect 430 403 436 404
rect 430 399 431 403
rect 435 399 436 403
rect 430 398 436 399
rect 215 386 219 387
rect 215 381 219 382
rect 263 386 267 387
rect 263 381 267 382
rect 271 386 275 387
rect 271 381 275 382
rect 327 386 331 387
rect 327 381 331 382
rect 335 386 339 387
rect 391 386 395 387
rect 335 381 339 382
rect 362 383 368 384
rect 198 375 204 376
rect 198 371 199 375
rect 203 371 204 375
rect 198 370 204 371
rect 216 369 218 381
rect 222 375 228 376
rect 222 371 223 375
rect 227 371 228 375
rect 222 370 228 371
rect 174 368 180 369
rect 174 364 175 368
rect 179 364 180 368
rect 174 363 180 364
rect 214 368 220 369
rect 214 364 215 368
rect 219 364 220 368
rect 214 363 220 364
rect 110 360 116 361
rect 110 356 111 360
rect 115 356 116 360
rect 224 356 226 370
rect 272 369 274 381
rect 336 369 338 381
rect 362 379 363 383
rect 367 379 368 383
rect 391 381 395 382
rect 407 386 411 387
rect 407 381 411 382
rect 362 378 368 379
rect 270 368 276 369
rect 270 364 271 368
rect 275 364 276 368
rect 270 363 276 364
rect 334 368 340 369
rect 334 364 335 368
rect 339 364 340 368
rect 334 363 340 364
rect 364 356 366 378
rect 408 369 410 381
rect 406 368 412 369
rect 406 364 407 368
rect 411 364 412 368
rect 406 363 412 364
rect 432 356 434 398
rect 464 387 466 407
rect 536 387 538 407
rect 552 404 554 418
rect 1094 416 1095 420
rect 1099 416 1100 420
rect 1134 417 1135 421
rect 1139 417 1140 421
rect 1158 420 1159 424
rect 1163 420 1164 424
rect 1158 419 1164 420
rect 1198 424 1204 425
rect 1198 420 1199 424
rect 1203 420 1204 424
rect 1198 419 1204 420
rect 1254 424 1260 425
rect 1254 420 1255 424
rect 1259 420 1260 424
rect 1254 419 1260 420
rect 1334 424 1340 425
rect 1334 420 1335 424
rect 1339 420 1340 424
rect 1334 419 1340 420
rect 1134 416 1140 417
rect 1094 415 1100 416
rect 606 412 612 413
rect 606 408 607 412
rect 611 408 612 412
rect 606 407 612 408
rect 678 412 684 413
rect 678 408 679 412
rect 683 408 684 412
rect 678 407 684 408
rect 742 412 748 413
rect 742 408 743 412
rect 747 408 748 412
rect 742 407 748 408
rect 806 412 812 413
rect 806 408 807 412
rect 811 408 812 412
rect 806 407 812 408
rect 870 412 876 413
rect 870 408 871 412
rect 875 408 876 412
rect 870 407 876 408
rect 942 412 948 413
rect 942 408 943 412
rect 947 408 948 412
rect 942 407 948 408
rect 550 403 556 404
rect 550 399 551 403
rect 555 399 556 403
rect 550 398 556 399
rect 608 387 610 407
rect 680 387 682 407
rect 744 387 746 407
rect 808 387 810 407
rect 872 387 874 407
rect 914 403 920 404
rect 914 399 915 403
rect 919 399 920 403
rect 914 398 920 399
rect 463 386 467 387
rect 463 381 467 382
rect 487 386 491 387
rect 487 381 491 382
rect 535 386 539 387
rect 535 381 539 382
rect 567 386 571 387
rect 567 381 571 382
rect 607 386 611 387
rect 607 381 611 382
rect 639 386 643 387
rect 639 381 643 382
rect 679 386 683 387
rect 679 381 683 382
rect 711 386 715 387
rect 711 381 715 382
rect 743 386 747 387
rect 743 381 747 382
rect 775 386 779 387
rect 775 381 779 382
rect 807 386 811 387
rect 807 381 811 382
rect 839 386 843 387
rect 839 381 843 382
rect 871 386 875 387
rect 871 381 875 382
rect 895 386 899 387
rect 895 381 899 382
rect 488 369 490 381
rect 502 375 508 376
rect 502 371 503 375
rect 507 371 508 375
rect 502 370 508 371
rect 486 368 492 369
rect 486 364 487 368
rect 491 364 492 368
rect 486 363 492 364
rect 504 356 506 370
rect 568 369 570 381
rect 582 375 588 376
rect 582 371 583 375
rect 587 371 588 375
rect 582 370 588 371
rect 566 368 572 369
rect 566 364 567 368
rect 571 364 572 368
rect 566 363 572 364
rect 584 356 586 370
rect 640 369 642 381
rect 712 369 714 381
rect 726 375 732 376
rect 726 371 727 375
rect 731 371 732 375
rect 726 370 732 371
rect 638 368 644 369
rect 638 364 639 368
rect 643 364 644 368
rect 710 368 716 369
rect 638 363 644 364
rect 667 364 671 365
rect 710 364 711 368
rect 715 364 716 368
rect 710 363 716 364
rect 667 359 671 360
rect 668 356 670 359
rect 728 356 730 370
rect 776 369 778 381
rect 790 375 796 376
rect 790 371 791 375
rect 795 371 796 375
rect 790 370 796 371
rect 774 368 780 369
rect 774 364 775 368
rect 779 364 780 368
rect 774 363 780 364
rect 792 356 794 370
rect 840 369 842 381
rect 854 375 860 376
rect 854 371 855 375
rect 859 371 860 375
rect 854 370 860 371
rect 886 375 892 376
rect 886 371 887 375
rect 891 371 892 375
rect 886 370 892 371
rect 838 368 844 369
rect 838 364 839 368
rect 843 364 844 368
rect 838 363 844 364
rect 856 356 858 370
rect 888 356 890 370
rect 896 369 898 381
rect 894 368 900 369
rect 894 364 895 368
rect 899 364 900 368
rect 916 365 918 398
rect 944 387 946 407
rect 1096 387 1098 415
rect 1206 407 1212 408
rect 1134 404 1140 405
rect 1134 400 1135 404
rect 1139 400 1140 404
rect 1206 403 1207 407
rect 1211 403 1212 407
rect 1206 402 1212 403
rect 1134 399 1140 400
rect 943 386 947 387
rect 943 381 947 382
rect 951 386 955 387
rect 951 381 955 382
rect 1007 386 1011 387
rect 1007 381 1011 382
rect 1047 386 1051 387
rect 1047 381 1051 382
rect 1095 386 1099 387
rect 1095 381 1099 382
rect 952 369 954 381
rect 966 375 972 376
rect 966 371 967 375
rect 971 371 972 375
rect 966 370 972 371
rect 950 368 956 369
rect 894 363 900 364
rect 915 364 919 365
rect 950 364 951 368
rect 955 364 956 368
rect 950 363 956 364
rect 915 359 919 360
rect 968 356 970 370
rect 1008 369 1010 381
rect 1022 375 1028 376
rect 1022 371 1023 375
rect 1027 371 1028 375
rect 1022 370 1028 371
rect 1030 375 1036 376
rect 1030 371 1031 375
rect 1035 371 1036 375
rect 1030 370 1036 371
rect 1006 368 1012 369
rect 1006 364 1007 368
rect 1011 364 1012 368
rect 1006 363 1012 364
rect 1024 356 1026 370
rect 110 355 116 356
rect 222 355 228 356
rect 222 351 223 355
rect 227 351 228 355
rect 222 350 228 351
rect 362 355 368 356
rect 362 351 363 355
rect 367 351 368 355
rect 362 350 368 351
rect 430 355 436 356
rect 430 351 431 355
rect 435 351 436 355
rect 430 350 436 351
rect 502 355 508 356
rect 502 351 503 355
rect 507 351 508 355
rect 502 350 508 351
rect 582 355 588 356
rect 582 351 583 355
rect 587 351 588 355
rect 582 350 588 351
rect 666 355 672 356
rect 666 351 667 355
rect 671 351 672 355
rect 666 350 672 351
rect 726 355 732 356
rect 726 351 727 355
rect 731 351 732 355
rect 726 350 732 351
rect 790 355 796 356
rect 790 351 791 355
rect 795 351 796 355
rect 790 350 796 351
rect 854 355 860 356
rect 854 351 855 355
rect 859 351 860 355
rect 854 350 860 351
rect 886 355 892 356
rect 886 351 887 355
rect 891 351 892 355
rect 886 350 892 351
rect 966 355 972 356
rect 966 351 967 355
rect 971 351 972 355
rect 966 350 972 351
rect 1022 355 1028 356
rect 1022 351 1023 355
rect 1027 351 1028 355
rect 1022 350 1028 351
rect 110 343 116 344
rect 110 339 111 343
rect 115 339 116 343
rect 110 338 116 339
rect 174 340 180 341
rect 112 331 114 338
rect 174 336 175 340
rect 179 336 180 340
rect 174 335 180 336
rect 214 340 220 341
rect 214 336 215 340
rect 219 336 220 340
rect 214 335 220 336
rect 270 340 276 341
rect 270 336 271 340
rect 275 336 276 340
rect 270 335 276 336
rect 334 340 340 341
rect 334 336 335 340
rect 339 336 340 340
rect 334 335 340 336
rect 406 340 412 341
rect 406 336 407 340
rect 411 336 412 340
rect 406 335 412 336
rect 486 340 492 341
rect 486 336 487 340
rect 491 336 492 340
rect 486 335 492 336
rect 566 340 572 341
rect 566 336 567 340
rect 571 336 572 340
rect 566 335 572 336
rect 638 340 644 341
rect 638 336 639 340
rect 643 336 644 340
rect 638 335 644 336
rect 710 340 716 341
rect 710 336 711 340
rect 715 336 716 340
rect 710 335 716 336
rect 774 340 780 341
rect 774 336 775 340
rect 779 336 780 340
rect 774 335 780 336
rect 838 340 844 341
rect 838 336 839 340
rect 843 336 844 340
rect 838 335 844 336
rect 894 340 900 341
rect 894 336 895 340
rect 899 336 900 340
rect 894 335 900 336
rect 950 340 956 341
rect 950 336 951 340
rect 955 336 956 340
rect 950 335 956 336
rect 1006 340 1012 341
rect 1006 336 1007 340
rect 1011 336 1012 340
rect 1006 335 1012 336
rect 176 331 178 335
rect 216 331 218 335
rect 272 331 274 335
rect 336 331 338 335
rect 408 331 410 335
rect 488 331 490 335
rect 568 331 570 335
rect 640 331 642 335
rect 712 331 714 335
rect 776 331 778 335
rect 840 331 842 335
rect 896 331 898 335
rect 952 331 954 335
rect 1008 331 1010 335
rect 111 330 115 331
rect 111 325 115 326
rect 175 330 179 331
rect 175 325 179 326
rect 215 330 219 331
rect 215 325 219 326
rect 271 330 275 331
rect 271 325 275 326
rect 335 330 339 331
rect 335 325 339 326
rect 383 330 387 331
rect 383 325 387 326
rect 407 330 411 331
rect 407 325 411 326
rect 423 330 427 331
rect 423 325 427 326
rect 463 330 467 331
rect 463 325 467 326
rect 487 330 491 331
rect 487 325 491 326
rect 503 330 507 331
rect 503 325 507 326
rect 543 330 547 331
rect 543 325 547 326
rect 567 330 571 331
rect 567 325 571 326
rect 591 330 595 331
rect 591 325 595 326
rect 639 330 643 331
rect 639 325 643 326
rect 687 330 691 331
rect 687 325 691 326
rect 711 330 715 331
rect 711 325 715 326
rect 735 330 739 331
rect 735 325 739 326
rect 775 330 779 331
rect 775 325 779 326
rect 783 330 787 331
rect 783 325 787 326
rect 831 330 835 331
rect 831 325 835 326
rect 839 330 843 331
rect 839 325 843 326
rect 879 330 883 331
rect 879 325 883 326
rect 895 330 899 331
rect 895 325 899 326
rect 927 330 931 331
rect 927 325 931 326
rect 951 330 955 331
rect 951 325 955 326
rect 967 330 971 331
rect 967 325 971 326
rect 1007 330 1011 331
rect 1007 325 1011 326
rect 112 322 114 325
rect 382 324 388 325
rect 110 321 116 322
rect 110 317 111 321
rect 115 317 116 321
rect 382 320 383 324
rect 387 320 388 324
rect 382 319 388 320
rect 422 324 428 325
rect 422 320 423 324
rect 427 320 428 324
rect 422 319 428 320
rect 462 324 468 325
rect 462 320 463 324
rect 467 320 468 324
rect 462 319 468 320
rect 502 324 508 325
rect 502 320 503 324
rect 507 320 508 324
rect 502 319 508 320
rect 542 324 548 325
rect 542 320 543 324
rect 547 320 548 324
rect 542 319 548 320
rect 590 324 596 325
rect 590 320 591 324
rect 595 320 596 324
rect 590 319 596 320
rect 638 324 644 325
rect 638 320 639 324
rect 643 320 644 324
rect 638 319 644 320
rect 686 324 692 325
rect 686 320 687 324
rect 691 320 692 324
rect 686 319 692 320
rect 734 324 740 325
rect 734 320 735 324
rect 739 320 740 324
rect 734 319 740 320
rect 782 324 788 325
rect 782 320 783 324
rect 787 320 788 324
rect 782 319 788 320
rect 830 324 836 325
rect 830 320 831 324
rect 835 320 836 324
rect 830 319 836 320
rect 878 324 884 325
rect 878 320 879 324
rect 883 320 884 324
rect 878 319 884 320
rect 926 324 932 325
rect 926 320 927 324
rect 931 320 932 324
rect 926 319 932 320
rect 966 324 972 325
rect 966 320 967 324
rect 971 320 972 324
rect 966 319 972 320
rect 1006 324 1012 325
rect 1006 320 1007 324
rect 1011 320 1012 324
rect 1006 319 1012 320
rect 110 316 116 317
rect 1032 316 1034 370
rect 1048 369 1050 381
rect 1046 368 1052 369
rect 1046 364 1047 368
rect 1051 364 1052 368
rect 1046 363 1052 364
rect 1096 361 1098 381
rect 1136 375 1138 399
rect 1158 396 1164 397
rect 1158 392 1159 396
rect 1163 392 1164 396
rect 1158 391 1164 392
rect 1198 396 1204 397
rect 1198 392 1199 396
rect 1203 392 1204 396
rect 1198 391 1204 392
rect 1160 375 1162 391
rect 1182 375 1188 376
rect 1200 375 1202 391
rect 1208 388 1210 402
rect 1254 396 1260 397
rect 1254 392 1255 396
rect 1259 392 1260 396
rect 1254 391 1260 392
rect 1334 396 1340 397
rect 1334 392 1335 396
rect 1339 392 1340 396
rect 1334 391 1340 392
rect 1206 387 1212 388
rect 1206 383 1207 387
rect 1211 383 1212 387
rect 1206 382 1212 383
rect 1256 375 1258 391
rect 1336 375 1338 391
rect 1344 380 1346 446
rect 1374 436 1380 437
rect 1374 432 1375 436
rect 1379 432 1380 436
rect 1374 431 1380 432
rect 1422 436 1428 437
rect 1422 432 1423 436
rect 1427 432 1428 436
rect 1422 431 1428 432
rect 1470 436 1476 437
rect 1470 432 1471 436
rect 1475 432 1476 436
rect 1470 431 1476 432
rect 1526 436 1532 437
rect 1526 432 1527 436
rect 1531 432 1532 436
rect 1526 431 1532 432
rect 1582 436 1588 437
rect 1582 432 1583 436
rect 1587 432 1588 436
rect 1582 431 1588 432
rect 1375 430 1379 431
rect 1375 425 1379 426
rect 1415 430 1419 431
rect 1415 425 1419 426
rect 1423 430 1427 431
rect 1423 425 1427 426
rect 1471 430 1475 431
rect 1471 425 1475 426
rect 1503 430 1507 431
rect 1503 425 1507 426
rect 1527 430 1531 431
rect 1527 425 1531 426
rect 1583 430 1587 431
rect 1583 425 1587 426
rect 1591 430 1595 431
rect 1591 425 1595 426
rect 1414 424 1420 425
rect 1414 420 1415 424
rect 1419 420 1420 424
rect 1414 419 1420 420
rect 1502 424 1508 425
rect 1502 420 1503 424
rect 1507 420 1508 424
rect 1502 419 1508 420
rect 1590 424 1596 425
rect 1590 420 1591 424
rect 1595 420 1596 424
rect 1590 419 1596 420
rect 1486 415 1492 416
rect 1486 411 1487 415
rect 1491 411 1492 415
rect 1486 410 1492 411
rect 1414 396 1420 397
rect 1414 392 1415 396
rect 1419 392 1420 396
rect 1414 391 1420 392
rect 1342 379 1348 380
rect 1342 375 1343 379
rect 1347 375 1348 379
rect 1416 375 1418 391
rect 1135 374 1139 375
rect 1135 369 1139 370
rect 1159 374 1163 375
rect 1182 371 1183 375
rect 1187 371 1188 375
rect 1182 370 1188 371
rect 1199 374 1203 375
rect 1159 369 1163 370
rect 1094 360 1100 361
rect 1094 356 1095 360
rect 1099 356 1100 360
rect 1070 355 1076 356
rect 1094 355 1100 356
rect 1070 351 1071 355
rect 1075 351 1076 355
rect 1070 350 1076 351
rect 1046 340 1052 341
rect 1046 336 1047 340
rect 1051 336 1052 340
rect 1046 335 1052 336
rect 1048 331 1050 335
rect 1047 330 1051 331
rect 1047 325 1051 326
rect 1046 324 1052 325
rect 1046 320 1047 324
rect 1051 320 1052 324
rect 1046 319 1052 320
rect 1030 315 1036 316
rect 1030 311 1031 315
rect 1035 311 1036 315
rect 1030 310 1036 311
rect 406 307 412 308
rect 110 304 116 305
rect 110 300 111 304
rect 115 300 116 304
rect 406 303 407 307
rect 411 303 412 307
rect 406 302 412 303
rect 430 307 436 308
rect 430 303 431 307
rect 435 303 436 307
rect 430 302 436 303
rect 470 307 476 308
rect 470 303 471 307
rect 475 303 476 307
rect 470 302 476 303
rect 510 307 516 308
rect 510 303 511 307
rect 515 303 516 307
rect 510 302 516 303
rect 550 307 556 308
rect 550 303 551 307
rect 555 303 556 307
rect 550 302 556 303
rect 762 307 768 308
rect 762 303 763 307
rect 767 303 768 307
rect 762 302 768 303
rect 770 307 776 308
rect 770 303 771 307
rect 775 303 776 307
rect 770 302 776 303
rect 974 307 980 308
rect 974 303 975 307
rect 979 303 980 307
rect 974 302 980 303
rect 1014 307 1020 308
rect 1014 303 1015 307
rect 1019 303 1020 307
rect 1014 302 1020 303
rect 1054 307 1060 308
rect 1054 303 1055 307
rect 1059 303 1060 307
rect 1054 302 1060 303
rect 110 299 116 300
rect 112 271 114 299
rect 382 296 388 297
rect 382 292 383 296
rect 387 292 388 296
rect 382 291 388 292
rect 384 271 386 291
rect 111 270 115 271
rect 111 265 115 266
rect 287 270 291 271
rect 287 265 291 266
rect 327 270 331 271
rect 327 265 331 266
rect 367 270 371 271
rect 367 265 371 266
rect 383 270 387 271
rect 408 268 410 302
rect 422 296 428 297
rect 422 292 423 296
rect 427 292 428 296
rect 422 291 428 292
rect 424 271 426 291
rect 432 288 434 302
rect 462 296 468 297
rect 462 292 463 296
rect 467 292 468 296
rect 462 291 468 292
rect 430 287 436 288
rect 430 283 431 287
rect 435 283 436 287
rect 430 282 436 283
rect 464 271 466 291
rect 472 288 474 302
rect 502 296 508 297
rect 502 292 503 296
rect 507 292 508 296
rect 502 291 508 292
rect 470 287 476 288
rect 470 283 471 287
rect 475 283 476 287
rect 470 282 476 283
rect 504 271 506 291
rect 512 288 514 302
rect 542 296 548 297
rect 542 292 543 296
rect 547 292 548 296
rect 542 291 548 292
rect 510 287 516 288
rect 510 283 511 287
rect 515 283 516 287
rect 510 282 516 283
rect 544 271 546 291
rect 552 288 554 302
rect 590 296 596 297
rect 590 292 591 296
rect 595 292 596 296
rect 590 291 596 292
rect 638 296 644 297
rect 638 292 639 296
rect 643 292 644 296
rect 638 291 644 292
rect 686 296 692 297
rect 686 292 687 296
rect 691 292 692 296
rect 686 291 692 292
rect 734 296 740 297
rect 734 292 735 296
rect 739 292 740 296
rect 734 291 740 292
rect 550 287 556 288
rect 550 283 551 287
rect 555 283 556 287
rect 550 282 556 283
rect 592 271 594 291
rect 640 271 642 291
rect 688 271 690 291
rect 706 287 712 288
rect 706 283 707 287
rect 711 283 712 287
rect 706 282 712 283
rect 415 270 419 271
rect 383 265 387 266
rect 406 267 412 268
rect 112 245 114 265
rect 288 253 290 265
rect 328 253 330 265
rect 342 259 348 260
rect 342 255 343 259
rect 347 255 348 259
rect 342 254 348 255
rect 286 252 292 253
rect 286 248 287 252
rect 291 248 292 252
rect 286 247 292 248
rect 326 252 332 253
rect 326 248 327 252
rect 331 248 332 252
rect 326 247 332 248
rect 110 244 116 245
rect 110 240 111 244
rect 115 240 116 244
rect 344 240 346 254
rect 368 253 370 265
rect 406 263 407 267
rect 411 263 412 267
rect 415 265 419 266
rect 423 270 427 271
rect 423 265 427 266
rect 463 270 467 271
rect 463 265 467 266
rect 471 270 475 271
rect 471 265 475 266
rect 503 270 507 271
rect 503 265 507 266
rect 535 270 539 271
rect 535 265 539 266
rect 543 270 547 271
rect 543 265 547 266
rect 591 270 595 271
rect 591 265 595 266
rect 607 270 611 271
rect 607 265 611 266
rect 639 270 643 271
rect 639 265 643 266
rect 679 270 683 271
rect 679 265 683 266
rect 687 270 691 271
rect 687 265 691 266
rect 406 262 412 263
rect 374 259 380 260
rect 374 255 375 259
rect 379 255 380 259
rect 374 254 380 255
rect 366 252 372 253
rect 366 248 367 252
rect 371 248 372 252
rect 366 247 372 248
rect 376 240 378 254
rect 416 253 418 265
rect 430 259 436 260
rect 430 255 431 259
rect 435 255 436 259
rect 430 254 436 255
rect 414 252 420 253
rect 414 248 415 252
rect 419 248 420 252
rect 414 247 420 248
rect 432 240 434 254
rect 472 253 474 265
rect 486 259 492 260
rect 486 255 487 259
rect 491 255 492 259
rect 486 254 492 255
rect 470 252 476 253
rect 470 248 471 252
rect 475 248 476 252
rect 470 247 476 248
rect 488 240 490 254
rect 536 253 538 265
rect 550 259 556 260
rect 550 255 551 259
rect 555 255 556 259
rect 550 254 556 255
rect 534 252 540 253
rect 534 248 535 252
rect 539 248 540 252
rect 534 247 540 248
rect 552 240 554 254
rect 608 253 610 265
rect 622 259 628 260
rect 622 255 623 259
rect 627 255 628 259
rect 622 254 628 255
rect 606 252 612 253
rect 606 248 607 252
rect 611 248 612 252
rect 606 247 612 248
rect 624 240 626 254
rect 680 253 682 265
rect 698 259 704 260
rect 698 255 699 259
rect 703 255 704 259
rect 698 254 704 255
rect 678 252 684 253
rect 678 248 679 252
rect 683 248 684 252
rect 678 247 684 248
rect 110 239 116 240
rect 334 239 340 240
rect 334 235 335 239
rect 339 235 340 239
rect 334 234 340 235
rect 342 239 348 240
rect 342 235 343 239
rect 347 235 348 239
rect 342 234 348 235
rect 374 239 380 240
rect 374 235 375 239
rect 379 235 380 239
rect 374 234 380 235
rect 430 239 436 240
rect 430 235 431 239
rect 435 235 436 239
rect 430 234 436 235
rect 486 239 492 240
rect 486 235 487 239
rect 491 235 492 239
rect 486 234 492 235
rect 550 239 556 240
rect 550 235 551 239
rect 555 235 556 239
rect 550 234 556 235
rect 622 239 628 240
rect 622 235 623 239
rect 627 235 628 239
rect 622 234 628 235
rect 110 227 116 228
rect 110 223 111 227
rect 115 223 116 227
rect 110 222 116 223
rect 286 224 292 225
rect 112 207 114 222
rect 286 220 287 224
rect 291 220 292 224
rect 286 219 292 220
rect 326 224 332 225
rect 326 220 327 224
rect 331 220 332 224
rect 326 219 332 220
rect 288 207 290 219
rect 328 207 330 219
rect 111 206 115 207
rect 111 201 115 202
rect 167 206 171 207
rect 167 201 171 202
rect 207 206 211 207
rect 207 201 211 202
rect 247 206 251 207
rect 247 201 251 202
rect 287 206 291 207
rect 287 201 291 202
rect 295 206 299 207
rect 295 201 299 202
rect 327 206 331 207
rect 327 201 331 202
rect 112 198 114 201
rect 166 200 172 201
rect 110 197 116 198
rect 110 193 111 197
rect 115 193 116 197
rect 166 196 167 200
rect 171 196 172 200
rect 166 195 172 196
rect 206 200 212 201
rect 206 196 207 200
rect 211 196 212 200
rect 206 195 212 196
rect 246 200 252 201
rect 246 196 247 200
rect 251 196 252 200
rect 246 195 252 196
rect 294 200 300 201
rect 294 196 295 200
rect 299 196 300 200
rect 294 195 300 196
rect 110 192 116 193
rect 194 183 200 184
rect 110 180 116 181
rect 110 176 111 180
rect 115 176 116 180
rect 194 179 195 183
rect 199 179 200 183
rect 194 178 200 179
rect 214 183 220 184
rect 214 179 215 183
rect 219 179 220 183
rect 214 178 220 179
rect 254 183 260 184
rect 254 179 255 183
rect 259 179 260 183
rect 254 178 260 179
rect 110 175 116 176
rect 112 139 114 175
rect 166 172 172 173
rect 166 168 167 172
rect 171 168 172 172
rect 166 167 172 168
rect 168 139 170 167
rect 111 138 115 139
rect 111 133 115 134
rect 135 138 139 139
rect 135 133 139 134
rect 167 138 171 139
rect 167 133 171 134
rect 175 138 179 139
rect 196 136 198 178
rect 206 172 212 173
rect 206 168 207 172
rect 211 168 212 172
rect 206 167 212 168
rect 208 139 210 167
rect 216 164 218 178
rect 246 172 252 173
rect 246 168 247 172
rect 251 168 252 172
rect 246 167 252 168
rect 214 163 220 164
rect 214 159 215 163
rect 219 159 220 163
rect 214 158 220 159
rect 248 139 250 167
rect 256 164 258 178
rect 294 172 300 173
rect 294 168 295 172
rect 299 168 300 172
rect 294 167 300 168
rect 254 163 260 164
rect 254 159 255 163
rect 259 159 260 163
rect 254 158 260 159
rect 296 139 298 167
rect 336 156 338 234
rect 366 224 372 225
rect 366 220 367 224
rect 371 220 372 224
rect 366 219 372 220
rect 414 224 420 225
rect 414 220 415 224
rect 419 220 420 224
rect 414 219 420 220
rect 470 224 476 225
rect 470 220 471 224
rect 475 220 476 224
rect 470 219 476 220
rect 534 224 540 225
rect 534 220 535 224
rect 539 220 540 224
rect 534 219 540 220
rect 606 224 612 225
rect 606 220 607 224
rect 611 220 612 224
rect 606 219 612 220
rect 678 224 684 225
rect 678 220 679 224
rect 683 220 684 224
rect 678 219 684 220
rect 368 207 370 219
rect 416 207 418 219
rect 472 207 474 219
rect 536 207 538 219
rect 608 207 610 219
rect 680 207 682 219
rect 343 206 347 207
rect 343 201 347 202
rect 367 206 371 207
rect 367 201 371 202
rect 399 206 403 207
rect 399 201 403 202
rect 415 206 419 207
rect 415 201 419 202
rect 463 206 467 207
rect 463 201 467 202
rect 471 206 475 207
rect 471 201 475 202
rect 527 206 531 207
rect 527 201 531 202
rect 535 206 539 207
rect 535 201 539 202
rect 599 206 603 207
rect 599 201 603 202
rect 607 206 611 207
rect 607 201 611 202
rect 671 206 675 207
rect 671 201 675 202
rect 679 206 683 207
rect 679 201 683 202
rect 342 200 348 201
rect 342 196 343 200
rect 347 196 348 200
rect 342 195 348 196
rect 398 200 404 201
rect 398 196 399 200
rect 403 196 404 200
rect 398 195 404 196
rect 462 200 468 201
rect 462 196 463 200
rect 467 196 468 200
rect 462 195 468 196
rect 526 200 532 201
rect 526 196 527 200
rect 531 196 532 200
rect 526 195 532 196
rect 598 200 604 201
rect 598 196 599 200
rect 603 196 604 200
rect 598 195 604 196
rect 670 200 676 201
rect 670 196 671 200
rect 675 196 676 200
rect 670 195 676 196
rect 700 184 702 254
rect 708 240 710 282
rect 736 271 738 291
rect 735 270 739 271
rect 735 265 739 266
rect 743 270 747 271
rect 743 265 747 266
rect 744 253 746 265
rect 764 260 766 302
rect 772 288 774 302
rect 782 296 788 297
rect 782 292 783 296
rect 787 292 788 296
rect 782 291 788 292
rect 830 296 836 297
rect 830 292 831 296
rect 835 292 836 296
rect 830 291 836 292
rect 878 296 884 297
rect 878 292 879 296
rect 883 292 884 296
rect 878 291 884 292
rect 926 296 932 297
rect 926 292 927 296
rect 931 292 932 296
rect 926 291 932 292
rect 966 296 972 297
rect 966 292 967 296
rect 971 292 972 296
rect 966 291 972 292
rect 770 287 776 288
rect 770 283 771 287
rect 775 283 776 287
rect 770 282 776 283
rect 784 271 786 291
rect 832 271 834 291
rect 880 271 882 291
rect 886 287 892 288
rect 886 283 887 287
rect 891 283 892 287
rect 886 282 892 283
rect 783 270 787 271
rect 783 265 787 266
rect 807 270 811 271
rect 807 265 811 266
rect 831 270 835 271
rect 831 265 835 266
rect 863 270 867 271
rect 863 265 867 266
rect 879 270 883 271
rect 879 265 883 266
rect 762 259 768 260
rect 762 255 763 259
rect 767 255 768 259
rect 762 254 768 255
rect 808 253 810 265
rect 864 253 866 265
rect 742 252 748 253
rect 742 248 743 252
rect 747 248 748 252
rect 742 247 748 248
rect 806 252 812 253
rect 806 248 807 252
rect 811 248 812 252
rect 806 247 812 248
rect 862 252 868 253
rect 862 248 863 252
rect 867 248 868 252
rect 862 247 868 248
rect 888 240 890 282
rect 928 271 930 291
rect 968 271 970 291
rect 976 288 978 302
rect 1006 296 1012 297
rect 1006 292 1007 296
rect 1011 292 1012 296
rect 1006 291 1012 292
rect 974 287 980 288
rect 974 283 975 287
rect 979 283 980 287
rect 974 282 980 283
rect 1008 271 1010 291
rect 1016 288 1018 302
rect 1046 296 1052 297
rect 1046 292 1047 296
rect 1051 292 1052 296
rect 1046 291 1052 292
rect 1014 287 1020 288
rect 1014 283 1015 287
rect 1019 283 1020 287
rect 1014 282 1020 283
rect 1048 271 1050 291
rect 1056 288 1058 302
rect 1072 288 1074 350
rect 1136 349 1138 369
rect 1160 357 1162 369
rect 1158 356 1164 357
rect 1158 352 1159 356
rect 1163 352 1164 356
rect 1158 351 1164 352
rect 1134 348 1140 349
rect 1134 344 1135 348
rect 1139 344 1140 348
rect 1184 344 1186 370
rect 1199 369 1203 370
rect 1247 374 1251 375
rect 1247 369 1251 370
rect 1255 374 1259 375
rect 1255 369 1259 370
rect 1335 374 1339 375
rect 1342 374 1348 375
rect 1359 374 1363 375
rect 1335 369 1339 370
rect 1359 369 1363 370
rect 1415 374 1419 375
rect 1415 369 1419 370
rect 1463 374 1467 375
rect 1463 369 1467 370
rect 1248 357 1250 369
rect 1262 363 1268 364
rect 1262 359 1263 363
rect 1267 359 1268 363
rect 1262 358 1268 359
rect 1326 363 1332 364
rect 1326 359 1327 363
rect 1331 359 1332 363
rect 1326 358 1332 359
rect 1246 356 1252 357
rect 1246 352 1247 356
rect 1251 352 1252 356
rect 1246 351 1252 352
rect 1264 344 1266 358
rect 1328 344 1330 358
rect 1360 357 1362 369
rect 1464 357 1466 369
rect 1488 364 1490 410
rect 1502 396 1508 397
rect 1502 392 1503 396
rect 1507 392 1508 396
rect 1502 391 1508 392
rect 1590 396 1596 397
rect 1590 392 1591 396
rect 1595 392 1596 396
rect 1590 391 1596 392
rect 1504 375 1506 391
rect 1592 375 1594 391
rect 1612 388 1614 446
rect 1646 436 1652 437
rect 1646 432 1647 436
rect 1651 432 1652 436
rect 1646 431 1652 432
rect 1718 436 1724 437
rect 1718 432 1719 436
rect 1723 432 1724 436
rect 1718 431 1724 432
rect 1806 436 1812 437
rect 1806 432 1807 436
rect 1811 432 1812 436
rect 1806 431 1812 432
rect 1894 436 1900 437
rect 1894 432 1895 436
rect 1899 432 1900 436
rect 1894 431 1900 432
rect 1990 436 1996 437
rect 1990 432 1991 436
rect 1995 432 1996 436
rect 1990 431 1996 432
rect 1647 430 1651 431
rect 1647 425 1651 426
rect 1671 430 1675 431
rect 1671 425 1675 426
rect 1719 430 1723 431
rect 1719 425 1723 426
rect 1751 430 1755 431
rect 1751 425 1755 426
rect 1807 430 1811 431
rect 1807 425 1811 426
rect 1831 430 1835 431
rect 1831 425 1835 426
rect 1895 430 1899 431
rect 1895 425 1899 426
rect 1911 430 1915 431
rect 1911 425 1915 426
rect 1991 430 1995 431
rect 1991 425 1995 426
rect 1999 430 2003 431
rect 1999 425 2003 426
rect 1670 424 1676 425
rect 1670 420 1671 424
rect 1675 420 1676 424
rect 1670 419 1676 420
rect 1750 424 1756 425
rect 1750 420 1751 424
rect 1755 420 1756 424
rect 1750 419 1756 420
rect 1830 424 1836 425
rect 1830 420 1831 424
rect 1835 420 1836 424
rect 1830 419 1836 420
rect 1910 424 1916 425
rect 1910 420 1911 424
rect 1915 420 1916 424
rect 1910 419 1916 420
rect 1998 424 2004 425
rect 1998 420 1999 424
rect 2003 420 2004 424
rect 1998 419 2004 420
rect 1854 415 1860 416
rect 1854 411 1855 415
rect 1859 411 1860 415
rect 1854 410 1860 411
rect 1686 407 1692 408
rect 1686 403 1687 407
rect 1691 403 1692 407
rect 1686 402 1692 403
rect 1706 407 1712 408
rect 1706 403 1707 407
rect 1711 403 1712 407
rect 1706 402 1712 403
rect 1670 396 1676 397
rect 1670 392 1671 396
rect 1675 392 1676 396
rect 1670 391 1676 392
rect 1610 387 1616 388
rect 1610 383 1611 387
rect 1615 383 1616 387
rect 1610 382 1616 383
rect 1672 375 1674 391
rect 1503 374 1507 375
rect 1503 369 1507 370
rect 1559 374 1563 375
rect 1559 369 1563 370
rect 1591 374 1595 375
rect 1591 369 1595 370
rect 1647 374 1651 375
rect 1647 369 1651 370
rect 1671 374 1675 375
rect 1671 369 1675 370
rect 1478 363 1484 364
rect 1478 359 1479 363
rect 1483 359 1484 363
rect 1478 358 1484 359
rect 1486 363 1492 364
rect 1486 359 1487 363
rect 1491 359 1492 363
rect 1486 358 1492 359
rect 1358 356 1364 357
rect 1358 352 1359 356
rect 1363 352 1364 356
rect 1358 351 1364 352
rect 1462 356 1468 357
rect 1462 352 1463 356
rect 1467 352 1468 356
rect 1462 351 1468 352
rect 1480 344 1482 358
rect 1560 357 1562 369
rect 1648 357 1650 369
rect 1688 368 1690 402
rect 1708 388 1710 402
rect 1750 396 1756 397
rect 1750 392 1751 396
rect 1755 392 1756 396
rect 1750 391 1756 392
rect 1830 396 1836 397
rect 1830 392 1831 396
rect 1835 392 1836 396
rect 1830 391 1836 392
rect 1706 387 1712 388
rect 1706 383 1707 387
rect 1711 383 1712 387
rect 1706 382 1712 383
rect 1752 375 1754 391
rect 1832 375 1834 391
rect 1856 388 1858 410
rect 2020 408 2022 466
rect 2072 465 2074 477
rect 2096 472 2098 506
rect 2118 504 2119 508
rect 2123 504 2124 508
rect 2118 503 2124 504
rect 2120 483 2122 503
rect 2119 482 2123 483
rect 2119 477 2123 478
rect 2094 471 2100 472
rect 2094 467 2095 471
rect 2099 467 2100 471
rect 2094 466 2100 467
rect 2070 464 2076 465
rect 2070 460 2071 464
rect 2075 460 2076 464
rect 2070 459 2076 460
rect 2120 457 2122 477
rect 2118 456 2124 457
rect 2118 452 2119 456
rect 2123 452 2124 456
rect 2094 451 2100 452
rect 2118 451 2124 452
rect 2094 447 2095 451
rect 2099 447 2100 451
rect 2094 446 2100 447
rect 2070 436 2076 437
rect 2070 432 2071 436
rect 2075 432 2076 436
rect 2070 431 2076 432
rect 2071 430 2075 431
rect 2071 425 2075 426
rect 2070 424 2076 425
rect 2070 420 2071 424
rect 2075 420 2076 424
rect 2070 419 2076 420
rect 2010 407 2016 408
rect 2010 403 2011 407
rect 2015 403 2016 407
rect 2010 402 2016 403
rect 2018 407 2024 408
rect 2018 403 2019 407
rect 2023 403 2024 407
rect 2018 402 2024 403
rect 1910 396 1916 397
rect 1910 392 1911 396
rect 1915 392 1916 396
rect 1910 391 1916 392
rect 1998 396 2004 397
rect 1998 392 1999 396
rect 2003 392 2004 396
rect 1998 391 2004 392
rect 1854 387 1860 388
rect 1854 383 1855 387
rect 1859 383 1860 387
rect 1854 382 1860 383
rect 1912 375 1914 391
rect 1938 387 1944 388
rect 1938 383 1939 387
rect 1943 383 1944 387
rect 1938 382 1944 383
rect 1727 374 1731 375
rect 1727 369 1731 370
rect 1751 374 1755 375
rect 1751 369 1755 370
rect 1799 374 1803 375
rect 1799 369 1803 370
rect 1831 374 1835 375
rect 1831 369 1835 370
rect 1863 374 1867 375
rect 1863 369 1867 370
rect 1911 374 1915 375
rect 1911 369 1915 370
rect 1919 374 1923 375
rect 1919 369 1923 370
rect 1686 367 1692 368
rect 1662 363 1668 364
rect 1662 359 1663 363
rect 1667 359 1668 363
rect 1686 363 1687 367
rect 1691 363 1692 367
rect 1686 362 1692 363
rect 1662 358 1668 359
rect 1558 356 1564 357
rect 1558 352 1559 356
rect 1563 352 1564 356
rect 1558 351 1564 352
rect 1646 356 1652 357
rect 1646 352 1647 356
rect 1651 352 1652 356
rect 1646 351 1652 352
rect 1664 344 1666 358
rect 1728 357 1730 369
rect 1800 357 1802 369
rect 1864 357 1866 369
rect 1920 357 1922 369
rect 1726 356 1732 357
rect 1726 352 1727 356
rect 1731 352 1732 356
rect 1726 351 1732 352
rect 1798 356 1804 357
rect 1798 352 1799 356
rect 1803 352 1804 356
rect 1798 351 1804 352
rect 1862 356 1868 357
rect 1862 352 1863 356
rect 1867 352 1868 356
rect 1862 351 1868 352
rect 1918 356 1924 357
rect 1918 352 1919 356
rect 1923 352 1924 356
rect 1918 351 1924 352
rect 1940 344 1942 382
rect 2000 375 2002 391
rect 2012 388 2014 402
rect 2070 396 2076 397
rect 2070 392 2071 396
rect 2075 392 2076 396
rect 2070 391 2076 392
rect 2010 387 2016 388
rect 2010 383 2011 387
rect 2015 383 2016 387
rect 2010 382 2016 383
rect 2072 375 2074 391
rect 2096 388 2098 446
rect 2118 439 2124 440
rect 2118 435 2119 439
rect 2123 435 2124 439
rect 2118 434 2124 435
rect 2120 431 2122 434
rect 2119 430 2123 431
rect 2119 425 2123 426
rect 2120 422 2122 425
rect 2118 421 2124 422
rect 2118 417 2119 421
rect 2123 417 2124 421
rect 2118 416 2124 417
rect 2118 404 2124 405
rect 2118 400 2119 404
rect 2123 400 2124 404
rect 2118 399 2124 400
rect 2094 387 2100 388
rect 2094 383 2095 387
rect 2099 383 2100 387
rect 2094 382 2100 383
rect 2120 375 2122 399
rect 1975 374 1979 375
rect 1975 369 1979 370
rect 1999 374 2003 375
rect 1999 369 2003 370
rect 2031 374 2035 375
rect 2031 369 2035 370
rect 2071 374 2075 375
rect 2071 369 2075 370
rect 2119 374 2123 375
rect 2119 369 2123 370
rect 1976 357 1978 369
rect 1990 363 1996 364
rect 1990 359 1991 363
rect 1995 359 1996 363
rect 1990 358 1996 359
rect 1974 356 1980 357
rect 1974 352 1975 356
rect 1979 352 1980 356
rect 1974 351 1980 352
rect 1992 344 1994 358
rect 2032 357 2034 369
rect 2046 363 2052 364
rect 2046 359 2047 363
rect 2051 359 2052 363
rect 2046 358 2052 359
rect 2030 356 2036 357
rect 2030 352 2031 356
rect 2035 352 2036 356
rect 2030 351 2036 352
rect 2048 344 2050 358
rect 2072 357 2074 369
rect 2086 363 2092 364
rect 2086 359 2087 363
rect 2091 359 2092 363
rect 2086 358 2092 359
rect 2070 356 2076 357
rect 2070 352 2071 356
rect 2075 352 2076 356
rect 2070 351 2076 352
rect 2088 344 2090 358
rect 2120 349 2122 369
rect 2118 348 2124 349
rect 2118 344 2119 348
rect 2123 344 2124 348
rect 1094 343 1100 344
rect 1134 343 1140 344
rect 1182 343 1188 344
rect 1094 339 1095 343
rect 1099 339 1100 343
rect 1094 338 1100 339
rect 1182 339 1183 343
rect 1187 339 1188 343
rect 1182 338 1188 339
rect 1262 343 1268 344
rect 1262 339 1263 343
rect 1267 339 1268 343
rect 1262 338 1268 339
rect 1326 343 1332 344
rect 1326 339 1327 343
rect 1331 339 1332 343
rect 1326 338 1332 339
rect 1478 343 1484 344
rect 1478 339 1479 343
rect 1483 339 1484 343
rect 1478 338 1484 339
rect 1662 343 1668 344
rect 1662 339 1663 343
rect 1667 339 1668 343
rect 1662 338 1668 339
rect 1910 343 1916 344
rect 1910 339 1911 343
rect 1915 339 1916 343
rect 1910 338 1916 339
rect 1938 343 1944 344
rect 1938 339 1939 343
rect 1943 339 1944 343
rect 1938 338 1944 339
rect 1990 343 1996 344
rect 1990 339 1991 343
rect 1995 339 1996 343
rect 1990 338 1996 339
rect 2046 343 2052 344
rect 2046 339 2047 343
rect 2051 339 2052 343
rect 2046 338 2052 339
rect 2086 343 2092 344
rect 2118 343 2124 344
rect 2086 339 2087 343
rect 2091 339 2092 343
rect 2086 338 2092 339
rect 1096 331 1098 338
rect 1134 331 1140 332
rect 1095 330 1099 331
rect 1134 327 1135 331
rect 1139 327 1140 331
rect 1134 326 1140 327
rect 1158 328 1164 329
rect 1095 325 1099 326
rect 1096 322 1098 325
rect 1094 321 1100 322
rect 1094 317 1095 321
rect 1099 317 1100 321
rect 1094 316 1100 317
rect 1136 315 1138 326
rect 1158 324 1159 328
rect 1163 324 1164 328
rect 1158 323 1164 324
rect 1246 328 1252 329
rect 1246 324 1247 328
rect 1251 324 1252 328
rect 1246 323 1252 324
rect 1358 328 1364 329
rect 1358 324 1359 328
rect 1363 324 1364 328
rect 1358 323 1364 324
rect 1462 328 1468 329
rect 1462 324 1463 328
rect 1467 324 1468 328
rect 1462 323 1468 324
rect 1558 328 1564 329
rect 1558 324 1559 328
rect 1563 324 1564 328
rect 1558 323 1564 324
rect 1646 328 1652 329
rect 1646 324 1647 328
rect 1651 324 1652 328
rect 1646 323 1652 324
rect 1726 328 1732 329
rect 1726 324 1727 328
rect 1731 324 1732 328
rect 1726 323 1732 324
rect 1798 328 1804 329
rect 1798 324 1799 328
rect 1803 324 1804 328
rect 1798 323 1804 324
rect 1862 328 1868 329
rect 1862 324 1863 328
rect 1867 324 1868 328
rect 1862 323 1868 324
rect 1160 315 1162 323
rect 1248 315 1250 323
rect 1360 315 1362 323
rect 1464 315 1466 323
rect 1560 315 1562 323
rect 1648 315 1650 323
rect 1728 315 1730 323
rect 1800 315 1802 323
rect 1864 315 1866 323
rect 1135 314 1139 315
rect 1135 309 1139 310
rect 1159 314 1163 315
rect 1159 309 1163 310
rect 1247 314 1251 315
rect 1247 309 1251 310
rect 1351 314 1355 315
rect 1351 309 1355 310
rect 1359 314 1363 315
rect 1359 309 1363 310
rect 1391 314 1395 315
rect 1391 309 1395 310
rect 1431 314 1435 315
rect 1431 309 1435 310
rect 1463 314 1467 315
rect 1463 309 1467 310
rect 1471 314 1475 315
rect 1471 309 1475 310
rect 1511 314 1515 315
rect 1511 309 1515 310
rect 1559 314 1563 315
rect 1559 309 1563 310
rect 1615 314 1619 315
rect 1615 309 1619 310
rect 1647 314 1651 315
rect 1647 309 1651 310
rect 1671 314 1675 315
rect 1671 309 1675 310
rect 1727 314 1731 315
rect 1727 309 1731 310
rect 1735 314 1739 315
rect 1735 309 1739 310
rect 1799 314 1803 315
rect 1799 309 1803 310
rect 1807 314 1811 315
rect 1807 309 1811 310
rect 1863 314 1867 315
rect 1863 309 1867 310
rect 1887 314 1891 315
rect 1887 309 1891 310
rect 1136 306 1138 309
rect 1350 308 1356 309
rect 1134 305 1140 306
rect 1094 304 1100 305
rect 1094 300 1095 304
rect 1099 300 1100 304
rect 1134 301 1135 305
rect 1139 301 1140 305
rect 1350 304 1351 308
rect 1355 304 1356 308
rect 1350 303 1356 304
rect 1390 308 1396 309
rect 1390 304 1391 308
rect 1395 304 1396 308
rect 1390 303 1396 304
rect 1430 308 1436 309
rect 1430 304 1431 308
rect 1435 304 1436 308
rect 1430 303 1436 304
rect 1470 308 1476 309
rect 1470 304 1471 308
rect 1475 304 1476 308
rect 1470 303 1476 304
rect 1510 308 1516 309
rect 1510 304 1511 308
rect 1515 304 1516 308
rect 1510 303 1516 304
rect 1558 308 1564 309
rect 1558 304 1559 308
rect 1563 304 1564 308
rect 1558 303 1564 304
rect 1614 308 1620 309
rect 1614 304 1615 308
rect 1619 304 1620 308
rect 1614 303 1620 304
rect 1670 308 1676 309
rect 1670 304 1671 308
rect 1675 304 1676 308
rect 1670 303 1676 304
rect 1734 308 1740 309
rect 1734 304 1735 308
rect 1739 304 1740 308
rect 1734 303 1740 304
rect 1806 308 1812 309
rect 1806 304 1807 308
rect 1811 304 1812 308
rect 1806 303 1812 304
rect 1886 308 1892 309
rect 1886 304 1887 308
rect 1891 304 1892 308
rect 1886 303 1892 304
rect 1134 300 1140 301
rect 1094 299 1100 300
rect 1054 287 1060 288
rect 1054 283 1055 287
rect 1059 283 1060 287
rect 1054 282 1060 283
rect 1070 287 1076 288
rect 1070 283 1071 287
rect 1075 283 1076 287
rect 1070 282 1076 283
rect 1096 271 1098 299
rect 1374 291 1380 292
rect 1134 288 1140 289
rect 1134 284 1135 288
rect 1139 284 1140 288
rect 1374 287 1375 291
rect 1379 287 1380 291
rect 1374 286 1380 287
rect 1398 291 1404 292
rect 1398 287 1399 291
rect 1403 287 1404 291
rect 1398 286 1404 287
rect 1438 291 1444 292
rect 1438 287 1439 291
rect 1443 287 1444 291
rect 1438 286 1444 287
rect 1478 291 1484 292
rect 1478 287 1479 291
rect 1483 287 1484 291
rect 1478 286 1484 287
rect 1518 291 1524 292
rect 1518 287 1519 291
rect 1523 287 1524 291
rect 1518 286 1524 287
rect 1722 291 1728 292
rect 1722 287 1723 291
rect 1727 287 1728 291
rect 1722 286 1728 287
rect 1134 283 1140 284
rect 927 270 931 271
rect 927 265 931 266
rect 967 270 971 271
rect 967 265 971 266
rect 991 270 995 271
rect 991 265 995 266
rect 1007 270 1011 271
rect 1007 265 1011 266
rect 1047 270 1051 271
rect 1047 265 1051 266
rect 1095 270 1099 271
rect 1095 265 1099 266
rect 928 253 930 265
rect 942 259 948 260
rect 942 255 943 259
rect 947 255 948 259
rect 942 254 948 255
rect 926 252 932 253
rect 926 248 927 252
rect 931 248 932 252
rect 926 247 932 248
rect 944 240 946 254
rect 992 253 994 265
rect 1006 259 1012 260
rect 1006 255 1007 259
rect 1011 255 1012 259
rect 1006 254 1012 255
rect 990 252 996 253
rect 990 248 991 252
rect 995 248 996 252
rect 990 247 996 248
rect 1008 240 1010 254
rect 1048 253 1050 265
rect 1062 259 1068 260
rect 1062 255 1063 259
rect 1067 255 1068 259
rect 1062 254 1068 255
rect 1070 259 1076 260
rect 1070 255 1071 259
rect 1075 255 1076 259
rect 1070 254 1076 255
rect 1046 252 1052 253
rect 1046 248 1047 252
rect 1051 248 1052 252
rect 1046 247 1052 248
rect 1064 240 1066 254
rect 706 239 712 240
rect 706 235 707 239
rect 711 235 712 239
rect 706 234 712 235
rect 778 239 784 240
rect 778 235 779 239
rect 783 235 784 239
rect 778 234 784 235
rect 886 239 892 240
rect 886 235 887 239
rect 891 235 892 239
rect 886 234 892 235
rect 942 239 948 240
rect 942 235 943 239
rect 947 235 948 239
rect 942 234 948 235
rect 1006 239 1012 240
rect 1006 235 1007 239
rect 1011 235 1012 239
rect 1006 234 1012 235
rect 1062 239 1068 240
rect 1062 235 1063 239
rect 1067 235 1068 239
rect 1062 234 1068 235
rect 742 224 748 225
rect 742 220 743 224
rect 747 220 748 224
rect 742 219 748 220
rect 744 207 746 219
rect 743 206 747 207
rect 743 201 747 202
rect 751 206 755 207
rect 751 201 755 202
rect 750 200 756 201
rect 750 196 751 200
rect 755 196 756 200
rect 750 195 756 196
rect 614 183 620 184
rect 614 179 615 183
rect 619 179 620 183
rect 614 178 620 179
rect 678 183 684 184
rect 678 179 679 183
rect 683 179 684 183
rect 678 178 684 179
rect 698 183 704 184
rect 698 179 699 183
rect 703 179 704 183
rect 698 178 704 179
rect 342 172 348 173
rect 342 168 343 172
rect 347 168 348 172
rect 342 167 348 168
rect 398 172 404 173
rect 398 168 399 172
rect 403 168 404 172
rect 398 167 404 168
rect 462 172 468 173
rect 462 168 463 172
rect 467 168 468 172
rect 462 167 468 168
rect 526 172 532 173
rect 526 168 527 172
rect 531 168 532 172
rect 526 167 532 168
rect 598 172 604 173
rect 598 168 599 172
rect 603 168 604 172
rect 598 167 604 168
rect 334 155 340 156
rect 334 151 335 155
rect 339 151 340 155
rect 334 150 340 151
rect 344 139 346 167
rect 400 139 402 167
rect 464 139 466 167
rect 528 139 530 167
rect 554 163 560 164
rect 554 159 555 163
rect 559 159 560 163
rect 554 158 560 159
rect 207 138 211 139
rect 175 133 179 134
rect 194 135 200 136
rect 112 113 114 133
rect 136 121 138 133
rect 176 121 178 133
rect 194 131 195 135
rect 199 131 200 135
rect 207 133 211 134
rect 215 138 219 139
rect 215 133 219 134
rect 247 138 251 139
rect 247 133 251 134
rect 255 138 259 139
rect 255 133 259 134
rect 295 138 299 139
rect 295 133 299 134
rect 335 138 339 139
rect 335 133 339 134
rect 343 138 347 139
rect 343 133 347 134
rect 375 138 379 139
rect 375 133 379 134
rect 399 138 403 139
rect 399 133 403 134
rect 415 138 419 139
rect 415 133 419 134
rect 455 138 459 139
rect 455 133 459 134
rect 463 138 467 139
rect 463 133 467 134
rect 495 138 499 139
rect 495 133 499 134
rect 527 138 531 139
rect 527 133 531 134
rect 535 138 539 139
rect 535 133 539 134
rect 194 130 200 131
rect 190 127 196 128
rect 190 123 191 127
rect 195 123 196 127
rect 190 122 196 123
rect 134 120 140 121
rect 134 116 135 120
rect 139 116 140 120
rect 134 115 140 116
rect 174 120 180 121
rect 174 116 175 120
rect 179 116 180 120
rect 174 115 180 116
rect 110 112 116 113
rect 110 108 111 112
rect 115 108 116 112
rect 192 108 194 122
rect 216 121 218 133
rect 230 127 236 128
rect 230 123 231 127
rect 235 123 236 127
rect 230 122 236 123
rect 214 120 220 121
rect 214 116 215 120
rect 219 116 220 120
rect 214 115 220 116
rect 232 108 234 122
rect 256 121 258 133
rect 270 127 276 128
rect 270 123 271 127
rect 275 123 276 127
rect 270 122 276 123
rect 254 120 260 121
rect 254 116 255 120
rect 259 116 260 120
rect 254 115 260 116
rect 272 108 274 122
rect 296 121 298 133
rect 302 127 308 128
rect 302 123 303 127
rect 307 123 308 127
rect 302 122 308 123
rect 294 120 300 121
rect 294 116 295 120
rect 299 116 300 120
rect 294 115 300 116
rect 304 108 306 122
rect 336 121 338 133
rect 350 127 356 128
rect 350 123 351 127
rect 355 123 356 127
rect 350 122 356 123
rect 334 120 340 121
rect 334 116 335 120
rect 339 116 340 120
rect 334 115 340 116
rect 352 108 354 122
rect 376 121 378 133
rect 390 127 396 128
rect 390 123 391 127
rect 395 123 396 127
rect 390 122 396 123
rect 374 120 380 121
rect 374 116 375 120
rect 379 116 380 120
rect 374 115 380 116
rect 392 108 394 122
rect 416 121 418 133
rect 430 127 436 128
rect 430 123 431 127
rect 435 123 436 127
rect 430 122 436 123
rect 414 120 420 121
rect 414 116 415 120
rect 419 116 420 120
rect 414 115 420 116
rect 432 108 434 122
rect 456 121 458 133
rect 470 127 476 128
rect 470 123 471 127
rect 475 123 476 127
rect 470 122 476 123
rect 454 120 460 121
rect 454 116 455 120
rect 459 116 460 120
rect 454 115 460 116
rect 472 108 474 122
rect 496 121 498 133
rect 510 127 516 128
rect 510 123 511 127
rect 515 123 516 127
rect 510 122 516 123
rect 494 120 500 121
rect 494 116 495 120
rect 499 116 500 120
rect 494 115 500 116
rect 512 108 514 122
rect 536 121 538 133
rect 534 120 540 121
rect 534 116 535 120
rect 539 116 540 120
rect 534 115 540 116
rect 556 108 558 158
rect 600 139 602 167
rect 616 164 618 178
rect 670 172 676 173
rect 670 168 671 172
rect 675 168 676 172
rect 670 167 676 168
rect 614 163 620 164
rect 614 159 615 163
rect 619 159 620 163
rect 614 158 620 159
rect 672 139 674 167
rect 680 164 682 178
rect 750 172 756 173
rect 750 168 751 172
rect 755 168 756 172
rect 750 167 756 168
rect 678 163 684 164
rect 678 159 679 163
rect 683 159 684 163
rect 678 158 684 159
rect 752 139 754 167
rect 780 164 782 234
rect 806 224 812 225
rect 806 220 807 224
rect 811 220 812 224
rect 806 219 812 220
rect 862 224 868 225
rect 862 220 863 224
rect 867 220 868 224
rect 862 219 868 220
rect 926 224 932 225
rect 926 220 927 224
rect 931 220 932 224
rect 926 219 932 220
rect 990 224 996 225
rect 990 220 991 224
rect 995 220 996 224
rect 990 219 996 220
rect 1046 224 1052 225
rect 1046 220 1047 224
rect 1051 220 1052 224
rect 1046 219 1052 220
rect 808 207 810 219
rect 864 207 866 219
rect 928 207 930 219
rect 992 207 994 219
rect 1048 207 1050 219
rect 807 206 811 207
rect 807 201 811 202
rect 831 206 835 207
rect 831 201 835 202
rect 863 206 867 207
rect 863 201 867 202
rect 911 206 915 207
rect 911 201 915 202
rect 927 206 931 207
rect 927 201 931 202
rect 991 206 995 207
rect 991 201 995 202
rect 1047 206 1051 207
rect 1047 201 1051 202
rect 830 200 836 201
rect 830 196 831 200
rect 835 196 836 200
rect 830 195 836 196
rect 910 200 916 201
rect 910 196 911 200
rect 915 196 916 200
rect 910 195 916 196
rect 990 200 996 201
rect 990 196 991 200
rect 995 196 996 200
rect 990 195 996 196
rect 1046 200 1052 201
rect 1046 196 1047 200
rect 1051 196 1052 200
rect 1046 195 1052 196
rect 1072 184 1074 254
rect 1096 245 1098 265
rect 1136 263 1138 283
rect 1350 280 1356 281
rect 1350 276 1351 280
rect 1355 276 1356 280
rect 1350 275 1356 276
rect 1352 263 1354 275
rect 1135 262 1139 263
rect 1135 257 1139 258
rect 1263 262 1267 263
rect 1263 257 1267 258
rect 1303 262 1307 263
rect 1303 257 1307 258
rect 1343 262 1347 263
rect 1343 257 1347 258
rect 1351 262 1355 263
rect 1376 260 1378 286
rect 1390 280 1396 281
rect 1390 276 1391 280
rect 1395 276 1396 280
rect 1390 275 1396 276
rect 1392 263 1394 275
rect 1400 272 1402 286
rect 1430 280 1436 281
rect 1430 276 1431 280
rect 1435 276 1436 280
rect 1430 275 1436 276
rect 1398 271 1404 272
rect 1398 267 1399 271
rect 1403 267 1404 271
rect 1398 266 1404 267
rect 1432 263 1434 275
rect 1440 272 1442 286
rect 1470 280 1476 281
rect 1470 276 1471 280
rect 1475 276 1476 280
rect 1470 275 1476 276
rect 1438 271 1444 272
rect 1438 267 1439 271
rect 1443 267 1444 271
rect 1438 266 1444 267
rect 1472 263 1474 275
rect 1480 272 1482 286
rect 1510 280 1516 281
rect 1510 276 1511 280
rect 1515 276 1516 280
rect 1510 275 1516 276
rect 1478 271 1484 272
rect 1478 267 1479 271
rect 1483 267 1484 271
rect 1478 266 1484 267
rect 1512 263 1514 275
rect 1520 272 1522 286
rect 1558 280 1564 281
rect 1558 276 1559 280
rect 1563 276 1564 280
rect 1558 275 1564 276
rect 1614 280 1620 281
rect 1614 276 1615 280
rect 1619 276 1620 280
rect 1614 275 1620 276
rect 1670 280 1676 281
rect 1670 276 1671 280
rect 1675 276 1676 280
rect 1670 275 1676 276
rect 1518 271 1524 272
rect 1518 267 1519 271
rect 1523 267 1524 271
rect 1518 266 1524 267
rect 1560 263 1562 275
rect 1570 263 1576 264
rect 1616 263 1618 275
rect 1672 263 1674 275
rect 1724 272 1726 286
rect 1734 280 1740 281
rect 1734 276 1735 280
rect 1739 276 1740 280
rect 1734 275 1740 276
rect 1806 280 1812 281
rect 1806 276 1807 280
rect 1811 276 1812 280
rect 1806 275 1812 276
rect 1886 280 1892 281
rect 1886 276 1887 280
rect 1891 276 1892 280
rect 1886 275 1892 276
rect 1722 271 1728 272
rect 1722 267 1723 271
rect 1727 267 1728 271
rect 1722 266 1728 267
rect 1736 263 1738 275
rect 1808 263 1810 275
rect 1888 263 1890 275
rect 1912 272 1914 338
rect 2118 331 2124 332
rect 1918 328 1924 329
rect 1918 324 1919 328
rect 1923 324 1924 328
rect 1918 323 1924 324
rect 1974 328 1980 329
rect 1974 324 1975 328
rect 1979 324 1980 328
rect 1974 323 1980 324
rect 2030 328 2036 329
rect 2030 324 2031 328
rect 2035 324 2036 328
rect 2030 323 2036 324
rect 2070 328 2076 329
rect 2070 324 2071 328
rect 2075 324 2076 328
rect 2118 327 2119 331
rect 2123 327 2124 331
rect 2118 326 2124 327
rect 2070 323 2076 324
rect 1920 315 1922 323
rect 1976 315 1978 323
rect 2032 315 2034 323
rect 2072 315 2074 323
rect 2120 315 2122 326
rect 1919 314 1923 315
rect 1919 309 1923 310
rect 1967 314 1971 315
rect 1967 309 1971 310
rect 1975 314 1979 315
rect 1975 309 1979 310
rect 2031 314 2035 315
rect 2031 309 2035 310
rect 2047 314 2051 315
rect 2047 309 2051 310
rect 2071 314 2075 315
rect 2071 309 2075 310
rect 2119 314 2123 315
rect 2119 309 2123 310
rect 1966 308 1972 309
rect 1966 304 1967 308
rect 1971 304 1972 308
rect 1966 303 1972 304
rect 2046 308 2052 309
rect 2046 304 2047 308
rect 2051 304 2052 308
rect 2120 306 2122 309
rect 2046 303 2052 304
rect 2118 305 2124 306
rect 2118 301 2119 305
rect 2123 301 2124 305
rect 2118 300 2124 301
rect 1982 291 1988 292
rect 1982 287 1983 291
rect 1987 287 1988 291
rect 1982 286 1988 287
rect 2062 291 2068 292
rect 2062 287 2063 291
rect 2067 287 2068 291
rect 2062 286 2068 287
rect 2094 291 2100 292
rect 2094 287 2095 291
rect 2099 287 2100 291
rect 2094 286 2100 287
rect 2118 288 2124 289
rect 1966 280 1972 281
rect 1966 276 1967 280
rect 1971 276 1972 280
rect 1966 275 1972 276
rect 1910 271 1916 272
rect 1910 267 1911 271
rect 1915 267 1916 271
rect 1910 266 1916 267
rect 1968 263 1970 275
rect 1984 272 1986 286
rect 2046 280 2052 281
rect 2046 276 2047 280
rect 2051 276 2052 280
rect 2046 275 2052 276
rect 1982 271 1988 272
rect 1982 267 1983 271
rect 1987 267 1988 271
rect 1982 266 1988 267
rect 2048 263 2050 275
rect 2064 272 2066 286
rect 2062 271 2068 272
rect 2062 267 2063 271
rect 2067 267 2068 271
rect 2062 266 2068 267
rect 1383 262 1387 263
rect 1351 257 1355 258
rect 1374 259 1380 260
rect 1094 244 1100 245
rect 1094 240 1095 244
rect 1099 240 1100 244
rect 1094 239 1100 240
rect 1136 237 1138 257
rect 1264 245 1266 257
rect 1304 245 1306 257
rect 1318 251 1324 252
rect 1318 247 1319 251
rect 1323 247 1324 251
rect 1318 246 1324 247
rect 1262 244 1268 245
rect 1262 240 1263 244
rect 1267 240 1268 244
rect 1262 239 1268 240
rect 1302 244 1308 245
rect 1302 240 1303 244
rect 1307 240 1308 244
rect 1302 239 1308 240
rect 1134 236 1140 237
rect 1134 232 1135 236
rect 1139 232 1140 236
rect 1320 232 1322 246
rect 1344 245 1346 257
rect 1374 255 1375 259
rect 1379 255 1380 259
rect 1383 257 1387 258
rect 1391 262 1395 263
rect 1391 257 1395 258
rect 1423 262 1427 263
rect 1423 257 1427 258
rect 1431 262 1435 263
rect 1431 257 1435 258
rect 1463 262 1467 263
rect 1463 257 1467 258
rect 1471 262 1475 263
rect 1471 257 1475 258
rect 1503 262 1507 263
rect 1503 257 1507 258
rect 1511 262 1515 263
rect 1511 257 1515 258
rect 1543 262 1547 263
rect 1543 257 1547 258
rect 1559 262 1563 263
rect 1570 259 1571 263
rect 1575 259 1576 263
rect 1570 258 1576 259
rect 1599 262 1603 263
rect 1559 257 1563 258
rect 1374 254 1380 255
rect 1358 251 1364 252
rect 1358 247 1359 251
rect 1363 247 1364 251
rect 1358 246 1364 247
rect 1342 244 1348 245
rect 1342 240 1343 244
rect 1347 240 1348 244
rect 1342 239 1348 240
rect 1360 232 1362 246
rect 1384 245 1386 257
rect 1398 251 1404 252
rect 1398 247 1399 251
rect 1403 247 1404 251
rect 1398 246 1404 247
rect 1382 244 1388 245
rect 1382 240 1383 244
rect 1387 240 1388 244
rect 1382 239 1388 240
rect 1400 232 1402 246
rect 1424 245 1426 257
rect 1438 251 1444 252
rect 1438 247 1439 251
rect 1443 247 1444 251
rect 1438 246 1444 247
rect 1422 244 1428 245
rect 1422 240 1423 244
rect 1427 240 1428 244
rect 1422 239 1428 240
rect 1440 232 1442 246
rect 1464 245 1466 257
rect 1478 251 1484 252
rect 1478 247 1479 251
rect 1483 247 1484 251
rect 1478 246 1484 247
rect 1462 244 1468 245
rect 1462 240 1463 244
rect 1467 240 1468 244
rect 1462 239 1468 240
rect 1480 232 1482 246
rect 1504 245 1506 257
rect 1518 251 1524 252
rect 1518 247 1519 251
rect 1523 247 1524 251
rect 1518 246 1524 247
rect 1502 244 1508 245
rect 1502 240 1503 244
rect 1507 240 1508 244
rect 1502 239 1508 240
rect 1520 232 1522 246
rect 1544 245 1546 257
rect 1542 244 1548 245
rect 1542 240 1543 244
rect 1547 240 1548 244
rect 1542 239 1548 240
rect 1572 232 1574 258
rect 1599 257 1603 258
rect 1615 262 1619 263
rect 1615 257 1619 258
rect 1671 262 1675 263
rect 1671 257 1675 258
rect 1735 262 1739 263
rect 1735 257 1739 258
rect 1759 262 1763 263
rect 1759 257 1763 258
rect 1807 262 1811 263
rect 1807 257 1811 258
rect 1863 262 1867 263
rect 1863 257 1867 258
rect 1887 262 1891 263
rect 1887 257 1891 258
rect 1967 262 1971 263
rect 1967 257 1971 258
rect 1975 262 1979 263
rect 1975 257 1979 258
rect 2047 262 2051 263
rect 2047 257 2051 258
rect 2071 262 2075 263
rect 2071 257 2075 258
rect 1600 245 1602 257
rect 1614 251 1620 252
rect 1614 247 1615 251
rect 1619 247 1620 251
rect 1614 246 1620 247
rect 1598 244 1604 245
rect 1598 240 1599 244
rect 1603 240 1604 244
rect 1598 239 1604 240
rect 1616 232 1618 246
rect 1672 245 1674 257
rect 1686 251 1692 252
rect 1686 247 1687 251
rect 1691 247 1692 251
rect 1686 246 1692 247
rect 1670 244 1676 245
rect 1670 240 1671 244
rect 1675 240 1676 244
rect 1670 239 1676 240
rect 1688 232 1690 246
rect 1760 245 1762 257
rect 1774 251 1780 252
rect 1774 247 1775 251
rect 1779 247 1780 251
rect 1774 246 1780 247
rect 1758 244 1764 245
rect 1758 240 1759 244
rect 1763 240 1764 244
rect 1758 239 1764 240
rect 1776 232 1778 246
rect 1864 245 1866 257
rect 1878 251 1884 252
rect 1878 247 1879 251
rect 1883 247 1884 251
rect 1878 246 1884 247
rect 1862 244 1868 245
rect 1862 240 1863 244
rect 1867 240 1868 244
rect 1862 239 1868 240
rect 1880 232 1882 246
rect 1976 245 1978 257
rect 1998 251 2004 252
rect 1998 247 1999 251
rect 2003 247 2004 251
rect 1998 246 2004 247
rect 1974 244 1980 245
rect 1974 240 1975 244
rect 1979 240 1980 244
rect 1974 239 1980 240
rect 1134 231 1140 232
rect 1310 231 1316 232
rect 1094 227 1100 228
rect 1094 223 1095 227
rect 1099 223 1100 227
rect 1310 227 1311 231
rect 1315 227 1316 231
rect 1310 226 1316 227
rect 1318 231 1324 232
rect 1318 227 1319 231
rect 1323 227 1324 231
rect 1318 226 1324 227
rect 1358 231 1364 232
rect 1358 227 1359 231
rect 1363 227 1364 231
rect 1358 226 1364 227
rect 1398 231 1404 232
rect 1398 227 1399 231
rect 1403 227 1404 231
rect 1398 226 1404 227
rect 1438 231 1444 232
rect 1438 227 1439 231
rect 1443 227 1444 231
rect 1438 226 1444 227
rect 1478 231 1484 232
rect 1478 227 1479 231
rect 1483 227 1484 231
rect 1478 226 1484 227
rect 1518 231 1524 232
rect 1518 227 1519 231
rect 1523 227 1524 231
rect 1518 226 1524 227
rect 1570 231 1576 232
rect 1570 227 1571 231
rect 1575 227 1576 231
rect 1570 226 1576 227
rect 1614 231 1620 232
rect 1614 227 1615 231
rect 1619 227 1620 231
rect 1614 226 1620 227
rect 1686 231 1692 232
rect 1686 227 1687 231
rect 1691 227 1692 231
rect 1686 226 1692 227
rect 1774 231 1780 232
rect 1774 227 1775 231
rect 1779 227 1780 231
rect 1774 226 1780 227
rect 1878 231 1884 232
rect 1878 227 1879 231
rect 1883 227 1884 231
rect 1878 226 1884 227
rect 1094 222 1100 223
rect 1096 207 1098 222
rect 1134 219 1140 220
rect 1134 215 1135 219
rect 1139 215 1140 219
rect 1134 214 1140 215
rect 1262 216 1268 217
rect 1136 207 1138 214
rect 1262 212 1263 216
rect 1267 212 1268 216
rect 1262 211 1268 212
rect 1302 216 1308 217
rect 1302 212 1303 216
rect 1307 212 1308 216
rect 1302 211 1308 212
rect 1264 207 1266 211
rect 1304 207 1306 211
rect 1095 206 1099 207
rect 1095 201 1099 202
rect 1135 206 1139 207
rect 1135 201 1139 202
rect 1183 206 1187 207
rect 1183 201 1187 202
rect 1231 206 1235 207
rect 1231 201 1235 202
rect 1263 206 1267 207
rect 1263 201 1267 202
rect 1295 206 1299 207
rect 1295 201 1299 202
rect 1303 206 1307 207
rect 1303 201 1307 202
rect 1096 198 1098 201
rect 1136 198 1138 201
rect 1182 200 1188 201
rect 1094 197 1100 198
rect 1094 193 1095 197
rect 1099 193 1100 197
rect 1094 192 1100 193
rect 1134 197 1140 198
rect 1134 193 1135 197
rect 1139 193 1140 197
rect 1182 196 1183 200
rect 1187 196 1188 200
rect 1182 195 1188 196
rect 1230 200 1236 201
rect 1230 196 1231 200
rect 1235 196 1236 200
rect 1230 195 1236 196
rect 1294 200 1300 201
rect 1294 196 1295 200
rect 1299 196 1300 200
rect 1294 195 1300 196
rect 1134 192 1140 193
rect 846 183 852 184
rect 846 179 847 183
rect 851 179 852 183
rect 846 178 852 179
rect 926 183 932 184
rect 926 179 927 183
rect 931 179 932 183
rect 926 178 932 179
rect 958 183 964 184
rect 958 179 959 183
rect 963 179 964 183
rect 958 178 964 179
rect 1062 183 1068 184
rect 1062 179 1063 183
rect 1067 179 1068 183
rect 1062 178 1068 179
rect 1070 183 1076 184
rect 1070 179 1071 183
rect 1075 179 1076 183
rect 1210 183 1216 184
rect 1070 178 1076 179
rect 1094 180 1100 181
rect 830 172 836 173
rect 830 168 831 172
rect 835 168 836 172
rect 830 167 836 168
rect 778 163 784 164
rect 778 159 779 163
rect 783 159 784 163
rect 778 158 784 159
rect 832 139 834 167
rect 848 164 850 178
rect 910 172 916 173
rect 910 168 911 172
rect 915 168 916 172
rect 910 167 916 168
rect 846 163 852 164
rect 846 159 847 163
rect 851 159 852 163
rect 846 158 852 159
rect 912 139 914 167
rect 928 164 930 178
rect 926 163 932 164
rect 926 159 927 163
rect 931 159 932 163
rect 926 158 932 159
rect 575 138 579 139
rect 575 133 579 134
rect 599 138 603 139
rect 599 133 603 134
rect 615 138 619 139
rect 615 133 619 134
rect 655 138 659 139
rect 655 133 659 134
rect 671 138 675 139
rect 671 133 675 134
rect 695 138 699 139
rect 695 133 699 134
rect 735 138 739 139
rect 735 133 739 134
rect 751 138 755 139
rect 751 133 755 134
rect 775 138 779 139
rect 775 133 779 134
rect 815 138 819 139
rect 815 133 819 134
rect 831 138 835 139
rect 831 133 835 134
rect 871 138 875 139
rect 871 133 875 134
rect 911 138 915 139
rect 911 133 915 134
rect 935 138 939 139
rect 935 133 939 134
rect 576 121 578 133
rect 590 127 596 128
rect 590 123 591 127
rect 595 123 596 127
rect 590 122 596 123
rect 574 120 580 121
rect 574 116 575 120
rect 579 116 580 120
rect 574 115 580 116
rect 592 108 594 122
rect 616 121 618 133
rect 630 127 636 128
rect 630 123 631 127
rect 635 123 636 127
rect 630 122 636 123
rect 614 120 620 121
rect 614 116 615 120
rect 619 116 620 120
rect 614 115 620 116
rect 632 108 634 122
rect 656 121 658 133
rect 670 127 676 128
rect 670 123 671 127
rect 675 123 676 127
rect 670 122 676 123
rect 654 120 660 121
rect 654 116 655 120
rect 659 116 660 120
rect 654 115 660 116
rect 672 108 674 122
rect 696 121 698 133
rect 710 127 716 128
rect 710 123 711 127
rect 715 123 716 127
rect 710 122 716 123
rect 694 120 700 121
rect 694 116 695 120
rect 699 116 700 120
rect 694 115 700 116
rect 712 108 714 122
rect 736 121 738 133
rect 750 127 756 128
rect 750 123 751 127
rect 755 123 756 127
rect 750 122 756 123
rect 734 120 740 121
rect 734 116 735 120
rect 739 116 740 120
rect 734 115 740 116
rect 752 108 754 122
rect 776 121 778 133
rect 790 127 796 128
rect 790 123 791 127
rect 795 123 796 127
rect 790 122 796 123
rect 774 120 780 121
rect 774 116 775 120
rect 779 116 780 120
rect 774 115 780 116
rect 792 108 794 122
rect 816 121 818 133
rect 830 127 836 128
rect 830 123 831 127
rect 835 123 836 127
rect 830 122 836 123
rect 814 120 820 121
rect 814 116 815 120
rect 819 116 820 120
rect 814 115 820 116
rect 832 108 834 122
rect 872 121 874 133
rect 886 127 892 128
rect 886 123 887 127
rect 891 123 892 127
rect 886 122 892 123
rect 870 120 876 121
rect 870 116 871 120
rect 875 116 876 120
rect 870 115 876 116
rect 888 108 890 122
rect 936 121 938 133
rect 960 128 962 178
rect 990 172 996 173
rect 990 168 991 172
rect 995 168 996 172
rect 990 167 996 168
rect 1046 172 1052 173
rect 1046 168 1047 172
rect 1051 168 1052 172
rect 1046 167 1052 168
rect 992 139 994 167
rect 1018 163 1024 164
rect 1018 159 1019 163
rect 1023 159 1024 163
rect 1018 158 1024 159
rect 991 138 995 139
rect 991 133 995 134
rect 999 138 1003 139
rect 999 133 1003 134
rect 942 127 948 128
rect 942 123 943 127
rect 947 123 948 127
rect 942 122 948 123
rect 958 127 964 128
rect 958 123 959 127
rect 963 123 964 127
rect 958 122 964 123
rect 934 120 940 121
rect 934 116 935 120
rect 939 116 940 120
rect 934 115 940 116
rect 944 108 946 122
rect 1000 121 1002 133
rect 998 120 1004 121
rect 998 116 999 120
rect 1003 116 1004 120
rect 998 115 1004 116
rect 1020 108 1022 158
rect 1048 139 1050 167
rect 1064 164 1066 178
rect 1094 176 1095 180
rect 1099 176 1100 180
rect 1094 175 1100 176
rect 1134 180 1140 181
rect 1134 176 1135 180
rect 1139 176 1140 180
rect 1210 179 1211 183
rect 1215 179 1216 183
rect 1210 178 1216 179
rect 1218 183 1224 184
rect 1218 179 1219 183
rect 1223 179 1224 183
rect 1218 178 1224 179
rect 1134 175 1140 176
rect 1062 163 1068 164
rect 1062 159 1063 163
rect 1067 159 1068 163
rect 1062 158 1068 159
rect 1096 139 1098 175
rect 1047 138 1051 139
rect 1047 133 1051 134
rect 1095 138 1099 139
rect 1095 133 1099 134
rect 1048 121 1050 133
rect 1062 127 1068 128
rect 1062 123 1063 127
rect 1067 123 1068 127
rect 1062 122 1068 123
rect 1046 120 1052 121
rect 1046 116 1047 120
rect 1051 116 1052 120
rect 1046 115 1052 116
rect 1064 108 1066 122
rect 1096 113 1098 133
rect 1136 131 1138 175
rect 1182 172 1188 173
rect 1182 168 1183 172
rect 1187 168 1188 172
rect 1182 167 1188 168
rect 1184 131 1186 167
rect 1135 130 1139 131
rect 1135 125 1139 126
rect 1159 130 1163 131
rect 1183 130 1187 131
rect 1159 125 1163 126
rect 1174 127 1180 128
rect 1094 112 1100 113
rect 1094 108 1095 112
rect 1099 108 1100 112
rect 110 107 116 108
rect 190 107 196 108
rect 190 103 191 107
rect 195 103 196 107
rect 190 102 196 103
rect 230 107 236 108
rect 230 103 231 107
rect 235 103 236 107
rect 230 102 236 103
rect 270 107 276 108
rect 270 103 271 107
rect 275 103 276 107
rect 270 102 276 103
rect 302 107 308 108
rect 302 103 303 107
rect 307 103 308 107
rect 302 102 308 103
rect 350 107 356 108
rect 350 103 351 107
rect 355 103 356 107
rect 350 102 356 103
rect 390 107 396 108
rect 390 103 391 107
rect 395 103 396 107
rect 390 102 396 103
rect 430 107 436 108
rect 430 103 431 107
rect 435 103 436 107
rect 430 102 436 103
rect 470 107 476 108
rect 470 103 471 107
rect 475 103 476 107
rect 470 102 476 103
rect 510 107 516 108
rect 510 103 511 107
rect 515 103 516 107
rect 510 102 516 103
rect 554 107 560 108
rect 554 103 555 107
rect 559 103 560 107
rect 554 102 560 103
rect 590 107 596 108
rect 590 103 591 107
rect 595 103 596 107
rect 590 102 596 103
rect 630 107 636 108
rect 630 103 631 107
rect 635 103 636 107
rect 630 102 636 103
rect 670 107 676 108
rect 670 103 671 107
rect 675 103 676 107
rect 670 102 676 103
rect 710 107 716 108
rect 710 103 711 107
rect 715 103 716 107
rect 710 102 716 103
rect 750 107 756 108
rect 750 103 751 107
rect 755 103 756 107
rect 750 102 756 103
rect 790 107 796 108
rect 790 103 791 107
rect 795 103 796 107
rect 790 102 796 103
rect 830 107 836 108
rect 830 103 831 107
rect 835 103 836 107
rect 830 102 836 103
rect 886 107 892 108
rect 886 103 887 107
rect 891 103 892 107
rect 886 102 892 103
rect 942 107 948 108
rect 942 103 943 107
rect 947 103 948 107
rect 942 102 948 103
rect 1018 107 1024 108
rect 1018 103 1019 107
rect 1023 103 1024 107
rect 1018 102 1024 103
rect 1062 107 1068 108
rect 1094 107 1100 108
rect 1062 103 1063 107
rect 1067 103 1068 107
rect 1136 105 1138 125
rect 1160 113 1162 125
rect 1174 123 1175 127
rect 1179 123 1180 127
rect 1183 125 1187 126
rect 1199 130 1203 131
rect 1212 128 1214 178
rect 1220 164 1222 178
rect 1230 172 1236 173
rect 1230 168 1231 172
rect 1235 168 1236 172
rect 1230 167 1236 168
rect 1294 172 1300 173
rect 1294 168 1295 172
rect 1299 168 1300 172
rect 1294 167 1300 168
rect 1218 163 1224 164
rect 1218 159 1219 163
rect 1223 159 1224 163
rect 1218 158 1224 159
rect 1232 131 1234 167
rect 1296 131 1298 167
rect 1312 156 1314 226
rect 1342 216 1348 217
rect 1342 212 1343 216
rect 1347 212 1348 216
rect 1342 211 1348 212
rect 1382 216 1388 217
rect 1382 212 1383 216
rect 1387 212 1388 216
rect 1382 211 1388 212
rect 1422 216 1428 217
rect 1422 212 1423 216
rect 1427 212 1428 216
rect 1422 211 1428 212
rect 1462 216 1468 217
rect 1462 212 1463 216
rect 1467 212 1468 216
rect 1462 211 1468 212
rect 1502 216 1508 217
rect 1502 212 1503 216
rect 1507 212 1508 216
rect 1502 211 1508 212
rect 1542 216 1548 217
rect 1542 212 1543 216
rect 1547 212 1548 216
rect 1542 211 1548 212
rect 1598 216 1604 217
rect 1598 212 1599 216
rect 1603 212 1604 216
rect 1598 211 1604 212
rect 1670 216 1676 217
rect 1670 212 1671 216
rect 1675 212 1676 216
rect 1670 211 1676 212
rect 1758 216 1764 217
rect 1758 212 1759 216
rect 1763 212 1764 216
rect 1758 211 1764 212
rect 1862 216 1868 217
rect 1862 212 1863 216
rect 1867 212 1868 216
rect 1862 211 1868 212
rect 1974 216 1980 217
rect 1974 212 1975 216
rect 1979 212 1980 216
rect 1974 211 1980 212
rect 1344 207 1346 211
rect 1384 207 1386 211
rect 1424 207 1426 211
rect 1464 207 1466 211
rect 1504 207 1506 211
rect 1544 207 1546 211
rect 1600 207 1602 211
rect 1614 207 1620 208
rect 1672 207 1674 211
rect 1760 207 1762 211
rect 1864 207 1866 211
rect 1976 207 1978 211
rect 2000 208 2002 246
rect 2072 245 2074 257
rect 2096 252 2098 286
rect 2118 284 2119 288
rect 2123 284 2124 288
rect 2118 283 2124 284
rect 2120 263 2122 283
rect 2119 262 2123 263
rect 2119 257 2123 258
rect 2094 251 2100 252
rect 2094 247 2095 251
rect 2099 247 2100 251
rect 2094 246 2100 247
rect 2070 244 2076 245
rect 2070 240 2071 244
rect 2075 240 2076 244
rect 2070 239 2076 240
rect 2120 237 2122 257
rect 2118 236 2124 237
rect 2118 232 2119 236
rect 2123 232 2124 236
rect 2062 231 2068 232
rect 2118 231 2124 232
rect 2062 227 2063 231
rect 2067 227 2068 231
rect 2062 226 2068 227
rect 1998 207 2004 208
rect 1343 206 1347 207
rect 1343 201 1347 202
rect 1359 206 1363 207
rect 1359 201 1363 202
rect 1383 206 1387 207
rect 1383 201 1387 202
rect 1423 206 1427 207
rect 1423 201 1427 202
rect 1431 206 1435 207
rect 1431 201 1435 202
rect 1463 206 1467 207
rect 1463 201 1467 202
rect 1503 206 1507 207
rect 1503 201 1507 202
rect 1511 206 1515 207
rect 1511 201 1515 202
rect 1543 206 1547 207
rect 1543 201 1547 202
rect 1591 206 1595 207
rect 1591 201 1595 202
rect 1599 206 1603 207
rect 1614 203 1615 207
rect 1619 203 1620 207
rect 1614 202 1620 203
rect 1663 206 1667 207
rect 1599 201 1603 202
rect 1358 200 1364 201
rect 1358 196 1359 200
rect 1363 196 1364 200
rect 1358 195 1364 196
rect 1430 200 1436 201
rect 1430 196 1431 200
rect 1435 196 1436 200
rect 1430 195 1436 196
rect 1510 200 1516 201
rect 1510 196 1511 200
rect 1515 196 1516 200
rect 1510 195 1516 196
rect 1590 200 1596 201
rect 1590 196 1591 200
rect 1595 196 1596 200
rect 1590 195 1596 196
rect 1616 184 1618 202
rect 1663 201 1667 202
rect 1671 206 1675 207
rect 1671 201 1675 202
rect 1735 206 1739 207
rect 1735 201 1739 202
rect 1759 206 1763 207
rect 1759 201 1763 202
rect 1807 206 1811 207
rect 1807 201 1811 202
rect 1863 206 1867 207
rect 1863 201 1867 202
rect 1879 206 1883 207
rect 1879 201 1883 202
rect 1951 206 1955 207
rect 1951 201 1955 202
rect 1975 206 1979 207
rect 1998 203 1999 207
rect 2003 203 2004 207
rect 1998 202 2004 203
rect 2023 206 2027 207
rect 1975 201 1979 202
rect 2023 201 2027 202
rect 1662 200 1668 201
rect 1662 196 1663 200
rect 1667 196 1668 200
rect 1662 195 1668 196
rect 1734 200 1740 201
rect 1734 196 1735 200
rect 1739 196 1740 200
rect 1734 195 1740 196
rect 1806 200 1812 201
rect 1806 196 1807 200
rect 1811 196 1812 200
rect 1806 195 1812 196
rect 1878 200 1884 201
rect 1878 196 1879 200
rect 1883 196 1884 200
rect 1878 195 1884 196
rect 1950 200 1956 201
rect 1950 196 1951 200
rect 1955 196 1956 200
rect 1950 195 1956 196
rect 2022 200 2028 201
rect 2022 196 2023 200
rect 2027 196 2028 200
rect 2022 195 2028 196
rect 1974 191 1980 192
rect 1974 187 1975 191
rect 1979 187 1980 191
rect 1974 186 1980 187
rect 1614 183 1620 184
rect 1614 179 1615 183
rect 1619 179 1620 183
rect 1614 178 1620 179
rect 1358 172 1364 173
rect 1358 168 1359 172
rect 1363 168 1364 172
rect 1358 167 1364 168
rect 1430 172 1436 173
rect 1430 168 1431 172
rect 1435 168 1436 172
rect 1430 167 1436 168
rect 1510 172 1516 173
rect 1510 168 1511 172
rect 1515 168 1516 172
rect 1510 167 1516 168
rect 1590 172 1596 173
rect 1590 168 1591 172
rect 1595 168 1596 172
rect 1590 167 1596 168
rect 1662 172 1668 173
rect 1662 168 1663 172
rect 1667 168 1668 172
rect 1662 167 1668 168
rect 1734 172 1740 173
rect 1734 168 1735 172
rect 1739 168 1740 172
rect 1734 167 1740 168
rect 1806 172 1812 173
rect 1806 168 1807 172
rect 1811 168 1812 172
rect 1806 167 1812 168
rect 1878 172 1884 173
rect 1878 168 1879 172
rect 1883 168 1884 172
rect 1878 167 1884 168
rect 1950 172 1956 173
rect 1950 168 1951 172
rect 1955 168 1956 172
rect 1950 167 1956 168
rect 1310 155 1316 156
rect 1310 151 1311 155
rect 1315 151 1316 155
rect 1310 150 1316 151
rect 1360 131 1362 167
rect 1432 131 1434 167
rect 1512 131 1514 167
rect 1592 131 1594 167
rect 1598 155 1604 156
rect 1598 151 1599 155
rect 1603 151 1604 155
rect 1598 150 1604 151
rect 1231 130 1235 131
rect 1199 125 1203 126
rect 1210 127 1216 128
rect 1174 122 1180 123
rect 1158 112 1164 113
rect 1158 108 1159 112
rect 1163 108 1164 112
rect 1158 107 1164 108
rect 1062 102 1068 103
rect 1134 104 1140 105
rect 1134 100 1135 104
rect 1139 100 1140 104
rect 1176 100 1178 122
rect 1200 113 1202 125
rect 1210 123 1211 127
rect 1215 123 1216 127
rect 1231 125 1235 126
rect 1239 130 1243 131
rect 1239 125 1243 126
rect 1279 130 1283 131
rect 1279 125 1283 126
rect 1295 130 1299 131
rect 1295 125 1299 126
rect 1319 130 1323 131
rect 1319 125 1323 126
rect 1359 130 1363 131
rect 1359 125 1363 126
rect 1367 130 1371 131
rect 1367 125 1371 126
rect 1431 130 1435 131
rect 1431 125 1435 126
rect 1495 130 1499 131
rect 1495 125 1499 126
rect 1511 130 1515 131
rect 1511 125 1515 126
rect 1559 130 1563 131
rect 1559 125 1563 126
rect 1591 130 1595 131
rect 1591 125 1595 126
rect 1210 122 1216 123
rect 1214 119 1220 120
rect 1214 115 1215 119
rect 1219 115 1220 119
rect 1214 114 1220 115
rect 1198 112 1204 113
rect 1198 108 1199 112
rect 1203 108 1204 112
rect 1198 107 1204 108
rect 1216 100 1218 114
rect 1240 113 1242 125
rect 1254 119 1260 120
rect 1254 115 1255 119
rect 1259 115 1260 119
rect 1254 114 1260 115
rect 1238 112 1244 113
rect 1238 108 1239 112
rect 1243 108 1244 112
rect 1238 107 1244 108
rect 1256 100 1258 114
rect 1280 113 1282 125
rect 1294 119 1300 120
rect 1294 115 1295 119
rect 1299 115 1300 119
rect 1294 114 1300 115
rect 1278 112 1284 113
rect 1278 108 1279 112
rect 1283 108 1284 112
rect 1278 107 1284 108
rect 1296 100 1298 114
rect 1320 113 1322 125
rect 1334 119 1340 120
rect 1334 115 1335 119
rect 1339 115 1340 119
rect 1334 114 1340 115
rect 1318 112 1324 113
rect 1318 108 1319 112
rect 1323 108 1324 112
rect 1318 107 1324 108
rect 1336 100 1338 114
rect 1368 113 1370 125
rect 1382 119 1388 120
rect 1382 115 1383 119
rect 1387 115 1388 119
rect 1382 114 1388 115
rect 1366 112 1372 113
rect 1366 108 1367 112
rect 1371 108 1372 112
rect 1366 107 1372 108
rect 1384 100 1386 114
rect 1432 113 1434 125
rect 1446 119 1452 120
rect 1446 115 1447 119
rect 1451 115 1452 119
rect 1446 114 1452 115
rect 1430 112 1436 113
rect 1430 108 1431 112
rect 1435 108 1436 112
rect 1430 107 1436 108
rect 1448 100 1450 114
rect 1496 113 1498 125
rect 1502 119 1508 120
rect 1502 115 1503 119
rect 1507 115 1508 119
rect 1502 114 1508 115
rect 1494 112 1500 113
rect 1494 108 1495 112
rect 1499 108 1500 112
rect 1494 107 1500 108
rect 1504 100 1506 114
rect 1560 113 1562 125
rect 1558 112 1564 113
rect 1558 108 1559 112
rect 1563 108 1564 112
rect 1558 107 1564 108
rect 1600 100 1602 150
rect 1664 131 1666 167
rect 1736 131 1738 167
rect 1808 131 1810 167
rect 1880 131 1882 167
rect 1952 131 1954 167
rect 1615 130 1619 131
rect 1615 125 1619 126
rect 1663 130 1667 131
rect 1663 125 1667 126
rect 1671 130 1675 131
rect 1671 125 1675 126
rect 1719 130 1723 131
rect 1719 125 1723 126
rect 1735 130 1739 131
rect 1735 125 1739 126
rect 1767 130 1771 131
rect 1767 125 1771 126
rect 1807 130 1811 131
rect 1807 125 1811 126
rect 1855 130 1859 131
rect 1855 125 1859 126
rect 1879 130 1883 131
rect 1879 125 1883 126
rect 1903 130 1907 131
rect 1903 125 1907 126
rect 1951 130 1955 131
rect 1951 125 1955 126
rect 1616 113 1618 125
rect 1630 119 1636 120
rect 1630 115 1631 119
rect 1635 115 1636 119
rect 1630 114 1636 115
rect 1614 112 1620 113
rect 1614 108 1615 112
rect 1619 108 1620 112
rect 1614 107 1620 108
rect 1632 100 1634 114
rect 1672 113 1674 125
rect 1686 119 1692 120
rect 1686 115 1687 119
rect 1691 115 1692 119
rect 1686 114 1692 115
rect 1670 112 1676 113
rect 1670 108 1671 112
rect 1675 108 1676 112
rect 1670 107 1676 108
rect 1688 100 1690 114
rect 1720 113 1722 125
rect 1734 119 1740 120
rect 1734 115 1735 119
rect 1739 115 1740 119
rect 1734 114 1740 115
rect 1718 112 1724 113
rect 1718 108 1719 112
rect 1723 108 1724 112
rect 1718 107 1724 108
rect 1736 100 1738 114
rect 1768 113 1770 125
rect 1782 119 1788 120
rect 1782 115 1783 119
rect 1787 115 1788 119
rect 1782 114 1788 115
rect 1766 112 1772 113
rect 1766 108 1767 112
rect 1771 108 1772 112
rect 1766 107 1772 108
rect 1784 100 1786 114
rect 1808 113 1810 125
rect 1822 119 1828 120
rect 1822 115 1823 119
rect 1827 115 1828 119
rect 1822 114 1828 115
rect 1806 112 1812 113
rect 1806 108 1807 112
rect 1811 108 1812 112
rect 1806 107 1812 108
rect 1824 100 1826 114
rect 1856 113 1858 125
rect 1870 119 1876 120
rect 1870 115 1871 119
rect 1875 115 1876 119
rect 1870 114 1876 115
rect 1854 112 1860 113
rect 1854 108 1855 112
rect 1859 108 1860 112
rect 1854 107 1860 108
rect 1872 100 1874 114
rect 1904 113 1906 125
rect 1918 119 1924 120
rect 1918 115 1919 119
rect 1923 115 1924 119
rect 1918 114 1924 115
rect 1902 112 1908 113
rect 1902 108 1903 112
rect 1907 108 1908 112
rect 1902 107 1908 108
rect 1920 100 1922 114
rect 1952 113 1954 125
rect 1976 120 1978 186
rect 2022 172 2028 173
rect 2022 168 2023 172
rect 2027 168 2028 172
rect 2022 167 2028 168
rect 2014 163 2020 164
rect 2014 159 2015 163
rect 2019 159 2020 163
rect 2014 158 2020 159
rect 1991 130 1995 131
rect 1991 125 1995 126
rect 1966 119 1972 120
rect 1966 115 1967 119
rect 1971 115 1972 119
rect 1966 114 1972 115
rect 1974 119 1980 120
rect 1974 115 1975 119
rect 1979 115 1980 119
rect 1974 114 1980 115
rect 1950 112 1956 113
rect 1950 108 1951 112
rect 1955 108 1956 112
rect 1950 107 1956 108
rect 1968 100 1970 114
rect 1992 113 1994 125
rect 1990 112 1996 113
rect 1990 108 1991 112
rect 1995 108 1996 112
rect 1990 107 1996 108
rect 2016 100 2018 158
rect 2024 131 2026 167
rect 2064 164 2066 226
rect 2118 219 2124 220
rect 2070 216 2076 217
rect 2070 212 2071 216
rect 2075 212 2076 216
rect 2118 215 2119 219
rect 2123 215 2124 219
rect 2118 214 2124 215
rect 2070 211 2076 212
rect 2072 207 2074 211
rect 2120 207 2122 214
rect 2071 206 2075 207
rect 2071 201 2075 202
rect 2119 206 2123 207
rect 2119 201 2123 202
rect 2070 200 2076 201
rect 2070 196 2071 200
rect 2075 196 2076 200
rect 2120 198 2122 201
rect 2070 195 2076 196
rect 2118 197 2124 198
rect 2118 193 2119 197
rect 2123 193 2124 197
rect 2118 192 2124 193
rect 2086 183 2092 184
rect 2086 179 2087 183
rect 2091 179 2092 183
rect 2086 178 2092 179
rect 2094 183 2100 184
rect 2094 179 2095 183
rect 2099 179 2100 183
rect 2094 178 2100 179
rect 2118 180 2124 181
rect 2070 172 2076 173
rect 2070 168 2071 172
rect 2075 168 2076 172
rect 2070 167 2076 168
rect 2062 163 2068 164
rect 2062 159 2063 163
rect 2067 159 2068 163
rect 2062 158 2068 159
rect 2072 131 2074 167
rect 2088 164 2090 178
rect 2086 163 2092 164
rect 2086 159 2087 163
rect 2091 159 2092 163
rect 2086 158 2092 159
rect 2023 130 2027 131
rect 2023 125 2027 126
rect 2031 130 2035 131
rect 2031 125 2035 126
rect 2071 130 2075 131
rect 2071 125 2075 126
rect 2032 113 2034 125
rect 2046 119 2052 120
rect 2046 115 2047 119
rect 2051 115 2052 119
rect 2046 114 2052 115
rect 2030 112 2036 113
rect 2030 108 2031 112
rect 2035 108 2036 112
rect 2030 107 2036 108
rect 2048 100 2050 114
rect 2072 113 2074 125
rect 2096 120 2098 178
rect 2118 176 2119 180
rect 2123 176 2124 180
rect 2118 175 2124 176
rect 2120 131 2122 175
rect 2119 130 2123 131
rect 2119 125 2123 126
rect 2086 119 2092 120
rect 2086 115 2087 119
rect 2091 115 2092 119
rect 2086 114 2092 115
rect 2094 119 2100 120
rect 2094 115 2095 119
rect 2099 115 2100 119
rect 2094 114 2100 115
rect 2070 112 2076 113
rect 2070 108 2071 112
rect 2075 108 2076 112
rect 2070 107 2076 108
rect 2088 100 2090 114
rect 2120 105 2122 125
rect 2118 104 2124 105
rect 2118 100 2119 104
rect 2123 100 2124 104
rect 1134 99 1140 100
rect 1174 99 1180 100
rect 110 95 116 96
rect 110 91 111 95
rect 115 91 116 95
rect 1094 95 1100 96
rect 110 90 116 91
rect 134 92 140 93
rect 112 87 114 90
rect 134 88 135 92
rect 139 88 140 92
rect 134 87 140 88
rect 174 92 180 93
rect 174 88 175 92
rect 179 88 180 92
rect 174 87 180 88
rect 214 92 220 93
rect 214 88 215 92
rect 219 88 220 92
rect 214 87 220 88
rect 254 92 260 93
rect 254 88 255 92
rect 259 88 260 92
rect 254 87 260 88
rect 294 92 300 93
rect 294 88 295 92
rect 299 88 300 92
rect 294 87 300 88
rect 334 92 340 93
rect 334 88 335 92
rect 339 88 340 92
rect 334 87 340 88
rect 374 92 380 93
rect 374 88 375 92
rect 379 88 380 92
rect 374 87 380 88
rect 414 92 420 93
rect 414 88 415 92
rect 419 88 420 92
rect 414 87 420 88
rect 454 92 460 93
rect 454 88 455 92
rect 459 88 460 92
rect 454 87 460 88
rect 494 92 500 93
rect 494 88 495 92
rect 499 88 500 92
rect 494 87 500 88
rect 534 92 540 93
rect 534 88 535 92
rect 539 88 540 92
rect 534 87 540 88
rect 574 92 580 93
rect 574 88 575 92
rect 579 88 580 92
rect 574 87 580 88
rect 614 92 620 93
rect 614 88 615 92
rect 619 88 620 92
rect 614 87 620 88
rect 654 92 660 93
rect 654 88 655 92
rect 659 88 660 92
rect 654 87 660 88
rect 694 92 700 93
rect 694 88 695 92
rect 699 88 700 92
rect 694 87 700 88
rect 734 92 740 93
rect 734 88 735 92
rect 739 88 740 92
rect 734 87 740 88
rect 774 92 780 93
rect 774 88 775 92
rect 779 88 780 92
rect 774 87 780 88
rect 814 92 820 93
rect 814 88 815 92
rect 819 88 820 92
rect 814 87 820 88
rect 870 92 876 93
rect 870 88 871 92
rect 875 88 876 92
rect 870 87 876 88
rect 934 92 940 93
rect 934 88 935 92
rect 939 88 940 92
rect 934 87 940 88
rect 998 92 1004 93
rect 998 88 999 92
rect 1003 88 1004 92
rect 998 87 1004 88
rect 1046 92 1052 93
rect 1046 88 1047 92
rect 1051 88 1052 92
rect 1094 91 1095 95
rect 1099 91 1100 95
rect 1174 95 1175 99
rect 1179 95 1180 99
rect 1174 94 1180 95
rect 1214 99 1220 100
rect 1214 95 1215 99
rect 1219 95 1220 99
rect 1214 94 1220 95
rect 1254 99 1260 100
rect 1254 95 1255 99
rect 1259 95 1260 99
rect 1254 94 1260 95
rect 1294 99 1300 100
rect 1294 95 1295 99
rect 1299 95 1300 99
rect 1294 94 1300 95
rect 1334 99 1340 100
rect 1334 95 1335 99
rect 1339 95 1340 99
rect 1334 94 1340 95
rect 1382 99 1388 100
rect 1382 95 1383 99
rect 1387 95 1388 99
rect 1382 94 1388 95
rect 1446 99 1452 100
rect 1446 95 1447 99
rect 1451 95 1452 99
rect 1446 94 1452 95
rect 1502 99 1508 100
rect 1502 95 1503 99
rect 1507 95 1508 99
rect 1502 94 1508 95
rect 1598 99 1604 100
rect 1598 95 1599 99
rect 1603 95 1604 99
rect 1598 94 1604 95
rect 1630 99 1636 100
rect 1630 95 1631 99
rect 1635 95 1636 99
rect 1630 94 1636 95
rect 1686 99 1692 100
rect 1686 95 1687 99
rect 1691 95 1692 99
rect 1686 94 1692 95
rect 1734 99 1740 100
rect 1734 95 1735 99
rect 1739 95 1740 99
rect 1734 94 1740 95
rect 1782 99 1788 100
rect 1782 95 1783 99
rect 1787 95 1788 99
rect 1782 94 1788 95
rect 1822 99 1828 100
rect 1822 95 1823 99
rect 1827 95 1828 99
rect 1822 94 1828 95
rect 1870 99 1876 100
rect 1870 95 1871 99
rect 1875 95 1876 99
rect 1870 94 1876 95
rect 1918 99 1924 100
rect 1918 95 1919 99
rect 1923 95 1924 99
rect 1918 94 1924 95
rect 1966 99 1972 100
rect 1966 95 1967 99
rect 1971 95 1972 99
rect 1966 94 1972 95
rect 2014 99 2020 100
rect 2014 95 2015 99
rect 2019 95 2020 99
rect 2014 94 2020 95
rect 2046 99 2052 100
rect 2046 95 2047 99
rect 2051 95 2052 99
rect 2046 94 2052 95
rect 2086 99 2092 100
rect 2118 99 2124 100
rect 2086 95 2087 99
rect 2091 95 2092 99
rect 2086 94 2092 95
rect 1094 90 1100 91
rect 1046 87 1052 88
rect 1096 87 1098 90
rect 1134 87 1140 88
rect 111 86 115 87
rect 111 81 115 82
rect 135 86 139 87
rect 135 81 139 82
rect 175 86 179 87
rect 175 81 179 82
rect 215 86 219 87
rect 215 81 219 82
rect 255 86 259 87
rect 255 81 259 82
rect 295 86 299 87
rect 295 81 299 82
rect 335 86 339 87
rect 335 81 339 82
rect 375 86 379 87
rect 375 81 379 82
rect 415 86 419 87
rect 415 81 419 82
rect 455 86 459 87
rect 455 81 459 82
rect 495 86 499 87
rect 495 81 499 82
rect 535 86 539 87
rect 535 81 539 82
rect 575 86 579 87
rect 575 81 579 82
rect 615 86 619 87
rect 615 81 619 82
rect 655 86 659 87
rect 655 81 659 82
rect 695 86 699 87
rect 695 81 699 82
rect 735 86 739 87
rect 735 81 739 82
rect 775 86 779 87
rect 775 81 779 82
rect 815 86 819 87
rect 815 81 819 82
rect 871 86 875 87
rect 871 81 875 82
rect 935 86 939 87
rect 935 81 939 82
rect 999 86 1003 87
rect 999 81 1003 82
rect 1047 86 1051 87
rect 1047 81 1051 82
rect 1095 86 1099 87
rect 1134 83 1135 87
rect 1139 83 1140 87
rect 2118 87 2124 88
rect 1134 82 1140 83
rect 1158 84 1164 85
rect 1095 81 1099 82
rect 1136 79 1138 82
rect 1158 80 1159 84
rect 1163 80 1164 84
rect 1158 79 1164 80
rect 1198 84 1204 85
rect 1198 80 1199 84
rect 1203 80 1204 84
rect 1198 79 1204 80
rect 1238 84 1244 85
rect 1238 80 1239 84
rect 1243 80 1244 84
rect 1238 79 1244 80
rect 1278 84 1284 85
rect 1278 80 1279 84
rect 1283 80 1284 84
rect 1278 79 1284 80
rect 1318 84 1324 85
rect 1318 80 1319 84
rect 1323 80 1324 84
rect 1318 79 1324 80
rect 1366 84 1372 85
rect 1366 80 1367 84
rect 1371 80 1372 84
rect 1366 79 1372 80
rect 1430 84 1436 85
rect 1430 80 1431 84
rect 1435 80 1436 84
rect 1430 79 1436 80
rect 1494 84 1500 85
rect 1494 80 1495 84
rect 1499 80 1500 84
rect 1494 79 1500 80
rect 1558 84 1564 85
rect 1558 80 1559 84
rect 1563 80 1564 84
rect 1558 79 1564 80
rect 1614 84 1620 85
rect 1614 80 1615 84
rect 1619 80 1620 84
rect 1614 79 1620 80
rect 1670 84 1676 85
rect 1670 80 1671 84
rect 1675 80 1676 84
rect 1670 79 1676 80
rect 1718 84 1724 85
rect 1718 80 1719 84
rect 1723 80 1724 84
rect 1718 79 1724 80
rect 1766 84 1772 85
rect 1766 80 1767 84
rect 1771 80 1772 84
rect 1766 79 1772 80
rect 1806 84 1812 85
rect 1806 80 1807 84
rect 1811 80 1812 84
rect 1806 79 1812 80
rect 1854 84 1860 85
rect 1854 80 1855 84
rect 1859 80 1860 84
rect 1854 79 1860 80
rect 1902 84 1908 85
rect 1902 80 1903 84
rect 1907 80 1908 84
rect 1902 79 1908 80
rect 1950 84 1956 85
rect 1950 80 1951 84
rect 1955 80 1956 84
rect 1950 79 1956 80
rect 1990 84 1996 85
rect 1990 80 1991 84
rect 1995 80 1996 84
rect 1990 79 1996 80
rect 2030 84 2036 85
rect 2030 80 2031 84
rect 2035 80 2036 84
rect 2030 79 2036 80
rect 2070 84 2076 85
rect 2070 80 2071 84
rect 2075 80 2076 84
rect 2118 83 2119 87
rect 2123 83 2124 87
rect 2118 82 2124 83
rect 2070 79 2076 80
rect 2120 79 2122 82
rect 1135 78 1139 79
rect 1135 73 1139 74
rect 1159 78 1163 79
rect 1159 73 1163 74
rect 1199 78 1203 79
rect 1199 73 1203 74
rect 1239 78 1243 79
rect 1239 73 1243 74
rect 1279 78 1283 79
rect 1279 73 1283 74
rect 1319 78 1323 79
rect 1319 73 1323 74
rect 1367 78 1371 79
rect 1367 73 1371 74
rect 1431 78 1435 79
rect 1431 73 1435 74
rect 1495 78 1499 79
rect 1495 73 1499 74
rect 1559 78 1563 79
rect 1559 73 1563 74
rect 1615 78 1619 79
rect 1615 73 1619 74
rect 1671 78 1675 79
rect 1671 73 1675 74
rect 1719 78 1723 79
rect 1719 73 1723 74
rect 1767 78 1771 79
rect 1767 73 1771 74
rect 1807 78 1811 79
rect 1807 73 1811 74
rect 1855 78 1859 79
rect 1855 73 1859 74
rect 1903 78 1907 79
rect 1903 73 1907 74
rect 1951 78 1955 79
rect 1951 73 1955 74
rect 1991 78 1995 79
rect 1991 73 1995 74
rect 2031 78 2035 79
rect 2031 73 2035 74
rect 2071 78 2075 79
rect 2071 73 2075 74
rect 2119 78 2123 79
rect 2119 73 2123 74
<< m4c >>
rect 1135 2210 1139 2214
rect 1343 2210 1347 2214
rect 1383 2210 1387 2214
rect 1423 2210 1427 2214
rect 1463 2210 1467 2214
rect 1503 2210 1507 2214
rect 1543 2210 1547 2214
rect 1583 2210 1587 2214
rect 1623 2210 1627 2214
rect 1663 2210 1667 2214
rect 1703 2210 1707 2214
rect 1743 2210 1747 2214
rect 1783 2210 1787 2214
rect 1823 2210 1827 2214
rect 2119 2210 2123 2214
rect 1135 2158 1139 2162
rect 1287 2158 1291 2162
rect 1327 2158 1331 2162
rect 1343 2158 1347 2162
rect 1367 2158 1371 2162
rect 1383 2158 1387 2162
rect 1315 2112 1319 2116
rect 1415 2158 1419 2162
rect 1423 2158 1427 2162
rect 1463 2158 1467 2162
rect 1503 2158 1507 2162
rect 1519 2158 1523 2162
rect 1543 2158 1547 2162
rect 1575 2158 1579 2162
rect 1583 2158 1587 2162
rect 1623 2158 1627 2162
rect 1663 2158 1667 2162
rect 1671 2158 1675 2162
rect 1703 2158 1707 2162
rect 1719 2158 1723 2162
rect 1743 2158 1747 2162
rect 1775 2158 1779 2162
rect 1783 2158 1787 2162
rect 1823 2158 1827 2162
rect 1831 2158 1835 2162
rect 1887 2158 1891 2162
rect 2119 2158 2123 2162
rect 1607 2112 1611 2116
rect 1135 2102 1139 2106
rect 1223 2102 1227 2106
rect 1279 2102 1283 2106
rect 1287 2102 1291 2106
rect 1327 2102 1331 2106
rect 1343 2102 1347 2106
rect 1367 2102 1371 2106
rect 1415 2102 1419 2106
rect 1423 2102 1427 2106
rect 1463 2102 1467 2106
rect 1503 2102 1507 2106
rect 1519 2102 1523 2106
rect 1575 2102 1579 2106
rect 1583 2102 1587 2106
rect 1623 2102 1627 2106
rect 1663 2102 1667 2106
rect 1671 2102 1675 2106
rect 1719 2102 1723 2106
rect 1743 2102 1747 2106
rect 1775 2102 1779 2106
rect 1831 2102 1835 2106
rect 1887 2102 1891 2106
rect 1919 2102 1923 2106
rect 2007 2102 2011 2106
rect 2071 2102 2075 2106
rect 2119 2102 2123 2106
rect 1135 2050 1139 2054
rect 1183 2050 1187 2054
rect 111 2030 115 2034
rect 191 2030 195 2034
rect 231 2030 235 2034
rect 287 2030 291 2034
rect 351 2030 355 2034
rect 423 2030 427 2034
rect 495 2030 499 2034
rect 575 2030 579 2034
rect 647 2030 651 2034
rect 719 2030 723 2034
rect 783 2030 787 2034
rect 839 2030 843 2034
rect 895 2030 899 2034
rect 951 2030 955 2034
rect 1007 2030 1011 2034
rect 1047 2030 1051 2034
rect 1095 2030 1099 2034
rect 111 1978 115 1982
rect 191 1978 195 1982
rect 231 1978 235 1982
rect 247 1978 251 1982
rect 287 1978 291 1982
rect 311 1978 315 1982
rect 351 1978 355 1982
rect 375 1978 379 1982
rect 423 1978 427 1982
rect 447 1978 451 1982
rect 495 1978 499 1982
rect 519 1978 523 1982
rect 575 1978 579 1982
rect 591 1978 595 1982
rect 647 1978 651 1982
rect 655 1978 659 1982
rect 719 1978 723 1982
rect 775 1978 779 1982
rect 783 1978 787 1982
rect 823 1978 827 1982
rect 839 1978 843 1982
rect 871 1978 875 1982
rect 895 1978 899 1982
rect 919 1978 923 1982
rect 951 1978 955 1982
rect 967 1978 971 1982
rect 1007 1978 1011 1982
rect 1047 1978 1051 1982
rect 1223 2050 1227 2054
rect 1239 2050 1243 2054
rect 1279 2050 1283 2054
rect 1311 2050 1315 2054
rect 1343 2050 1347 2054
rect 1399 2050 1403 2054
rect 1423 2050 1427 2054
rect 1487 2050 1491 2054
rect 1503 2050 1507 2054
rect 1583 2050 1587 2054
rect 1663 2050 1667 2054
rect 1671 2050 1675 2054
rect 1743 2050 1747 2054
rect 1759 2050 1763 2054
rect 1831 2050 1835 2054
rect 1839 2050 1843 2054
rect 1919 2050 1923 2054
rect 2007 2050 2011 2054
rect 1135 1998 1139 2002
rect 1183 1998 1187 2002
rect 1239 1998 1243 2002
rect 1303 1998 1307 2002
rect 1311 1998 1315 2002
rect 1383 1998 1387 2002
rect 1399 1998 1403 2002
rect 1463 1998 1467 2002
rect 1487 1998 1491 2002
rect 1543 1998 1547 2002
rect 1095 1978 1099 1982
rect 1583 1998 1587 2002
rect 1615 1998 1619 2002
rect 1671 1998 1675 2002
rect 1687 1998 1691 2002
rect 1751 1998 1755 2002
rect 1759 1998 1763 2002
rect 1815 1998 1819 2002
rect 1643 1976 1647 1980
rect 111 1926 115 1930
rect 135 1926 139 1930
rect 175 1926 179 1930
rect 191 1926 195 1930
rect 231 1926 235 1930
rect 247 1926 251 1930
rect 295 1926 299 1930
rect 311 1926 315 1930
rect 367 1926 371 1930
rect 375 1926 379 1930
rect 431 1926 435 1930
rect 447 1926 451 1930
rect 495 1926 499 1930
rect 519 1926 523 1930
rect 559 1926 563 1930
rect 591 1926 595 1930
rect 1135 1942 1139 1946
rect 1159 1942 1163 1946
rect 1223 1942 1227 1946
rect 1303 1942 1307 1946
rect 111 1870 115 1874
rect 135 1870 139 1874
rect 175 1870 179 1874
rect 199 1870 203 1874
rect 231 1870 235 1874
rect 271 1870 275 1874
rect 295 1870 299 1874
rect 335 1870 339 1874
rect 367 1870 371 1874
rect 399 1870 403 1874
rect 431 1870 435 1874
rect 455 1870 459 1874
rect 495 1870 499 1874
rect 503 1870 507 1874
rect 111 1810 115 1814
rect 135 1810 139 1814
rect 151 1810 155 1814
rect 199 1810 203 1814
rect 215 1810 219 1814
rect 271 1810 275 1814
rect 327 1810 331 1814
rect 335 1810 339 1814
rect 383 1810 387 1814
rect 399 1810 403 1814
rect 431 1810 435 1814
rect 111 1758 115 1762
rect 151 1758 155 1762
rect 215 1758 219 1762
rect 231 1758 235 1762
rect 271 1758 275 1762
rect 295 1758 299 1762
rect 327 1758 331 1762
rect 351 1758 355 1762
rect 615 1926 619 1930
rect 655 1926 659 1930
rect 671 1926 675 1930
rect 719 1926 723 1930
rect 727 1926 731 1930
rect 775 1926 779 1930
rect 783 1926 787 1930
rect 823 1926 827 1930
rect 847 1926 851 1930
rect 871 1926 875 1930
rect 919 1926 923 1930
rect 967 1926 971 1930
rect 1007 1926 1011 1930
rect 1047 1926 1051 1930
rect 1095 1926 1099 1930
rect 551 1870 555 1874
rect 559 1870 563 1874
rect 599 1870 603 1874
rect 615 1870 619 1874
rect 455 1810 459 1814
rect 479 1810 483 1814
rect 503 1810 507 1814
rect 1135 1886 1139 1890
rect 1159 1886 1163 1890
rect 1199 1886 1203 1890
rect 647 1870 651 1874
rect 671 1870 675 1874
rect 695 1870 699 1874
rect 727 1870 731 1874
rect 751 1870 755 1874
rect 783 1870 787 1874
rect 847 1870 851 1874
rect 1095 1870 1099 1874
rect 1383 1942 1387 1946
rect 1463 1942 1467 1946
rect 1535 1942 1539 1946
rect 1543 1942 1547 1946
rect 1615 1942 1619 1946
rect 1687 1942 1691 1946
rect 1695 1942 1699 1946
rect 1751 1942 1755 1946
rect 1783 1942 1787 1946
rect 2071 2050 2075 2054
rect 2119 2050 2123 2054
rect 1839 1998 1843 2002
rect 1879 1998 1883 2002
rect 1919 1998 1923 2002
rect 1951 1998 1955 2002
rect 2007 1998 2011 2002
rect 2023 1998 2027 2002
rect 2071 1998 2075 2002
rect 2119 1998 2123 2002
rect 1975 1976 1979 1980
rect 1815 1942 1819 1946
rect 1879 1942 1883 1946
rect 1951 1942 1955 1946
rect 1983 1942 1987 1946
rect 2023 1942 2027 1946
rect 2071 1942 2075 1946
rect 1223 1886 1227 1890
rect 1263 1886 1267 1890
rect 1303 1886 1307 1890
rect 1327 1886 1331 1890
rect 1383 1886 1387 1890
rect 1391 1886 1395 1890
rect 1447 1886 1451 1890
rect 1463 1886 1467 1890
rect 1135 1834 1139 1838
rect 1159 1834 1163 1838
rect 1199 1834 1203 1838
rect 1231 1834 1235 1838
rect 1263 1834 1267 1838
rect 1303 1834 1307 1838
rect 1503 1886 1507 1890
rect 1535 1886 1539 1890
rect 1559 1886 1563 1890
rect 1615 1886 1619 1890
rect 1631 1886 1635 1890
rect 1695 1886 1699 1890
rect 1711 1886 1715 1890
rect 1327 1834 1331 1838
rect 1383 1834 1387 1838
rect 1391 1834 1395 1838
rect 527 1810 531 1814
rect 551 1810 555 1814
rect 575 1810 579 1814
rect 599 1810 603 1814
rect 623 1810 627 1814
rect 647 1810 651 1814
rect 671 1810 675 1814
rect 695 1810 699 1814
rect 727 1810 731 1814
rect 751 1810 755 1814
rect 1095 1810 1099 1814
rect 1135 1782 1139 1786
rect 1159 1782 1163 1786
rect 1191 1782 1195 1786
rect 383 1758 387 1762
rect 415 1758 419 1762
rect 431 1758 435 1762
rect 479 1758 483 1762
rect 527 1758 531 1762
rect 543 1758 547 1762
rect 575 1758 579 1762
rect 615 1758 619 1762
rect 623 1758 627 1762
rect 671 1758 675 1762
rect 687 1758 691 1762
rect 727 1758 731 1762
rect 759 1758 763 1762
rect 111 1702 115 1706
rect 135 1702 139 1706
rect 199 1702 203 1706
rect 231 1702 235 1706
rect 279 1702 283 1706
rect 295 1702 299 1706
rect 351 1702 355 1706
rect 367 1702 371 1706
rect 415 1702 419 1706
rect 463 1702 467 1706
rect 479 1702 483 1706
rect 543 1702 547 1706
rect 551 1702 555 1706
rect 111 1646 115 1650
rect 135 1646 139 1650
rect 183 1646 187 1650
rect 111 1594 115 1598
rect 135 1594 139 1598
rect 199 1646 203 1650
rect 263 1646 267 1650
rect 279 1646 283 1650
rect 615 1702 619 1706
rect 639 1702 643 1706
rect 831 1758 835 1762
rect 911 1758 915 1762
rect 991 1758 995 1762
rect 1095 1758 1099 1762
rect 1447 1834 1451 1838
rect 1463 1834 1467 1838
rect 1503 1834 1507 1838
rect 1551 1834 1555 1838
rect 1559 1834 1563 1838
rect 1631 1834 1635 1838
rect 1647 1834 1651 1838
rect 2119 1942 2123 1946
rect 1783 1886 1787 1890
rect 1799 1886 1803 1890
rect 1879 1886 1883 1890
rect 1895 1886 1899 1890
rect 1983 1886 1987 1890
rect 1991 1886 1995 1890
rect 2071 1886 2075 1890
rect 2119 1886 2123 1890
rect 1711 1834 1715 1838
rect 1751 1834 1755 1838
rect 1799 1834 1803 1838
rect 1855 1834 1859 1838
rect 1895 1834 1899 1838
rect 1967 1834 1971 1838
rect 1991 1834 1995 1838
rect 2071 1834 2075 1838
rect 1231 1782 1235 1786
rect 1255 1782 1259 1786
rect 1303 1782 1307 1786
rect 1319 1782 1323 1786
rect 1383 1782 1387 1786
rect 1455 1782 1459 1786
rect 1463 1782 1467 1786
rect 1527 1782 1531 1786
rect 1551 1782 1555 1786
rect 687 1702 691 1706
rect 719 1702 723 1706
rect 759 1702 763 1706
rect 791 1702 795 1706
rect 831 1702 835 1706
rect 855 1702 859 1706
rect 911 1702 915 1706
rect 919 1702 923 1706
rect 983 1702 987 1706
rect 991 1702 995 1706
rect 343 1646 347 1650
rect 367 1646 371 1650
rect 423 1646 427 1650
rect 463 1646 467 1650
rect 503 1646 507 1650
rect 551 1646 555 1650
rect 583 1646 587 1650
rect 175 1594 179 1598
rect 183 1594 187 1598
rect 231 1594 235 1598
rect 263 1594 267 1598
rect 303 1594 307 1598
rect 343 1594 347 1598
rect 375 1594 379 1598
rect 423 1594 427 1598
rect 455 1594 459 1598
rect 639 1646 643 1650
rect 655 1646 659 1650
rect 719 1646 723 1650
rect 727 1646 731 1650
rect 791 1646 795 1650
rect 847 1646 851 1650
rect 855 1646 859 1650
rect 1135 1730 1139 1734
rect 1191 1730 1195 1734
rect 1247 1730 1251 1734
rect 1255 1730 1259 1734
rect 1295 1730 1299 1734
rect 1319 1730 1323 1734
rect 1343 1730 1347 1734
rect 1607 1782 1611 1786
rect 1647 1782 1651 1786
rect 1687 1782 1691 1786
rect 1383 1730 1387 1734
rect 1399 1730 1403 1734
rect 1047 1702 1051 1706
rect 1095 1702 1099 1706
rect 1135 1674 1139 1678
rect 1247 1674 1251 1678
rect 1263 1674 1267 1678
rect 903 1646 907 1650
rect 919 1646 923 1650
rect 959 1646 963 1650
rect 983 1646 987 1650
rect 1007 1646 1011 1650
rect 503 1594 507 1598
rect 527 1594 531 1598
rect 583 1594 587 1598
rect 599 1594 603 1598
rect 655 1594 659 1598
rect 671 1594 675 1598
rect 727 1594 731 1598
rect 743 1594 747 1598
rect 111 1542 115 1546
rect 135 1542 139 1546
rect 175 1542 179 1546
rect 231 1542 235 1546
rect 303 1542 307 1546
rect 311 1542 315 1546
rect 375 1542 379 1546
rect 391 1542 395 1546
rect 455 1542 459 1546
rect 479 1542 483 1546
rect 527 1542 531 1546
rect 567 1542 571 1546
rect 1047 1646 1051 1650
rect 1095 1646 1099 1650
rect 1455 1730 1459 1734
rect 1463 1730 1467 1734
rect 1527 1730 1531 1734
rect 1599 1730 1603 1734
rect 1607 1730 1611 1734
rect 1671 1730 1675 1734
rect 1687 1730 1691 1734
rect 1751 1782 1755 1786
rect 1767 1782 1771 1786
rect 1847 1782 1851 1786
rect 1855 1782 1859 1786
rect 1927 1782 1931 1786
rect 1967 1782 1971 1786
rect 2007 1782 2011 1786
rect 1743 1730 1747 1734
rect 1767 1730 1771 1734
rect 1295 1674 1299 1678
rect 1303 1674 1307 1678
rect 1343 1674 1347 1678
rect 1391 1674 1395 1678
rect 1399 1674 1403 1678
rect 1447 1674 1451 1678
rect 1463 1674 1467 1678
rect 1503 1674 1507 1678
rect 1527 1674 1531 1678
rect 1567 1674 1571 1678
rect 1599 1674 1603 1678
rect 1807 1730 1811 1734
rect 1847 1730 1851 1734
rect 1879 1730 1883 1734
rect 1927 1730 1931 1734
rect 1951 1730 1955 1734
rect 2007 1730 2011 1734
rect 2119 1834 2123 1838
rect 2071 1782 2075 1786
rect 2119 1782 2123 1786
rect 2023 1730 2027 1734
rect 2071 1730 2075 1734
rect 1631 1674 1635 1678
rect 1671 1674 1675 1678
rect 1695 1674 1699 1678
rect 1743 1674 1747 1678
rect 1759 1674 1763 1678
rect 1807 1674 1811 1678
rect 1831 1674 1835 1678
rect 1879 1674 1883 1678
rect 1911 1674 1915 1678
rect 791 1594 795 1598
rect 815 1594 819 1598
rect 847 1594 851 1598
rect 887 1594 891 1598
rect 903 1594 907 1598
rect 959 1594 963 1598
rect 1007 1594 1011 1598
rect 1047 1594 1051 1598
rect 1095 1594 1099 1598
rect 1135 1610 1139 1614
rect 1159 1610 1163 1614
rect 1215 1610 1219 1614
rect 1263 1610 1267 1614
rect 1303 1610 1307 1614
rect 1343 1610 1347 1614
rect 1383 1610 1387 1614
rect 1391 1610 1395 1614
rect 1447 1610 1451 1614
rect 1463 1610 1467 1614
rect 1503 1610 1507 1614
rect 1543 1610 1547 1614
rect 1567 1610 1571 1614
rect 1623 1610 1627 1614
rect 1631 1610 1635 1614
rect 599 1542 603 1546
rect 655 1542 659 1546
rect 671 1542 675 1546
rect 743 1542 747 1546
rect 815 1542 819 1546
rect 823 1542 827 1546
rect 111 1490 115 1494
rect 135 1490 139 1494
rect 175 1490 179 1494
rect 199 1490 203 1494
rect 231 1490 235 1494
rect 279 1490 283 1494
rect 311 1490 315 1494
rect 359 1490 363 1494
rect 391 1490 395 1494
rect 111 1438 115 1442
rect 135 1438 139 1442
rect 111 1386 115 1390
rect 135 1386 139 1390
rect 191 1438 195 1442
rect 199 1438 203 1442
rect 263 1438 267 1442
rect 279 1438 283 1442
rect 439 1490 443 1494
rect 479 1490 483 1494
rect 519 1490 523 1494
rect 567 1490 571 1494
rect 599 1490 603 1494
rect 655 1490 659 1494
rect 679 1490 683 1494
rect 335 1438 339 1442
rect 359 1438 363 1442
rect 407 1438 411 1442
rect 439 1438 443 1442
rect 175 1386 179 1390
rect 191 1386 195 1390
rect 479 1438 483 1442
rect 519 1438 523 1442
rect 551 1438 555 1442
rect 599 1438 603 1442
rect 631 1438 635 1442
rect 1135 1558 1139 1562
rect 1159 1558 1163 1562
rect 1199 1558 1203 1562
rect 1215 1558 1219 1562
rect 1247 1558 1251 1562
rect 1303 1558 1307 1562
rect 1319 1558 1323 1562
rect 1383 1558 1387 1562
rect 1399 1558 1403 1562
rect 1463 1558 1467 1562
rect 1479 1558 1483 1562
rect 887 1542 891 1546
rect 911 1542 915 1546
rect 999 1542 1003 1546
rect 1095 1542 1099 1546
rect 1951 1674 1955 1678
rect 1999 1674 2003 1678
rect 2023 1674 2027 1678
rect 2119 1730 2123 1734
rect 2071 1674 2075 1678
rect 2119 1674 2123 1678
rect 1695 1610 1699 1614
rect 1711 1610 1715 1614
rect 1543 1558 1547 1562
rect 1559 1558 1563 1562
rect 1759 1610 1763 1614
rect 1799 1610 1803 1614
rect 1831 1610 1835 1614
rect 1887 1610 1891 1614
rect 1911 1610 1915 1614
rect 1983 1610 1987 1614
rect 1999 1610 2003 1614
rect 2071 1610 2075 1614
rect 1623 1558 1627 1562
rect 1647 1558 1651 1562
rect 1711 1558 1715 1562
rect 1735 1558 1739 1562
rect 1799 1558 1803 1562
rect 1823 1558 1827 1562
rect 1887 1558 1891 1562
rect 1911 1558 1915 1562
rect 743 1490 747 1494
rect 767 1490 771 1494
rect 823 1490 827 1494
rect 855 1490 859 1494
rect 911 1490 915 1494
rect 943 1490 947 1494
rect 679 1438 683 1442
rect 711 1438 715 1442
rect 767 1438 771 1442
rect 799 1438 803 1442
rect 1135 1506 1139 1510
rect 1159 1506 1163 1510
rect 999 1490 1003 1494
rect 1031 1490 1035 1494
rect 1095 1490 1099 1494
rect 855 1438 859 1442
rect 887 1438 891 1442
rect 943 1438 947 1442
rect 975 1438 979 1442
rect 1031 1438 1035 1442
rect 1047 1438 1051 1442
rect 239 1386 243 1390
rect 263 1386 267 1390
rect 303 1386 307 1390
rect 335 1386 339 1390
rect 367 1386 371 1390
rect 407 1386 411 1390
rect 439 1386 443 1390
rect 479 1386 483 1390
rect 503 1386 507 1390
rect 111 1326 115 1330
rect 135 1326 139 1330
rect 175 1326 179 1330
rect 215 1326 219 1330
rect 239 1326 243 1330
rect 255 1326 259 1330
rect 303 1326 307 1330
rect 319 1326 323 1330
rect 111 1270 115 1274
rect 135 1270 139 1274
rect 175 1270 179 1274
rect 215 1270 219 1274
rect 255 1270 259 1274
rect 551 1386 555 1390
rect 575 1386 579 1390
rect 631 1386 635 1390
rect 647 1386 651 1390
rect 711 1386 715 1390
rect 783 1386 787 1390
rect 799 1386 803 1390
rect 855 1386 859 1390
rect 887 1386 891 1390
rect 927 1386 931 1390
rect 367 1326 371 1330
rect 391 1326 395 1330
rect 439 1326 443 1330
rect 463 1326 467 1330
rect 503 1326 507 1330
rect 543 1326 547 1330
rect 575 1326 579 1330
rect 623 1326 627 1330
rect 647 1326 651 1330
rect 703 1326 707 1330
rect 711 1326 715 1330
rect 783 1326 787 1330
rect 975 1386 979 1390
rect 999 1386 1003 1390
rect 1199 1506 1203 1510
rect 1239 1506 1243 1510
rect 1247 1506 1251 1510
rect 1303 1506 1307 1510
rect 1319 1506 1323 1510
rect 1375 1506 1379 1510
rect 1399 1506 1403 1510
rect 1455 1506 1459 1510
rect 1479 1506 1483 1510
rect 1543 1506 1547 1510
rect 1559 1506 1563 1510
rect 1623 1506 1627 1510
rect 1647 1506 1651 1510
rect 1703 1506 1707 1510
rect 1735 1506 1739 1510
rect 1775 1506 1779 1510
rect 1823 1506 1827 1510
rect 1847 1506 1851 1510
rect 1911 1506 1915 1510
rect 1919 1506 1923 1510
rect 2119 1610 2123 1614
rect 1983 1558 1987 1562
rect 1999 1558 2003 1562
rect 2071 1558 2075 1562
rect 2119 1558 2123 1562
rect 1991 1506 1995 1510
rect 1999 1506 2003 1510
rect 1135 1450 1139 1454
rect 1159 1450 1163 1454
rect 1199 1450 1203 1454
rect 1239 1450 1243 1454
rect 1279 1450 1283 1454
rect 1303 1450 1307 1454
rect 1327 1450 1331 1454
rect 1375 1450 1379 1454
rect 1383 1450 1387 1454
rect 1439 1450 1443 1454
rect 1455 1450 1459 1454
rect 1495 1450 1499 1454
rect 1095 1438 1099 1442
rect 1543 1450 1547 1454
rect 1551 1450 1555 1454
rect 1607 1450 1611 1454
rect 1623 1450 1627 1454
rect 1671 1450 1675 1454
rect 1703 1450 1707 1454
rect 1735 1450 1739 1454
rect 1775 1450 1779 1454
rect 1807 1450 1811 1454
rect 1847 1450 1851 1454
rect 1887 1450 1891 1454
rect 1135 1394 1139 1398
rect 1279 1394 1283 1398
rect 1327 1394 1331 1398
rect 1335 1394 1339 1398
rect 1375 1394 1379 1398
rect 1383 1394 1387 1398
rect 1415 1394 1419 1398
rect 1439 1394 1443 1398
rect 1455 1394 1459 1398
rect 1495 1394 1499 1398
rect 1535 1394 1539 1398
rect 1551 1394 1555 1398
rect 1583 1394 1587 1398
rect 1607 1394 1611 1398
rect 1647 1394 1651 1398
rect 1671 1394 1675 1398
rect 1719 1394 1723 1398
rect 1735 1394 1739 1398
rect 1047 1386 1051 1390
rect 1095 1386 1099 1390
rect 2063 1506 2067 1510
rect 2071 1506 2075 1510
rect 2119 1506 2123 1510
rect 1919 1450 1923 1454
rect 1975 1450 1979 1454
rect 1991 1450 1995 1454
rect 2063 1450 2067 1454
rect 2119 1450 2123 1454
rect 1807 1394 1811 1398
rect 1887 1394 1891 1398
rect 1895 1394 1899 1398
rect 1975 1394 1979 1398
rect 1991 1394 1995 1398
rect 1135 1342 1139 1346
rect 1159 1342 1163 1346
rect 1223 1342 1227 1346
rect 1311 1342 1315 1346
rect 1335 1342 1339 1346
rect 1375 1342 1379 1346
rect 1407 1342 1411 1346
rect 1415 1342 1419 1346
rect 855 1326 859 1330
rect 863 1326 867 1330
rect 927 1326 931 1330
rect 943 1326 947 1330
rect 999 1326 1003 1330
rect 1023 1326 1027 1330
rect 1047 1326 1051 1330
rect 1095 1326 1099 1330
rect 1455 1342 1459 1346
rect 1495 1342 1499 1346
rect 1503 1342 1507 1346
rect 1535 1342 1539 1346
rect 1583 1342 1587 1346
rect 2063 1394 2067 1398
rect 2071 1394 2075 1398
rect 2119 1394 2123 1398
rect 1599 1342 1603 1346
rect 1647 1342 1651 1346
rect 1679 1342 1683 1346
rect 1719 1342 1723 1346
rect 1759 1342 1763 1346
rect 1807 1342 1811 1346
rect 1831 1342 1835 1346
rect 1895 1342 1899 1346
rect 1959 1342 1963 1346
rect 1991 1342 1995 1346
rect 2023 1342 2027 1346
rect 2071 1342 2075 1346
rect 319 1270 323 1274
rect 391 1270 395 1274
rect 399 1270 403 1274
rect 463 1270 467 1274
rect 487 1270 491 1274
rect 543 1270 547 1274
rect 583 1270 587 1274
rect 623 1270 627 1274
rect 687 1270 691 1274
rect 703 1270 707 1274
rect 783 1270 787 1274
rect 799 1270 803 1274
rect 863 1270 867 1274
rect 919 1270 923 1274
rect 943 1270 947 1274
rect 1023 1270 1027 1274
rect 1047 1270 1051 1274
rect 111 1214 115 1218
rect 135 1214 139 1218
rect 175 1214 179 1218
rect 215 1214 219 1218
rect 255 1214 259 1218
rect 271 1214 275 1218
rect 311 1214 315 1218
rect 319 1214 323 1218
rect 351 1214 355 1218
rect 399 1214 403 1218
rect 447 1214 451 1218
rect 487 1214 491 1218
rect 495 1214 499 1218
rect 551 1214 555 1218
rect 583 1214 587 1218
rect 607 1214 611 1218
rect 671 1214 675 1218
rect 687 1214 691 1218
rect 743 1214 747 1218
rect 799 1214 803 1218
rect 815 1214 819 1218
rect 895 1214 899 1218
rect 919 1214 923 1218
rect 983 1214 987 1218
rect 1135 1290 1139 1294
rect 1159 1290 1163 1294
rect 1175 1290 1179 1294
rect 1223 1290 1227 1294
rect 1231 1290 1235 1294
rect 1303 1290 1307 1294
rect 1311 1290 1315 1294
rect 1095 1270 1099 1274
rect 1199 1256 1203 1260
rect 1391 1290 1395 1294
rect 1407 1290 1411 1294
rect 1479 1290 1483 1294
rect 1503 1290 1507 1294
rect 1567 1290 1571 1294
rect 1599 1290 1603 1294
rect 1655 1290 1659 1294
rect 1679 1290 1683 1294
rect 1743 1290 1747 1294
rect 1759 1290 1763 1294
rect 1135 1234 1139 1238
rect 1175 1234 1179 1238
rect 1231 1234 1235 1238
rect 1287 1234 1291 1238
rect 1303 1234 1307 1238
rect 1047 1214 1051 1218
rect 1095 1214 1099 1218
rect 1327 1234 1331 1238
rect 1375 1234 1379 1238
rect 1391 1234 1395 1238
rect 1591 1256 1595 1260
rect 1431 1234 1435 1238
rect 1479 1234 1483 1238
rect 1495 1234 1499 1238
rect 1559 1234 1563 1238
rect 1567 1234 1571 1238
rect 1623 1234 1627 1238
rect 1655 1234 1659 1238
rect 1831 1290 1835 1294
rect 1895 1290 1899 1294
rect 1919 1290 1923 1294
rect 1959 1290 1963 1294
rect 2007 1290 2011 1294
rect 2023 1290 2027 1294
rect 2119 1342 2123 1346
rect 2071 1290 2075 1294
rect 1679 1234 1683 1238
rect 1735 1234 1739 1238
rect 1743 1234 1747 1238
rect 1791 1234 1795 1238
rect 1831 1234 1835 1238
rect 1847 1234 1851 1238
rect 1903 1234 1907 1238
rect 1919 1234 1923 1238
rect 1967 1234 1971 1238
rect 2119 1290 2123 1294
rect 2007 1234 2011 1238
rect 2031 1234 2035 1238
rect 2071 1234 2075 1238
rect 2119 1234 2123 1238
rect 111 1158 115 1162
rect 271 1158 275 1162
rect 311 1158 315 1162
rect 351 1158 355 1162
rect 399 1158 403 1162
rect 439 1158 443 1162
rect 447 1158 451 1162
rect 479 1158 483 1162
rect 495 1158 499 1162
rect 527 1158 531 1162
rect 551 1158 555 1162
rect 575 1158 579 1162
rect 607 1158 611 1162
rect 623 1158 627 1162
rect 671 1158 675 1162
rect 111 1106 115 1110
rect 159 1106 163 1110
rect 199 1106 203 1110
rect 255 1106 259 1110
rect 319 1106 323 1110
rect 399 1106 403 1110
rect 111 1050 115 1054
rect 135 1050 139 1054
rect 159 1050 163 1054
rect 175 1050 179 1054
rect 439 1106 443 1110
rect 479 1106 483 1110
rect 527 1106 531 1110
rect 559 1106 563 1110
rect 575 1106 579 1110
rect 623 1106 627 1110
rect 639 1106 643 1110
rect 719 1158 723 1162
rect 743 1158 747 1162
rect 775 1158 779 1162
rect 815 1158 819 1162
rect 831 1158 835 1162
rect 887 1158 891 1162
rect 895 1158 899 1162
rect 943 1158 947 1162
rect 1135 1182 1139 1186
rect 1159 1182 1163 1186
rect 1207 1182 1211 1186
rect 1279 1182 1283 1186
rect 1287 1182 1291 1186
rect 1327 1182 1331 1186
rect 1351 1182 1355 1186
rect 1375 1182 1379 1186
rect 1423 1182 1427 1186
rect 1431 1182 1435 1186
rect 1487 1182 1491 1186
rect 1495 1182 1499 1186
rect 983 1158 987 1162
rect 1007 1158 1011 1162
rect 1047 1158 1051 1162
rect 1095 1158 1099 1162
rect 671 1106 675 1110
rect 711 1106 715 1110
rect 719 1106 723 1110
rect 775 1106 779 1110
rect 783 1106 787 1110
rect 831 1106 835 1110
rect 855 1106 859 1110
rect 887 1106 891 1110
rect 927 1106 931 1110
rect 943 1106 947 1110
rect 999 1106 1003 1110
rect 1007 1106 1011 1110
rect 1135 1126 1139 1130
rect 1047 1106 1051 1110
rect 199 1050 203 1054
rect 215 1050 219 1054
rect 255 1050 259 1054
rect 319 1050 323 1054
rect 383 1050 387 1054
rect 399 1050 403 1054
rect 447 1050 451 1054
rect 479 1050 483 1054
rect 511 1050 515 1054
rect 559 1050 563 1054
rect 575 1050 579 1054
rect 111 994 115 998
rect 135 994 139 998
rect 175 994 179 998
rect 215 994 219 998
rect 223 994 227 998
rect 255 994 259 998
rect 279 994 283 998
rect 319 994 323 998
rect 343 994 347 998
rect 383 994 387 998
rect 407 994 411 998
rect 447 994 451 998
rect 471 994 475 998
rect 511 994 515 998
rect 527 994 531 998
rect 631 1050 635 1054
rect 639 1050 643 1054
rect 687 1050 691 1054
rect 711 1050 715 1054
rect 743 1050 747 1054
rect 783 1050 787 1054
rect 799 1050 803 1054
rect 855 1050 859 1054
rect 863 1050 867 1054
rect 575 994 579 998
rect 583 994 587 998
rect 1159 1126 1163 1130
rect 1191 1126 1195 1130
rect 1207 1126 1211 1130
rect 1271 1126 1275 1130
rect 1279 1126 1283 1130
rect 1343 1126 1347 1130
rect 1351 1126 1355 1130
rect 1095 1106 1099 1110
rect 927 1050 931 1054
rect 999 1050 1003 1054
rect 1047 1050 1051 1054
rect 1135 1074 1139 1078
rect 1159 1074 1163 1078
rect 1191 1074 1195 1078
rect 1199 1074 1203 1078
rect 1247 1074 1251 1078
rect 1271 1074 1275 1078
rect 1303 1074 1307 1078
rect 1559 1182 1563 1186
rect 1623 1182 1627 1186
rect 1631 1182 1635 1186
rect 1415 1126 1419 1130
rect 1423 1126 1427 1130
rect 1487 1126 1491 1130
rect 1559 1126 1563 1130
rect 1567 1126 1571 1130
rect 1679 1182 1683 1186
rect 1711 1182 1715 1186
rect 1735 1182 1739 1186
rect 1791 1182 1795 1186
rect 1799 1182 1803 1186
rect 1847 1182 1851 1186
rect 1887 1182 1891 1186
rect 1903 1182 1907 1186
rect 1967 1182 1971 1186
rect 1983 1182 1987 1186
rect 2031 1182 2035 1186
rect 2071 1182 2075 1186
rect 1343 1074 1347 1078
rect 1351 1074 1355 1078
rect 1095 1050 1099 1054
rect 1135 1018 1139 1022
rect 1159 1018 1163 1022
rect 1199 1018 1203 1022
rect 631 994 635 998
rect 687 994 691 998
rect 743 994 747 998
rect 799 994 803 998
rect 863 994 867 998
rect 1095 994 1099 998
rect 1239 1018 1243 1022
rect 1247 1018 1251 1022
rect 1399 1074 1403 1078
rect 1415 1074 1419 1078
rect 1455 1074 1459 1078
rect 1295 1018 1299 1022
rect 1303 1018 1307 1022
rect 1351 1018 1355 1022
rect 1399 1018 1403 1022
rect 1407 1018 1411 1022
rect 111 938 115 942
rect 135 938 139 942
rect 175 938 179 942
rect 223 938 227 942
rect 263 938 267 942
rect 279 938 283 942
rect 303 938 307 942
rect 343 938 347 942
rect 351 938 355 942
rect 399 938 403 942
rect 407 938 411 942
rect 455 938 459 942
rect 471 938 475 942
rect 1135 958 1139 962
rect 1159 958 1163 962
rect 1199 958 1203 962
rect 1207 958 1211 962
rect 511 938 515 942
rect 527 938 531 942
rect 567 938 571 942
rect 583 938 587 942
rect 623 938 627 942
rect 631 938 635 942
rect 687 938 691 942
rect 111 882 115 886
rect 263 882 267 886
rect 303 882 307 886
rect 351 882 355 886
rect 399 882 403 886
rect 415 882 419 886
rect 455 882 459 886
rect 479 882 483 886
rect 511 882 515 886
rect 551 882 555 886
rect 567 882 571 886
rect 623 882 627 886
rect 743 938 747 942
rect 751 938 755 942
rect 799 938 803 942
rect 815 938 819 942
rect 879 938 883 942
rect 943 938 947 942
rect 1007 938 1011 942
rect 1047 938 1051 942
rect 1095 938 1099 942
rect 687 882 691 886
rect 695 882 699 886
rect 751 882 755 886
rect 767 882 771 886
rect 815 882 819 886
rect 831 882 835 886
rect 879 882 883 886
rect 887 882 891 886
rect 943 882 947 886
rect 1239 958 1243 962
rect 1287 958 1291 962
rect 1295 958 1299 962
rect 1351 958 1355 962
rect 1375 958 1379 962
rect 1631 1126 1635 1130
rect 1655 1126 1659 1130
rect 1711 1126 1715 1130
rect 1751 1126 1755 1130
rect 1799 1126 1803 1130
rect 1855 1126 1859 1130
rect 1887 1126 1891 1130
rect 1959 1126 1963 1130
rect 1983 1126 1987 1130
rect 1487 1074 1491 1078
rect 1511 1074 1515 1078
rect 1567 1074 1571 1078
rect 1583 1074 1587 1078
rect 1655 1074 1659 1078
rect 1663 1074 1667 1078
rect 1751 1074 1755 1078
rect 1759 1074 1763 1078
rect 1855 1074 1859 1078
rect 1863 1074 1867 1078
rect 1959 1074 1963 1078
rect 1967 1074 1971 1078
rect 1455 1018 1459 1022
rect 1463 1018 1467 1022
rect 1511 1018 1515 1022
rect 1519 1018 1523 1022
rect 1575 1018 1579 1022
rect 1583 1018 1587 1022
rect 1639 1018 1643 1022
rect 1663 1018 1667 1022
rect 1711 1018 1715 1022
rect 1759 1018 1763 1022
rect 1791 1018 1795 1022
rect 1863 1018 1867 1022
rect 1879 1018 1883 1022
rect 1967 1018 1971 1022
rect 2119 1182 2123 1186
rect 2071 1126 2075 1130
rect 2119 1126 2123 1130
rect 2071 1074 2075 1078
rect 2119 1074 2123 1078
rect 2063 1018 2067 1022
rect 2071 1018 2075 1022
rect 2119 1018 2123 1022
rect 1407 958 1411 962
rect 1455 958 1459 962
rect 1463 958 1467 962
rect 1135 906 1139 910
rect 1007 882 1011 886
rect 1047 882 1051 886
rect 1159 906 1163 910
rect 1207 906 1211 910
rect 1239 906 1243 910
rect 1095 882 1099 886
rect 1519 958 1523 962
rect 1535 958 1539 962
rect 1575 958 1579 962
rect 1615 958 1619 962
rect 1639 958 1643 962
rect 1687 958 1691 962
rect 1711 958 1715 962
rect 1751 958 1755 962
rect 1287 906 1291 910
rect 1319 906 1323 910
rect 1375 906 1379 910
rect 1407 906 1411 910
rect 1455 906 1459 910
rect 1495 906 1499 910
rect 1535 906 1539 910
rect 1583 906 1587 910
rect 111 830 115 834
rect 279 830 283 834
rect 303 830 307 834
rect 343 830 347 834
rect 351 830 355 834
rect 415 830 419 834
rect 479 830 483 834
rect 487 830 491 834
rect 551 830 555 834
rect 567 830 571 834
rect 623 830 627 834
rect 647 830 651 834
rect 695 830 699 834
rect 727 830 731 834
rect 767 830 771 834
rect 111 778 115 782
rect 215 778 219 782
rect 279 778 283 782
rect 343 778 347 782
rect 351 778 355 782
rect 415 778 419 782
rect 423 778 427 782
rect 111 726 115 730
rect 175 726 179 730
rect 487 778 491 782
rect 495 778 499 782
rect 567 778 571 782
rect 639 778 643 782
rect 647 778 651 782
rect 799 830 803 834
rect 831 830 835 834
rect 863 830 867 834
rect 887 830 891 834
rect 927 830 931 834
rect 1135 854 1139 858
rect 1159 854 1163 858
rect 1239 854 1243 858
rect 1247 854 1251 858
rect 1319 854 1323 858
rect 1359 854 1363 858
rect 1791 958 1795 962
rect 1815 958 1819 962
rect 1879 958 1883 962
rect 1951 958 1955 962
rect 1967 958 1971 962
rect 2023 958 2027 962
rect 2063 958 2067 962
rect 2071 958 2075 962
rect 2119 958 2123 962
rect 1615 906 1619 910
rect 1663 906 1667 910
rect 1687 906 1691 910
rect 1743 906 1747 910
rect 1751 906 1755 910
rect 1815 906 1819 910
rect 1879 906 1883 910
rect 1887 906 1891 910
rect 1951 906 1955 910
rect 2023 906 2027 910
rect 1407 854 1411 858
rect 1455 854 1459 858
rect 703 778 707 782
rect 727 778 731 782
rect 759 778 763 782
rect 799 778 803 782
rect 815 778 819 782
rect 863 778 867 782
rect 943 830 947 834
rect 999 830 1003 834
rect 1007 830 1011 834
rect 1047 830 1051 834
rect 1095 830 1099 834
rect 911 778 915 782
rect 927 778 931 782
rect 959 778 963 782
rect 999 778 1003 782
rect 1007 778 1011 782
rect 215 726 219 730
rect 239 726 243 730
rect 279 726 283 730
rect 311 726 315 730
rect 351 726 355 730
rect 391 726 395 730
rect 423 726 427 730
rect 471 726 475 730
rect 495 726 499 730
rect 543 726 547 730
rect 111 674 115 678
rect 135 674 139 678
rect 175 674 179 678
rect 215 674 219 678
rect 239 674 243 678
rect 271 674 275 678
rect 111 614 115 618
rect 135 614 139 618
rect 311 674 315 678
rect 335 674 339 678
rect 391 674 395 678
rect 399 674 403 678
rect 567 726 571 730
rect 615 726 619 730
rect 639 726 643 730
rect 679 726 683 730
rect 703 726 707 730
rect 735 726 739 730
rect 759 726 763 730
rect 799 726 803 730
rect 815 726 819 730
rect 463 674 467 678
rect 471 674 475 678
rect 527 674 531 678
rect 543 674 547 678
rect 591 674 595 678
rect 615 674 619 678
rect 647 674 651 678
rect 679 674 683 678
rect 703 674 707 678
rect 1047 778 1051 782
rect 1135 802 1139 806
rect 1159 802 1163 806
rect 1095 778 1099 782
rect 1247 802 1251 806
rect 1279 802 1283 806
rect 1359 802 1363 806
rect 1407 802 1411 806
rect 1455 802 1459 806
rect 1495 854 1499 858
rect 1543 854 1547 858
rect 1583 854 1587 858
rect 1631 854 1635 858
rect 1663 854 1667 858
rect 1711 854 1715 858
rect 1519 802 1523 806
rect 1543 802 1547 806
rect 1743 854 1747 858
rect 1783 854 1787 858
rect 2071 906 2075 910
rect 2119 906 2123 910
rect 1815 854 1819 858
rect 1855 854 1859 858
rect 1887 854 1891 858
rect 1935 854 1939 858
rect 1951 854 1955 858
rect 2015 854 2019 858
rect 2023 854 2027 858
rect 2071 854 2075 858
rect 1623 802 1627 806
rect 1631 802 1635 806
rect 1711 802 1715 806
rect 1719 802 1723 806
rect 1783 802 1787 806
rect 1815 802 1819 806
rect 1855 802 1859 806
rect 1903 802 1907 806
rect 2119 854 2123 858
rect 1935 802 1939 806
rect 1999 802 2003 806
rect 2015 802 2019 806
rect 2071 802 2075 806
rect 2119 802 2123 806
rect 1135 746 1139 750
rect 1159 746 1163 750
rect 1279 746 1283 750
rect 1335 746 1339 750
rect 1375 746 1379 750
rect 1407 746 1411 750
rect 1415 746 1419 750
rect 1455 746 1459 750
rect 1503 746 1507 750
rect 1519 746 1523 750
rect 1551 746 1555 750
rect 1599 746 1603 750
rect 1623 746 1627 750
rect 1655 746 1659 750
rect 1711 746 1715 750
rect 1719 746 1723 750
rect 1767 746 1771 750
rect 1815 746 1819 750
rect 863 726 867 730
rect 911 726 915 730
rect 927 726 931 730
rect 959 726 963 730
rect 1007 726 1011 730
rect 1047 726 1051 730
rect 1095 726 1099 730
rect 1135 694 1139 698
rect 1247 694 1251 698
rect 1287 694 1291 698
rect 1335 694 1339 698
rect 735 674 739 678
rect 759 674 763 678
rect 799 674 803 678
rect 823 674 827 678
rect 863 674 867 678
rect 927 674 931 678
rect 1095 674 1099 678
rect 1375 694 1379 698
rect 1391 694 1395 698
rect 1415 694 1419 698
rect 1447 694 1451 698
rect 1455 694 1459 698
rect 1503 694 1507 698
rect 1511 694 1515 698
rect 1551 694 1555 698
rect 1583 694 1587 698
rect 1599 694 1603 698
rect 1655 694 1659 698
rect 1831 746 1835 750
rect 1895 746 1899 750
rect 1903 746 1907 750
rect 1959 746 1963 750
rect 1999 746 2003 750
rect 2023 746 2027 750
rect 2071 746 2075 750
rect 1711 694 1715 698
rect 1735 694 1739 698
rect 1767 694 1771 698
rect 1823 694 1827 698
rect 1831 694 1835 698
rect 1895 694 1899 698
rect 1911 694 1915 698
rect 1959 694 1963 698
rect 1999 694 2003 698
rect 2023 694 2027 698
rect 175 614 179 618
rect 215 614 219 618
rect 255 614 259 618
rect 271 614 275 618
rect 303 614 307 618
rect 335 614 339 618
rect 351 614 355 618
rect 399 614 403 618
rect 439 614 443 618
rect 463 614 467 618
rect 487 614 491 618
rect 527 614 531 618
rect 535 614 539 618
rect 583 614 587 618
rect 591 614 595 618
rect 111 558 115 562
rect 135 558 139 562
rect 175 558 179 562
rect 215 558 219 562
rect 223 558 227 562
rect 255 558 259 562
rect 279 558 283 562
rect 303 558 307 562
rect 327 558 331 562
rect 351 558 355 562
rect 375 558 379 562
rect 399 558 403 562
rect 423 558 427 562
rect 439 558 443 562
rect 463 558 467 562
rect 631 614 635 618
rect 647 614 651 618
rect 1135 642 1139 646
rect 1159 642 1163 646
rect 1199 642 1203 646
rect 1239 642 1243 646
rect 1247 642 1251 646
rect 1279 642 1283 646
rect 1287 642 1291 646
rect 679 614 683 618
rect 703 614 707 618
rect 727 614 731 618
rect 759 614 763 618
rect 823 614 827 618
rect 1095 614 1099 618
rect 1135 586 1139 590
rect 1159 586 1163 590
rect 1335 642 1339 646
rect 1343 642 1347 646
rect 1391 642 1395 646
rect 1415 642 1419 646
rect 1447 642 1451 646
rect 1495 642 1499 646
rect 1511 642 1515 646
rect 1583 642 1587 646
rect 1655 642 1659 646
rect 1199 586 1203 590
rect 1239 586 1243 590
rect 1279 586 1283 590
rect 1319 586 1323 590
rect 1343 586 1347 590
rect 1359 586 1363 590
rect 1415 586 1419 590
rect 1487 586 1491 590
rect 1495 586 1499 590
rect 1671 642 1675 646
rect 1735 642 1739 646
rect 1759 642 1763 646
rect 1823 642 1827 646
rect 1839 642 1843 646
rect 1911 642 1915 646
rect 1919 642 1923 646
rect 2119 746 2123 750
rect 2071 694 2075 698
rect 2119 694 2123 698
rect 1999 642 2003 646
rect 2007 642 2011 646
rect 2071 642 2075 646
rect 487 558 491 562
rect 511 558 515 562
rect 535 558 539 562
rect 559 558 563 562
rect 583 558 587 562
rect 607 558 611 562
rect 631 558 635 562
rect 655 558 659 562
rect 679 558 683 562
rect 703 558 707 562
rect 727 558 731 562
rect 751 558 755 562
rect 1095 558 1099 562
rect 1567 586 1571 590
rect 1583 586 1587 590
rect 1655 586 1659 590
rect 1671 586 1675 590
rect 1751 586 1755 590
rect 1759 586 1763 590
rect 1839 586 1843 590
rect 1855 586 1859 590
rect 1919 586 1923 590
rect 1967 586 1971 590
rect 2007 586 2011 590
rect 111 498 115 502
rect 135 498 139 502
rect 175 498 179 502
rect 223 498 227 502
rect 231 498 235 502
rect 279 498 283 502
rect 295 498 299 502
rect 327 498 331 502
rect 359 498 363 502
rect 375 498 379 502
rect 423 498 427 502
rect 463 498 467 502
rect 479 498 483 502
rect 511 498 515 502
rect 535 498 539 502
rect 559 498 563 502
rect 111 442 115 446
rect 135 442 139 446
rect 175 442 179 446
rect 215 442 219 446
rect 231 442 235 446
rect 263 442 267 446
rect 295 442 299 446
rect 327 442 331 446
rect 359 442 363 446
rect 391 442 395 446
rect 423 442 427 446
rect 463 442 467 446
rect 479 442 483 446
rect 535 442 539 446
rect 1135 530 1139 534
rect 1159 530 1163 534
rect 1199 530 1203 534
rect 1239 530 1243 534
rect 1279 530 1283 534
rect 1303 530 1307 534
rect 1319 530 1323 534
rect 1343 530 1347 534
rect 1359 530 1363 534
rect 1383 530 1387 534
rect 1415 530 1419 534
rect 1423 530 1427 534
rect 591 498 595 502
rect 607 498 611 502
rect 639 498 643 502
rect 655 498 659 502
rect 687 498 691 502
rect 703 498 707 502
rect 735 498 739 502
rect 751 498 755 502
rect 791 498 795 502
rect 847 498 851 502
rect 1095 498 1099 502
rect 591 442 595 446
rect 607 442 611 446
rect 639 442 643 446
rect 679 442 683 446
rect 687 442 691 446
rect 735 442 739 446
rect 743 442 747 446
rect 791 442 795 446
rect 807 442 811 446
rect 847 442 851 446
rect 1463 530 1467 534
rect 1487 530 1491 534
rect 1503 530 1507 534
rect 1543 530 1547 534
rect 1567 530 1571 534
rect 1591 530 1595 534
rect 1647 530 1651 534
rect 1655 530 1659 534
rect 1703 530 1707 534
rect 1751 530 1755 534
rect 1767 530 1771 534
rect 1839 530 1843 534
rect 1855 530 1859 534
rect 1919 530 1923 534
rect 2119 642 2123 646
rect 2071 586 2075 590
rect 2119 586 2123 590
rect 1967 530 1971 534
rect 2007 530 2011 534
rect 2071 530 2075 534
rect 2119 530 2123 534
rect 1135 478 1139 482
rect 1295 478 1299 482
rect 1303 478 1307 482
rect 1335 478 1339 482
rect 1343 478 1347 482
rect 1375 478 1379 482
rect 1383 478 1387 482
rect 1423 478 1427 482
rect 1463 478 1467 482
rect 1471 478 1475 482
rect 1503 478 1507 482
rect 1527 478 1531 482
rect 1543 478 1547 482
rect 1583 478 1587 482
rect 1591 478 1595 482
rect 1647 478 1651 482
rect 1703 478 1707 482
rect 1719 478 1723 482
rect 1767 478 1771 482
rect 1807 478 1811 482
rect 1839 478 1843 482
rect 1895 478 1899 482
rect 1919 478 1923 482
rect 1991 478 1995 482
rect 2007 478 2011 482
rect 2071 478 2075 482
rect 871 442 875 446
rect 943 442 947 446
rect 1095 442 1099 446
rect 1135 426 1139 430
rect 1159 426 1163 430
rect 1199 426 1203 430
rect 1255 426 1259 430
rect 1295 426 1299 430
rect 1335 426 1339 430
rect 111 382 115 386
rect 175 382 179 386
rect 215 382 219 386
rect 263 382 267 386
rect 271 382 275 386
rect 327 382 331 386
rect 335 382 339 386
rect 391 382 395 386
rect 407 382 411 386
rect 463 382 467 386
rect 487 382 491 386
rect 535 382 539 386
rect 567 382 571 386
rect 607 382 611 386
rect 639 382 643 386
rect 679 382 683 386
rect 711 382 715 386
rect 743 382 747 386
rect 775 382 779 386
rect 807 382 811 386
rect 839 382 843 386
rect 871 382 875 386
rect 895 382 899 386
rect 667 360 671 364
rect 943 382 947 386
rect 951 382 955 386
rect 1007 382 1011 386
rect 1047 382 1051 386
rect 1095 382 1099 386
rect 915 360 919 364
rect 111 326 115 330
rect 175 326 179 330
rect 215 326 219 330
rect 271 326 275 330
rect 335 326 339 330
rect 383 326 387 330
rect 407 326 411 330
rect 423 326 427 330
rect 463 326 467 330
rect 487 326 491 330
rect 503 326 507 330
rect 543 326 547 330
rect 567 326 571 330
rect 591 326 595 330
rect 639 326 643 330
rect 687 326 691 330
rect 711 326 715 330
rect 735 326 739 330
rect 775 326 779 330
rect 783 326 787 330
rect 831 326 835 330
rect 839 326 843 330
rect 879 326 883 330
rect 895 326 899 330
rect 927 326 931 330
rect 951 326 955 330
rect 967 326 971 330
rect 1007 326 1011 330
rect 1375 426 1379 430
rect 1415 426 1419 430
rect 1423 426 1427 430
rect 1471 426 1475 430
rect 1503 426 1507 430
rect 1527 426 1531 430
rect 1583 426 1587 430
rect 1591 426 1595 430
rect 1135 370 1139 374
rect 1159 370 1163 374
rect 1199 370 1203 374
rect 1047 326 1051 330
rect 111 266 115 270
rect 287 266 291 270
rect 327 266 331 270
rect 367 266 371 270
rect 383 266 387 270
rect 415 266 419 270
rect 423 266 427 270
rect 463 266 467 270
rect 471 266 475 270
rect 503 266 507 270
rect 535 266 539 270
rect 543 266 547 270
rect 591 266 595 270
rect 607 266 611 270
rect 639 266 643 270
rect 679 266 683 270
rect 687 266 691 270
rect 111 202 115 206
rect 167 202 171 206
rect 207 202 211 206
rect 247 202 251 206
rect 287 202 291 206
rect 295 202 299 206
rect 327 202 331 206
rect 111 134 115 138
rect 135 134 139 138
rect 167 134 171 138
rect 175 134 179 138
rect 343 202 347 206
rect 367 202 371 206
rect 399 202 403 206
rect 415 202 419 206
rect 463 202 467 206
rect 471 202 475 206
rect 527 202 531 206
rect 535 202 539 206
rect 599 202 603 206
rect 607 202 611 206
rect 671 202 675 206
rect 679 202 683 206
rect 735 266 739 270
rect 743 266 747 270
rect 783 266 787 270
rect 807 266 811 270
rect 831 266 835 270
rect 863 266 867 270
rect 879 266 883 270
rect 1247 370 1251 374
rect 1255 370 1259 374
rect 1335 370 1339 374
rect 1359 370 1363 374
rect 1415 370 1419 374
rect 1463 370 1467 374
rect 1647 426 1651 430
rect 1671 426 1675 430
rect 1719 426 1723 430
rect 1751 426 1755 430
rect 1807 426 1811 430
rect 1831 426 1835 430
rect 1895 426 1899 430
rect 1911 426 1915 430
rect 1991 426 1995 430
rect 1999 426 2003 430
rect 1503 370 1507 374
rect 1559 370 1563 374
rect 1591 370 1595 374
rect 1647 370 1651 374
rect 1671 370 1675 374
rect 2119 478 2123 482
rect 2071 426 2075 430
rect 1727 370 1731 374
rect 1751 370 1755 374
rect 1799 370 1803 374
rect 1831 370 1835 374
rect 1863 370 1867 374
rect 1911 370 1915 374
rect 1919 370 1923 374
rect 2119 426 2123 430
rect 1975 370 1979 374
rect 1999 370 2003 374
rect 2031 370 2035 374
rect 2071 370 2075 374
rect 2119 370 2123 374
rect 1095 326 1099 330
rect 1135 310 1139 314
rect 1159 310 1163 314
rect 1247 310 1251 314
rect 1351 310 1355 314
rect 1359 310 1363 314
rect 1391 310 1395 314
rect 1431 310 1435 314
rect 1463 310 1467 314
rect 1471 310 1475 314
rect 1511 310 1515 314
rect 1559 310 1563 314
rect 1615 310 1619 314
rect 1647 310 1651 314
rect 1671 310 1675 314
rect 1727 310 1731 314
rect 1735 310 1739 314
rect 1799 310 1803 314
rect 1807 310 1811 314
rect 1863 310 1867 314
rect 1887 310 1891 314
rect 927 266 931 270
rect 967 266 971 270
rect 991 266 995 270
rect 1007 266 1011 270
rect 1047 266 1051 270
rect 1095 266 1099 270
rect 743 202 747 206
rect 751 202 755 206
rect 207 134 211 138
rect 215 134 219 138
rect 247 134 251 138
rect 255 134 259 138
rect 295 134 299 138
rect 335 134 339 138
rect 343 134 347 138
rect 375 134 379 138
rect 399 134 403 138
rect 415 134 419 138
rect 455 134 459 138
rect 463 134 467 138
rect 495 134 499 138
rect 527 134 531 138
rect 535 134 539 138
rect 807 202 811 206
rect 831 202 835 206
rect 863 202 867 206
rect 911 202 915 206
rect 927 202 931 206
rect 991 202 995 206
rect 1047 202 1051 206
rect 1135 258 1139 262
rect 1263 258 1267 262
rect 1303 258 1307 262
rect 1343 258 1347 262
rect 1351 258 1355 262
rect 1919 310 1923 314
rect 1967 310 1971 314
rect 1975 310 1979 314
rect 2031 310 2035 314
rect 2047 310 2051 314
rect 2071 310 2075 314
rect 2119 310 2123 314
rect 1383 258 1387 262
rect 1391 258 1395 262
rect 1423 258 1427 262
rect 1431 258 1435 262
rect 1463 258 1467 262
rect 1471 258 1475 262
rect 1503 258 1507 262
rect 1511 258 1515 262
rect 1543 258 1547 262
rect 1559 258 1563 262
rect 1599 258 1603 262
rect 1615 258 1619 262
rect 1671 258 1675 262
rect 1735 258 1739 262
rect 1759 258 1763 262
rect 1807 258 1811 262
rect 1863 258 1867 262
rect 1887 258 1891 262
rect 1967 258 1971 262
rect 1975 258 1979 262
rect 2047 258 2051 262
rect 2071 258 2075 262
rect 1095 202 1099 206
rect 1135 202 1139 206
rect 1183 202 1187 206
rect 1231 202 1235 206
rect 1263 202 1267 206
rect 1295 202 1299 206
rect 1303 202 1307 206
rect 575 134 579 138
rect 599 134 603 138
rect 615 134 619 138
rect 655 134 659 138
rect 671 134 675 138
rect 695 134 699 138
rect 735 134 739 138
rect 751 134 755 138
rect 775 134 779 138
rect 815 134 819 138
rect 831 134 835 138
rect 871 134 875 138
rect 911 134 915 138
rect 935 134 939 138
rect 991 134 995 138
rect 999 134 1003 138
rect 1047 134 1051 138
rect 1095 134 1099 138
rect 1135 126 1139 130
rect 1159 126 1163 130
rect 1183 126 1187 130
rect 1199 126 1203 130
rect 2119 258 2123 262
rect 1343 202 1347 206
rect 1359 202 1363 206
rect 1383 202 1387 206
rect 1423 202 1427 206
rect 1431 202 1435 206
rect 1463 202 1467 206
rect 1503 202 1507 206
rect 1511 202 1515 206
rect 1543 202 1547 206
rect 1591 202 1595 206
rect 1599 202 1603 206
rect 1663 202 1667 206
rect 1671 202 1675 206
rect 1735 202 1739 206
rect 1759 202 1763 206
rect 1807 202 1811 206
rect 1863 202 1867 206
rect 1879 202 1883 206
rect 1951 202 1955 206
rect 1975 202 1979 206
rect 2023 202 2027 206
rect 1231 126 1235 130
rect 1239 126 1243 130
rect 1279 126 1283 130
rect 1295 126 1299 130
rect 1319 126 1323 130
rect 1359 126 1363 130
rect 1367 126 1371 130
rect 1431 126 1435 130
rect 1495 126 1499 130
rect 1511 126 1515 130
rect 1559 126 1563 130
rect 1591 126 1595 130
rect 1615 126 1619 130
rect 1663 126 1667 130
rect 1671 126 1675 130
rect 1719 126 1723 130
rect 1735 126 1739 130
rect 1767 126 1771 130
rect 1807 126 1811 130
rect 1855 126 1859 130
rect 1879 126 1883 130
rect 1903 126 1907 130
rect 1951 126 1955 130
rect 1991 126 1995 130
rect 2071 202 2075 206
rect 2119 202 2123 206
rect 2023 126 2027 130
rect 2031 126 2035 130
rect 2071 126 2075 130
rect 2119 126 2123 130
rect 111 82 115 86
rect 135 82 139 86
rect 175 82 179 86
rect 215 82 219 86
rect 255 82 259 86
rect 295 82 299 86
rect 335 82 339 86
rect 375 82 379 86
rect 415 82 419 86
rect 455 82 459 86
rect 495 82 499 86
rect 535 82 539 86
rect 575 82 579 86
rect 615 82 619 86
rect 655 82 659 86
rect 695 82 699 86
rect 735 82 739 86
rect 775 82 779 86
rect 815 82 819 86
rect 871 82 875 86
rect 935 82 939 86
rect 999 82 1003 86
rect 1047 82 1051 86
rect 1095 82 1099 86
rect 1135 74 1139 78
rect 1159 74 1163 78
rect 1199 74 1203 78
rect 1239 74 1243 78
rect 1279 74 1283 78
rect 1319 74 1323 78
rect 1367 74 1371 78
rect 1431 74 1435 78
rect 1495 74 1499 78
rect 1559 74 1563 78
rect 1615 74 1619 78
rect 1671 74 1675 78
rect 1719 74 1723 78
rect 1767 74 1771 78
rect 1807 74 1811 78
rect 1855 74 1859 78
rect 1903 74 1907 78
rect 1951 74 1955 78
rect 1991 74 1995 78
rect 2031 74 2035 78
rect 2071 74 2075 78
rect 2119 74 2123 78
<< m4 >>
rect 1118 2209 1119 2215
rect 1125 2214 2155 2215
rect 1125 2210 1135 2214
rect 1139 2210 1343 2214
rect 1347 2210 1383 2214
rect 1387 2210 1423 2214
rect 1427 2210 1463 2214
rect 1467 2210 1503 2214
rect 1507 2210 1543 2214
rect 1547 2210 1583 2214
rect 1587 2210 1623 2214
rect 1627 2210 1663 2214
rect 1667 2210 1703 2214
rect 1707 2210 1743 2214
rect 1747 2210 1783 2214
rect 1787 2210 1823 2214
rect 1827 2210 2119 2214
rect 2123 2210 2155 2214
rect 1125 2209 2155 2210
rect 2161 2209 2162 2215
rect 1106 2157 1107 2163
rect 1113 2162 2143 2163
rect 1113 2158 1135 2162
rect 1139 2158 1287 2162
rect 1291 2158 1327 2162
rect 1331 2158 1343 2162
rect 1347 2158 1367 2162
rect 1371 2158 1383 2162
rect 1387 2158 1415 2162
rect 1419 2158 1423 2162
rect 1427 2158 1463 2162
rect 1467 2158 1503 2162
rect 1507 2158 1519 2162
rect 1523 2158 1543 2162
rect 1547 2158 1575 2162
rect 1579 2158 1583 2162
rect 1587 2158 1623 2162
rect 1627 2158 1663 2162
rect 1667 2158 1671 2162
rect 1675 2158 1703 2162
rect 1707 2158 1719 2162
rect 1723 2158 1743 2162
rect 1747 2158 1775 2162
rect 1779 2158 1783 2162
rect 1787 2158 1823 2162
rect 1827 2158 1831 2162
rect 1835 2158 1887 2162
rect 1891 2158 2119 2162
rect 2123 2158 2143 2162
rect 1113 2157 2143 2158
rect 2149 2157 2150 2163
rect 1314 2116 1320 2117
rect 1606 2116 1612 2117
rect 1314 2112 1315 2116
rect 1319 2112 1607 2116
rect 1611 2112 1612 2116
rect 1314 2111 1320 2112
rect 1606 2111 1612 2112
rect 1118 2101 1119 2107
rect 1125 2106 2155 2107
rect 1125 2102 1135 2106
rect 1139 2102 1223 2106
rect 1227 2102 1279 2106
rect 1283 2102 1287 2106
rect 1291 2102 1327 2106
rect 1331 2102 1343 2106
rect 1347 2102 1367 2106
rect 1371 2102 1415 2106
rect 1419 2102 1423 2106
rect 1427 2102 1463 2106
rect 1467 2102 1503 2106
rect 1507 2102 1519 2106
rect 1523 2102 1575 2106
rect 1579 2102 1583 2106
rect 1587 2102 1623 2106
rect 1627 2102 1663 2106
rect 1667 2102 1671 2106
rect 1675 2102 1719 2106
rect 1723 2102 1743 2106
rect 1747 2102 1775 2106
rect 1779 2102 1831 2106
rect 1835 2102 1887 2106
rect 1891 2102 1919 2106
rect 1923 2102 2007 2106
rect 2011 2102 2071 2106
rect 2075 2102 2119 2106
rect 2123 2102 2155 2106
rect 1125 2101 2155 2102
rect 2161 2101 2162 2107
rect 1106 2049 1107 2055
rect 1113 2054 2143 2055
rect 1113 2050 1135 2054
rect 1139 2050 1183 2054
rect 1187 2050 1223 2054
rect 1227 2050 1239 2054
rect 1243 2050 1279 2054
rect 1283 2050 1311 2054
rect 1315 2050 1343 2054
rect 1347 2050 1399 2054
rect 1403 2050 1423 2054
rect 1427 2050 1487 2054
rect 1491 2050 1503 2054
rect 1507 2050 1583 2054
rect 1587 2050 1663 2054
rect 1667 2050 1671 2054
rect 1675 2050 1743 2054
rect 1747 2050 1759 2054
rect 1763 2050 1831 2054
rect 1835 2050 1839 2054
rect 1843 2050 1919 2054
rect 1923 2050 2007 2054
rect 2011 2050 2071 2054
rect 2075 2050 2119 2054
rect 2123 2050 2143 2054
rect 1113 2049 2143 2050
rect 2149 2049 2150 2055
rect 96 2029 97 2035
rect 103 2034 1119 2035
rect 103 2030 111 2034
rect 115 2030 191 2034
rect 195 2030 231 2034
rect 235 2030 287 2034
rect 291 2030 351 2034
rect 355 2030 423 2034
rect 427 2030 495 2034
rect 499 2030 575 2034
rect 579 2030 647 2034
rect 651 2030 719 2034
rect 723 2030 783 2034
rect 787 2030 839 2034
rect 843 2030 895 2034
rect 899 2030 951 2034
rect 955 2030 1007 2034
rect 1011 2030 1047 2034
rect 1051 2030 1095 2034
rect 1099 2030 1119 2034
rect 103 2029 1119 2030
rect 1125 2029 1126 2035
rect 1118 1997 1119 2003
rect 1125 2002 2155 2003
rect 1125 1998 1135 2002
rect 1139 1998 1183 2002
rect 1187 1998 1239 2002
rect 1243 1998 1303 2002
rect 1307 1998 1311 2002
rect 1315 1998 1383 2002
rect 1387 1998 1399 2002
rect 1403 1998 1463 2002
rect 1467 1998 1487 2002
rect 1491 1998 1543 2002
rect 1547 1998 1583 2002
rect 1587 1998 1615 2002
rect 1619 1998 1671 2002
rect 1675 1998 1687 2002
rect 1691 1998 1751 2002
rect 1755 1998 1759 2002
rect 1763 1998 1815 2002
rect 1819 1998 1839 2002
rect 1843 1998 1879 2002
rect 1883 1998 1919 2002
rect 1923 1998 1951 2002
rect 1955 1998 2007 2002
rect 2011 1998 2023 2002
rect 2027 1998 2071 2002
rect 2075 1998 2119 2002
rect 2123 1998 2155 2002
rect 1125 1997 2155 1998
rect 2161 1997 2162 2003
rect 84 1977 85 1983
rect 91 1982 1107 1983
rect 91 1978 111 1982
rect 115 1978 191 1982
rect 195 1978 231 1982
rect 235 1978 247 1982
rect 251 1978 287 1982
rect 291 1978 311 1982
rect 315 1978 351 1982
rect 355 1978 375 1982
rect 379 1978 423 1982
rect 427 1978 447 1982
rect 451 1978 495 1982
rect 499 1978 519 1982
rect 523 1978 575 1982
rect 579 1978 591 1982
rect 595 1978 647 1982
rect 651 1978 655 1982
rect 659 1978 719 1982
rect 723 1978 775 1982
rect 779 1978 783 1982
rect 787 1978 823 1982
rect 827 1978 839 1982
rect 843 1978 871 1982
rect 875 1978 895 1982
rect 899 1978 919 1982
rect 923 1978 951 1982
rect 955 1978 967 1982
rect 971 1978 1007 1982
rect 1011 1978 1047 1982
rect 1051 1978 1095 1982
rect 1099 1978 1107 1982
rect 91 1977 1107 1978
rect 1113 1977 1114 1983
rect 1642 1980 1648 1981
rect 1974 1980 1980 1981
rect 1642 1976 1643 1980
rect 1647 1976 1975 1980
rect 1979 1976 1980 1980
rect 1642 1975 1648 1976
rect 1974 1975 1980 1976
rect 1106 1941 1107 1947
rect 1113 1946 2143 1947
rect 1113 1942 1135 1946
rect 1139 1942 1159 1946
rect 1163 1942 1223 1946
rect 1227 1942 1303 1946
rect 1307 1942 1383 1946
rect 1387 1942 1463 1946
rect 1467 1942 1535 1946
rect 1539 1942 1543 1946
rect 1547 1942 1615 1946
rect 1619 1942 1687 1946
rect 1691 1942 1695 1946
rect 1699 1942 1751 1946
rect 1755 1942 1783 1946
rect 1787 1942 1815 1946
rect 1819 1942 1879 1946
rect 1883 1942 1951 1946
rect 1955 1942 1983 1946
rect 1987 1942 2023 1946
rect 2027 1942 2071 1946
rect 2075 1942 2119 1946
rect 2123 1942 2143 1946
rect 1113 1941 2143 1942
rect 2149 1941 2150 1947
rect 96 1925 97 1931
rect 103 1930 1119 1931
rect 103 1926 111 1930
rect 115 1926 135 1930
rect 139 1926 175 1930
rect 179 1926 191 1930
rect 195 1926 231 1930
rect 235 1926 247 1930
rect 251 1926 295 1930
rect 299 1926 311 1930
rect 315 1926 367 1930
rect 371 1926 375 1930
rect 379 1926 431 1930
rect 435 1926 447 1930
rect 451 1926 495 1930
rect 499 1926 519 1930
rect 523 1926 559 1930
rect 563 1926 591 1930
rect 595 1926 615 1930
rect 619 1926 655 1930
rect 659 1926 671 1930
rect 675 1926 719 1930
rect 723 1926 727 1930
rect 731 1926 775 1930
rect 779 1926 783 1930
rect 787 1926 823 1930
rect 827 1926 847 1930
rect 851 1926 871 1930
rect 875 1926 919 1930
rect 923 1926 967 1930
rect 971 1926 1007 1930
rect 1011 1926 1047 1930
rect 1051 1926 1095 1930
rect 1099 1926 1119 1930
rect 103 1925 1119 1926
rect 1125 1925 1126 1931
rect 1118 1885 1119 1891
rect 1125 1890 2155 1891
rect 1125 1886 1135 1890
rect 1139 1886 1159 1890
rect 1163 1886 1199 1890
rect 1203 1886 1223 1890
rect 1227 1886 1263 1890
rect 1267 1886 1303 1890
rect 1307 1886 1327 1890
rect 1331 1886 1383 1890
rect 1387 1886 1391 1890
rect 1395 1886 1447 1890
rect 1451 1886 1463 1890
rect 1467 1886 1503 1890
rect 1507 1886 1535 1890
rect 1539 1886 1559 1890
rect 1563 1886 1615 1890
rect 1619 1886 1631 1890
rect 1635 1886 1695 1890
rect 1699 1886 1711 1890
rect 1715 1886 1783 1890
rect 1787 1886 1799 1890
rect 1803 1886 1879 1890
rect 1883 1886 1895 1890
rect 1899 1886 1983 1890
rect 1987 1886 1991 1890
rect 1995 1886 2071 1890
rect 2075 1886 2119 1890
rect 2123 1886 2155 1890
rect 1125 1885 2155 1886
rect 2161 1885 2162 1891
rect 84 1869 85 1875
rect 91 1874 1107 1875
rect 91 1870 111 1874
rect 115 1870 135 1874
rect 139 1870 175 1874
rect 179 1870 199 1874
rect 203 1870 231 1874
rect 235 1870 271 1874
rect 275 1870 295 1874
rect 299 1870 335 1874
rect 339 1870 367 1874
rect 371 1870 399 1874
rect 403 1870 431 1874
rect 435 1870 455 1874
rect 459 1870 495 1874
rect 499 1870 503 1874
rect 507 1870 551 1874
rect 555 1870 559 1874
rect 563 1870 599 1874
rect 603 1870 615 1874
rect 619 1870 647 1874
rect 651 1870 671 1874
rect 675 1870 695 1874
rect 699 1870 727 1874
rect 731 1870 751 1874
rect 755 1870 783 1874
rect 787 1870 847 1874
rect 851 1870 1095 1874
rect 1099 1870 1107 1874
rect 91 1869 1107 1870
rect 1113 1869 1114 1875
rect 1106 1833 1107 1839
rect 1113 1838 2143 1839
rect 1113 1834 1135 1838
rect 1139 1834 1159 1838
rect 1163 1834 1199 1838
rect 1203 1834 1231 1838
rect 1235 1834 1263 1838
rect 1267 1834 1303 1838
rect 1307 1834 1327 1838
rect 1331 1834 1383 1838
rect 1387 1834 1391 1838
rect 1395 1834 1447 1838
rect 1451 1834 1463 1838
rect 1467 1834 1503 1838
rect 1507 1834 1551 1838
rect 1555 1834 1559 1838
rect 1563 1834 1631 1838
rect 1635 1834 1647 1838
rect 1651 1834 1711 1838
rect 1715 1834 1751 1838
rect 1755 1834 1799 1838
rect 1803 1834 1855 1838
rect 1859 1834 1895 1838
rect 1899 1834 1967 1838
rect 1971 1834 1991 1838
rect 1995 1834 2071 1838
rect 2075 1834 2119 1838
rect 2123 1834 2143 1838
rect 1113 1833 2143 1834
rect 2149 1833 2150 1839
rect 96 1809 97 1815
rect 103 1814 1119 1815
rect 103 1810 111 1814
rect 115 1810 135 1814
rect 139 1810 151 1814
rect 155 1810 199 1814
rect 203 1810 215 1814
rect 219 1810 271 1814
rect 275 1810 327 1814
rect 331 1810 335 1814
rect 339 1810 383 1814
rect 387 1810 399 1814
rect 403 1810 431 1814
rect 435 1810 455 1814
rect 459 1810 479 1814
rect 483 1810 503 1814
rect 507 1810 527 1814
rect 531 1810 551 1814
rect 555 1810 575 1814
rect 579 1810 599 1814
rect 603 1810 623 1814
rect 627 1810 647 1814
rect 651 1810 671 1814
rect 675 1810 695 1814
rect 699 1810 727 1814
rect 731 1810 751 1814
rect 755 1810 1095 1814
rect 1099 1810 1119 1814
rect 103 1809 1119 1810
rect 1125 1809 1126 1815
rect 1118 1781 1119 1787
rect 1125 1786 2155 1787
rect 1125 1782 1135 1786
rect 1139 1782 1159 1786
rect 1163 1782 1191 1786
rect 1195 1782 1231 1786
rect 1235 1782 1255 1786
rect 1259 1782 1303 1786
rect 1307 1782 1319 1786
rect 1323 1782 1383 1786
rect 1387 1782 1455 1786
rect 1459 1782 1463 1786
rect 1467 1782 1527 1786
rect 1531 1782 1551 1786
rect 1555 1782 1607 1786
rect 1611 1782 1647 1786
rect 1651 1782 1687 1786
rect 1691 1782 1751 1786
rect 1755 1782 1767 1786
rect 1771 1782 1847 1786
rect 1851 1782 1855 1786
rect 1859 1782 1927 1786
rect 1931 1782 1967 1786
rect 1971 1782 2007 1786
rect 2011 1782 2071 1786
rect 2075 1782 2119 1786
rect 2123 1782 2155 1786
rect 1125 1781 2155 1782
rect 2161 1781 2162 1787
rect 84 1757 85 1763
rect 91 1762 1107 1763
rect 91 1758 111 1762
rect 115 1758 151 1762
rect 155 1758 215 1762
rect 219 1758 231 1762
rect 235 1758 271 1762
rect 275 1758 295 1762
rect 299 1758 327 1762
rect 331 1758 351 1762
rect 355 1758 383 1762
rect 387 1758 415 1762
rect 419 1758 431 1762
rect 435 1758 479 1762
rect 483 1758 527 1762
rect 531 1758 543 1762
rect 547 1758 575 1762
rect 579 1758 615 1762
rect 619 1758 623 1762
rect 627 1758 671 1762
rect 675 1758 687 1762
rect 691 1758 727 1762
rect 731 1758 759 1762
rect 763 1758 831 1762
rect 835 1758 911 1762
rect 915 1758 991 1762
rect 995 1758 1095 1762
rect 1099 1758 1107 1762
rect 91 1757 1107 1758
rect 1113 1757 1114 1763
rect 1106 1729 1107 1735
rect 1113 1734 2143 1735
rect 1113 1730 1135 1734
rect 1139 1730 1191 1734
rect 1195 1730 1247 1734
rect 1251 1730 1255 1734
rect 1259 1730 1295 1734
rect 1299 1730 1319 1734
rect 1323 1730 1343 1734
rect 1347 1730 1383 1734
rect 1387 1730 1399 1734
rect 1403 1730 1455 1734
rect 1459 1730 1463 1734
rect 1467 1730 1527 1734
rect 1531 1730 1599 1734
rect 1603 1730 1607 1734
rect 1611 1730 1671 1734
rect 1675 1730 1687 1734
rect 1691 1730 1743 1734
rect 1747 1730 1767 1734
rect 1771 1730 1807 1734
rect 1811 1730 1847 1734
rect 1851 1730 1879 1734
rect 1883 1730 1927 1734
rect 1931 1730 1951 1734
rect 1955 1730 2007 1734
rect 2011 1730 2023 1734
rect 2027 1730 2071 1734
rect 2075 1730 2119 1734
rect 2123 1730 2143 1734
rect 1113 1729 2143 1730
rect 2149 1729 2150 1735
rect 96 1701 97 1707
rect 103 1706 1119 1707
rect 103 1702 111 1706
rect 115 1702 135 1706
rect 139 1702 199 1706
rect 203 1702 231 1706
rect 235 1702 279 1706
rect 283 1702 295 1706
rect 299 1702 351 1706
rect 355 1702 367 1706
rect 371 1702 415 1706
rect 419 1702 463 1706
rect 467 1702 479 1706
rect 483 1702 543 1706
rect 547 1702 551 1706
rect 555 1702 615 1706
rect 619 1702 639 1706
rect 643 1702 687 1706
rect 691 1702 719 1706
rect 723 1702 759 1706
rect 763 1702 791 1706
rect 795 1702 831 1706
rect 835 1702 855 1706
rect 859 1702 911 1706
rect 915 1702 919 1706
rect 923 1702 983 1706
rect 987 1702 991 1706
rect 995 1702 1047 1706
rect 1051 1702 1095 1706
rect 1099 1702 1119 1706
rect 103 1701 1119 1702
rect 1125 1701 1126 1707
rect 1118 1673 1119 1679
rect 1125 1678 2155 1679
rect 1125 1674 1135 1678
rect 1139 1674 1247 1678
rect 1251 1674 1263 1678
rect 1267 1674 1295 1678
rect 1299 1674 1303 1678
rect 1307 1674 1343 1678
rect 1347 1674 1391 1678
rect 1395 1674 1399 1678
rect 1403 1674 1447 1678
rect 1451 1674 1463 1678
rect 1467 1674 1503 1678
rect 1507 1674 1527 1678
rect 1531 1674 1567 1678
rect 1571 1674 1599 1678
rect 1603 1674 1631 1678
rect 1635 1674 1671 1678
rect 1675 1674 1695 1678
rect 1699 1674 1743 1678
rect 1747 1674 1759 1678
rect 1763 1674 1807 1678
rect 1811 1674 1831 1678
rect 1835 1674 1879 1678
rect 1883 1674 1911 1678
rect 1915 1674 1951 1678
rect 1955 1674 1999 1678
rect 2003 1674 2023 1678
rect 2027 1674 2071 1678
rect 2075 1674 2119 1678
rect 2123 1674 2155 1678
rect 1125 1673 2155 1674
rect 2161 1673 2162 1679
rect 84 1645 85 1651
rect 91 1650 1107 1651
rect 91 1646 111 1650
rect 115 1646 135 1650
rect 139 1646 183 1650
rect 187 1646 199 1650
rect 203 1646 263 1650
rect 267 1646 279 1650
rect 283 1646 343 1650
rect 347 1646 367 1650
rect 371 1646 423 1650
rect 427 1646 463 1650
rect 467 1646 503 1650
rect 507 1646 551 1650
rect 555 1646 583 1650
rect 587 1646 639 1650
rect 643 1646 655 1650
rect 659 1646 719 1650
rect 723 1646 727 1650
rect 731 1646 791 1650
rect 795 1646 847 1650
rect 851 1646 855 1650
rect 859 1646 903 1650
rect 907 1646 919 1650
rect 923 1646 959 1650
rect 963 1646 983 1650
rect 987 1646 1007 1650
rect 1011 1646 1047 1650
rect 1051 1646 1095 1650
rect 1099 1646 1107 1650
rect 91 1645 1107 1646
rect 1113 1645 1114 1651
rect 1106 1609 1107 1615
rect 1113 1614 2143 1615
rect 1113 1610 1135 1614
rect 1139 1610 1159 1614
rect 1163 1610 1215 1614
rect 1219 1610 1263 1614
rect 1267 1610 1303 1614
rect 1307 1610 1343 1614
rect 1347 1610 1383 1614
rect 1387 1610 1391 1614
rect 1395 1610 1447 1614
rect 1451 1610 1463 1614
rect 1467 1610 1503 1614
rect 1507 1610 1543 1614
rect 1547 1610 1567 1614
rect 1571 1610 1623 1614
rect 1627 1610 1631 1614
rect 1635 1610 1695 1614
rect 1699 1610 1711 1614
rect 1715 1610 1759 1614
rect 1763 1610 1799 1614
rect 1803 1610 1831 1614
rect 1835 1610 1887 1614
rect 1891 1610 1911 1614
rect 1915 1610 1983 1614
rect 1987 1610 1999 1614
rect 2003 1610 2071 1614
rect 2075 1610 2119 1614
rect 2123 1610 2143 1614
rect 1113 1609 2143 1610
rect 2149 1609 2150 1615
rect 96 1593 97 1599
rect 103 1598 1119 1599
rect 103 1594 111 1598
rect 115 1594 135 1598
rect 139 1594 175 1598
rect 179 1594 183 1598
rect 187 1594 231 1598
rect 235 1594 263 1598
rect 267 1594 303 1598
rect 307 1594 343 1598
rect 347 1594 375 1598
rect 379 1594 423 1598
rect 427 1594 455 1598
rect 459 1594 503 1598
rect 507 1594 527 1598
rect 531 1594 583 1598
rect 587 1594 599 1598
rect 603 1594 655 1598
rect 659 1594 671 1598
rect 675 1594 727 1598
rect 731 1594 743 1598
rect 747 1594 791 1598
rect 795 1594 815 1598
rect 819 1594 847 1598
rect 851 1594 887 1598
rect 891 1594 903 1598
rect 907 1594 959 1598
rect 963 1594 1007 1598
rect 1011 1594 1047 1598
rect 1051 1594 1095 1598
rect 1099 1594 1119 1598
rect 103 1593 1119 1594
rect 1125 1593 1126 1599
rect 1118 1557 1119 1563
rect 1125 1562 2155 1563
rect 1125 1558 1135 1562
rect 1139 1558 1159 1562
rect 1163 1558 1199 1562
rect 1203 1558 1215 1562
rect 1219 1558 1247 1562
rect 1251 1558 1303 1562
rect 1307 1558 1319 1562
rect 1323 1558 1383 1562
rect 1387 1558 1399 1562
rect 1403 1558 1463 1562
rect 1467 1558 1479 1562
rect 1483 1558 1543 1562
rect 1547 1558 1559 1562
rect 1563 1558 1623 1562
rect 1627 1558 1647 1562
rect 1651 1558 1711 1562
rect 1715 1558 1735 1562
rect 1739 1558 1799 1562
rect 1803 1558 1823 1562
rect 1827 1558 1887 1562
rect 1891 1558 1911 1562
rect 1915 1558 1983 1562
rect 1987 1558 1999 1562
rect 2003 1558 2071 1562
rect 2075 1558 2119 1562
rect 2123 1558 2155 1562
rect 1125 1557 2155 1558
rect 2161 1557 2162 1563
rect 84 1541 85 1547
rect 91 1546 1107 1547
rect 91 1542 111 1546
rect 115 1542 135 1546
rect 139 1542 175 1546
rect 179 1542 231 1546
rect 235 1542 303 1546
rect 307 1542 311 1546
rect 315 1542 375 1546
rect 379 1542 391 1546
rect 395 1542 455 1546
rect 459 1542 479 1546
rect 483 1542 527 1546
rect 531 1542 567 1546
rect 571 1542 599 1546
rect 603 1542 655 1546
rect 659 1542 671 1546
rect 675 1542 743 1546
rect 747 1542 815 1546
rect 819 1542 823 1546
rect 827 1542 887 1546
rect 891 1542 911 1546
rect 915 1542 999 1546
rect 1003 1542 1095 1546
rect 1099 1542 1107 1546
rect 91 1541 1107 1542
rect 1113 1541 1114 1547
rect 1106 1505 1107 1511
rect 1113 1510 2143 1511
rect 1113 1506 1135 1510
rect 1139 1506 1159 1510
rect 1163 1506 1199 1510
rect 1203 1506 1239 1510
rect 1243 1506 1247 1510
rect 1251 1506 1303 1510
rect 1307 1506 1319 1510
rect 1323 1506 1375 1510
rect 1379 1506 1399 1510
rect 1403 1506 1455 1510
rect 1459 1506 1479 1510
rect 1483 1506 1543 1510
rect 1547 1506 1559 1510
rect 1563 1506 1623 1510
rect 1627 1506 1647 1510
rect 1651 1506 1703 1510
rect 1707 1506 1735 1510
rect 1739 1506 1775 1510
rect 1779 1506 1823 1510
rect 1827 1506 1847 1510
rect 1851 1506 1911 1510
rect 1915 1506 1919 1510
rect 1923 1506 1991 1510
rect 1995 1506 1999 1510
rect 2003 1506 2063 1510
rect 2067 1506 2071 1510
rect 2075 1506 2119 1510
rect 2123 1506 2143 1510
rect 1113 1505 2143 1506
rect 2149 1505 2150 1511
rect 96 1489 97 1495
rect 103 1494 1119 1495
rect 103 1490 111 1494
rect 115 1490 135 1494
rect 139 1490 175 1494
rect 179 1490 199 1494
rect 203 1490 231 1494
rect 235 1490 279 1494
rect 283 1490 311 1494
rect 315 1490 359 1494
rect 363 1490 391 1494
rect 395 1490 439 1494
rect 443 1490 479 1494
rect 483 1490 519 1494
rect 523 1490 567 1494
rect 571 1490 599 1494
rect 603 1490 655 1494
rect 659 1490 679 1494
rect 683 1490 743 1494
rect 747 1490 767 1494
rect 771 1490 823 1494
rect 827 1490 855 1494
rect 859 1490 911 1494
rect 915 1490 943 1494
rect 947 1490 999 1494
rect 1003 1490 1031 1494
rect 1035 1490 1095 1494
rect 1099 1490 1119 1494
rect 103 1489 1119 1490
rect 1125 1489 1126 1495
rect 1118 1449 1119 1455
rect 1125 1454 2155 1455
rect 1125 1450 1135 1454
rect 1139 1450 1159 1454
rect 1163 1450 1199 1454
rect 1203 1450 1239 1454
rect 1243 1450 1279 1454
rect 1283 1450 1303 1454
rect 1307 1450 1327 1454
rect 1331 1450 1375 1454
rect 1379 1450 1383 1454
rect 1387 1450 1439 1454
rect 1443 1450 1455 1454
rect 1459 1450 1495 1454
rect 1499 1450 1543 1454
rect 1547 1450 1551 1454
rect 1555 1450 1607 1454
rect 1611 1450 1623 1454
rect 1627 1450 1671 1454
rect 1675 1450 1703 1454
rect 1707 1450 1735 1454
rect 1739 1450 1775 1454
rect 1779 1450 1807 1454
rect 1811 1450 1847 1454
rect 1851 1450 1887 1454
rect 1891 1450 1919 1454
rect 1923 1450 1975 1454
rect 1979 1450 1991 1454
rect 1995 1450 2063 1454
rect 2067 1450 2119 1454
rect 2123 1450 2155 1454
rect 1125 1449 2155 1450
rect 2161 1449 2162 1455
rect 84 1437 85 1443
rect 91 1442 1107 1443
rect 91 1438 111 1442
rect 115 1438 135 1442
rect 139 1438 191 1442
rect 195 1438 199 1442
rect 203 1438 263 1442
rect 267 1438 279 1442
rect 283 1438 335 1442
rect 339 1438 359 1442
rect 363 1438 407 1442
rect 411 1438 439 1442
rect 443 1438 479 1442
rect 483 1438 519 1442
rect 523 1438 551 1442
rect 555 1438 599 1442
rect 603 1438 631 1442
rect 635 1438 679 1442
rect 683 1438 711 1442
rect 715 1438 767 1442
rect 771 1438 799 1442
rect 803 1438 855 1442
rect 859 1438 887 1442
rect 891 1438 943 1442
rect 947 1438 975 1442
rect 979 1438 1031 1442
rect 1035 1438 1047 1442
rect 1051 1438 1095 1442
rect 1099 1438 1107 1442
rect 91 1437 1107 1438
rect 1113 1437 1114 1443
rect 1106 1395 1107 1401
rect 1113 1399 1138 1401
rect 1113 1398 2143 1399
rect 1113 1395 1135 1398
rect 1132 1394 1135 1395
rect 1139 1394 1279 1398
rect 1283 1394 1327 1398
rect 1331 1394 1335 1398
rect 1339 1394 1375 1398
rect 1379 1394 1383 1398
rect 1387 1394 1415 1398
rect 1419 1394 1439 1398
rect 1443 1394 1455 1398
rect 1459 1394 1495 1398
rect 1499 1394 1535 1398
rect 1539 1394 1551 1398
rect 1555 1394 1583 1398
rect 1587 1394 1607 1398
rect 1611 1394 1647 1398
rect 1651 1394 1671 1398
rect 1675 1394 1719 1398
rect 1723 1394 1735 1398
rect 1739 1394 1807 1398
rect 1811 1394 1887 1398
rect 1891 1394 1895 1398
rect 1899 1394 1975 1398
rect 1979 1394 1991 1398
rect 1995 1394 2063 1398
rect 2067 1394 2071 1398
rect 2075 1394 2119 1398
rect 2123 1394 2143 1398
rect 1132 1393 2143 1394
rect 2149 1393 2150 1399
rect 96 1385 97 1391
rect 103 1390 1119 1391
rect 103 1386 111 1390
rect 115 1386 135 1390
rect 139 1386 175 1390
rect 179 1386 191 1390
rect 195 1386 239 1390
rect 243 1386 263 1390
rect 267 1386 303 1390
rect 307 1386 335 1390
rect 339 1386 367 1390
rect 371 1386 407 1390
rect 411 1386 439 1390
rect 443 1386 479 1390
rect 483 1386 503 1390
rect 507 1386 551 1390
rect 555 1386 575 1390
rect 579 1386 631 1390
rect 635 1386 647 1390
rect 651 1386 711 1390
rect 715 1386 783 1390
rect 787 1386 799 1390
rect 803 1386 855 1390
rect 859 1386 887 1390
rect 891 1386 927 1390
rect 931 1386 975 1390
rect 979 1386 999 1390
rect 1003 1386 1047 1390
rect 1051 1386 1095 1390
rect 1099 1386 1119 1390
rect 103 1385 1119 1386
rect 1125 1385 1126 1391
rect 1118 1341 1119 1347
rect 1125 1346 2155 1347
rect 1125 1342 1135 1346
rect 1139 1342 1159 1346
rect 1163 1342 1223 1346
rect 1227 1342 1311 1346
rect 1315 1342 1335 1346
rect 1339 1342 1375 1346
rect 1379 1342 1407 1346
rect 1411 1342 1415 1346
rect 1419 1342 1455 1346
rect 1459 1342 1495 1346
rect 1499 1342 1503 1346
rect 1507 1342 1535 1346
rect 1539 1342 1583 1346
rect 1587 1342 1599 1346
rect 1603 1342 1647 1346
rect 1651 1342 1679 1346
rect 1683 1342 1719 1346
rect 1723 1342 1759 1346
rect 1763 1342 1807 1346
rect 1811 1342 1831 1346
rect 1835 1342 1895 1346
rect 1899 1342 1959 1346
rect 1963 1342 1991 1346
rect 1995 1342 2023 1346
rect 2027 1342 2071 1346
rect 2075 1342 2119 1346
rect 2123 1342 2155 1346
rect 1125 1341 2155 1342
rect 2161 1341 2162 1347
rect 84 1325 85 1331
rect 91 1330 1107 1331
rect 91 1326 111 1330
rect 115 1326 135 1330
rect 139 1326 175 1330
rect 179 1326 215 1330
rect 219 1326 239 1330
rect 243 1326 255 1330
rect 259 1326 303 1330
rect 307 1326 319 1330
rect 323 1326 367 1330
rect 371 1326 391 1330
rect 395 1326 439 1330
rect 443 1326 463 1330
rect 467 1326 503 1330
rect 507 1326 543 1330
rect 547 1326 575 1330
rect 579 1326 623 1330
rect 627 1326 647 1330
rect 651 1326 703 1330
rect 707 1326 711 1330
rect 715 1326 783 1330
rect 787 1326 855 1330
rect 859 1326 863 1330
rect 867 1326 927 1330
rect 931 1326 943 1330
rect 947 1326 999 1330
rect 1003 1326 1023 1330
rect 1027 1326 1047 1330
rect 1051 1326 1095 1330
rect 1099 1326 1107 1330
rect 91 1325 1107 1326
rect 1113 1325 1114 1331
rect 1106 1289 1107 1295
rect 1113 1294 2143 1295
rect 1113 1290 1135 1294
rect 1139 1290 1159 1294
rect 1163 1290 1175 1294
rect 1179 1290 1223 1294
rect 1227 1290 1231 1294
rect 1235 1290 1303 1294
rect 1307 1290 1311 1294
rect 1315 1290 1391 1294
rect 1395 1290 1407 1294
rect 1411 1290 1479 1294
rect 1483 1290 1503 1294
rect 1507 1290 1567 1294
rect 1571 1290 1599 1294
rect 1603 1290 1655 1294
rect 1659 1290 1679 1294
rect 1683 1290 1743 1294
rect 1747 1290 1759 1294
rect 1763 1290 1831 1294
rect 1835 1290 1895 1294
rect 1899 1290 1919 1294
rect 1923 1290 1959 1294
rect 1963 1290 2007 1294
rect 2011 1290 2023 1294
rect 2027 1290 2071 1294
rect 2075 1290 2119 1294
rect 2123 1290 2143 1294
rect 1113 1289 2143 1290
rect 2149 1289 2150 1295
rect 96 1269 97 1275
rect 103 1274 1119 1275
rect 103 1270 111 1274
rect 115 1270 135 1274
rect 139 1270 175 1274
rect 179 1270 215 1274
rect 219 1270 255 1274
rect 259 1270 319 1274
rect 323 1270 391 1274
rect 395 1270 399 1274
rect 403 1270 463 1274
rect 467 1270 487 1274
rect 491 1270 543 1274
rect 547 1270 583 1274
rect 587 1270 623 1274
rect 627 1270 687 1274
rect 691 1270 703 1274
rect 707 1270 783 1274
rect 787 1270 799 1274
rect 803 1270 863 1274
rect 867 1270 919 1274
rect 923 1270 943 1274
rect 947 1270 1023 1274
rect 1027 1270 1047 1274
rect 1051 1270 1095 1274
rect 1099 1270 1119 1274
rect 103 1269 1119 1270
rect 1125 1269 1126 1275
rect 1198 1260 1204 1261
rect 1590 1260 1596 1261
rect 1198 1256 1199 1260
rect 1203 1256 1591 1260
rect 1595 1256 1596 1260
rect 1198 1255 1204 1256
rect 1590 1255 1596 1256
rect 1118 1233 1119 1239
rect 1125 1238 2155 1239
rect 1125 1234 1135 1238
rect 1139 1234 1175 1238
rect 1179 1234 1231 1238
rect 1235 1234 1287 1238
rect 1291 1234 1303 1238
rect 1307 1234 1327 1238
rect 1331 1234 1375 1238
rect 1379 1234 1391 1238
rect 1395 1234 1431 1238
rect 1435 1234 1479 1238
rect 1483 1234 1495 1238
rect 1499 1234 1559 1238
rect 1563 1234 1567 1238
rect 1571 1234 1623 1238
rect 1627 1234 1655 1238
rect 1659 1234 1679 1238
rect 1683 1234 1735 1238
rect 1739 1234 1743 1238
rect 1747 1234 1791 1238
rect 1795 1234 1831 1238
rect 1835 1234 1847 1238
rect 1851 1234 1903 1238
rect 1907 1234 1919 1238
rect 1923 1234 1967 1238
rect 1971 1234 2007 1238
rect 2011 1234 2031 1238
rect 2035 1234 2071 1238
rect 2075 1234 2119 1238
rect 2123 1234 2155 1238
rect 1125 1233 2155 1234
rect 2161 1233 2162 1239
rect 84 1213 85 1219
rect 91 1218 1107 1219
rect 91 1214 111 1218
rect 115 1214 135 1218
rect 139 1214 175 1218
rect 179 1214 215 1218
rect 219 1214 255 1218
rect 259 1214 271 1218
rect 275 1214 311 1218
rect 315 1214 319 1218
rect 323 1214 351 1218
rect 355 1214 399 1218
rect 403 1214 447 1218
rect 451 1214 487 1218
rect 491 1214 495 1218
rect 499 1214 551 1218
rect 555 1214 583 1218
rect 587 1214 607 1218
rect 611 1214 671 1218
rect 675 1214 687 1218
rect 691 1214 743 1218
rect 747 1214 799 1218
rect 803 1214 815 1218
rect 819 1214 895 1218
rect 899 1214 919 1218
rect 923 1214 983 1218
rect 987 1214 1047 1218
rect 1051 1214 1095 1218
rect 1099 1214 1107 1218
rect 91 1213 1107 1214
rect 1113 1213 1114 1219
rect 1106 1181 1107 1187
rect 1113 1186 2143 1187
rect 1113 1182 1135 1186
rect 1139 1182 1159 1186
rect 1163 1182 1207 1186
rect 1211 1182 1279 1186
rect 1283 1182 1287 1186
rect 1291 1182 1327 1186
rect 1331 1182 1351 1186
rect 1355 1182 1375 1186
rect 1379 1182 1423 1186
rect 1427 1182 1431 1186
rect 1435 1182 1487 1186
rect 1491 1182 1495 1186
rect 1499 1182 1559 1186
rect 1563 1182 1623 1186
rect 1627 1182 1631 1186
rect 1635 1182 1679 1186
rect 1683 1182 1711 1186
rect 1715 1182 1735 1186
rect 1739 1182 1791 1186
rect 1795 1182 1799 1186
rect 1803 1182 1847 1186
rect 1851 1182 1887 1186
rect 1891 1182 1903 1186
rect 1907 1182 1967 1186
rect 1971 1182 1983 1186
rect 1987 1182 2031 1186
rect 2035 1182 2071 1186
rect 2075 1182 2119 1186
rect 2123 1182 2143 1186
rect 1113 1181 2143 1182
rect 2149 1181 2150 1187
rect 96 1157 97 1163
rect 103 1162 1119 1163
rect 103 1158 111 1162
rect 115 1158 271 1162
rect 275 1158 311 1162
rect 315 1158 351 1162
rect 355 1158 399 1162
rect 403 1158 439 1162
rect 443 1158 447 1162
rect 451 1158 479 1162
rect 483 1158 495 1162
rect 499 1158 527 1162
rect 531 1158 551 1162
rect 555 1158 575 1162
rect 579 1158 607 1162
rect 611 1158 623 1162
rect 627 1158 671 1162
rect 675 1158 719 1162
rect 723 1158 743 1162
rect 747 1158 775 1162
rect 779 1158 815 1162
rect 819 1158 831 1162
rect 835 1158 887 1162
rect 891 1158 895 1162
rect 899 1158 943 1162
rect 947 1158 983 1162
rect 987 1158 1007 1162
rect 1011 1158 1047 1162
rect 1051 1158 1095 1162
rect 1099 1158 1119 1162
rect 103 1157 1119 1158
rect 1125 1157 1126 1163
rect 1118 1125 1119 1131
rect 1125 1130 2155 1131
rect 1125 1126 1135 1130
rect 1139 1126 1159 1130
rect 1163 1126 1191 1130
rect 1195 1126 1207 1130
rect 1211 1126 1271 1130
rect 1275 1126 1279 1130
rect 1283 1126 1343 1130
rect 1347 1126 1351 1130
rect 1355 1126 1415 1130
rect 1419 1126 1423 1130
rect 1427 1126 1487 1130
rect 1491 1126 1559 1130
rect 1563 1126 1567 1130
rect 1571 1126 1631 1130
rect 1635 1126 1655 1130
rect 1659 1126 1711 1130
rect 1715 1126 1751 1130
rect 1755 1126 1799 1130
rect 1803 1126 1855 1130
rect 1859 1126 1887 1130
rect 1891 1126 1959 1130
rect 1963 1126 1983 1130
rect 1987 1126 2071 1130
rect 2075 1126 2119 1130
rect 2123 1126 2155 1130
rect 1125 1125 2155 1126
rect 2161 1125 2162 1131
rect 84 1105 85 1111
rect 91 1110 1107 1111
rect 91 1106 111 1110
rect 115 1106 159 1110
rect 163 1106 199 1110
rect 203 1106 255 1110
rect 259 1106 319 1110
rect 323 1106 399 1110
rect 403 1106 439 1110
rect 443 1106 479 1110
rect 483 1106 527 1110
rect 531 1106 559 1110
rect 563 1106 575 1110
rect 579 1106 623 1110
rect 627 1106 639 1110
rect 643 1106 671 1110
rect 675 1106 711 1110
rect 715 1106 719 1110
rect 723 1106 775 1110
rect 779 1106 783 1110
rect 787 1106 831 1110
rect 835 1106 855 1110
rect 859 1106 887 1110
rect 891 1106 927 1110
rect 931 1106 943 1110
rect 947 1106 999 1110
rect 1003 1106 1007 1110
rect 1011 1106 1047 1110
rect 1051 1106 1095 1110
rect 1099 1106 1107 1110
rect 91 1105 1107 1106
rect 1113 1105 1114 1111
rect 1106 1073 1107 1079
rect 1113 1078 2143 1079
rect 1113 1074 1135 1078
rect 1139 1074 1159 1078
rect 1163 1074 1191 1078
rect 1195 1074 1199 1078
rect 1203 1074 1247 1078
rect 1251 1074 1271 1078
rect 1275 1074 1303 1078
rect 1307 1074 1343 1078
rect 1347 1074 1351 1078
rect 1355 1074 1399 1078
rect 1403 1074 1415 1078
rect 1419 1074 1455 1078
rect 1459 1074 1487 1078
rect 1491 1074 1511 1078
rect 1515 1074 1567 1078
rect 1571 1074 1583 1078
rect 1587 1074 1655 1078
rect 1659 1074 1663 1078
rect 1667 1074 1751 1078
rect 1755 1074 1759 1078
rect 1763 1074 1855 1078
rect 1859 1074 1863 1078
rect 1867 1074 1959 1078
rect 1963 1074 1967 1078
rect 1971 1074 2071 1078
rect 2075 1074 2119 1078
rect 2123 1074 2143 1078
rect 1113 1073 2143 1074
rect 2149 1073 2150 1079
rect 96 1049 97 1055
rect 103 1054 1119 1055
rect 103 1050 111 1054
rect 115 1050 135 1054
rect 139 1050 159 1054
rect 163 1050 175 1054
rect 179 1050 199 1054
rect 203 1050 215 1054
rect 219 1050 255 1054
rect 259 1050 319 1054
rect 323 1050 383 1054
rect 387 1050 399 1054
rect 403 1050 447 1054
rect 451 1050 479 1054
rect 483 1050 511 1054
rect 515 1050 559 1054
rect 563 1050 575 1054
rect 579 1050 631 1054
rect 635 1050 639 1054
rect 643 1050 687 1054
rect 691 1050 711 1054
rect 715 1050 743 1054
rect 747 1050 783 1054
rect 787 1050 799 1054
rect 803 1050 855 1054
rect 859 1050 863 1054
rect 867 1050 927 1054
rect 931 1050 999 1054
rect 1003 1050 1047 1054
rect 1051 1050 1095 1054
rect 1099 1050 1119 1054
rect 103 1049 1119 1050
rect 1125 1049 1126 1055
rect 1118 1017 1119 1023
rect 1125 1022 2155 1023
rect 1125 1018 1135 1022
rect 1139 1018 1159 1022
rect 1163 1018 1199 1022
rect 1203 1018 1239 1022
rect 1243 1018 1247 1022
rect 1251 1018 1295 1022
rect 1299 1018 1303 1022
rect 1307 1018 1351 1022
rect 1355 1018 1399 1022
rect 1403 1018 1407 1022
rect 1411 1018 1455 1022
rect 1459 1018 1463 1022
rect 1467 1018 1511 1022
rect 1515 1018 1519 1022
rect 1523 1018 1575 1022
rect 1579 1018 1583 1022
rect 1587 1018 1639 1022
rect 1643 1018 1663 1022
rect 1667 1018 1711 1022
rect 1715 1018 1759 1022
rect 1763 1018 1791 1022
rect 1795 1018 1863 1022
rect 1867 1018 1879 1022
rect 1883 1018 1967 1022
rect 1971 1018 2063 1022
rect 2067 1018 2071 1022
rect 2075 1018 2119 1022
rect 2123 1018 2155 1022
rect 1125 1017 2155 1018
rect 2161 1017 2162 1023
rect 84 993 85 999
rect 91 998 1107 999
rect 91 994 111 998
rect 115 994 135 998
rect 139 994 175 998
rect 179 994 215 998
rect 219 994 223 998
rect 227 994 255 998
rect 259 994 279 998
rect 283 994 319 998
rect 323 994 343 998
rect 347 994 383 998
rect 387 994 407 998
rect 411 994 447 998
rect 451 994 471 998
rect 475 994 511 998
rect 515 994 527 998
rect 531 994 575 998
rect 579 994 583 998
rect 587 994 631 998
rect 635 994 687 998
rect 691 994 743 998
rect 747 994 799 998
rect 803 994 863 998
rect 867 994 1095 998
rect 1099 994 1107 998
rect 91 993 1107 994
rect 1113 993 1114 999
rect 1106 957 1107 963
rect 1113 962 2143 963
rect 1113 958 1135 962
rect 1139 958 1159 962
rect 1163 958 1199 962
rect 1203 958 1207 962
rect 1211 958 1239 962
rect 1243 958 1287 962
rect 1291 958 1295 962
rect 1299 958 1351 962
rect 1355 958 1375 962
rect 1379 958 1407 962
rect 1411 958 1455 962
rect 1459 958 1463 962
rect 1467 958 1519 962
rect 1523 958 1535 962
rect 1539 958 1575 962
rect 1579 958 1615 962
rect 1619 958 1639 962
rect 1643 958 1687 962
rect 1691 958 1711 962
rect 1715 958 1751 962
rect 1755 958 1791 962
rect 1795 958 1815 962
rect 1819 958 1879 962
rect 1883 958 1951 962
rect 1955 958 1967 962
rect 1971 958 2023 962
rect 2027 958 2063 962
rect 2067 958 2071 962
rect 2075 958 2119 962
rect 2123 958 2143 962
rect 1113 957 2143 958
rect 2149 957 2150 963
rect 96 937 97 943
rect 103 942 1119 943
rect 103 938 111 942
rect 115 938 135 942
rect 139 938 175 942
rect 179 938 223 942
rect 227 938 263 942
rect 267 938 279 942
rect 283 938 303 942
rect 307 938 343 942
rect 347 938 351 942
rect 355 938 399 942
rect 403 938 407 942
rect 411 938 455 942
rect 459 938 471 942
rect 475 938 511 942
rect 515 938 527 942
rect 531 938 567 942
rect 571 938 583 942
rect 587 938 623 942
rect 627 938 631 942
rect 635 938 687 942
rect 691 938 743 942
rect 747 938 751 942
rect 755 938 799 942
rect 803 938 815 942
rect 819 938 879 942
rect 883 938 943 942
rect 947 938 1007 942
rect 1011 938 1047 942
rect 1051 938 1095 942
rect 1099 938 1119 942
rect 103 937 1119 938
rect 1125 937 1126 943
rect 1118 905 1119 911
rect 1125 910 2155 911
rect 1125 906 1135 910
rect 1139 906 1159 910
rect 1163 906 1207 910
rect 1211 906 1239 910
rect 1243 906 1287 910
rect 1291 906 1319 910
rect 1323 906 1375 910
rect 1379 906 1407 910
rect 1411 906 1455 910
rect 1459 906 1495 910
rect 1499 906 1535 910
rect 1539 906 1583 910
rect 1587 906 1615 910
rect 1619 906 1663 910
rect 1667 906 1687 910
rect 1691 906 1743 910
rect 1747 906 1751 910
rect 1755 906 1815 910
rect 1819 906 1879 910
rect 1883 906 1887 910
rect 1891 906 1951 910
rect 1955 906 2023 910
rect 2027 906 2071 910
rect 2075 906 2119 910
rect 2123 906 2155 910
rect 1125 905 2155 906
rect 2161 905 2162 911
rect 84 881 85 887
rect 91 886 1107 887
rect 91 882 111 886
rect 115 882 263 886
rect 267 882 303 886
rect 307 882 351 886
rect 355 882 399 886
rect 403 882 415 886
rect 419 882 455 886
rect 459 882 479 886
rect 483 882 511 886
rect 515 882 551 886
rect 555 882 567 886
rect 571 882 623 886
rect 627 882 687 886
rect 691 882 695 886
rect 699 882 751 886
rect 755 882 767 886
rect 771 882 815 886
rect 819 882 831 886
rect 835 882 879 886
rect 883 882 887 886
rect 891 882 943 886
rect 947 882 1007 886
rect 1011 882 1047 886
rect 1051 882 1095 886
rect 1099 882 1107 886
rect 91 881 1107 882
rect 1113 881 1114 887
rect 1106 853 1107 859
rect 1113 858 2143 859
rect 1113 854 1135 858
rect 1139 854 1159 858
rect 1163 854 1239 858
rect 1243 854 1247 858
rect 1251 854 1319 858
rect 1323 854 1359 858
rect 1363 854 1407 858
rect 1411 854 1455 858
rect 1459 854 1495 858
rect 1499 854 1543 858
rect 1547 854 1583 858
rect 1587 854 1631 858
rect 1635 854 1663 858
rect 1667 854 1711 858
rect 1715 854 1743 858
rect 1747 854 1783 858
rect 1787 854 1815 858
rect 1819 854 1855 858
rect 1859 854 1887 858
rect 1891 854 1935 858
rect 1939 854 1951 858
rect 1955 854 2015 858
rect 2019 854 2023 858
rect 2027 854 2071 858
rect 2075 854 2119 858
rect 2123 854 2143 858
rect 1113 853 2143 854
rect 2149 853 2150 859
rect 96 829 97 835
rect 103 834 1119 835
rect 103 830 111 834
rect 115 830 279 834
rect 283 830 303 834
rect 307 830 343 834
rect 347 830 351 834
rect 355 830 415 834
rect 419 830 479 834
rect 483 830 487 834
rect 491 830 551 834
rect 555 830 567 834
rect 571 830 623 834
rect 627 830 647 834
rect 651 830 695 834
rect 699 830 727 834
rect 731 830 767 834
rect 771 830 799 834
rect 803 830 831 834
rect 835 830 863 834
rect 867 830 887 834
rect 891 830 927 834
rect 931 830 943 834
rect 947 830 999 834
rect 1003 830 1007 834
rect 1011 830 1047 834
rect 1051 830 1095 834
rect 1099 830 1119 834
rect 103 829 1119 830
rect 1125 829 1126 835
rect 1118 801 1119 807
rect 1125 806 2155 807
rect 1125 802 1135 806
rect 1139 802 1159 806
rect 1163 802 1247 806
rect 1251 802 1279 806
rect 1283 802 1359 806
rect 1363 802 1407 806
rect 1411 802 1455 806
rect 1459 802 1519 806
rect 1523 802 1543 806
rect 1547 802 1623 806
rect 1627 802 1631 806
rect 1635 802 1711 806
rect 1715 802 1719 806
rect 1723 802 1783 806
rect 1787 802 1815 806
rect 1819 802 1855 806
rect 1859 802 1903 806
rect 1907 802 1935 806
rect 1939 802 1999 806
rect 2003 802 2015 806
rect 2019 802 2071 806
rect 2075 802 2119 806
rect 2123 802 2155 806
rect 1125 801 2155 802
rect 2161 801 2162 807
rect 84 777 85 783
rect 91 782 1107 783
rect 91 778 111 782
rect 115 778 215 782
rect 219 778 279 782
rect 283 778 343 782
rect 347 778 351 782
rect 355 778 415 782
rect 419 778 423 782
rect 427 778 487 782
rect 491 778 495 782
rect 499 778 567 782
rect 571 778 639 782
rect 643 778 647 782
rect 651 778 703 782
rect 707 778 727 782
rect 731 778 759 782
rect 763 778 799 782
rect 803 778 815 782
rect 819 778 863 782
rect 867 778 911 782
rect 915 778 927 782
rect 931 778 959 782
rect 963 778 999 782
rect 1003 778 1007 782
rect 1011 778 1047 782
rect 1051 778 1095 782
rect 1099 778 1107 782
rect 91 777 1107 778
rect 1113 777 1114 783
rect 1106 745 1107 751
rect 1113 750 2143 751
rect 1113 746 1135 750
rect 1139 746 1159 750
rect 1163 746 1279 750
rect 1283 746 1335 750
rect 1339 746 1375 750
rect 1379 746 1407 750
rect 1411 746 1415 750
rect 1419 746 1455 750
rect 1459 746 1503 750
rect 1507 746 1519 750
rect 1523 746 1551 750
rect 1555 746 1599 750
rect 1603 746 1623 750
rect 1627 746 1655 750
rect 1659 746 1711 750
rect 1715 746 1719 750
rect 1723 746 1767 750
rect 1771 746 1815 750
rect 1819 746 1831 750
rect 1835 746 1895 750
rect 1899 746 1903 750
rect 1907 746 1959 750
rect 1963 746 1999 750
rect 2003 746 2023 750
rect 2027 746 2071 750
rect 2075 746 2119 750
rect 2123 746 2143 750
rect 1113 745 2143 746
rect 2149 745 2150 751
rect 96 725 97 731
rect 103 730 1119 731
rect 103 726 111 730
rect 115 726 175 730
rect 179 726 215 730
rect 219 726 239 730
rect 243 726 279 730
rect 283 726 311 730
rect 315 726 351 730
rect 355 726 391 730
rect 395 726 423 730
rect 427 726 471 730
rect 475 726 495 730
rect 499 726 543 730
rect 547 726 567 730
rect 571 726 615 730
rect 619 726 639 730
rect 643 726 679 730
rect 683 726 703 730
rect 707 726 735 730
rect 739 726 759 730
rect 763 726 799 730
rect 803 726 815 730
rect 819 726 863 730
rect 867 726 911 730
rect 915 726 927 730
rect 931 726 959 730
rect 963 726 1007 730
rect 1011 726 1047 730
rect 1051 726 1095 730
rect 1099 726 1119 730
rect 103 725 1119 726
rect 1125 725 1126 731
rect 1118 693 1119 699
rect 1125 698 2155 699
rect 1125 694 1135 698
rect 1139 694 1247 698
rect 1251 694 1287 698
rect 1291 694 1335 698
rect 1339 694 1375 698
rect 1379 694 1391 698
rect 1395 694 1415 698
rect 1419 694 1447 698
rect 1451 694 1455 698
rect 1459 694 1503 698
rect 1507 694 1511 698
rect 1515 694 1551 698
rect 1555 694 1583 698
rect 1587 694 1599 698
rect 1603 694 1655 698
rect 1659 694 1711 698
rect 1715 694 1735 698
rect 1739 694 1767 698
rect 1771 694 1823 698
rect 1827 694 1831 698
rect 1835 694 1895 698
rect 1899 694 1911 698
rect 1915 694 1959 698
rect 1963 694 1999 698
rect 2003 694 2023 698
rect 2027 694 2071 698
rect 2075 694 2119 698
rect 2123 694 2155 698
rect 1125 693 2155 694
rect 2161 693 2162 699
rect 84 673 85 679
rect 91 678 1107 679
rect 91 674 111 678
rect 115 674 135 678
rect 139 674 175 678
rect 179 674 215 678
rect 219 674 239 678
rect 243 674 271 678
rect 275 674 311 678
rect 315 674 335 678
rect 339 674 391 678
rect 395 674 399 678
rect 403 674 463 678
rect 467 674 471 678
rect 475 674 527 678
rect 531 674 543 678
rect 547 674 591 678
rect 595 674 615 678
rect 619 674 647 678
rect 651 674 679 678
rect 683 674 703 678
rect 707 674 735 678
rect 739 674 759 678
rect 763 674 799 678
rect 803 674 823 678
rect 827 674 863 678
rect 867 674 927 678
rect 931 674 1095 678
rect 1099 674 1107 678
rect 91 673 1107 674
rect 1113 673 1114 679
rect 1106 641 1107 647
rect 1113 646 2143 647
rect 1113 642 1135 646
rect 1139 642 1159 646
rect 1163 642 1199 646
rect 1203 642 1239 646
rect 1243 642 1247 646
rect 1251 642 1279 646
rect 1283 642 1287 646
rect 1291 642 1335 646
rect 1339 642 1343 646
rect 1347 642 1391 646
rect 1395 642 1415 646
rect 1419 642 1447 646
rect 1451 642 1495 646
rect 1499 642 1511 646
rect 1515 642 1583 646
rect 1587 642 1655 646
rect 1659 642 1671 646
rect 1675 642 1735 646
rect 1739 642 1759 646
rect 1763 642 1823 646
rect 1827 642 1839 646
rect 1843 642 1911 646
rect 1915 642 1919 646
rect 1923 642 1999 646
rect 2003 642 2007 646
rect 2011 642 2071 646
rect 2075 642 2119 646
rect 2123 642 2143 646
rect 1113 641 2143 642
rect 2149 641 2150 647
rect 96 613 97 619
rect 103 618 1119 619
rect 103 614 111 618
rect 115 614 135 618
rect 139 614 175 618
rect 179 614 215 618
rect 219 614 255 618
rect 259 614 271 618
rect 275 614 303 618
rect 307 614 335 618
rect 339 614 351 618
rect 355 614 399 618
rect 403 614 439 618
rect 443 614 463 618
rect 467 614 487 618
rect 491 614 527 618
rect 531 614 535 618
rect 539 614 583 618
rect 587 614 591 618
rect 595 614 631 618
rect 635 614 647 618
rect 651 614 679 618
rect 683 614 703 618
rect 707 614 727 618
rect 731 614 759 618
rect 763 614 823 618
rect 827 614 1095 618
rect 1099 614 1119 618
rect 103 613 1119 614
rect 1125 613 1126 619
rect 1118 585 1119 591
rect 1125 590 2155 591
rect 1125 586 1135 590
rect 1139 586 1159 590
rect 1163 586 1199 590
rect 1203 586 1239 590
rect 1243 586 1279 590
rect 1283 586 1319 590
rect 1323 586 1343 590
rect 1347 586 1359 590
rect 1363 586 1415 590
rect 1419 586 1487 590
rect 1491 586 1495 590
rect 1499 586 1567 590
rect 1571 586 1583 590
rect 1587 586 1655 590
rect 1659 586 1671 590
rect 1675 586 1751 590
rect 1755 586 1759 590
rect 1763 586 1839 590
rect 1843 586 1855 590
rect 1859 586 1919 590
rect 1923 586 1967 590
rect 1971 586 2007 590
rect 2011 586 2071 590
rect 2075 586 2119 590
rect 2123 586 2155 590
rect 1125 585 2155 586
rect 2161 585 2162 591
rect 84 557 85 563
rect 91 562 1107 563
rect 91 558 111 562
rect 115 558 135 562
rect 139 558 175 562
rect 179 558 215 562
rect 219 558 223 562
rect 227 558 255 562
rect 259 558 279 562
rect 283 558 303 562
rect 307 558 327 562
rect 331 558 351 562
rect 355 558 375 562
rect 379 558 399 562
rect 403 558 423 562
rect 427 558 439 562
rect 443 558 463 562
rect 467 558 487 562
rect 491 558 511 562
rect 515 558 535 562
rect 539 558 559 562
rect 563 558 583 562
rect 587 558 607 562
rect 611 558 631 562
rect 635 558 655 562
rect 659 558 679 562
rect 683 558 703 562
rect 707 558 727 562
rect 731 558 751 562
rect 755 558 1095 562
rect 1099 558 1107 562
rect 91 557 1107 558
rect 1113 557 1114 563
rect 1106 529 1107 535
rect 1113 534 2143 535
rect 1113 530 1135 534
rect 1139 530 1159 534
rect 1163 530 1199 534
rect 1203 530 1239 534
rect 1243 530 1279 534
rect 1283 530 1303 534
rect 1307 530 1319 534
rect 1323 530 1343 534
rect 1347 530 1359 534
rect 1363 530 1383 534
rect 1387 530 1415 534
rect 1419 530 1423 534
rect 1427 530 1463 534
rect 1467 530 1487 534
rect 1491 530 1503 534
rect 1507 530 1543 534
rect 1547 530 1567 534
rect 1571 530 1591 534
rect 1595 530 1647 534
rect 1651 530 1655 534
rect 1659 530 1703 534
rect 1707 530 1751 534
rect 1755 530 1767 534
rect 1771 530 1839 534
rect 1843 530 1855 534
rect 1859 530 1919 534
rect 1923 530 1967 534
rect 1971 530 2007 534
rect 2011 530 2071 534
rect 2075 530 2119 534
rect 2123 530 2143 534
rect 1113 529 2143 530
rect 2149 529 2150 535
rect 96 497 97 503
rect 103 502 1119 503
rect 103 498 111 502
rect 115 498 135 502
rect 139 498 175 502
rect 179 498 223 502
rect 227 498 231 502
rect 235 498 279 502
rect 283 498 295 502
rect 299 498 327 502
rect 331 498 359 502
rect 363 498 375 502
rect 379 498 423 502
rect 427 498 463 502
rect 467 498 479 502
rect 483 498 511 502
rect 515 498 535 502
rect 539 498 559 502
rect 563 498 591 502
rect 595 498 607 502
rect 611 498 639 502
rect 643 498 655 502
rect 659 498 687 502
rect 691 498 703 502
rect 707 498 735 502
rect 739 498 751 502
rect 755 498 791 502
rect 795 498 847 502
rect 851 498 1095 502
rect 1099 498 1119 502
rect 103 497 1119 498
rect 1125 497 1126 503
rect 1118 477 1119 483
rect 1125 482 2155 483
rect 1125 478 1135 482
rect 1139 478 1295 482
rect 1299 478 1303 482
rect 1307 478 1335 482
rect 1339 478 1343 482
rect 1347 478 1375 482
rect 1379 478 1383 482
rect 1387 478 1423 482
rect 1427 478 1463 482
rect 1467 478 1471 482
rect 1475 478 1503 482
rect 1507 478 1527 482
rect 1531 478 1543 482
rect 1547 478 1583 482
rect 1587 478 1591 482
rect 1595 478 1647 482
rect 1651 478 1703 482
rect 1707 478 1719 482
rect 1723 478 1767 482
rect 1771 478 1807 482
rect 1811 478 1839 482
rect 1843 478 1895 482
rect 1899 478 1919 482
rect 1923 478 1991 482
rect 1995 478 2007 482
rect 2011 478 2071 482
rect 2075 478 2119 482
rect 2123 478 2155 482
rect 1125 477 2155 478
rect 2161 477 2162 483
rect 84 441 85 447
rect 91 446 1107 447
rect 91 442 111 446
rect 115 442 135 446
rect 139 442 175 446
rect 179 442 215 446
rect 219 442 231 446
rect 235 442 263 446
rect 267 442 295 446
rect 299 442 327 446
rect 331 442 359 446
rect 363 442 391 446
rect 395 442 423 446
rect 427 442 463 446
rect 467 442 479 446
rect 483 442 535 446
rect 539 442 591 446
rect 595 442 607 446
rect 611 442 639 446
rect 643 442 679 446
rect 683 442 687 446
rect 691 442 735 446
rect 739 442 743 446
rect 747 442 791 446
rect 795 442 807 446
rect 811 442 847 446
rect 851 442 871 446
rect 875 442 943 446
rect 947 442 1095 446
rect 1099 442 1107 446
rect 91 441 1107 442
rect 1113 441 1114 447
rect 1106 425 1107 431
rect 1113 430 2143 431
rect 1113 426 1135 430
rect 1139 426 1159 430
rect 1163 426 1199 430
rect 1203 426 1255 430
rect 1259 426 1295 430
rect 1299 426 1335 430
rect 1339 426 1375 430
rect 1379 426 1415 430
rect 1419 426 1423 430
rect 1427 426 1471 430
rect 1475 426 1503 430
rect 1507 426 1527 430
rect 1531 426 1583 430
rect 1587 426 1591 430
rect 1595 426 1647 430
rect 1651 426 1671 430
rect 1675 426 1719 430
rect 1723 426 1751 430
rect 1755 426 1807 430
rect 1811 426 1831 430
rect 1835 426 1895 430
rect 1899 426 1911 430
rect 1915 426 1991 430
rect 1995 426 1999 430
rect 2003 426 2071 430
rect 2075 426 2119 430
rect 2123 426 2143 430
rect 1113 425 2143 426
rect 2149 425 2150 431
rect 96 381 97 387
rect 103 386 1119 387
rect 103 382 111 386
rect 115 382 175 386
rect 179 382 215 386
rect 219 382 263 386
rect 267 382 271 386
rect 275 382 327 386
rect 331 382 335 386
rect 339 382 391 386
rect 395 382 407 386
rect 411 382 463 386
rect 467 382 487 386
rect 491 382 535 386
rect 539 382 567 386
rect 571 382 607 386
rect 611 382 639 386
rect 643 382 679 386
rect 683 382 711 386
rect 715 382 743 386
rect 747 382 775 386
rect 779 382 807 386
rect 811 382 839 386
rect 843 382 871 386
rect 875 382 895 386
rect 899 382 943 386
rect 947 382 951 386
rect 955 382 1007 386
rect 1011 382 1047 386
rect 1051 382 1095 386
rect 1099 382 1119 386
rect 103 381 1119 382
rect 1125 381 1126 387
rect 1118 369 1119 375
rect 1125 374 2155 375
rect 1125 370 1135 374
rect 1139 370 1159 374
rect 1163 370 1199 374
rect 1203 370 1247 374
rect 1251 370 1255 374
rect 1259 370 1335 374
rect 1339 370 1359 374
rect 1363 370 1415 374
rect 1419 370 1463 374
rect 1467 370 1503 374
rect 1507 370 1559 374
rect 1563 370 1591 374
rect 1595 370 1647 374
rect 1651 370 1671 374
rect 1675 370 1727 374
rect 1731 370 1751 374
rect 1755 370 1799 374
rect 1803 370 1831 374
rect 1835 370 1863 374
rect 1867 370 1911 374
rect 1915 370 1919 374
rect 1923 370 1975 374
rect 1979 370 1999 374
rect 2003 370 2031 374
rect 2035 370 2071 374
rect 2075 370 2119 374
rect 2123 370 2155 374
rect 1125 369 2155 370
rect 2161 369 2162 375
rect 666 364 672 365
rect 914 364 920 365
rect 666 360 667 364
rect 671 360 915 364
rect 919 360 920 364
rect 666 359 672 360
rect 914 359 920 360
rect 84 325 85 331
rect 91 330 1107 331
rect 91 326 111 330
rect 115 326 175 330
rect 179 326 215 330
rect 219 326 271 330
rect 275 326 335 330
rect 339 326 383 330
rect 387 326 407 330
rect 411 326 423 330
rect 427 326 463 330
rect 467 326 487 330
rect 491 326 503 330
rect 507 326 543 330
rect 547 326 567 330
rect 571 326 591 330
rect 595 326 639 330
rect 643 326 687 330
rect 691 326 711 330
rect 715 326 735 330
rect 739 326 775 330
rect 779 326 783 330
rect 787 326 831 330
rect 835 326 839 330
rect 843 326 879 330
rect 883 326 895 330
rect 899 326 927 330
rect 931 326 951 330
rect 955 326 967 330
rect 971 326 1007 330
rect 1011 326 1047 330
rect 1051 326 1095 330
rect 1099 326 1107 330
rect 91 325 1107 326
rect 1113 325 1114 331
rect 1106 309 1107 315
rect 1113 314 2143 315
rect 1113 310 1135 314
rect 1139 310 1159 314
rect 1163 310 1247 314
rect 1251 310 1351 314
rect 1355 310 1359 314
rect 1363 310 1391 314
rect 1395 310 1431 314
rect 1435 310 1463 314
rect 1467 310 1471 314
rect 1475 310 1511 314
rect 1515 310 1559 314
rect 1563 310 1615 314
rect 1619 310 1647 314
rect 1651 310 1671 314
rect 1675 310 1727 314
rect 1731 310 1735 314
rect 1739 310 1799 314
rect 1803 310 1807 314
rect 1811 310 1863 314
rect 1867 310 1887 314
rect 1891 310 1919 314
rect 1923 310 1967 314
rect 1971 310 1975 314
rect 1979 310 2031 314
rect 2035 310 2047 314
rect 2051 310 2071 314
rect 2075 310 2119 314
rect 2123 310 2143 314
rect 1113 309 2143 310
rect 2149 309 2150 315
rect 96 265 97 271
rect 103 270 1119 271
rect 103 266 111 270
rect 115 266 287 270
rect 291 266 327 270
rect 331 266 367 270
rect 371 266 383 270
rect 387 266 415 270
rect 419 266 423 270
rect 427 266 463 270
rect 467 266 471 270
rect 475 266 503 270
rect 507 266 535 270
rect 539 266 543 270
rect 547 266 591 270
rect 595 266 607 270
rect 611 266 639 270
rect 643 266 679 270
rect 683 266 687 270
rect 691 266 735 270
rect 739 266 743 270
rect 747 266 783 270
rect 787 266 807 270
rect 811 266 831 270
rect 835 266 863 270
rect 867 266 879 270
rect 883 266 927 270
rect 931 266 967 270
rect 971 266 991 270
rect 995 266 1007 270
rect 1011 266 1047 270
rect 1051 266 1095 270
rect 1099 266 1119 270
rect 103 265 1119 266
rect 1125 265 1126 271
rect 1118 263 1126 265
rect 1118 257 1119 263
rect 1125 262 2155 263
rect 1125 258 1135 262
rect 1139 258 1263 262
rect 1267 258 1303 262
rect 1307 258 1343 262
rect 1347 258 1351 262
rect 1355 258 1383 262
rect 1387 258 1391 262
rect 1395 258 1423 262
rect 1427 258 1431 262
rect 1435 258 1463 262
rect 1467 258 1471 262
rect 1475 258 1503 262
rect 1507 258 1511 262
rect 1515 258 1543 262
rect 1547 258 1559 262
rect 1563 258 1599 262
rect 1603 258 1615 262
rect 1619 258 1671 262
rect 1675 258 1735 262
rect 1739 258 1759 262
rect 1763 258 1807 262
rect 1811 258 1863 262
rect 1867 258 1887 262
rect 1891 258 1967 262
rect 1971 258 1975 262
rect 1979 258 2047 262
rect 2051 258 2071 262
rect 2075 258 2119 262
rect 2123 258 2155 262
rect 1125 257 2155 258
rect 2161 257 2162 263
rect 84 201 85 207
rect 91 206 1107 207
rect 91 202 111 206
rect 115 202 167 206
rect 171 202 207 206
rect 211 202 247 206
rect 251 202 287 206
rect 291 202 295 206
rect 299 202 327 206
rect 331 202 343 206
rect 347 202 367 206
rect 371 202 399 206
rect 403 202 415 206
rect 419 202 463 206
rect 467 202 471 206
rect 475 202 527 206
rect 531 202 535 206
rect 539 202 599 206
rect 603 202 607 206
rect 611 202 671 206
rect 675 202 679 206
rect 683 202 743 206
rect 747 202 751 206
rect 755 202 807 206
rect 811 202 831 206
rect 835 202 863 206
rect 867 202 911 206
rect 915 202 927 206
rect 931 202 991 206
rect 995 202 1047 206
rect 1051 202 1095 206
rect 1099 202 1107 206
rect 91 201 1107 202
rect 1113 206 2150 207
rect 1113 202 1135 206
rect 1139 202 1183 206
rect 1187 202 1231 206
rect 1235 202 1263 206
rect 1267 202 1295 206
rect 1299 202 1303 206
rect 1307 202 1343 206
rect 1347 202 1359 206
rect 1363 202 1383 206
rect 1387 202 1423 206
rect 1427 202 1431 206
rect 1435 202 1463 206
rect 1467 202 1503 206
rect 1507 202 1511 206
rect 1515 202 1543 206
rect 1547 202 1591 206
rect 1595 202 1599 206
rect 1603 202 1663 206
rect 1667 202 1671 206
rect 1675 202 1735 206
rect 1739 202 1759 206
rect 1763 202 1807 206
rect 1811 202 1863 206
rect 1867 202 1879 206
rect 1883 202 1951 206
rect 1955 202 1975 206
rect 1979 202 2023 206
rect 2027 202 2071 206
rect 2075 202 2119 206
rect 2123 202 2150 206
rect 1113 201 2150 202
rect 96 133 97 139
rect 103 138 1119 139
rect 103 134 111 138
rect 115 134 135 138
rect 139 134 167 138
rect 171 134 175 138
rect 179 134 207 138
rect 211 134 215 138
rect 219 134 247 138
rect 251 134 255 138
rect 259 134 295 138
rect 299 134 335 138
rect 339 134 343 138
rect 347 134 375 138
rect 379 134 399 138
rect 403 134 415 138
rect 419 134 455 138
rect 459 134 463 138
rect 467 134 495 138
rect 499 134 527 138
rect 531 134 535 138
rect 539 134 575 138
rect 579 134 599 138
rect 603 134 615 138
rect 619 134 655 138
rect 659 134 671 138
rect 675 134 695 138
rect 699 134 735 138
rect 739 134 751 138
rect 755 134 775 138
rect 779 134 815 138
rect 819 134 831 138
rect 835 134 871 138
rect 875 134 911 138
rect 915 134 935 138
rect 939 134 991 138
rect 995 134 999 138
rect 1003 134 1047 138
rect 1051 134 1095 138
rect 1099 134 1119 138
rect 103 133 1119 134
rect 1125 133 1126 139
rect 1118 131 1126 133
rect 1118 125 1119 131
rect 1125 130 2155 131
rect 1125 126 1135 130
rect 1139 126 1159 130
rect 1163 126 1183 130
rect 1187 126 1199 130
rect 1203 126 1231 130
rect 1235 126 1239 130
rect 1243 126 1279 130
rect 1283 126 1295 130
rect 1299 126 1319 130
rect 1323 126 1359 130
rect 1363 126 1367 130
rect 1371 126 1431 130
rect 1435 126 1495 130
rect 1499 126 1511 130
rect 1515 126 1559 130
rect 1563 126 1591 130
rect 1595 126 1615 130
rect 1619 126 1663 130
rect 1667 126 1671 130
rect 1675 126 1719 130
rect 1723 126 1735 130
rect 1739 126 1767 130
rect 1771 126 1807 130
rect 1811 126 1855 130
rect 1859 126 1879 130
rect 1883 126 1903 130
rect 1907 126 1951 130
rect 1955 126 1991 130
rect 1995 126 2023 130
rect 2027 126 2031 130
rect 2035 126 2071 130
rect 2075 126 2119 130
rect 2123 126 2155 130
rect 1125 125 2155 126
rect 2161 125 2162 131
rect 84 81 85 87
rect 91 86 1107 87
rect 91 82 111 86
rect 115 82 135 86
rect 139 82 175 86
rect 179 82 215 86
rect 219 82 255 86
rect 259 82 295 86
rect 299 82 335 86
rect 339 82 375 86
rect 379 82 415 86
rect 419 82 455 86
rect 459 82 495 86
rect 499 82 535 86
rect 539 82 575 86
rect 579 82 615 86
rect 619 82 655 86
rect 659 82 695 86
rect 699 82 735 86
rect 739 82 775 86
rect 779 82 815 86
rect 819 82 871 86
rect 875 82 935 86
rect 939 82 999 86
rect 1003 82 1047 86
rect 1051 82 1095 86
rect 1099 82 1107 86
rect 91 81 1107 82
rect 1113 81 1114 87
rect 1106 79 1114 81
rect 1106 73 1107 79
rect 1113 78 2143 79
rect 1113 74 1135 78
rect 1139 74 1159 78
rect 1163 74 1199 78
rect 1203 74 1239 78
rect 1243 74 1279 78
rect 1283 74 1319 78
rect 1323 74 1367 78
rect 1371 74 1431 78
rect 1435 74 1495 78
rect 1499 74 1559 78
rect 1563 74 1615 78
rect 1619 74 1671 78
rect 1675 74 1719 78
rect 1723 74 1767 78
rect 1771 74 1807 78
rect 1811 74 1855 78
rect 1859 74 1903 78
rect 1907 74 1951 78
rect 1955 74 1991 78
rect 1995 74 2031 78
rect 2035 74 2071 78
rect 2075 74 2119 78
rect 2123 74 2143 78
rect 1113 73 2143 74
rect 2149 73 2150 79
<< m5c >>
rect 1119 2209 1125 2215
rect 2155 2209 2161 2215
rect 1107 2157 1113 2163
rect 2143 2157 2149 2163
rect 1119 2101 1125 2107
rect 2155 2101 2161 2107
rect 1107 2049 1113 2055
rect 2143 2049 2149 2055
rect 97 2029 103 2035
rect 1119 2029 1125 2035
rect 1119 1997 1125 2003
rect 2155 1997 2161 2003
rect 85 1977 91 1983
rect 1107 1977 1113 1983
rect 1107 1941 1113 1947
rect 2143 1941 2149 1947
rect 97 1925 103 1931
rect 1119 1925 1125 1931
rect 1119 1885 1125 1891
rect 2155 1885 2161 1891
rect 85 1869 91 1875
rect 1107 1869 1113 1875
rect 1107 1833 1113 1839
rect 2143 1833 2149 1839
rect 97 1809 103 1815
rect 1119 1809 1125 1815
rect 1119 1781 1125 1787
rect 2155 1781 2161 1787
rect 85 1757 91 1763
rect 1107 1757 1113 1763
rect 1107 1729 1113 1735
rect 2143 1729 2149 1735
rect 97 1701 103 1707
rect 1119 1701 1125 1707
rect 1119 1673 1125 1679
rect 2155 1673 2161 1679
rect 85 1645 91 1651
rect 1107 1645 1113 1651
rect 1107 1609 1113 1615
rect 2143 1609 2149 1615
rect 97 1593 103 1599
rect 1119 1593 1125 1599
rect 1119 1557 1125 1563
rect 2155 1557 2161 1563
rect 85 1541 91 1547
rect 1107 1541 1113 1547
rect 1107 1505 1113 1511
rect 2143 1505 2149 1511
rect 97 1489 103 1495
rect 1119 1489 1125 1495
rect 1119 1449 1125 1455
rect 2155 1449 2161 1455
rect 85 1437 91 1443
rect 1107 1437 1113 1443
rect 1107 1395 1113 1401
rect 2143 1393 2149 1399
rect 97 1385 103 1391
rect 1119 1385 1125 1391
rect 1119 1341 1125 1347
rect 2155 1341 2161 1347
rect 85 1325 91 1331
rect 1107 1325 1113 1331
rect 1107 1289 1113 1295
rect 2143 1289 2149 1295
rect 97 1269 103 1275
rect 1119 1269 1125 1275
rect 1119 1233 1125 1239
rect 2155 1233 2161 1239
rect 85 1213 91 1219
rect 1107 1213 1113 1219
rect 1107 1181 1113 1187
rect 2143 1181 2149 1187
rect 97 1157 103 1163
rect 1119 1157 1125 1163
rect 1119 1125 1125 1131
rect 2155 1125 2161 1131
rect 85 1105 91 1111
rect 1107 1105 1113 1111
rect 1107 1073 1113 1079
rect 2143 1073 2149 1079
rect 97 1049 103 1055
rect 1119 1049 1125 1055
rect 1119 1017 1125 1023
rect 2155 1017 2161 1023
rect 85 993 91 999
rect 1107 993 1113 999
rect 1107 957 1113 963
rect 2143 957 2149 963
rect 97 937 103 943
rect 1119 937 1125 943
rect 1119 905 1125 911
rect 2155 905 2161 911
rect 85 881 91 887
rect 1107 881 1113 887
rect 1107 853 1113 859
rect 2143 853 2149 859
rect 97 829 103 835
rect 1119 829 1125 835
rect 1119 801 1125 807
rect 2155 801 2161 807
rect 85 777 91 783
rect 1107 777 1113 783
rect 1107 745 1113 751
rect 2143 745 2149 751
rect 97 725 103 731
rect 1119 725 1125 731
rect 1119 693 1125 699
rect 2155 693 2161 699
rect 85 673 91 679
rect 1107 673 1113 679
rect 1107 641 1113 647
rect 2143 641 2149 647
rect 97 613 103 619
rect 1119 613 1125 619
rect 1119 585 1125 591
rect 2155 585 2161 591
rect 85 557 91 563
rect 1107 557 1113 563
rect 1107 529 1113 535
rect 2143 529 2149 535
rect 97 497 103 503
rect 1119 497 1125 503
rect 1119 477 1125 483
rect 2155 477 2161 483
rect 85 441 91 447
rect 1107 441 1113 447
rect 1107 425 1113 431
rect 2143 425 2149 431
rect 97 381 103 387
rect 1119 381 1125 387
rect 1119 369 1125 375
rect 2155 369 2161 375
rect 85 325 91 331
rect 1107 325 1113 331
rect 1107 309 1113 315
rect 2143 309 2149 315
rect 97 265 103 271
rect 1119 265 1125 271
rect 1119 257 1125 263
rect 2155 257 2161 263
rect 85 201 91 207
rect 1107 201 1113 207
rect 97 133 103 139
rect 1119 133 1125 139
rect 1119 125 1125 131
rect 2155 125 2161 131
rect 85 81 91 87
rect 1107 81 1113 87
rect 1107 73 1113 79
rect 2143 73 2149 79
<< m5 >>
rect 84 1983 92 2232
rect 84 1977 85 1983
rect 91 1977 92 1983
rect 84 1875 92 1977
rect 84 1869 85 1875
rect 91 1869 92 1875
rect 84 1763 92 1869
rect 84 1757 85 1763
rect 91 1757 92 1763
rect 84 1651 92 1757
rect 84 1645 85 1651
rect 91 1645 92 1651
rect 84 1547 92 1645
rect 84 1541 85 1547
rect 91 1541 92 1547
rect 84 1443 92 1541
rect 84 1437 85 1443
rect 91 1437 92 1443
rect 84 1331 92 1437
rect 84 1325 85 1331
rect 91 1325 92 1331
rect 84 1219 92 1325
rect 84 1213 85 1219
rect 91 1213 92 1219
rect 84 1111 92 1213
rect 84 1105 85 1111
rect 91 1105 92 1111
rect 84 999 92 1105
rect 84 993 85 999
rect 91 993 92 999
rect 84 887 92 993
rect 84 881 85 887
rect 91 881 92 887
rect 84 783 92 881
rect 84 777 85 783
rect 91 777 92 783
rect 84 679 92 777
rect 84 673 85 679
rect 91 673 92 679
rect 84 563 92 673
rect 84 557 85 563
rect 91 557 92 563
rect 84 447 92 557
rect 84 441 85 447
rect 91 441 92 447
rect 84 331 92 441
rect 84 325 85 331
rect 91 325 92 331
rect 84 207 92 325
rect 84 201 85 207
rect 91 201 92 207
rect 84 87 92 201
rect 84 81 85 87
rect 91 81 92 87
rect 84 72 92 81
rect 96 2035 104 2232
rect 96 2029 97 2035
rect 103 2029 104 2035
rect 96 1931 104 2029
rect 96 1925 97 1931
rect 103 1925 104 1931
rect 96 1815 104 1925
rect 96 1809 97 1815
rect 103 1809 104 1815
rect 96 1707 104 1809
rect 96 1701 97 1707
rect 103 1701 104 1707
rect 96 1599 104 1701
rect 96 1593 97 1599
rect 103 1593 104 1599
rect 96 1495 104 1593
rect 96 1489 97 1495
rect 103 1489 104 1495
rect 96 1391 104 1489
rect 96 1385 97 1391
rect 103 1385 104 1391
rect 96 1275 104 1385
rect 96 1269 97 1275
rect 103 1269 104 1275
rect 96 1163 104 1269
rect 96 1157 97 1163
rect 103 1157 104 1163
rect 96 1055 104 1157
rect 96 1049 97 1055
rect 103 1049 104 1055
rect 96 943 104 1049
rect 96 937 97 943
rect 103 937 104 943
rect 96 835 104 937
rect 96 829 97 835
rect 103 829 104 835
rect 96 731 104 829
rect 96 725 97 731
rect 103 725 104 731
rect 96 619 104 725
rect 96 613 97 619
rect 103 613 104 619
rect 96 503 104 613
rect 96 497 97 503
rect 103 497 104 503
rect 96 387 104 497
rect 96 381 97 387
rect 103 381 104 387
rect 96 271 104 381
rect 96 265 97 271
rect 103 265 104 271
rect 96 139 104 265
rect 96 133 97 139
rect 103 133 104 139
rect 96 72 104 133
rect 1106 2163 1114 2232
rect 1106 2157 1107 2163
rect 1113 2157 1114 2163
rect 1106 2055 1114 2157
rect 1106 2049 1107 2055
rect 1113 2049 1114 2055
rect 1106 1983 1114 2049
rect 1106 1977 1107 1983
rect 1113 1977 1114 1983
rect 1106 1947 1114 1977
rect 1106 1941 1107 1947
rect 1113 1941 1114 1947
rect 1106 1875 1114 1941
rect 1106 1869 1107 1875
rect 1113 1869 1114 1875
rect 1106 1839 1114 1869
rect 1106 1833 1107 1839
rect 1113 1833 1114 1839
rect 1106 1763 1114 1833
rect 1106 1757 1107 1763
rect 1113 1757 1114 1763
rect 1106 1735 1114 1757
rect 1106 1729 1107 1735
rect 1113 1729 1114 1735
rect 1106 1651 1114 1729
rect 1106 1645 1107 1651
rect 1113 1645 1114 1651
rect 1106 1615 1114 1645
rect 1106 1609 1107 1615
rect 1113 1609 1114 1615
rect 1106 1547 1114 1609
rect 1106 1541 1107 1547
rect 1113 1541 1114 1547
rect 1106 1511 1114 1541
rect 1106 1505 1107 1511
rect 1113 1505 1114 1511
rect 1106 1443 1114 1505
rect 1106 1437 1107 1443
rect 1113 1437 1114 1443
rect 1106 1401 1114 1437
rect 1106 1395 1107 1401
rect 1113 1395 1114 1401
rect 1106 1331 1114 1395
rect 1106 1325 1107 1331
rect 1113 1325 1114 1331
rect 1106 1295 1114 1325
rect 1106 1289 1107 1295
rect 1113 1289 1114 1295
rect 1106 1219 1114 1289
rect 1106 1213 1107 1219
rect 1113 1213 1114 1219
rect 1106 1187 1114 1213
rect 1106 1181 1107 1187
rect 1113 1181 1114 1187
rect 1106 1111 1114 1181
rect 1106 1105 1107 1111
rect 1113 1105 1114 1111
rect 1106 1079 1114 1105
rect 1106 1073 1107 1079
rect 1113 1073 1114 1079
rect 1106 999 1114 1073
rect 1106 993 1107 999
rect 1113 993 1114 999
rect 1106 963 1114 993
rect 1106 957 1107 963
rect 1113 957 1114 963
rect 1106 887 1114 957
rect 1106 881 1107 887
rect 1113 881 1114 887
rect 1106 859 1114 881
rect 1106 853 1107 859
rect 1113 853 1114 859
rect 1106 783 1114 853
rect 1106 777 1107 783
rect 1113 777 1114 783
rect 1106 751 1114 777
rect 1106 745 1107 751
rect 1113 745 1114 751
rect 1106 679 1114 745
rect 1106 673 1107 679
rect 1113 673 1114 679
rect 1106 647 1114 673
rect 1106 641 1107 647
rect 1113 641 1114 647
rect 1106 563 1114 641
rect 1106 557 1107 563
rect 1113 557 1114 563
rect 1106 535 1114 557
rect 1106 529 1107 535
rect 1113 529 1114 535
rect 1106 447 1114 529
rect 1106 441 1107 447
rect 1113 441 1114 447
rect 1106 431 1114 441
rect 1106 425 1107 431
rect 1113 425 1114 431
rect 1106 331 1114 425
rect 1106 325 1107 331
rect 1113 325 1114 331
rect 1106 315 1114 325
rect 1106 309 1107 315
rect 1113 309 1114 315
rect 1106 207 1114 309
rect 1106 201 1107 207
rect 1113 201 1114 207
rect 1106 87 1114 201
rect 1106 81 1107 87
rect 1113 81 1114 87
rect 1106 79 1114 81
rect 1106 73 1107 79
rect 1113 73 1114 79
rect 1106 72 1114 73
rect 1118 2215 1126 2232
rect 1118 2209 1119 2215
rect 1125 2209 1126 2215
rect 1118 2107 1126 2209
rect 1118 2101 1119 2107
rect 1125 2101 1126 2107
rect 1118 2035 1126 2101
rect 1118 2029 1119 2035
rect 1125 2029 1126 2035
rect 1118 2003 1126 2029
rect 1118 1997 1119 2003
rect 1125 1997 1126 2003
rect 1118 1931 1126 1997
rect 1118 1925 1119 1931
rect 1125 1925 1126 1931
rect 1118 1891 1126 1925
rect 1118 1885 1119 1891
rect 1125 1885 1126 1891
rect 1118 1815 1126 1885
rect 1118 1809 1119 1815
rect 1125 1809 1126 1815
rect 1118 1787 1126 1809
rect 1118 1781 1119 1787
rect 1125 1781 1126 1787
rect 1118 1707 1126 1781
rect 1118 1701 1119 1707
rect 1125 1701 1126 1707
rect 1118 1679 1126 1701
rect 1118 1673 1119 1679
rect 1125 1673 1126 1679
rect 1118 1599 1126 1673
rect 1118 1593 1119 1599
rect 1125 1593 1126 1599
rect 1118 1563 1126 1593
rect 1118 1557 1119 1563
rect 1125 1557 1126 1563
rect 1118 1495 1126 1557
rect 1118 1489 1119 1495
rect 1125 1489 1126 1495
rect 1118 1455 1126 1489
rect 1118 1449 1119 1455
rect 1125 1449 1126 1455
rect 1118 1391 1126 1449
rect 1118 1385 1119 1391
rect 1125 1385 1126 1391
rect 1118 1347 1126 1385
rect 1118 1341 1119 1347
rect 1125 1341 1126 1347
rect 1118 1275 1126 1341
rect 1118 1269 1119 1275
rect 1125 1269 1126 1275
rect 1118 1239 1126 1269
rect 1118 1233 1119 1239
rect 1125 1233 1126 1239
rect 1118 1163 1126 1233
rect 1118 1157 1119 1163
rect 1125 1157 1126 1163
rect 1118 1131 1126 1157
rect 1118 1125 1119 1131
rect 1125 1125 1126 1131
rect 1118 1055 1126 1125
rect 1118 1049 1119 1055
rect 1125 1049 1126 1055
rect 1118 1023 1126 1049
rect 1118 1017 1119 1023
rect 1125 1017 1126 1023
rect 1118 943 1126 1017
rect 1118 937 1119 943
rect 1125 937 1126 943
rect 1118 911 1126 937
rect 1118 905 1119 911
rect 1125 905 1126 911
rect 1118 835 1126 905
rect 1118 829 1119 835
rect 1125 829 1126 835
rect 1118 807 1126 829
rect 1118 801 1119 807
rect 1125 801 1126 807
rect 1118 731 1126 801
rect 1118 725 1119 731
rect 1125 725 1126 731
rect 1118 699 1126 725
rect 1118 693 1119 699
rect 1125 693 1126 699
rect 1118 619 1126 693
rect 1118 613 1119 619
rect 1125 613 1126 619
rect 1118 591 1126 613
rect 1118 585 1119 591
rect 1125 585 1126 591
rect 1118 503 1126 585
rect 1118 497 1119 503
rect 1125 497 1126 503
rect 1118 483 1126 497
rect 1118 477 1119 483
rect 1125 477 1126 483
rect 1118 387 1126 477
rect 1118 381 1119 387
rect 1125 381 1126 387
rect 1118 375 1126 381
rect 1118 369 1119 375
rect 1125 369 1126 375
rect 1118 271 1126 369
rect 1118 265 1119 271
rect 1125 265 1126 271
rect 1118 263 1126 265
rect 1118 257 1119 263
rect 1125 257 1126 263
rect 1118 139 1126 257
rect 1118 133 1119 139
rect 1125 133 1126 139
rect 1118 131 1126 133
rect 1118 125 1119 131
rect 1125 125 1126 131
rect 1118 72 1126 125
rect 2142 2163 2150 2232
rect 2142 2157 2143 2163
rect 2149 2157 2150 2163
rect 2142 2055 2150 2157
rect 2142 2049 2143 2055
rect 2149 2049 2150 2055
rect 2142 1947 2150 2049
rect 2142 1941 2143 1947
rect 2149 1941 2150 1947
rect 2142 1839 2150 1941
rect 2142 1833 2143 1839
rect 2149 1833 2150 1839
rect 2142 1735 2150 1833
rect 2142 1729 2143 1735
rect 2149 1729 2150 1735
rect 2142 1615 2150 1729
rect 2142 1609 2143 1615
rect 2149 1609 2150 1615
rect 2142 1511 2150 1609
rect 2142 1505 2143 1511
rect 2149 1505 2150 1511
rect 2142 1399 2150 1505
rect 2142 1393 2143 1399
rect 2149 1393 2150 1399
rect 2142 1295 2150 1393
rect 2142 1289 2143 1295
rect 2149 1289 2150 1295
rect 2142 1187 2150 1289
rect 2142 1181 2143 1187
rect 2149 1181 2150 1187
rect 2142 1079 2150 1181
rect 2142 1073 2143 1079
rect 2149 1073 2150 1079
rect 2142 963 2150 1073
rect 2142 957 2143 963
rect 2149 957 2150 963
rect 2142 859 2150 957
rect 2142 853 2143 859
rect 2149 853 2150 859
rect 2142 751 2150 853
rect 2142 745 2143 751
rect 2149 745 2150 751
rect 2142 647 2150 745
rect 2142 641 2143 647
rect 2149 641 2150 647
rect 2142 535 2150 641
rect 2142 529 2143 535
rect 2149 529 2150 535
rect 2142 431 2150 529
rect 2142 425 2143 431
rect 2149 425 2150 431
rect 2142 315 2150 425
rect 2142 309 2143 315
rect 2149 309 2150 315
rect 2142 79 2150 309
rect 2142 73 2143 79
rect 2149 73 2150 79
rect 2142 72 2150 73
rect 2154 2215 2162 2232
rect 2154 2209 2155 2215
rect 2161 2209 2162 2215
rect 2154 2107 2162 2209
rect 2154 2101 2155 2107
rect 2161 2101 2162 2107
rect 2154 2003 2162 2101
rect 2154 1997 2155 2003
rect 2161 1997 2162 2003
rect 2154 1891 2162 1997
rect 2154 1885 2155 1891
rect 2161 1885 2162 1891
rect 2154 1787 2162 1885
rect 2154 1781 2155 1787
rect 2161 1781 2162 1787
rect 2154 1679 2162 1781
rect 2154 1673 2155 1679
rect 2161 1673 2162 1679
rect 2154 1563 2162 1673
rect 2154 1557 2155 1563
rect 2161 1557 2162 1563
rect 2154 1455 2162 1557
rect 2154 1449 2155 1455
rect 2161 1449 2162 1455
rect 2154 1347 2162 1449
rect 2154 1341 2155 1347
rect 2161 1341 2162 1347
rect 2154 1239 2162 1341
rect 2154 1233 2155 1239
rect 2161 1233 2162 1239
rect 2154 1131 2162 1233
rect 2154 1125 2155 1131
rect 2161 1125 2162 1131
rect 2154 1023 2162 1125
rect 2154 1017 2155 1023
rect 2161 1017 2162 1023
rect 2154 911 2162 1017
rect 2154 905 2155 911
rect 2161 905 2162 911
rect 2154 807 2162 905
rect 2154 801 2155 807
rect 2161 801 2162 807
rect 2154 699 2162 801
rect 2154 693 2155 699
rect 2161 693 2162 699
rect 2154 591 2162 693
rect 2154 585 2155 591
rect 2161 585 2162 591
rect 2154 483 2162 585
rect 2154 477 2155 483
rect 2161 477 2162 483
rect 2154 375 2162 477
rect 2154 369 2155 375
rect 2161 369 2162 375
rect 2154 263 2162 369
rect 2154 257 2155 263
rect 2161 257 2162 263
rect 2154 131 2162 257
rect 2154 125 2155 131
rect 2161 125 2162 131
rect 2154 72 2162 125
use circuitwell  npwells
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use circuitppnp  ppnps
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use welltap_svt  __well_tap__147
timestamp 1731220634
transform 1 0 2112 0 1 2164
box 7 3 12 24
use welltap_svt  __well_tap__146
timestamp 1731220634
transform 1 0 1128 0 1 2164
box 7 3 12 24
use welltap_svt  __well_tap__145
timestamp 1731220634
transform 1 0 2112 0 -1 2156
box 7 3 12 24
use welltap_svt  __well_tap__144
timestamp 1731220634
transform 1 0 1128 0 -1 2156
box 7 3 12 24
use welltap_svt  __well_tap__143
timestamp 1731220634
transform 1 0 2112 0 1 2056
box 7 3 12 24
use welltap_svt  __well_tap__142
timestamp 1731220634
transform 1 0 1128 0 1 2056
box 7 3 12 24
use welltap_svt  __well_tap__141
timestamp 1731220634
transform 1 0 2112 0 -1 2048
box 7 3 12 24
use welltap_svt  __well_tap__140
timestamp 1731220634
transform 1 0 1128 0 -1 2048
box 7 3 12 24
use welltap_svt  __well_tap__139
timestamp 1731220634
transform 1 0 2112 0 1 1952
box 7 3 12 24
use welltap_svt  __well_tap__138
timestamp 1731220634
transform 1 0 1128 0 1 1952
box 7 3 12 24
use welltap_svt  __well_tap__137
timestamp 1731220634
transform 1 0 2112 0 -1 1940
box 7 3 12 24
use welltap_svt  __well_tap__136
timestamp 1731220634
transform 1 0 1128 0 -1 1940
box 7 3 12 24
use welltap_svt  __well_tap__135
timestamp 1731220634
transform 1 0 2112 0 1 1840
box 7 3 12 24
use welltap_svt  __well_tap__134
timestamp 1731220634
transform 1 0 1128 0 1 1840
box 7 3 12 24
use welltap_svt  __well_tap__133
timestamp 1731220634
transform 1 0 2112 0 -1 1832
box 7 3 12 24
use welltap_svt  __well_tap__132
timestamp 1731220634
transform 1 0 1128 0 -1 1832
box 7 3 12 24
use welltap_svt  __well_tap__131
timestamp 1731220634
transform 1 0 2112 0 1 1736
box 7 3 12 24
use welltap_svt  __well_tap__130
timestamp 1731220634
transform 1 0 1128 0 1 1736
box 7 3 12 24
use welltap_svt  __well_tap__129
timestamp 1731220634
transform 1 0 2112 0 -1 1728
box 7 3 12 24
use welltap_svt  __well_tap__128
timestamp 1731220634
transform 1 0 1128 0 -1 1728
box 7 3 12 24
use welltap_svt  __well_tap__127
timestamp 1731220634
transform 1 0 2112 0 1 1628
box 7 3 12 24
use welltap_svt  __well_tap__126
timestamp 1731220634
transform 1 0 1128 0 1 1628
box 7 3 12 24
use welltap_svt  __well_tap__125
timestamp 1731220634
transform 1 0 2112 0 -1 1608
box 7 3 12 24
use welltap_svt  __well_tap__124
timestamp 1731220634
transform 1 0 1128 0 -1 1608
box 7 3 12 24
use welltap_svt  __well_tap__123
timestamp 1731220634
transform 1 0 2112 0 1 1512
box 7 3 12 24
use welltap_svt  __well_tap__122
timestamp 1731220634
transform 1 0 1128 0 1 1512
box 7 3 12 24
use welltap_svt  __well_tap__121
timestamp 1731220634
transform 1 0 2112 0 -1 1504
box 7 3 12 24
use welltap_svt  __well_tap__120
timestamp 1731220634
transform 1 0 1128 0 -1 1504
box 7 3 12 24
use welltap_svt  __well_tap__119
timestamp 1731220634
transform 1 0 2112 0 1 1404
box 7 3 12 24
use welltap_svt  __well_tap__118
timestamp 1731220634
transform 1 0 1128 0 1 1404
box 7 3 12 24
use welltap_svt  __well_tap__117
timestamp 1731220634
transform 1 0 2112 0 -1 1392
box 7 3 12 24
use welltap_svt  __well_tap__116
timestamp 1731220634
transform 1 0 1128 0 -1 1392
box 7 3 12 24
use welltap_svt  __well_tap__115
timestamp 1731220634
transform 1 0 2112 0 1 1296
box 7 3 12 24
use welltap_svt  __well_tap__114
timestamp 1731220634
transform 1 0 1128 0 1 1296
box 7 3 12 24
use welltap_svt  __well_tap__113
timestamp 1731220634
transform 1 0 2112 0 -1 1288
box 7 3 12 24
use welltap_svt  __well_tap__112
timestamp 1731220634
transform 1 0 1128 0 -1 1288
box 7 3 12 24
use welltap_svt  __well_tap__111
timestamp 1731220634
transform 1 0 2112 0 1 1188
box 7 3 12 24
use welltap_svt  __well_tap__110
timestamp 1731220634
transform 1 0 1128 0 1 1188
box 7 3 12 24
use welltap_svt  __well_tap__109
timestamp 1731220634
transform 1 0 2112 0 -1 1180
box 7 3 12 24
use welltap_svt  __well_tap__108
timestamp 1731220634
transform 1 0 1128 0 -1 1180
box 7 3 12 24
use welltap_svt  __well_tap__107
timestamp 1731220634
transform 1 0 2112 0 1 1080
box 7 3 12 24
use welltap_svt  __well_tap__106
timestamp 1731220634
transform 1 0 1128 0 1 1080
box 7 3 12 24
use welltap_svt  __well_tap__105
timestamp 1731220634
transform 1 0 2112 0 -1 1072
box 7 3 12 24
use welltap_svt  __well_tap__104
timestamp 1731220634
transform 1 0 1128 0 -1 1072
box 7 3 12 24
use welltap_svt  __well_tap__103
timestamp 1731220634
transform 1 0 2112 0 1 972
box 7 3 12 24
use welltap_svt  __well_tap__102
timestamp 1731220634
transform 1 0 1128 0 1 972
box 7 3 12 24
use welltap_svt  __well_tap__101
timestamp 1731220634
transform 1 0 2112 0 -1 956
box 7 3 12 24
use welltap_svt  __well_tap__100
timestamp 1731220634
transform 1 0 1128 0 -1 956
box 7 3 12 24
use welltap_svt  __well_tap__99
timestamp 1731220634
transform 1 0 2112 0 1 860
box 7 3 12 24
use welltap_svt  __well_tap__98
timestamp 1731220634
transform 1 0 1128 0 1 860
box 7 3 12 24
use welltap_svt  __well_tap__97
timestamp 1731220634
transform 1 0 2112 0 -1 852
box 7 3 12 24
use welltap_svt  __well_tap__96
timestamp 1731220634
transform 1 0 1128 0 -1 852
box 7 3 12 24
use welltap_svt  __well_tap__95
timestamp 1731220634
transform 1 0 2112 0 1 756
box 7 3 12 24
use welltap_svt  __well_tap__94
timestamp 1731220634
transform 1 0 1128 0 1 756
box 7 3 12 24
use welltap_svt  __well_tap__93
timestamp 1731220634
transform 1 0 2112 0 -1 744
box 7 3 12 24
use welltap_svt  __well_tap__92
timestamp 1731220634
transform 1 0 1128 0 -1 744
box 7 3 12 24
use welltap_svt  __well_tap__91
timestamp 1731220634
transform 1 0 2112 0 1 648
box 7 3 12 24
use welltap_svt  __well_tap__90
timestamp 1731220634
transform 1 0 1128 0 1 648
box 7 3 12 24
use welltap_svt  __well_tap__89
timestamp 1731220634
transform 1 0 2112 0 -1 640
box 7 3 12 24
use welltap_svt  __well_tap__88
timestamp 1731220634
transform 1 0 1128 0 -1 640
box 7 3 12 24
use welltap_svt  __well_tap__87
timestamp 1731220634
transform 1 0 2112 0 1 540
box 7 3 12 24
use welltap_svt  __well_tap__86
timestamp 1731220634
transform 1 0 1128 0 1 540
box 7 3 12 24
use welltap_svt  __well_tap__85
timestamp 1731220634
transform 1 0 2112 0 -1 528
box 7 3 12 24
use welltap_svt  __well_tap__84
timestamp 1731220634
transform 1 0 1128 0 -1 528
box 7 3 12 24
use welltap_svt  __well_tap__83
timestamp 1731220634
transform 1 0 2112 0 1 432
box 7 3 12 24
use welltap_svt  __well_tap__82
timestamp 1731220634
transform 1 0 1128 0 1 432
box 7 3 12 24
use welltap_svt  __well_tap__81
timestamp 1731220634
transform 1 0 2112 0 -1 424
box 7 3 12 24
use welltap_svt  __well_tap__80
timestamp 1731220634
transform 1 0 1128 0 -1 424
box 7 3 12 24
use welltap_svt  __well_tap__79
timestamp 1731220634
transform 1 0 2112 0 1 324
box 7 3 12 24
use welltap_svt  __well_tap__78
timestamp 1731220634
transform 1 0 1128 0 1 324
box 7 3 12 24
use welltap_svt  __well_tap__77
timestamp 1731220634
transform 1 0 2112 0 -1 308
box 7 3 12 24
use welltap_svt  __well_tap__76
timestamp 1731220634
transform 1 0 1128 0 -1 308
box 7 3 12 24
use welltap_svt  __well_tap__75
timestamp 1731220634
transform 1 0 2112 0 1 212
box 7 3 12 24
use welltap_svt  __well_tap__74
timestamp 1731220634
transform 1 0 1128 0 1 212
box 7 3 12 24
use welltap_svt  __well_tap__73
timestamp 1731220634
transform 1 0 2112 0 -1 200
box 7 3 12 24
use welltap_svt  __well_tap__72
timestamp 1731220634
transform 1 0 1128 0 -1 200
box 7 3 12 24
use welltap_svt  __well_tap__71
timestamp 1731220634
transform 1 0 2112 0 1 80
box 7 3 12 24
use welltap_svt  __well_tap__70
timestamp 1731220634
transform 1 0 1128 0 1 80
box 7 3 12 24
use welltap_svt  __well_tap__69
timestamp 1731220634
transform 1 0 1088 0 1 1984
box 7 3 12 24
use welltap_svt  __well_tap__68
timestamp 1731220634
transform 1 0 104 0 1 1984
box 7 3 12 24
use welltap_svt  __well_tap__67
timestamp 1731220634
transform 1 0 1088 0 -1 1976
box 7 3 12 24
use welltap_svt  __well_tap__66
timestamp 1731220634
transform 1 0 104 0 -1 1976
box 7 3 12 24
use welltap_svt  __well_tap__65
timestamp 1731220634
transform 1 0 1088 0 1 1880
box 7 3 12 24
use welltap_svt  __well_tap__64
timestamp 1731220634
transform 1 0 104 0 1 1880
box 7 3 12 24
use welltap_svt  __well_tap__63
timestamp 1731220634
transform 1 0 1088 0 -1 1868
box 7 3 12 24
use welltap_svt  __well_tap__62
timestamp 1731220634
transform 1 0 104 0 -1 1868
box 7 3 12 24
use welltap_svt  __well_tap__61
timestamp 1731220634
transform 1 0 1088 0 1 1764
box 7 3 12 24
use welltap_svt  __well_tap__60
timestamp 1731220634
transform 1 0 104 0 1 1764
box 7 3 12 24
use welltap_svt  __well_tap__59
timestamp 1731220634
transform 1 0 1088 0 -1 1756
box 7 3 12 24
use welltap_svt  __well_tap__58
timestamp 1731220634
transform 1 0 104 0 -1 1756
box 7 3 12 24
use welltap_svt  __well_tap__57
timestamp 1731220634
transform 1 0 1088 0 1 1656
box 7 3 12 24
use welltap_svt  __well_tap__56
timestamp 1731220634
transform 1 0 104 0 1 1656
box 7 3 12 24
use welltap_svt  __well_tap__55
timestamp 1731220634
transform 1 0 1088 0 -1 1644
box 7 3 12 24
use welltap_svt  __well_tap__54
timestamp 1731220634
transform 1 0 104 0 -1 1644
box 7 3 12 24
use welltap_svt  __well_tap__53
timestamp 1731220634
transform 1 0 1088 0 1 1548
box 7 3 12 24
use welltap_svt  __well_tap__52
timestamp 1731220634
transform 1 0 104 0 1 1548
box 7 3 12 24
use welltap_svt  __well_tap__51
timestamp 1731220634
transform 1 0 1088 0 -1 1540
box 7 3 12 24
use welltap_svt  __well_tap__50
timestamp 1731220634
transform 1 0 104 0 -1 1540
box 7 3 12 24
use welltap_svt  __well_tap__49
timestamp 1731220634
transform 1 0 1088 0 1 1444
box 7 3 12 24
use welltap_svt  __well_tap__48
timestamp 1731220634
transform 1 0 104 0 1 1444
box 7 3 12 24
use welltap_svt  __well_tap__47
timestamp 1731220634
transform 1 0 1088 0 -1 1436
box 7 3 12 24
use welltap_svt  __well_tap__46
timestamp 1731220634
transform 1 0 104 0 -1 1436
box 7 3 12 24
use welltap_svt  __well_tap__45
timestamp 1731220634
transform 1 0 1088 0 1 1340
box 7 3 12 24
use welltap_svt  __well_tap__44
timestamp 1731220634
transform 1 0 104 0 1 1340
box 7 3 12 24
use welltap_svt  __well_tap__43
timestamp 1731220634
transform 1 0 1088 0 -1 1324
box 7 3 12 24
use welltap_svt  __well_tap__42
timestamp 1731220634
transform 1 0 104 0 -1 1324
box 7 3 12 24
use welltap_svt  __well_tap__41
timestamp 1731220634
transform 1 0 1088 0 1 1224
box 7 3 12 24
use welltap_svt  __well_tap__40
timestamp 1731220634
transform 1 0 104 0 1 1224
box 7 3 12 24
use welltap_svt  __well_tap__39
timestamp 1731220634
transform 1 0 1088 0 -1 1212
box 7 3 12 24
use welltap_svt  __well_tap__38
timestamp 1731220634
transform 1 0 104 0 -1 1212
box 7 3 12 24
use welltap_svt  __well_tap__37
timestamp 1731220634
transform 1 0 1088 0 1 1112
box 7 3 12 24
use welltap_svt  __well_tap__36
timestamp 1731220634
transform 1 0 104 0 1 1112
box 7 3 12 24
use welltap_svt  __well_tap__35
timestamp 1731220634
transform 1 0 1088 0 -1 1104
box 7 3 12 24
use welltap_svt  __well_tap__34
timestamp 1731220634
transform 1 0 104 0 -1 1104
box 7 3 12 24
use welltap_svt  __well_tap__33
timestamp 1731220634
transform 1 0 1088 0 1 1004
box 7 3 12 24
use welltap_svt  __well_tap__32
timestamp 1731220634
transform 1 0 104 0 1 1004
box 7 3 12 24
use welltap_svt  __well_tap__31
timestamp 1731220634
transform 1 0 1088 0 -1 992
box 7 3 12 24
use welltap_svt  __well_tap__30
timestamp 1731220634
transform 1 0 104 0 -1 992
box 7 3 12 24
use welltap_svt  __well_tap__29
timestamp 1731220634
transform 1 0 1088 0 1 892
box 7 3 12 24
use welltap_svt  __well_tap__28
timestamp 1731220634
transform 1 0 104 0 1 892
box 7 3 12 24
use welltap_svt  __well_tap__27
timestamp 1731220634
transform 1 0 1088 0 -1 880
box 7 3 12 24
use welltap_svt  __well_tap__26
timestamp 1731220634
transform 1 0 104 0 -1 880
box 7 3 12 24
use welltap_svt  __well_tap__25
timestamp 1731220634
transform 1 0 1088 0 1 784
box 7 3 12 24
use welltap_svt  __well_tap__24
timestamp 1731220634
transform 1 0 104 0 1 784
box 7 3 12 24
use welltap_svt  __well_tap__23
timestamp 1731220634
transform 1 0 1088 0 -1 776
box 7 3 12 24
use welltap_svt  __well_tap__22
timestamp 1731220634
transform 1 0 104 0 -1 776
box 7 3 12 24
use welltap_svt  __well_tap__21
timestamp 1731220634
transform 1 0 1088 0 1 680
box 7 3 12 24
use welltap_svt  __well_tap__20
timestamp 1731220634
transform 1 0 104 0 1 680
box 7 3 12 24
use welltap_svt  __well_tap__19
timestamp 1731220634
transform 1 0 1088 0 -1 672
box 7 3 12 24
use welltap_svt  __well_tap__18
timestamp 1731220634
transform 1 0 104 0 -1 672
box 7 3 12 24
use welltap_svt  __well_tap__17
timestamp 1731220634
transform 1 0 1088 0 1 568
box 7 3 12 24
use welltap_svt  __well_tap__16
timestamp 1731220634
transform 1 0 104 0 1 568
box 7 3 12 24
use welltap_svt  __well_tap__15
timestamp 1731220634
transform 1 0 1088 0 -1 556
box 7 3 12 24
use welltap_svt  __well_tap__14
timestamp 1731220634
transform 1 0 104 0 -1 556
box 7 3 12 24
use welltap_svt  __well_tap__13
timestamp 1731220634
transform 1 0 1088 0 1 452
box 7 3 12 24
use welltap_svt  __well_tap__12
timestamp 1731220634
transform 1 0 104 0 1 452
box 7 3 12 24
use welltap_svt  __well_tap__11
timestamp 1731220634
transform 1 0 1088 0 -1 440
box 7 3 12 24
use welltap_svt  __well_tap__10
timestamp 1731220634
transform 1 0 104 0 -1 440
box 7 3 12 24
use welltap_svt  __well_tap__9
timestamp 1731220634
transform 1 0 1088 0 1 336
box 7 3 12 24
use welltap_svt  __well_tap__8
timestamp 1731220634
transform 1 0 104 0 1 336
box 7 3 12 24
use welltap_svt  __well_tap__7
timestamp 1731220634
transform 1 0 1088 0 -1 324
box 7 3 12 24
use welltap_svt  __well_tap__6
timestamp 1731220634
transform 1 0 104 0 -1 324
box 7 3 12 24
use welltap_svt  __well_tap__5
timestamp 1731220634
transform 1 0 1088 0 1 220
box 7 3 12 24
use welltap_svt  __well_tap__4
timestamp 1731220634
transform 1 0 104 0 1 220
box 7 3 12 24
use welltap_svt  __well_tap__3
timestamp 1731220634
transform 1 0 1088 0 -1 200
box 7 3 12 24
use welltap_svt  __well_tap__2
timestamp 1731220634
transform 1 0 104 0 -1 200
box 7 3 12 24
use welltap_svt  __well_tap__1
timestamp 1731220634
transform 1 0 1088 0 1 88
box 7 3 12 24
use welltap_svt  __well_tap__0
timestamp 1731220634
transform 1 0 104 0 1 88
box 7 3 12 24
use _0_0std_0_0cells_0_0NOR2X1  tst_5999_6
timestamp 1731220634
transform 1 0 128 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5998_6
timestamp 1731220634
transform 1 0 168 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5997_6
timestamp 1731220634
transform 1 0 208 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5996_6
timestamp 1731220634
transform 1 0 248 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5995_6
timestamp 1731220634
transform 1 0 288 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5994_6
timestamp 1731220634
transform 1 0 328 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5993_6
timestamp 1731220634
transform 1 0 368 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5992_6
timestamp 1731220634
transform 1 0 408 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5991_6
timestamp 1731220634
transform 1 0 448 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5990_6
timestamp 1731220634
transform 1 0 488 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5989_6
timestamp 1731220634
transform 1 0 160 0 -1 204
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5988_6
timestamp 1731220634
transform 1 0 200 0 -1 204
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5987_6
timestamp 1731220634
transform 1 0 240 0 -1 204
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5986_6
timestamp 1731220634
transform 1 0 288 0 -1 204
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5985_6
timestamp 1731220634
transform 1 0 336 0 -1 204
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5984_6
timestamp 1731220634
transform 1 0 392 0 -1 204
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5983_6
timestamp 1731220634
transform 1 0 456 0 -1 204
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5982_6
timestamp 1731220634
transform 1 0 280 0 1 216
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5981_6
timestamp 1731220634
transform 1 0 320 0 1 216
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5980_6
timestamp 1731220634
transform 1 0 360 0 1 216
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5979_6
timestamp 1731220634
transform 1 0 408 0 1 216
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5978_6
timestamp 1731220634
transform 1 0 464 0 1 216
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5977_6
timestamp 1731220634
transform 1 0 528 0 1 216
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5976_6
timestamp 1731220634
transform 1 0 600 0 1 216
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5975_6
timestamp 1731220634
transform 1 0 376 0 -1 328
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5974_6
timestamp 1731220634
transform 1 0 416 0 -1 328
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5973_6
timestamp 1731220634
transform 1 0 456 0 -1 328
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5972_6
timestamp 1731220634
transform 1 0 496 0 -1 328
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5971_6
timestamp 1731220634
transform 1 0 536 0 -1 328
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5970_6
timestamp 1731220634
transform 1 0 584 0 -1 328
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5969_6
timestamp 1731220634
transform 1 0 632 0 -1 328
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5968_6
timestamp 1731220634
transform 1 0 680 0 -1 328
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5967_6
timestamp 1731220634
transform 1 0 672 0 1 216
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5966_6
timestamp 1731220634
transform 1 0 664 0 -1 204
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5965_6
timestamp 1731220634
transform 1 0 592 0 -1 204
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5964_6
timestamp 1731220634
transform 1 0 520 0 -1 204
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5963_6
timestamp 1731220634
transform 1 0 528 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5962_6
timestamp 1731220634
transform 1 0 568 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5961_6
timestamp 1731220634
transform 1 0 608 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5960_6
timestamp 1731220634
transform 1 0 648 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5959_6
timestamp 1731220634
transform 1 0 688 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5958_6
timestamp 1731220634
transform 1 0 728 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5957_6
timestamp 1731220634
transform 1 0 768 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5956_6
timestamp 1731220634
transform 1 0 808 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5955_6
timestamp 1731220634
transform 1 0 864 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5954_6
timestamp 1731220634
transform 1 0 928 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5953_6
timestamp 1731220634
transform 1 0 904 0 -1 204
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5952_6
timestamp 1731220634
transform 1 0 824 0 -1 204
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5951_6
timestamp 1731220634
transform 1 0 744 0 -1 204
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5950_6
timestamp 1731220634
transform 1 0 800 0 1 216
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5949_6
timestamp 1731220634
transform 1 0 736 0 1 216
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5948_6
timestamp 1731220634
transform 1 0 728 0 -1 328
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5947_6
timestamp 1731220634
transform 1 0 776 0 -1 328
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5946_6
timestamp 1731220634
transform 1 0 824 0 -1 328
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5945_6
timestamp 1731220634
transform 1 0 872 0 -1 328
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5944_6
timestamp 1731220634
transform 1 0 856 0 1 216
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5943_6
timestamp 1731220634
transform 1 0 920 0 1 216
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5942_6
timestamp 1731220634
transform 1 0 984 0 1 216
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5941_6
timestamp 1731220634
transform 1 0 1040 0 1 216
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5940_6
timestamp 1731220634
transform 1 0 1040 0 -1 204
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5939_6
timestamp 1731220634
transform 1 0 984 0 -1 204
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5938_6
timestamp 1731220634
transform 1 0 992 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5937_6
timestamp 1731220634
transform 1 0 1040 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5936_6
timestamp 1731220634
transform 1 0 1152 0 1 76
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5935_6
timestamp 1731220634
transform 1 0 1192 0 1 76
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5934_6
timestamp 1731220634
transform 1 0 1232 0 1 76
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5933_6
timestamp 1731220634
transform 1 0 1272 0 1 76
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5932_6
timestamp 1731220634
transform 1 0 1312 0 1 76
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5931_6
timestamp 1731220634
transform 1 0 1360 0 1 76
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5930_6
timestamp 1731220634
transform 1 0 1424 0 1 76
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5929_6
timestamp 1731220634
transform 1 0 1488 0 1 76
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5928_6
timestamp 1731220634
transform 1 0 1176 0 -1 204
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5927_6
timestamp 1731220634
transform 1 0 1224 0 -1 204
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5926_6
timestamp 1731220634
transform 1 0 1288 0 -1 204
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5925_6
timestamp 1731220634
transform 1 0 1352 0 -1 204
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5924_6
timestamp 1731220634
transform 1 0 1424 0 -1 204
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5923_6
timestamp 1731220634
transform 1 0 1504 0 -1 204
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5922_6
timestamp 1731220634
transform 1 0 1256 0 1 208
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5921_6
timestamp 1731220634
transform 1 0 1296 0 1 208
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5920_6
timestamp 1731220634
transform 1 0 1336 0 1 208
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5919_6
timestamp 1731220634
transform 1 0 1376 0 1 208
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5918_6
timestamp 1731220634
transform 1 0 1416 0 1 208
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5917_6
timestamp 1731220634
transform 1 0 1456 0 1 208
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5916_6
timestamp 1731220634
transform 1 0 1496 0 1 208
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5915_6
timestamp 1731220634
transform 1 0 1344 0 -1 312
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5914_6
timestamp 1731220634
transform 1 0 1384 0 -1 312
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5913_6
timestamp 1731220634
transform 1 0 1424 0 -1 312
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5912_6
timestamp 1731220634
transform 1 0 1464 0 -1 312
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5911_6
timestamp 1731220634
transform 1 0 1504 0 -1 312
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5910_6
timestamp 1731220634
transform 1 0 1552 0 -1 312
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5909_6
timestamp 1731220634
transform 1 0 1608 0 -1 312
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5908_6
timestamp 1731220634
transform 1 0 1664 0 -1 312
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5907_6
timestamp 1731220634
transform 1 0 1728 0 -1 312
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5906_6
timestamp 1731220634
transform 1 0 1800 0 -1 312
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5905_6
timestamp 1731220634
transform 1 0 1536 0 1 208
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5904_6
timestamp 1731220634
transform 1 0 1592 0 1 208
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5903_6
timestamp 1731220634
transform 1 0 1664 0 1 208
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5902_6
timestamp 1731220634
transform 1 0 1752 0 1 208
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5901_6
timestamp 1731220634
transform 1 0 1856 0 1 208
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5900_6
timestamp 1731220634
transform 1 0 1968 0 1 208
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5899_6
timestamp 1731220634
transform 1 0 1584 0 -1 204
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5898_6
timestamp 1731220634
transform 1 0 1656 0 -1 204
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5897_6
timestamp 1731220634
transform 1 0 1728 0 -1 204
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5896_6
timestamp 1731220634
transform 1 0 1800 0 -1 204
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5895_6
timestamp 1731220634
transform 1 0 1552 0 1 76
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5894_6
timestamp 1731220634
transform 1 0 1608 0 1 76
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5893_6
timestamp 1731220634
transform 1 0 1664 0 1 76
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5892_6
timestamp 1731220634
transform 1 0 1712 0 1 76
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5891_6
timestamp 1731220634
transform 1 0 1760 0 1 76
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5890_6
timestamp 1731220634
transform 1 0 1800 0 1 76
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5889_6
timestamp 1731220634
transform 1 0 1848 0 1 76
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5888_6
timestamp 1731220634
transform 1 0 1896 0 1 76
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5887_6
timestamp 1731220634
transform 1 0 1944 0 1 76
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5886_6
timestamp 1731220634
transform 1 0 1872 0 -1 204
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5885_6
timestamp 1731220634
transform 1 0 1944 0 -1 204
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5884_6
timestamp 1731220634
transform 1 0 1984 0 1 76
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5883_6
timestamp 1731220634
transform 1 0 2024 0 1 76
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5882_6
timestamp 1731220634
transform 1 0 2064 0 1 76
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5881_6
timestamp 1731220634
transform 1 0 2064 0 -1 204
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5880_6
timestamp 1731220634
transform 1 0 2016 0 -1 204
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5879_6
timestamp 1731220634
transform 1 0 2064 0 1 208
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5878_6
timestamp 1731220634
transform 1 0 2040 0 -1 312
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5877_6
timestamp 1731220634
transform 1 0 1960 0 -1 312
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5876_6
timestamp 1731220634
transform 1 0 1880 0 -1 312
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5875_6
timestamp 1731220634
transform 1 0 1856 0 1 320
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5874_6
timestamp 1731220634
transform 1 0 1792 0 1 320
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5873_6
timestamp 1731220634
transform 1 0 1720 0 1 320
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5872_6
timestamp 1731220634
transform 1 0 1552 0 1 320
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5871_6
timestamp 1731220634
transform 1 0 1640 0 1 320
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5870_6
timestamp 1731220634
transform 1 0 1664 0 -1 428
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5869_6
timestamp 1731220634
transform 1 0 1744 0 -1 428
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5868_6
timestamp 1731220634
transform 1 0 1824 0 -1 428
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5867_6
timestamp 1731220634
transform 1 0 1584 0 -1 428
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5866_6
timestamp 1731220634
transform 1 0 1576 0 1 428
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5865_6
timestamp 1731220634
transform 1 0 1640 0 1 428
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5864_6
timestamp 1731220634
transform 1 0 1712 0 1 428
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5863_6
timestamp 1731220634
transform 1 0 1800 0 1 428
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5862_6
timestamp 1731220634
transform 1 0 1888 0 1 428
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5861_6
timestamp 1731220634
transform 1 0 1832 0 -1 532
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5860_6
timestamp 1731220634
transform 1 0 1760 0 -1 532
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5859_6
timestamp 1731220634
transform 1 0 1696 0 -1 532
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5858_6
timestamp 1731220634
transform 1 0 1640 0 -1 532
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5857_6
timestamp 1731220634
transform 1 0 1584 0 -1 532
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5856_6
timestamp 1731220634
transform 1 0 1480 0 1 536
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5855_6
timestamp 1731220634
transform 1 0 1560 0 1 536
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5854_6
timestamp 1731220634
transform 1 0 1648 0 1 536
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5853_6
timestamp 1731220634
transform 1 0 1744 0 1 536
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5852_6
timestamp 1731220634
transform 1 0 1488 0 -1 644
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5851_6
timestamp 1731220634
transform 1 0 1576 0 -1 644
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5850_6
timestamp 1731220634
transform 1 0 1664 0 -1 644
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5849_6
timestamp 1731220634
transform 1 0 1752 0 -1 644
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5848_6
timestamp 1731220634
transform 1 0 1576 0 1 644
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5847_6
timestamp 1731220634
transform 1 0 1648 0 1 644
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5846_6
timestamp 1731220634
transform 1 0 1728 0 1 644
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5845_6
timestamp 1731220634
transform 1 0 1816 0 1 644
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5844_6
timestamp 1731220634
transform 1 0 1648 0 -1 748
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5843_6
timestamp 1731220634
transform 1 0 1704 0 -1 748
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5842_6
timestamp 1731220634
transform 1 0 1760 0 -1 748
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5841_6
timestamp 1731220634
transform 1 0 1824 0 -1 748
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5840_6
timestamp 1731220634
transform 1 0 1712 0 1 752
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5839_6
timestamp 1731220634
transform 1 0 1616 0 1 752
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5838_6
timestamp 1731220634
transform 1 0 1512 0 1 752
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5837_6
timestamp 1731220634
transform 1 0 1536 0 -1 856
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5836_6
timestamp 1731220634
transform 1 0 1624 0 -1 856
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5835_6
timestamp 1731220634
transform 1 0 1704 0 -1 856
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5834_6
timestamp 1731220634
transform 1 0 1656 0 1 856
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5833_6
timestamp 1731220634
transform 1 0 1736 0 1 856
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5832_6
timestamp 1731220634
transform 1 0 1776 0 -1 856
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5831_6
timestamp 1731220634
transform 1 0 1848 0 -1 856
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5830_6
timestamp 1731220634
transform 1 0 1928 0 -1 856
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5829_6
timestamp 1731220634
transform 1 0 1808 0 1 752
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5828_6
timestamp 1731220634
transform 1 0 1896 0 1 752
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5827_6
timestamp 1731220634
transform 1 0 1992 0 1 752
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5826_6
timestamp 1731220634
transform 1 0 1952 0 -1 748
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5825_6
timestamp 1731220634
transform 1 0 1888 0 -1 748
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5824_6
timestamp 1731220634
transform 1 0 1904 0 1 644
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5823_6
timestamp 1731220634
transform 1 0 1992 0 1 644
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5822_6
timestamp 1731220634
transform 1 0 1912 0 -1 644
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5821_6
timestamp 1731220634
transform 1 0 1832 0 -1 644
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5820_6
timestamp 1731220634
transform 1 0 1848 0 1 536
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5819_6
timestamp 1731220634
transform 1 0 1960 0 1 536
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5818_6
timestamp 1731220634
transform 1 0 1912 0 -1 532
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5817_6
timestamp 1731220634
transform 1 0 1984 0 1 428
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5816_6
timestamp 1731220634
transform 1 0 1992 0 -1 428
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5815_6
timestamp 1731220634
transform 1 0 1904 0 -1 428
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5814_6
timestamp 1731220634
transform 1 0 1912 0 1 320
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5813_6
timestamp 1731220634
transform 1 0 1968 0 1 320
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5812_6
timestamp 1731220634
transform 1 0 2024 0 1 320
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5811_6
timestamp 1731220634
transform 1 0 2064 0 1 320
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5810_6
timestamp 1731220634
transform 1 0 2064 0 -1 428
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5809_6
timestamp 1731220634
transform 1 0 2064 0 1 428
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5808_6
timestamp 1731220634
transform 1 0 2064 0 -1 532
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5807_6
timestamp 1731220634
transform 1 0 2000 0 -1 532
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5806_6
timestamp 1731220634
transform 1 0 2064 0 1 536
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5805_6
timestamp 1731220634
transform 1 0 2000 0 -1 644
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5804_6
timestamp 1731220634
transform 1 0 2064 0 -1 644
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5803_6
timestamp 1731220634
transform 1 0 2064 0 1 644
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5802_6
timestamp 1731220634
transform 1 0 2016 0 -1 748
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5801_6
timestamp 1731220634
transform 1 0 2064 0 -1 748
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5800_6
timestamp 1731220634
transform 1 0 2064 0 1 752
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5799_6
timestamp 1731220634
transform 1 0 2064 0 -1 856
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5798_6
timestamp 1731220634
transform 1 0 2064 0 1 856
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5797_6
timestamp 1731220634
transform 1 0 2064 0 -1 960
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5796_6
timestamp 1731220634
transform 1 0 2008 0 -1 856
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5795_6
timestamp 1731220634
transform 1 0 1808 0 1 856
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5794_6
timestamp 1731220634
transform 1 0 1880 0 1 856
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5793_6
timestamp 1731220634
transform 1 0 1944 0 1 856
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5792_6
timestamp 1731220634
transform 1 0 2016 0 1 856
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5791_6
timestamp 1731220634
transform 1 0 2016 0 -1 960
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5790_6
timestamp 1731220634
transform 1 0 1944 0 -1 960
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5789_6
timestamp 1731220634
transform 1 0 1872 0 -1 960
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5788_6
timestamp 1731220634
transform 1 0 1808 0 -1 960
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5787_6
timestamp 1731220634
transform 1 0 1608 0 -1 960
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5786_6
timestamp 1731220634
transform 1 0 1680 0 -1 960
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5785_6
timestamp 1731220634
transform 1 0 1744 0 -1 960
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5784_6
timestamp 1731220634
transform 1 0 1784 0 1 968
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5783_6
timestamp 1731220634
transform 1 0 1872 0 1 968
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5782_6
timestamp 1731220634
transform 1 0 1704 0 1 968
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5781_6
timestamp 1731220634
transform 1 0 1512 0 1 968
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5780_6
timestamp 1731220634
transform 1 0 1568 0 1 968
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5779_6
timestamp 1731220634
transform 1 0 1632 0 1 968
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5778_6
timestamp 1731220634
transform 1 0 1656 0 -1 1076
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5777_6
timestamp 1731220634
transform 1 0 1752 0 -1 1076
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5776_6
timestamp 1731220634
transform 1 0 1856 0 -1 1076
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5775_6
timestamp 1731220634
transform 1 0 1576 0 -1 1076
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5774_6
timestamp 1731220634
transform 1 0 1504 0 -1 1076
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5773_6
timestamp 1731220634
transform 1 0 1408 0 1 1076
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5772_6
timestamp 1731220634
transform 1 0 1448 0 -1 1076
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5771_6
timestamp 1731220634
transform 1 0 1480 0 1 1076
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5770_6
timestamp 1731220634
transform 1 0 1560 0 1 1076
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5769_6
timestamp 1731220634
transform 1 0 1648 0 1 1076
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5768_6
timestamp 1731220634
transform 1 0 1744 0 1 1076
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5767_6
timestamp 1731220634
transform 1 0 1848 0 1 1076
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5766_6
timestamp 1731220634
transform 1 0 1552 0 -1 1184
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5765_6
timestamp 1731220634
transform 1 0 1624 0 -1 1184
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5764_6
timestamp 1731220634
transform 1 0 1704 0 -1 1184
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5763_6
timestamp 1731220634
transform 1 0 1792 0 -1 1184
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5762_6
timestamp 1731220634
transform 1 0 1880 0 -1 1184
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5761_6
timestamp 1731220634
transform 1 0 1616 0 1 1184
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5760_6
timestamp 1731220634
transform 1 0 1672 0 1 1184
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5759_6
timestamp 1731220634
transform 1 0 1728 0 1 1184
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5758_6
timestamp 1731220634
transform 1 0 1784 0 1 1184
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5757_6
timestamp 1731220634
transform 1 0 1840 0 1 1184
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5756_6
timestamp 1731220634
transform 1 0 1896 0 1 1184
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5755_6
timestamp 1731220634
transform 1 0 1648 0 -1 1292
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5754_6
timestamp 1731220634
transform 1 0 1736 0 -1 1292
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5753_6
timestamp 1731220634
transform 1 0 1824 0 -1 1292
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5752_6
timestamp 1731220634
transform 1 0 1912 0 -1 1292
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5751_6
timestamp 1731220634
transform 1 0 1672 0 1 1292
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5750_6
timestamp 1731220634
transform 1 0 1752 0 1 1292
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5749_6
timestamp 1731220634
transform 1 0 1824 0 1 1292
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5748_6
timestamp 1731220634
transform 1 0 1888 0 1 1292
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5747_6
timestamp 1731220634
transform 1 0 1952 0 1 1292
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5746_6
timestamp 1731220634
transform 1 0 2016 0 1 1292
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5745_6
timestamp 1731220634
transform 1 0 2000 0 -1 1292
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5744_6
timestamp 1731220634
transform 1 0 1960 0 1 1184
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5743_6
timestamp 1731220634
transform 1 0 1976 0 -1 1184
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5742_6
timestamp 1731220634
transform 1 0 1952 0 1 1076
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5741_6
timestamp 1731220634
transform 1 0 1960 0 1 968
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5740_6
timestamp 1731220634
transform 1 0 2056 0 1 968
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5739_6
timestamp 1731220634
transform 1 0 1960 0 -1 1076
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5738_6
timestamp 1731220634
transform 1 0 2064 0 -1 1076
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5737_6
timestamp 1731220634
transform 1 0 2064 0 1 1076
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5736_6
timestamp 1731220634
transform 1 0 2064 0 -1 1184
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5735_6
timestamp 1731220634
transform 1 0 2024 0 1 1184
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5734_6
timestamp 1731220634
transform 1 0 2064 0 1 1184
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5733_6
timestamp 1731220634
transform 1 0 2064 0 -1 1292
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5732_6
timestamp 1731220634
transform 1 0 2064 0 1 1292
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5731_6
timestamp 1731220634
transform 1 0 2064 0 -1 1396
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5730_6
timestamp 1731220634
transform 1 0 1984 0 -1 1396
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5729_6
timestamp 1731220634
transform 1 0 1968 0 1 1400
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5728_6
timestamp 1731220634
transform 1 0 2056 0 1 1400
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5727_6
timestamp 1731220634
transform 1 0 2056 0 -1 1508
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5726_6
timestamp 1731220634
transform 1 0 1984 0 -1 1508
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5725_6
timestamp 1731220634
transform 1 0 1992 0 1 1508
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5724_6
timestamp 1731220634
transform 1 0 1904 0 1 1508
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5723_6
timestamp 1731220634
transform 1 0 1816 0 1 1508
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5722_6
timestamp 1731220634
transform 1 0 1616 0 -1 1508
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5721_6
timestamp 1731220634
transform 1 0 1696 0 -1 1508
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5720_6
timestamp 1731220634
transform 1 0 1768 0 -1 1508
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5719_6
timestamp 1731220634
transform 1 0 1840 0 -1 1508
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5718_6
timestamp 1731220634
transform 1 0 1880 0 1 1400
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5717_6
timestamp 1731220634
transform 1 0 1800 0 1 1400
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5716_6
timestamp 1731220634
transform 1 0 1728 0 1 1400
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5715_6
timestamp 1731220634
transform 1 0 1544 0 1 1400
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5714_6
timestamp 1731220634
transform 1 0 1600 0 1 1400
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5713_6
timestamp 1731220634
transform 1 0 1664 0 1 1400
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5712_6
timestamp 1731220634
transform 1 0 1712 0 -1 1396
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5711_6
timestamp 1731220634
transform 1 0 1800 0 -1 1396
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5710_6
timestamp 1731220634
transform 1 0 1888 0 -1 1396
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5709_6
timestamp 1731220634
transform 1 0 1640 0 -1 1396
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5708_6
timestamp 1731220634
transform 1 0 1576 0 -1 1396
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5707_6
timestamp 1731220634
transform 1 0 1448 0 -1 1396
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5706_6
timestamp 1731220634
transform 1 0 1488 0 -1 1396
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5705_6
timestamp 1731220634
transform 1 0 1528 0 -1 1396
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5704_6
timestamp 1731220634
transform 1 0 1592 0 1 1292
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5703_6
timestamp 1731220634
transform 1 0 1496 0 1 1292
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5702_6
timestamp 1731220634
transform 1 0 1400 0 1 1292
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5701_6
timestamp 1731220634
transform 1 0 1408 0 -1 1396
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5700_6
timestamp 1731220634
transform 1 0 1368 0 -1 1396
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5699_6
timestamp 1731220634
transform 1 0 1328 0 -1 1396
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5698_6
timestamp 1731220634
transform 1 0 1272 0 1 1400
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5697_6
timestamp 1731220634
transform 1 0 1320 0 1 1400
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5696_6
timestamp 1731220634
transform 1 0 1376 0 1 1400
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5695_6
timestamp 1731220634
transform 1 0 1432 0 1 1400
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5694_6
timestamp 1731220634
transform 1 0 1488 0 1 1400
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5693_6
timestamp 1731220634
transform 1 0 1536 0 -1 1508
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5692_6
timestamp 1731220634
transform 1 0 1448 0 -1 1508
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5691_6
timestamp 1731220634
transform 1 0 1368 0 -1 1508
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5690_6
timestamp 1731220634
transform 1 0 1296 0 -1 1508
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5689_6
timestamp 1731220634
transform 1 0 1232 0 -1 1508
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5688_6
timestamp 1731220634
transform 1 0 1192 0 -1 1508
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5687_6
timestamp 1731220634
transform 1 0 1152 0 -1 1508
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5686_6
timestamp 1731220634
transform 1 0 1152 0 1 1508
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5685_6
timestamp 1731220634
transform 1 0 1192 0 1 1508
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5684_6
timestamp 1731220634
transform 1 0 1240 0 1 1508
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5683_6
timestamp 1731220634
transform 1 0 1312 0 1 1508
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5682_6
timestamp 1731220634
transform 1 0 1392 0 1 1508
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5681_6
timestamp 1731220634
transform 1 0 1472 0 1 1508
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5680_6
timestamp 1731220634
transform 1 0 1376 0 -1 1612
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5679_6
timestamp 1731220634
transform 1 0 1296 0 -1 1612
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5678_6
timestamp 1731220634
transform 1 0 1208 0 -1 1612
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5677_6
timestamp 1731220634
transform 1 0 1152 0 -1 1612
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5676_6
timestamp 1731220634
transform 1 0 1040 0 -1 1648
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5675_6
timestamp 1731220634
transform 1 0 896 0 -1 1648
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5674_6
timestamp 1731220634
transform 1 0 952 0 -1 1648
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5673_6
timestamp 1731220634
transform 1 0 1000 0 -1 1648
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5672_6
timestamp 1731220634
transform 1 0 1040 0 1 1652
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5671_6
timestamp 1731220634
transform 1 0 912 0 1 1652
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5670_6
timestamp 1731220634
transform 1 0 976 0 1 1652
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5669_6
timestamp 1731220634
transform 1 0 984 0 -1 1760
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5668_6
timestamp 1731220634
transform 1 0 904 0 -1 1760
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5667_6
timestamp 1731220634
transform 1 0 824 0 -1 1760
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5666_6
timestamp 1731220634
transform 1 0 712 0 1 1652
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5665_6
timestamp 1731220634
transform 1 0 784 0 1 1652
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5664_6
timestamp 1731220634
transform 1 0 848 0 1 1652
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5663_6
timestamp 1731220634
transform 1 0 840 0 -1 1648
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5662_6
timestamp 1731220634
transform 1 0 784 0 -1 1648
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5661_6
timestamp 1731220634
transform 1 0 720 0 -1 1648
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5660_6
timestamp 1731220634
transform 1 0 736 0 1 1544
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5659_6
timestamp 1731220634
transform 1 0 664 0 1 1544
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5658_6
timestamp 1731220634
transform 1 0 592 0 1 1544
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5657_6
timestamp 1731220634
transform 1 0 520 0 1 1544
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5656_6
timestamp 1731220634
transform 1 0 560 0 -1 1544
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5655_6
timestamp 1731220634
transform 1 0 648 0 -1 1544
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5654_6
timestamp 1731220634
transform 1 0 736 0 -1 1544
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5653_6
timestamp 1731220634
transform 1 0 672 0 1 1440
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5652_6
timestamp 1731220634
transform 1 0 760 0 1 1440
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5651_6
timestamp 1731220634
transform 1 0 848 0 1 1440
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5650_6
timestamp 1731220634
transform 1 0 792 0 -1 1440
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5649_6
timestamp 1731220634
transform 1 0 880 0 -1 1440
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5648_6
timestamp 1731220634
transform 1 0 920 0 1 1336
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5647_6
timestamp 1731220634
transform 1 0 848 0 1 1336
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5646_6
timestamp 1731220634
transform 1 0 776 0 1 1336
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5645_6
timestamp 1731220634
transform 1 0 776 0 -1 1328
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5644_6
timestamp 1731220634
transform 1 0 856 0 -1 1328
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5643_6
timestamp 1731220634
transform 1 0 936 0 -1 1328
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5642_6
timestamp 1731220634
transform 1 0 1016 0 -1 1328
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5641_6
timestamp 1731220634
transform 1 0 1040 0 1 1220
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5640_6
timestamp 1731220634
transform 1 0 912 0 1 1220
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5639_6
timestamp 1731220634
transform 1 0 976 0 -1 1216
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5638_6
timestamp 1731220634
transform 1 0 936 0 1 1108
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5637_6
timestamp 1731220634
transform 1 0 992 0 -1 1108
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5636_6
timestamp 1731220634
transform 1 0 920 0 -1 1108
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5635_6
timestamp 1731220634
transform 1 0 568 0 1 1000
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5634_6
timestamp 1731220634
transform 1 0 504 0 1 1000
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5633_6
timestamp 1731220634
transform 1 0 520 0 -1 996
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5632_6
timestamp 1731220634
transform 1 0 464 0 -1 996
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5631_6
timestamp 1731220634
transform 1 0 448 0 1 888
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5630_6
timestamp 1731220634
transform 1 0 504 0 1 888
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5629_6
timestamp 1731220634
transform 1 0 560 0 1 888
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5628_6
timestamp 1731220634
transform 1 0 616 0 1 888
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5627_6
timestamp 1731220634
transform 1 0 616 0 -1 884
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5626_6
timestamp 1731220634
transform 1 0 544 0 -1 884
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5625_6
timestamp 1731220634
transform 1 0 472 0 -1 884
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5624_6
timestamp 1731220634
transform 1 0 480 0 1 780
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5623_6
timestamp 1731220634
transform 1 0 560 0 1 780
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5622_6
timestamp 1731220634
transform 1 0 640 0 1 780
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5621_6
timestamp 1731220634
transform 1 0 560 0 -1 780
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5620_6
timestamp 1731220634
transform 1 0 488 0 -1 780
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5619_6
timestamp 1731220634
transform 1 0 536 0 1 676
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5618_6
timestamp 1731220634
transform 1 0 464 0 1 676
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5617_6
timestamp 1731220634
transform 1 0 384 0 1 676
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5616_6
timestamp 1731220634
transform 1 0 392 0 -1 676
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5615_6
timestamp 1731220634
transform 1 0 456 0 -1 676
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5614_6
timestamp 1731220634
transform 1 0 328 0 -1 676
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5613_6
timestamp 1731220634
transform 1 0 296 0 1 564
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5612_6
timestamp 1731220634
transform 1 0 344 0 1 564
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5611_6
timestamp 1731220634
transform 1 0 392 0 1 564
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5610_6
timestamp 1731220634
transform 1 0 416 0 -1 560
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5609_6
timestamp 1731220634
transform 1 0 368 0 -1 560
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5608_6
timestamp 1731220634
transform 1 0 320 0 -1 560
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5607_6
timestamp 1731220634
transform 1 0 352 0 1 448
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5606_6
timestamp 1731220634
transform 1 0 416 0 1 448
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5605_6
timestamp 1731220634
transform 1 0 472 0 1 448
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5604_6
timestamp 1731220634
transform 1 0 528 0 -1 444
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5603_6
timestamp 1731220634
transform 1 0 456 0 -1 444
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5602_6
timestamp 1731220634
transform 1 0 320 0 -1 444
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5601_6
timestamp 1731220634
transform 1 0 384 0 -1 444
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5600_6
timestamp 1731220634
transform 1 0 400 0 1 332
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5599_6
timestamp 1731220634
transform 1 0 480 0 1 332
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5598_6
timestamp 1731220634
transform 1 0 560 0 1 332
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5597_6
timestamp 1731220634
transform 1 0 328 0 1 332
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5596_6
timestamp 1731220634
transform 1 0 264 0 1 332
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5595_6
timestamp 1731220634
transform 1 0 208 0 1 332
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5594_6
timestamp 1731220634
transform 1 0 168 0 1 332
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5593_6
timestamp 1731220634
transform 1 0 168 0 -1 444
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5592_6
timestamp 1731220634
transform 1 0 208 0 -1 444
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5591_6
timestamp 1731220634
transform 1 0 256 0 -1 444
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5590_6
timestamp 1731220634
transform 1 0 128 0 1 448
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5589_6
timestamp 1731220634
transform 1 0 168 0 1 448
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5588_6
timestamp 1731220634
transform 1 0 224 0 1 448
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5587_6
timestamp 1731220634
transform 1 0 288 0 1 448
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5586_6
timestamp 1731220634
transform 1 0 272 0 -1 560
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5585_6
timestamp 1731220634
transform 1 0 216 0 -1 560
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5584_6
timestamp 1731220634
transform 1 0 168 0 -1 560
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5583_6
timestamp 1731220634
transform 1 0 128 0 -1 560
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5582_6
timestamp 1731220634
transform 1 0 128 0 1 564
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5581_6
timestamp 1731220634
transform 1 0 168 0 1 564
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5580_6
timestamp 1731220634
transform 1 0 208 0 1 564
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5579_6
timestamp 1731220634
transform 1 0 248 0 1 564
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5578_6
timestamp 1731220634
transform 1 0 128 0 -1 676
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5577_6
timestamp 1731220634
transform 1 0 168 0 -1 676
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5576_6
timestamp 1731220634
transform 1 0 208 0 -1 676
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5575_6
timestamp 1731220634
transform 1 0 264 0 -1 676
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5574_6
timestamp 1731220634
transform 1 0 304 0 1 676
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5573_6
timestamp 1731220634
transform 1 0 232 0 1 676
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5572_6
timestamp 1731220634
transform 1 0 168 0 1 676
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5571_6
timestamp 1731220634
transform 1 0 208 0 -1 780
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5570_6
timestamp 1731220634
transform 1 0 272 0 -1 780
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5569_6
timestamp 1731220634
transform 1 0 344 0 -1 780
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5568_6
timestamp 1731220634
transform 1 0 416 0 -1 780
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5567_6
timestamp 1731220634
transform 1 0 408 0 1 780
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5566_6
timestamp 1731220634
transform 1 0 336 0 1 780
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5565_6
timestamp 1731220634
transform 1 0 272 0 1 780
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5564_6
timestamp 1731220634
transform 1 0 296 0 -1 884
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5563_6
timestamp 1731220634
transform 1 0 344 0 -1 884
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5562_6
timestamp 1731220634
transform 1 0 408 0 -1 884
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5561_6
timestamp 1731220634
transform 1 0 256 0 1 888
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5560_6
timestamp 1731220634
transform 1 0 296 0 1 888
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5559_6
timestamp 1731220634
transform 1 0 344 0 1 888
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5558_6
timestamp 1731220634
transform 1 0 392 0 1 888
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5557_6
timestamp 1731220634
transform 1 0 400 0 -1 996
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5556_6
timestamp 1731220634
transform 1 0 336 0 -1 996
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5555_6
timestamp 1731220634
transform 1 0 272 0 -1 996
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5554_6
timestamp 1731220634
transform 1 0 128 0 -1 996
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5553_6
timestamp 1731220634
transform 1 0 168 0 -1 996
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5552_6
timestamp 1731220634
transform 1 0 216 0 -1 996
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5551_6
timestamp 1731220634
transform 1 0 312 0 1 1000
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5550_6
timestamp 1731220634
transform 1 0 376 0 1 1000
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5549_6
timestamp 1731220634
transform 1 0 440 0 1 1000
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5548_6
timestamp 1731220634
transform 1 0 128 0 1 1000
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5547_6
timestamp 1731220634
transform 1 0 168 0 1 1000
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5546_6
timestamp 1731220634
transform 1 0 208 0 1 1000
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5545_6
timestamp 1731220634
transform 1 0 248 0 1 1000
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5544_6
timestamp 1731220634
transform 1 0 152 0 -1 1108
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5543_6
timestamp 1731220634
transform 1 0 192 0 -1 1108
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5542_6
timestamp 1731220634
transform 1 0 248 0 -1 1108
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5541_6
timestamp 1731220634
transform 1 0 312 0 -1 1108
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5540_6
timestamp 1731220634
transform 1 0 392 0 -1 1108
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5539_6
timestamp 1731220634
transform 1 0 472 0 -1 1108
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5538_6
timestamp 1731220634
transform 1 0 552 0 -1 1108
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5537_6
timestamp 1731220634
transform 1 0 392 0 1 1108
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5536_6
timestamp 1731220634
transform 1 0 432 0 1 1108
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5535_6
timestamp 1731220634
transform 1 0 472 0 1 1108
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5534_6
timestamp 1731220634
transform 1 0 520 0 1 1108
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5533_6
timestamp 1731220634
transform 1 0 568 0 1 1108
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5532_6
timestamp 1731220634
transform 1 0 616 0 1 1108
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5531_6
timestamp 1731220634
transform 1 0 488 0 -1 1216
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5530_6
timestamp 1731220634
transform 1 0 440 0 -1 1216
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5529_6
timestamp 1731220634
transform 1 0 392 0 -1 1216
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5528_6
timestamp 1731220634
transform 1 0 264 0 -1 1216
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5527_6
timestamp 1731220634
transform 1 0 304 0 -1 1216
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5526_6
timestamp 1731220634
transform 1 0 344 0 -1 1216
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5525_6
timestamp 1731220634
transform 1 0 392 0 1 1220
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5524_6
timestamp 1731220634
transform 1 0 312 0 1 1220
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5523_6
timestamp 1731220634
transform 1 0 248 0 1 1220
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5522_6
timestamp 1731220634
transform 1 0 128 0 1 1220
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5521_6
timestamp 1731220634
transform 1 0 168 0 1 1220
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5520_6
timestamp 1731220634
transform 1 0 208 0 1 1220
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5519_6
timestamp 1731220634
transform 1 0 248 0 -1 1328
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5518_6
timestamp 1731220634
transform 1 0 312 0 -1 1328
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5517_6
timestamp 1731220634
transform 1 0 208 0 -1 1328
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5516_6
timestamp 1731220634
transform 1 0 168 0 -1 1328
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5515_6
timestamp 1731220634
transform 1 0 128 0 -1 1328
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5514_6
timestamp 1731220634
transform 1 0 128 0 1 1336
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5513_6
timestamp 1731220634
transform 1 0 128 0 -1 1440
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5512_6
timestamp 1731220634
transform 1 0 128 0 1 1440
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5511_6
timestamp 1731220634
transform 1 0 192 0 1 1440
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5510_6
timestamp 1731220634
transform 1 0 128 0 -1 1544
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5509_6
timestamp 1731220634
transform 1 0 168 0 -1 1544
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5508_6
timestamp 1731220634
transform 1 0 224 0 1 1544
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5507_6
timestamp 1731220634
transform 1 0 168 0 1 1544
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5506_6
timestamp 1731220634
transform 1 0 128 0 1 1544
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5505_6
timestamp 1731220634
transform 1 0 128 0 -1 1648
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5504_6
timestamp 1731220634
transform 1 0 176 0 -1 1648
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5503_6
timestamp 1731220634
transform 1 0 128 0 1 1652
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5502_6
timestamp 1731220634
transform 1 0 192 0 1 1652
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5501_6
timestamp 1731220634
transform 1 0 272 0 1 1652
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5500_6
timestamp 1731220634
transform 1 0 288 0 -1 1760
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5499_6
timestamp 1731220634
transform 1 0 224 0 -1 1760
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5498_6
timestamp 1731220634
transform 1 0 264 0 1 1760
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5497_6
timestamp 1731220634
transform 1 0 208 0 1 1760
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5496_6
timestamp 1731220634
transform 1 0 144 0 1 1760
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5495_6
timestamp 1731220634
transform 1 0 192 0 -1 1872
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5494_6
timestamp 1731220634
transform 1 0 264 0 -1 1872
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5493_6
timestamp 1731220634
transform 1 0 128 0 -1 1872
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5492_6
timestamp 1731220634
transform 1 0 128 0 1 1876
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5491_6
timestamp 1731220634
transform 1 0 168 0 1 1876
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5490_6
timestamp 1731220634
transform 1 0 224 0 1 1876
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5489_6
timestamp 1731220634
transform 1 0 288 0 1 1876
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5488_6
timestamp 1731220634
transform 1 0 304 0 -1 1980
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5487_6
timestamp 1731220634
transform 1 0 240 0 -1 1980
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5486_6
timestamp 1731220634
transform 1 0 184 0 -1 1980
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5485_6
timestamp 1731220634
transform 1 0 184 0 1 1980
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5484_6
timestamp 1731220634
transform 1 0 224 0 1 1980
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5483_6
timestamp 1731220634
transform 1 0 280 0 1 1980
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5482_6
timestamp 1731220634
transform 1 0 344 0 1 1980
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5481_6
timestamp 1731220634
transform 1 0 416 0 1 1980
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5480_6
timestamp 1731220634
transform 1 0 488 0 1 1980
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5479_6
timestamp 1731220634
transform 1 0 568 0 1 1980
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5478_6
timestamp 1731220634
transform 1 0 512 0 -1 1980
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5477_6
timestamp 1731220634
transform 1 0 440 0 -1 1980
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5476_6
timestamp 1731220634
transform 1 0 368 0 -1 1980
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5475_6
timestamp 1731220634
transform 1 0 360 0 1 1876
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5474_6
timestamp 1731220634
transform 1 0 424 0 1 1876
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5473_6
timestamp 1731220634
transform 1 0 488 0 1 1876
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5472_6
timestamp 1731220634
transform 1 0 448 0 -1 1872
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5471_6
timestamp 1731220634
transform 1 0 328 0 -1 1872
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5470_6
timestamp 1731220634
transform 1 0 392 0 -1 1872
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5469_6
timestamp 1731220634
transform 1 0 424 0 1 1760
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5468_6
timestamp 1731220634
transform 1 0 376 0 1 1760
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5467_6
timestamp 1731220634
transform 1 0 320 0 1 1760
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5466_6
timestamp 1731220634
transform 1 0 344 0 -1 1760
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5465_6
timestamp 1731220634
transform 1 0 408 0 -1 1760
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5464_6
timestamp 1731220634
transform 1 0 472 0 -1 1760
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5463_6
timestamp 1731220634
transform 1 0 536 0 -1 1760
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5462_6
timestamp 1731220634
transform 1 0 544 0 1 1652
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5461_6
timestamp 1731220634
transform 1 0 456 0 1 1652
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5460_6
timestamp 1731220634
transform 1 0 360 0 1 1652
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5459_6
timestamp 1731220634
transform 1 0 256 0 -1 1648
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5458_6
timestamp 1731220634
transform 1 0 336 0 -1 1648
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5457_6
timestamp 1731220634
transform 1 0 416 0 -1 1648
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5456_6
timestamp 1731220634
transform 1 0 496 0 -1 1648
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5455_6
timestamp 1731220634
transform 1 0 448 0 1 1544
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5454_6
timestamp 1731220634
transform 1 0 368 0 1 1544
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5453_6
timestamp 1731220634
transform 1 0 296 0 1 1544
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5452_6
timestamp 1731220634
transform 1 0 224 0 -1 1544
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5451_6
timestamp 1731220634
transform 1 0 304 0 -1 1544
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5450_6
timestamp 1731220634
transform 1 0 384 0 -1 1544
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5449_6
timestamp 1731220634
transform 1 0 472 0 -1 1544
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5448_6
timestamp 1731220634
transform 1 0 352 0 1 1440
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5447_6
timestamp 1731220634
transform 1 0 272 0 1 1440
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5446_6
timestamp 1731220634
transform 1 0 256 0 -1 1440
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5445_6
timestamp 1731220634
transform 1 0 184 0 -1 1440
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5444_6
timestamp 1731220634
transform 1 0 168 0 1 1336
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5443_6
timestamp 1731220634
transform 1 0 232 0 1 1336
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5442_6
timestamp 1731220634
transform 1 0 384 0 -1 1328
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5441_6
timestamp 1731220634
transform 1 0 456 0 -1 1328
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5440_6
timestamp 1731220634
transform 1 0 296 0 1 1336
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5439_6
timestamp 1731220634
transform 1 0 360 0 1 1336
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5438_6
timestamp 1731220634
transform 1 0 432 0 1 1336
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5437_6
timestamp 1731220634
transform 1 0 496 0 1 1336
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5436_6
timestamp 1731220634
transform 1 0 472 0 -1 1440
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5435_6
timestamp 1731220634
transform 1 0 328 0 -1 1440
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5434_6
timestamp 1731220634
transform 1 0 400 0 -1 1440
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5433_6
timestamp 1731220634
transform 1 0 432 0 1 1440
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5432_6
timestamp 1731220634
transform 1 0 512 0 1 1440
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5431_6
timestamp 1731220634
transform 1 0 592 0 1 1440
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5430_6
timestamp 1731220634
transform 1 0 624 0 -1 1440
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5429_6
timestamp 1731220634
transform 1 0 704 0 -1 1440
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5428_6
timestamp 1731220634
transform 1 0 544 0 -1 1440
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5427_6
timestamp 1731220634
transform 1 0 568 0 1 1336
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5426_6
timestamp 1731220634
transform 1 0 640 0 1 1336
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5425_6
timestamp 1731220634
transform 1 0 704 0 1 1336
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5424_6
timestamp 1731220634
transform 1 0 696 0 -1 1328
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5423_6
timestamp 1731220634
transform 1 0 616 0 -1 1328
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5422_6
timestamp 1731220634
transform 1 0 536 0 -1 1328
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5421_6
timestamp 1731220634
transform 1 0 480 0 1 1220
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5420_6
timestamp 1731220634
transform 1 0 576 0 1 1220
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5419_6
timestamp 1731220634
transform 1 0 680 0 1 1220
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5418_6
timestamp 1731220634
transform 1 0 792 0 1 1220
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5417_6
timestamp 1731220634
transform 1 0 544 0 -1 1216
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5416_6
timestamp 1731220634
transform 1 0 600 0 -1 1216
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5415_6
timestamp 1731220634
transform 1 0 664 0 -1 1216
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5414_6
timestamp 1731220634
transform 1 0 736 0 -1 1216
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5413_6
timestamp 1731220634
transform 1 0 808 0 -1 1216
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5412_6
timestamp 1731220634
transform 1 0 888 0 -1 1216
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5411_6
timestamp 1731220634
transform 1 0 664 0 1 1108
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5410_6
timestamp 1731220634
transform 1 0 712 0 1 1108
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5409_6
timestamp 1731220634
transform 1 0 768 0 1 1108
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5408_6
timestamp 1731220634
transform 1 0 824 0 1 1108
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5407_6
timestamp 1731220634
transform 1 0 880 0 1 1108
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5406_6
timestamp 1731220634
transform 1 0 632 0 -1 1108
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5405_6
timestamp 1731220634
transform 1 0 704 0 -1 1108
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5404_6
timestamp 1731220634
transform 1 0 776 0 -1 1108
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5403_6
timestamp 1731220634
transform 1 0 848 0 -1 1108
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5402_6
timestamp 1731220634
transform 1 0 856 0 1 1000
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5401_6
timestamp 1731220634
transform 1 0 792 0 1 1000
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5400_6
timestamp 1731220634
transform 1 0 736 0 1 1000
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5399_6
timestamp 1731220634
transform 1 0 680 0 1 1000
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5398_6
timestamp 1731220634
transform 1 0 624 0 1 1000
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5397_6
timestamp 1731220634
transform 1 0 576 0 -1 996
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5396_6
timestamp 1731220634
transform 1 0 624 0 -1 996
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5395_6
timestamp 1731220634
transform 1 0 680 0 -1 996
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5394_6
timestamp 1731220634
transform 1 0 736 0 -1 996
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5393_6
timestamp 1731220634
transform 1 0 792 0 -1 996
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5392_6
timestamp 1731220634
transform 1 0 680 0 1 888
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5391_6
timestamp 1731220634
transform 1 0 744 0 1 888
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5390_6
timestamp 1731220634
transform 1 0 808 0 1 888
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5389_6
timestamp 1731220634
transform 1 0 872 0 1 888
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5388_6
timestamp 1731220634
transform 1 0 936 0 1 888
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5387_6
timestamp 1731220634
transform 1 0 688 0 -1 884
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5386_6
timestamp 1731220634
transform 1 0 760 0 -1 884
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5385_6
timestamp 1731220634
transform 1 0 824 0 -1 884
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5384_6
timestamp 1731220634
transform 1 0 880 0 -1 884
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5383_6
timestamp 1731220634
transform 1 0 720 0 1 780
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5382_6
timestamp 1731220634
transform 1 0 792 0 1 780
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5381_6
timestamp 1731220634
transform 1 0 936 0 -1 884
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5380_6
timestamp 1731220634
transform 1 0 1000 0 -1 884
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5379_6
timestamp 1731220634
transform 1 0 1040 0 -1 884
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5378_6
timestamp 1731220634
transform 1 0 1000 0 1 888
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5377_6
timestamp 1731220634
transform 1 0 1040 0 1 888
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5376_6
timestamp 1731220634
transform 1 0 1152 0 -1 960
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5375_6
timestamp 1731220634
transform 1 0 1200 0 -1 960
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5374_6
timestamp 1731220634
transform 1 0 1152 0 1 968
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5373_6
timestamp 1731220634
transform 1 0 1192 0 1 968
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5372_6
timestamp 1731220634
transform 1 0 1192 0 -1 1076
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5371_6
timestamp 1731220634
transform 1 0 1152 0 -1 1076
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5370_6
timestamp 1731220634
transform 1 0 1040 0 -1 1108
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5369_6
timestamp 1731220634
transform 1 0 1000 0 1 1108
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5368_6
timestamp 1731220634
transform 1 0 1040 0 1 1108
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5367_6
timestamp 1731220634
transform 1 0 1152 0 -1 1184
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5366_6
timestamp 1731220634
transform 1 0 1200 0 -1 1184
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5365_6
timestamp 1731220634
transform 1 0 1272 0 -1 1184
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5364_6
timestamp 1731220634
transform 1 0 1184 0 1 1076
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5363_6
timestamp 1731220634
transform 1 0 1264 0 1 1076
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5362_6
timestamp 1731220634
transform 1 0 1296 0 -1 1076
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5361_6
timestamp 1731220634
transform 1 0 1240 0 -1 1076
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5360_6
timestamp 1731220634
transform 1 0 1232 0 1 968
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5359_6
timestamp 1731220634
transform 1 0 1288 0 1 968
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5358_6
timestamp 1731220634
transform 1 0 1344 0 1 968
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5357_6
timestamp 1731220634
transform 1 0 1368 0 -1 960
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5356_6
timestamp 1731220634
transform 1 0 1280 0 -1 960
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5355_6
timestamp 1731220634
transform 1 0 1232 0 1 856
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5354_6
timestamp 1731220634
transform 1 0 1312 0 1 856
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5353_6
timestamp 1731220634
transform 1 0 1400 0 1 856
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5352_6
timestamp 1731220634
transform 1 0 1352 0 -1 856
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5351_6
timestamp 1731220634
transform 1 0 1240 0 -1 856
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5350_6
timestamp 1731220634
transform 1 0 1152 0 -1 856
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5349_6
timestamp 1731220634
transform 1 0 1152 0 1 752
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5348_6
timestamp 1731220634
transform 1 0 1040 0 1 780
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5347_6
timestamp 1731220634
transform 1 0 1040 0 -1 780
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5346_6
timestamp 1731220634
transform 1 0 1000 0 -1 780
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5345_6
timestamp 1731220634
transform 1 0 952 0 -1 780
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5344_6
timestamp 1731220634
transform 1 0 992 0 1 780
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5343_6
timestamp 1731220634
transform 1 0 920 0 1 780
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5342_6
timestamp 1731220634
transform 1 0 856 0 1 780
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5341_6
timestamp 1731220634
transform 1 0 904 0 -1 780
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5340_6
timestamp 1731220634
transform 1 0 856 0 -1 780
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5339_6
timestamp 1731220634
transform 1 0 808 0 -1 780
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5338_6
timestamp 1731220634
transform 1 0 632 0 -1 780
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5337_6
timestamp 1731220634
transform 1 0 696 0 -1 780
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5336_6
timestamp 1731220634
transform 1 0 752 0 -1 780
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5335_6
timestamp 1731220634
transform 1 0 792 0 1 676
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5334_6
timestamp 1731220634
transform 1 0 856 0 1 676
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5333_6
timestamp 1731220634
transform 1 0 920 0 1 676
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5332_6
timestamp 1731220634
transform 1 0 728 0 1 676
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5331_6
timestamp 1731220634
transform 1 0 608 0 1 676
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5330_6
timestamp 1731220634
transform 1 0 672 0 1 676
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5329_6
timestamp 1731220634
transform 1 0 696 0 -1 676
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5328_6
timestamp 1731220634
transform 1 0 752 0 -1 676
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5327_6
timestamp 1731220634
transform 1 0 816 0 -1 676
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5326_6
timestamp 1731220634
transform 1 0 640 0 -1 676
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5325_6
timestamp 1731220634
transform 1 0 520 0 -1 676
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5324_6
timestamp 1731220634
transform 1 0 584 0 -1 676
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5323_6
timestamp 1731220634
transform 1 0 624 0 1 564
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5322_6
timestamp 1731220634
transform 1 0 672 0 1 564
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5321_6
timestamp 1731220634
transform 1 0 720 0 1 564
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5320_6
timestamp 1731220634
transform 1 0 576 0 1 564
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5319_6
timestamp 1731220634
transform 1 0 528 0 1 564
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5318_6
timestamp 1731220634
transform 1 0 480 0 1 564
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5317_6
timestamp 1731220634
transform 1 0 432 0 1 564
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5316_6
timestamp 1731220634
transform 1 0 456 0 -1 560
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5315_6
timestamp 1731220634
transform 1 0 504 0 -1 560
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5314_6
timestamp 1731220634
transform 1 0 552 0 -1 560
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5313_6
timestamp 1731220634
transform 1 0 600 0 -1 560
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5312_6
timestamp 1731220634
transform 1 0 648 0 -1 560
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5311_6
timestamp 1731220634
transform 1 0 696 0 -1 560
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5310_6
timestamp 1731220634
transform 1 0 744 0 -1 560
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5309_6
timestamp 1731220634
transform 1 0 528 0 1 448
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5308_6
timestamp 1731220634
transform 1 0 584 0 1 448
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5307_6
timestamp 1731220634
transform 1 0 632 0 1 448
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5306_6
timestamp 1731220634
transform 1 0 680 0 1 448
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5305_6
timestamp 1731220634
transform 1 0 728 0 1 448
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5304_6
timestamp 1731220634
transform 1 0 784 0 1 448
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5303_6
timestamp 1731220634
transform 1 0 840 0 1 448
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5302_6
timestamp 1731220634
transform 1 0 600 0 -1 444
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5301_6
timestamp 1731220634
transform 1 0 672 0 -1 444
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5300_6
timestamp 1731220634
transform 1 0 736 0 -1 444
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5299_6
timestamp 1731220634
transform 1 0 800 0 -1 444
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5298_6
timestamp 1731220634
transform 1 0 864 0 -1 444
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5297_6
timestamp 1731220634
transform 1 0 936 0 -1 444
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5296_6
timestamp 1731220634
transform 1 0 632 0 1 332
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5295_6
timestamp 1731220634
transform 1 0 704 0 1 332
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5294_6
timestamp 1731220634
transform 1 0 768 0 1 332
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5293_6
timestamp 1731220634
transform 1 0 832 0 1 332
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5292_6
timestamp 1731220634
transform 1 0 888 0 1 332
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5291_6
timestamp 1731220634
transform 1 0 944 0 1 332
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5290_6
timestamp 1731220634
transform 1 0 1000 0 1 332
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5289_6
timestamp 1731220634
transform 1 0 920 0 -1 328
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5288_6
timestamp 1731220634
transform 1 0 960 0 -1 328
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5287_6
timestamp 1731220634
transform 1 0 1000 0 -1 328
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5286_6
timestamp 1731220634
transform 1 0 1040 0 -1 328
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5285_6
timestamp 1731220634
transform 1 0 1040 0 1 332
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5284_6
timestamp 1731220634
transform 1 0 1152 0 1 320
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5283_6
timestamp 1731220634
transform 1 0 1240 0 1 320
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5282_6
timestamp 1731220634
transform 1 0 1352 0 1 320
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5281_6
timestamp 1731220634
transform 1 0 1456 0 1 320
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5280_6
timestamp 1731220634
transform 1 0 1152 0 -1 428
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5279_6
timestamp 1731220634
transform 1 0 1192 0 -1 428
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5278_6
timestamp 1731220634
transform 1 0 1248 0 -1 428
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5277_6
timestamp 1731220634
transform 1 0 1328 0 -1 428
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5276_6
timestamp 1731220634
transform 1 0 1408 0 -1 428
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5275_6
timestamp 1731220634
transform 1 0 1496 0 -1 428
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5274_6
timestamp 1731220634
transform 1 0 1288 0 1 428
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5273_6
timestamp 1731220634
transform 1 0 1328 0 1 428
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5272_6
timestamp 1731220634
transform 1 0 1368 0 1 428
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5271_6
timestamp 1731220634
transform 1 0 1416 0 1 428
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5270_6
timestamp 1731220634
transform 1 0 1464 0 1 428
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5269_6
timestamp 1731220634
transform 1 0 1520 0 1 428
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5268_6
timestamp 1731220634
transform 1 0 1536 0 -1 532
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5267_6
timestamp 1731220634
transform 1 0 1496 0 -1 532
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5266_6
timestamp 1731220634
transform 1 0 1456 0 -1 532
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5265_6
timestamp 1731220634
transform 1 0 1416 0 -1 532
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5264_6
timestamp 1731220634
transform 1 0 1296 0 -1 532
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5263_6
timestamp 1731220634
transform 1 0 1336 0 -1 532
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5262_6
timestamp 1731220634
transform 1 0 1376 0 -1 532
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5261_6
timestamp 1731220634
transform 1 0 1408 0 1 536
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5260_6
timestamp 1731220634
transform 1 0 1352 0 1 536
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5259_6
timestamp 1731220634
transform 1 0 1312 0 1 536
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5258_6
timestamp 1731220634
transform 1 0 1272 0 1 536
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5257_6
timestamp 1731220634
transform 1 0 1232 0 1 536
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5256_6
timestamp 1731220634
transform 1 0 1192 0 1 536
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5255_6
timestamp 1731220634
transform 1 0 1152 0 1 536
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5254_6
timestamp 1731220634
transform 1 0 1152 0 -1 644
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5253_6
timestamp 1731220634
transform 1 0 1192 0 -1 644
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5252_6
timestamp 1731220634
transform 1 0 1232 0 -1 644
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5251_6
timestamp 1731220634
transform 1 0 1272 0 -1 644
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5250_6
timestamp 1731220634
transform 1 0 1336 0 -1 644
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5249_6
timestamp 1731220634
transform 1 0 1408 0 -1 644
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5248_6
timestamp 1731220634
transform 1 0 1240 0 1 644
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5247_6
timestamp 1731220634
transform 1 0 1280 0 1 644
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5246_6
timestamp 1731220634
transform 1 0 1328 0 1 644
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5245_6
timestamp 1731220634
transform 1 0 1384 0 1 644
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5244_6
timestamp 1731220634
transform 1 0 1440 0 1 644
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5243_6
timestamp 1731220634
transform 1 0 1504 0 1 644
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5242_6
timestamp 1731220634
transform 1 0 1328 0 -1 748
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5241_6
timestamp 1731220634
transform 1 0 1368 0 -1 748
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5240_6
timestamp 1731220634
transform 1 0 1408 0 -1 748
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5239_6
timestamp 1731220634
transform 1 0 1448 0 -1 748
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5238_6
timestamp 1731220634
transform 1 0 1496 0 -1 748
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5237_6
timestamp 1731220634
transform 1 0 1544 0 -1 748
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5236_6
timestamp 1731220634
transform 1 0 1592 0 -1 748
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5235_6
timestamp 1731220634
transform 1 0 1272 0 1 752
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5234_6
timestamp 1731220634
transform 1 0 1400 0 1 752
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5233_6
timestamp 1731220634
transform 1 0 1448 0 -1 856
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5232_6
timestamp 1731220634
transform 1 0 1488 0 1 856
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5231_6
timestamp 1731220634
transform 1 0 1576 0 1 856
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5230_6
timestamp 1731220634
transform 1 0 1528 0 -1 960
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5229_6
timestamp 1731220634
transform 1 0 1448 0 -1 960
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5228_6
timestamp 1731220634
transform 1 0 1456 0 1 968
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5227_6
timestamp 1731220634
transform 1 0 1400 0 1 968
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5226_6
timestamp 1731220634
transform 1 0 1392 0 -1 1076
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5225_6
timestamp 1731220634
transform 1 0 1344 0 -1 1076
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5224_6
timestamp 1731220634
transform 1 0 1336 0 1 1076
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5223_6
timestamp 1731220634
transform 1 0 1344 0 -1 1184
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5222_6
timestamp 1731220634
transform 1 0 1416 0 -1 1184
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5221_6
timestamp 1731220634
transform 1 0 1480 0 -1 1184
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5220_6
timestamp 1731220634
transform 1 0 1488 0 1 1184
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5219_6
timestamp 1731220634
transform 1 0 1552 0 1 1184
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5218_6
timestamp 1731220634
transform 1 0 1424 0 1 1184
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5217_6
timestamp 1731220634
transform 1 0 1280 0 1 1184
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5216_6
timestamp 1731220634
transform 1 0 1320 0 1 1184
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5215_6
timestamp 1731220634
transform 1 0 1368 0 1 1184
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5214_6
timestamp 1731220634
transform 1 0 1384 0 -1 1292
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5213_6
timestamp 1731220634
transform 1 0 1472 0 -1 1292
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5212_6
timestamp 1731220634
transform 1 0 1560 0 -1 1292
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5211_6
timestamp 1731220634
transform 1 0 1168 0 -1 1292
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5210_6
timestamp 1731220634
transform 1 0 1224 0 -1 1292
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5209_6
timestamp 1731220634
transform 1 0 1296 0 -1 1292
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5208_6
timestamp 1731220634
transform 1 0 1304 0 1 1292
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5207_6
timestamp 1731220634
transform 1 0 1216 0 1 1292
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5206_6
timestamp 1731220634
transform 1 0 1152 0 1 1292
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5205_6
timestamp 1731220634
transform 1 0 1040 0 1 1336
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5204_6
timestamp 1731220634
transform 1 0 992 0 1 1336
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5203_6
timestamp 1731220634
transform 1 0 968 0 -1 1440
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5202_6
timestamp 1731220634
transform 1 0 1040 0 -1 1440
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5201_6
timestamp 1731220634
transform 1 0 1024 0 1 1440
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5200_6
timestamp 1731220634
transform 1 0 936 0 1 1440
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5199_6
timestamp 1731220634
transform 1 0 992 0 -1 1544
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5198_6
timestamp 1731220634
transform 1 0 904 0 -1 1544
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5197_6
timestamp 1731220634
transform 1 0 816 0 -1 1544
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5196_6
timestamp 1731220634
transform 1 0 880 0 1 1544
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5195_6
timestamp 1731220634
transform 1 0 808 0 1 1544
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5194_6
timestamp 1731220634
transform 1 0 648 0 -1 1648
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5193_6
timestamp 1731220634
transform 1 0 576 0 -1 1648
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5192_6
timestamp 1731220634
transform 1 0 632 0 1 1652
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5191_6
timestamp 1731220634
transform 1 0 608 0 -1 1760
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5190_6
timestamp 1731220634
transform 1 0 680 0 -1 1760
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5189_6
timestamp 1731220634
transform 1 0 752 0 -1 1760
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5188_6
timestamp 1731220634
transform 1 0 720 0 1 1760
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5187_6
timestamp 1731220634
transform 1 0 664 0 1 1760
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5186_6
timestamp 1731220634
transform 1 0 472 0 1 1760
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5185_6
timestamp 1731220634
transform 1 0 520 0 1 1760
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5184_6
timestamp 1731220634
transform 1 0 568 0 1 1760
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5183_6
timestamp 1731220634
transform 1 0 616 0 1 1760
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5182_6
timestamp 1731220634
transform 1 0 496 0 -1 1872
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5181_6
timestamp 1731220634
transform 1 0 544 0 -1 1872
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5180_6
timestamp 1731220634
transform 1 0 592 0 -1 1872
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5179_6
timestamp 1731220634
transform 1 0 640 0 -1 1872
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5178_6
timestamp 1731220634
transform 1 0 688 0 -1 1872
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5177_6
timestamp 1731220634
transform 1 0 744 0 -1 1872
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5176_6
timestamp 1731220634
transform 1 0 552 0 1 1876
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5175_6
timestamp 1731220634
transform 1 0 608 0 1 1876
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5174_6
timestamp 1731220634
transform 1 0 664 0 1 1876
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5173_6
timestamp 1731220634
transform 1 0 720 0 1 1876
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5172_6
timestamp 1731220634
transform 1 0 776 0 1 1876
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5171_6
timestamp 1731220634
transform 1 0 840 0 1 1876
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5170_6
timestamp 1731220634
transform 1 0 584 0 -1 1980
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5169_6
timestamp 1731220634
transform 1 0 648 0 -1 1980
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5168_6
timestamp 1731220634
transform 1 0 712 0 -1 1980
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5167_6
timestamp 1731220634
transform 1 0 768 0 -1 1980
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5166_6
timestamp 1731220634
transform 1 0 816 0 -1 1980
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5165_6
timestamp 1731220634
transform 1 0 864 0 -1 1980
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5164_6
timestamp 1731220634
transform 1 0 640 0 1 1980
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5163_6
timestamp 1731220634
transform 1 0 712 0 1 1980
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5162_6
timestamp 1731220634
transform 1 0 776 0 1 1980
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5161_6
timestamp 1731220634
transform 1 0 832 0 1 1980
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5160_6
timestamp 1731220634
transform 1 0 888 0 1 1980
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5159_6
timestamp 1731220634
transform 1 0 944 0 1 1980
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5158_6
timestamp 1731220634
transform 1 0 1000 0 1 1980
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5157_6
timestamp 1731220634
transform 1 0 1040 0 1 1980
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5156_6
timestamp 1731220634
transform 1 0 912 0 -1 1980
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5155_6
timestamp 1731220634
transform 1 0 960 0 -1 1980
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5154_6
timestamp 1731220634
transform 1 0 1000 0 -1 1980
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5153_6
timestamp 1731220634
transform 1 0 1040 0 -1 1980
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5152_6
timestamp 1731220634
transform 1 0 1152 0 -1 1944
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5151_6
timestamp 1731220634
transform 1 0 1216 0 -1 1944
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5150_6
timestamp 1731220634
transform 1 0 1152 0 1 1836
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5149_6
timestamp 1731220634
transform 1 0 1192 0 1 1836
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5148_6
timestamp 1731220634
transform 1 0 1256 0 1 1836
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5147_6
timestamp 1731220634
transform 1 0 1296 0 -1 1836
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5146_6
timestamp 1731220634
transform 1 0 1224 0 -1 1836
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5145_6
timestamp 1731220634
transform 1 0 1152 0 -1 1836
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5144_6
timestamp 1731220634
transform 1 0 1184 0 1 1732
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5143_6
timestamp 1731220634
transform 1 0 1248 0 1 1732
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5142_6
timestamp 1731220634
transform 1 0 1312 0 1 1732
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5141_6
timestamp 1731220634
transform 1 0 1336 0 -1 1732
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5140_6
timestamp 1731220634
transform 1 0 1288 0 -1 1732
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5139_6
timestamp 1731220634
transform 1 0 1240 0 -1 1732
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5138_6
timestamp 1731220634
transform 1 0 1256 0 1 1624
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5137_6
timestamp 1731220634
transform 1 0 1296 0 1 1624
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5136_6
timestamp 1731220634
transform 1 0 1336 0 1 1624
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5135_6
timestamp 1731220634
transform 1 0 1384 0 1 1624
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5134_6
timestamp 1731220634
transform 1 0 1440 0 1 1624
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5133_6
timestamp 1731220634
transform 1 0 1496 0 1 1624
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5132_6
timestamp 1731220634
transform 1 0 1520 0 -1 1732
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5131_6
timestamp 1731220634
transform 1 0 1456 0 -1 1732
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5130_6
timestamp 1731220634
transform 1 0 1392 0 -1 1732
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5129_6
timestamp 1731220634
transform 1 0 1376 0 1 1732
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5128_6
timestamp 1731220634
transform 1 0 1448 0 1 1732
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5127_6
timestamp 1731220634
transform 1 0 1520 0 1 1732
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5126_6
timestamp 1731220634
transform 1 0 1544 0 -1 1836
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5125_6
timestamp 1731220634
transform 1 0 1456 0 -1 1836
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5124_6
timestamp 1731220634
transform 1 0 1376 0 -1 1836
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5123_6
timestamp 1731220634
transform 1 0 1320 0 1 1836
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5122_6
timestamp 1731220634
transform 1 0 1384 0 1 1836
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5121_6
timestamp 1731220634
transform 1 0 1440 0 1 1836
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5120_6
timestamp 1731220634
transform 1 0 1456 0 -1 1944
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5119_6
timestamp 1731220634
transform 1 0 1376 0 -1 1944
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5118_6
timestamp 1731220634
transform 1 0 1296 0 -1 1944
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5117_6
timestamp 1731220634
transform 1 0 1296 0 1 1948
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5116_6
timestamp 1731220634
transform 1 0 1376 0 1 1948
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5115_6
timestamp 1731220634
transform 1 0 1456 0 1 1948
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5114_6
timestamp 1731220634
transform 1 0 1536 0 1 1948
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5113_6
timestamp 1731220634
transform 1 0 1576 0 -1 2052
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5112_6
timestamp 1731220634
transform 1 0 1480 0 -1 2052
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5111_6
timestamp 1731220634
transform 1 0 1392 0 -1 2052
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5110_6
timestamp 1731220634
transform 1 0 1304 0 -1 2052
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5109_6
timestamp 1731220634
transform 1 0 1232 0 -1 2052
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5108_6
timestamp 1731220634
transform 1 0 1176 0 -1 2052
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5107_6
timestamp 1731220634
transform 1 0 1216 0 1 2052
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5106_6
timestamp 1731220634
transform 1 0 1272 0 1 2052
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5105_6
timestamp 1731220634
transform 1 0 1336 0 1 2052
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5104_6
timestamp 1731220634
transform 1 0 1416 0 1 2052
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5103_6
timestamp 1731220634
transform 1 0 1496 0 1 2052
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5102_6
timestamp 1731220634
transform 1 0 1576 0 1 2052
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5101_6
timestamp 1731220634
transform 1 0 1280 0 -1 2160
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5100_6
timestamp 1731220634
transform 1 0 1320 0 -1 2160
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_599_6
timestamp 1731220634
transform 1 0 1360 0 -1 2160
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_598_6
timestamp 1731220634
transform 1 0 1408 0 -1 2160
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_597_6
timestamp 1731220634
transform 1 0 1456 0 -1 2160
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_596_6
timestamp 1731220634
transform 1 0 1512 0 -1 2160
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_595_6
timestamp 1731220634
transform 1 0 1568 0 -1 2160
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_594_6
timestamp 1731220634
transform 1 0 1336 0 1 2160
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_593_6
timestamp 1731220634
transform 1 0 1376 0 1 2160
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_592_6
timestamp 1731220634
transform 1 0 1416 0 1 2160
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_591_6
timestamp 1731220634
transform 1 0 1456 0 1 2160
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_590_6
timestamp 1731220634
transform 1 0 1496 0 1 2160
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_589_6
timestamp 1731220634
transform 1 0 1536 0 1 2160
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_588_6
timestamp 1731220634
transform 1 0 1576 0 1 2160
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_587_6
timestamp 1731220634
transform 1 0 1616 0 1 2160
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_586_6
timestamp 1731220634
transform 1 0 1656 0 1 2160
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_585_6
timestamp 1731220634
transform 1 0 1696 0 1 2160
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_584_6
timestamp 1731220634
transform 1 0 1736 0 1 2160
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_583_6
timestamp 1731220634
transform 1 0 1776 0 1 2160
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_582_6
timestamp 1731220634
transform 1 0 1816 0 1 2160
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_581_6
timestamp 1731220634
transform 1 0 1616 0 -1 2160
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_580_6
timestamp 1731220634
transform 1 0 1664 0 -1 2160
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_579_6
timestamp 1731220634
transform 1 0 1712 0 -1 2160
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_578_6
timestamp 1731220634
transform 1 0 1768 0 -1 2160
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_577_6
timestamp 1731220634
transform 1 0 1824 0 -1 2160
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_576_6
timestamp 1731220634
transform 1 0 1880 0 -1 2160
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_575_6
timestamp 1731220634
transform 1 0 1656 0 1 2052
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_574_6
timestamp 1731220634
transform 1 0 1736 0 1 2052
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_573_6
timestamp 1731220634
transform 1 0 1824 0 1 2052
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_572_6
timestamp 1731220634
transform 1 0 1912 0 1 2052
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_571_6
timestamp 1731220634
transform 1 0 2000 0 1 2052
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_570_6
timestamp 1731220634
transform 1 0 2000 0 -1 2052
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_569_6
timestamp 1731220634
transform 1 0 1912 0 -1 2052
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_568_6
timestamp 1731220634
transform 1 0 1832 0 -1 2052
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_567_6
timestamp 1731220634
transform 1 0 1664 0 -1 2052
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_566_6
timestamp 1731220634
transform 1 0 1752 0 -1 2052
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_565_6
timestamp 1731220634
transform 1 0 1808 0 1 1948
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_564_6
timestamp 1731220634
transform 1 0 1872 0 1 1948
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_563_6
timestamp 1731220634
transform 1 0 1944 0 1 1948
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_562_6
timestamp 1731220634
transform 1 0 1608 0 1 1948
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_561_6
timestamp 1731220634
transform 1 0 1680 0 1 1948
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_560_6
timestamp 1731220634
transform 1 0 1744 0 1 1948
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_559_6
timestamp 1731220634
transform 1 0 1776 0 -1 1944
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_558_6
timestamp 1731220634
transform 1 0 1872 0 -1 1944
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_557_6
timestamp 1731220634
transform 1 0 1976 0 -1 1944
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_556_6
timestamp 1731220634
transform 1 0 1528 0 -1 1944
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_555_6
timestamp 1731220634
transform 1 0 1608 0 -1 1944
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_554_6
timestamp 1731220634
transform 1 0 1688 0 -1 1944
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_553_6
timestamp 1731220634
transform 1 0 1704 0 1 1836
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_552_6
timestamp 1731220634
transform 1 0 1792 0 1 1836
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_551_6
timestamp 1731220634
transform 1 0 1888 0 1 1836
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_550_6
timestamp 1731220634
transform 1 0 1496 0 1 1836
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_549_6
timestamp 1731220634
transform 1 0 1552 0 1 1836
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_548_6
timestamp 1731220634
transform 1 0 1624 0 1 1836
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_547_6
timestamp 1731220634
transform 1 0 1640 0 -1 1836
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_546_6
timestamp 1731220634
transform 1 0 1744 0 -1 1836
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_545_6
timestamp 1731220634
transform 1 0 1680 0 1 1732
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_544_6
timestamp 1731220634
transform 1 0 1600 0 1 1732
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_543_6
timestamp 1731220634
transform 1 0 1664 0 -1 1732
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_542_6
timestamp 1731220634
transform 1 0 1592 0 -1 1732
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_541_6
timestamp 1731220634
transform 1 0 1560 0 1 1624
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_540_6
timestamp 1731220634
transform 1 0 1624 0 1 1624
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_539_6
timestamp 1731220634
transform 1 0 1616 0 -1 1612
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_538_6
timestamp 1731220634
transform 1 0 1456 0 -1 1612
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_537_6
timestamp 1731220634
transform 1 0 1536 0 -1 1612
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_536_6
timestamp 1731220634
transform 1 0 1552 0 1 1508
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_535_6
timestamp 1731220634
transform 1 0 1640 0 1 1508
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_534_6
timestamp 1731220634
transform 1 0 1728 0 1 1508
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_533_6
timestamp 1731220634
transform 1 0 1792 0 -1 1612
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_532_6
timestamp 1731220634
transform 1 0 1880 0 -1 1612
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_531_6
timestamp 1731220634
transform 1 0 1704 0 -1 1612
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_530_6
timestamp 1731220634
transform 1 0 1688 0 1 1624
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_529_6
timestamp 1731220634
transform 1 0 1752 0 1 1624
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_528_6
timestamp 1731220634
transform 1 0 1824 0 1 1624
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_527_6
timestamp 1731220634
transform 1 0 1904 0 1 1624
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_526_6
timestamp 1731220634
transform 1 0 1872 0 -1 1732
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_525_6
timestamp 1731220634
transform 1 0 1800 0 -1 1732
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_524_6
timestamp 1731220634
transform 1 0 1736 0 -1 1732
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_523_6
timestamp 1731220634
transform 1 0 1760 0 1 1732
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_522_6
timestamp 1731220634
transform 1 0 1840 0 1 1732
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_521_6
timestamp 1731220634
transform 1 0 1920 0 1 1732
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_520_6
timestamp 1731220634
transform 1 0 1848 0 -1 1836
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_519_6
timestamp 1731220634
transform 1 0 1960 0 -1 1836
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_518_6
timestamp 1731220634
transform 1 0 2000 0 1 1732
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_517_6
timestamp 1731220634
transform 1 0 1944 0 -1 1732
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_516_6
timestamp 1731220634
transform 1 0 1992 0 1 1624
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_515_6
timestamp 1731220634
transform 1 0 1976 0 -1 1612
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_514_6
timestamp 1731220634
transform 1 0 1912 0 -1 1508
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_513_6
timestamp 1731220634
transform 1 0 2064 0 1 1508
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_512_6
timestamp 1731220634
transform 1 0 2064 0 -1 1612
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_511_6
timestamp 1731220634
transform 1 0 2064 0 1 1624
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_510_6
timestamp 1731220634
transform 1 0 2016 0 -1 1732
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_59_6
timestamp 1731220634
transform 1 0 2064 0 -1 1732
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_58_6
timestamp 1731220634
transform 1 0 2064 0 1 1732
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_57_6
timestamp 1731220634
transform 1 0 2064 0 -1 1836
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_56_6
timestamp 1731220634
transform 1 0 1984 0 1 1836
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_55_6
timestamp 1731220634
transform 1 0 2064 0 1 1836
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_54_6
timestamp 1731220634
transform 1 0 2064 0 -1 1944
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_53_6
timestamp 1731220634
transform 1 0 2016 0 1 1948
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_52_6
timestamp 1731220634
transform 1 0 2064 0 1 1948
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_51_6
timestamp 1731220634
transform 1 0 2064 0 -1 2052
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_50_6
timestamp 1731220634
transform 1 0 2064 0 1 2052
box 4 6 36 48
<< end >>
