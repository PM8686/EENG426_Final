magic
tech sky130l
timestamp 1730254790
<< ndiffusion >>
rect 8 27 13 32
rect 8 24 9 27
rect 12 24 13 27
rect 8 22 13 24
rect 15 26 22 32
rect 15 23 17 26
rect 20 23 22 26
rect 15 22 22 23
rect 24 22 29 32
rect 31 30 36 32
rect 31 27 32 30
rect 35 27 36 30
rect 31 22 36 27
rect 38 27 43 32
rect 38 24 39 27
rect 42 24 43 27
rect 38 22 43 24
rect 45 30 52 32
rect 45 27 47 30
rect 50 27 52 30
rect 45 22 52 27
rect 48 12 52 22
rect 54 24 59 32
rect 54 21 55 24
rect 58 21 59 24
rect 54 12 59 21
rect 61 30 68 32
rect 61 27 63 30
rect 66 27 68 30
rect 61 12 68 27
rect 70 24 75 32
rect 70 21 71 24
rect 74 21 75 24
rect 70 12 75 21
rect 77 23 84 32
rect 77 20 80 23
rect 83 20 84 23
rect 77 12 84 20
rect 86 12 89 32
rect 91 12 94 32
rect 96 30 101 32
rect 96 27 97 30
rect 100 27 101 30
rect 96 26 101 27
rect 103 31 108 32
rect 103 28 104 31
rect 107 28 108 31
rect 103 26 108 28
rect 114 30 119 32
rect 114 27 115 30
rect 118 27 119 30
rect 114 26 119 27
rect 121 31 126 32
rect 121 28 122 31
rect 125 28 126 31
rect 121 26 126 28
rect 96 12 100 26
<< ndc >>
rect 9 24 12 27
rect 17 23 20 26
rect 32 27 35 30
rect 39 24 42 27
rect 47 27 50 30
rect 55 21 58 24
rect 63 27 66 30
rect 71 21 74 24
rect 80 20 83 23
rect 97 27 100 30
rect 104 28 107 31
rect 115 27 118 30
rect 122 28 125 31
<< ntransistor >>
rect 13 22 15 32
rect 22 22 24 32
rect 29 22 31 32
rect 36 22 38 32
rect 43 22 45 32
rect 52 12 54 32
rect 59 12 61 32
rect 68 12 70 32
rect 75 12 77 32
rect 84 12 86 32
rect 89 12 91 32
rect 94 12 96 32
rect 101 26 103 32
rect 119 26 121 32
<< pdiffusion >>
rect 64 75 68 79
rect 48 62 52 75
rect 18 50 22 62
rect 8 44 13 50
rect 8 41 9 44
rect 12 41 13 44
rect 8 39 13 41
rect 15 49 22 50
rect 15 46 16 49
rect 19 46 22 49
rect 15 39 22 46
rect 24 43 29 62
rect 24 40 25 43
rect 28 40 29 43
rect 24 39 29 40
rect 31 49 36 62
rect 31 46 32 49
rect 35 46 36 49
rect 31 39 36 46
rect 38 39 43 62
rect 45 44 52 62
rect 45 41 47 44
rect 50 41 52 44
rect 45 39 52 41
rect 54 50 59 75
rect 54 47 55 50
rect 58 47 59 50
rect 54 39 59 47
rect 61 44 68 75
rect 61 41 63 44
rect 66 41 68 44
rect 61 39 68 41
rect 70 75 74 79
rect 80 75 84 87
rect 70 50 75 75
rect 70 47 71 50
rect 74 47 75 50
rect 70 39 75 47
rect 77 43 84 75
rect 77 40 80 43
rect 83 40 84 43
rect 77 39 84 40
rect 86 39 89 87
rect 91 39 94 87
rect 96 47 100 87
rect 96 44 101 47
rect 96 41 97 44
rect 100 41 101 44
rect 96 39 101 41
rect 103 46 108 47
rect 103 43 104 46
rect 107 43 108 46
rect 103 39 108 43
rect 114 46 119 47
rect 114 43 115 46
rect 118 43 119 46
rect 114 39 119 43
rect 121 44 126 47
rect 121 41 122 44
rect 125 41 126 44
rect 121 39 126 41
<< pdc >>
rect 9 41 12 44
rect 16 46 19 49
rect 25 40 28 43
rect 32 46 35 49
rect 47 41 50 44
rect 55 47 58 50
rect 63 41 66 44
rect 71 47 74 50
rect 80 40 83 43
rect 97 41 100 44
rect 104 43 107 46
rect 115 43 118 46
rect 122 41 125 44
<< ptransistor >>
rect 13 39 15 50
rect 22 39 24 62
rect 29 39 31 62
rect 36 39 38 62
rect 43 39 45 62
rect 52 39 54 75
rect 59 39 61 75
rect 68 39 70 79
rect 75 39 77 75
rect 84 39 86 87
rect 89 39 91 87
rect 94 39 96 87
rect 101 39 103 47
rect 119 39 121 47
<< polysilicon >>
rect 29 97 34 98
rect 29 94 30 97
rect 33 94 34 97
rect 29 93 34 94
rect 43 97 48 98
rect 43 94 44 97
rect 47 94 48 97
rect 43 93 48 94
rect 68 97 73 98
rect 68 94 69 97
rect 72 94 73 97
rect 68 93 73 94
rect 80 97 85 98
rect 80 94 81 97
rect 84 94 85 97
rect 21 89 26 90
rect 21 86 22 89
rect 25 86 26 89
rect 21 85 26 86
rect 13 81 19 82
rect 13 78 15 81
rect 18 78 19 81
rect 13 77 19 78
rect 13 50 15 77
rect 22 62 24 85
rect 29 62 31 93
rect 35 89 40 90
rect 35 86 36 89
rect 39 86 40 89
rect 35 85 40 86
rect 36 62 38 85
rect 43 62 45 93
rect 49 89 54 90
rect 49 86 50 89
rect 53 86 54 89
rect 49 85 54 86
rect 52 75 54 85
rect 57 86 62 87
rect 57 83 58 86
rect 61 83 62 86
rect 57 82 62 83
rect 59 75 61 82
rect 68 79 70 93
rect 80 90 85 94
rect 88 97 93 98
rect 88 94 89 97
rect 92 94 93 97
rect 88 93 93 94
rect 96 97 101 98
rect 96 94 97 97
rect 100 94 101 97
rect 80 88 86 90
rect 84 87 86 88
rect 89 87 91 93
rect 96 90 101 94
rect 94 88 101 90
rect 94 87 96 88
rect 75 75 77 77
rect 101 47 103 49
rect 119 47 121 49
rect 13 32 15 39
rect 22 32 24 39
rect 29 32 31 39
rect 36 32 38 39
rect 43 32 45 39
rect 52 32 54 39
rect 59 32 61 39
rect 68 32 70 39
rect 75 32 77 39
rect 84 32 86 39
rect 89 32 91 39
rect 94 32 96 39
rect 101 32 103 39
rect 119 32 121 39
rect 13 20 15 22
rect 22 20 24 22
rect 29 20 31 22
rect 36 20 38 22
rect 43 20 45 22
rect 52 10 54 12
rect 59 10 61 12
rect 68 10 70 12
rect 75 10 77 12
rect 84 10 86 12
rect 89 10 91 12
rect 94 10 96 12
rect 101 10 103 26
rect 119 24 121 26
rect 116 23 121 24
rect 116 20 117 23
rect 120 20 121 23
rect 116 19 121 20
rect 75 9 80 10
rect 75 6 76 9
rect 79 6 80 9
rect 75 5 80 6
rect 101 9 106 10
rect 101 6 102 9
rect 105 6 106 9
rect 101 5 106 6
<< pc >>
rect 30 94 33 97
rect 44 94 47 97
rect 69 94 72 97
rect 81 94 84 97
rect 22 86 25 89
rect 15 78 18 81
rect 36 86 39 89
rect 50 86 53 89
rect 58 83 61 86
rect 89 94 92 97
rect 97 94 100 97
rect 117 20 120 23
rect 76 6 79 9
rect 102 6 105 9
<< m1 >>
rect 8 97 12 98
rect 8 94 9 97
rect 8 72 12 94
rect 30 97 33 98
rect 30 93 33 94
rect 44 97 47 98
rect 44 93 47 94
rect 69 97 72 98
rect 69 93 72 94
rect 81 97 84 98
rect 22 89 25 90
rect 22 85 25 86
rect 36 89 39 90
rect 36 85 39 86
rect 50 89 53 90
rect 64 89 68 90
rect 50 85 53 86
rect 58 86 61 87
rect 15 81 18 82
rect 15 77 18 78
rect 58 81 61 83
rect 58 77 61 78
rect 67 86 68 89
rect 64 72 68 86
rect 72 81 76 82
rect 75 78 76 81
rect 72 72 76 78
rect 81 81 84 94
rect 89 97 92 98
rect 89 89 92 94
rect 97 97 100 98
rect 97 93 100 94
rect 81 77 84 78
rect 8 44 12 52
rect 15 46 16 49
rect 19 46 32 49
rect 35 46 36 49
rect 54 47 55 50
rect 58 47 71 50
rect 74 47 75 50
rect 104 46 108 52
rect 8 41 9 44
rect 47 44 50 45
rect 97 44 100 45
rect 8 40 12 41
rect 24 40 25 43
rect 28 40 29 43
rect 62 41 63 44
rect 66 41 67 44
rect 80 43 83 44
rect 47 40 50 41
rect 97 40 100 41
rect 107 43 108 46
rect 9 27 12 28
rect 9 23 12 24
rect 9 19 12 20
rect 17 26 20 27
rect 17 9 20 23
rect 17 5 20 6
rect 24 9 29 40
rect 32 30 35 31
rect 47 30 50 31
rect 32 16 35 27
rect 39 27 42 28
rect 62 27 63 30
rect 66 27 67 30
rect 47 26 50 27
rect 39 23 42 24
rect 54 21 55 24
rect 58 21 71 24
rect 74 21 75 24
rect 80 23 83 40
rect 104 31 108 43
rect 112 46 118 52
rect 112 43 115 46
rect 112 37 118 43
rect 122 44 125 45
rect 122 40 125 41
rect 112 34 125 37
rect 122 31 125 34
rect 97 30 100 31
rect 107 28 108 31
rect 104 27 108 28
rect 115 30 118 31
rect 122 27 125 28
rect 97 26 100 27
rect 115 26 118 27
rect 39 19 42 20
rect 116 20 117 23
rect 120 20 121 23
rect 80 19 83 20
rect 32 12 36 16
rect 24 6 25 9
rect 28 6 29 9
rect 75 6 76 9
rect 79 6 80 9
rect 101 6 102 9
rect 105 6 106 9
rect 24 5 29 6
<< m2c >>
rect 9 94 12 97
rect 30 94 33 97
rect 44 94 47 97
rect 69 94 72 97
rect 22 86 25 89
rect 36 86 39 89
rect 50 86 53 89
rect 15 78 18 81
rect 58 78 61 81
rect 64 86 67 89
rect 72 78 75 81
rect 97 94 100 97
rect 89 86 92 89
rect 81 78 84 81
rect 9 41 12 44
rect 47 41 50 44
rect 63 41 66 44
rect 97 41 100 44
rect 9 20 12 23
rect 17 6 20 9
rect 32 27 35 30
rect 47 27 50 30
rect 63 27 66 30
rect 39 20 42 23
rect 122 41 125 44
rect 97 27 100 30
rect 115 27 118 30
rect 80 20 83 23
rect 117 20 120 23
rect 25 6 28 9
rect 76 6 79 9
rect 102 6 105 9
<< m2 >>
rect 8 97 101 98
rect 8 94 9 97
rect 12 94 30 97
rect 33 94 44 97
rect 47 94 69 97
rect 72 94 97 97
rect 100 94 101 97
rect 8 93 101 94
rect 21 89 93 90
rect 21 86 22 89
rect 25 86 36 89
rect 39 86 50 89
rect 53 86 64 89
rect 67 86 89 89
rect 92 86 93 89
rect 21 85 93 86
rect 14 81 85 82
rect 14 78 15 81
rect 18 78 58 81
rect 61 78 72 81
rect 75 78 81 81
rect 84 78 85 81
rect 14 77 85 78
rect 8 44 126 45
rect 8 41 9 44
rect 12 41 47 44
rect 50 41 63 44
rect 66 41 97 44
rect 100 41 122 44
rect 125 41 126 44
rect 8 40 126 41
rect 31 30 119 31
rect 31 27 32 30
rect 35 27 47 30
rect 50 27 63 30
rect 66 27 97 30
rect 100 27 115 30
rect 118 27 119 30
rect 31 26 119 27
rect 8 23 43 24
rect 8 20 9 23
rect 12 20 39 23
rect 42 20 43 23
rect 8 19 43 20
rect 79 23 121 24
rect 79 20 80 23
rect 83 20 117 23
rect 120 20 121 23
rect 79 19 121 20
rect 16 9 106 10
rect 16 6 17 9
rect 20 6 25 9
rect 28 6 76 9
rect 79 6 102 9
rect 105 6 106 9
rect 16 5 106 6
<< labels >>
rlabel m2 s 100 94 101 97 6 A
port 1 nsew signal input
rlabel m2 s 97 94 100 97 6 A
port 1 nsew signal input
rlabel m2 s 72 94 97 97 6 A
port 1 nsew signal input
rlabel m2 s 69 94 72 97 6 A
port 1 nsew signal input
rlabel m2 s 47 94 69 97 6 A
port 1 nsew signal input
rlabel m2 s 44 94 47 97 6 A
port 1 nsew signal input
rlabel m2 s 33 94 44 97 6 A
port 1 nsew signal input
rlabel m2 s 30 94 33 97 6 A
port 1 nsew signal input
rlabel m2 s 12 94 30 97 6 A
port 1 nsew signal input
rlabel m2 s 9 94 12 97 6 A
port 1 nsew signal input
rlabel m2 s 8 93 101 94 6 A
port 1 nsew signal input
rlabel m2 s 8 94 9 97 6 A
port 1 nsew signal input
rlabel m2 s 8 97 101 98 6 A
port 1 nsew signal input
rlabel m2c s 97 94 100 97 6 A
port 1 nsew signal input
rlabel m2c s 69 94 72 97 6 A
port 1 nsew signal input
rlabel m2c s 44 94 47 97 6 A
port 1 nsew signal input
rlabel m2c s 30 94 33 97 6 A
port 1 nsew signal input
rlabel m2c s 9 94 12 97 6 A
port 1 nsew signal input
rlabel m1 s 97 93 100 94 6 A
port 1 nsew signal input
rlabel m1 s 97 94 100 97 6 A
port 1 nsew signal input
rlabel m1 s 97 97 100 98 6 A
port 1 nsew signal input
rlabel m1 s 69 93 72 94 6 A
port 1 nsew signal input
rlabel m1 s 69 94 72 97 6 A
port 1 nsew signal input
rlabel m1 s 69 97 72 98 6 A
port 1 nsew signal input
rlabel m1 s 44 93 47 94 6 A
port 1 nsew signal input
rlabel m1 s 44 94 47 97 6 A
port 1 nsew signal input
rlabel m1 s 44 97 47 98 6 A
port 1 nsew signal input
rlabel m1 s 30 93 33 94 6 A
port 1 nsew signal input
rlabel m1 s 30 94 33 97 6 A
port 1 nsew signal input
rlabel m1 s 30 97 33 98 6 A
port 1 nsew signal input
rlabel m1 s 9 94 12 97 6 A
port 1 nsew signal input
rlabel m1 s 8 72 12 94 6 A
port 1 nsew signal input
rlabel m1 s 8 94 9 97 6 A
port 1 nsew signal input
rlabel m1 s 8 97 12 98 6 A
port 1 nsew signal input
rlabel m2 s 92 86 93 89 6 B
port 2 nsew signal input
rlabel m2 s 89 86 92 89 6 B
port 2 nsew signal input
rlabel m2 s 67 86 89 89 6 B
port 2 nsew signal input
rlabel m2 s 64 86 67 89 6 B
port 2 nsew signal input
rlabel m2 s 53 86 64 89 6 B
port 2 nsew signal input
rlabel m2 s 50 86 53 89 6 B
port 2 nsew signal input
rlabel m2 s 39 86 50 89 6 B
port 2 nsew signal input
rlabel m2 s 36 86 39 89 6 B
port 2 nsew signal input
rlabel m2 s 25 86 36 89 6 B
port 2 nsew signal input
rlabel m2 s 22 86 25 89 6 B
port 2 nsew signal input
rlabel m2 s 21 85 93 86 6 B
port 2 nsew signal input
rlabel m2 s 21 86 22 89 6 B
port 2 nsew signal input
rlabel m2 s 21 89 93 90 6 B
port 2 nsew signal input
rlabel m2c s 89 86 92 89 6 B
port 2 nsew signal input
rlabel m2c s 64 86 67 89 6 B
port 2 nsew signal input
rlabel m2c s 50 86 53 89 6 B
port 2 nsew signal input
rlabel m2c s 36 86 39 89 6 B
port 2 nsew signal input
rlabel m2c s 22 86 25 89 6 B
port 2 nsew signal input
rlabel m1 s 89 86 92 89 6 B
port 2 nsew signal input
rlabel m1 s 89 89 92 94 6 B
port 2 nsew signal input
rlabel m1 s 89 94 92 97 6 B
port 2 nsew signal input
rlabel m1 s 89 97 92 98 6 B
port 2 nsew signal input
rlabel m1 s 67 86 68 89 6 B
port 2 nsew signal input
rlabel m1 s 64 72 68 86 6 B
port 2 nsew signal input
rlabel m1 s 64 86 67 89 6 B
port 2 nsew signal input
rlabel m1 s 64 89 68 90 6 B
port 2 nsew signal input
rlabel m1 s 36 85 39 86 6 B
port 2 nsew signal input
rlabel m1 s 36 86 39 89 6 B
port 2 nsew signal input
rlabel m1 s 36 89 39 90 6 B
port 2 nsew signal input
rlabel m1 s 50 85 53 86 6 B
port 2 nsew signal input
rlabel m1 s 50 86 53 89 6 B
port 2 nsew signal input
rlabel m1 s 50 89 53 90 6 B
port 2 nsew signal input
rlabel m1 s 22 85 25 86 6 B
port 2 nsew signal input
rlabel m1 s 22 86 25 89 6 B
port 2 nsew signal input
rlabel m1 s 22 89 25 90 6 B
port 2 nsew signal input
rlabel m2 s 84 78 85 81 6 C
port 3 nsew signal input
rlabel m2 s 81 78 84 81 6 C
port 3 nsew signal input
rlabel m2 s 75 78 81 81 6 C
port 3 nsew signal input
rlabel m2 s 72 78 75 81 6 C
port 3 nsew signal input
rlabel m2 s 61 78 72 81 6 C
port 3 nsew signal input
rlabel m2 s 58 78 61 81 6 C
port 3 nsew signal input
rlabel m2 s 18 78 58 81 6 C
port 3 nsew signal input
rlabel m2 s 15 78 18 81 6 C
port 3 nsew signal input
rlabel m2 s 14 77 85 78 6 C
port 3 nsew signal input
rlabel m2 s 14 78 15 81 6 C
port 3 nsew signal input
rlabel m2 s 14 81 85 82 6 C
port 3 nsew signal input
rlabel m2c s 81 78 84 81 6 C
port 3 nsew signal input
rlabel m2c s 72 78 75 81 6 C
port 3 nsew signal input
rlabel m2c s 58 78 61 81 6 C
port 3 nsew signal input
rlabel m2c s 15 78 18 81 6 C
port 3 nsew signal input
rlabel m1 s 81 78 84 81 6 C
port 3 nsew signal input
rlabel m1 s 81 77 84 78 6 C
port 3 nsew signal input
rlabel m1 s 81 81 84 94 6 C
port 3 nsew signal input
rlabel m1 s 81 94 84 97 6 C
port 3 nsew signal input
rlabel m1 s 81 97 84 98 6 C
port 3 nsew signal input
rlabel m1 s 75 78 76 81 6 C
port 3 nsew signal input
rlabel m1 s 72 72 76 78 6 C
port 3 nsew signal input
rlabel m1 s 72 78 75 81 6 C
port 3 nsew signal input
rlabel m1 s 72 81 76 82 6 C
port 3 nsew signal input
rlabel m1 s 58 77 61 78 6 C
port 3 nsew signal input
rlabel m1 s 58 78 61 81 6 C
port 3 nsew signal input
rlabel m1 s 58 81 61 83 6 C
port 3 nsew signal input
rlabel m1 s 58 83 61 86 6 C
port 3 nsew signal input
rlabel m1 s 58 86 61 87 6 C
port 3 nsew signal input
rlabel m1 s 15 77 18 78 6 C
port 3 nsew signal input
rlabel m1 s 15 78 18 81 6 C
port 3 nsew signal input
rlabel m1 s 15 81 18 82 6 C
port 3 nsew signal input
rlabel m1 s 107 28 108 31 6 YC
port 4 nsew signal output
rlabel m1 s 107 43 108 46 6 YC
port 4 nsew signal output
rlabel m1 s 104 27 108 28 6 YC
port 4 nsew signal output
rlabel m1 s 104 28 107 31 6 YC
port 4 nsew signal output
rlabel m1 s 104 31 108 43 6 YC
port 4 nsew signal output
rlabel m1 s 104 43 107 46 6 YC
port 4 nsew signal output
rlabel m1 s 104 46 108 52 6 YC
port 4 nsew signal output
rlabel m1 s 122 27 125 28 6 YS
port 5 nsew signal output
rlabel m1 s 122 28 125 31 6 YS
port 5 nsew signal output
rlabel m1 s 122 31 125 34 6 YS
port 5 nsew signal output
rlabel m1 s 115 43 118 46 6 YS
port 5 nsew signal output
rlabel m1 s 112 43 115 46 6 YS
port 5 nsew signal output
rlabel m1 s 112 34 125 37 6 YS
port 5 nsew signal output
rlabel m1 s 112 37 118 43 6 YS
port 5 nsew signal output
rlabel m1 s 112 46 118 52 6 YS
port 5 nsew signal output
rlabel m2 s 125 41 126 44 6 Vdd
port 6 nsew power input
rlabel m2 s 122 41 125 44 6 Vdd
port 6 nsew power input
rlabel m2 s 100 41 122 44 6 Vdd
port 6 nsew power input
rlabel m2 s 97 41 100 44 6 Vdd
port 6 nsew power input
rlabel m2 s 66 41 97 44 6 Vdd
port 6 nsew power input
rlabel m2 s 63 41 66 44 6 Vdd
port 6 nsew power input
rlabel m2 s 50 41 63 44 6 Vdd
port 6 nsew power input
rlabel m2 s 47 41 50 44 6 Vdd
port 6 nsew power input
rlabel m2 s 12 41 47 44 6 Vdd
port 6 nsew power input
rlabel m2 s 9 41 12 44 6 Vdd
port 6 nsew power input
rlabel m2 s 8 40 126 41 6 Vdd
port 6 nsew power input
rlabel m2 s 8 41 9 44 6 Vdd
port 6 nsew power input
rlabel m2 s 8 44 126 45 6 Vdd
port 6 nsew power input
rlabel m2c s 122 41 125 44 6 Vdd
port 6 nsew power input
rlabel m2c s 97 41 100 44 6 Vdd
port 6 nsew power input
rlabel m2c s 63 41 66 44 6 Vdd
port 6 nsew power input
rlabel m2c s 47 41 50 44 6 Vdd
port 6 nsew power input
rlabel m2c s 9 41 12 44 6 Vdd
port 6 nsew power input
rlabel m1 s 122 40 125 41 6 Vdd
port 6 nsew power input
rlabel m1 s 122 41 125 44 6 Vdd
port 6 nsew power input
rlabel m1 s 122 44 125 45 6 Vdd
port 6 nsew power input
rlabel m1 s 97 40 100 41 6 Vdd
port 6 nsew power input
rlabel m1 s 97 41 100 44 6 Vdd
port 6 nsew power input
rlabel m1 s 97 44 100 45 6 Vdd
port 6 nsew power input
rlabel m1 s 66 41 67 44 6 Vdd
port 6 nsew power input
rlabel m1 s 63 41 66 44 6 Vdd
port 6 nsew power input
rlabel m1 s 62 41 63 44 6 Vdd
port 6 nsew power input
rlabel m1 s 47 40 50 41 6 Vdd
port 6 nsew power input
rlabel m1 s 47 41 50 44 6 Vdd
port 6 nsew power input
rlabel m1 s 47 44 50 45 6 Vdd
port 6 nsew power input
rlabel m1 s 9 41 12 44 6 Vdd
port 6 nsew power input
rlabel m1 s 8 40 12 41 6 Vdd
port 6 nsew power input
rlabel m1 s 8 41 9 44 6 Vdd
port 6 nsew power input
rlabel m1 s 8 44 12 52 6 Vdd
port 6 nsew power input
rlabel m2 s 118 27 119 30 6 GND
port 7 nsew ground input
rlabel m2 s 115 27 118 30 6 GND
port 7 nsew ground input
rlabel m2 s 100 27 115 30 6 GND
port 7 nsew ground output
rlabel m2 s 97 27 100 30 6 GND
port 7 nsew ground output
rlabel m2 s 66 27 97 30 6 GND
port 7 nsew ground output
rlabel m2 s 63 27 66 30 6 GND
port 7 nsew ground output
rlabel m2 s 50 27 63 30 6 GND
port 7 nsew ground output
rlabel m2 s 47 27 50 30 6 GND
port 7 nsew ground output
rlabel m2 s 35 27 47 30 6 GND
port 7 nsew ground output
rlabel m2 s 32 27 35 30 6 GND
port 7 nsew ground output
rlabel m2 s 31 26 119 27 6 GND
port 7 nsew ground output
rlabel m2 s 31 27 32 30 6 GND
port 7 nsew ground output
rlabel m2 s 31 30 119 31 6 GND
port 7 nsew ground output
rlabel m2c s 115 27 118 30 6 GND
port 7 nsew ground output
rlabel m2c s 97 27 100 30 6 GND
port 7 nsew ground output
rlabel m2c s 63 27 66 30 6 GND
port 7 nsew ground output
rlabel m2c s 47 27 50 30 6 GND
port 7 nsew ground output
rlabel m2c s 32 27 35 30 6 GND
port 7 nsew ground output
rlabel m1 s 115 30 118 31 6 GND
port 7 nsew ground output
rlabel m1 s 115 27 118 30 6 GND
port 7 nsew ground output
rlabel m1 s 115 26 118 27 6 GND
port 7 nsew ground output
rlabel m1 s 97 26 100 27 6 GND
port 7 nsew ground output
rlabel m1 s 97 27 100 30 6 GND
port 7 nsew ground output
rlabel m1 s 97 30 100 31 6 GND
port 7 nsew ground output
rlabel m1 s 66 27 67 30 6 GND
port 7 nsew ground output
rlabel m1 s 63 27 66 30 6 GND
port 7 nsew ground output
rlabel m1 s 62 27 63 30 6 GND
port 7 nsew ground output
rlabel m1 s 47 27 50 30 6 GND
port 7 nsew ground output
rlabel m1 s 47 30 50 31 6 GND
port 7 nsew ground output
rlabel m1 s 47 26 50 27 6 GND
port 7 nsew ground output
rlabel m1 s 32 12 36 16 6 GND
port 7 nsew ground output
rlabel m1 s 32 16 35 27 6 GND
port 7 nsew ground output
rlabel m1 s 32 27 35 30 6 GND
port 7 nsew ground output
rlabel m1 s 32 30 35 31 6 GND
port 7 nsew ground output
rlabel space 0 0 136 100 1 prboundary
rlabel polysilicon 102 33 102 33 3 _YC
rlabel polysilicon 95 33 95 33 3 A
rlabel polysilicon 90 33 90 33 3 B
rlabel polysilicon 97 91 97 91 3 A
rlabel polysilicon 97 95 97 95 3 A
rlabel polysilicon 97 98 97 98 3 A
rlabel polysilicon 85 33 85 33 3 C
rlabel polysilicon 95 88 95 88 3 A
rlabel polysilicon 95 89 95 89 3 A
rlabel pdiffusion 104 40 104 40 3 YC
rlabel pdiffusion 104 44 104 44 3 YC
rlabel pdiffusion 104 47 104 47 3 YC
rlabel polysilicon 102 48 102 48 3 _YC
rlabel polysilicon 69 80 69 80 3 A
rlabel polysilicon 69 94 69 94 3 A
rlabel polysilicon 69 95 69 95 3 A
rlabel polysilicon 69 98 69 98 3 A
rlabel ptransistor 102 40 102 40 3 _YC
rlabel polysilicon 93 95 93 95 3 B
rlabel pdiffusion 65 76 65 76 3 Vdd
rlabel ndiffusion 126 29 126 29 3 YS
rlabel pdiffusion 97 40 97 40 3 Vdd
rlabel pdiffusion 97 42 97 42 3 Vdd
rlabel pdiffusion 97 45 97 45 3 Vdd
rlabel pdiffusion 97 48 97 48 3 Vdd
rlabel polysilicon 90 88 90 88 3 B
rlabel polysilicon 62 84 62 84 3 C
rlabel polysilicon 76 33 76 33 3 _YC
rlabel ptransistor 95 40 95 40 3 A
rlabel polysilicon 89 94 89 94 3 B
rlabel polysilicon 89 95 89 95 3 B
rlabel polysilicon 89 98 89 98 3 B
rlabel polysilicon 60 76 60 76 3 C
rlabel ndiffusion 122 27 122 27 3 YS
rlabel ndiffusion 122 29 122 29 3 YS
rlabel ndiffusion 122 32 122 32 3 YS
rlabel ndiffusion 115 31 115 31 3 GND
rlabel pdiffusion 122 40 122 40 3 Vdd
rlabel pdiffusion 122 42 122 42 3 Vdd
rlabel pdiffusion 122 45 122 45 3 Vdd
rlabel pdiffusion 119 44 119 44 3 YS
rlabel polysilicon 85 95 85 95 3 C
rlabel polysilicon 58 83 58 83 3 C
rlabel polysilicon 58 84 58 84 3 C
rlabel polysilicon 58 87 58 87 3 C
rlabel ntransistor 120 27 120 27 3 _YS
rlabel polysilicon 120 33 120 33 3 _YS
rlabel ptransistor 120 40 120 40 3 _YS
rlabel polysilicon 120 48 120 48 3 _YS
rlabel polysilicon 69 33 69 33 3 A
rlabel ptransistor 90 40 90 40 3 B
rlabel polysilicon 85 88 85 88 3 C
rlabel ndiffusion 115 27 115 27 3 GND
rlabel ndiffusion 115 28 115 28 3 GND
rlabel pdiffusion 115 40 115 40 3 YS
rlabel pdiffusion 115 44 115 44 3 YS
rlabel pdiffusion 115 47 115 47 3 YS
rlabel pdiffusion 84 41 84 41 3 _YS
rlabel pdiffusion 81 76 81 76 3 _YS
rlabel polysilicon 81 89 81 89 3 C
rlabel polysilicon 81 91 81 91 3 C
rlabel polysilicon 81 95 81 95 3 C
rlabel polysilicon 81 98 81 98 3 C
rlabel polysilicon 53 76 53 76 3 B
rlabel polysilicon 117 20 117 20 3 _YS
rlabel polysilicon 117 24 117 24 3 _YS
rlabel polysilicon 120 25 120 25 3 _YS
rlabel ptransistor 85 40 85 40 3 C
rlabel polysilicon 50 86 50 86 3 B
rlabel polysilicon 50 87 50 87 3 B
rlabel polysilicon 50 90 50 90 3 B
rlabel ndiffusion 104 27 104 27 3 YC
rlabel ndiffusion 104 29 104 29 3 YC
rlabel ndiffusion 104 32 104 32 3 YC
rlabel pdiffusion 78 40 78 40 3 _YS
rlabel pdiffusion 78 41 78 41 3 _YS
rlabel pdiffusion 78 44 78 44 3 _YS
rlabel polysilicon 76 76 76 76 3 _YC
rlabel pdiffusion 49 63 49 63 3 Vdd
rlabel polysilicon 102 11 102 11 3 _YC
rlabel ntransistor 102 27 102 27 3 _YC
rlabel polysilicon 60 33 60 33 3 C
rlabel ptransistor 76 40 76 40 3 _YC
rlabel ndiffusion 97 13 97 13 3 GND
rlabel ndiffusion 97 27 97 27 3 GND
rlabel ndiffusion 97 28 97 28 3 GND
rlabel ndiffusion 97 31 97 31 3 GND
rlabel pdiffusion 71 40 71 40 3 #12
rlabel pdiffusion 71 48 71 48 3 #12
rlabel pdiffusion 71 51 71 51 3 #12
rlabel pdiffusion 71 76 71 76 3 #12
rlabel polysilicon 95 11 95 11 3 A
rlabel ntransistor 95 13 95 13 3 A
rlabel polysilicon 53 33 53 33 3 B
rlabel ptransistor 69 40 69 40 3 A
rlabel polysilicon 44 63 44 63 3 A
rlabel pdiffusion 62 40 62 40 3 Vdd
rlabel pdiffusion 62 42 62 42 3 Vdd
rlabel pdiffusion 62 45 62 45 3 Vdd
rlabel polysilicon 90 11 90 11 3 B
rlabel ntransistor 90 13 90 13 3 B
rlabel ptransistor 60 40 60 40 3 C
rlabel polysilicon 44 94 44 94 3 A
rlabel polysilicon 44 95 44 95 3 A
rlabel polysilicon 44 98 44 98 3 A
rlabel pdiffusion 55 40 55 40 3 #12
rlabel pdiffusion 55 51 55 51 3 #12
rlabel polysilicon 37 63 37 63 3 B
rlabel polysilicon 85 11 85 11 3 C
rlabel ntransistor 85 13 85 13 3 C
rlabel polysilicon 44 33 44 33 3 A
rlabel ptransistor 53 40 53 40 3 B
rlabel polysilicon 36 86 36 86 3 B
rlabel polysilicon 36 87 36 87 3 B
rlabel polysilicon 36 90 36 90 3 B
rlabel ndiffusion 78 13 78 13 3 _YS
rlabel ndiffusion 78 21 78 21 3 _YS
rlabel ndiffusion 78 24 78 24 3 _YS
rlabel ndiffusion 46 23 46 23 3 GND
rlabel ndiffusion 46 28 46 28 3 GND
rlabel ndiffusion 46 31 46 31 3 GND
rlabel ndiffusion 43 25 43 25 3 #3
rlabel pdiffusion 46 40 46 40 3 Vdd
rlabel pdiffusion 46 42 46 42 3 Vdd
rlabel pdiffusion 46 45 46 45 3 Vdd
rlabel polysilicon 76 11 76 11 3 _YC
rlabel ntransistor 76 13 76 13 3 _YC
rlabel polysilicon 44 21 44 21 3 A
rlabel ntransistor 44 23 44 23 3 A
rlabel polysilicon 37 33 37 33 3 B
rlabel ptransistor 44 40 44 40 3 A
rlabel ndiffusion 71 13 71 13 3 #15
rlabel ndiffusion 71 22 71 22 3 #15
rlabel ndiffusion 71 25 71 25 3 #15
rlabel ndiffusion 39 23 39 23 3 #3
rlabel ndiffusion 39 25 39 25 3 #3
rlabel ndiffusion 39 28 39 28 3 #3
rlabel polysilicon 30 63 30 63 3 A
rlabel polysilicon 69 11 69 11 3 A
rlabel ntransistor 69 13 69 13 3 A
rlabel polysilicon 37 21 37 21 3 B
rlabel ntransistor 37 23 37 23 3 B
rlabel polysilicon 30 33 30 33 3 A
rlabel ptransistor 37 40 37 40 3 B
rlabel polysilicon 102 6 102 6 3 _YC
rlabel polysilicon 102 10 102 10 3 _YC
rlabel ndiffusion 62 13 62 13 3 GND
rlabel ndiffusion 62 28 62 28 3 GND
rlabel ndiffusion 62 31 62 31 3 GND
rlabel ndiffusion 32 23 32 23 3 GND
rlabel pdiffusion 32 40 32 40 3 #8
rlabel pdiffusion 32 47 32 47 3 #8
rlabel pdiffusion 32 50 32 50 3 #8
rlabel polysilicon 60 11 60 11 3 C
rlabel ntransistor 60 13 60 13 3 C
rlabel polysilicon 30 21 30 21 3 A
rlabel ntransistor 30 23 30 23 3 A
rlabel polysilicon 23 33 23 33 3 B
rlabel ptransistor 30 40 30 40 3 A
rlabel polysilicon 23 63 23 63 3 B
rlabel polysilicon 30 94 30 94 3 A
rlabel polysilicon 30 95 30 95 3 A
rlabel polysilicon 30 98 30 98 3 A
rlabel polysilicon 76 6 76 6 3 _YC
rlabel polysilicon 76 10 76 10 3 _YC
rlabel ndiffusion 55 13 55 13 3 #15
rlabel ndiffusion 55 25 55 25 3 #15
rlabel ndiffusion 21 24 21 24 3 _YC
rlabel pdiffusion 25 40 25 40 3 _YC
rlabel pdiffusion 25 44 25 44 3 _YC
rlabel polysilicon 53 11 53 11 3 B
rlabel ntransistor 53 13 53 13 3 B
rlabel polysilicon 23 21 23 21 3 B
rlabel ntransistor 23 23 23 23 3 B
rlabel ptransistor 23 40 23 40 3 B
rlabel pdiffusion 19 51 19 51 3 #8
rlabel ndiffusion 49 13 49 13 3 GND
rlabel ndiffusion 16 23 16 23 3 _YC
rlabel ndiffusion 16 24 16 24 3 _YC
rlabel ndiffusion 16 27 16 27 3 _YC
rlabel ndiffusion 13 25 13 25 3 #3
rlabel pdiffusion 16 40 16 40 3 #8
rlabel pdiffusion 16 50 16 50 3 #8
rlabel polysilicon 14 21 14 21 3 C
rlabel ntransistor 14 23 14 23 3 C
rlabel polysilicon 14 33 14 33 3 C
rlabel ptransistor 14 40 14 40 3 C
rlabel polysilicon 14 51 14 51 3 C
rlabel polysilicon 14 78 14 78 3 C
rlabel polysilicon 14 79 14 79 3 C
rlabel polysilicon 14 82 14 82 3 C
rlabel ndiffusion 9 23 9 23 3 #3
rlabel ndiffusion 9 25 9 25 3 #3
rlabel ndiffusion 9 28 9 28 3 #3
rlabel pdiffusion 9 40 9 40 3 Vdd
rlabel m1 98 94 98 94 3 A
port 1 e default input
rlabel m1 98 98 98 98 3 A
port 1 e default input
rlabel m1 90 90 90 90 3 B
port 2 e default input
rlabel pc 90 95 90 95 3 B
port 2 e default input
rlabel m1 90 98 90 98 3 B
port 2 e default input
rlabel m1 82 78 82 78 3 C
port 3 e default input
rlabel m1 82 82 82 82 3 C
port 3 e default input
rlabel pc 82 95 82 95 3 C
port 3 e default input
rlabel m1 82 98 82 98 3 C
port 3 e default input
rlabel m1 123 28 123 28 3 YS
port 5 e default output
rlabel ndc 123 29 123 29 3 YS
port 5 e default output
rlabel m1 123 32 123 32 3 YS
port 5 e default output
rlabel m1 123 41 123 41 3 Vdd
rlabel m1 123 45 123 45 3 Vdd
rlabel pdc 116 44 116 44 3 YS
port 5 e default output
rlabel m1 98 41 98 41 3 Vdd
rlabel m1 98 45 98 45 3 Vdd
rlabel m1 116 31 116 31 3 GND
rlabel m1 113 44 113 44 3 YS
port 5 e default output
rlabel m1 73 73 73 73 3 C
port 3 e default input
rlabel m1 73 82 73 82 3 C
port 3 e default input
rlabel m1 113 35 113 35 3 YS
port 5 e default output
rlabel m1 113 38 113 38 3 YS
port 5 e default output
rlabel m1 113 47 113 47 3 YS
port 5 e
rlabel pdc 81 41 81 41 3 _YS
rlabel m1 81 44 81 44 3 _YS
rlabel m1 108 29 108 29 3 YC
port 4 e default output
rlabel m1 108 44 108 44 3 YC
port 4 e default output
rlabel m1 116 27 116 27 3 GND
rlabel m1 105 28 105 28 3 YC
port 4 e default output
rlabel ndc 105 29 105 29 3 YC
port 4 e default output
rlabel m1 105 32 105 32 3 YC
port 4 e default output
rlabel pdc 105 44 105 44 3 YC
port 4 e default output
rlabel m1 105 47 105 47 3 YC
port 4 e
rlabel m1 70 94 70 94 3 A
port 1 e default input
rlabel m1 70 98 70 98 3 A
port 1 e default input
rlabel m1 98 27 98 27 3 GND
rlabel m1 98 31 98 31 3 GND
rlabel m1 75 48 75 48 3 #12
rlabel m1 65 73 65 73 3 B
port 2 e default input
rlabel m1 65 90 65 90 3 B
port 2 e default input
rlabel pdc 72 48 72 48 3 #12
rlabel m1 81 24 81 24 3 _YS
rlabel m1 63 28 63 28 3 GND
rlabel m1 63 42 63 42 3 Vdd
rlabel m1 59 48 59 48 3 #12
rlabel m1 59 78 59 78 3 C
port 3 e default input
rlabel m1 59 82 59 82 3 C
port 3 e default input
rlabel pc 59 84 59 84 3 C
port 3 e default input
rlabel m1 59 87 59 87 3 C
port 3 e default input
rlabel m1 45 94 45 94 3 A
port 1 e default input
rlabel m1 45 98 45 98 3 A
port 1 e default input
rlabel pdc 56 48 56 48 3 #12
rlabel m1 75 22 75 22 3 #15
rlabel m1 55 48 55 48 3 #12
rlabel m1 37 86 37 86 3 B
port 2 e default input
rlabel m1 37 90 37 90 3 B
port 2 e default input
rlabel ndc 72 22 72 22 3 #15
rlabel m1 51 86 51 86 3 B
port 2 e default input
rlabel m1 51 90 51 90 3 B
port 2 e default input
rlabel m1 59 22 59 22 3 #15
rlabel m1 48 31 48 31 3 GND
rlabel m1 48 41 48 41 3 Vdd
rlabel m1 48 45 48 45 3 Vdd
rlabel ndc 56 22 56 22 3 #15
rlabel m1 31 94 31 94 3 A
port 1 e default input
rlabel m1 31 98 31 98 3 A
port 1 e default input
rlabel m1 55 22 55 22 3 #15
rlabel m1 48 27 48 27 3 GND
rlabel m1 117 21 117 21 3 _YS
rlabel m1 40 28 40 28 3 #3
rlabel m1 40 20 40 20 3 #3
rlabel m1 40 24 40 24 3 #3
rlabel ndc 40 25 40 25 3 #3
rlabel m1 29 41 29 41 3 _YC
rlabel m1 23 86 23 86 3 B
port 2 e default input
rlabel m1 23 90 23 90 3 B
port 2 e default input
rlabel m1 102 7 102 7 3 _YC
rlabel m1 81 20 81 20 3 _YS
rlabel pdc 26 41 26 41 3 _YC
rlabel m1 36 47 36 47 3 #8
rlabel m1 33 13 33 13 3 GND
rlabel m1 33 17 33 17 3 GND
rlabel m1 33 31 33 31 3 GND
rlabel m1 25 41 25 41 3 _YC
rlabel pdc 33 47 33 47 3 #8
rlabel m1 18 27 18 27 3 _YC
rlabel m1 20 47 20 47 3 #8
rlabel m1 76 7 76 7 3 _YC
rlabel m1 25 6 25 6 3 _YC
rlabel m1 25 7 25 7 3 _YC
rlabel m1 25 10 25 10 3 _YC
rlabel pdc 17 47 17 47 3 #8
rlabel ndc 18 24 18 24 3 _YC
rlabel m1 16 47 16 47 3 #8
rlabel m1 16 78 16 78 3 C
port 3 e default input
rlabel m1 16 82 16 82 3 C
port 3 e default input
rlabel m1 18 6 18 6 3 _YC
rlabel m1 18 10 18 10 3 _YC
rlabel m1 10 20 10 20 3 #3
rlabel m1 10 24 10 24 3 #3
rlabel ndc 10 25 10 25 3 #3
rlabel m1 10 28 10 28 3 #3
rlabel m1 9 73 9 73 3 A
port 1 e default input
rlabel m2 121 21 121 21 3 _YS
rlabel m2c 118 21 118 21 3 _YS
rlabel m2 119 28 119 28 3 GND
rlabel m2 84 21 84 21 3 _YS
rlabel m2c 116 28 116 28 3 GND
rlabel m2c 81 21 81 21 3 _YS
rlabel m2 101 28 101 28 3 GND
rlabel m2 80 20 80 20 3 _YS
rlabel m2 80 21 80 21 3 _YS
rlabel m2 80 24 80 24 3 _YS
rlabel m2c 98 28 98 28 3 GND
rlabel m2 93 87 93 87 3 B
port 2 e default input
rlabel m2 67 28 67 28 3 GND
rlabel m2c 90 87 90 87 3 B
port 2 e default input
rlabel m2c 64 28 64 28 3 GND
rlabel m2 68 87 68 87 3 B
port 2 e default input
rlabel m2 51 28 51 28 3 GND
rlabel m2c 65 87 65 87 3 B
port 2 e default input
rlabel m2c 48 28 48 28 3 GND
rlabel m2 54 87 54 87 3 B
port 2 e default input
rlabel m2 106 7 106 7 3 _YC
rlabel m2 36 28 36 28 3 GND
rlabel m2 85 79 85 79 3 C
port 3 e default input
rlabel m2c 51 87 51 87 3 B
port 2 e default input
rlabel m2c 103 7 103 7 3 _YC
rlabel m2c 33 28 33 28 3 GND
rlabel m2 126 42 126 42 3 Vdd
rlabel m2c 82 79 82 79 3 C
port 3 e default input
rlabel m2 40 87 40 87 3 B
port 2 e default input
rlabel m2 101 95 101 95 3 A
port 1 e default input
rlabel m2 80 7 80 7 3 _YC
rlabel m2 32 27 32 27 3 GND
rlabel m2 32 28 32 28 3 GND
rlabel m2 32 31 32 31 3 GND
rlabel m2c 123 42 123 42 3 Vdd
rlabel m2 76 79 76 79 3 C
port 3 e default input
rlabel m2c 37 87 37 87 3 B
port 2 e default input
rlabel m2c 98 95 98 95 3 A
port 1 e default input
rlabel m2c 77 7 77 7 3 _YC
rlabel m2 101 42 101 42 3 Vdd
rlabel m2c 73 79 73 79 3 C
port 3 e default input
rlabel m2 26 87 26 87 3 B
port 2 e
rlabel m2 73 95 73 95 3 A
port 1 e default input
rlabel m2 29 7 29 7 3 _YC
rlabel m2c 98 42 98 42 3 Vdd
rlabel m2 62 79 62 79 3 C
port 3 e default input
rlabel m2c 23 87 23 87 3 B
port 2 e
rlabel m2c 70 95 70 95 3 A
port 1 e default input
rlabel m2c 26 7 26 7 3 _YC
rlabel m2 67 42 67 42 3 Vdd
rlabel m2c 59 79 59 79 3 C
port 3 e default input
rlabel m2 22 86 22 86 3 B
port 2 e
rlabel m2 22 87 22 87 3 B
port 2 e
rlabel m2 22 90 22 90 3 B
port 2 e
rlabel m2 48 95 48 95 3 A
port 1 e default input
rlabel m2 21 7 21 7 3 _YC
rlabel m2c 64 42 64 42 3 Vdd
rlabel m2 19 79 19 79 3 C
port 3 e
rlabel m2c 45 95 45 95 3 A
port 1 e default input
rlabel m2c 18 7 18 7 3 _YC
rlabel m2 43 21 43 21 3 #3
rlabel m2 51 42 51 42 3 Vdd
rlabel m2c 16 79 16 79 3 C
port 3 e
rlabel m2 34 95 34 95 3 A
port 1 e default input
rlabel m2 17 6 17 6 3 _YC
rlabel m2 17 7 17 7 3 _YC
rlabel m2 17 10 17 10 3 _YC
rlabel m2c 40 21 40 21 3 #3
rlabel m2c 48 42 48 42 3 Vdd
rlabel m2 15 78 15 78 3 C
port 3 e
rlabel m2 15 79 15 79 3 C
port 3 e
rlabel m2 15 82 15 82 3 C
port 3 e
rlabel m2c 31 95 31 95 3 A
port 1 e default input
rlabel m2 13 21 13 21 3 #3
rlabel m2 13 42 13 42 3 Vdd
rlabel m2 13 95 13 95 3 A
port 1 e
rlabel m2c 10 21 10 21 3 #3
rlabel m2c 10 42 10 42 3 Vdd
rlabel m2c 10 95 10 95 3 A
port 1 e
rlabel m2 9 20 9 20 3 #3
rlabel m2 9 21 9 21 3 #3
rlabel m2 9 24 9 24 3 #3
rlabel m2 9 41 9 41 3 Vdd
rlabel m2 9 42 9 42 3 Vdd
rlabel m2 9 45 9 45 3 Vdd
rlabel m2 9 94 9 94 3 A
port 1 e
rlabel m2 9 95 9 95 3 A
port 1 e
rlabel m2 9 98 9 98 3 A
port 1 e
<< properties >>
string LEFsite CoreSite
string LEFclass CORE
string FIXED_BBOX 0 0 136 100
string LEFsymmetry X Y
string LEFview TRUE
<< end >>
