magic
tech sky130l
timestamp 1731220421
<< m2 >>
rect 110 5692 116 5693
rect 1934 5692 1940 5693
rect 110 5688 111 5692
rect 115 5688 116 5692
rect 110 5687 116 5688
rect 130 5691 136 5692
rect 130 5687 131 5691
rect 135 5687 136 5691
rect 130 5686 136 5687
rect 266 5691 272 5692
rect 266 5687 267 5691
rect 271 5687 272 5691
rect 266 5686 272 5687
rect 402 5691 408 5692
rect 402 5687 403 5691
rect 407 5687 408 5691
rect 1934 5688 1935 5692
rect 1939 5688 1940 5692
rect 1934 5687 1940 5688
rect 402 5686 408 5687
rect 158 5676 164 5677
rect 110 5675 116 5676
rect 110 5671 111 5675
rect 115 5671 116 5675
rect 158 5672 159 5676
rect 163 5672 164 5676
rect 158 5671 164 5672
rect 294 5676 300 5677
rect 294 5672 295 5676
rect 299 5672 300 5676
rect 294 5671 300 5672
rect 430 5676 436 5677
rect 430 5672 431 5676
rect 435 5672 436 5676
rect 430 5671 436 5672
rect 1934 5675 1940 5676
rect 1934 5671 1935 5675
rect 1939 5671 1940 5675
rect 110 5670 116 5671
rect 1934 5670 1940 5671
rect 3838 5628 3844 5629
rect 5662 5628 5668 5629
rect 1974 5624 1980 5625
rect 3798 5624 3804 5625
rect 1974 5620 1975 5624
rect 1979 5620 1980 5624
rect 1974 5619 1980 5620
rect 1994 5623 2000 5624
rect 1994 5619 1995 5623
rect 1999 5619 2000 5623
rect 1994 5618 2000 5619
rect 2170 5623 2176 5624
rect 2170 5619 2171 5623
rect 2175 5619 2176 5623
rect 2170 5618 2176 5619
rect 2370 5623 2376 5624
rect 2370 5619 2371 5623
rect 2375 5619 2376 5623
rect 2370 5618 2376 5619
rect 2562 5623 2568 5624
rect 2562 5619 2563 5623
rect 2567 5619 2568 5623
rect 2562 5618 2568 5619
rect 2746 5623 2752 5624
rect 2746 5619 2747 5623
rect 2751 5619 2752 5623
rect 2746 5618 2752 5619
rect 2930 5623 2936 5624
rect 2930 5619 2931 5623
rect 2935 5619 2936 5623
rect 2930 5618 2936 5619
rect 3106 5623 3112 5624
rect 3106 5619 3107 5623
rect 3111 5619 3112 5623
rect 3106 5618 3112 5619
rect 3274 5623 3280 5624
rect 3274 5619 3275 5623
rect 3279 5619 3280 5623
rect 3274 5618 3280 5619
rect 3442 5623 3448 5624
rect 3442 5619 3443 5623
rect 3447 5619 3448 5623
rect 3442 5618 3448 5619
rect 3618 5623 3624 5624
rect 3618 5619 3619 5623
rect 3623 5619 3624 5623
rect 3798 5620 3799 5624
rect 3803 5620 3804 5624
rect 3838 5624 3839 5628
rect 3843 5624 3844 5628
rect 3838 5623 3844 5624
rect 4466 5627 4472 5628
rect 4466 5623 4467 5627
rect 4471 5623 4472 5627
rect 4466 5622 4472 5623
rect 4602 5627 4608 5628
rect 4602 5623 4603 5627
rect 4607 5623 4608 5627
rect 4602 5622 4608 5623
rect 4738 5627 4744 5628
rect 4738 5623 4739 5627
rect 4743 5623 4744 5627
rect 4738 5622 4744 5623
rect 4874 5627 4880 5628
rect 4874 5623 4875 5627
rect 4879 5623 4880 5627
rect 5662 5624 5663 5628
rect 5667 5624 5668 5628
rect 5662 5623 5668 5624
rect 4874 5622 4880 5623
rect 3798 5619 3804 5620
rect 3618 5618 3624 5619
rect 110 5617 116 5618
rect 1934 5617 1940 5618
rect 110 5613 111 5617
rect 115 5613 116 5617
rect 110 5612 116 5613
rect 342 5616 348 5617
rect 342 5612 343 5616
rect 347 5612 348 5616
rect 342 5611 348 5612
rect 534 5616 540 5617
rect 534 5612 535 5616
rect 539 5612 540 5616
rect 534 5611 540 5612
rect 734 5616 740 5617
rect 734 5612 735 5616
rect 739 5612 740 5616
rect 734 5611 740 5612
rect 942 5616 948 5617
rect 942 5612 943 5616
rect 947 5612 948 5616
rect 942 5611 948 5612
rect 1158 5616 1164 5617
rect 1158 5612 1159 5616
rect 1163 5612 1164 5616
rect 1158 5611 1164 5612
rect 1382 5616 1388 5617
rect 1382 5612 1383 5616
rect 1387 5612 1388 5616
rect 1382 5611 1388 5612
rect 1606 5616 1612 5617
rect 1606 5612 1607 5616
rect 1611 5612 1612 5616
rect 1606 5611 1612 5612
rect 1814 5616 1820 5617
rect 1814 5612 1815 5616
rect 1819 5612 1820 5616
rect 1934 5613 1935 5617
rect 1939 5613 1940 5617
rect 1934 5612 1940 5613
rect 4494 5612 4500 5613
rect 1814 5611 1820 5612
rect 3838 5611 3844 5612
rect 2022 5608 2028 5609
rect 1974 5607 1980 5608
rect 1974 5603 1975 5607
rect 1979 5603 1980 5607
rect 2022 5604 2023 5608
rect 2027 5604 2028 5608
rect 2022 5603 2028 5604
rect 2198 5608 2204 5609
rect 2198 5604 2199 5608
rect 2203 5604 2204 5608
rect 2198 5603 2204 5604
rect 2398 5608 2404 5609
rect 2398 5604 2399 5608
rect 2403 5604 2404 5608
rect 2398 5603 2404 5604
rect 2590 5608 2596 5609
rect 2590 5604 2591 5608
rect 2595 5604 2596 5608
rect 2590 5603 2596 5604
rect 2774 5608 2780 5609
rect 2774 5604 2775 5608
rect 2779 5604 2780 5608
rect 2774 5603 2780 5604
rect 2958 5608 2964 5609
rect 2958 5604 2959 5608
rect 2963 5604 2964 5608
rect 2958 5603 2964 5604
rect 3134 5608 3140 5609
rect 3134 5604 3135 5608
rect 3139 5604 3140 5608
rect 3134 5603 3140 5604
rect 3302 5608 3308 5609
rect 3302 5604 3303 5608
rect 3307 5604 3308 5608
rect 3302 5603 3308 5604
rect 3470 5608 3476 5609
rect 3470 5604 3471 5608
rect 3475 5604 3476 5608
rect 3470 5603 3476 5604
rect 3646 5608 3652 5609
rect 3646 5604 3647 5608
rect 3651 5604 3652 5608
rect 3646 5603 3652 5604
rect 3798 5607 3804 5608
rect 3798 5603 3799 5607
rect 3803 5603 3804 5607
rect 3838 5607 3839 5611
rect 3843 5607 3844 5611
rect 4494 5608 4495 5612
rect 4499 5608 4500 5612
rect 4494 5607 4500 5608
rect 4630 5612 4636 5613
rect 4630 5608 4631 5612
rect 4635 5608 4636 5612
rect 4630 5607 4636 5608
rect 4766 5612 4772 5613
rect 4766 5608 4767 5612
rect 4771 5608 4772 5612
rect 4766 5607 4772 5608
rect 4902 5612 4908 5613
rect 4902 5608 4903 5612
rect 4907 5608 4908 5612
rect 4902 5607 4908 5608
rect 5662 5611 5668 5612
rect 5662 5607 5663 5611
rect 5667 5607 5668 5611
rect 3838 5606 3844 5607
rect 5662 5606 5668 5607
rect 1974 5602 1980 5603
rect 3798 5602 3804 5603
rect 314 5601 320 5602
rect 110 5600 116 5601
rect 110 5596 111 5600
rect 115 5596 116 5600
rect 314 5597 315 5601
rect 319 5597 320 5601
rect 314 5596 320 5597
rect 506 5601 512 5602
rect 506 5597 507 5601
rect 511 5597 512 5601
rect 506 5596 512 5597
rect 706 5601 712 5602
rect 706 5597 707 5601
rect 711 5597 712 5601
rect 706 5596 712 5597
rect 914 5601 920 5602
rect 914 5597 915 5601
rect 919 5597 920 5601
rect 914 5596 920 5597
rect 1130 5601 1136 5602
rect 1130 5597 1131 5601
rect 1135 5597 1136 5601
rect 1130 5596 1136 5597
rect 1354 5601 1360 5602
rect 1354 5597 1355 5601
rect 1359 5597 1360 5601
rect 1354 5596 1360 5597
rect 1578 5601 1584 5602
rect 1578 5597 1579 5601
rect 1583 5597 1584 5601
rect 1578 5596 1584 5597
rect 1786 5601 1792 5602
rect 1786 5597 1787 5601
rect 1791 5597 1792 5601
rect 1786 5596 1792 5597
rect 1934 5600 1940 5601
rect 1934 5596 1935 5600
rect 1939 5596 1940 5600
rect 110 5595 116 5596
rect 1934 5595 1940 5596
rect 3838 5553 3844 5554
rect 5662 5553 5668 5554
rect 1974 5549 1980 5550
rect 3798 5549 3804 5550
rect 1974 5545 1975 5549
rect 1979 5545 1980 5549
rect 1974 5544 1980 5545
rect 2374 5548 2380 5549
rect 2374 5544 2375 5548
rect 2379 5544 2380 5548
rect 2374 5543 2380 5544
rect 2606 5548 2612 5549
rect 2606 5544 2607 5548
rect 2611 5544 2612 5548
rect 2606 5543 2612 5544
rect 2830 5548 2836 5549
rect 2830 5544 2831 5548
rect 2835 5544 2836 5548
rect 2830 5543 2836 5544
rect 3046 5548 3052 5549
rect 3046 5544 3047 5548
rect 3051 5544 3052 5548
rect 3046 5543 3052 5544
rect 3262 5548 3268 5549
rect 3262 5544 3263 5548
rect 3267 5544 3268 5548
rect 3262 5543 3268 5544
rect 3478 5548 3484 5549
rect 3478 5544 3479 5548
rect 3483 5544 3484 5548
rect 3478 5543 3484 5544
rect 3678 5548 3684 5549
rect 3678 5544 3679 5548
rect 3683 5544 3684 5548
rect 3798 5545 3799 5549
rect 3803 5545 3804 5549
rect 3838 5549 3839 5553
rect 3843 5549 3844 5553
rect 3838 5548 3844 5549
rect 4430 5552 4436 5553
rect 4430 5548 4431 5552
rect 4435 5548 4436 5552
rect 4430 5547 4436 5548
rect 4566 5552 4572 5553
rect 4566 5548 4567 5552
rect 4571 5548 4572 5552
rect 4566 5547 4572 5548
rect 4702 5552 4708 5553
rect 4702 5548 4703 5552
rect 4707 5548 4708 5552
rect 4702 5547 4708 5548
rect 4838 5552 4844 5553
rect 4838 5548 4839 5552
rect 4843 5548 4844 5552
rect 4838 5547 4844 5548
rect 4974 5552 4980 5553
rect 4974 5548 4975 5552
rect 4979 5548 4980 5552
rect 4974 5547 4980 5548
rect 5110 5552 5116 5553
rect 5110 5548 5111 5552
rect 5115 5548 5116 5552
rect 5662 5549 5663 5553
rect 5667 5549 5668 5553
rect 5662 5548 5668 5549
rect 5110 5547 5116 5548
rect 3798 5544 3804 5545
rect 3678 5543 3684 5544
rect 4402 5537 4408 5538
rect 3838 5536 3844 5537
rect 2346 5533 2352 5534
rect 1974 5532 1980 5533
rect 1974 5528 1975 5532
rect 1979 5528 1980 5532
rect 2346 5529 2347 5533
rect 2351 5529 2352 5533
rect 2346 5528 2352 5529
rect 2578 5533 2584 5534
rect 2578 5529 2579 5533
rect 2583 5529 2584 5533
rect 2578 5528 2584 5529
rect 2802 5533 2808 5534
rect 2802 5529 2803 5533
rect 2807 5529 2808 5533
rect 2802 5528 2808 5529
rect 3018 5533 3024 5534
rect 3018 5529 3019 5533
rect 3023 5529 3024 5533
rect 3018 5528 3024 5529
rect 3234 5533 3240 5534
rect 3234 5529 3235 5533
rect 3239 5529 3240 5533
rect 3234 5528 3240 5529
rect 3450 5533 3456 5534
rect 3450 5529 3451 5533
rect 3455 5529 3456 5533
rect 3450 5528 3456 5529
rect 3650 5533 3656 5534
rect 3650 5529 3651 5533
rect 3655 5529 3656 5533
rect 3650 5528 3656 5529
rect 3798 5532 3804 5533
rect 3798 5528 3799 5532
rect 3803 5528 3804 5532
rect 3838 5532 3839 5536
rect 3843 5532 3844 5536
rect 4402 5533 4403 5537
rect 4407 5533 4408 5537
rect 4402 5532 4408 5533
rect 4538 5537 4544 5538
rect 4538 5533 4539 5537
rect 4543 5533 4544 5537
rect 4538 5532 4544 5533
rect 4674 5537 4680 5538
rect 4674 5533 4675 5537
rect 4679 5533 4680 5537
rect 4674 5532 4680 5533
rect 4810 5537 4816 5538
rect 4810 5533 4811 5537
rect 4815 5533 4816 5537
rect 4810 5532 4816 5533
rect 4946 5537 4952 5538
rect 4946 5533 4947 5537
rect 4951 5533 4952 5537
rect 4946 5532 4952 5533
rect 5082 5537 5088 5538
rect 5082 5533 5083 5537
rect 5087 5533 5088 5537
rect 5082 5532 5088 5533
rect 5662 5536 5668 5537
rect 5662 5532 5663 5536
rect 5667 5532 5668 5536
rect 3838 5531 3844 5532
rect 5662 5531 5668 5532
rect 1974 5527 1980 5528
rect 3798 5527 3804 5528
rect 110 5468 116 5469
rect 1934 5468 1940 5469
rect 110 5464 111 5468
rect 115 5464 116 5468
rect 110 5463 116 5464
rect 874 5467 880 5468
rect 874 5463 875 5467
rect 879 5463 880 5467
rect 874 5462 880 5463
rect 1010 5467 1016 5468
rect 1010 5463 1011 5467
rect 1015 5463 1016 5467
rect 1010 5462 1016 5463
rect 1146 5467 1152 5468
rect 1146 5463 1147 5467
rect 1151 5463 1152 5467
rect 1146 5462 1152 5463
rect 1290 5467 1296 5468
rect 1290 5463 1291 5467
rect 1295 5463 1296 5467
rect 1290 5462 1296 5463
rect 1434 5467 1440 5468
rect 1434 5463 1435 5467
rect 1439 5463 1440 5467
rect 1434 5462 1440 5463
rect 1578 5467 1584 5468
rect 1578 5463 1579 5467
rect 1583 5463 1584 5467
rect 1578 5462 1584 5463
rect 1722 5467 1728 5468
rect 1722 5463 1723 5467
rect 1727 5463 1728 5467
rect 1934 5464 1935 5468
rect 1939 5464 1940 5468
rect 1934 5463 1940 5464
rect 1722 5462 1728 5463
rect 902 5452 908 5453
rect 110 5451 116 5452
rect 110 5447 111 5451
rect 115 5447 116 5451
rect 902 5448 903 5452
rect 907 5448 908 5452
rect 902 5447 908 5448
rect 1038 5452 1044 5453
rect 1038 5448 1039 5452
rect 1043 5448 1044 5452
rect 1038 5447 1044 5448
rect 1174 5452 1180 5453
rect 1174 5448 1175 5452
rect 1179 5448 1180 5452
rect 1174 5447 1180 5448
rect 1318 5452 1324 5453
rect 1318 5448 1319 5452
rect 1323 5448 1324 5452
rect 1318 5447 1324 5448
rect 1462 5452 1468 5453
rect 1462 5448 1463 5452
rect 1467 5448 1468 5452
rect 1462 5447 1468 5448
rect 1606 5452 1612 5453
rect 1606 5448 1607 5452
rect 1611 5448 1612 5452
rect 1606 5447 1612 5448
rect 1750 5452 1756 5453
rect 1750 5448 1751 5452
rect 1755 5448 1756 5452
rect 1750 5447 1756 5448
rect 1934 5451 1940 5452
rect 1934 5447 1935 5451
rect 1939 5447 1940 5451
rect 110 5446 116 5447
rect 1934 5446 1940 5447
rect 3838 5404 3844 5405
rect 5662 5404 5668 5405
rect 3838 5400 3839 5404
rect 3843 5400 3844 5404
rect 3838 5399 3844 5400
rect 4426 5403 4432 5404
rect 4426 5399 4427 5403
rect 4431 5399 4432 5403
rect 4426 5398 4432 5399
rect 4586 5403 4592 5404
rect 4586 5399 4587 5403
rect 4591 5399 4592 5403
rect 4586 5398 4592 5399
rect 4746 5403 4752 5404
rect 4746 5399 4747 5403
rect 4751 5399 4752 5403
rect 4746 5398 4752 5399
rect 4906 5403 4912 5404
rect 4906 5399 4907 5403
rect 4911 5399 4912 5403
rect 4906 5398 4912 5399
rect 5074 5403 5080 5404
rect 5074 5399 5075 5403
rect 5079 5399 5080 5403
rect 5662 5400 5663 5404
rect 5667 5400 5668 5404
rect 5662 5399 5668 5400
rect 5074 5398 5080 5399
rect 1974 5396 1980 5397
rect 3798 5396 3804 5397
rect 110 5393 116 5394
rect 1934 5393 1940 5394
rect 110 5389 111 5393
rect 115 5389 116 5393
rect 110 5388 116 5389
rect 718 5392 724 5393
rect 718 5388 719 5392
rect 723 5388 724 5392
rect 718 5387 724 5388
rect 854 5392 860 5393
rect 854 5388 855 5392
rect 859 5388 860 5392
rect 854 5387 860 5388
rect 990 5392 996 5393
rect 990 5388 991 5392
rect 995 5388 996 5392
rect 990 5387 996 5388
rect 1126 5392 1132 5393
rect 1126 5388 1127 5392
rect 1131 5388 1132 5392
rect 1126 5387 1132 5388
rect 1262 5392 1268 5393
rect 1262 5388 1263 5392
rect 1267 5388 1268 5392
rect 1262 5387 1268 5388
rect 1398 5392 1404 5393
rect 1398 5388 1399 5392
rect 1403 5388 1404 5392
rect 1398 5387 1404 5388
rect 1534 5392 1540 5393
rect 1534 5388 1535 5392
rect 1539 5388 1540 5392
rect 1534 5387 1540 5388
rect 1670 5392 1676 5393
rect 1670 5388 1671 5392
rect 1675 5388 1676 5392
rect 1670 5387 1676 5388
rect 1806 5392 1812 5393
rect 1806 5388 1807 5392
rect 1811 5388 1812 5392
rect 1934 5389 1935 5393
rect 1939 5389 1940 5393
rect 1974 5392 1975 5396
rect 1979 5392 1980 5396
rect 1974 5391 1980 5392
rect 2450 5395 2456 5396
rect 2450 5391 2451 5395
rect 2455 5391 2456 5395
rect 2450 5390 2456 5391
rect 2698 5395 2704 5396
rect 2698 5391 2699 5395
rect 2703 5391 2704 5395
rect 2698 5390 2704 5391
rect 2946 5395 2952 5396
rect 2946 5391 2947 5395
rect 2951 5391 2952 5395
rect 2946 5390 2952 5391
rect 3186 5395 3192 5396
rect 3186 5391 3187 5395
rect 3191 5391 3192 5395
rect 3186 5390 3192 5391
rect 3426 5395 3432 5396
rect 3426 5391 3427 5395
rect 3431 5391 3432 5395
rect 3426 5390 3432 5391
rect 3650 5395 3656 5396
rect 3650 5391 3651 5395
rect 3655 5391 3656 5395
rect 3798 5392 3799 5396
rect 3803 5392 3804 5396
rect 3798 5391 3804 5392
rect 3650 5390 3656 5391
rect 1934 5388 1940 5389
rect 4454 5388 4460 5389
rect 1806 5387 1812 5388
rect 3838 5387 3844 5388
rect 3838 5383 3839 5387
rect 3843 5383 3844 5387
rect 4454 5384 4455 5388
rect 4459 5384 4460 5388
rect 4454 5383 4460 5384
rect 4614 5388 4620 5389
rect 4614 5384 4615 5388
rect 4619 5384 4620 5388
rect 4614 5383 4620 5384
rect 4774 5388 4780 5389
rect 4774 5384 4775 5388
rect 4779 5384 4780 5388
rect 4774 5383 4780 5384
rect 4934 5388 4940 5389
rect 4934 5384 4935 5388
rect 4939 5384 4940 5388
rect 4934 5383 4940 5384
rect 5102 5388 5108 5389
rect 5102 5384 5103 5388
rect 5107 5384 5108 5388
rect 5102 5383 5108 5384
rect 5662 5387 5668 5388
rect 5662 5383 5663 5387
rect 5667 5383 5668 5387
rect 3838 5382 3844 5383
rect 5662 5382 5668 5383
rect 2478 5380 2484 5381
rect 1974 5379 1980 5380
rect 690 5377 696 5378
rect 110 5376 116 5377
rect 110 5372 111 5376
rect 115 5372 116 5376
rect 690 5373 691 5377
rect 695 5373 696 5377
rect 690 5372 696 5373
rect 826 5377 832 5378
rect 826 5373 827 5377
rect 831 5373 832 5377
rect 826 5372 832 5373
rect 962 5377 968 5378
rect 962 5373 963 5377
rect 967 5373 968 5377
rect 962 5372 968 5373
rect 1098 5377 1104 5378
rect 1098 5373 1099 5377
rect 1103 5373 1104 5377
rect 1098 5372 1104 5373
rect 1234 5377 1240 5378
rect 1234 5373 1235 5377
rect 1239 5373 1240 5377
rect 1234 5372 1240 5373
rect 1370 5377 1376 5378
rect 1370 5373 1371 5377
rect 1375 5373 1376 5377
rect 1370 5372 1376 5373
rect 1506 5377 1512 5378
rect 1506 5373 1507 5377
rect 1511 5373 1512 5377
rect 1506 5372 1512 5373
rect 1642 5377 1648 5378
rect 1642 5373 1643 5377
rect 1647 5373 1648 5377
rect 1642 5372 1648 5373
rect 1778 5377 1784 5378
rect 1778 5373 1779 5377
rect 1783 5373 1784 5377
rect 1778 5372 1784 5373
rect 1934 5376 1940 5377
rect 1934 5372 1935 5376
rect 1939 5372 1940 5376
rect 1974 5375 1975 5379
rect 1979 5375 1980 5379
rect 2478 5376 2479 5380
rect 2483 5376 2484 5380
rect 2478 5375 2484 5376
rect 2726 5380 2732 5381
rect 2726 5376 2727 5380
rect 2731 5376 2732 5380
rect 2726 5375 2732 5376
rect 2974 5380 2980 5381
rect 2974 5376 2975 5380
rect 2979 5376 2980 5380
rect 2974 5375 2980 5376
rect 3214 5380 3220 5381
rect 3214 5376 3215 5380
rect 3219 5376 3220 5380
rect 3214 5375 3220 5376
rect 3454 5380 3460 5381
rect 3454 5376 3455 5380
rect 3459 5376 3460 5380
rect 3454 5375 3460 5376
rect 3678 5380 3684 5381
rect 3678 5376 3679 5380
rect 3683 5376 3684 5380
rect 3678 5375 3684 5376
rect 3798 5379 3804 5380
rect 3798 5375 3799 5379
rect 3803 5375 3804 5379
rect 1974 5374 1980 5375
rect 3798 5374 3804 5375
rect 110 5371 116 5372
rect 1934 5371 1940 5372
rect 1974 5321 1980 5322
rect 3798 5321 3804 5322
rect 1974 5317 1975 5321
rect 1979 5317 1980 5321
rect 1974 5316 1980 5317
rect 2318 5320 2324 5321
rect 2318 5316 2319 5320
rect 2323 5316 2324 5320
rect 2318 5315 2324 5316
rect 2518 5320 2524 5321
rect 2518 5316 2519 5320
rect 2523 5316 2524 5320
rect 2518 5315 2524 5316
rect 2718 5320 2724 5321
rect 2718 5316 2719 5320
rect 2723 5316 2724 5320
rect 2718 5315 2724 5316
rect 2918 5320 2924 5321
rect 2918 5316 2919 5320
rect 2923 5316 2924 5320
rect 2918 5315 2924 5316
rect 3118 5320 3124 5321
rect 3118 5316 3119 5320
rect 3123 5316 3124 5320
rect 3118 5315 3124 5316
rect 3326 5320 3332 5321
rect 3326 5316 3327 5320
rect 3331 5316 3332 5320
rect 3326 5315 3332 5316
rect 3534 5320 3540 5321
rect 3534 5316 3535 5320
rect 3539 5316 3540 5320
rect 3798 5317 3799 5321
rect 3803 5317 3804 5321
rect 3798 5316 3804 5317
rect 3838 5321 3844 5322
rect 5662 5321 5668 5322
rect 3838 5317 3839 5321
rect 3843 5317 3844 5321
rect 3838 5316 3844 5317
rect 4430 5320 4436 5321
rect 4430 5316 4431 5320
rect 4435 5316 4436 5320
rect 3534 5315 3540 5316
rect 4430 5315 4436 5316
rect 4614 5320 4620 5321
rect 4614 5316 4615 5320
rect 4619 5316 4620 5320
rect 4614 5315 4620 5316
rect 4798 5320 4804 5321
rect 4798 5316 4799 5320
rect 4803 5316 4804 5320
rect 4798 5315 4804 5316
rect 4982 5320 4988 5321
rect 4982 5316 4983 5320
rect 4987 5316 4988 5320
rect 4982 5315 4988 5316
rect 5174 5320 5180 5321
rect 5174 5316 5175 5320
rect 5179 5316 5180 5320
rect 5662 5317 5663 5321
rect 5667 5317 5668 5321
rect 5662 5316 5668 5317
rect 5174 5315 5180 5316
rect 2290 5305 2296 5306
rect 1974 5304 1980 5305
rect 1974 5300 1975 5304
rect 1979 5300 1980 5304
rect 2290 5301 2291 5305
rect 2295 5301 2296 5305
rect 2290 5300 2296 5301
rect 2490 5305 2496 5306
rect 2490 5301 2491 5305
rect 2495 5301 2496 5305
rect 2490 5300 2496 5301
rect 2690 5305 2696 5306
rect 2690 5301 2691 5305
rect 2695 5301 2696 5305
rect 2690 5300 2696 5301
rect 2890 5305 2896 5306
rect 2890 5301 2891 5305
rect 2895 5301 2896 5305
rect 2890 5300 2896 5301
rect 3090 5305 3096 5306
rect 3090 5301 3091 5305
rect 3095 5301 3096 5305
rect 3090 5300 3096 5301
rect 3298 5305 3304 5306
rect 3298 5301 3299 5305
rect 3303 5301 3304 5305
rect 3298 5300 3304 5301
rect 3506 5305 3512 5306
rect 4402 5305 4408 5306
rect 3506 5301 3507 5305
rect 3511 5301 3512 5305
rect 3506 5300 3512 5301
rect 3798 5304 3804 5305
rect 3798 5300 3799 5304
rect 3803 5300 3804 5304
rect 1974 5299 1980 5300
rect 3798 5299 3804 5300
rect 3838 5304 3844 5305
rect 3838 5300 3839 5304
rect 3843 5300 3844 5304
rect 4402 5301 4403 5305
rect 4407 5301 4408 5305
rect 4402 5300 4408 5301
rect 4586 5305 4592 5306
rect 4586 5301 4587 5305
rect 4591 5301 4592 5305
rect 4586 5300 4592 5301
rect 4770 5305 4776 5306
rect 4770 5301 4771 5305
rect 4775 5301 4776 5305
rect 4770 5300 4776 5301
rect 4954 5305 4960 5306
rect 4954 5301 4955 5305
rect 4959 5301 4960 5305
rect 4954 5300 4960 5301
rect 5146 5305 5152 5306
rect 5146 5301 5147 5305
rect 5151 5301 5152 5305
rect 5146 5300 5152 5301
rect 5662 5304 5668 5305
rect 5662 5300 5663 5304
rect 5667 5300 5668 5304
rect 3838 5299 3844 5300
rect 5662 5299 5668 5300
rect 110 5244 116 5245
rect 1934 5244 1940 5245
rect 110 5240 111 5244
rect 115 5240 116 5244
rect 110 5239 116 5240
rect 722 5243 728 5244
rect 722 5239 723 5243
rect 727 5239 728 5243
rect 722 5238 728 5239
rect 874 5243 880 5244
rect 874 5239 875 5243
rect 879 5239 880 5243
rect 874 5238 880 5239
rect 1026 5243 1032 5244
rect 1026 5239 1027 5243
rect 1031 5239 1032 5243
rect 1026 5238 1032 5239
rect 1186 5243 1192 5244
rect 1186 5239 1187 5243
rect 1191 5239 1192 5243
rect 1186 5238 1192 5239
rect 1354 5243 1360 5244
rect 1354 5239 1355 5243
rect 1359 5239 1360 5243
rect 1354 5238 1360 5239
rect 1522 5243 1528 5244
rect 1522 5239 1523 5243
rect 1527 5239 1528 5243
rect 1934 5240 1935 5244
rect 1939 5240 1940 5244
rect 1934 5239 1940 5240
rect 1522 5238 1528 5239
rect 750 5228 756 5229
rect 110 5227 116 5228
rect 110 5223 111 5227
rect 115 5223 116 5227
rect 750 5224 751 5228
rect 755 5224 756 5228
rect 750 5223 756 5224
rect 902 5228 908 5229
rect 902 5224 903 5228
rect 907 5224 908 5228
rect 902 5223 908 5224
rect 1054 5228 1060 5229
rect 1054 5224 1055 5228
rect 1059 5224 1060 5228
rect 1054 5223 1060 5224
rect 1214 5228 1220 5229
rect 1214 5224 1215 5228
rect 1219 5224 1220 5228
rect 1214 5223 1220 5224
rect 1382 5228 1388 5229
rect 1382 5224 1383 5228
rect 1387 5224 1388 5228
rect 1382 5223 1388 5224
rect 1550 5228 1556 5229
rect 1550 5224 1551 5228
rect 1555 5224 1556 5228
rect 1550 5223 1556 5224
rect 1934 5227 1940 5228
rect 1934 5223 1935 5227
rect 1939 5223 1940 5227
rect 110 5222 116 5223
rect 1934 5222 1940 5223
rect 110 5169 116 5170
rect 1934 5169 1940 5170
rect 110 5165 111 5169
rect 115 5165 116 5169
rect 110 5164 116 5165
rect 446 5168 452 5169
rect 446 5164 447 5168
rect 451 5164 452 5168
rect 446 5163 452 5164
rect 622 5168 628 5169
rect 622 5164 623 5168
rect 627 5164 628 5168
rect 622 5163 628 5164
rect 806 5168 812 5169
rect 806 5164 807 5168
rect 811 5164 812 5168
rect 806 5163 812 5164
rect 998 5168 1004 5169
rect 998 5164 999 5168
rect 1003 5164 1004 5168
rect 998 5163 1004 5164
rect 1198 5168 1204 5169
rect 1198 5164 1199 5168
rect 1203 5164 1204 5168
rect 1198 5163 1204 5164
rect 1398 5168 1404 5169
rect 1398 5164 1399 5168
rect 1403 5164 1404 5168
rect 1398 5163 1404 5164
rect 1606 5168 1612 5169
rect 1606 5164 1607 5168
rect 1611 5164 1612 5168
rect 1606 5163 1612 5164
rect 1814 5168 1820 5169
rect 1814 5164 1815 5168
rect 1819 5164 1820 5168
rect 1934 5165 1935 5169
rect 1939 5165 1940 5169
rect 1934 5164 1940 5165
rect 1974 5168 1980 5169
rect 3798 5168 3804 5169
rect 1974 5164 1975 5168
rect 1979 5164 1980 5168
rect 1814 5163 1820 5164
rect 1974 5163 1980 5164
rect 2274 5167 2280 5168
rect 2274 5163 2275 5167
rect 2279 5163 2280 5167
rect 2274 5162 2280 5163
rect 2474 5167 2480 5168
rect 2474 5163 2475 5167
rect 2479 5163 2480 5167
rect 2474 5162 2480 5163
rect 2682 5167 2688 5168
rect 2682 5163 2683 5167
rect 2687 5163 2688 5167
rect 2682 5162 2688 5163
rect 2890 5167 2896 5168
rect 2890 5163 2891 5167
rect 2895 5163 2896 5167
rect 2890 5162 2896 5163
rect 3098 5167 3104 5168
rect 3098 5163 3099 5167
rect 3103 5163 3104 5167
rect 3098 5162 3104 5163
rect 3306 5167 3312 5168
rect 3306 5163 3307 5167
rect 3311 5163 3312 5167
rect 3798 5164 3799 5168
rect 3803 5164 3804 5168
rect 3798 5163 3804 5164
rect 3306 5162 3312 5163
rect 3838 5156 3844 5157
rect 5662 5156 5668 5157
rect 418 5153 424 5154
rect 110 5152 116 5153
rect 110 5148 111 5152
rect 115 5148 116 5152
rect 418 5149 419 5153
rect 423 5149 424 5153
rect 418 5148 424 5149
rect 594 5153 600 5154
rect 594 5149 595 5153
rect 599 5149 600 5153
rect 594 5148 600 5149
rect 778 5153 784 5154
rect 778 5149 779 5153
rect 783 5149 784 5153
rect 778 5148 784 5149
rect 970 5153 976 5154
rect 970 5149 971 5153
rect 975 5149 976 5153
rect 970 5148 976 5149
rect 1170 5153 1176 5154
rect 1170 5149 1171 5153
rect 1175 5149 1176 5153
rect 1170 5148 1176 5149
rect 1370 5153 1376 5154
rect 1370 5149 1371 5153
rect 1375 5149 1376 5153
rect 1370 5148 1376 5149
rect 1578 5153 1584 5154
rect 1578 5149 1579 5153
rect 1583 5149 1584 5153
rect 1578 5148 1584 5149
rect 1786 5153 1792 5154
rect 1786 5149 1787 5153
rect 1791 5149 1792 5153
rect 1786 5148 1792 5149
rect 1934 5152 1940 5153
rect 2302 5152 2308 5153
rect 1934 5148 1935 5152
rect 1939 5148 1940 5152
rect 110 5147 116 5148
rect 1934 5147 1940 5148
rect 1974 5151 1980 5152
rect 1974 5147 1975 5151
rect 1979 5147 1980 5151
rect 2302 5148 2303 5152
rect 2307 5148 2308 5152
rect 2302 5147 2308 5148
rect 2502 5152 2508 5153
rect 2502 5148 2503 5152
rect 2507 5148 2508 5152
rect 2502 5147 2508 5148
rect 2710 5152 2716 5153
rect 2710 5148 2711 5152
rect 2715 5148 2716 5152
rect 2710 5147 2716 5148
rect 2918 5152 2924 5153
rect 2918 5148 2919 5152
rect 2923 5148 2924 5152
rect 2918 5147 2924 5148
rect 3126 5152 3132 5153
rect 3126 5148 3127 5152
rect 3131 5148 3132 5152
rect 3126 5147 3132 5148
rect 3334 5152 3340 5153
rect 3838 5152 3839 5156
rect 3843 5152 3844 5156
rect 3334 5148 3335 5152
rect 3339 5148 3340 5152
rect 3334 5147 3340 5148
rect 3798 5151 3804 5152
rect 3838 5151 3844 5152
rect 4434 5155 4440 5156
rect 4434 5151 4435 5155
rect 4439 5151 4440 5155
rect 3798 5147 3799 5151
rect 3803 5147 3804 5151
rect 4434 5150 4440 5151
rect 4594 5155 4600 5156
rect 4594 5151 4595 5155
rect 4599 5151 4600 5155
rect 4594 5150 4600 5151
rect 4754 5155 4760 5156
rect 4754 5151 4755 5155
rect 4759 5151 4760 5155
rect 4754 5150 4760 5151
rect 4914 5155 4920 5156
rect 4914 5151 4915 5155
rect 4919 5151 4920 5155
rect 4914 5150 4920 5151
rect 5066 5155 5072 5156
rect 5066 5151 5067 5155
rect 5071 5151 5072 5155
rect 5066 5150 5072 5151
rect 5218 5155 5224 5156
rect 5218 5151 5219 5155
rect 5223 5151 5224 5155
rect 5218 5150 5224 5151
rect 5378 5155 5384 5156
rect 5378 5151 5379 5155
rect 5383 5151 5384 5155
rect 5378 5150 5384 5151
rect 5514 5155 5520 5156
rect 5514 5151 5515 5155
rect 5519 5151 5520 5155
rect 5662 5152 5663 5156
rect 5667 5152 5668 5156
rect 5662 5151 5668 5152
rect 5514 5150 5520 5151
rect 1974 5146 1980 5147
rect 3798 5146 3804 5147
rect 4462 5140 4468 5141
rect 3838 5139 3844 5140
rect 3838 5135 3839 5139
rect 3843 5135 3844 5139
rect 4462 5136 4463 5140
rect 4467 5136 4468 5140
rect 4462 5135 4468 5136
rect 4622 5140 4628 5141
rect 4622 5136 4623 5140
rect 4627 5136 4628 5140
rect 4622 5135 4628 5136
rect 4782 5140 4788 5141
rect 4782 5136 4783 5140
rect 4787 5136 4788 5140
rect 4782 5135 4788 5136
rect 4942 5140 4948 5141
rect 4942 5136 4943 5140
rect 4947 5136 4948 5140
rect 4942 5135 4948 5136
rect 5094 5140 5100 5141
rect 5094 5136 5095 5140
rect 5099 5136 5100 5140
rect 5094 5135 5100 5136
rect 5246 5140 5252 5141
rect 5246 5136 5247 5140
rect 5251 5136 5252 5140
rect 5246 5135 5252 5136
rect 5406 5140 5412 5141
rect 5406 5136 5407 5140
rect 5411 5136 5412 5140
rect 5406 5135 5412 5136
rect 5542 5140 5548 5141
rect 5542 5136 5543 5140
rect 5547 5136 5548 5140
rect 5542 5135 5548 5136
rect 5662 5139 5668 5140
rect 5662 5135 5663 5139
rect 5667 5135 5668 5139
rect 3838 5134 3844 5135
rect 5662 5134 5668 5135
rect 1974 5077 1980 5078
rect 3798 5077 3804 5078
rect 1974 5073 1975 5077
rect 1979 5073 1980 5077
rect 1974 5072 1980 5073
rect 2118 5076 2124 5077
rect 2118 5072 2119 5076
rect 2123 5072 2124 5076
rect 2118 5071 2124 5072
rect 2326 5076 2332 5077
rect 2326 5072 2327 5076
rect 2331 5072 2332 5076
rect 2326 5071 2332 5072
rect 2534 5076 2540 5077
rect 2534 5072 2535 5076
rect 2539 5072 2540 5076
rect 2534 5071 2540 5072
rect 2750 5076 2756 5077
rect 2750 5072 2751 5076
rect 2755 5072 2756 5076
rect 2750 5071 2756 5072
rect 2974 5076 2980 5077
rect 2974 5072 2975 5076
rect 2979 5072 2980 5076
rect 2974 5071 2980 5072
rect 3206 5076 3212 5077
rect 3206 5072 3207 5076
rect 3211 5072 3212 5076
rect 3798 5073 3799 5077
rect 3803 5073 3804 5077
rect 3798 5072 3804 5073
rect 3838 5073 3844 5074
rect 5662 5073 5668 5074
rect 3206 5071 3212 5072
rect 3838 5069 3839 5073
rect 3843 5069 3844 5073
rect 3838 5068 3844 5069
rect 3886 5072 3892 5073
rect 3886 5068 3887 5072
rect 3891 5068 3892 5072
rect 3886 5067 3892 5068
rect 4086 5072 4092 5073
rect 4086 5068 4087 5072
rect 4091 5068 4092 5072
rect 4086 5067 4092 5068
rect 4326 5072 4332 5073
rect 4326 5068 4327 5072
rect 4331 5068 4332 5072
rect 4326 5067 4332 5068
rect 4566 5072 4572 5073
rect 4566 5068 4567 5072
rect 4571 5068 4572 5072
rect 4566 5067 4572 5068
rect 4814 5072 4820 5073
rect 4814 5068 4815 5072
rect 4819 5068 4820 5072
rect 4814 5067 4820 5068
rect 5062 5072 5068 5073
rect 5062 5068 5063 5072
rect 5067 5068 5068 5072
rect 5062 5067 5068 5068
rect 5310 5072 5316 5073
rect 5310 5068 5311 5072
rect 5315 5068 5316 5072
rect 5310 5067 5316 5068
rect 5542 5072 5548 5073
rect 5542 5068 5543 5072
rect 5547 5068 5548 5072
rect 5662 5069 5663 5073
rect 5667 5069 5668 5073
rect 5662 5068 5668 5069
rect 5542 5067 5548 5068
rect 2090 5061 2096 5062
rect 1974 5060 1980 5061
rect 1974 5056 1975 5060
rect 1979 5056 1980 5060
rect 2090 5057 2091 5061
rect 2095 5057 2096 5061
rect 2090 5056 2096 5057
rect 2298 5061 2304 5062
rect 2298 5057 2299 5061
rect 2303 5057 2304 5061
rect 2298 5056 2304 5057
rect 2506 5061 2512 5062
rect 2506 5057 2507 5061
rect 2511 5057 2512 5061
rect 2506 5056 2512 5057
rect 2722 5061 2728 5062
rect 2722 5057 2723 5061
rect 2727 5057 2728 5061
rect 2722 5056 2728 5057
rect 2946 5061 2952 5062
rect 2946 5057 2947 5061
rect 2951 5057 2952 5061
rect 2946 5056 2952 5057
rect 3178 5061 3184 5062
rect 3178 5057 3179 5061
rect 3183 5057 3184 5061
rect 3178 5056 3184 5057
rect 3798 5060 3804 5061
rect 3798 5056 3799 5060
rect 3803 5056 3804 5060
rect 3858 5057 3864 5058
rect 1974 5055 1980 5056
rect 3798 5055 3804 5056
rect 3838 5056 3844 5057
rect 3838 5052 3839 5056
rect 3843 5052 3844 5056
rect 3858 5053 3859 5057
rect 3863 5053 3864 5057
rect 3858 5052 3864 5053
rect 4058 5057 4064 5058
rect 4058 5053 4059 5057
rect 4063 5053 4064 5057
rect 4058 5052 4064 5053
rect 4298 5057 4304 5058
rect 4298 5053 4299 5057
rect 4303 5053 4304 5057
rect 4298 5052 4304 5053
rect 4538 5057 4544 5058
rect 4538 5053 4539 5057
rect 4543 5053 4544 5057
rect 4538 5052 4544 5053
rect 4786 5057 4792 5058
rect 4786 5053 4787 5057
rect 4791 5053 4792 5057
rect 4786 5052 4792 5053
rect 5034 5057 5040 5058
rect 5034 5053 5035 5057
rect 5039 5053 5040 5057
rect 5034 5052 5040 5053
rect 5282 5057 5288 5058
rect 5282 5053 5283 5057
rect 5287 5053 5288 5057
rect 5282 5052 5288 5053
rect 5514 5057 5520 5058
rect 5514 5053 5515 5057
rect 5519 5053 5520 5057
rect 5514 5052 5520 5053
rect 5662 5056 5668 5057
rect 5662 5052 5663 5056
rect 5667 5052 5668 5056
rect 3838 5051 3844 5052
rect 5662 5051 5668 5052
rect 110 5012 116 5013
rect 1934 5012 1940 5013
rect 110 5008 111 5012
rect 115 5008 116 5012
rect 110 5007 116 5008
rect 154 5011 160 5012
rect 154 5007 155 5011
rect 159 5007 160 5011
rect 154 5006 160 5007
rect 378 5011 384 5012
rect 378 5007 379 5011
rect 383 5007 384 5011
rect 378 5006 384 5007
rect 626 5011 632 5012
rect 626 5007 627 5011
rect 631 5007 632 5011
rect 626 5006 632 5007
rect 898 5011 904 5012
rect 898 5007 899 5011
rect 903 5007 904 5011
rect 898 5006 904 5007
rect 1194 5011 1200 5012
rect 1194 5007 1195 5011
rect 1199 5007 1200 5011
rect 1194 5006 1200 5007
rect 1498 5011 1504 5012
rect 1498 5007 1499 5011
rect 1503 5007 1504 5011
rect 1498 5006 1504 5007
rect 1786 5011 1792 5012
rect 1786 5007 1787 5011
rect 1791 5007 1792 5011
rect 1934 5008 1935 5012
rect 1939 5008 1940 5012
rect 1934 5007 1940 5008
rect 1786 5006 1792 5007
rect 182 4996 188 4997
rect 110 4995 116 4996
rect 110 4991 111 4995
rect 115 4991 116 4995
rect 182 4992 183 4996
rect 187 4992 188 4996
rect 182 4991 188 4992
rect 406 4996 412 4997
rect 406 4992 407 4996
rect 411 4992 412 4996
rect 406 4991 412 4992
rect 654 4996 660 4997
rect 654 4992 655 4996
rect 659 4992 660 4996
rect 654 4991 660 4992
rect 926 4996 932 4997
rect 926 4992 927 4996
rect 931 4992 932 4996
rect 926 4991 932 4992
rect 1222 4996 1228 4997
rect 1222 4992 1223 4996
rect 1227 4992 1228 4996
rect 1222 4991 1228 4992
rect 1526 4996 1532 4997
rect 1526 4992 1527 4996
rect 1531 4992 1532 4996
rect 1526 4991 1532 4992
rect 1814 4996 1820 4997
rect 1814 4992 1815 4996
rect 1819 4992 1820 4996
rect 1814 4991 1820 4992
rect 1934 4995 1940 4996
rect 1934 4991 1935 4995
rect 1939 4991 1940 4995
rect 110 4990 116 4991
rect 1934 4990 1940 4991
rect 3838 4924 3844 4925
rect 5662 4924 5668 4925
rect 1974 4920 1980 4921
rect 3798 4920 3804 4921
rect 1974 4916 1975 4920
rect 1979 4916 1980 4920
rect 1974 4915 1980 4916
rect 1994 4919 2000 4920
rect 1994 4915 1995 4919
rect 1999 4915 2000 4919
rect 1994 4914 2000 4915
rect 2130 4919 2136 4920
rect 2130 4915 2131 4919
rect 2135 4915 2136 4919
rect 2130 4914 2136 4915
rect 2266 4919 2272 4920
rect 2266 4915 2267 4919
rect 2271 4915 2272 4919
rect 2266 4914 2272 4915
rect 2418 4919 2424 4920
rect 2418 4915 2419 4919
rect 2423 4915 2424 4919
rect 2418 4914 2424 4915
rect 2618 4919 2624 4920
rect 2618 4915 2619 4919
rect 2623 4915 2624 4919
rect 2618 4914 2624 4915
rect 2858 4919 2864 4920
rect 2858 4915 2859 4919
rect 2863 4915 2864 4919
rect 2858 4914 2864 4915
rect 3122 4919 3128 4920
rect 3122 4915 3123 4919
rect 3127 4915 3128 4919
rect 3122 4914 3128 4915
rect 3394 4919 3400 4920
rect 3394 4915 3395 4919
rect 3399 4915 3400 4919
rect 3394 4914 3400 4915
rect 3650 4919 3656 4920
rect 3650 4915 3651 4919
rect 3655 4915 3656 4919
rect 3798 4916 3799 4920
rect 3803 4916 3804 4920
rect 3838 4920 3839 4924
rect 3843 4920 3844 4924
rect 3838 4919 3844 4920
rect 3858 4923 3864 4924
rect 3858 4919 3859 4923
rect 3863 4919 3864 4923
rect 3858 4918 3864 4919
rect 3994 4923 4000 4924
rect 3994 4919 3995 4923
rect 3999 4919 4000 4923
rect 3994 4918 4000 4919
rect 4130 4923 4136 4924
rect 4130 4919 4131 4923
rect 4135 4919 4136 4923
rect 4130 4918 4136 4919
rect 4266 4923 4272 4924
rect 4266 4919 4267 4923
rect 4271 4919 4272 4923
rect 4266 4918 4272 4919
rect 4402 4923 4408 4924
rect 4402 4919 4403 4923
rect 4407 4919 4408 4923
rect 4402 4918 4408 4919
rect 4538 4923 4544 4924
rect 4538 4919 4539 4923
rect 4543 4919 4544 4923
rect 4538 4918 4544 4919
rect 4674 4923 4680 4924
rect 4674 4919 4675 4923
rect 4679 4919 4680 4923
rect 4674 4918 4680 4919
rect 4810 4923 4816 4924
rect 4810 4919 4811 4923
rect 4815 4919 4816 4923
rect 4810 4918 4816 4919
rect 4946 4923 4952 4924
rect 4946 4919 4947 4923
rect 4951 4919 4952 4923
rect 4946 4918 4952 4919
rect 5082 4923 5088 4924
rect 5082 4919 5083 4923
rect 5087 4919 5088 4923
rect 5082 4918 5088 4919
rect 5226 4923 5232 4924
rect 5226 4919 5227 4923
rect 5231 4919 5232 4923
rect 5226 4918 5232 4919
rect 5378 4923 5384 4924
rect 5378 4919 5379 4923
rect 5383 4919 5384 4923
rect 5378 4918 5384 4919
rect 5514 4923 5520 4924
rect 5514 4919 5515 4923
rect 5519 4919 5520 4923
rect 5662 4920 5663 4924
rect 5667 4920 5668 4924
rect 5662 4919 5668 4920
rect 5514 4918 5520 4919
rect 3798 4915 3804 4916
rect 3650 4914 3656 4915
rect 110 4909 116 4910
rect 1934 4909 1940 4910
rect 110 4905 111 4909
rect 115 4905 116 4909
rect 110 4904 116 4905
rect 158 4908 164 4909
rect 158 4904 159 4908
rect 163 4904 164 4908
rect 158 4903 164 4904
rect 294 4908 300 4909
rect 294 4904 295 4908
rect 299 4904 300 4908
rect 294 4903 300 4904
rect 430 4908 436 4909
rect 430 4904 431 4908
rect 435 4904 436 4908
rect 430 4903 436 4904
rect 566 4908 572 4909
rect 566 4904 567 4908
rect 571 4904 572 4908
rect 566 4903 572 4904
rect 702 4908 708 4909
rect 702 4904 703 4908
rect 707 4904 708 4908
rect 1934 4905 1935 4909
rect 1939 4905 1940 4909
rect 3886 4908 3892 4909
rect 3838 4907 3844 4908
rect 1934 4904 1940 4905
rect 2022 4904 2028 4905
rect 702 4903 708 4904
rect 1974 4903 1980 4904
rect 1974 4899 1975 4903
rect 1979 4899 1980 4903
rect 2022 4900 2023 4904
rect 2027 4900 2028 4904
rect 2022 4899 2028 4900
rect 2158 4904 2164 4905
rect 2158 4900 2159 4904
rect 2163 4900 2164 4904
rect 2158 4899 2164 4900
rect 2294 4904 2300 4905
rect 2294 4900 2295 4904
rect 2299 4900 2300 4904
rect 2294 4899 2300 4900
rect 2446 4904 2452 4905
rect 2446 4900 2447 4904
rect 2451 4900 2452 4904
rect 2446 4899 2452 4900
rect 2646 4904 2652 4905
rect 2646 4900 2647 4904
rect 2651 4900 2652 4904
rect 2646 4899 2652 4900
rect 2886 4904 2892 4905
rect 2886 4900 2887 4904
rect 2891 4900 2892 4904
rect 2886 4899 2892 4900
rect 3150 4904 3156 4905
rect 3150 4900 3151 4904
rect 3155 4900 3156 4904
rect 3150 4899 3156 4900
rect 3422 4904 3428 4905
rect 3422 4900 3423 4904
rect 3427 4900 3428 4904
rect 3422 4899 3428 4900
rect 3678 4904 3684 4905
rect 3678 4900 3679 4904
rect 3683 4900 3684 4904
rect 3678 4899 3684 4900
rect 3798 4903 3804 4904
rect 3798 4899 3799 4903
rect 3803 4899 3804 4903
rect 3838 4903 3839 4907
rect 3843 4903 3844 4907
rect 3886 4904 3887 4908
rect 3891 4904 3892 4908
rect 3886 4903 3892 4904
rect 4022 4908 4028 4909
rect 4022 4904 4023 4908
rect 4027 4904 4028 4908
rect 4022 4903 4028 4904
rect 4158 4908 4164 4909
rect 4158 4904 4159 4908
rect 4163 4904 4164 4908
rect 4158 4903 4164 4904
rect 4294 4908 4300 4909
rect 4294 4904 4295 4908
rect 4299 4904 4300 4908
rect 4294 4903 4300 4904
rect 4430 4908 4436 4909
rect 4430 4904 4431 4908
rect 4435 4904 4436 4908
rect 4430 4903 4436 4904
rect 4566 4908 4572 4909
rect 4566 4904 4567 4908
rect 4571 4904 4572 4908
rect 4566 4903 4572 4904
rect 4702 4908 4708 4909
rect 4702 4904 4703 4908
rect 4707 4904 4708 4908
rect 4702 4903 4708 4904
rect 4838 4908 4844 4909
rect 4838 4904 4839 4908
rect 4843 4904 4844 4908
rect 4838 4903 4844 4904
rect 4974 4908 4980 4909
rect 4974 4904 4975 4908
rect 4979 4904 4980 4908
rect 4974 4903 4980 4904
rect 5110 4908 5116 4909
rect 5110 4904 5111 4908
rect 5115 4904 5116 4908
rect 5110 4903 5116 4904
rect 5254 4908 5260 4909
rect 5254 4904 5255 4908
rect 5259 4904 5260 4908
rect 5254 4903 5260 4904
rect 5406 4908 5412 4909
rect 5406 4904 5407 4908
rect 5411 4904 5412 4908
rect 5406 4903 5412 4904
rect 5542 4908 5548 4909
rect 5542 4904 5543 4908
rect 5547 4904 5548 4908
rect 5542 4903 5548 4904
rect 5662 4907 5668 4908
rect 5662 4903 5663 4907
rect 5667 4903 5668 4907
rect 3838 4902 3844 4903
rect 5662 4902 5668 4903
rect 1974 4898 1980 4899
rect 3798 4898 3804 4899
rect 130 4893 136 4894
rect 110 4892 116 4893
rect 110 4888 111 4892
rect 115 4888 116 4892
rect 130 4889 131 4893
rect 135 4889 136 4893
rect 130 4888 136 4889
rect 266 4893 272 4894
rect 266 4889 267 4893
rect 271 4889 272 4893
rect 266 4888 272 4889
rect 402 4893 408 4894
rect 402 4889 403 4893
rect 407 4889 408 4893
rect 402 4888 408 4889
rect 538 4893 544 4894
rect 538 4889 539 4893
rect 543 4889 544 4893
rect 538 4888 544 4889
rect 674 4893 680 4894
rect 674 4889 675 4893
rect 679 4889 680 4893
rect 674 4888 680 4889
rect 1934 4892 1940 4893
rect 1934 4888 1935 4892
rect 1939 4888 1940 4892
rect 110 4887 116 4888
rect 1934 4887 1940 4888
rect 1974 4837 1980 4838
rect 3798 4837 3804 4838
rect 1974 4833 1975 4837
rect 1979 4833 1980 4837
rect 1974 4832 1980 4833
rect 2326 4836 2332 4837
rect 2326 4832 2327 4836
rect 2331 4832 2332 4836
rect 2326 4831 2332 4832
rect 2558 4836 2564 4837
rect 2558 4832 2559 4836
rect 2563 4832 2564 4836
rect 2558 4831 2564 4832
rect 2822 4836 2828 4837
rect 2822 4832 2823 4836
rect 2827 4832 2828 4836
rect 2822 4831 2828 4832
rect 3102 4836 3108 4837
rect 3102 4832 3103 4836
rect 3107 4832 3108 4836
rect 3102 4831 3108 4832
rect 3398 4836 3404 4837
rect 3398 4832 3399 4836
rect 3403 4832 3404 4836
rect 3398 4831 3404 4832
rect 3678 4836 3684 4837
rect 3678 4832 3679 4836
rect 3683 4832 3684 4836
rect 3798 4833 3799 4837
rect 3803 4833 3804 4837
rect 3798 4832 3804 4833
rect 3678 4831 3684 4832
rect 2298 4821 2304 4822
rect 1974 4820 1980 4821
rect 1974 4816 1975 4820
rect 1979 4816 1980 4820
rect 2298 4817 2299 4821
rect 2303 4817 2304 4821
rect 2298 4816 2304 4817
rect 2530 4821 2536 4822
rect 2530 4817 2531 4821
rect 2535 4817 2536 4821
rect 2530 4816 2536 4817
rect 2794 4821 2800 4822
rect 2794 4817 2795 4821
rect 2799 4817 2800 4821
rect 2794 4816 2800 4817
rect 3074 4821 3080 4822
rect 3074 4817 3075 4821
rect 3079 4817 3080 4821
rect 3074 4816 3080 4817
rect 3370 4821 3376 4822
rect 3370 4817 3371 4821
rect 3375 4817 3376 4821
rect 3370 4816 3376 4817
rect 3650 4821 3656 4822
rect 3650 4817 3651 4821
rect 3655 4817 3656 4821
rect 3650 4816 3656 4817
rect 3798 4820 3804 4821
rect 3798 4816 3799 4820
rect 3803 4816 3804 4820
rect 1974 4815 1980 4816
rect 3798 4815 3804 4816
rect 3838 4773 3844 4774
rect 5662 4773 5668 4774
rect 3838 4769 3839 4773
rect 3843 4769 3844 4773
rect 3838 4768 3844 4769
rect 3886 4772 3892 4773
rect 3886 4768 3887 4772
rect 3891 4768 3892 4772
rect 3886 4767 3892 4768
rect 4070 4772 4076 4773
rect 4070 4768 4071 4772
rect 4075 4768 4076 4772
rect 4070 4767 4076 4768
rect 4294 4772 4300 4773
rect 4294 4768 4295 4772
rect 4299 4768 4300 4772
rect 4294 4767 4300 4768
rect 4534 4772 4540 4773
rect 4534 4768 4535 4772
rect 4539 4768 4540 4772
rect 4534 4767 4540 4768
rect 4782 4772 4788 4773
rect 4782 4768 4783 4772
rect 4787 4768 4788 4772
rect 4782 4767 4788 4768
rect 5038 4772 5044 4773
rect 5038 4768 5039 4772
rect 5043 4768 5044 4772
rect 5038 4767 5044 4768
rect 5302 4772 5308 4773
rect 5302 4768 5303 4772
rect 5307 4768 5308 4772
rect 5302 4767 5308 4768
rect 5542 4772 5548 4773
rect 5542 4768 5543 4772
rect 5547 4768 5548 4772
rect 5662 4769 5663 4773
rect 5667 4769 5668 4773
rect 5662 4768 5668 4769
rect 5542 4767 5548 4768
rect 3858 4757 3864 4758
rect 3838 4756 3844 4757
rect 3838 4752 3839 4756
rect 3843 4752 3844 4756
rect 3858 4753 3859 4757
rect 3863 4753 3864 4757
rect 3858 4752 3864 4753
rect 4042 4757 4048 4758
rect 4042 4753 4043 4757
rect 4047 4753 4048 4757
rect 4042 4752 4048 4753
rect 4266 4757 4272 4758
rect 4266 4753 4267 4757
rect 4271 4753 4272 4757
rect 4266 4752 4272 4753
rect 4506 4757 4512 4758
rect 4506 4753 4507 4757
rect 4511 4753 4512 4757
rect 4506 4752 4512 4753
rect 4754 4757 4760 4758
rect 4754 4753 4755 4757
rect 4759 4753 4760 4757
rect 4754 4752 4760 4753
rect 5010 4757 5016 4758
rect 5010 4753 5011 4757
rect 5015 4753 5016 4757
rect 5010 4752 5016 4753
rect 5274 4757 5280 4758
rect 5274 4753 5275 4757
rect 5279 4753 5280 4757
rect 5274 4752 5280 4753
rect 5514 4757 5520 4758
rect 5514 4753 5515 4757
rect 5519 4753 5520 4757
rect 5514 4752 5520 4753
rect 5662 4756 5668 4757
rect 5662 4752 5663 4756
rect 5667 4752 5668 4756
rect 3838 4751 3844 4752
rect 5662 4751 5668 4752
rect 110 4748 116 4749
rect 1934 4748 1940 4749
rect 110 4744 111 4748
rect 115 4744 116 4748
rect 110 4743 116 4744
rect 130 4747 136 4748
rect 130 4743 131 4747
rect 135 4743 136 4747
rect 130 4742 136 4743
rect 266 4747 272 4748
rect 266 4743 267 4747
rect 271 4743 272 4747
rect 266 4742 272 4743
rect 402 4747 408 4748
rect 402 4743 403 4747
rect 407 4743 408 4747
rect 402 4742 408 4743
rect 538 4747 544 4748
rect 538 4743 539 4747
rect 543 4743 544 4747
rect 538 4742 544 4743
rect 674 4747 680 4748
rect 674 4743 675 4747
rect 679 4743 680 4747
rect 1934 4744 1935 4748
rect 1939 4744 1940 4748
rect 1934 4743 1940 4744
rect 674 4742 680 4743
rect 158 4732 164 4733
rect 110 4731 116 4732
rect 110 4727 111 4731
rect 115 4727 116 4731
rect 158 4728 159 4732
rect 163 4728 164 4732
rect 158 4727 164 4728
rect 294 4732 300 4733
rect 294 4728 295 4732
rect 299 4728 300 4732
rect 294 4727 300 4728
rect 430 4732 436 4733
rect 430 4728 431 4732
rect 435 4728 436 4732
rect 430 4727 436 4728
rect 566 4732 572 4733
rect 566 4728 567 4732
rect 571 4728 572 4732
rect 566 4727 572 4728
rect 702 4732 708 4733
rect 702 4728 703 4732
rect 707 4728 708 4732
rect 702 4727 708 4728
rect 1934 4731 1940 4732
rect 1934 4727 1935 4731
rect 1939 4727 1940 4731
rect 110 4726 116 4727
rect 1934 4726 1940 4727
rect 1974 4676 1980 4677
rect 3798 4676 3804 4677
rect 1974 4672 1975 4676
rect 1979 4672 1980 4676
rect 1974 4671 1980 4672
rect 2018 4675 2024 4676
rect 2018 4671 2019 4675
rect 2023 4671 2024 4675
rect 2018 4670 2024 4671
rect 2194 4675 2200 4676
rect 2194 4671 2195 4675
rect 2199 4671 2200 4675
rect 2194 4670 2200 4671
rect 2370 4675 2376 4676
rect 2370 4671 2371 4675
rect 2375 4671 2376 4675
rect 2370 4670 2376 4671
rect 2546 4675 2552 4676
rect 2546 4671 2547 4675
rect 2551 4671 2552 4675
rect 2546 4670 2552 4671
rect 2722 4675 2728 4676
rect 2722 4671 2723 4675
rect 2727 4671 2728 4675
rect 3798 4672 3799 4676
rect 3803 4672 3804 4676
rect 3798 4671 3804 4672
rect 2722 4670 2728 4671
rect 110 4669 116 4670
rect 1934 4669 1940 4670
rect 110 4665 111 4669
rect 115 4665 116 4669
rect 110 4664 116 4665
rect 158 4668 164 4669
rect 158 4664 159 4668
rect 163 4664 164 4668
rect 158 4663 164 4664
rect 294 4668 300 4669
rect 294 4664 295 4668
rect 299 4664 300 4668
rect 294 4663 300 4664
rect 430 4668 436 4669
rect 430 4664 431 4668
rect 435 4664 436 4668
rect 430 4663 436 4664
rect 566 4668 572 4669
rect 566 4664 567 4668
rect 571 4664 572 4668
rect 566 4663 572 4664
rect 702 4668 708 4669
rect 702 4664 703 4668
rect 707 4664 708 4668
rect 1934 4665 1935 4669
rect 1939 4665 1940 4669
rect 1934 4664 1940 4665
rect 702 4663 708 4664
rect 2046 4660 2052 4661
rect 1974 4659 1980 4660
rect 1974 4655 1975 4659
rect 1979 4655 1980 4659
rect 2046 4656 2047 4660
rect 2051 4656 2052 4660
rect 2046 4655 2052 4656
rect 2222 4660 2228 4661
rect 2222 4656 2223 4660
rect 2227 4656 2228 4660
rect 2222 4655 2228 4656
rect 2398 4660 2404 4661
rect 2398 4656 2399 4660
rect 2403 4656 2404 4660
rect 2398 4655 2404 4656
rect 2574 4660 2580 4661
rect 2574 4656 2575 4660
rect 2579 4656 2580 4660
rect 2574 4655 2580 4656
rect 2750 4660 2756 4661
rect 2750 4656 2751 4660
rect 2755 4656 2756 4660
rect 2750 4655 2756 4656
rect 3798 4659 3804 4660
rect 3798 4655 3799 4659
rect 3803 4655 3804 4659
rect 1974 4654 1980 4655
rect 3798 4654 3804 4655
rect 130 4653 136 4654
rect 110 4652 116 4653
rect 110 4648 111 4652
rect 115 4648 116 4652
rect 130 4649 131 4653
rect 135 4649 136 4653
rect 130 4648 136 4649
rect 266 4653 272 4654
rect 266 4649 267 4653
rect 271 4649 272 4653
rect 266 4648 272 4649
rect 402 4653 408 4654
rect 402 4649 403 4653
rect 407 4649 408 4653
rect 402 4648 408 4649
rect 538 4653 544 4654
rect 538 4649 539 4653
rect 543 4649 544 4653
rect 538 4648 544 4649
rect 674 4653 680 4654
rect 674 4649 675 4653
rect 679 4649 680 4653
rect 674 4648 680 4649
rect 1934 4652 1940 4653
rect 1934 4648 1935 4652
rect 1939 4648 1940 4652
rect 110 4647 116 4648
rect 1934 4647 1940 4648
rect 3838 4624 3844 4625
rect 5662 4624 5668 4625
rect 3838 4620 3839 4624
rect 3843 4620 3844 4624
rect 3838 4619 3844 4620
rect 3858 4623 3864 4624
rect 3858 4619 3859 4623
rect 3863 4619 3864 4623
rect 3858 4618 3864 4619
rect 3994 4623 4000 4624
rect 3994 4619 3995 4623
rect 3999 4619 4000 4623
rect 3994 4618 4000 4619
rect 4130 4623 4136 4624
rect 4130 4619 4131 4623
rect 4135 4619 4136 4623
rect 4130 4618 4136 4619
rect 4266 4623 4272 4624
rect 4266 4619 4267 4623
rect 4271 4619 4272 4623
rect 4266 4618 4272 4619
rect 4402 4623 4408 4624
rect 4402 4619 4403 4623
rect 4407 4619 4408 4623
rect 4402 4618 4408 4619
rect 4538 4623 4544 4624
rect 4538 4619 4539 4623
rect 4543 4619 4544 4623
rect 4538 4618 4544 4619
rect 4674 4623 4680 4624
rect 4674 4619 4675 4623
rect 4679 4619 4680 4623
rect 4674 4618 4680 4619
rect 4818 4623 4824 4624
rect 4818 4619 4819 4623
rect 4823 4619 4824 4623
rect 4818 4618 4824 4619
rect 4962 4623 4968 4624
rect 4962 4619 4963 4623
rect 4967 4619 4968 4623
rect 4962 4618 4968 4619
rect 5106 4623 5112 4624
rect 5106 4619 5107 4623
rect 5111 4619 5112 4623
rect 5106 4618 5112 4619
rect 5242 4623 5248 4624
rect 5242 4619 5243 4623
rect 5247 4619 5248 4623
rect 5242 4618 5248 4619
rect 5378 4623 5384 4624
rect 5378 4619 5379 4623
rect 5383 4619 5384 4623
rect 5378 4618 5384 4619
rect 5514 4623 5520 4624
rect 5514 4619 5515 4623
rect 5519 4619 5520 4623
rect 5662 4620 5663 4624
rect 5667 4620 5668 4624
rect 5662 4619 5668 4620
rect 5514 4618 5520 4619
rect 3886 4608 3892 4609
rect 3838 4607 3844 4608
rect 3838 4603 3839 4607
rect 3843 4603 3844 4607
rect 3886 4604 3887 4608
rect 3891 4604 3892 4608
rect 3886 4603 3892 4604
rect 4022 4608 4028 4609
rect 4022 4604 4023 4608
rect 4027 4604 4028 4608
rect 4022 4603 4028 4604
rect 4158 4608 4164 4609
rect 4158 4604 4159 4608
rect 4163 4604 4164 4608
rect 4158 4603 4164 4604
rect 4294 4608 4300 4609
rect 4294 4604 4295 4608
rect 4299 4604 4300 4608
rect 4294 4603 4300 4604
rect 4430 4608 4436 4609
rect 4430 4604 4431 4608
rect 4435 4604 4436 4608
rect 4430 4603 4436 4604
rect 4566 4608 4572 4609
rect 4566 4604 4567 4608
rect 4571 4604 4572 4608
rect 4566 4603 4572 4604
rect 4702 4608 4708 4609
rect 4702 4604 4703 4608
rect 4707 4604 4708 4608
rect 4702 4603 4708 4604
rect 4846 4608 4852 4609
rect 4846 4604 4847 4608
rect 4851 4604 4852 4608
rect 4846 4603 4852 4604
rect 4990 4608 4996 4609
rect 4990 4604 4991 4608
rect 4995 4604 4996 4608
rect 4990 4603 4996 4604
rect 5134 4608 5140 4609
rect 5134 4604 5135 4608
rect 5139 4604 5140 4608
rect 5134 4603 5140 4604
rect 5270 4608 5276 4609
rect 5270 4604 5271 4608
rect 5275 4604 5276 4608
rect 5270 4603 5276 4604
rect 5406 4608 5412 4609
rect 5406 4604 5407 4608
rect 5411 4604 5412 4608
rect 5406 4603 5412 4604
rect 5542 4608 5548 4609
rect 5542 4604 5543 4608
rect 5547 4604 5548 4608
rect 5542 4603 5548 4604
rect 5662 4607 5668 4608
rect 5662 4603 5663 4607
rect 5667 4603 5668 4607
rect 3838 4602 3844 4603
rect 5662 4602 5668 4603
rect 1974 4597 1980 4598
rect 3798 4597 3804 4598
rect 1974 4593 1975 4597
rect 1979 4593 1980 4597
rect 1974 4592 1980 4593
rect 2022 4596 2028 4597
rect 2022 4592 2023 4596
rect 2027 4592 2028 4596
rect 2022 4591 2028 4592
rect 2262 4596 2268 4597
rect 2262 4592 2263 4596
rect 2267 4592 2268 4596
rect 2262 4591 2268 4592
rect 2526 4596 2532 4597
rect 2526 4592 2527 4596
rect 2531 4592 2532 4596
rect 2526 4591 2532 4592
rect 2774 4596 2780 4597
rect 2774 4592 2775 4596
rect 2779 4592 2780 4596
rect 2774 4591 2780 4592
rect 3014 4596 3020 4597
rect 3014 4592 3015 4596
rect 3019 4592 3020 4596
rect 3014 4591 3020 4592
rect 3246 4596 3252 4597
rect 3246 4592 3247 4596
rect 3251 4592 3252 4596
rect 3246 4591 3252 4592
rect 3470 4596 3476 4597
rect 3470 4592 3471 4596
rect 3475 4592 3476 4596
rect 3470 4591 3476 4592
rect 3678 4596 3684 4597
rect 3678 4592 3679 4596
rect 3683 4592 3684 4596
rect 3798 4593 3799 4597
rect 3803 4593 3804 4597
rect 3798 4592 3804 4593
rect 3678 4591 3684 4592
rect 1994 4581 2000 4582
rect 1974 4580 1980 4581
rect 1974 4576 1975 4580
rect 1979 4576 1980 4580
rect 1994 4577 1995 4581
rect 1999 4577 2000 4581
rect 1994 4576 2000 4577
rect 2234 4581 2240 4582
rect 2234 4577 2235 4581
rect 2239 4577 2240 4581
rect 2234 4576 2240 4577
rect 2498 4581 2504 4582
rect 2498 4577 2499 4581
rect 2503 4577 2504 4581
rect 2498 4576 2504 4577
rect 2746 4581 2752 4582
rect 2746 4577 2747 4581
rect 2751 4577 2752 4581
rect 2746 4576 2752 4577
rect 2986 4581 2992 4582
rect 2986 4577 2987 4581
rect 2991 4577 2992 4581
rect 2986 4576 2992 4577
rect 3218 4581 3224 4582
rect 3218 4577 3219 4581
rect 3223 4577 3224 4581
rect 3218 4576 3224 4577
rect 3442 4581 3448 4582
rect 3442 4577 3443 4581
rect 3447 4577 3448 4581
rect 3442 4576 3448 4577
rect 3650 4581 3656 4582
rect 3650 4577 3651 4581
rect 3655 4577 3656 4581
rect 3650 4576 3656 4577
rect 3798 4580 3804 4581
rect 3798 4576 3799 4580
rect 3803 4576 3804 4580
rect 1974 4575 1980 4576
rect 3798 4575 3804 4576
rect 3838 4549 3844 4550
rect 5662 4549 5668 4550
rect 3838 4545 3839 4549
rect 3843 4545 3844 4549
rect 3838 4544 3844 4545
rect 4670 4548 4676 4549
rect 4670 4544 4671 4548
rect 4675 4544 4676 4548
rect 4670 4543 4676 4544
rect 4806 4548 4812 4549
rect 4806 4544 4807 4548
rect 4811 4544 4812 4548
rect 4806 4543 4812 4544
rect 4942 4548 4948 4549
rect 4942 4544 4943 4548
rect 4947 4544 4948 4548
rect 4942 4543 4948 4544
rect 5078 4548 5084 4549
rect 5078 4544 5079 4548
rect 5083 4544 5084 4548
rect 5662 4545 5663 4549
rect 5667 4545 5668 4549
rect 5662 4544 5668 4545
rect 5078 4543 5084 4544
rect 4642 4533 4648 4534
rect 3838 4532 3844 4533
rect 3838 4528 3839 4532
rect 3843 4528 3844 4532
rect 4642 4529 4643 4533
rect 4647 4529 4648 4533
rect 4642 4528 4648 4529
rect 4778 4533 4784 4534
rect 4778 4529 4779 4533
rect 4783 4529 4784 4533
rect 4778 4528 4784 4529
rect 4914 4533 4920 4534
rect 4914 4529 4915 4533
rect 4919 4529 4920 4533
rect 4914 4528 4920 4529
rect 5050 4533 5056 4534
rect 5050 4529 5051 4533
rect 5055 4529 5056 4533
rect 5050 4528 5056 4529
rect 5662 4532 5668 4533
rect 5662 4528 5663 4532
rect 5667 4528 5668 4532
rect 3838 4527 3844 4528
rect 5662 4527 5668 4528
rect 110 4508 116 4509
rect 1934 4508 1940 4509
rect 110 4504 111 4508
rect 115 4504 116 4508
rect 110 4503 116 4504
rect 250 4507 256 4508
rect 250 4503 251 4507
rect 255 4503 256 4507
rect 250 4502 256 4503
rect 442 4507 448 4508
rect 442 4503 443 4507
rect 447 4503 448 4507
rect 442 4502 448 4503
rect 650 4507 656 4508
rect 650 4503 651 4507
rect 655 4503 656 4507
rect 650 4502 656 4503
rect 874 4507 880 4508
rect 874 4503 875 4507
rect 879 4503 880 4507
rect 874 4502 880 4503
rect 1098 4507 1104 4508
rect 1098 4503 1099 4507
rect 1103 4503 1104 4507
rect 1098 4502 1104 4503
rect 1330 4507 1336 4508
rect 1330 4503 1331 4507
rect 1335 4503 1336 4507
rect 1330 4502 1336 4503
rect 1570 4507 1576 4508
rect 1570 4503 1571 4507
rect 1575 4503 1576 4507
rect 1570 4502 1576 4503
rect 1786 4507 1792 4508
rect 1786 4503 1787 4507
rect 1791 4503 1792 4507
rect 1934 4504 1935 4508
rect 1939 4504 1940 4508
rect 1934 4503 1940 4504
rect 1786 4502 1792 4503
rect 278 4492 284 4493
rect 110 4491 116 4492
rect 110 4487 111 4491
rect 115 4487 116 4491
rect 278 4488 279 4492
rect 283 4488 284 4492
rect 278 4487 284 4488
rect 470 4492 476 4493
rect 470 4488 471 4492
rect 475 4488 476 4492
rect 470 4487 476 4488
rect 678 4492 684 4493
rect 678 4488 679 4492
rect 683 4488 684 4492
rect 678 4487 684 4488
rect 902 4492 908 4493
rect 902 4488 903 4492
rect 907 4488 908 4492
rect 902 4487 908 4488
rect 1126 4492 1132 4493
rect 1126 4488 1127 4492
rect 1131 4488 1132 4492
rect 1126 4487 1132 4488
rect 1358 4492 1364 4493
rect 1358 4488 1359 4492
rect 1363 4488 1364 4492
rect 1358 4487 1364 4488
rect 1598 4492 1604 4493
rect 1598 4488 1599 4492
rect 1603 4488 1604 4492
rect 1598 4487 1604 4488
rect 1814 4492 1820 4493
rect 1814 4488 1815 4492
rect 1819 4488 1820 4492
rect 1814 4487 1820 4488
rect 1934 4491 1940 4492
rect 1934 4487 1935 4491
rect 1939 4487 1940 4491
rect 110 4486 116 4487
rect 1934 4486 1940 4487
rect 1974 4436 1980 4437
rect 3798 4436 3804 4437
rect 110 4433 116 4434
rect 1934 4433 1940 4434
rect 110 4429 111 4433
rect 115 4429 116 4433
rect 110 4428 116 4429
rect 510 4432 516 4433
rect 510 4428 511 4432
rect 515 4428 516 4432
rect 510 4427 516 4428
rect 686 4432 692 4433
rect 686 4428 687 4432
rect 691 4428 692 4432
rect 686 4427 692 4428
rect 870 4432 876 4433
rect 870 4428 871 4432
rect 875 4428 876 4432
rect 870 4427 876 4428
rect 1070 4432 1076 4433
rect 1070 4428 1071 4432
rect 1075 4428 1076 4432
rect 1070 4427 1076 4428
rect 1278 4432 1284 4433
rect 1278 4428 1279 4432
rect 1283 4428 1284 4432
rect 1278 4427 1284 4428
rect 1494 4432 1500 4433
rect 1494 4428 1495 4432
rect 1499 4428 1500 4432
rect 1494 4427 1500 4428
rect 1718 4432 1724 4433
rect 1718 4428 1719 4432
rect 1723 4428 1724 4432
rect 1934 4429 1935 4433
rect 1939 4429 1940 4433
rect 1974 4432 1975 4436
rect 1979 4432 1980 4436
rect 1974 4431 1980 4432
rect 2266 4435 2272 4436
rect 2266 4431 2267 4435
rect 2271 4431 2272 4435
rect 2266 4430 2272 4431
rect 2514 4435 2520 4436
rect 2514 4431 2515 4435
rect 2519 4431 2520 4435
rect 2514 4430 2520 4431
rect 2746 4435 2752 4436
rect 2746 4431 2747 4435
rect 2751 4431 2752 4435
rect 2746 4430 2752 4431
rect 2970 4435 2976 4436
rect 2970 4431 2971 4435
rect 2975 4431 2976 4435
rect 2970 4430 2976 4431
rect 3186 4435 3192 4436
rect 3186 4431 3187 4435
rect 3191 4431 3192 4435
rect 3186 4430 3192 4431
rect 3394 4435 3400 4436
rect 3394 4431 3395 4435
rect 3399 4431 3400 4435
rect 3394 4430 3400 4431
rect 3610 4435 3616 4436
rect 3610 4431 3611 4435
rect 3615 4431 3616 4435
rect 3798 4432 3799 4436
rect 3803 4432 3804 4436
rect 3798 4431 3804 4432
rect 3610 4430 3616 4431
rect 1934 4428 1940 4429
rect 1718 4427 1724 4428
rect 2294 4420 2300 4421
rect 1974 4419 1980 4420
rect 482 4417 488 4418
rect 110 4416 116 4417
rect 110 4412 111 4416
rect 115 4412 116 4416
rect 482 4413 483 4417
rect 487 4413 488 4417
rect 482 4412 488 4413
rect 658 4417 664 4418
rect 658 4413 659 4417
rect 663 4413 664 4417
rect 658 4412 664 4413
rect 842 4417 848 4418
rect 842 4413 843 4417
rect 847 4413 848 4417
rect 842 4412 848 4413
rect 1042 4417 1048 4418
rect 1042 4413 1043 4417
rect 1047 4413 1048 4417
rect 1042 4412 1048 4413
rect 1250 4417 1256 4418
rect 1250 4413 1251 4417
rect 1255 4413 1256 4417
rect 1250 4412 1256 4413
rect 1466 4417 1472 4418
rect 1466 4413 1467 4417
rect 1471 4413 1472 4417
rect 1466 4412 1472 4413
rect 1690 4417 1696 4418
rect 1690 4413 1691 4417
rect 1695 4413 1696 4417
rect 1690 4412 1696 4413
rect 1934 4416 1940 4417
rect 1934 4412 1935 4416
rect 1939 4412 1940 4416
rect 1974 4415 1975 4419
rect 1979 4415 1980 4419
rect 2294 4416 2295 4420
rect 2299 4416 2300 4420
rect 2294 4415 2300 4416
rect 2542 4420 2548 4421
rect 2542 4416 2543 4420
rect 2547 4416 2548 4420
rect 2542 4415 2548 4416
rect 2774 4420 2780 4421
rect 2774 4416 2775 4420
rect 2779 4416 2780 4420
rect 2774 4415 2780 4416
rect 2998 4420 3004 4421
rect 2998 4416 2999 4420
rect 3003 4416 3004 4420
rect 2998 4415 3004 4416
rect 3214 4420 3220 4421
rect 3214 4416 3215 4420
rect 3219 4416 3220 4420
rect 3214 4415 3220 4416
rect 3422 4420 3428 4421
rect 3422 4416 3423 4420
rect 3427 4416 3428 4420
rect 3422 4415 3428 4416
rect 3638 4420 3644 4421
rect 3638 4416 3639 4420
rect 3643 4416 3644 4420
rect 3638 4415 3644 4416
rect 3798 4419 3804 4420
rect 3798 4415 3799 4419
rect 3803 4415 3804 4419
rect 1974 4414 1980 4415
rect 3798 4414 3804 4415
rect 110 4411 116 4412
rect 1934 4411 1940 4412
rect 3838 4396 3844 4397
rect 5662 4396 5668 4397
rect 3838 4392 3839 4396
rect 3843 4392 3844 4396
rect 3838 4391 3844 4392
rect 4346 4395 4352 4396
rect 4346 4391 4347 4395
rect 4351 4391 4352 4395
rect 4346 4390 4352 4391
rect 4482 4395 4488 4396
rect 4482 4391 4483 4395
rect 4487 4391 4488 4395
rect 4482 4390 4488 4391
rect 4618 4395 4624 4396
rect 4618 4391 4619 4395
rect 4623 4391 4624 4395
rect 4618 4390 4624 4391
rect 4754 4395 4760 4396
rect 4754 4391 4755 4395
rect 4759 4391 4760 4395
rect 4754 4390 4760 4391
rect 4890 4395 4896 4396
rect 4890 4391 4891 4395
rect 4895 4391 4896 4395
rect 5662 4392 5663 4396
rect 5667 4392 5668 4396
rect 5662 4391 5668 4392
rect 4890 4390 4896 4391
rect 4374 4380 4380 4381
rect 3838 4379 3844 4380
rect 3838 4375 3839 4379
rect 3843 4375 3844 4379
rect 4374 4376 4375 4380
rect 4379 4376 4380 4380
rect 4374 4375 4380 4376
rect 4510 4380 4516 4381
rect 4510 4376 4511 4380
rect 4515 4376 4516 4380
rect 4510 4375 4516 4376
rect 4646 4380 4652 4381
rect 4646 4376 4647 4380
rect 4651 4376 4652 4380
rect 4646 4375 4652 4376
rect 4782 4380 4788 4381
rect 4782 4376 4783 4380
rect 4787 4376 4788 4380
rect 4782 4375 4788 4376
rect 4918 4380 4924 4381
rect 4918 4376 4919 4380
rect 4923 4376 4924 4380
rect 4918 4375 4924 4376
rect 5662 4379 5668 4380
rect 5662 4375 5663 4379
rect 5667 4375 5668 4379
rect 3838 4374 3844 4375
rect 5662 4374 5668 4375
rect 1974 4349 1980 4350
rect 3798 4349 3804 4350
rect 1974 4345 1975 4349
rect 1979 4345 1980 4349
rect 1974 4344 1980 4345
rect 2022 4348 2028 4349
rect 2022 4344 2023 4348
rect 2027 4344 2028 4348
rect 2022 4343 2028 4344
rect 2198 4348 2204 4349
rect 2198 4344 2199 4348
rect 2203 4344 2204 4348
rect 2198 4343 2204 4344
rect 2398 4348 2404 4349
rect 2398 4344 2399 4348
rect 2403 4344 2404 4348
rect 2398 4343 2404 4344
rect 2590 4348 2596 4349
rect 2590 4344 2591 4348
rect 2595 4344 2596 4348
rect 2590 4343 2596 4344
rect 2774 4348 2780 4349
rect 2774 4344 2775 4348
rect 2779 4344 2780 4348
rect 2774 4343 2780 4344
rect 2950 4348 2956 4349
rect 2950 4344 2951 4348
rect 2955 4344 2956 4348
rect 2950 4343 2956 4344
rect 3134 4348 3140 4349
rect 3134 4344 3135 4348
rect 3139 4344 3140 4348
rect 3134 4343 3140 4344
rect 3318 4348 3324 4349
rect 3318 4344 3319 4348
rect 3323 4344 3324 4348
rect 3798 4345 3799 4349
rect 3803 4345 3804 4349
rect 3798 4344 3804 4345
rect 3318 4343 3324 4344
rect 1994 4333 2000 4334
rect 1974 4332 1980 4333
rect 1974 4328 1975 4332
rect 1979 4328 1980 4332
rect 1994 4329 1995 4333
rect 1999 4329 2000 4333
rect 1994 4328 2000 4329
rect 2170 4333 2176 4334
rect 2170 4329 2171 4333
rect 2175 4329 2176 4333
rect 2170 4328 2176 4329
rect 2370 4333 2376 4334
rect 2370 4329 2371 4333
rect 2375 4329 2376 4333
rect 2370 4328 2376 4329
rect 2562 4333 2568 4334
rect 2562 4329 2563 4333
rect 2567 4329 2568 4333
rect 2562 4328 2568 4329
rect 2746 4333 2752 4334
rect 2746 4329 2747 4333
rect 2751 4329 2752 4333
rect 2746 4328 2752 4329
rect 2922 4333 2928 4334
rect 2922 4329 2923 4333
rect 2927 4329 2928 4333
rect 2922 4328 2928 4329
rect 3106 4333 3112 4334
rect 3106 4329 3107 4333
rect 3111 4329 3112 4333
rect 3106 4328 3112 4329
rect 3290 4333 3296 4334
rect 3290 4329 3291 4333
rect 3295 4329 3296 4333
rect 3290 4328 3296 4329
rect 3798 4332 3804 4333
rect 3798 4328 3799 4332
rect 3803 4328 3804 4332
rect 1974 4327 1980 4328
rect 3798 4327 3804 4328
rect 3838 4305 3844 4306
rect 5662 4305 5668 4306
rect 3838 4301 3839 4305
rect 3843 4301 3844 4305
rect 3838 4300 3844 4301
rect 4134 4304 4140 4305
rect 4134 4300 4135 4304
rect 4139 4300 4140 4304
rect 4134 4299 4140 4300
rect 4270 4304 4276 4305
rect 4270 4300 4271 4304
rect 4275 4300 4276 4304
rect 4270 4299 4276 4300
rect 4406 4304 4412 4305
rect 4406 4300 4407 4304
rect 4411 4300 4412 4304
rect 4406 4299 4412 4300
rect 4542 4304 4548 4305
rect 4542 4300 4543 4304
rect 4547 4300 4548 4304
rect 4542 4299 4548 4300
rect 4678 4304 4684 4305
rect 4678 4300 4679 4304
rect 4683 4300 4684 4304
rect 5662 4301 5663 4305
rect 5667 4301 5668 4305
rect 5662 4300 5668 4301
rect 4678 4299 4684 4300
rect 4106 4289 4112 4290
rect 3838 4288 3844 4289
rect 3838 4284 3839 4288
rect 3843 4284 3844 4288
rect 4106 4285 4107 4289
rect 4111 4285 4112 4289
rect 4106 4284 4112 4285
rect 4242 4289 4248 4290
rect 4242 4285 4243 4289
rect 4247 4285 4248 4289
rect 4242 4284 4248 4285
rect 4378 4289 4384 4290
rect 4378 4285 4379 4289
rect 4383 4285 4384 4289
rect 4378 4284 4384 4285
rect 4514 4289 4520 4290
rect 4514 4285 4515 4289
rect 4519 4285 4520 4289
rect 4514 4284 4520 4285
rect 4650 4289 4656 4290
rect 4650 4285 4651 4289
rect 4655 4285 4656 4289
rect 4650 4284 4656 4285
rect 5662 4288 5668 4289
rect 5662 4284 5663 4288
rect 5667 4284 5668 4288
rect 3838 4283 3844 4284
rect 5662 4283 5668 4284
rect 110 4280 116 4281
rect 1934 4280 1940 4281
rect 110 4276 111 4280
rect 115 4276 116 4280
rect 110 4275 116 4276
rect 714 4279 720 4280
rect 714 4275 715 4279
rect 719 4275 720 4279
rect 714 4274 720 4275
rect 850 4279 856 4280
rect 850 4275 851 4279
rect 855 4275 856 4279
rect 850 4274 856 4275
rect 986 4279 992 4280
rect 986 4275 987 4279
rect 991 4275 992 4279
rect 986 4274 992 4275
rect 1122 4279 1128 4280
rect 1122 4275 1123 4279
rect 1127 4275 1128 4279
rect 1122 4274 1128 4275
rect 1258 4279 1264 4280
rect 1258 4275 1259 4279
rect 1263 4275 1264 4279
rect 1258 4274 1264 4275
rect 1394 4279 1400 4280
rect 1394 4275 1395 4279
rect 1399 4275 1400 4279
rect 1394 4274 1400 4275
rect 1530 4279 1536 4280
rect 1530 4275 1531 4279
rect 1535 4275 1536 4279
rect 1530 4274 1536 4275
rect 1666 4279 1672 4280
rect 1666 4275 1667 4279
rect 1671 4275 1672 4279
rect 1934 4276 1935 4280
rect 1939 4276 1940 4280
rect 1934 4275 1940 4276
rect 1666 4274 1672 4275
rect 742 4264 748 4265
rect 110 4263 116 4264
rect 110 4259 111 4263
rect 115 4259 116 4263
rect 742 4260 743 4264
rect 747 4260 748 4264
rect 742 4259 748 4260
rect 878 4264 884 4265
rect 878 4260 879 4264
rect 883 4260 884 4264
rect 878 4259 884 4260
rect 1014 4264 1020 4265
rect 1014 4260 1015 4264
rect 1019 4260 1020 4264
rect 1014 4259 1020 4260
rect 1150 4264 1156 4265
rect 1150 4260 1151 4264
rect 1155 4260 1156 4264
rect 1150 4259 1156 4260
rect 1286 4264 1292 4265
rect 1286 4260 1287 4264
rect 1291 4260 1292 4264
rect 1286 4259 1292 4260
rect 1422 4264 1428 4265
rect 1422 4260 1423 4264
rect 1427 4260 1428 4264
rect 1422 4259 1428 4260
rect 1558 4264 1564 4265
rect 1558 4260 1559 4264
rect 1563 4260 1564 4264
rect 1558 4259 1564 4260
rect 1694 4264 1700 4265
rect 1694 4260 1695 4264
rect 1699 4260 1700 4264
rect 1694 4259 1700 4260
rect 1934 4263 1940 4264
rect 1934 4259 1935 4263
rect 1939 4259 1940 4263
rect 110 4258 116 4259
rect 1934 4258 1940 4259
rect 110 4197 116 4198
rect 1934 4197 1940 4198
rect 110 4193 111 4197
rect 115 4193 116 4197
rect 110 4192 116 4193
rect 726 4196 732 4197
rect 726 4192 727 4196
rect 731 4192 732 4196
rect 726 4191 732 4192
rect 862 4196 868 4197
rect 862 4192 863 4196
rect 867 4192 868 4196
rect 862 4191 868 4192
rect 998 4196 1004 4197
rect 998 4192 999 4196
rect 1003 4192 1004 4196
rect 998 4191 1004 4192
rect 1134 4196 1140 4197
rect 1134 4192 1135 4196
rect 1139 4192 1140 4196
rect 1134 4191 1140 4192
rect 1270 4196 1276 4197
rect 1270 4192 1271 4196
rect 1275 4192 1276 4196
rect 1270 4191 1276 4192
rect 1406 4196 1412 4197
rect 1406 4192 1407 4196
rect 1411 4192 1412 4196
rect 1406 4191 1412 4192
rect 1542 4196 1548 4197
rect 1542 4192 1543 4196
rect 1547 4192 1548 4196
rect 1542 4191 1548 4192
rect 1678 4196 1684 4197
rect 1678 4192 1679 4196
rect 1683 4192 1684 4196
rect 1678 4191 1684 4192
rect 1814 4196 1820 4197
rect 1814 4192 1815 4196
rect 1819 4192 1820 4196
rect 1934 4193 1935 4197
rect 1939 4193 1940 4197
rect 1934 4192 1940 4193
rect 1974 4196 1980 4197
rect 3798 4196 3804 4197
rect 1974 4192 1975 4196
rect 1979 4192 1980 4196
rect 1814 4191 1820 4192
rect 1974 4191 1980 4192
rect 1994 4195 2000 4196
rect 1994 4191 1995 4195
rect 1999 4191 2000 4195
rect 1994 4190 2000 4191
rect 2242 4195 2248 4196
rect 2242 4191 2243 4195
rect 2247 4191 2248 4195
rect 2242 4190 2248 4191
rect 2506 4195 2512 4196
rect 2506 4191 2507 4195
rect 2511 4191 2512 4195
rect 2506 4190 2512 4191
rect 2762 4195 2768 4196
rect 2762 4191 2763 4195
rect 2767 4191 2768 4195
rect 2762 4190 2768 4191
rect 3018 4195 3024 4196
rect 3018 4191 3019 4195
rect 3023 4191 3024 4195
rect 3018 4190 3024 4191
rect 3282 4195 3288 4196
rect 3282 4191 3283 4195
rect 3287 4191 3288 4195
rect 3798 4192 3799 4196
rect 3803 4192 3804 4196
rect 3798 4191 3804 4192
rect 3282 4190 3288 4191
rect 698 4181 704 4182
rect 110 4180 116 4181
rect 110 4176 111 4180
rect 115 4176 116 4180
rect 698 4177 699 4181
rect 703 4177 704 4181
rect 698 4176 704 4177
rect 834 4181 840 4182
rect 834 4177 835 4181
rect 839 4177 840 4181
rect 834 4176 840 4177
rect 970 4181 976 4182
rect 970 4177 971 4181
rect 975 4177 976 4181
rect 970 4176 976 4177
rect 1106 4181 1112 4182
rect 1106 4177 1107 4181
rect 1111 4177 1112 4181
rect 1106 4176 1112 4177
rect 1242 4181 1248 4182
rect 1242 4177 1243 4181
rect 1247 4177 1248 4181
rect 1242 4176 1248 4177
rect 1378 4181 1384 4182
rect 1378 4177 1379 4181
rect 1383 4177 1384 4181
rect 1378 4176 1384 4177
rect 1514 4181 1520 4182
rect 1514 4177 1515 4181
rect 1519 4177 1520 4181
rect 1514 4176 1520 4177
rect 1650 4181 1656 4182
rect 1650 4177 1651 4181
rect 1655 4177 1656 4181
rect 1650 4176 1656 4177
rect 1786 4181 1792 4182
rect 1786 4177 1787 4181
rect 1791 4177 1792 4181
rect 1786 4176 1792 4177
rect 1934 4180 1940 4181
rect 2022 4180 2028 4181
rect 1934 4176 1935 4180
rect 1939 4176 1940 4180
rect 110 4175 116 4176
rect 1934 4175 1940 4176
rect 1974 4179 1980 4180
rect 1974 4175 1975 4179
rect 1979 4175 1980 4179
rect 2022 4176 2023 4180
rect 2027 4176 2028 4180
rect 2022 4175 2028 4176
rect 2270 4180 2276 4181
rect 2270 4176 2271 4180
rect 2275 4176 2276 4180
rect 2270 4175 2276 4176
rect 2534 4180 2540 4181
rect 2534 4176 2535 4180
rect 2539 4176 2540 4180
rect 2534 4175 2540 4176
rect 2790 4180 2796 4181
rect 2790 4176 2791 4180
rect 2795 4176 2796 4180
rect 2790 4175 2796 4176
rect 3046 4180 3052 4181
rect 3046 4176 3047 4180
rect 3051 4176 3052 4180
rect 3046 4175 3052 4176
rect 3310 4180 3316 4181
rect 3310 4176 3311 4180
rect 3315 4176 3316 4180
rect 3310 4175 3316 4176
rect 3798 4179 3804 4180
rect 3798 4175 3799 4179
rect 3803 4175 3804 4179
rect 1974 4174 1980 4175
rect 3798 4174 3804 4175
rect 3838 4144 3844 4145
rect 5662 4144 5668 4145
rect 3838 4140 3839 4144
rect 3843 4140 3844 4144
rect 3838 4139 3844 4140
rect 3970 4143 3976 4144
rect 3970 4139 3971 4143
rect 3975 4139 3976 4143
rect 3970 4138 3976 4139
rect 4106 4143 4112 4144
rect 4106 4139 4107 4143
rect 4111 4139 4112 4143
rect 4106 4138 4112 4139
rect 4242 4143 4248 4144
rect 4242 4139 4243 4143
rect 4247 4139 4248 4143
rect 4242 4138 4248 4139
rect 4378 4143 4384 4144
rect 4378 4139 4379 4143
rect 4383 4139 4384 4143
rect 4378 4138 4384 4139
rect 4514 4143 4520 4144
rect 4514 4139 4515 4143
rect 4519 4139 4520 4143
rect 5662 4140 5663 4144
rect 5667 4140 5668 4144
rect 5662 4139 5668 4140
rect 4514 4138 4520 4139
rect 3998 4128 4004 4129
rect 3838 4127 3844 4128
rect 3838 4123 3839 4127
rect 3843 4123 3844 4127
rect 3998 4124 3999 4128
rect 4003 4124 4004 4128
rect 3998 4123 4004 4124
rect 4134 4128 4140 4129
rect 4134 4124 4135 4128
rect 4139 4124 4140 4128
rect 4134 4123 4140 4124
rect 4270 4128 4276 4129
rect 4270 4124 4271 4128
rect 4275 4124 4276 4128
rect 4270 4123 4276 4124
rect 4406 4128 4412 4129
rect 4406 4124 4407 4128
rect 4411 4124 4412 4128
rect 4406 4123 4412 4124
rect 4542 4128 4548 4129
rect 4542 4124 4543 4128
rect 4547 4124 4548 4128
rect 4542 4123 4548 4124
rect 5662 4127 5668 4128
rect 5662 4123 5663 4127
rect 5667 4123 5668 4127
rect 3838 4122 3844 4123
rect 5662 4122 5668 4123
rect 1974 4109 1980 4110
rect 3798 4109 3804 4110
rect 1974 4105 1975 4109
rect 1979 4105 1980 4109
rect 1974 4104 1980 4105
rect 3134 4108 3140 4109
rect 3134 4104 3135 4108
rect 3139 4104 3140 4108
rect 3134 4103 3140 4104
rect 3270 4108 3276 4109
rect 3270 4104 3271 4108
rect 3275 4104 3276 4108
rect 3270 4103 3276 4104
rect 3406 4108 3412 4109
rect 3406 4104 3407 4108
rect 3411 4104 3412 4108
rect 3406 4103 3412 4104
rect 3542 4108 3548 4109
rect 3542 4104 3543 4108
rect 3547 4104 3548 4108
rect 3542 4103 3548 4104
rect 3678 4108 3684 4109
rect 3678 4104 3679 4108
rect 3683 4104 3684 4108
rect 3798 4105 3799 4109
rect 3803 4105 3804 4109
rect 3798 4104 3804 4105
rect 3678 4103 3684 4104
rect 3106 4093 3112 4094
rect 1974 4092 1980 4093
rect 1974 4088 1975 4092
rect 1979 4088 1980 4092
rect 3106 4089 3107 4093
rect 3111 4089 3112 4093
rect 3106 4088 3112 4089
rect 3242 4093 3248 4094
rect 3242 4089 3243 4093
rect 3247 4089 3248 4093
rect 3242 4088 3248 4089
rect 3378 4093 3384 4094
rect 3378 4089 3379 4093
rect 3383 4089 3384 4093
rect 3378 4088 3384 4089
rect 3514 4093 3520 4094
rect 3514 4089 3515 4093
rect 3519 4089 3520 4093
rect 3514 4088 3520 4089
rect 3650 4093 3656 4094
rect 3650 4089 3651 4093
rect 3655 4089 3656 4093
rect 3650 4088 3656 4089
rect 3798 4092 3804 4093
rect 3798 4088 3799 4092
rect 3803 4088 3804 4092
rect 1974 4087 1980 4088
rect 3798 4087 3804 4088
rect 110 4048 116 4049
rect 1934 4048 1940 4049
rect 110 4044 111 4048
rect 115 4044 116 4048
rect 110 4043 116 4044
rect 562 4047 568 4048
rect 562 4043 563 4047
rect 567 4043 568 4047
rect 562 4042 568 4043
rect 698 4047 704 4048
rect 698 4043 699 4047
rect 703 4043 704 4047
rect 698 4042 704 4043
rect 834 4047 840 4048
rect 834 4043 835 4047
rect 839 4043 840 4047
rect 834 4042 840 4043
rect 970 4047 976 4048
rect 970 4043 971 4047
rect 975 4043 976 4047
rect 970 4042 976 4043
rect 1106 4047 1112 4048
rect 1106 4043 1107 4047
rect 1111 4043 1112 4047
rect 1106 4042 1112 4043
rect 1242 4047 1248 4048
rect 1242 4043 1243 4047
rect 1247 4043 1248 4047
rect 1242 4042 1248 4043
rect 1378 4047 1384 4048
rect 1378 4043 1379 4047
rect 1383 4043 1384 4047
rect 1378 4042 1384 4043
rect 1514 4047 1520 4048
rect 1514 4043 1515 4047
rect 1519 4043 1520 4047
rect 1514 4042 1520 4043
rect 1650 4047 1656 4048
rect 1650 4043 1651 4047
rect 1655 4043 1656 4047
rect 1650 4042 1656 4043
rect 1786 4047 1792 4048
rect 1786 4043 1787 4047
rect 1791 4043 1792 4047
rect 1934 4044 1935 4048
rect 1939 4044 1940 4048
rect 1934 4043 1940 4044
rect 3838 4045 3844 4046
rect 5662 4045 5668 4046
rect 1786 4042 1792 4043
rect 3838 4041 3839 4045
rect 3843 4041 3844 4045
rect 3838 4040 3844 4041
rect 3886 4044 3892 4045
rect 3886 4040 3887 4044
rect 3891 4040 3892 4044
rect 3886 4039 3892 4040
rect 4022 4044 4028 4045
rect 4022 4040 4023 4044
rect 4027 4040 4028 4044
rect 4022 4039 4028 4040
rect 4158 4044 4164 4045
rect 4158 4040 4159 4044
rect 4163 4040 4164 4044
rect 4158 4039 4164 4040
rect 4294 4044 4300 4045
rect 4294 4040 4295 4044
rect 4299 4040 4300 4044
rect 4294 4039 4300 4040
rect 4430 4044 4436 4045
rect 4430 4040 4431 4044
rect 4435 4040 4436 4044
rect 4430 4039 4436 4040
rect 4566 4044 4572 4045
rect 4566 4040 4567 4044
rect 4571 4040 4572 4044
rect 4566 4039 4572 4040
rect 4702 4044 4708 4045
rect 4702 4040 4703 4044
rect 4707 4040 4708 4044
rect 4702 4039 4708 4040
rect 4838 4044 4844 4045
rect 4838 4040 4839 4044
rect 4843 4040 4844 4044
rect 5662 4041 5663 4045
rect 5667 4041 5668 4045
rect 5662 4040 5668 4041
rect 4838 4039 4844 4040
rect 590 4032 596 4033
rect 110 4031 116 4032
rect 110 4027 111 4031
rect 115 4027 116 4031
rect 590 4028 591 4032
rect 595 4028 596 4032
rect 590 4027 596 4028
rect 726 4032 732 4033
rect 726 4028 727 4032
rect 731 4028 732 4032
rect 726 4027 732 4028
rect 862 4032 868 4033
rect 862 4028 863 4032
rect 867 4028 868 4032
rect 862 4027 868 4028
rect 998 4032 1004 4033
rect 998 4028 999 4032
rect 1003 4028 1004 4032
rect 998 4027 1004 4028
rect 1134 4032 1140 4033
rect 1134 4028 1135 4032
rect 1139 4028 1140 4032
rect 1134 4027 1140 4028
rect 1270 4032 1276 4033
rect 1270 4028 1271 4032
rect 1275 4028 1276 4032
rect 1270 4027 1276 4028
rect 1406 4032 1412 4033
rect 1406 4028 1407 4032
rect 1411 4028 1412 4032
rect 1406 4027 1412 4028
rect 1542 4032 1548 4033
rect 1542 4028 1543 4032
rect 1547 4028 1548 4032
rect 1542 4027 1548 4028
rect 1678 4032 1684 4033
rect 1678 4028 1679 4032
rect 1683 4028 1684 4032
rect 1678 4027 1684 4028
rect 1814 4032 1820 4033
rect 1814 4028 1815 4032
rect 1819 4028 1820 4032
rect 1814 4027 1820 4028
rect 1934 4031 1940 4032
rect 1934 4027 1935 4031
rect 1939 4027 1940 4031
rect 3858 4029 3864 4030
rect 110 4026 116 4027
rect 1934 4026 1940 4027
rect 3838 4028 3844 4029
rect 3838 4024 3839 4028
rect 3843 4024 3844 4028
rect 3858 4025 3859 4029
rect 3863 4025 3864 4029
rect 3858 4024 3864 4025
rect 3994 4029 4000 4030
rect 3994 4025 3995 4029
rect 3999 4025 4000 4029
rect 3994 4024 4000 4025
rect 4130 4029 4136 4030
rect 4130 4025 4131 4029
rect 4135 4025 4136 4029
rect 4130 4024 4136 4025
rect 4266 4029 4272 4030
rect 4266 4025 4267 4029
rect 4271 4025 4272 4029
rect 4266 4024 4272 4025
rect 4402 4029 4408 4030
rect 4402 4025 4403 4029
rect 4407 4025 4408 4029
rect 4402 4024 4408 4025
rect 4538 4029 4544 4030
rect 4538 4025 4539 4029
rect 4543 4025 4544 4029
rect 4538 4024 4544 4025
rect 4674 4029 4680 4030
rect 4674 4025 4675 4029
rect 4679 4025 4680 4029
rect 4674 4024 4680 4025
rect 4810 4029 4816 4030
rect 4810 4025 4811 4029
rect 4815 4025 4816 4029
rect 4810 4024 4816 4025
rect 5662 4028 5668 4029
rect 5662 4024 5663 4028
rect 5667 4024 5668 4028
rect 3838 4023 3844 4024
rect 5662 4023 5668 4024
rect 110 3973 116 3974
rect 1934 3973 1940 3974
rect 110 3969 111 3973
rect 115 3969 116 3973
rect 110 3968 116 3969
rect 158 3972 164 3973
rect 158 3968 159 3972
rect 163 3968 164 3972
rect 158 3967 164 3968
rect 326 3972 332 3973
rect 326 3968 327 3972
rect 331 3968 332 3972
rect 326 3967 332 3968
rect 534 3972 540 3973
rect 534 3968 535 3972
rect 539 3968 540 3972
rect 534 3967 540 3968
rect 750 3972 756 3973
rect 750 3968 751 3972
rect 755 3968 756 3972
rect 750 3967 756 3968
rect 966 3972 972 3973
rect 966 3968 967 3972
rect 971 3968 972 3972
rect 966 3967 972 3968
rect 1182 3972 1188 3973
rect 1182 3968 1183 3972
rect 1187 3968 1188 3972
rect 1182 3967 1188 3968
rect 1398 3972 1404 3973
rect 1398 3968 1399 3972
rect 1403 3968 1404 3972
rect 1398 3967 1404 3968
rect 1614 3972 1620 3973
rect 1614 3968 1615 3972
rect 1619 3968 1620 3972
rect 1614 3967 1620 3968
rect 1814 3972 1820 3973
rect 1814 3968 1815 3972
rect 1819 3968 1820 3972
rect 1934 3969 1935 3973
rect 1939 3969 1940 3973
rect 1934 3968 1940 3969
rect 1814 3967 1820 3968
rect 130 3957 136 3958
rect 110 3956 116 3957
rect 110 3952 111 3956
rect 115 3952 116 3956
rect 130 3953 131 3957
rect 135 3953 136 3957
rect 130 3952 136 3953
rect 298 3957 304 3958
rect 298 3953 299 3957
rect 303 3953 304 3957
rect 298 3952 304 3953
rect 506 3957 512 3958
rect 506 3953 507 3957
rect 511 3953 512 3957
rect 506 3952 512 3953
rect 722 3957 728 3958
rect 722 3953 723 3957
rect 727 3953 728 3957
rect 722 3952 728 3953
rect 938 3957 944 3958
rect 938 3953 939 3957
rect 943 3953 944 3957
rect 938 3952 944 3953
rect 1154 3957 1160 3958
rect 1154 3953 1155 3957
rect 1159 3953 1160 3957
rect 1154 3952 1160 3953
rect 1370 3957 1376 3958
rect 1370 3953 1371 3957
rect 1375 3953 1376 3957
rect 1370 3952 1376 3953
rect 1586 3957 1592 3958
rect 1586 3953 1587 3957
rect 1591 3953 1592 3957
rect 1586 3952 1592 3953
rect 1786 3957 1792 3958
rect 1786 3953 1787 3957
rect 1791 3953 1792 3957
rect 1786 3952 1792 3953
rect 1934 3956 1940 3957
rect 1934 3952 1935 3956
rect 1939 3952 1940 3956
rect 110 3951 116 3952
rect 1934 3951 1940 3952
rect 3838 3896 3844 3897
rect 5662 3896 5668 3897
rect 3838 3892 3839 3896
rect 3843 3892 3844 3896
rect 3838 3891 3844 3892
rect 3858 3895 3864 3896
rect 3858 3891 3859 3895
rect 3863 3891 3864 3895
rect 3858 3890 3864 3891
rect 3994 3895 4000 3896
rect 3994 3891 3995 3895
rect 3999 3891 4000 3895
rect 3994 3890 4000 3891
rect 4146 3895 4152 3896
rect 4146 3891 4147 3895
rect 4151 3891 4152 3895
rect 4146 3890 4152 3891
rect 4298 3895 4304 3896
rect 4298 3891 4299 3895
rect 4303 3891 4304 3895
rect 4298 3890 4304 3891
rect 4458 3895 4464 3896
rect 4458 3891 4459 3895
rect 4463 3891 4464 3895
rect 4458 3890 4464 3891
rect 4618 3895 4624 3896
rect 4618 3891 4619 3895
rect 4623 3891 4624 3895
rect 4618 3890 4624 3891
rect 4778 3895 4784 3896
rect 4778 3891 4779 3895
rect 4783 3891 4784 3895
rect 5662 3892 5663 3896
rect 5667 3892 5668 3896
rect 5662 3891 5668 3892
rect 4778 3890 4784 3891
rect 3886 3880 3892 3881
rect 3838 3879 3844 3880
rect 3838 3875 3839 3879
rect 3843 3875 3844 3879
rect 3886 3876 3887 3880
rect 3891 3876 3892 3880
rect 3886 3875 3892 3876
rect 4022 3880 4028 3881
rect 4022 3876 4023 3880
rect 4027 3876 4028 3880
rect 4022 3875 4028 3876
rect 4174 3880 4180 3881
rect 4174 3876 4175 3880
rect 4179 3876 4180 3880
rect 4174 3875 4180 3876
rect 4326 3880 4332 3881
rect 4326 3876 4327 3880
rect 4331 3876 4332 3880
rect 4326 3875 4332 3876
rect 4486 3880 4492 3881
rect 4486 3876 4487 3880
rect 4491 3876 4492 3880
rect 4486 3875 4492 3876
rect 4646 3880 4652 3881
rect 4646 3876 4647 3880
rect 4651 3876 4652 3880
rect 4646 3875 4652 3876
rect 4806 3880 4812 3881
rect 4806 3876 4807 3880
rect 4811 3876 4812 3880
rect 4806 3875 4812 3876
rect 5662 3879 5668 3880
rect 5662 3875 5663 3879
rect 5667 3875 5668 3879
rect 3838 3874 3844 3875
rect 5662 3874 5668 3875
rect 1974 3868 1980 3869
rect 3798 3868 3804 3869
rect 1974 3864 1975 3868
rect 1979 3864 1980 3868
rect 1974 3863 1980 3864
rect 1994 3867 2000 3868
rect 1994 3863 1995 3867
rect 1999 3863 2000 3867
rect 1994 3862 2000 3863
rect 2402 3867 2408 3868
rect 2402 3863 2403 3867
rect 2407 3863 2408 3867
rect 2402 3862 2408 3863
rect 2826 3867 2832 3868
rect 2826 3863 2827 3867
rect 2831 3863 2832 3867
rect 2826 3862 2832 3863
rect 3250 3867 3256 3868
rect 3250 3863 3251 3867
rect 3255 3863 3256 3867
rect 3250 3862 3256 3863
rect 3650 3867 3656 3868
rect 3650 3863 3651 3867
rect 3655 3863 3656 3867
rect 3798 3864 3799 3868
rect 3803 3864 3804 3868
rect 3798 3863 3804 3864
rect 3650 3862 3656 3863
rect 2022 3852 2028 3853
rect 1974 3851 1980 3852
rect 1974 3847 1975 3851
rect 1979 3847 1980 3851
rect 2022 3848 2023 3852
rect 2027 3848 2028 3852
rect 2022 3847 2028 3848
rect 2430 3852 2436 3853
rect 2430 3848 2431 3852
rect 2435 3848 2436 3852
rect 2430 3847 2436 3848
rect 2854 3852 2860 3853
rect 2854 3848 2855 3852
rect 2859 3848 2860 3852
rect 2854 3847 2860 3848
rect 3278 3852 3284 3853
rect 3278 3848 3279 3852
rect 3283 3848 3284 3852
rect 3278 3847 3284 3848
rect 3678 3852 3684 3853
rect 3678 3848 3679 3852
rect 3683 3848 3684 3852
rect 3678 3847 3684 3848
rect 3798 3851 3804 3852
rect 3798 3847 3799 3851
rect 3803 3847 3804 3851
rect 1974 3846 1980 3847
rect 3798 3846 3804 3847
rect 110 3824 116 3825
rect 1934 3824 1940 3825
rect 110 3820 111 3824
rect 115 3820 116 3824
rect 110 3819 116 3820
rect 130 3823 136 3824
rect 130 3819 131 3823
rect 135 3819 136 3823
rect 130 3818 136 3819
rect 354 3823 360 3824
rect 354 3819 355 3823
rect 359 3819 360 3823
rect 354 3818 360 3819
rect 618 3823 624 3824
rect 618 3819 619 3823
rect 623 3819 624 3823
rect 618 3818 624 3819
rect 898 3823 904 3824
rect 898 3819 899 3823
rect 903 3819 904 3823
rect 898 3818 904 3819
rect 1194 3823 1200 3824
rect 1194 3819 1195 3823
rect 1199 3819 1200 3823
rect 1194 3818 1200 3819
rect 1498 3823 1504 3824
rect 1498 3819 1499 3823
rect 1503 3819 1504 3823
rect 1498 3818 1504 3819
rect 1786 3823 1792 3824
rect 1786 3819 1787 3823
rect 1791 3819 1792 3823
rect 1934 3820 1935 3824
rect 1939 3820 1940 3824
rect 1934 3819 1940 3820
rect 1786 3818 1792 3819
rect 158 3808 164 3809
rect 110 3807 116 3808
rect 110 3803 111 3807
rect 115 3803 116 3807
rect 158 3804 159 3808
rect 163 3804 164 3808
rect 158 3803 164 3804
rect 382 3808 388 3809
rect 382 3804 383 3808
rect 387 3804 388 3808
rect 382 3803 388 3804
rect 646 3808 652 3809
rect 646 3804 647 3808
rect 651 3804 652 3808
rect 646 3803 652 3804
rect 926 3808 932 3809
rect 926 3804 927 3808
rect 931 3804 932 3808
rect 926 3803 932 3804
rect 1222 3808 1228 3809
rect 1222 3804 1223 3808
rect 1227 3804 1228 3808
rect 1222 3803 1228 3804
rect 1526 3808 1532 3809
rect 1526 3804 1527 3808
rect 1531 3804 1532 3808
rect 1526 3803 1532 3804
rect 1814 3808 1820 3809
rect 1814 3804 1815 3808
rect 1819 3804 1820 3808
rect 1814 3803 1820 3804
rect 1934 3807 1940 3808
rect 1934 3803 1935 3807
rect 1939 3803 1940 3807
rect 110 3802 116 3803
rect 1934 3802 1940 3803
rect 1974 3793 1980 3794
rect 3798 3793 3804 3794
rect 1974 3789 1975 3793
rect 1979 3789 1980 3793
rect 1974 3788 1980 3789
rect 2022 3792 2028 3793
rect 2022 3788 2023 3792
rect 2027 3788 2028 3792
rect 2022 3787 2028 3788
rect 2174 3792 2180 3793
rect 2174 3788 2175 3792
rect 2179 3788 2180 3792
rect 2174 3787 2180 3788
rect 2350 3792 2356 3793
rect 2350 3788 2351 3792
rect 2355 3788 2356 3792
rect 2350 3787 2356 3788
rect 2534 3792 2540 3793
rect 2534 3788 2535 3792
rect 2539 3788 2540 3792
rect 2534 3787 2540 3788
rect 2718 3792 2724 3793
rect 2718 3788 2719 3792
rect 2723 3788 2724 3792
rect 2718 3787 2724 3788
rect 2894 3792 2900 3793
rect 2894 3788 2895 3792
rect 2899 3788 2900 3792
rect 2894 3787 2900 3788
rect 3070 3792 3076 3793
rect 3070 3788 3071 3792
rect 3075 3788 3076 3792
rect 3070 3787 3076 3788
rect 3246 3792 3252 3793
rect 3246 3788 3247 3792
rect 3251 3788 3252 3792
rect 3246 3787 3252 3788
rect 3422 3792 3428 3793
rect 3422 3788 3423 3792
rect 3427 3788 3428 3792
rect 3422 3787 3428 3788
rect 3606 3792 3612 3793
rect 3606 3788 3607 3792
rect 3611 3788 3612 3792
rect 3798 3789 3799 3793
rect 3803 3789 3804 3793
rect 3798 3788 3804 3789
rect 3838 3793 3844 3794
rect 5662 3793 5668 3794
rect 3838 3789 3839 3793
rect 3843 3789 3844 3793
rect 3838 3788 3844 3789
rect 4502 3792 4508 3793
rect 4502 3788 4503 3792
rect 4507 3788 4508 3792
rect 3606 3787 3612 3788
rect 4502 3787 4508 3788
rect 4638 3792 4644 3793
rect 4638 3788 4639 3792
rect 4643 3788 4644 3792
rect 4638 3787 4644 3788
rect 4774 3792 4780 3793
rect 4774 3788 4775 3792
rect 4779 3788 4780 3792
rect 4774 3787 4780 3788
rect 4910 3792 4916 3793
rect 4910 3788 4911 3792
rect 4915 3788 4916 3792
rect 4910 3787 4916 3788
rect 5046 3792 5052 3793
rect 5046 3788 5047 3792
rect 5051 3788 5052 3792
rect 5662 3789 5663 3793
rect 5667 3789 5668 3793
rect 5662 3788 5668 3789
rect 5046 3787 5052 3788
rect 1994 3777 2000 3778
rect 1974 3776 1980 3777
rect 1974 3772 1975 3776
rect 1979 3772 1980 3776
rect 1994 3773 1995 3777
rect 1999 3773 2000 3777
rect 1994 3772 2000 3773
rect 2146 3777 2152 3778
rect 2146 3773 2147 3777
rect 2151 3773 2152 3777
rect 2146 3772 2152 3773
rect 2322 3777 2328 3778
rect 2322 3773 2323 3777
rect 2327 3773 2328 3777
rect 2322 3772 2328 3773
rect 2506 3777 2512 3778
rect 2506 3773 2507 3777
rect 2511 3773 2512 3777
rect 2506 3772 2512 3773
rect 2690 3777 2696 3778
rect 2690 3773 2691 3777
rect 2695 3773 2696 3777
rect 2690 3772 2696 3773
rect 2866 3777 2872 3778
rect 2866 3773 2867 3777
rect 2871 3773 2872 3777
rect 2866 3772 2872 3773
rect 3042 3777 3048 3778
rect 3042 3773 3043 3777
rect 3047 3773 3048 3777
rect 3042 3772 3048 3773
rect 3218 3777 3224 3778
rect 3218 3773 3219 3777
rect 3223 3773 3224 3777
rect 3218 3772 3224 3773
rect 3394 3777 3400 3778
rect 3394 3773 3395 3777
rect 3399 3773 3400 3777
rect 3394 3772 3400 3773
rect 3578 3777 3584 3778
rect 4474 3777 4480 3778
rect 3578 3773 3579 3777
rect 3583 3773 3584 3777
rect 3578 3772 3584 3773
rect 3798 3776 3804 3777
rect 3798 3772 3799 3776
rect 3803 3772 3804 3776
rect 1974 3771 1980 3772
rect 3798 3771 3804 3772
rect 3838 3776 3844 3777
rect 3838 3772 3839 3776
rect 3843 3772 3844 3776
rect 4474 3773 4475 3777
rect 4479 3773 4480 3777
rect 4474 3772 4480 3773
rect 4610 3777 4616 3778
rect 4610 3773 4611 3777
rect 4615 3773 4616 3777
rect 4610 3772 4616 3773
rect 4746 3777 4752 3778
rect 4746 3773 4747 3777
rect 4751 3773 4752 3777
rect 4746 3772 4752 3773
rect 4882 3777 4888 3778
rect 4882 3773 4883 3777
rect 4887 3773 4888 3777
rect 4882 3772 4888 3773
rect 5018 3777 5024 3778
rect 5018 3773 5019 3777
rect 5023 3773 5024 3777
rect 5018 3772 5024 3773
rect 5662 3776 5668 3777
rect 5662 3772 5663 3776
rect 5667 3772 5668 3776
rect 3838 3771 3844 3772
rect 5662 3771 5668 3772
rect 110 3737 116 3738
rect 1934 3737 1940 3738
rect 110 3733 111 3737
rect 115 3733 116 3737
rect 110 3732 116 3733
rect 246 3736 252 3737
rect 246 3732 247 3736
rect 251 3732 252 3736
rect 246 3731 252 3732
rect 518 3736 524 3737
rect 518 3732 519 3736
rect 523 3732 524 3736
rect 518 3731 524 3732
rect 790 3736 796 3737
rect 790 3732 791 3736
rect 795 3732 796 3736
rect 790 3731 796 3732
rect 1062 3736 1068 3737
rect 1062 3732 1063 3736
rect 1067 3732 1068 3736
rect 1062 3731 1068 3732
rect 1342 3736 1348 3737
rect 1342 3732 1343 3736
rect 1347 3732 1348 3736
rect 1934 3733 1935 3737
rect 1939 3733 1940 3737
rect 1934 3732 1940 3733
rect 1342 3731 1348 3732
rect 218 3721 224 3722
rect 110 3720 116 3721
rect 110 3716 111 3720
rect 115 3716 116 3720
rect 218 3717 219 3721
rect 223 3717 224 3721
rect 218 3716 224 3717
rect 490 3721 496 3722
rect 490 3717 491 3721
rect 495 3717 496 3721
rect 490 3716 496 3717
rect 762 3721 768 3722
rect 762 3717 763 3721
rect 767 3717 768 3721
rect 762 3716 768 3717
rect 1034 3721 1040 3722
rect 1034 3717 1035 3721
rect 1039 3717 1040 3721
rect 1034 3716 1040 3717
rect 1314 3721 1320 3722
rect 1314 3717 1315 3721
rect 1319 3717 1320 3721
rect 1314 3716 1320 3717
rect 1934 3720 1940 3721
rect 1934 3716 1935 3720
rect 1939 3716 1940 3720
rect 110 3715 116 3716
rect 1934 3715 1940 3716
rect 1974 3636 1980 3637
rect 3798 3636 3804 3637
rect 1974 3632 1975 3636
rect 1979 3632 1980 3636
rect 1974 3631 1980 3632
rect 2010 3635 2016 3636
rect 2010 3631 2011 3635
rect 2015 3631 2016 3635
rect 2010 3630 2016 3631
rect 2146 3635 2152 3636
rect 2146 3631 2147 3635
rect 2151 3631 2152 3635
rect 2146 3630 2152 3631
rect 2290 3635 2296 3636
rect 2290 3631 2291 3635
rect 2295 3631 2296 3635
rect 2290 3630 2296 3631
rect 2434 3635 2440 3636
rect 2434 3631 2435 3635
rect 2439 3631 2440 3635
rect 2434 3630 2440 3631
rect 2578 3635 2584 3636
rect 2578 3631 2579 3635
rect 2583 3631 2584 3635
rect 2578 3630 2584 3631
rect 2722 3635 2728 3636
rect 2722 3631 2723 3635
rect 2727 3631 2728 3635
rect 2722 3630 2728 3631
rect 2866 3635 2872 3636
rect 2866 3631 2867 3635
rect 2871 3631 2872 3635
rect 2866 3630 2872 3631
rect 3010 3635 3016 3636
rect 3010 3631 3011 3635
rect 3015 3631 3016 3635
rect 3010 3630 3016 3631
rect 3154 3635 3160 3636
rect 3154 3631 3155 3635
rect 3159 3631 3160 3635
rect 3154 3630 3160 3631
rect 3298 3635 3304 3636
rect 3298 3631 3299 3635
rect 3303 3631 3304 3635
rect 3798 3632 3799 3636
rect 3803 3632 3804 3636
rect 3798 3631 3804 3632
rect 3298 3630 3304 3631
rect 3838 3624 3844 3625
rect 5662 3624 5668 3625
rect 2038 3620 2044 3621
rect 1974 3619 1980 3620
rect 1974 3615 1975 3619
rect 1979 3615 1980 3619
rect 2038 3616 2039 3620
rect 2043 3616 2044 3620
rect 2038 3615 2044 3616
rect 2174 3620 2180 3621
rect 2174 3616 2175 3620
rect 2179 3616 2180 3620
rect 2174 3615 2180 3616
rect 2318 3620 2324 3621
rect 2318 3616 2319 3620
rect 2323 3616 2324 3620
rect 2318 3615 2324 3616
rect 2462 3620 2468 3621
rect 2462 3616 2463 3620
rect 2467 3616 2468 3620
rect 2462 3615 2468 3616
rect 2606 3620 2612 3621
rect 2606 3616 2607 3620
rect 2611 3616 2612 3620
rect 2606 3615 2612 3616
rect 2750 3620 2756 3621
rect 2750 3616 2751 3620
rect 2755 3616 2756 3620
rect 2750 3615 2756 3616
rect 2894 3620 2900 3621
rect 2894 3616 2895 3620
rect 2899 3616 2900 3620
rect 2894 3615 2900 3616
rect 3038 3620 3044 3621
rect 3038 3616 3039 3620
rect 3043 3616 3044 3620
rect 3038 3615 3044 3616
rect 3182 3620 3188 3621
rect 3182 3616 3183 3620
rect 3187 3616 3188 3620
rect 3182 3615 3188 3616
rect 3326 3620 3332 3621
rect 3838 3620 3839 3624
rect 3843 3620 3844 3624
rect 3326 3616 3327 3620
rect 3331 3616 3332 3620
rect 3326 3615 3332 3616
rect 3798 3619 3804 3620
rect 3838 3619 3844 3620
rect 4018 3623 4024 3624
rect 4018 3619 4019 3623
rect 4023 3619 4024 3623
rect 3798 3615 3799 3619
rect 3803 3615 3804 3619
rect 4018 3618 4024 3619
rect 4154 3623 4160 3624
rect 4154 3619 4155 3623
rect 4159 3619 4160 3623
rect 4154 3618 4160 3619
rect 4290 3623 4296 3624
rect 4290 3619 4291 3623
rect 4295 3619 4296 3623
rect 4290 3618 4296 3619
rect 4426 3623 4432 3624
rect 4426 3619 4427 3623
rect 4431 3619 4432 3623
rect 4426 3618 4432 3619
rect 4562 3623 4568 3624
rect 4562 3619 4563 3623
rect 4567 3619 4568 3623
rect 4562 3618 4568 3619
rect 4698 3623 4704 3624
rect 4698 3619 4699 3623
rect 4703 3619 4704 3623
rect 4698 3618 4704 3619
rect 4834 3623 4840 3624
rect 4834 3619 4835 3623
rect 4839 3619 4840 3623
rect 4834 3618 4840 3619
rect 4970 3623 4976 3624
rect 4970 3619 4971 3623
rect 4975 3619 4976 3623
rect 4970 3618 4976 3619
rect 5106 3623 5112 3624
rect 5106 3619 5107 3623
rect 5111 3619 5112 3623
rect 5106 3618 5112 3619
rect 5242 3623 5248 3624
rect 5242 3619 5243 3623
rect 5247 3619 5248 3623
rect 5242 3618 5248 3619
rect 5378 3623 5384 3624
rect 5378 3619 5379 3623
rect 5383 3619 5384 3623
rect 5378 3618 5384 3619
rect 5514 3623 5520 3624
rect 5514 3619 5515 3623
rect 5519 3619 5520 3623
rect 5662 3620 5663 3624
rect 5667 3620 5668 3624
rect 5662 3619 5668 3620
rect 5514 3618 5520 3619
rect 1974 3614 1980 3615
rect 3798 3614 3804 3615
rect 4046 3608 4052 3609
rect 3838 3607 3844 3608
rect 3838 3603 3839 3607
rect 3843 3603 3844 3607
rect 4046 3604 4047 3608
rect 4051 3604 4052 3608
rect 4046 3603 4052 3604
rect 4182 3608 4188 3609
rect 4182 3604 4183 3608
rect 4187 3604 4188 3608
rect 4182 3603 4188 3604
rect 4318 3608 4324 3609
rect 4318 3604 4319 3608
rect 4323 3604 4324 3608
rect 4318 3603 4324 3604
rect 4454 3608 4460 3609
rect 4454 3604 4455 3608
rect 4459 3604 4460 3608
rect 4454 3603 4460 3604
rect 4590 3608 4596 3609
rect 4590 3604 4591 3608
rect 4595 3604 4596 3608
rect 4590 3603 4596 3604
rect 4726 3608 4732 3609
rect 4726 3604 4727 3608
rect 4731 3604 4732 3608
rect 4726 3603 4732 3604
rect 4862 3608 4868 3609
rect 4862 3604 4863 3608
rect 4867 3604 4868 3608
rect 4862 3603 4868 3604
rect 4998 3608 5004 3609
rect 4998 3604 4999 3608
rect 5003 3604 5004 3608
rect 4998 3603 5004 3604
rect 5134 3608 5140 3609
rect 5134 3604 5135 3608
rect 5139 3604 5140 3608
rect 5134 3603 5140 3604
rect 5270 3608 5276 3609
rect 5270 3604 5271 3608
rect 5275 3604 5276 3608
rect 5270 3603 5276 3604
rect 5406 3608 5412 3609
rect 5406 3604 5407 3608
rect 5411 3604 5412 3608
rect 5406 3603 5412 3604
rect 5542 3608 5548 3609
rect 5542 3604 5543 3608
rect 5547 3604 5548 3608
rect 5542 3603 5548 3604
rect 5662 3607 5668 3608
rect 5662 3603 5663 3607
rect 5667 3603 5668 3607
rect 3838 3602 3844 3603
rect 5662 3602 5668 3603
rect 110 3572 116 3573
rect 1934 3572 1940 3573
rect 110 3568 111 3572
rect 115 3568 116 3572
rect 110 3567 116 3568
rect 490 3571 496 3572
rect 490 3567 491 3571
rect 495 3567 496 3571
rect 490 3566 496 3567
rect 634 3571 640 3572
rect 634 3567 635 3571
rect 639 3567 640 3571
rect 634 3566 640 3567
rect 778 3571 784 3572
rect 778 3567 779 3571
rect 783 3567 784 3571
rect 778 3566 784 3567
rect 922 3571 928 3572
rect 922 3567 923 3571
rect 927 3567 928 3571
rect 922 3566 928 3567
rect 1066 3571 1072 3572
rect 1066 3567 1067 3571
rect 1071 3567 1072 3571
rect 1066 3566 1072 3567
rect 1210 3571 1216 3572
rect 1210 3567 1211 3571
rect 1215 3567 1216 3571
rect 1934 3568 1935 3572
rect 1939 3568 1940 3572
rect 1934 3567 1940 3568
rect 1210 3566 1216 3567
rect 518 3556 524 3557
rect 110 3555 116 3556
rect 110 3551 111 3555
rect 115 3551 116 3555
rect 518 3552 519 3556
rect 523 3552 524 3556
rect 518 3551 524 3552
rect 662 3556 668 3557
rect 662 3552 663 3556
rect 667 3552 668 3556
rect 662 3551 668 3552
rect 806 3556 812 3557
rect 806 3552 807 3556
rect 811 3552 812 3556
rect 806 3551 812 3552
rect 950 3556 956 3557
rect 950 3552 951 3556
rect 955 3552 956 3556
rect 950 3551 956 3552
rect 1094 3556 1100 3557
rect 1094 3552 1095 3556
rect 1099 3552 1100 3556
rect 1094 3551 1100 3552
rect 1238 3556 1244 3557
rect 1238 3552 1239 3556
rect 1243 3552 1244 3556
rect 1238 3551 1244 3552
rect 1934 3555 1940 3556
rect 1934 3551 1935 3555
rect 1939 3551 1940 3555
rect 110 3550 116 3551
rect 1934 3550 1940 3551
rect 1974 3553 1980 3554
rect 3798 3553 3804 3554
rect 1974 3549 1975 3553
rect 1979 3549 1980 3553
rect 1974 3548 1980 3549
rect 2238 3552 2244 3553
rect 2238 3548 2239 3552
rect 2243 3548 2244 3552
rect 2238 3547 2244 3548
rect 2374 3552 2380 3553
rect 2374 3548 2375 3552
rect 2379 3548 2380 3552
rect 2374 3547 2380 3548
rect 2510 3552 2516 3553
rect 2510 3548 2511 3552
rect 2515 3548 2516 3552
rect 2510 3547 2516 3548
rect 2646 3552 2652 3553
rect 2646 3548 2647 3552
rect 2651 3548 2652 3552
rect 2646 3547 2652 3548
rect 2782 3552 2788 3553
rect 2782 3548 2783 3552
rect 2787 3548 2788 3552
rect 2782 3547 2788 3548
rect 2918 3552 2924 3553
rect 2918 3548 2919 3552
rect 2923 3548 2924 3552
rect 2918 3547 2924 3548
rect 3054 3552 3060 3553
rect 3054 3548 3055 3552
rect 3059 3548 3060 3552
rect 3054 3547 3060 3548
rect 3190 3552 3196 3553
rect 3190 3548 3191 3552
rect 3195 3548 3196 3552
rect 3190 3547 3196 3548
rect 3326 3552 3332 3553
rect 3326 3548 3327 3552
rect 3331 3548 3332 3552
rect 3326 3547 3332 3548
rect 3462 3552 3468 3553
rect 3462 3548 3463 3552
rect 3467 3548 3468 3552
rect 3798 3549 3799 3553
rect 3803 3549 3804 3553
rect 3798 3548 3804 3549
rect 3462 3547 3468 3548
rect 2210 3537 2216 3538
rect 1974 3536 1980 3537
rect 1974 3532 1975 3536
rect 1979 3532 1980 3536
rect 2210 3533 2211 3537
rect 2215 3533 2216 3537
rect 2210 3532 2216 3533
rect 2346 3537 2352 3538
rect 2346 3533 2347 3537
rect 2351 3533 2352 3537
rect 2346 3532 2352 3533
rect 2482 3537 2488 3538
rect 2482 3533 2483 3537
rect 2487 3533 2488 3537
rect 2482 3532 2488 3533
rect 2618 3537 2624 3538
rect 2618 3533 2619 3537
rect 2623 3533 2624 3537
rect 2618 3532 2624 3533
rect 2754 3537 2760 3538
rect 2754 3533 2755 3537
rect 2759 3533 2760 3537
rect 2754 3532 2760 3533
rect 2890 3537 2896 3538
rect 2890 3533 2891 3537
rect 2895 3533 2896 3537
rect 2890 3532 2896 3533
rect 3026 3537 3032 3538
rect 3026 3533 3027 3537
rect 3031 3533 3032 3537
rect 3026 3532 3032 3533
rect 3162 3537 3168 3538
rect 3162 3533 3163 3537
rect 3167 3533 3168 3537
rect 3162 3532 3168 3533
rect 3298 3537 3304 3538
rect 3298 3533 3299 3537
rect 3303 3533 3304 3537
rect 3298 3532 3304 3533
rect 3434 3537 3440 3538
rect 3434 3533 3435 3537
rect 3439 3533 3440 3537
rect 3434 3532 3440 3533
rect 3798 3536 3804 3537
rect 3798 3532 3799 3536
rect 3803 3532 3804 3536
rect 1974 3531 1980 3532
rect 3798 3531 3804 3532
rect 3838 3501 3844 3502
rect 5662 3501 5668 3502
rect 3838 3497 3839 3501
rect 3843 3497 3844 3501
rect 3838 3496 3844 3497
rect 5406 3500 5412 3501
rect 5406 3496 5407 3500
rect 5411 3496 5412 3500
rect 5406 3495 5412 3496
rect 5542 3500 5548 3501
rect 5542 3496 5543 3500
rect 5547 3496 5548 3500
rect 5662 3497 5663 3501
rect 5667 3497 5668 3501
rect 5662 3496 5668 3497
rect 5542 3495 5548 3496
rect 5378 3485 5384 3486
rect 3838 3484 3844 3485
rect 3838 3480 3839 3484
rect 3843 3480 3844 3484
rect 5378 3481 5379 3485
rect 5383 3481 5384 3485
rect 5378 3480 5384 3481
rect 5514 3485 5520 3486
rect 5514 3481 5515 3485
rect 5519 3481 5520 3485
rect 5514 3480 5520 3481
rect 5662 3484 5668 3485
rect 5662 3480 5663 3484
rect 5667 3480 5668 3484
rect 3838 3479 3844 3480
rect 5662 3479 5668 3480
rect 110 3477 116 3478
rect 1934 3477 1940 3478
rect 110 3473 111 3477
rect 115 3473 116 3477
rect 110 3472 116 3473
rect 430 3476 436 3477
rect 430 3472 431 3476
rect 435 3472 436 3476
rect 430 3471 436 3472
rect 566 3476 572 3477
rect 566 3472 567 3476
rect 571 3472 572 3476
rect 566 3471 572 3472
rect 702 3476 708 3477
rect 702 3472 703 3476
rect 707 3472 708 3476
rect 702 3471 708 3472
rect 838 3476 844 3477
rect 838 3472 839 3476
rect 843 3472 844 3476
rect 838 3471 844 3472
rect 974 3476 980 3477
rect 974 3472 975 3476
rect 979 3472 980 3476
rect 1934 3473 1935 3477
rect 1939 3473 1940 3477
rect 1934 3472 1940 3473
rect 974 3471 980 3472
rect 402 3461 408 3462
rect 110 3460 116 3461
rect 110 3456 111 3460
rect 115 3456 116 3460
rect 402 3457 403 3461
rect 407 3457 408 3461
rect 402 3456 408 3457
rect 538 3461 544 3462
rect 538 3457 539 3461
rect 543 3457 544 3461
rect 538 3456 544 3457
rect 674 3461 680 3462
rect 674 3457 675 3461
rect 679 3457 680 3461
rect 674 3456 680 3457
rect 810 3461 816 3462
rect 810 3457 811 3461
rect 815 3457 816 3461
rect 810 3456 816 3457
rect 946 3461 952 3462
rect 946 3457 947 3461
rect 951 3457 952 3461
rect 946 3456 952 3457
rect 1934 3460 1940 3461
rect 1934 3456 1935 3460
rect 1939 3456 1940 3460
rect 110 3455 116 3456
rect 1934 3455 1940 3456
rect 1974 3400 1980 3401
rect 3798 3400 3804 3401
rect 1974 3396 1975 3400
rect 1979 3396 1980 3400
rect 1974 3395 1980 3396
rect 2170 3399 2176 3400
rect 2170 3395 2171 3399
rect 2175 3395 2176 3399
rect 2170 3394 2176 3395
rect 2346 3399 2352 3400
rect 2346 3395 2347 3399
rect 2351 3395 2352 3399
rect 2346 3394 2352 3395
rect 2530 3399 2536 3400
rect 2530 3395 2531 3399
rect 2535 3395 2536 3399
rect 2530 3394 2536 3395
rect 2714 3399 2720 3400
rect 2714 3395 2715 3399
rect 2719 3395 2720 3399
rect 2714 3394 2720 3395
rect 2906 3399 2912 3400
rect 2906 3395 2907 3399
rect 2911 3395 2912 3399
rect 2906 3394 2912 3395
rect 3098 3399 3104 3400
rect 3098 3395 3099 3399
rect 3103 3395 3104 3399
rect 3098 3394 3104 3395
rect 3290 3399 3296 3400
rect 3290 3395 3291 3399
rect 3295 3395 3296 3399
rect 3290 3394 3296 3395
rect 3482 3399 3488 3400
rect 3482 3395 3483 3399
rect 3487 3395 3488 3399
rect 3482 3394 3488 3395
rect 3650 3399 3656 3400
rect 3650 3395 3651 3399
rect 3655 3395 3656 3399
rect 3798 3396 3799 3400
rect 3803 3396 3804 3400
rect 3798 3395 3804 3396
rect 3650 3394 3656 3395
rect 2198 3384 2204 3385
rect 1974 3383 1980 3384
rect 1974 3379 1975 3383
rect 1979 3379 1980 3383
rect 2198 3380 2199 3384
rect 2203 3380 2204 3384
rect 2198 3379 2204 3380
rect 2374 3384 2380 3385
rect 2374 3380 2375 3384
rect 2379 3380 2380 3384
rect 2374 3379 2380 3380
rect 2558 3384 2564 3385
rect 2558 3380 2559 3384
rect 2563 3380 2564 3384
rect 2558 3379 2564 3380
rect 2742 3384 2748 3385
rect 2742 3380 2743 3384
rect 2747 3380 2748 3384
rect 2742 3379 2748 3380
rect 2934 3384 2940 3385
rect 2934 3380 2935 3384
rect 2939 3380 2940 3384
rect 2934 3379 2940 3380
rect 3126 3384 3132 3385
rect 3126 3380 3127 3384
rect 3131 3380 3132 3384
rect 3126 3379 3132 3380
rect 3318 3384 3324 3385
rect 3318 3380 3319 3384
rect 3323 3380 3324 3384
rect 3318 3379 3324 3380
rect 3510 3384 3516 3385
rect 3510 3380 3511 3384
rect 3515 3380 3516 3384
rect 3510 3379 3516 3380
rect 3678 3384 3684 3385
rect 3678 3380 3679 3384
rect 3683 3380 3684 3384
rect 3678 3379 3684 3380
rect 3798 3383 3804 3384
rect 3798 3379 3799 3383
rect 3803 3379 3804 3383
rect 1974 3378 1980 3379
rect 3798 3378 3804 3379
rect 3838 3344 3844 3345
rect 5662 3344 5668 3345
rect 3838 3340 3839 3344
rect 3843 3340 3844 3344
rect 3838 3339 3844 3340
rect 3858 3343 3864 3344
rect 3858 3339 3859 3343
rect 3863 3339 3864 3343
rect 3858 3338 3864 3339
rect 4098 3343 4104 3344
rect 4098 3339 4099 3343
rect 4103 3339 4104 3343
rect 4098 3338 4104 3339
rect 4346 3343 4352 3344
rect 4346 3339 4347 3343
rect 4351 3339 4352 3343
rect 4346 3338 4352 3339
rect 4586 3343 4592 3344
rect 4586 3339 4587 3343
rect 4591 3339 4592 3343
rect 4586 3338 4592 3339
rect 4810 3343 4816 3344
rect 4810 3339 4811 3343
rect 4815 3339 4816 3343
rect 4810 3338 4816 3339
rect 5026 3343 5032 3344
rect 5026 3339 5027 3343
rect 5031 3339 5032 3343
rect 5026 3338 5032 3339
rect 5234 3343 5240 3344
rect 5234 3339 5235 3343
rect 5239 3339 5240 3343
rect 5234 3338 5240 3339
rect 5450 3343 5456 3344
rect 5450 3339 5451 3343
rect 5455 3339 5456 3343
rect 5662 3340 5663 3344
rect 5667 3340 5668 3344
rect 5662 3339 5668 3340
rect 5450 3338 5456 3339
rect 3886 3328 3892 3329
rect 3838 3327 3844 3328
rect 3838 3323 3839 3327
rect 3843 3323 3844 3327
rect 3886 3324 3887 3328
rect 3891 3324 3892 3328
rect 3886 3323 3892 3324
rect 4126 3328 4132 3329
rect 4126 3324 4127 3328
rect 4131 3324 4132 3328
rect 4126 3323 4132 3324
rect 4374 3328 4380 3329
rect 4374 3324 4375 3328
rect 4379 3324 4380 3328
rect 4374 3323 4380 3324
rect 4614 3328 4620 3329
rect 4614 3324 4615 3328
rect 4619 3324 4620 3328
rect 4614 3323 4620 3324
rect 4838 3328 4844 3329
rect 4838 3324 4839 3328
rect 4843 3324 4844 3328
rect 4838 3323 4844 3324
rect 5054 3328 5060 3329
rect 5054 3324 5055 3328
rect 5059 3324 5060 3328
rect 5054 3323 5060 3324
rect 5262 3328 5268 3329
rect 5262 3324 5263 3328
rect 5267 3324 5268 3328
rect 5262 3323 5268 3324
rect 5478 3328 5484 3329
rect 5478 3324 5479 3328
rect 5483 3324 5484 3328
rect 5478 3323 5484 3324
rect 5662 3327 5668 3328
rect 5662 3323 5663 3327
rect 5667 3323 5668 3327
rect 3838 3322 3844 3323
rect 5662 3322 5668 3323
rect 110 3320 116 3321
rect 1934 3320 1940 3321
rect 110 3316 111 3320
rect 115 3316 116 3320
rect 110 3315 116 3316
rect 322 3319 328 3320
rect 322 3315 323 3319
rect 327 3315 328 3319
rect 322 3314 328 3315
rect 458 3319 464 3320
rect 458 3315 459 3319
rect 463 3315 464 3319
rect 458 3314 464 3315
rect 594 3319 600 3320
rect 594 3315 595 3319
rect 599 3315 600 3319
rect 594 3314 600 3315
rect 730 3319 736 3320
rect 730 3315 731 3319
rect 735 3315 736 3319
rect 730 3314 736 3315
rect 866 3319 872 3320
rect 866 3315 867 3319
rect 871 3315 872 3319
rect 1934 3316 1935 3320
rect 1939 3316 1940 3320
rect 1934 3315 1940 3316
rect 866 3314 872 3315
rect 350 3304 356 3305
rect 110 3303 116 3304
rect 110 3299 111 3303
rect 115 3299 116 3303
rect 350 3300 351 3304
rect 355 3300 356 3304
rect 350 3299 356 3300
rect 486 3304 492 3305
rect 486 3300 487 3304
rect 491 3300 492 3304
rect 486 3299 492 3300
rect 622 3304 628 3305
rect 622 3300 623 3304
rect 627 3300 628 3304
rect 622 3299 628 3300
rect 758 3304 764 3305
rect 758 3300 759 3304
rect 763 3300 764 3304
rect 758 3299 764 3300
rect 894 3304 900 3305
rect 894 3300 895 3304
rect 899 3300 900 3304
rect 894 3299 900 3300
rect 1934 3303 1940 3304
rect 1934 3299 1935 3303
rect 1939 3299 1940 3303
rect 110 3298 116 3299
rect 1934 3298 1940 3299
rect 1974 3301 1980 3302
rect 3798 3301 3804 3302
rect 1974 3297 1975 3301
rect 1979 3297 1980 3301
rect 1974 3296 1980 3297
rect 2150 3300 2156 3301
rect 2150 3296 2151 3300
rect 2155 3296 2156 3300
rect 2150 3295 2156 3296
rect 2398 3300 2404 3301
rect 2398 3296 2399 3300
rect 2403 3296 2404 3300
rect 2398 3295 2404 3296
rect 2686 3300 2692 3301
rect 2686 3296 2687 3300
rect 2691 3296 2692 3300
rect 2686 3295 2692 3296
rect 3014 3300 3020 3301
rect 3014 3296 3015 3300
rect 3019 3296 3020 3300
rect 3014 3295 3020 3296
rect 3358 3300 3364 3301
rect 3358 3296 3359 3300
rect 3363 3296 3364 3300
rect 3358 3295 3364 3296
rect 3678 3300 3684 3301
rect 3678 3296 3679 3300
rect 3683 3296 3684 3300
rect 3798 3297 3799 3301
rect 3803 3297 3804 3301
rect 3798 3296 3804 3297
rect 3678 3295 3684 3296
rect 2122 3285 2128 3286
rect 1974 3284 1980 3285
rect 1974 3280 1975 3284
rect 1979 3280 1980 3284
rect 2122 3281 2123 3285
rect 2127 3281 2128 3285
rect 2122 3280 2128 3281
rect 2370 3285 2376 3286
rect 2370 3281 2371 3285
rect 2375 3281 2376 3285
rect 2370 3280 2376 3281
rect 2658 3285 2664 3286
rect 2658 3281 2659 3285
rect 2663 3281 2664 3285
rect 2658 3280 2664 3281
rect 2986 3285 2992 3286
rect 2986 3281 2987 3285
rect 2991 3281 2992 3285
rect 2986 3280 2992 3281
rect 3330 3285 3336 3286
rect 3330 3281 3331 3285
rect 3335 3281 3336 3285
rect 3330 3280 3336 3281
rect 3650 3285 3656 3286
rect 3650 3281 3651 3285
rect 3655 3281 3656 3285
rect 3650 3280 3656 3281
rect 3798 3284 3804 3285
rect 3798 3280 3799 3284
rect 3803 3280 3804 3284
rect 1974 3279 1980 3280
rect 3798 3279 3804 3280
rect 3838 3269 3844 3270
rect 5662 3269 5668 3270
rect 3838 3265 3839 3269
rect 3843 3265 3844 3269
rect 3838 3264 3844 3265
rect 3886 3268 3892 3269
rect 3886 3264 3887 3268
rect 3891 3264 3892 3268
rect 3886 3263 3892 3264
rect 4126 3268 4132 3269
rect 4126 3264 4127 3268
rect 4131 3264 4132 3268
rect 4126 3263 4132 3264
rect 4374 3268 4380 3269
rect 4374 3264 4375 3268
rect 4379 3264 4380 3268
rect 4374 3263 4380 3264
rect 4606 3268 4612 3269
rect 4606 3264 4607 3268
rect 4611 3264 4612 3268
rect 4606 3263 4612 3264
rect 4814 3268 4820 3269
rect 4814 3264 4815 3268
rect 4819 3264 4820 3268
rect 4814 3263 4820 3264
rect 5014 3268 5020 3269
rect 5014 3264 5015 3268
rect 5019 3264 5020 3268
rect 5014 3263 5020 3264
rect 5198 3268 5204 3269
rect 5198 3264 5199 3268
rect 5203 3264 5204 3268
rect 5198 3263 5204 3264
rect 5382 3268 5388 3269
rect 5382 3264 5383 3268
rect 5387 3264 5388 3268
rect 5382 3263 5388 3264
rect 5542 3268 5548 3269
rect 5542 3264 5543 3268
rect 5547 3264 5548 3268
rect 5662 3265 5663 3269
rect 5667 3265 5668 3269
rect 5662 3264 5668 3265
rect 5542 3263 5548 3264
rect 3858 3253 3864 3254
rect 3838 3252 3844 3253
rect 3838 3248 3839 3252
rect 3843 3248 3844 3252
rect 3858 3249 3859 3253
rect 3863 3249 3864 3253
rect 3858 3248 3864 3249
rect 4098 3253 4104 3254
rect 4098 3249 4099 3253
rect 4103 3249 4104 3253
rect 4098 3248 4104 3249
rect 4346 3253 4352 3254
rect 4346 3249 4347 3253
rect 4351 3249 4352 3253
rect 4346 3248 4352 3249
rect 4578 3253 4584 3254
rect 4578 3249 4579 3253
rect 4583 3249 4584 3253
rect 4578 3248 4584 3249
rect 4786 3253 4792 3254
rect 4786 3249 4787 3253
rect 4791 3249 4792 3253
rect 4786 3248 4792 3249
rect 4986 3253 4992 3254
rect 4986 3249 4987 3253
rect 4991 3249 4992 3253
rect 4986 3248 4992 3249
rect 5170 3253 5176 3254
rect 5170 3249 5171 3253
rect 5175 3249 5176 3253
rect 5170 3248 5176 3249
rect 5354 3253 5360 3254
rect 5354 3249 5355 3253
rect 5359 3249 5360 3253
rect 5354 3248 5360 3249
rect 5514 3253 5520 3254
rect 5514 3249 5515 3253
rect 5519 3249 5520 3253
rect 5514 3248 5520 3249
rect 5662 3252 5668 3253
rect 5662 3248 5663 3252
rect 5667 3248 5668 3252
rect 3838 3247 3844 3248
rect 5662 3247 5668 3248
rect 110 3237 116 3238
rect 1934 3237 1940 3238
rect 110 3233 111 3237
rect 115 3233 116 3237
rect 110 3232 116 3233
rect 158 3236 164 3237
rect 158 3232 159 3236
rect 163 3232 164 3236
rect 158 3231 164 3232
rect 334 3236 340 3237
rect 334 3232 335 3236
rect 339 3232 340 3236
rect 334 3231 340 3232
rect 542 3236 548 3237
rect 542 3232 543 3236
rect 547 3232 548 3236
rect 542 3231 548 3232
rect 750 3236 756 3237
rect 750 3232 751 3236
rect 755 3232 756 3236
rect 750 3231 756 3232
rect 958 3236 964 3237
rect 958 3232 959 3236
rect 963 3232 964 3236
rect 1934 3233 1935 3237
rect 1939 3233 1940 3237
rect 1934 3232 1940 3233
rect 958 3231 964 3232
rect 130 3221 136 3222
rect 110 3220 116 3221
rect 110 3216 111 3220
rect 115 3216 116 3220
rect 130 3217 131 3221
rect 135 3217 136 3221
rect 130 3216 136 3217
rect 306 3221 312 3222
rect 306 3217 307 3221
rect 311 3217 312 3221
rect 306 3216 312 3217
rect 514 3221 520 3222
rect 514 3217 515 3221
rect 519 3217 520 3221
rect 514 3216 520 3217
rect 722 3221 728 3222
rect 722 3217 723 3221
rect 727 3217 728 3221
rect 722 3216 728 3217
rect 930 3221 936 3222
rect 930 3217 931 3221
rect 935 3217 936 3221
rect 930 3216 936 3217
rect 1934 3220 1940 3221
rect 1934 3216 1935 3220
rect 1939 3216 1940 3220
rect 110 3215 116 3216
rect 1934 3215 1940 3216
rect 1974 3152 1980 3153
rect 3798 3152 3804 3153
rect 1974 3148 1975 3152
rect 1979 3148 1980 3152
rect 1974 3147 1980 3148
rect 1994 3151 2000 3152
rect 1994 3147 1995 3151
rect 1999 3147 2000 3151
rect 1994 3146 2000 3147
rect 2146 3151 2152 3152
rect 2146 3147 2147 3151
rect 2151 3147 2152 3151
rect 2146 3146 2152 3147
rect 2346 3151 2352 3152
rect 2346 3147 2347 3151
rect 2351 3147 2352 3151
rect 2346 3146 2352 3147
rect 2554 3151 2560 3152
rect 2554 3147 2555 3151
rect 2559 3147 2560 3151
rect 2554 3146 2560 3147
rect 2770 3151 2776 3152
rect 2770 3147 2771 3151
rect 2775 3147 2776 3151
rect 2770 3146 2776 3147
rect 2986 3151 2992 3152
rect 2986 3147 2987 3151
rect 2991 3147 2992 3151
rect 2986 3146 2992 3147
rect 3210 3151 3216 3152
rect 3210 3147 3211 3151
rect 3215 3147 3216 3151
rect 3210 3146 3216 3147
rect 3442 3151 3448 3152
rect 3442 3147 3443 3151
rect 3447 3147 3448 3151
rect 3442 3146 3448 3147
rect 3650 3151 3656 3152
rect 3650 3147 3651 3151
rect 3655 3147 3656 3151
rect 3798 3148 3799 3152
rect 3803 3148 3804 3152
rect 3798 3147 3804 3148
rect 3650 3146 3656 3147
rect 2022 3136 2028 3137
rect 1974 3135 1980 3136
rect 1974 3131 1975 3135
rect 1979 3131 1980 3135
rect 2022 3132 2023 3136
rect 2027 3132 2028 3136
rect 2022 3131 2028 3132
rect 2174 3136 2180 3137
rect 2174 3132 2175 3136
rect 2179 3132 2180 3136
rect 2174 3131 2180 3132
rect 2374 3136 2380 3137
rect 2374 3132 2375 3136
rect 2379 3132 2380 3136
rect 2374 3131 2380 3132
rect 2582 3136 2588 3137
rect 2582 3132 2583 3136
rect 2587 3132 2588 3136
rect 2582 3131 2588 3132
rect 2798 3136 2804 3137
rect 2798 3132 2799 3136
rect 2803 3132 2804 3136
rect 2798 3131 2804 3132
rect 3014 3136 3020 3137
rect 3014 3132 3015 3136
rect 3019 3132 3020 3136
rect 3014 3131 3020 3132
rect 3238 3136 3244 3137
rect 3238 3132 3239 3136
rect 3243 3132 3244 3136
rect 3238 3131 3244 3132
rect 3470 3136 3476 3137
rect 3470 3132 3471 3136
rect 3475 3132 3476 3136
rect 3470 3131 3476 3132
rect 3678 3136 3684 3137
rect 3678 3132 3679 3136
rect 3683 3132 3684 3136
rect 3678 3131 3684 3132
rect 3798 3135 3804 3136
rect 3798 3131 3799 3135
rect 3803 3131 3804 3135
rect 1974 3130 1980 3131
rect 3798 3130 3804 3131
rect 3838 3104 3844 3105
rect 5662 3104 5668 3105
rect 3838 3100 3839 3104
rect 3843 3100 3844 3104
rect 3838 3099 3844 3100
rect 4466 3103 4472 3104
rect 4466 3099 4467 3103
rect 4471 3099 4472 3103
rect 4466 3098 4472 3099
rect 4650 3103 4656 3104
rect 4650 3099 4651 3103
rect 4655 3099 4656 3103
rect 4650 3098 4656 3099
rect 4858 3103 4864 3104
rect 4858 3099 4859 3103
rect 4863 3099 4864 3103
rect 4858 3098 4864 3099
rect 5074 3103 5080 3104
rect 5074 3099 5075 3103
rect 5079 3099 5080 3103
rect 5074 3098 5080 3099
rect 5306 3103 5312 3104
rect 5306 3099 5307 3103
rect 5311 3099 5312 3103
rect 5306 3098 5312 3099
rect 5514 3103 5520 3104
rect 5514 3099 5515 3103
rect 5519 3099 5520 3103
rect 5662 3100 5663 3104
rect 5667 3100 5668 3104
rect 5662 3099 5668 3100
rect 5514 3098 5520 3099
rect 4494 3088 4500 3089
rect 3838 3087 3844 3088
rect 3838 3083 3839 3087
rect 3843 3083 3844 3087
rect 4494 3084 4495 3088
rect 4499 3084 4500 3088
rect 4494 3083 4500 3084
rect 4678 3088 4684 3089
rect 4678 3084 4679 3088
rect 4683 3084 4684 3088
rect 4678 3083 4684 3084
rect 4886 3088 4892 3089
rect 4886 3084 4887 3088
rect 4891 3084 4892 3088
rect 4886 3083 4892 3084
rect 5102 3088 5108 3089
rect 5102 3084 5103 3088
rect 5107 3084 5108 3088
rect 5102 3083 5108 3084
rect 5334 3088 5340 3089
rect 5334 3084 5335 3088
rect 5339 3084 5340 3088
rect 5334 3083 5340 3084
rect 5542 3088 5548 3089
rect 5542 3084 5543 3088
rect 5547 3084 5548 3088
rect 5542 3083 5548 3084
rect 5662 3087 5668 3088
rect 5662 3083 5663 3087
rect 5667 3083 5668 3087
rect 3838 3082 3844 3083
rect 5662 3082 5668 3083
rect 1974 3077 1980 3078
rect 3798 3077 3804 3078
rect 1974 3073 1975 3077
rect 1979 3073 1980 3077
rect 110 3072 116 3073
rect 1934 3072 1940 3073
rect 1974 3072 1980 3073
rect 2646 3076 2652 3077
rect 2646 3072 2647 3076
rect 2651 3072 2652 3076
rect 110 3068 111 3072
rect 115 3068 116 3072
rect 110 3067 116 3068
rect 130 3071 136 3072
rect 130 3067 131 3071
rect 135 3067 136 3071
rect 130 3066 136 3067
rect 370 3071 376 3072
rect 370 3067 371 3071
rect 375 3067 376 3071
rect 370 3066 376 3067
rect 626 3071 632 3072
rect 626 3067 627 3071
rect 631 3067 632 3071
rect 626 3066 632 3067
rect 874 3071 880 3072
rect 874 3067 875 3071
rect 879 3067 880 3071
rect 874 3066 880 3067
rect 1114 3071 1120 3072
rect 1114 3067 1115 3071
rect 1119 3067 1120 3071
rect 1114 3066 1120 3067
rect 1346 3071 1352 3072
rect 1346 3067 1347 3071
rect 1351 3067 1352 3071
rect 1346 3066 1352 3067
rect 1578 3071 1584 3072
rect 1578 3067 1579 3071
rect 1583 3067 1584 3071
rect 1578 3066 1584 3067
rect 1786 3071 1792 3072
rect 1786 3067 1787 3071
rect 1791 3067 1792 3071
rect 1934 3068 1935 3072
rect 1939 3068 1940 3072
rect 2646 3071 2652 3072
rect 2782 3076 2788 3077
rect 2782 3072 2783 3076
rect 2787 3072 2788 3076
rect 2782 3071 2788 3072
rect 2926 3076 2932 3077
rect 2926 3072 2927 3076
rect 2931 3072 2932 3076
rect 2926 3071 2932 3072
rect 3078 3076 3084 3077
rect 3078 3072 3079 3076
rect 3083 3072 3084 3076
rect 3078 3071 3084 3072
rect 3238 3076 3244 3077
rect 3238 3072 3239 3076
rect 3243 3072 3244 3076
rect 3238 3071 3244 3072
rect 3398 3076 3404 3077
rect 3398 3072 3399 3076
rect 3403 3072 3404 3076
rect 3398 3071 3404 3072
rect 3566 3076 3572 3077
rect 3566 3072 3567 3076
rect 3571 3072 3572 3076
rect 3798 3073 3799 3077
rect 3803 3073 3804 3077
rect 3798 3072 3804 3073
rect 3566 3071 3572 3072
rect 1934 3067 1940 3068
rect 1786 3066 1792 3067
rect 2618 3061 2624 3062
rect 1974 3060 1980 3061
rect 158 3056 164 3057
rect 110 3055 116 3056
rect 110 3051 111 3055
rect 115 3051 116 3055
rect 158 3052 159 3056
rect 163 3052 164 3056
rect 158 3051 164 3052
rect 398 3056 404 3057
rect 398 3052 399 3056
rect 403 3052 404 3056
rect 398 3051 404 3052
rect 654 3056 660 3057
rect 654 3052 655 3056
rect 659 3052 660 3056
rect 654 3051 660 3052
rect 902 3056 908 3057
rect 902 3052 903 3056
rect 907 3052 908 3056
rect 902 3051 908 3052
rect 1142 3056 1148 3057
rect 1142 3052 1143 3056
rect 1147 3052 1148 3056
rect 1142 3051 1148 3052
rect 1374 3056 1380 3057
rect 1374 3052 1375 3056
rect 1379 3052 1380 3056
rect 1374 3051 1380 3052
rect 1606 3056 1612 3057
rect 1606 3052 1607 3056
rect 1611 3052 1612 3056
rect 1606 3051 1612 3052
rect 1814 3056 1820 3057
rect 1974 3056 1975 3060
rect 1979 3056 1980 3060
rect 2618 3057 2619 3061
rect 2623 3057 2624 3061
rect 2618 3056 2624 3057
rect 2754 3061 2760 3062
rect 2754 3057 2755 3061
rect 2759 3057 2760 3061
rect 2754 3056 2760 3057
rect 2898 3061 2904 3062
rect 2898 3057 2899 3061
rect 2903 3057 2904 3061
rect 2898 3056 2904 3057
rect 3050 3061 3056 3062
rect 3050 3057 3051 3061
rect 3055 3057 3056 3061
rect 3050 3056 3056 3057
rect 3210 3061 3216 3062
rect 3210 3057 3211 3061
rect 3215 3057 3216 3061
rect 3210 3056 3216 3057
rect 3370 3061 3376 3062
rect 3370 3057 3371 3061
rect 3375 3057 3376 3061
rect 3370 3056 3376 3057
rect 3538 3061 3544 3062
rect 3538 3057 3539 3061
rect 3543 3057 3544 3061
rect 3538 3056 3544 3057
rect 3798 3060 3804 3061
rect 3798 3056 3799 3060
rect 3803 3056 3804 3060
rect 1814 3052 1815 3056
rect 1819 3052 1820 3056
rect 1814 3051 1820 3052
rect 1934 3055 1940 3056
rect 1974 3055 1980 3056
rect 3798 3055 3804 3056
rect 1934 3051 1935 3055
rect 1939 3051 1940 3055
rect 110 3050 116 3051
rect 1934 3050 1940 3051
rect 3838 3029 3844 3030
rect 5662 3029 5668 3030
rect 3838 3025 3839 3029
rect 3843 3025 3844 3029
rect 3838 3024 3844 3025
rect 4254 3028 4260 3029
rect 4254 3024 4255 3028
rect 4259 3024 4260 3028
rect 4254 3023 4260 3024
rect 4454 3028 4460 3029
rect 4454 3024 4455 3028
rect 4459 3024 4460 3028
rect 4454 3023 4460 3024
rect 4670 3028 4676 3029
rect 4670 3024 4671 3028
rect 4675 3024 4676 3028
rect 4670 3023 4676 3024
rect 4910 3028 4916 3029
rect 4910 3024 4911 3028
rect 4915 3024 4916 3028
rect 4910 3023 4916 3024
rect 5166 3028 5172 3029
rect 5166 3024 5167 3028
rect 5171 3024 5172 3028
rect 5166 3023 5172 3024
rect 5422 3028 5428 3029
rect 5422 3024 5423 3028
rect 5427 3024 5428 3028
rect 5662 3025 5663 3029
rect 5667 3025 5668 3029
rect 5662 3024 5668 3025
rect 5422 3023 5428 3024
rect 4226 3013 4232 3014
rect 3838 3012 3844 3013
rect 3838 3008 3839 3012
rect 3843 3008 3844 3012
rect 4226 3009 4227 3013
rect 4231 3009 4232 3013
rect 4226 3008 4232 3009
rect 4426 3013 4432 3014
rect 4426 3009 4427 3013
rect 4431 3009 4432 3013
rect 4426 3008 4432 3009
rect 4642 3013 4648 3014
rect 4642 3009 4643 3013
rect 4647 3009 4648 3013
rect 4642 3008 4648 3009
rect 4882 3013 4888 3014
rect 4882 3009 4883 3013
rect 4887 3009 4888 3013
rect 4882 3008 4888 3009
rect 5138 3013 5144 3014
rect 5138 3009 5139 3013
rect 5143 3009 5144 3013
rect 5138 3008 5144 3009
rect 5394 3013 5400 3014
rect 5394 3009 5395 3013
rect 5399 3009 5400 3013
rect 5394 3008 5400 3009
rect 5662 3012 5668 3013
rect 5662 3008 5663 3012
rect 5667 3008 5668 3012
rect 3838 3007 3844 3008
rect 5662 3007 5668 3008
rect 110 2997 116 2998
rect 1934 2997 1940 2998
rect 110 2993 111 2997
rect 115 2993 116 2997
rect 110 2992 116 2993
rect 174 2996 180 2997
rect 174 2992 175 2996
rect 179 2992 180 2996
rect 174 2991 180 2992
rect 406 2996 412 2997
rect 406 2992 407 2996
rect 411 2992 412 2996
rect 406 2991 412 2992
rect 622 2996 628 2997
rect 622 2992 623 2996
rect 627 2992 628 2996
rect 622 2991 628 2992
rect 822 2996 828 2997
rect 822 2992 823 2996
rect 827 2992 828 2996
rect 822 2991 828 2992
rect 1006 2996 1012 2997
rect 1006 2992 1007 2996
rect 1011 2992 1012 2996
rect 1006 2991 1012 2992
rect 1182 2996 1188 2997
rect 1182 2992 1183 2996
rect 1187 2992 1188 2996
rect 1182 2991 1188 2992
rect 1350 2996 1356 2997
rect 1350 2992 1351 2996
rect 1355 2992 1356 2996
rect 1350 2991 1356 2992
rect 1510 2996 1516 2997
rect 1510 2992 1511 2996
rect 1515 2992 1516 2996
rect 1510 2991 1516 2992
rect 1670 2996 1676 2997
rect 1670 2992 1671 2996
rect 1675 2992 1676 2996
rect 1670 2991 1676 2992
rect 1814 2996 1820 2997
rect 1814 2992 1815 2996
rect 1819 2992 1820 2996
rect 1934 2993 1935 2997
rect 1939 2993 1940 2997
rect 1934 2992 1940 2993
rect 1814 2991 1820 2992
rect 146 2981 152 2982
rect 110 2980 116 2981
rect 110 2976 111 2980
rect 115 2976 116 2980
rect 146 2977 147 2981
rect 151 2977 152 2981
rect 146 2976 152 2977
rect 378 2981 384 2982
rect 378 2977 379 2981
rect 383 2977 384 2981
rect 378 2976 384 2977
rect 594 2981 600 2982
rect 594 2977 595 2981
rect 599 2977 600 2981
rect 594 2976 600 2977
rect 794 2981 800 2982
rect 794 2977 795 2981
rect 799 2977 800 2981
rect 794 2976 800 2977
rect 978 2981 984 2982
rect 978 2977 979 2981
rect 983 2977 984 2981
rect 978 2976 984 2977
rect 1154 2981 1160 2982
rect 1154 2977 1155 2981
rect 1159 2977 1160 2981
rect 1154 2976 1160 2977
rect 1322 2981 1328 2982
rect 1322 2977 1323 2981
rect 1327 2977 1328 2981
rect 1322 2976 1328 2977
rect 1482 2981 1488 2982
rect 1482 2977 1483 2981
rect 1487 2977 1488 2981
rect 1482 2976 1488 2977
rect 1642 2981 1648 2982
rect 1642 2977 1643 2981
rect 1647 2977 1648 2981
rect 1642 2976 1648 2977
rect 1786 2981 1792 2982
rect 1786 2977 1787 2981
rect 1791 2977 1792 2981
rect 1786 2976 1792 2977
rect 1934 2980 1940 2981
rect 1934 2976 1935 2980
rect 1939 2976 1940 2980
rect 110 2975 116 2976
rect 1934 2975 1940 2976
rect 1974 2928 1980 2929
rect 3798 2928 3804 2929
rect 1974 2924 1975 2928
rect 1979 2924 1980 2928
rect 1974 2923 1980 2924
rect 2802 2927 2808 2928
rect 2802 2923 2803 2927
rect 2807 2923 2808 2927
rect 2802 2922 2808 2923
rect 2938 2927 2944 2928
rect 2938 2923 2939 2927
rect 2943 2923 2944 2927
rect 2938 2922 2944 2923
rect 3074 2927 3080 2928
rect 3074 2923 3075 2927
rect 3079 2923 3080 2927
rect 3074 2922 3080 2923
rect 3210 2927 3216 2928
rect 3210 2923 3211 2927
rect 3215 2923 3216 2927
rect 3210 2922 3216 2923
rect 3346 2927 3352 2928
rect 3346 2923 3347 2927
rect 3351 2923 3352 2927
rect 3346 2922 3352 2923
rect 3482 2927 3488 2928
rect 3482 2923 3483 2927
rect 3487 2923 3488 2927
rect 3798 2924 3799 2928
rect 3803 2924 3804 2928
rect 3798 2923 3804 2924
rect 3482 2922 3488 2923
rect 2830 2912 2836 2913
rect 1974 2911 1980 2912
rect 1974 2907 1975 2911
rect 1979 2907 1980 2911
rect 2830 2908 2831 2912
rect 2835 2908 2836 2912
rect 2830 2907 2836 2908
rect 2966 2912 2972 2913
rect 2966 2908 2967 2912
rect 2971 2908 2972 2912
rect 2966 2907 2972 2908
rect 3102 2912 3108 2913
rect 3102 2908 3103 2912
rect 3107 2908 3108 2912
rect 3102 2907 3108 2908
rect 3238 2912 3244 2913
rect 3238 2908 3239 2912
rect 3243 2908 3244 2912
rect 3238 2907 3244 2908
rect 3374 2912 3380 2913
rect 3374 2908 3375 2912
rect 3379 2908 3380 2912
rect 3374 2907 3380 2908
rect 3510 2912 3516 2913
rect 3510 2908 3511 2912
rect 3515 2908 3516 2912
rect 3510 2907 3516 2908
rect 3798 2911 3804 2912
rect 3798 2907 3799 2911
rect 3803 2907 3804 2911
rect 1974 2906 1980 2907
rect 3798 2906 3804 2907
rect 3838 2856 3844 2857
rect 5662 2856 5668 2857
rect 3838 2852 3839 2856
rect 3843 2852 3844 2856
rect 3838 2851 3844 2852
rect 3994 2855 4000 2856
rect 3994 2851 3995 2855
rect 3999 2851 4000 2855
rect 3994 2850 4000 2851
rect 4210 2855 4216 2856
rect 4210 2851 4211 2855
rect 4215 2851 4216 2855
rect 4210 2850 4216 2851
rect 4442 2855 4448 2856
rect 4442 2851 4443 2855
rect 4447 2851 4448 2855
rect 4442 2850 4448 2851
rect 4698 2855 4704 2856
rect 4698 2851 4699 2855
rect 4703 2851 4704 2855
rect 4698 2850 4704 2851
rect 4970 2855 4976 2856
rect 4970 2851 4971 2855
rect 4975 2851 4976 2855
rect 4970 2850 4976 2851
rect 5250 2855 5256 2856
rect 5250 2851 5251 2855
rect 5255 2851 5256 2855
rect 5250 2850 5256 2851
rect 5514 2855 5520 2856
rect 5514 2851 5515 2855
rect 5519 2851 5520 2855
rect 5662 2852 5663 2856
rect 5667 2852 5668 2856
rect 5662 2851 5668 2852
rect 5514 2850 5520 2851
rect 110 2844 116 2845
rect 1934 2844 1940 2845
rect 110 2840 111 2844
rect 115 2840 116 2844
rect 110 2839 116 2840
rect 394 2843 400 2844
rect 394 2839 395 2843
rect 399 2839 400 2843
rect 394 2838 400 2839
rect 594 2843 600 2844
rect 594 2839 595 2843
rect 599 2839 600 2843
rect 594 2838 600 2839
rect 786 2843 792 2844
rect 786 2839 787 2843
rect 791 2839 792 2843
rect 786 2838 792 2839
rect 970 2843 976 2844
rect 970 2839 971 2843
rect 975 2839 976 2843
rect 970 2838 976 2839
rect 1146 2843 1152 2844
rect 1146 2839 1147 2843
rect 1151 2839 1152 2843
rect 1146 2838 1152 2839
rect 1314 2843 1320 2844
rect 1314 2839 1315 2843
rect 1319 2839 1320 2843
rect 1314 2838 1320 2839
rect 1482 2843 1488 2844
rect 1482 2839 1483 2843
rect 1487 2839 1488 2843
rect 1482 2838 1488 2839
rect 1642 2843 1648 2844
rect 1642 2839 1643 2843
rect 1647 2839 1648 2843
rect 1642 2838 1648 2839
rect 1786 2843 1792 2844
rect 1786 2839 1787 2843
rect 1791 2839 1792 2843
rect 1934 2840 1935 2844
rect 1939 2840 1940 2844
rect 4022 2840 4028 2841
rect 1934 2839 1940 2840
rect 3838 2839 3844 2840
rect 1786 2838 1792 2839
rect 3838 2835 3839 2839
rect 3843 2835 3844 2839
rect 4022 2836 4023 2840
rect 4027 2836 4028 2840
rect 4022 2835 4028 2836
rect 4238 2840 4244 2841
rect 4238 2836 4239 2840
rect 4243 2836 4244 2840
rect 4238 2835 4244 2836
rect 4470 2840 4476 2841
rect 4470 2836 4471 2840
rect 4475 2836 4476 2840
rect 4470 2835 4476 2836
rect 4726 2840 4732 2841
rect 4726 2836 4727 2840
rect 4731 2836 4732 2840
rect 4726 2835 4732 2836
rect 4998 2840 5004 2841
rect 4998 2836 4999 2840
rect 5003 2836 5004 2840
rect 4998 2835 5004 2836
rect 5278 2840 5284 2841
rect 5278 2836 5279 2840
rect 5283 2836 5284 2840
rect 5278 2835 5284 2836
rect 5542 2840 5548 2841
rect 5542 2836 5543 2840
rect 5547 2836 5548 2840
rect 5542 2835 5548 2836
rect 5662 2839 5668 2840
rect 5662 2835 5663 2839
rect 5667 2835 5668 2839
rect 3838 2834 3844 2835
rect 5662 2834 5668 2835
rect 422 2828 428 2829
rect 110 2827 116 2828
rect 110 2823 111 2827
rect 115 2823 116 2827
rect 422 2824 423 2828
rect 427 2824 428 2828
rect 422 2823 428 2824
rect 622 2828 628 2829
rect 622 2824 623 2828
rect 627 2824 628 2828
rect 622 2823 628 2824
rect 814 2828 820 2829
rect 814 2824 815 2828
rect 819 2824 820 2828
rect 814 2823 820 2824
rect 998 2828 1004 2829
rect 998 2824 999 2828
rect 1003 2824 1004 2828
rect 998 2823 1004 2824
rect 1174 2828 1180 2829
rect 1174 2824 1175 2828
rect 1179 2824 1180 2828
rect 1174 2823 1180 2824
rect 1342 2828 1348 2829
rect 1342 2824 1343 2828
rect 1347 2824 1348 2828
rect 1342 2823 1348 2824
rect 1510 2828 1516 2829
rect 1510 2824 1511 2828
rect 1515 2824 1516 2828
rect 1510 2823 1516 2824
rect 1670 2828 1676 2829
rect 1670 2824 1671 2828
rect 1675 2824 1676 2828
rect 1670 2823 1676 2824
rect 1814 2828 1820 2829
rect 1814 2824 1815 2828
rect 1819 2824 1820 2828
rect 1814 2823 1820 2824
rect 1934 2827 1940 2828
rect 1934 2823 1935 2827
rect 1939 2823 1940 2827
rect 110 2822 116 2823
rect 1934 2822 1940 2823
rect 1974 2801 1980 2802
rect 3798 2801 3804 2802
rect 1974 2797 1975 2801
rect 1979 2797 1980 2801
rect 1974 2796 1980 2797
rect 2022 2800 2028 2801
rect 2022 2796 2023 2800
rect 2027 2796 2028 2800
rect 2022 2795 2028 2796
rect 2166 2800 2172 2801
rect 2166 2796 2167 2800
rect 2171 2796 2172 2800
rect 2166 2795 2172 2796
rect 2334 2800 2340 2801
rect 2334 2796 2335 2800
rect 2339 2796 2340 2800
rect 2334 2795 2340 2796
rect 2494 2800 2500 2801
rect 2494 2796 2495 2800
rect 2499 2796 2500 2800
rect 2494 2795 2500 2796
rect 2662 2800 2668 2801
rect 2662 2796 2663 2800
rect 2667 2796 2668 2800
rect 2662 2795 2668 2796
rect 2830 2800 2836 2801
rect 2830 2796 2831 2800
rect 2835 2796 2836 2800
rect 2830 2795 2836 2796
rect 2998 2800 3004 2801
rect 2998 2796 2999 2800
rect 3003 2796 3004 2800
rect 2998 2795 3004 2796
rect 3166 2800 3172 2801
rect 3166 2796 3167 2800
rect 3171 2796 3172 2800
rect 3798 2797 3799 2801
rect 3803 2797 3804 2801
rect 3798 2796 3804 2797
rect 3166 2795 3172 2796
rect 1994 2785 2000 2786
rect 1974 2784 1980 2785
rect 1974 2780 1975 2784
rect 1979 2780 1980 2784
rect 1994 2781 1995 2785
rect 1999 2781 2000 2785
rect 1994 2780 2000 2781
rect 2138 2785 2144 2786
rect 2138 2781 2139 2785
rect 2143 2781 2144 2785
rect 2138 2780 2144 2781
rect 2306 2785 2312 2786
rect 2306 2781 2307 2785
rect 2311 2781 2312 2785
rect 2306 2780 2312 2781
rect 2466 2785 2472 2786
rect 2466 2781 2467 2785
rect 2471 2781 2472 2785
rect 2466 2780 2472 2781
rect 2634 2785 2640 2786
rect 2634 2781 2635 2785
rect 2639 2781 2640 2785
rect 2634 2780 2640 2781
rect 2802 2785 2808 2786
rect 2802 2781 2803 2785
rect 2807 2781 2808 2785
rect 2802 2780 2808 2781
rect 2970 2785 2976 2786
rect 2970 2781 2971 2785
rect 2975 2781 2976 2785
rect 2970 2780 2976 2781
rect 3138 2785 3144 2786
rect 3138 2781 3139 2785
rect 3143 2781 3144 2785
rect 3138 2780 3144 2781
rect 3798 2784 3804 2785
rect 3798 2780 3799 2784
rect 3803 2780 3804 2784
rect 1974 2779 1980 2780
rect 3798 2779 3804 2780
rect 3838 2777 3844 2778
rect 5662 2777 5668 2778
rect 3838 2773 3839 2777
rect 3843 2773 3844 2777
rect 3838 2772 3844 2773
rect 3918 2776 3924 2777
rect 3918 2772 3919 2776
rect 3923 2772 3924 2776
rect 3918 2771 3924 2772
rect 4054 2776 4060 2777
rect 4054 2772 4055 2776
rect 4059 2772 4060 2776
rect 4054 2771 4060 2772
rect 4190 2776 4196 2777
rect 4190 2772 4191 2776
rect 4195 2772 4196 2776
rect 4190 2771 4196 2772
rect 4326 2776 4332 2777
rect 4326 2772 4327 2776
rect 4331 2772 4332 2776
rect 4326 2771 4332 2772
rect 4462 2776 4468 2777
rect 4462 2772 4463 2776
rect 4467 2772 4468 2776
rect 5662 2773 5663 2777
rect 5667 2773 5668 2777
rect 5662 2772 5668 2773
rect 4462 2771 4468 2772
rect 3890 2761 3896 2762
rect 3838 2760 3844 2761
rect 110 2757 116 2758
rect 1934 2757 1940 2758
rect 110 2753 111 2757
rect 115 2753 116 2757
rect 110 2752 116 2753
rect 654 2756 660 2757
rect 654 2752 655 2756
rect 659 2752 660 2756
rect 654 2751 660 2752
rect 814 2756 820 2757
rect 814 2752 815 2756
rect 819 2752 820 2756
rect 814 2751 820 2752
rect 974 2756 980 2757
rect 974 2752 975 2756
rect 979 2752 980 2756
rect 974 2751 980 2752
rect 1142 2756 1148 2757
rect 1142 2752 1143 2756
rect 1147 2752 1148 2756
rect 1142 2751 1148 2752
rect 1310 2756 1316 2757
rect 1310 2752 1311 2756
rect 1315 2752 1316 2756
rect 1310 2751 1316 2752
rect 1478 2756 1484 2757
rect 1478 2752 1479 2756
rect 1483 2752 1484 2756
rect 1934 2753 1935 2757
rect 1939 2753 1940 2757
rect 3838 2756 3839 2760
rect 3843 2756 3844 2760
rect 3890 2757 3891 2761
rect 3895 2757 3896 2761
rect 3890 2756 3896 2757
rect 4026 2761 4032 2762
rect 4026 2757 4027 2761
rect 4031 2757 4032 2761
rect 4026 2756 4032 2757
rect 4162 2761 4168 2762
rect 4162 2757 4163 2761
rect 4167 2757 4168 2761
rect 4162 2756 4168 2757
rect 4298 2761 4304 2762
rect 4298 2757 4299 2761
rect 4303 2757 4304 2761
rect 4298 2756 4304 2757
rect 4434 2761 4440 2762
rect 4434 2757 4435 2761
rect 4439 2757 4440 2761
rect 4434 2756 4440 2757
rect 5662 2760 5668 2761
rect 5662 2756 5663 2760
rect 5667 2756 5668 2760
rect 3838 2755 3844 2756
rect 5662 2755 5668 2756
rect 1934 2752 1940 2753
rect 1478 2751 1484 2752
rect 626 2741 632 2742
rect 110 2740 116 2741
rect 110 2736 111 2740
rect 115 2736 116 2740
rect 626 2737 627 2741
rect 631 2737 632 2741
rect 626 2736 632 2737
rect 786 2741 792 2742
rect 786 2737 787 2741
rect 791 2737 792 2741
rect 786 2736 792 2737
rect 946 2741 952 2742
rect 946 2737 947 2741
rect 951 2737 952 2741
rect 946 2736 952 2737
rect 1114 2741 1120 2742
rect 1114 2737 1115 2741
rect 1119 2737 1120 2741
rect 1114 2736 1120 2737
rect 1282 2741 1288 2742
rect 1282 2737 1283 2741
rect 1287 2737 1288 2741
rect 1282 2736 1288 2737
rect 1450 2741 1456 2742
rect 1450 2737 1451 2741
rect 1455 2737 1456 2741
rect 1450 2736 1456 2737
rect 1934 2740 1940 2741
rect 1934 2736 1935 2740
rect 1939 2736 1940 2740
rect 110 2735 116 2736
rect 1934 2735 1940 2736
rect 1974 2652 1980 2653
rect 3798 2652 3804 2653
rect 1974 2648 1975 2652
rect 1979 2648 1980 2652
rect 1974 2647 1980 2648
rect 2378 2651 2384 2652
rect 2378 2647 2379 2651
rect 2383 2647 2384 2651
rect 2378 2646 2384 2647
rect 2514 2651 2520 2652
rect 2514 2647 2515 2651
rect 2519 2647 2520 2651
rect 2514 2646 2520 2647
rect 2658 2651 2664 2652
rect 2658 2647 2659 2651
rect 2663 2647 2664 2651
rect 2658 2646 2664 2647
rect 2802 2651 2808 2652
rect 2802 2647 2803 2651
rect 2807 2647 2808 2651
rect 2802 2646 2808 2647
rect 2946 2651 2952 2652
rect 2946 2647 2947 2651
rect 2951 2647 2952 2651
rect 2946 2646 2952 2647
rect 3090 2651 3096 2652
rect 3090 2647 3091 2651
rect 3095 2647 3096 2651
rect 3090 2646 3096 2647
rect 3234 2651 3240 2652
rect 3234 2647 3235 2651
rect 3239 2647 3240 2651
rect 3798 2648 3799 2652
rect 3803 2648 3804 2652
rect 3798 2647 3804 2648
rect 3234 2646 3240 2647
rect 2406 2636 2412 2637
rect 1974 2635 1980 2636
rect 1974 2631 1975 2635
rect 1979 2631 1980 2635
rect 2406 2632 2407 2636
rect 2411 2632 2412 2636
rect 2406 2631 2412 2632
rect 2542 2636 2548 2637
rect 2542 2632 2543 2636
rect 2547 2632 2548 2636
rect 2542 2631 2548 2632
rect 2686 2636 2692 2637
rect 2686 2632 2687 2636
rect 2691 2632 2692 2636
rect 2686 2631 2692 2632
rect 2830 2636 2836 2637
rect 2830 2632 2831 2636
rect 2835 2632 2836 2636
rect 2830 2631 2836 2632
rect 2974 2636 2980 2637
rect 2974 2632 2975 2636
rect 2979 2632 2980 2636
rect 2974 2631 2980 2632
rect 3118 2636 3124 2637
rect 3118 2632 3119 2636
rect 3123 2632 3124 2636
rect 3118 2631 3124 2632
rect 3262 2636 3268 2637
rect 3262 2632 3263 2636
rect 3267 2632 3268 2636
rect 3262 2631 3268 2632
rect 3798 2635 3804 2636
rect 3798 2631 3799 2635
rect 3803 2631 3804 2635
rect 1974 2630 1980 2631
rect 3798 2630 3804 2631
rect 3838 2616 3844 2617
rect 5662 2616 5668 2617
rect 3838 2612 3839 2616
rect 3843 2612 3844 2616
rect 3838 2611 3844 2612
rect 4098 2615 4104 2616
rect 4098 2611 4099 2615
rect 4103 2611 4104 2615
rect 4098 2610 4104 2611
rect 4298 2615 4304 2616
rect 4298 2611 4299 2615
rect 4303 2611 4304 2615
rect 4298 2610 4304 2611
rect 4514 2615 4520 2616
rect 4514 2611 4515 2615
rect 4519 2611 4520 2615
rect 4514 2610 4520 2611
rect 4754 2615 4760 2616
rect 4754 2611 4755 2615
rect 4759 2611 4760 2615
rect 4754 2610 4760 2611
rect 5010 2615 5016 2616
rect 5010 2611 5011 2615
rect 5015 2611 5016 2615
rect 5010 2610 5016 2611
rect 5274 2615 5280 2616
rect 5274 2611 5275 2615
rect 5279 2611 5280 2615
rect 5274 2610 5280 2611
rect 5514 2615 5520 2616
rect 5514 2611 5515 2615
rect 5519 2611 5520 2615
rect 5662 2612 5663 2616
rect 5667 2612 5668 2616
rect 5662 2611 5668 2612
rect 5514 2610 5520 2611
rect 110 2608 116 2609
rect 1934 2608 1940 2609
rect 110 2604 111 2608
rect 115 2604 116 2608
rect 110 2603 116 2604
rect 770 2607 776 2608
rect 770 2603 771 2607
rect 775 2603 776 2607
rect 770 2602 776 2603
rect 906 2607 912 2608
rect 906 2603 907 2607
rect 911 2603 912 2607
rect 906 2602 912 2603
rect 1042 2607 1048 2608
rect 1042 2603 1043 2607
rect 1047 2603 1048 2607
rect 1042 2602 1048 2603
rect 1178 2607 1184 2608
rect 1178 2603 1179 2607
rect 1183 2603 1184 2607
rect 1178 2602 1184 2603
rect 1314 2607 1320 2608
rect 1314 2603 1315 2607
rect 1319 2603 1320 2607
rect 1314 2602 1320 2603
rect 1450 2607 1456 2608
rect 1450 2603 1451 2607
rect 1455 2603 1456 2607
rect 1450 2602 1456 2603
rect 1586 2607 1592 2608
rect 1586 2603 1587 2607
rect 1591 2603 1592 2607
rect 1586 2602 1592 2603
rect 1722 2607 1728 2608
rect 1722 2603 1723 2607
rect 1727 2603 1728 2607
rect 1934 2604 1935 2608
rect 1939 2604 1940 2608
rect 1934 2603 1940 2604
rect 1722 2602 1728 2603
rect 4126 2600 4132 2601
rect 3838 2599 3844 2600
rect 3838 2595 3839 2599
rect 3843 2595 3844 2599
rect 4126 2596 4127 2600
rect 4131 2596 4132 2600
rect 4126 2595 4132 2596
rect 4326 2600 4332 2601
rect 4326 2596 4327 2600
rect 4331 2596 4332 2600
rect 4326 2595 4332 2596
rect 4542 2600 4548 2601
rect 4542 2596 4543 2600
rect 4547 2596 4548 2600
rect 4542 2595 4548 2596
rect 4782 2600 4788 2601
rect 4782 2596 4783 2600
rect 4787 2596 4788 2600
rect 4782 2595 4788 2596
rect 5038 2600 5044 2601
rect 5038 2596 5039 2600
rect 5043 2596 5044 2600
rect 5038 2595 5044 2596
rect 5302 2600 5308 2601
rect 5302 2596 5303 2600
rect 5307 2596 5308 2600
rect 5302 2595 5308 2596
rect 5542 2600 5548 2601
rect 5542 2596 5543 2600
rect 5547 2596 5548 2600
rect 5542 2595 5548 2596
rect 5662 2599 5668 2600
rect 5662 2595 5663 2599
rect 5667 2595 5668 2599
rect 3838 2594 3844 2595
rect 5662 2594 5668 2595
rect 798 2592 804 2593
rect 110 2591 116 2592
rect 110 2587 111 2591
rect 115 2587 116 2591
rect 798 2588 799 2592
rect 803 2588 804 2592
rect 798 2587 804 2588
rect 934 2592 940 2593
rect 934 2588 935 2592
rect 939 2588 940 2592
rect 934 2587 940 2588
rect 1070 2592 1076 2593
rect 1070 2588 1071 2592
rect 1075 2588 1076 2592
rect 1070 2587 1076 2588
rect 1206 2592 1212 2593
rect 1206 2588 1207 2592
rect 1211 2588 1212 2592
rect 1206 2587 1212 2588
rect 1342 2592 1348 2593
rect 1342 2588 1343 2592
rect 1347 2588 1348 2592
rect 1342 2587 1348 2588
rect 1478 2592 1484 2593
rect 1478 2588 1479 2592
rect 1483 2588 1484 2592
rect 1478 2587 1484 2588
rect 1614 2592 1620 2593
rect 1614 2588 1615 2592
rect 1619 2588 1620 2592
rect 1614 2587 1620 2588
rect 1750 2592 1756 2593
rect 1750 2588 1751 2592
rect 1755 2588 1756 2592
rect 1750 2587 1756 2588
rect 1934 2591 1940 2592
rect 1934 2587 1935 2591
rect 1939 2587 1940 2591
rect 110 2586 116 2587
rect 1934 2586 1940 2587
rect 1974 2573 1980 2574
rect 3798 2573 3804 2574
rect 1974 2569 1975 2573
rect 1979 2569 1980 2573
rect 1974 2568 1980 2569
rect 2510 2572 2516 2573
rect 2510 2568 2511 2572
rect 2515 2568 2516 2572
rect 2510 2567 2516 2568
rect 2646 2572 2652 2573
rect 2646 2568 2647 2572
rect 2651 2568 2652 2572
rect 2646 2567 2652 2568
rect 2782 2572 2788 2573
rect 2782 2568 2783 2572
rect 2787 2568 2788 2572
rect 2782 2567 2788 2568
rect 2918 2572 2924 2573
rect 2918 2568 2919 2572
rect 2923 2568 2924 2572
rect 2918 2567 2924 2568
rect 3054 2572 3060 2573
rect 3054 2568 3055 2572
rect 3059 2568 3060 2572
rect 3054 2567 3060 2568
rect 3190 2572 3196 2573
rect 3190 2568 3191 2572
rect 3195 2568 3196 2572
rect 3190 2567 3196 2568
rect 3326 2572 3332 2573
rect 3326 2568 3327 2572
rect 3331 2568 3332 2572
rect 3326 2567 3332 2568
rect 3462 2572 3468 2573
rect 3462 2568 3463 2572
rect 3467 2568 3468 2572
rect 3798 2569 3799 2573
rect 3803 2569 3804 2573
rect 3798 2568 3804 2569
rect 3462 2567 3468 2568
rect 2482 2557 2488 2558
rect 1974 2556 1980 2557
rect 1974 2552 1975 2556
rect 1979 2552 1980 2556
rect 2482 2553 2483 2557
rect 2487 2553 2488 2557
rect 2482 2552 2488 2553
rect 2618 2557 2624 2558
rect 2618 2553 2619 2557
rect 2623 2553 2624 2557
rect 2618 2552 2624 2553
rect 2754 2557 2760 2558
rect 2754 2553 2755 2557
rect 2759 2553 2760 2557
rect 2754 2552 2760 2553
rect 2890 2557 2896 2558
rect 2890 2553 2891 2557
rect 2895 2553 2896 2557
rect 2890 2552 2896 2553
rect 3026 2557 3032 2558
rect 3026 2553 3027 2557
rect 3031 2553 3032 2557
rect 3026 2552 3032 2553
rect 3162 2557 3168 2558
rect 3162 2553 3163 2557
rect 3167 2553 3168 2557
rect 3162 2552 3168 2553
rect 3298 2557 3304 2558
rect 3298 2553 3299 2557
rect 3303 2553 3304 2557
rect 3298 2552 3304 2553
rect 3434 2557 3440 2558
rect 3434 2553 3435 2557
rect 3439 2553 3440 2557
rect 3434 2552 3440 2553
rect 3798 2556 3804 2557
rect 3798 2552 3799 2556
rect 3803 2552 3804 2556
rect 1974 2551 1980 2552
rect 3798 2551 3804 2552
rect 3838 2537 3844 2538
rect 5662 2537 5668 2538
rect 3838 2533 3839 2537
rect 3843 2533 3844 2537
rect 3838 2532 3844 2533
rect 4494 2536 4500 2537
rect 4494 2532 4495 2536
rect 4499 2532 4500 2536
rect 4494 2531 4500 2532
rect 4630 2536 4636 2537
rect 4630 2532 4631 2536
rect 4635 2532 4636 2536
rect 4630 2531 4636 2532
rect 4766 2536 4772 2537
rect 4766 2532 4767 2536
rect 4771 2532 4772 2536
rect 4766 2531 4772 2532
rect 4902 2536 4908 2537
rect 4902 2532 4903 2536
rect 4907 2532 4908 2536
rect 4902 2531 4908 2532
rect 5038 2536 5044 2537
rect 5038 2532 5039 2536
rect 5043 2532 5044 2536
rect 5662 2533 5663 2537
rect 5667 2533 5668 2537
rect 5662 2532 5668 2533
rect 5038 2531 5044 2532
rect 4466 2521 4472 2522
rect 3838 2520 3844 2521
rect 110 2517 116 2518
rect 1934 2517 1940 2518
rect 110 2513 111 2517
rect 115 2513 116 2517
rect 110 2512 116 2513
rect 550 2516 556 2517
rect 550 2512 551 2516
rect 555 2512 556 2516
rect 550 2511 556 2512
rect 686 2516 692 2517
rect 686 2512 687 2516
rect 691 2512 692 2516
rect 686 2511 692 2512
rect 830 2516 836 2517
rect 830 2512 831 2516
rect 835 2512 836 2516
rect 830 2511 836 2512
rect 982 2516 988 2517
rect 982 2512 983 2516
rect 987 2512 988 2516
rect 982 2511 988 2512
rect 1134 2516 1140 2517
rect 1134 2512 1135 2516
rect 1139 2512 1140 2516
rect 1134 2511 1140 2512
rect 1294 2516 1300 2517
rect 1294 2512 1295 2516
rect 1299 2512 1300 2516
rect 1294 2511 1300 2512
rect 1454 2516 1460 2517
rect 1454 2512 1455 2516
rect 1459 2512 1460 2516
rect 1454 2511 1460 2512
rect 1614 2516 1620 2517
rect 1614 2512 1615 2516
rect 1619 2512 1620 2516
rect 1614 2511 1620 2512
rect 1782 2516 1788 2517
rect 1782 2512 1783 2516
rect 1787 2512 1788 2516
rect 1934 2513 1935 2517
rect 1939 2513 1940 2517
rect 3838 2516 3839 2520
rect 3843 2516 3844 2520
rect 4466 2517 4467 2521
rect 4471 2517 4472 2521
rect 4466 2516 4472 2517
rect 4602 2521 4608 2522
rect 4602 2517 4603 2521
rect 4607 2517 4608 2521
rect 4602 2516 4608 2517
rect 4738 2521 4744 2522
rect 4738 2517 4739 2521
rect 4743 2517 4744 2521
rect 4738 2516 4744 2517
rect 4874 2521 4880 2522
rect 4874 2517 4875 2521
rect 4879 2517 4880 2521
rect 4874 2516 4880 2517
rect 5010 2521 5016 2522
rect 5010 2517 5011 2521
rect 5015 2517 5016 2521
rect 5010 2516 5016 2517
rect 5662 2520 5668 2521
rect 5662 2516 5663 2520
rect 5667 2516 5668 2520
rect 3838 2515 3844 2516
rect 5662 2515 5668 2516
rect 1934 2512 1940 2513
rect 1782 2511 1788 2512
rect 522 2501 528 2502
rect 110 2500 116 2501
rect 110 2496 111 2500
rect 115 2496 116 2500
rect 522 2497 523 2501
rect 527 2497 528 2501
rect 522 2496 528 2497
rect 658 2501 664 2502
rect 658 2497 659 2501
rect 663 2497 664 2501
rect 658 2496 664 2497
rect 802 2501 808 2502
rect 802 2497 803 2501
rect 807 2497 808 2501
rect 802 2496 808 2497
rect 954 2501 960 2502
rect 954 2497 955 2501
rect 959 2497 960 2501
rect 954 2496 960 2497
rect 1106 2501 1112 2502
rect 1106 2497 1107 2501
rect 1111 2497 1112 2501
rect 1106 2496 1112 2497
rect 1266 2501 1272 2502
rect 1266 2497 1267 2501
rect 1271 2497 1272 2501
rect 1266 2496 1272 2497
rect 1426 2501 1432 2502
rect 1426 2497 1427 2501
rect 1431 2497 1432 2501
rect 1426 2496 1432 2497
rect 1586 2501 1592 2502
rect 1586 2497 1587 2501
rect 1591 2497 1592 2501
rect 1586 2496 1592 2497
rect 1754 2501 1760 2502
rect 1754 2497 1755 2501
rect 1759 2497 1760 2501
rect 1754 2496 1760 2497
rect 1934 2500 1940 2501
rect 1934 2496 1935 2500
rect 1939 2496 1940 2500
rect 110 2495 116 2496
rect 1934 2495 1940 2496
rect 1974 2408 1980 2409
rect 3798 2408 3804 2409
rect 1974 2404 1975 2408
rect 1979 2404 1980 2408
rect 1974 2403 1980 2404
rect 2306 2407 2312 2408
rect 2306 2403 2307 2407
rect 2311 2403 2312 2407
rect 2306 2402 2312 2403
rect 2514 2407 2520 2408
rect 2514 2403 2515 2407
rect 2519 2403 2520 2407
rect 2514 2402 2520 2403
rect 2714 2407 2720 2408
rect 2714 2403 2715 2407
rect 2719 2403 2720 2407
rect 2714 2402 2720 2403
rect 2906 2407 2912 2408
rect 2906 2403 2907 2407
rect 2911 2403 2912 2407
rect 2906 2402 2912 2403
rect 3098 2407 3104 2408
rect 3098 2403 3099 2407
rect 3103 2403 3104 2407
rect 3098 2402 3104 2403
rect 3282 2407 3288 2408
rect 3282 2403 3283 2407
rect 3287 2403 3288 2407
rect 3282 2402 3288 2403
rect 3466 2407 3472 2408
rect 3466 2403 3467 2407
rect 3471 2403 3472 2407
rect 3466 2402 3472 2403
rect 3650 2407 3656 2408
rect 3650 2403 3651 2407
rect 3655 2403 3656 2407
rect 3798 2404 3799 2408
rect 3803 2404 3804 2408
rect 3798 2403 3804 2404
rect 3650 2402 3656 2403
rect 2334 2392 2340 2393
rect 1974 2391 1980 2392
rect 1974 2387 1975 2391
rect 1979 2387 1980 2391
rect 2334 2388 2335 2392
rect 2339 2388 2340 2392
rect 2334 2387 2340 2388
rect 2542 2392 2548 2393
rect 2542 2388 2543 2392
rect 2547 2388 2548 2392
rect 2542 2387 2548 2388
rect 2742 2392 2748 2393
rect 2742 2388 2743 2392
rect 2747 2388 2748 2392
rect 2742 2387 2748 2388
rect 2934 2392 2940 2393
rect 2934 2388 2935 2392
rect 2939 2388 2940 2392
rect 2934 2387 2940 2388
rect 3126 2392 3132 2393
rect 3126 2388 3127 2392
rect 3131 2388 3132 2392
rect 3126 2387 3132 2388
rect 3310 2392 3316 2393
rect 3310 2388 3311 2392
rect 3315 2388 3316 2392
rect 3310 2387 3316 2388
rect 3494 2392 3500 2393
rect 3494 2388 3495 2392
rect 3499 2388 3500 2392
rect 3494 2387 3500 2388
rect 3678 2392 3684 2393
rect 3678 2388 3679 2392
rect 3683 2388 3684 2392
rect 3678 2387 3684 2388
rect 3798 2391 3804 2392
rect 3798 2387 3799 2391
rect 3803 2387 3804 2391
rect 1974 2386 1980 2387
rect 3798 2386 3804 2387
rect 3838 2372 3844 2373
rect 5662 2372 5668 2373
rect 3838 2368 3839 2372
rect 3843 2368 3844 2372
rect 3838 2367 3844 2368
rect 4698 2371 4704 2372
rect 4698 2367 4699 2371
rect 4703 2367 4704 2371
rect 4698 2366 4704 2367
rect 4834 2371 4840 2372
rect 4834 2367 4835 2371
rect 4839 2367 4840 2371
rect 4834 2366 4840 2367
rect 4970 2371 4976 2372
rect 4970 2367 4971 2371
rect 4975 2367 4976 2371
rect 4970 2366 4976 2367
rect 5106 2371 5112 2372
rect 5106 2367 5107 2371
rect 5111 2367 5112 2371
rect 5106 2366 5112 2367
rect 5242 2371 5248 2372
rect 5242 2367 5243 2371
rect 5247 2367 5248 2371
rect 5242 2366 5248 2367
rect 5378 2371 5384 2372
rect 5378 2367 5379 2371
rect 5383 2367 5384 2371
rect 5378 2366 5384 2367
rect 5514 2371 5520 2372
rect 5514 2367 5515 2371
rect 5519 2367 5520 2371
rect 5662 2368 5663 2372
rect 5667 2368 5668 2372
rect 5662 2367 5668 2368
rect 5514 2366 5520 2367
rect 110 2356 116 2357
rect 1934 2356 1940 2357
rect 4726 2356 4732 2357
rect 110 2352 111 2356
rect 115 2352 116 2356
rect 110 2351 116 2352
rect 130 2355 136 2356
rect 130 2351 131 2355
rect 135 2351 136 2355
rect 130 2350 136 2351
rect 338 2355 344 2356
rect 338 2351 339 2355
rect 343 2351 344 2355
rect 338 2350 344 2351
rect 562 2355 568 2356
rect 562 2351 563 2355
rect 567 2351 568 2355
rect 562 2350 568 2351
rect 802 2355 808 2356
rect 802 2351 803 2355
rect 807 2351 808 2355
rect 802 2350 808 2351
rect 1042 2355 1048 2356
rect 1042 2351 1043 2355
rect 1047 2351 1048 2355
rect 1042 2350 1048 2351
rect 1290 2355 1296 2356
rect 1290 2351 1291 2355
rect 1295 2351 1296 2355
rect 1290 2350 1296 2351
rect 1546 2355 1552 2356
rect 1546 2351 1547 2355
rect 1551 2351 1552 2355
rect 1546 2350 1552 2351
rect 1786 2355 1792 2356
rect 1786 2351 1787 2355
rect 1791 2351 1792 2355
rect 1934 2352 1935 2356
rect 1939 2352 1940 2356
rect 1934 2351 1940 2352
rect 3838 2355 3844 2356
rect 3838 2351 3839 2355
rect 3843 2351 3844 2355
rect 4726 2352 4727 2356
rect 4731 2352 4732 2356
rect 4726 2351 4732 2352
rect 4862 2356 4868 2357
rect 4862 2352 4863 2356
rect 4867 2352 4868 2356
rect 4862 2351 4868 2352
rect 4998 2356 5004 2357
rect 4998 2352 4999 2356
rect 5003 2352 5004 2356
rect 4998 2351 5004 2352
rect 5134 2356 5140 2357
rect 5134 2352 5135 2356
rect 5139 2352 5140 2356
rect 5134 2351 5140 2352
rect 5270 2356 5276 2357
rect 5270 2352 5271 2356
rect 5275 2352 5276 2356
rect 5270 2351 5276 2352
rect 5406 2356 5412 2357
rect 5406 2352 5407 2356
rect 5411 2352 5412 2356
rect 5406 2351 5412 2352
rect 5542 2356 5548 2357
rect 5542 2352 5543 2356
rect 5547 2352 5548 2356
rect 5542 2351 5548 2352
rect 5662 2355 5668 2356
rect 5662 2351 5663 2355
rect 5667 2351 5668 2355
rect 1786 2350 1792 2351
rect 3838 2350 3844 2351
rect 5662 2350 5668 2351
rect 158 2340 164 2341
rect 110 2339 116 2340
rect 110 2335 111 2339
rect 115 2335 116 2339
rect 158 2336 159 2340
rect 163 2336 164 2340
rect 158 2335 164 2336
rect 366 2340 372 2341
rect 366 2336 367 2340
rect 371 2336 372 2340
rect 366 2335 372 2336
rect 590 2340 596 2341
rect 590 2336 591 2340
rect 595 2336 596 2340
rect 590 2335 596 2336
rect 830 2340 836 2341
rect 830 2336 831 2340
rect 835 2336 836 2340
rect 830 2335 836 2336
rect 1070 2340 1076 2341
rect 1070 2336 1071 2340
rect 1075 2336 1076 2340
rect 1070 2335 1076 2336
rect 1318 2340 1324 2341
rect 1318 2336 1319 2340
rect 1323 2336 1324 2340
rect 1318 2335 1324 2336
rect 1574 2340 1580 2341
rect 1574 2336 1575 2340
rect 1579 2336 1580 2340
rect 1574 2335 1580 2336
rect 1814 2340 1820 2341
rect 1814 2336 1815 2340
rect 1819 2336 1820 2340
rect 1814 2335 1820 2336
rect 1934 2339 1940 2340
rect 1934 2335 1935 2339
rect 1939 2335 1940 2339
rect 110 2334 116 2335
rect 1934 2334 1940 2335
rect 1974 2325 1980 2326
rect 3798 2325 3804 2326
rect 1974 2321 1975 2325
rect 1979 2321 1980 2325
rect 1974 2320 1980 2321
rect 2222 2324 2228 2325
rect 2222 2320 2223 2324
rect 2227 2320 2228 2324
rect 2222 2319 2228 2320
rect 2502 2324 2508 2325
rect 2502 2320 2503 2324
rect 2507 2320 2508 2324
rect 2502 2319 2508 2320
rect 2766 2324 2772 2325
rect 2766 2320 2767 2324
rect 2771 2320 2772 2324
rect 2766 2319 2772 2320
rect 3006 2324 3012 2325
rect 3006 2320 3007 2324
rect 3011 2320 3012 2324
rect 3006 2319 3012 2320
rect 3238 2324 3244 2325
rect 3238 2320 3239 2324
rect 3243 2320 3244 2324
rect 3238 2319 3244 2320
rect 3470 2324 3476 2325
rect 3470 2320 3471 2324
rect 3475 2320 3476 2324
rect 3470 2319 3476 2320
rect 3678 2324 3684 2325
rect 3678 2320 3679 2324
rect 3683 2320 3684 2324
rect 3798 2321 3799 2325
rect 3803 2321 3804 2325
rect 3798 2320 3804 2321
rect 3678 2319 3684 2320
rect 2194 2309 2200 2310
rect 1974 2308 1980 2309
rect 1974 2304 1975 2308
rect 1979 2304 1980 2308
rect 2194 2305 2195 2309
rect 2199 2305 2200 2309
rect 2194 2304 2200 2305
rect 2474 2309 2480 2310
rect 2474 2305 2475 2309
rect 2479 2305 2480 2309
rect 2474 2304 2480 2305
rect 2738 2309 2744 2310
rect 2738 2305 2739 2309
rect 2743 2305 2744 2309
rect 2738 2304 2744 2305
rect 2978 2309 2984 2310
rect 2978 2305 2979 2309
rect 2983 2305 2984 2309
rect 2978 2304 2984 2305
rect 3210 2309 3216 2310
rect 3210 2305 3211 2309
rect 3215 2305 3216 2309
rect 3210 2304 3216 2305
rect 3442 2309 3448 2310
rect 3442 2305 3443 2309
rect 3447 2305 3448 2309
rect 3442 2304 3448 2305
rect 3650 2309 3656 2310
rect 3650 2305 3651 2309
rect 3655 2305 3656 2309
rect 3650 2304 3656 2305
rect 3798 2308 3804 2309
rect 3798 2304 3799 2308
rect 3803 2304 3804 2308
rect 1974 2303 1980 2304
rect 3798 2303 3804 2304
rect 3838 2285 3844 2286
rect 5662 2285 5668 2286
rect 3838 2281 3839 2285
rect 3843 2281 3844 2285
rect 3838 2280 3844 2281
rect 3886 2284 3892 2285
rect 3886 2280 3887 2284
rect 3891 2280 3892 2284
rect 3886 2279 3892 2280
rect 4182 2284 4188 2285
rect 4182 2280 4183 2284
rect 4187 2280 4188 2284
rect 4182 2279 4188 2280
rect 4494 2284 4500 2285
rect 4494 2280 4495 2284
rect 4499 2280 4500 2284
rect 4494 2279 4500 2280
rect 4790 2284 4796 2285
rect 4790 2280 4791 2284
rect 4795 2280 4796 2284
rect 4790 2279 4796 2280
rect 5086 2284 5092 2285
rect 5086 2280 5087 2284
rect 5091 2280 5092 2284
rect 5086 2279 5092 2280
rect 5382 2284 5388 2285
rect 5382 2280 5383 2284
rect 5387 2280 5388 2284
rect 5662 2281 5663 2285
rect 5667 2281 5668 2285
rect 5662 2280 5668 2281
rect 5382 2279 5388 2280
rect 110 2277 116 2278
rect 1934 2277 1940 2278
rect 110 2273 111 2277
rect 115 2273 116 2277
rect 110 2272 116 2273
rect 158 2276 164 2277
rect 158 2272 159 2276
rect 163 2272 164 2276
rect 158 2271 164 2272
rect 318 2276 324 2277
rect 318 2272 319 2276
rect 323 2272 324 2276
rect 318 2271 324 2272
rect 550 2276 556 2277
rect 550 2272 551 2276
rect 555 2272 556 2276
rect 550 2271 556 2272
rect 830 2276 836 2277
rect 830 2272 831 2276
rect 835 2272 836 2276
rect 830 2271 836 2272
rect 1150 2276 1156 2277
rect 1150 2272 1151 2276
rect 1155 2272 1156 2276
rect 1150 2271 1156 2272
rect 1494 2276 1500 2277
rect 1494 2272 1495 2276
rect 1499 2272 1500 2276
rect 1494 2271 1500 2272
rect 1814 2276 1820 2277
rect 1814 2272 1815 2276
rect 1819 2272 1820 2276
rect 1934 2273 1935 2277
rect 1939 2273 1940 2277
rect 1934 2272 1940 2273
rect 1814 2271 1820 2272
rect 3858 2269 3864 2270
rect 3838 2268 3844 2269
rect 3838 2264 3839 2268
rect 3843 2264 3844 2268
rect 3858 2265 3859 2269
rect 3863 2265 3864 2269
rect 3858 2264 3864 2265
rect 4154 2269 4160 2270
rect 4154 2265 4155 2269
rect 4159 2265 4160 2269
rect 4154 2264 4160 2265
rect 4466 2269 4472 2270
rect 4466 2265 4467 2269
rect 4471 2265 4472 2269
rect 4466 2264 4472 2265
rect 4762 2269 4768 2270
rect 4762 2265 4763 2269
rect 4767 2265 4768 2269
rect 4762 2264 4768 2265
rect 5058 2269 5064 2270
rect 5058 2265 5059 2269
rect 5063 2265 5064 2269
rect 5058 2264 5064 2265
rect 5354 2269 5360 2270
rect 5354 2265 5355 2269
rect 5359 2265 5360 2269
rect 5354 2264 5360 2265
rect 5662 2268 5668 2269
rect 5662 2264 5663 2268
rect 5667 2264 5668 2268
rect 3838 2263 3844 2264
rect 5662 2263 5668 2264
rect 130 2261 136 2262
rect 110 2260 116 2261
rect 110 2256 111 2260
rect 115 2256 116 2260
rect 130 2257 131 2261
rect 135 2257 136 2261
rect 130 2256 136 2257
rect 290 2261 296 2262
rect 290 2257 291 2261
rect 295 2257 296 2261
rect 290 2256 296 2257
rect 522 2261 528 2262
rect 522 2257 523 2261
rect 527 2257 528 2261
rect 522 2256 528 2257
rect 802 2261 808 2262
rect 802 2257 803 2261
rect 807 2257 808 2261
rect 802 2256 808 2257
rect 1122 2261 1128 2262
rect 1122 2257 1123 2261
rect 1127 2257 1128 2261
rect 1122 2256 1128 2257
rect 1466 2261 1472 2262
rect 1466 2257 1467 2261
rect 1471 2257 1472 2261
rect 1466 2256 1472 2257
rect 1786 2261 1792 2262
rect 1786 2257 1787 2261
rect 1791 2257 1792 2261
rect 1786 2256 1792 2257
rect 1934 2260 1940 2261
rect 1934 2256 1935 2260
rect 1939 2256 1940 2260
rect 110 2255 116 2256
rect 1934 2255 1940 2256
rect 1974 2176 1980 2177
rect 3798 2176 3804 2177
rect 1974 2172 1975 2176
rect 1979 2172 1980 2176
rect 1974 2171 1980 2172
rect 1994 2175 2000 2176
rect 1994 2171 1995 2175
rect 1999 2171 2000 2175
rect 1994 2170 2000 2171
rect 2154 2175 2160 2176
rect 2154 2171 2155 2175
rect 2159 2171 2160 2175
rect 2154 2170 2160 2171
rect 2386 2175 2392 2176
rect 2386 2171 2387 2175
rect 2391 2171 2392 2175
rect 2386 2170 2392 2171
rect 2666 2175 2672 2176
rect 2666 2171 2667 2175
rect 2671 2171 2672 2175
rect 2666 2170 2672 2171
rect 2986 2175 2992 2176
rect 2986 2171 2987 2175
rect 2991 2171 2992 2175
rect 2986 2170 2992 2171
rect 3330 2175 3336 2176
rect 3330 2171 3331 2175
rect 3335 2171 3336 2175
rect 3330 2170 3336 2171
rect 3650 2175 3656 2176
rect 3650 2171 3651 2175
rect 3655 2171 3656 2175
rect 3798 2172 3799 2176
rect 3803 2172 3804 2176
rect 3798 2171 3804 2172
rect 3650 2170 3656 2171
rect 2022 2160 2028 2161
rect 1974 2159 1980 2160
rect 1974 2155 1975 2159
rect 1979 2155 1980 2159
rect 2022 2156 2023 2160
rect 2027 2156 2028 2160
rect 2022 2155 2028 2156
rect 2182 2160 2188 2161
rect 2182 2156 2183 2160
rect 2187 2156 2188 2160
rect 2182 2155 2188 2156
rect 2414 2160 2420 2161
rect 2414 2156 2415 2160
rect 2419 2156 2420 2160
rect 2414 2155 2420 2156
rect 2694 2160 2700 2161
rect 2694 2156 2695 2160
rect 2699 2156 2700 2160
rect 2694 2155 2700 2156
rect 3014 2160 3020 2161
rect 3014 2156 3015 2160
rect 3019 2156 3020 2160
rect 3014 2155 3020 2156
rect 3358 2160 3364 2161
rect 3358 2156 3359 2160
rect 3363 2156 3364 2160
rect 3358 2155 3364 2156
rect 3678 2160 3684 2161
rect 3678 2156 3679 2160
rect 3683 2156 3684 2160
rect 3678 2155 3684 2156
rect 3798 2159 3804 2160
rect 3798 2155 3799 2159
rect 3803 2155 3804 2159
rect 1974 2154 1980 2155
rect 3798 2154 3804 2155
rect 3838 2132 3844 2133
rect 5662 2132 5668 2133
rect 3838 2128 3839 2132
rect 3843 2128 3844 2132
rect 3838 2127 3844 2128
rect 3858 2131 3864 2132
rect 3858 2127 3859 2131
rect 3863 2127 3864 2131
rect 3858 2126 3864 2127
rect 3994 2131 4000 2132
rect 3994 2127 3995 2131
rect 3999 2127 4000 2131
rect 3994 2126 4000 2127
rect 4130 2131 4136 2132
rect 4130 2127 4131 2131
rect 4135 2127 4136 2131
rect 4130 2126 4136 2127
rect 4266 2131 4272 2132
rect 4266 2127 4267 2131
rect 4271 2127 4272 2131
rect 4266 2126 4272 2127
rect 4402 2131 4408 2132
rect 4402 2127 4403 2131
rect 4407 2127 4408 2131
rect 4402 2126 4408 2127
rect 4538 2131 4544 2132
rect 4538 2127 4539 2131
rect 4543 2127 4544 2131
rect 4538 2126 4544 2127
rect 4698 2131 4704 2132
rect 4698 2127 4699 2131
rect 4703 2127 4704 2131
rect 4698 2126 4704 2127
rect 4890 2131 4896 2132
rect 4890 2127 4891 2131
rect 4895 2127 4896 2131
rect 4890 2126 4896 2127
rect 5098 2131 5104 2132
rect 5098 2127 5099 2131
rect 5103 2127 5104 2131
rect 5098 2126 5104 2127
rect 5314 2131 5320 2132
rect 5314 2127 5315 2131
rect 5319 2127 5320 2131
rect 5314 2126 5320 2127
rect 5514 2131 5520 2132
rect 5514 2127 5515 2131
rect 5519 2127 5520 2131
rect 5662 2128 5663 2132
rect 5667 2128 5668 2132
rect 5662 2127 5668 2128
rect 5514 2126 5520 2127
rect 3886 2116 3892 2117
rect 3838 2115 3844 2116
rect 3838 2111 3839 2115
rect 3843 2111 3844 2115
rect 3886 2112 3887 2116
rect 3891 2112 3892 2116
rect 3886 2111 3892 2112
rect 4022 2116 4028 2117
rect 4022 2112 4023 2116
rect 4027 2112 4028 2116
rect 4022 2111 4028 2112
rect 4158 2116 4164 2117
rect 4158 2112 4159 2116
rect 4163 2112 4164 2116
rect 4158 2111 4164 2112
rect 4294 2116 4300 2117
rect 4294 2112 4295 2116
rect 4299 2112 4300 2116
rect 4294 2111 4300 2112
rect 4430 2116 4436 2117
rect 4430 2112 4431 2116
rect 4435 2112 4436 2116
rect 4430 2111 4436 2112
rect 4566 2116 4572 2117
rect 4566 2112 4567 2116
rect 4571 2112 4572 2116
rect 4566 2111 4572 2112
rect 4726 2116 4732 2117
rect 4726 2112 4727 2116
rect 4731 2112 4732 2116
rect 4726 2111 4732 2112
rect 4918 2116 4924 2117
rect 4918 2112 4919 2116
rect 4923 2112 4924 2116
rect 4918 2111 4924 2112
rect 5126 2116 5132 2117
rect 5126 2112 5127 2116
rect 5131 2112 5132 2116
rect 5126 2111 5132 2112
rect 5342 2116 5348 2117
rect 5342 2112 5343 2116
rect 5347 2112 5348 2116
rect 5342 2111 5348 2112
rect 5542 2116 5548 2117
rect 5542 2112 5543 2116
rect 5547 2112 5548 2116
rect 5542 2111 5548 2112
rect 5662 2115 5668 2116
rect 5662 2111 5663 2115
rect 5667 2111 5668 2115
rect 3838 2110 3844 2111
rect 5662 2110 5668 2111
rect 110 2104 116 2105
rect 1934 2104 1940 2105
rect 110 2100 111 2104
rect 115 2100 116 2104
rect 110 2099 116 2100
rect 290 2103 296 2104
rect 290 2099 291 2103
rect 295 2099 296 2103
rect 290 2098 296 2099
rect 482 2103 488 2104
rect 482 2099 483 2103
rect 487 2099 488 2103
rect 482 2098 488 2099
rect 690 2103 696 2104
rect 690 2099 691 2103
rect 695 2099 696 2103
rect 690 2098 696 2099
rect 914 2103 920 2104
rect 914 2099 915 2103
rect 919 2099 920 2103
rect 914 2098 920 2099
rect 1146 2103 1152 2104
rect 1146 2099 1147 2103
rect 1151 2099 1152 2103
rect 1146 2098 1152 2099
rect 1386 2103 1392 2104
rect 1386 2099 1387 2103
rect 1391 2099 1392 2103
rect 1386 2098 1392 2099
rect 1634 2103 1640 2104
rect 1634 2099 1635 2103
rect 1639 2099 1640 2103
rect 1934 2100 1935 2104
rect 1939 2100 1940 2104
rect 1934 2099 1940 2100
rect 1634 2098 1640 2099
rect 318 2088 324 2089
rect 110 2087 116 2088
rect 110 2083 111 2087
rect 115 2083 116 2087
rect 318 2084 319 2088
rect 323 2084 324 2088
rect 318 2083 324 2084
rect 510 2088 516 2089
rect 510 2084 511 2088
rect 515 2084 516 2088
rect 510 2083 516 2084
rect 718 2088 724 2089
rect 718 2084 719 2088
rect 723 2084 724 2088
rect 718 2083 724 2084
rect 942 2088 948 2089
rect 942 2084 943 2088
rect 947 2084 948 2088
rect 942 2083 948 2084
rect 1174 2088 1180 2089
rect 1174 2084 1175 2088
rect 1179 2084 1180 2088
rect 1174 2083 1180 2084
rect 1414 2088 1420 2089
rect 1414 2084 1415 2088
rect 1419 2084 1420 2088
rect 1414 2083 1420 2084
rect 1662 2088 1668 2089
rect 1662 2084 1663 2088
rect 1667 2084 1668 2088
rect 1662 2083 1668 2084
rect 1934 2087 1940 2088
rect 1934 2083 1935 2087
rect 1939 2083 1940 2087
rect 110 2082 116 2083
rect 1934 2082 1940 2083
rect 3838 2037 3844 2038
rect 5662 2037 5668 2038
rect 3838 2033 3839 2037
rect 3843 2033 3844 2037
rect 3838 2032 3844 2033
rect 3886 2036 3892 2037
rect 3886 2032 3887 2036
rect 3891 2032 3892 2036
rect 3886 2031 3892 2032
rect 4022 2036 4028 2037
rect 4022 2032 4023 2036
rect 4027 2032 4028 2036
rect 4022 2031 4028 2032
rect 4158 2036 4164 2037
rect 4158 2032 4159 2036
rect 4163 2032 4164 2036
rect 4158 2031 4164 2032
rect 4294 2036 4300 2037
rect 4294 2032 4295 2036
rect 4299 2032 4300 2036
rect 4294 2031 4300 2032
rect 4430 2036 4436 2037
rect 4430 2032 4431 2036
rect 4435 2032 4436 2036
rect 4430 2031 4436 2032
rect 4566 2036 4572 2037
rect 4566 2032 4567 2036
rect 4571 2032 4572 2036
rect 4566 2031 4572 2032
rect 4718 2036 4724 2037
rect 4718 2032 4719 2036
rect 4723 2032 4724 2036
rect 4718 2031 4724 2032
rect 4894 2036 4900 2037
rect 4894 2032 4895 2036
rect 4899 2032 4900 2036
rect 4894 2031 4900 2032
rect 5086 2036 5092 2037
rect 5086 2032 5087 2036
rect 5091 2032 5092 2036
rect 5086 2031 5092 2032
rect 5278 2036 5284 2037
rect 5278 2032 5279 2036
rect 5283 2032 5284 2036
rect 5278 2031 5284 2032
rect 5478 2036 5484 2037
rect 5478 2032 5479 2036
rect 5483 2032 5484 2036
rect 5662 2033 5663 2037
rect 5667 2033 5668 2037
rect 5662 2032 5668 2033
rect 5478 2031 5484 2032
rect 110 2025 116 2026
rect 1934 2025 1940 2026
rect 110 2021 111 2025
rect 115 2021 116 2025
rect 110 2020 116 2021
rect 262 2024 268 2025
rect 262 2020 263 2024
rect 267 2020 268 2024
rect 262 2019 268 2020
rect 398 2024 404 2025
rect 398 2020 399 2024
rect 403 2020 404 2024
rect 398 2019 404 2020
rect 534 2024 540 2025
rect 534 2020 535 2024
rect 539 2020 540 2024
rect 534 2019 540 2020
rect 678 2024 684 2025
rect 678 2020 679 2024
rect 683 2020 684 2024
rect 678 2019 684 2020
rect 822 2024 828 2025
rect 822 2020 823 2024
rect 827 2020 828 2024
rect 822 2019 828 2020
rect 966 2024 972 2025
rect 966 2020 967 2024
rect 971 2020 972 2024
rect 966 2019 972 2020
rect 1110 2024 1116 2025
rect 1110 2020 1111 2024
rect 1115 2020 1116 2024
rect 1110 2019 1116 2020
rect 1254 2024 1260 2025
rect 1254 2020 1255 2024
rect 1259 2020 1260 2024
rect 1254 2019 1260 2020
rect 1398 2024 1404 2025
rect 1398 2020 1399 2024
rect 1403 2020 1404 2024
rect 1398 2019 1404 2020
rect 1542 2024 1548 2025
rect 1542 2020 1543 2024
rect 1547 2020 1548 2024
rect 1542 2019 1548 2020
rect 1678 2024 1684 2025
rect 1678 2020 1679 2024
rect 1683 2020 1684 2024
rect 1678 2019 1684 2020
rect 1814 2024 1820 2025
rect 1814 2020 1815 2024
rect 1819 2020 1820 2024
rect 1934 2021 1935 2025
rect 1939 2021 1940 2025
rect 3858 2021 3864 2022
rect 1934 2020 1940 2021
rect 3838 2020 3844 2021
rect 1814 2019 1820 2020
rect 3838 2016 3839 2020
rect 3843 2016 3844 2020
rect 3858 2017 3859 2021
rect 3863 2017 3864 2021
rect 3858 2016 3864 2017
rect 3994 2021 4000 2022
rect 3994 2017 3995 2021
rect 3999 2017 4000 2021
rect 3994 2016 4000 2017
rect 4130 2021 4136 2022
rect 4130 2017 4131 2021
rect 4135 2017 4136 2021
rect 4130 2016 4136 2017
rect 4266 2021 4272 2022
rect 4266 2017 4267 2021
rect 4271 2017 4272 2021
rect 4266 2016 4272 2017
rect 4402 2021 4408 2022
rect 4402 2017 4403 2021
rect 4407 2017 4408 2021
rect 4402 2016 4408 2017
rect 4538 2021 4544 2022
rect 4538 2017 4539 2021
rect 4543 2017 4544 2021
rect 4538 2016 4544 2017
rect 4690 2021 4696 2022
rect 4690 2017 4691 2021
rect 4695 2017 4696 2021
rect 4690 2016 4696 2017
rect 4866 2021 4872 2022
rect 4866 2017 4867 2021
rect 4871 2017 4872 2021
rect 4866 2016 4872 2017
rect 5058 2021 5064 2022
rect 5058 2017 5059 2021
rect 5063 2017 5064 2021
rect 5058 2016 5064 2017
rect 5250 2021 5256 2022
rect 5250 2017 5251 2021
rect 5255 2017 5256 2021
rect 5250 2016 5256 2017
rect 5450 2021 5456 2022
rect 5450 2017 5451 2021
rect 5455 2017 5456 2021
rect 5450 2016 5456 2017
rect 5662 2020 5668 2021
rect 5662 2016 5663 2020
rect 5667 2016 5668 2020
rect 3838 2015 3844 2016
rect 5662 2015 5668 2016
rect 234 2009 240 2010
rect 110 2008 116 2009
rect 110 2004 111 2008
rect 115 2004 116 2008
rect 234 2005 235 2009
rect 239 2005 240 2009
rect 234 2004 240 2005
rect 370 2009 376 2010
rect 370 2005 371 2009
rect 375 2005 376 2009
rect 370 2004 376 2005
rect 506 2009 512 2010
rect 506 2005 507 2009
rect 511 2005 512 2009
rect 506 2004 512 2005
rect 650 2009 656 2010
rect 650 2005 651 2009
rect 655 2005 656 2009
rect 650 2004 656 2005
rect 794 2009 800 2010
rect 794 2005 795 2009
rect 799 2005 800 2009
rect 794 2004 800 2005
rect 938 2009 944 2010
rect 938 2005 939 2009
rect 943 2005 944 2009
rect 938 2004 944 2005
rect 1082 2009 1088 2010
rect 1082 2005 1083 2009
rect 1087 2005 1088 2009
rect 1082 2004 1088 2005
rect 1226 2009 1232 2010
rect 1226 2005 1227 2009
rect 1231 2005 1232 2009
rect 1226 2004 1232 2005
rect 1370 2009 1376 2010
rect 1370 2005 1371 2009
rect 1375 2005 1376 2009
rect 1370 2004 1376 2005
rect 1514 2009 1520 2010
rect 1514 2005 1515 2009
rect 1519 2005 1520 2009
rect 1514 2004 1520 2005
rect 1650 2009 1656 2010
rect 1650 2005 1651 2009
rect 1655 2005 1656 2009
rect 1650 2004 1656 2005
rect 1786 2009 1792 2010
rect 1786 2005 1787 2009
rect 1791 2005 1792 2009
rect 1786 2004 1792 2005
rect 1934 2008 1940 2009
rect 1934 2004 1935 2008
rect 1939 2004 1940 2008
rect 110 2003 116 2004
rect 1934 2003 1940 2004
rect 1974 1901 1980 1902
rect 3798 1901 3804 1902
rect 1974 1897 1975 1901
rect 1979 1897 1980 1901
rect 1974 1896 1980 1897
rect 3134 1900 3140 1901
rect 3134 1896 3135 1900
rect 3139 1896 3140 1900
rect 3134 1895 3140 1896
rect 3270 1900 3276 1901
rect 3270 1896 3271 1900
rect 3275 1896 3276 1900
rect 3270 1895 3276 1896
rect 3406 1900 3412 1901
rect 3406 1896 3407 1900
rect 3411 1896 3412 1900
rect 3406 1895 3412 1896
rect 3542 1900 3548 1901
rect 3542 1896 3543 1900
rect 3547 1896 3548 1900
rect 3542 1895 3548 1896
rect 3678 1900 3684 1901
rect 3678 1896 3679 1900
rect 3683 1896 3684 1900
rect 3798 1897 3799 1901
rect 3803 1897 3804 1901
rect 3798 1896 3804 1897
rect 3678 1895 3684 1896
rect 3838 1888 3844 1889
rect 5662 1888 5668 1889
rect 3106 1885 3112 1886
rect 1974 1884 1980 1885
rect 1974 1880 1975 1884
rect 1979 1880 1980 1884
rect 3106 1881 3107 1885
rect 3111 1881 3112 1885
rect 3106 1880 3112 1881
rect 3242 1885 3248 1886
rect 3242 1881 3243 1885
rect 3247 1881 3248 1885
rect 3242 1880 3248 1881
rect 3378 1885 3384 1886
rect 3378 1881 3379 1885
rect 3383 1881 3384 1885
rect 3378 1880 3384 1881
rect 3514 1885 3520 1886
rect 3514 1881 3515 1885
rect 3519 1881 3520 1885
rect 3514 1880 3520 1881
rect 3650 1885 3656 1886
rect 3650 1881 3651 1885
rect 3655 1881 3656 1885
rect 3650 1880 3656 1881
rect 3798 1884 3804 1885
rect 3798 1880 3799 1884
rect 3803 1880 3804 1884
rect 3838 1884 3839 1888
rect 3843 1884 3844 1888
rect 3838 1883 3844 1884
rect 3858 1887 3864 1888
rect 3858 1883 3859 1887
rect 3863 1883 3864 1887
rect 3858 1882 3864 1883
rect 4042 1887 4048 1888
rect 4042 1883 4043 1887
rect 4047 1883 4048 1887
rect 4042 1882 4048 1883
rect 4282 1887 4288 1888
rect 4282 1883 4283 1887
rect 4287 1883 4288 1887
rect 4282 1882 4288 1883
rect 4562 1887 4568 1888
rect 4562 1883 4563 1887
rect 4567 1883 4568 1887
rect 4562 1882 4568 1883
rect 4874 1887 4880 1888
rect 4874 1883 4875 1887
rect 4879 1883 4880 1887
rect 4874 1882 4880 1883
rect 5202 1887 5208 1888
rect 5202 1883 5203 1887
rect 5207 1883 5208 1887
rect 5202 1882 5208 1883
rect 5514 1887 5520 1888
rect 5514 1883 5515 1887
rect 5519 1883 5520 1887
rect 5662 1884 5663 1888
rect 5667 1884 5668 1888
rect 5662 1883 5668 1884
rect 5514 1882 5520 1883
rect 1974 1879 1980 1880
rect 3798 1879 3804 1880
rect 3886 1872 3892 1873
rect 3838 1871 3844 1872
rect 3838 1867 3839 1871
rect 3843 1867 3844 1871
rect 3886 1868 3887 1872
rect 3891 1868 3892 1872
rect 3886 1867 3892 1868
rect 4070 1872 4076 1873
rect 4070 1868 4071 1872
rect 4075 1868 4076 1872
rect 4070 1867 4076 1868
rect 4310 1872 4316 1873
rect 4310 1868 4311 1872
rect 4315 1868 4316 1872
rect 4310 1867 4316 1868
rect 4590 1872 4596 1873
rect 4590 1868 4591 1872
rect 4595 1868 4596 1872
rect 4590 1867 4596 1868
rect 4902 1872 4908 1873
rect 4902 1868 4903 1872
rect 4907 1868 4908 1872
rect 4902 1867 4908 1868
rect 5230 1872 5236 1873
rect 5230 1868 5231 1872
rect 5235 1868 5236 1872
rect 5230 1867 5236 1868
rect 5542 1872 5548 1873
rect 5542 1868 5543 1872
rect 5547 1868 5548 1872
rect 5542 1867 5548 1868
rect 5662 1871 5668 1872
rect 5662 1867 5663 1871
rect 5667 1867 5668 1871
rect 3838 1866 3844 1867
rect 5662 1866 5668 1867
rect 110 1864 116 1865
rect 1934 1864 1940 1865
rect 110 1860 111 1864
rect 115 1860 116 1864
rect 110 1859 116 1860
rect 234 1863 240 1864
rect 234 1859 235 1863
rect 239 1859 240 1863
rect 234 1858 240 1859
rect 434 1863 440 1864
rect 434 1859 435 1863
rect 439 1859 440 1863
rect 434 1858 440 1859
rect 626 1863 632 1864
rect 626 1859 627 1863
rect 631 1859 632 1863
rect 626 1858 632 1859
rect 810 1863 816 1864
rect 810 1859 811 1863
rect 815 1859 816 1863
rect 810 1858 816 1859
rect 986 1863 992 1864
rect 986 1859 987 1863
rect 991 1859 992 1863
rect 986 1858 992 1859
rect 1154 1863 1160 1864
rect 1154 1859 1155 1863
rect 1159 1859 1160 1863
rect 1154 1858 1160 1859
rect 1322 1863 1328 1864
rect 1322 1859 1323 1863
rect 1327 1859 1328 1863
rect 1322 1858 1328 1859
rect 1482 1863 1488 1864
rect 1482 1859 1483 1863
rect 1487 1859 1488 1863
rect 1482 1858 1488 1859
rect 1642 1863 1648 1864
rect 1642 1859 1643 1863
rect 1647 1859 1648 1863
rect 1642 1858 1648 1859
rect 1786 1863 1792 1864
rect 1786 1859 1787 1863
rect 1791 1859 1792 1863
rect 1934 1860 1935 1864
rect 1939 1860 1940 1864
rect 1934 1859 1940 1860
rect 1786 1858 1792 1859
rect 262 1848 268 1849
rect 110 1847 116 1848
rect 110 1843 111 1847
rect 115 1843 116 1847
rect 262 1844 263 1848
rect 267 1844 268 1848
rect 262 1843 268 1844
rect 462 1848 468 1849
rect 462 1844 463 1848
rect 467 1844 468 1848
rect 462 1843 468 1844
rect 654 1848 660 1849
rect 654 1844 655 1848
rect 659 1844 660 1848
rect 654 1843 660 1844
rect 838 1848 844 1849
rect 838 1844 839 1848
rect 843 1844 844 1848
rect 838 1843 844 1844
rect 1014 1848 1020 1849
rect 1014 1844 1015 1848
rect 1019 1844 1020 1848
rect 1014 1843 1020 1844
rect 1182 1848 1188 1849
rect 1182 1844 1183 1848
rect 1187 1844 1188 1848
rect 1182 1843 1188 1844
rect 1350 1848 1356 1849
rect 1350 1844 1351 1848
rect 1355 1844 1356 1848
rect 1350 1843 1356 1844
rect 1510 1848 1516 1849
rect 1510 1844 1511 1848
rect 1515 1844 1516 1848
rect 1510 1843 1516 1844
rect 1670 1848 1676 1849
rect 1670 1844 1671 1848
rect 1675 1844 1676 1848
rect 1670 1843 1676 1844
rect 1814 1848 1820 1849
rect 1814 1844 1815 1848
rect 1819 1844 1820 1848
rect 1814 1843 1820 1844
rect 1934 1847 1940 1848
rect 1934 1843 1935 1847
rect 1939 1843 1940 1847
rect 110 1842 116 1843
rect 1934 1842 1940 1843
rect 3838 1813 3844 1814
rect 5662 1813 5668 1814
rect 3838 1809 3839 1813
rect 3843 1809 3844 1813
rect 3838 1808 3844 1809
rect 4406 1812 4412 1813
rect 4406 1808 4407 1812
rect 4411 1808 4412 1812
rect 4406 1807 4412 1808
rect 4542 1812 4548 1813
rect 4542 1808 4543 1812
rect 4547 1808 4548 1812
rect 4542 1807 4548 1808
rect 4678 1812 4684 1813
rect 4678 1808 4679 1812
rect 4683 1808 4684 1812
rect 4678 1807 4684 1808
rect 4814 1812 4820 1813
rect 4814 1808 4815 1812
rect 4819 1808 4820 1812
rect 4814 1807 4820 1808
rect 4950 1812 4956 1813
rect 4950 1808 4951 1812
rect 4955 1808 4956 1812
rect 5662 1809 5663 1813
rect 5667 1809 5668 1813
rect 5662 1808 5668 1809
rect 4950 1807 4956 1808
rect 4378 1797 4384 1798
rect 3838 1796 3844 1797
rect 3838 1792 3839 1796
rect 3843 1792 3844 1796
rect 4378 1793 4379 1797
rect 4383 1793 4384 1797
rect 4378 1792 4384 1793
rect 4514 1797 4520 1798
rect 4514 1793 4515 1797
rect 4519 1793 4520 1797
rect 4514 1792 4520 1793
rect 4650 1797 4656 1798
rect 4650 1793 4651 1797
rect 4655 1793 4656 1797
rect 4650 1792 4656 1793
rect 4786 1797 4792 1798
rect 4786 1793 4787 1797
rect 4791 1793 4792 1797
rect 4786 1792 4792 1793
rect 4922 1797 4928 1798
rect 4922 1793 4923 1797
rect 4927 1793 4928 1797
rect 4922 1792 4928 1793
rect 5662 1796 5668 1797
rect 5662 1792 5663 1796
rect 5667 1792 5668 1796
rect 3838 1791 3844 1792
rect 5662 1791 5668 1792
rect 110 1777 116 1778
rect 1934 1777 1940 1778
rect 110 1773 111 1777
rect 115 1773 116 1777
rect 110 1772 116 1773
rect 222 1776 228 1777
rect 222 1772 223 1776
rect 227 1772 228 1776
rect 222 1771 228 1772
rect 462 1776 468 1777
rect 462 1772 463 1776
rect 467 1772 468 1776
rect 462 1771 468 1772
rect 694 1776 700 1777
rect 694 1772 695 1776
rect 699 1772 700 1776
rect 694 1771 700 1772
rect 926 1776 932 1777
rect 926 1772 927 1776
rect 931 1772 932 1776
rect 926 1771 932 1772
rect 1158 1776 1164 1777
rect 1158 1772 1159 1776
rect 1163 1772 1164 1776
rect 1158 1771 1164 1772
rect 1390 1776 1396 1777
rect 1390 1772 1391 1776
rect 1395 1772 1396 1776
rect 1934 1773 1935 1777
rect 1939 1773 1940 1777
rect 1934 1772 1940 1773
rect 1390 1771 1396 1772
rect 194 1761 200 1762
rect 110 1760 116 1761
rect 110 1756 111 1760
rect 115 1756 116 1760
rect 194 1757 195 1761
rect 199 1757 200 1761
rect 194 1756 200 1757
rect 434 1761 440 1762
rect 434 1757 435 1761
rect 439 1757 440 1761
rect 434 1756 440 1757
rect 666 1761 672 1762
rect 666 1757 667 1761
rect 671 1757 672 1761
rect 666 1756 672 1757
rect 898 1761 904 1762
rect 898 1757 899 1761
rect 903 1757 904 1761
rect 898 1756 904 1757
rect 1130 1761 1136 1762
rect 1130 1757 1131 1761
rect 1135 1757 1136 1761
rect 1130 1756 1136 1757
rect 1362 1761 1368 1762
rect 1362 1757 1363 1761
rect 1367 1757 1368 1761
rect 1362 1756 1368 1757
rect 1934 1760 1940 1761
rect 1934 1756 1935 1760
rect 1939 1756 1940 1760
rect 110 1755 116 1756
rect 1934 1755 1940 1756
rect 1974 1740 1980 1741
rect 3798 1740 3804 1741
rect 1974 1736 1975 1740
rect 1979 1736 1980 1740
rect 1974 1735 1980 1736
rect 1994 1739 2000 1740
rect 1994 1735 1995 1739
rect 1999 1735 2000 1739
rect 1994 1734 2000 1735
rect 2130 1739 2136 1740
rect 2130 1735 2131 1739
rect 2135 1735 2136 1739
rect 2130 1734 2136 1735
rect 2266 1739 2272 1740
rect 2266 1735 2267 1739
rect 2271 1735 2272 1739
rect 2266 1734 2272 1735
rect 2418 1739 2424 1740
rect 2418 1735 2419 1739
rect 2423 1735 2424 1739
rect 2418 1734 2424 1735
rect 2578 1739 2584 1740
rect 2578 1735 2579 1739
rect 2583 1735 2584 1739
rect 2578 1734 2584 1735
rect 2738 1739 2744 1740
rect 2738 1735 2739 1739
rect 2743 1735 2744 1739
rect 2738 1734 2744 1735
rect 2898 1739 2904 1740
rect 2898 1735 2899 1739
rect 2903 1735 2904 1739
rect 2898 1734 2904 1735
rect 3050 1739 3056 1740
rect 3050 1735 3051 1739
rect 3055 1735 3056 1739
rect 3050 1734 3056 1735
rect 3202 1739 3208 1740
rect 3202 1735 3203 1739
rect 3207 1735 3208 1739
rect 3202 1734 3208 1735
rect 3354 1739 3360 1740
rect 3354 1735 3355 1739
rect 3359 1735 3360 1739
rect 3354 1734 3360 1735
rect 3514 1739 3520 1740
rect 3514 1735 3515 1739
rect 3519 1735 3520 1739
rect 3514 1734 3520 1735
rect 3650 1739 3656 1740
rect 3650 1735 3651 1739
rect 3655 1735 3656 1739
rect 3798 1736 3799 1740
rect 3803 1736 3804 1740
rect 3798 1735 3804 1736
rect 3650 1734 3656 1735
rect 2022 1724 2028 1725
rect 1974 1723 1980 1724
rect 1974 1719 1975 1723
rect 1979 1719 1980 1723
rect 2022 1720 2023 1724
rect 2027 1720 2028 1724
rect 2022 1719 2028 1720
rect 2158 1724 2164 1725
rect 2158 1720 2159 1724
rect 2163 1720 2164 1724
rect 2158 1719 2164 1720
rect 2294 1724 2300 1725
rect 2294 1720 2295 1724
rect 2299 1720 2300 1724
rect 2294 1719 2300 1720
rect 2446 1724 2452 1725
rect 2446 1720 2447 1724
rect 2451 1720 2452 1724
rect 2446 1719 2452 1720
rect 2606 1724 2612 1725
rect 2606 1720 2607 1724
rect 2611 1720 2612 1724
rect 2606 1719 2612 1720
rect 2766 1724 2772 1725
rect 2766 1720 2767 1724
rect 2771 1720 2772 1724
rect 2766 1719 2772 1720
rect 2926 1724 2932 1725
rect 2926 1720 2927 1724
rect 2931 1720 2932 1724
rect 2926 1719 2932 1720
rect 3078 1724 3084 1725
rect 3078 1720 3079 1724
rect 3083 1720 3084 1724
rect 3078 1719 3084 1720
rect 3230 1724 3236 1725
rect 3230 1720 3231 1724
rect 3235 1720 3236 1724
rect 3230 1719 3236 1720
rect 3382 1724 3388 1725
rect 3382 1720 3383 1724
rect 3387 1720 3388 1724
rect 3382 1719 3388 1720
rect 3542 1724 3548 1725
rect 3542 1720 3543 1724
rect 3547 1720 3548 1724
rect 3542 1719 3548 1720
rect 3678 1724 3684 1725
rect 3678 1720 3679 1724
rect 3683 1720 3684 1724
rect 3678 1719 3684 1720
rect 3798 1723 3804 1724
rect 3798 1719 3799 1723
rect 3803 1719 3804 1723
rect 1974 1718 1980 1719
rect 3798 1718 3804 1719
rect 1974 1653 1980 1654
rect 3798 1653 3804 1654
rect 1974 1649 1975 1653
rect 1979 1649 1980 1653
rect 1974 1648 1980 1649
rect 2022 1652 2028 1653
rect 2022 1648 2023 1652
rect 2027 1648 2028 1652
rect 2022 1647 2028 1648
rect 2166 1652 2172 1653
rect 2166 1648 2167 1652
rect 2171 1648 2172 1652
rect 2166 1647 2172 1648
rect 2318 1652 2324 1653
rect 2318 1648 2319 1652
rect 2323 1648 2324 1652
rect 2318 1647 2324 1648
rect 2478 1652 2484 1653
rect 2478 1648 2479 1652
rect 2483 1648 2484 1652
rect 2478 1647 2484 1648
rect 2638 1652 2644 1653
rect 2638 1648 2639 1652
rect 2643 1648 2644 1652
rect 2638 1647 2644 1648
rect 2790 1652 2796 1653
rect 2790 1648 2791 1652
rect 2795 1648 2796 1652
rect 2790 1647 2796 1648
rect 2942 1652 2948 1653
rect 2942 1648 2943 1652
rect 2947 1648 2948 1652
rect 2942 1647 2948 1648
rect 3102 1652 3108 1653
rect 3102 1648 3103 1652
rect 3107 1648 3108 1652
rect 3102 1647 3108 1648
rect 3262 1652 3268 1653
rect 3262 1648 3263 1652
rect 3267 1648 3268 1652
rect 3262 1647 3268 1648
rect 3422 1652 3428 1653
rect 3422 1648 3423 1652
rect 3427 1648 3428 1652
rect 3798 1649 3799 1653
rect 3803 1649 3804 1653
rect 3798 1648 3804 1649
rect 3838 1648 3844 1649
rect 5662 1648 5668 1649
rect 3422 1647 3428 1648
rect 3838 1644 3839 1648
rect 3843 1644 3844 1648
rect 3838 1643 3844 1644
rect 4562 1647 4568 1648
rect 4562 1643 4563 1647
rect 4567 1643 4568 1647
rect 4562 1642 4568 1643
rect 4698 1647 4704 1648
rect 4698 1643 4699 1647
rect 4703 1643 4704 1647
rect 4698 1642 4704 1643
rect 4834 1647 4840 1648
rect 4834 1643 4835 1647
rect 4839 1643 4840 1647
rect 4834 1642 4840 1643
rect 4970 1647 4976 1648
rect 4970 1643 4971 1647
rect 4975 1643 4976 1647
rect 4970 1642 4976 1643
rect 5106 1647 5112 1648
rect 5106 1643 5107 1647
rect 5111 1643 5112 1647
rect 5106 1642 5112 1643
rect 5242 1647 5248 1648
rect 5242 1643 5243 1647
rect 5247 1643 5248 1647
rect 5242 1642 5248 1643
rect 5378 1647 5384 1648
rect 5378 1643 5379 1647
rect 5383 1643 5384 1647
rect 5378 1642 5384 1643
rect 5514 1647 5520 1648
rect 5514 1643 5515 1647
rect 5519 1643 5520 1647
rect 5662 1644 5663 1648
rect 5667 1644 5668 1648
rect 5662 1643 5668 1644
rect 5514 1642 5520 1643
rect 1994 1637 2000 1638
rect 1974 1636 1980 1637
rect 1974 1632 1975 1636
rect 1979 1632 1980 1636
rect 1994 1633 1995 1637
rect 1999 1633 2000 1637
rect 1994 1632 2000 1633
rect 2138 1637 2144 1638
rect 2138 1633 2139 1637
rect 2143 1633 2144 1637
rect 2138 1632 2144 1633
rect 2290 1637 2296 1638
rect 2290 1633 2291 1637
rect 2295 1633 2296 1637
rect 2290 1632 2296 1633
rect 2450 1637 2456 1638
rect 2450 1633 2451 1637
rect 2455 1633 2456 1637
rect 2450 1632 2456 1633
rect 2610 1637 2616 1638
rect 2610 1633 2611 1637
rect 2615 1633 2616 1637
rect 2610 1632 2616 1633
rect 2762 1637 2768 1638
rect 2762 1633 2763 1637
rect 2767 1633 2768 1637
rect 2762 1632 2768 1633
rect 2914 1637 2920 1638
rect 2914 1633 2915 1637
rect 2919 1633 2920 1637
rect 2914 1632 2920 1633
rect 3074 1637 3080 1638
rect 3074 1633 3075 1637
rect 3079 1633 3080 1637
rect 3074 1632 3080 1633
rect 3234 1637 3240 1638
rect 3234 1633 3235 1637
rect 3239 1633 3240 1637
rect 3234 1632 3240 1633
rect 3394 1637 3400 1638
rect 3394 1633 3395 1637
rect 3399 1633 3400 1637
rect 3394 1632 3400 1633
rect 3798 1636 3804 1637
rect 3798 1632 3799 1636
rect 3803 1632 3804 1636
rect 4590 1632 4596 1633
rect 1974 1631 1980 1632
rect 3798 1631 3804 1632
rect 3838 1631 3844 1632
rect 3838 1627 3839 1631
rect 3843 1627 3844 1631
rect 4590 1628 4591 1632
rect 4595 1628 4596 1632
rect 4590 1627 4596 1628
rect 4726 1632 4732 1633
rect 4726 1628 4727 1632
rect 4731 1628 4732 1632
rect 4726 1627 4732 1628
rect 4862 1632 4868 1633
rect 4862 1628 4863 1632
rect 4867 1628 4868 1632
rect 4862 1627 4868 1628
rect 4998 1632 5004 1633
rect 4998 1628 4999 1632
rect 5003 1628 5004 1632
rect 4998 1627 5004 1628
rect 5134 1632 5140 1633
rect 5134 1628 5135 1632
rect 5139 1628 5140 1632
rect 5134 1627 5140 1628
rect 5270 1632 5276 1633
rect 5270 1628 5271 1632
rect 5275 1628 5276 1632
rect 5270 1627 5276 1628
rect 5406 1632 5412 1633
rect 5406 1628 5407 1632
rect 5411 1628 5412 1632
rect 5406 1627 5412 1628
rect 5542 1632 5548 1633
rect 5542 1628 5543 1632
rect 5547 1628 5548 1632
rect 5542 1627 5548 1628
rect 5662 1631 5668 1632
rect 5662 1627 5663 1631
rect 5667 1627 5668 1631
rect 3838 1626 3844 1627
rect 5662 1626 5668 1627
rect 110 1616 116 1617
rect 1934 1616 1940 1617
rect 110 1612 111 1616
rect 115 1612 116 1616
rect 110 1611 116 1612
rect 130 1615 136 1616
rect 130 1611 131 1615
rect 135 1611 136 1615
rect 130 1610 136 1611
rect 362 1615 368 1616
rect 362 1611 363 1615
rect 367 1611 368 1615
rect 362 1610 368 1611
rect 618 1615 624 1616
rect 618 1611 619 1615
rect 623 1611 624 1615
rect 618 1610 624 1611
rect 874 1615 880 1616
rect 874 1611 875 1615
rect 879 1611 880 1615
rect 874 1610 880 1611
rect 1138 1615 1144 1616
rect 1138 1611 1139 1615
rect 1143 1611 1144 1615
rect 1934 1612 1935 1616
rect 1939 1612 1940 1616
rect 1934 1611 1940 1612
rect 1138 1610 1144 1611
rect 158 1600 164 1601
rect 110 1599 116 1600
rect 110 1595 111 1599
rect 115 1595 116 1599
rect 158 1596 159 1600
rect 163 1596 164 1600
rect 158 1595 164 1596
rect 390 1600 396 1601
rect 390 1596 391 1600
rect 395 1596 396 1600
rect 390 1595 396 1596
rect 646 1600 652 1601
rect 646 1596 647 1600
rect 651 1596 652 1600
rect 646 1595 652 1596
rect 902 1600 908 1601
rect 902 1596 903 1600
rect 907 1596 908 1600
rect 902 1595 908 1596
rect 1166 1600 1172 1601
rect 1166 1596 1167 1600
rect 1171 1596 1172 1600
rect 1166 1595 1172 1596
rect 1934 1599 1940 1600
rect 1934 1595 1935 1599
rect 1939 1595 1940 1599
rect 110 1594 116 1595
rect 1934 1594 1940 1595
rect 3838 1557 3844 1558
rect 5662 1557 5668 1558
rect 3838 1553 3839 1557
rect 3843 1553 3844 1557
rect 3838 1552 3844 1553
rect 4590 1556 4596 1557
rect 4590 1552 4591 1556
rect 4595 1552 4596 1556
rect 4590 1551 4596 1552
rect 4726 1556 4732 1557
rect 4726 1552 4727 1556
rect 4731 1552 4732 1556
rect 4726 1551 4732 1552
rect 4862 1556 4868 1557
rect 4862 1552 4863 1556
rect 4867 1552 4868 1556
rect 4862 1551 4868 1552
rect 4998 1556 5004 1557
rect 4998 1552 4999 1556
rect 5003 1552 5004 1556
rect 4998 1551 5004 1552
rect 5134 1556 5140 1557
rect 5134 1552 5135 1556
rect 5139 1552 5140 1556
rect 5134 1551 5140 1552
rect 5270 1556 5276 1557
rect 5270 1552 5271 1556
rect 5275 1552 5276 1556
rect 5270 1551 5276 1552
rect 5406 1556 5412 1557
rect 5406 1552 5407 1556
rect 5411 1552 5412 1556
rect 5406 1551 5412 1552
rect 5542 1556 5548 1557
rect 5542 1552 5543 1556
rect 5547 1552 5548 1556
rect 5662 1553 5663 1557
rect 5667 1553 5668 1557
rect 5662 1552 5668 1553
rect 5542 1551 5548 1552
rect 4562 1541 4568 1542
rect 3838 1540 3844 1541
rect 3838 1536 3839 1540
rect 3843 1536 3844 1540
rect 4562 1537 4563 1541
rect 4567 1537 4568 1541
rect 4562 1536 4568 1537
rect 4698 1541 4704 1542
rect 4698 1537 4699 1541
rect 4703 1537 4704 1541
rect 4698 1536 4704 1537
rect 4834 1541 4840 1542
rect 4834 1537 4835 1541
rect 4839 1537 4840 1541
rect 4834 1536 4840 1537
rect 4970 1541 4976 1542
rect 4970 1537 4971 1541
rect 4975 1537 4976 1541
rect 4970 1536 4976 1537
rect 5106 1541 5112 1542
rect 5106 1537 5107 1541
rect 5111 1537 5112 1541
rect 5106 1536 5112 1537
rect 5242 1541 5248 1542
rect 5242 1537 5243 1541
rect 5247 1537 5248 1541
rect 5242 1536 5248 1537
rect 5378 1541 5384 1542
rect 5378 1537 5379 1541
rect 5383 1537 5384 1541
rect 5378 1536 5384 1537
rect 5514 1541 5520 1542
rect 5514 1537 5515 1541
rect 5519 1537 5520 1541
rect 5514 1536 5520 1537
rect 5662 1540 5668 1541
rect 5662 1536 5663 1540
rect 5667 1536 5668 1540
rect 3838 1535 3844 1536
rect 5662 1535 5668 1536
rect 110 1529 116 1530
rect 1934 1529 1940 1530
rect 110 1525 111 1529
rect 115 1525 116 1529
rect 110 1524 116 1525
rect 158 1528 164 1529
rect 158 1524 159 1528
rect 163 1524 164 1528
rect 158 1523 164 1524
rect 326 1528 332 1529
rect 326 1524 327 1528
rect 331 1524 332 1528
rect 326 1523 332 1524
rect 510 1528 516 1529
rect 510 1524 511 1528
rect 515 1524 516 1528
rect 510 1523 516 1524
rect 694 1528 700 1529
rect 694 1524 695 1528
rect 699 1524 700 1528
rect 694 1523 700 1524
rect 886 1528 892 1529
rect 886 1524 887 1528
rect 891 1524 892 1528
rect 886 1523 892 1524
rect 1078 1528 1084 1529
rect 1078 1524 1079 1528
rect 1083 1524 1084 1528
rect 1934 1525 1935 1529
rect 1939 1525 1940 1529
rect 1934 1524 1940 1525
rect 1078 1523 1084 1524
rect 130 1513 136 1514
rect 110 1512 116 1513
rect 110 1508 111 1512
rect 115 1508 116 1512
rect 130 1509 131 1513
rect 135 1509 136 1513
rect 130 1508 136 1509
rect 298 1513 304 1514
rect 298 1509 299 1513
rect 303 1509 304 1513
rect 298 1508 304 1509
rect 482 1513 488 1514
rect 482 1509 483 1513
rect 487 1509 488 1513
rect 482 1508 488 1509
rect 666 1513 672 1514
rect 666 1509 667 1513
rect 671 1509 672 1513
rect 666 1508 672 1509
rect 858 1513 864 1514
rect 858 1509 859 1513
rect 863 1509 864 1513
rect 858 1508 864 1509
rect 1050 1513 1056 1514
rect 1050 1509 1051 1513
rect 1055 1509 1056 1513
rect 1050 1508 1056 1509
rect 1934 1512 1940 1513
rect 1934 1508 1935 1512
rect 1939 1508 1940 1512
rect 110 1507 116 1508
rect 1934 1507 1940 1508
rect 1974 1492 1980 1493
rect 3798 1492 3804 1493
rect 1974 1488 1975 1492
rect 1979 1488 1980 1492
rect 1974 1487 1980 1488
rect 1994 1491 2000 1492
rect 1994 1487 1995 1491
rect 1999 1487 2000 1491
rect 1994 1486 2000 1487
rect 2130 1491 2136 1492
rect 2130 1487 2131 1491
rect 2135 1487 2136 1491
rect 2130 1486 2136 1487
rect 2266 1491 2272 1492
rect 2266 1487 2267 1491
rect 2271 1487 2272 1491
rect 2266 1486 2272 1487
rect 2402 1491 2408 1492
rect 2402 1487 2403 1491
rect 2407 1487 2408 1491
rect 2402 1486 2408 1487
rect 2538 1491 2544 1492
rect 2538 1487 2539 1491
rect 2543 1487 2544 1491
rect 2538 1486 2544 1487
rect 2674 1491 2680 1492
rect 2674 1487 2675 1491
rect 2679 1487 2680 1491
rect 2674 1486 2680 1487
rect 2810 1491 2816 1492
rect 2810 1487 2811 1491
rect 2815 1487 2816 1491
rect 2810 1486 2816 1487
rect 2946 1491 2952 1492
rect 2946 1487 2947 1491
rect 2951 1487 2952 1491
rect 2946 1486 2952 1487
rect 3082 1491 3088 1492
rect 3082 1487 3083 1491
rect 3087 1487 3088 1491
rect 3082 1486 3088 1487
rect 3218 1491 3224 1492
rect 3218 1487 3219 1491
rect 3223 1487 3224 1491
rect 3218 1486 3224 1487
rect 3354 1491 3360 1492
rect 3354 1487 3355 1491
rect 3359 1487 3360 1491
rect 3354 1486 3360 1487
rect 3490 1491 3496 1492
rect 3490 1487 3491 1491
rect 3495 1487 3496 1491
rect 3798 1488 3799 1492
rect 3803 1488 3804 1492
rect 3798 1487 3804 1488
rect 3490 1486 3496 1487
rect 2022 1476 2028 1477
rect 1974 1475 1980 1476
rect 1974 1471 1975 1475
rect 1979 1471 1980 1475
rect 2022 1472 2023 1476
rect 2027 1472 2028 1476
rect 2022 1471 2028 1472
rect 2158 1476 2164 1477
rect 2158 1472 2159 1476
rect 2163 1472 2164 1476
rect 2158 1471 2164 1472
rect 2294 1476 2300 1477
rect 2294 1472 2295 1476
rect 2299 1472 2300 1476
rect 2294 1471 2300 1472
rect 2430 1476 2436 1477
rect 2430 1472 2431 1476
rect 2435 1472 2436 1476
rect 2430 1471 2436 1472
rect 2566 1476 2572 1477
rect 2566 1472 2567 1476
rect 2571 1472 2572 1476
rect 2566 1471 2572 1472
rect 2702 1476 2708 1477
rect 2702 1472 2703 1476
rect 2707 1472 2708 1476
rect 2702 1471 2708 1472
rect 2838 1476 2844 1477
rect 2838 1472 2839 1476
rect 2843 1472 2844 1476
rect 2838 1471 2844 1472
rect 2974 1476 2980 1477
rect 2974 1472 2975 1476
rect 2979 1472 2980 1476
rect 2974 1471 2980 1472
rect 3110 1476 3116 1477
rect 3110 1472 3111 1476
rect 3115 1472 3116 1476
rect 3110 1471 3116 1472
rect 3246 1476 3252 1477
rect 3246 1472 3247 1476
rect 3251 1472 3252 1476
rect 3246 1471 3252 1472
rect 3382 1476 3388 1477
rect 3382 1472 3383 1476
rect 3387 1472 3388 1476
rect 3382 1471 3388 1472
rect 3518 1476 3524 1477
rect 3518 1472 3519 1476
rect 3523 1472 3524 1476
rect 3518 1471 3524 1472
rect 3798 1475 3804 1476
rect 3798 1471 3799 1475
rect 3803 1471 3804 1475
rect 1974 1470 1980 1471
rect 3798 1470 3804 1471
rect 1974 1405 1980 1406
rect 3798 1405 3804 1406
rect 1974 1401 1975 1405
rect 1979 1401 1980 1405
rect 1974 1400 1980 1401
rect 2166 1404 2172 1405
rect 2166 1400 2167 1404
rect 2171 1400 2172 1404
rect 2166 1399 2172 1400
rect 2302 1404 2308 1405
rect 2302 1400 2303 1404
rect 2307 1400 2308 1404
rect 2302 1399 2308 1400
rect 2438 1404 2444 1405
rect 2438 1400 2439 1404
rect 2443 1400 2444 1404
rect 2438 1399 2444 1400
rect 2574 1404 2580 1405
rect 2574 1400 2575 1404
rect 2579 1400 2580 1404
rect 2574 1399 2580 1400
rect 2710 1404 2716 1405
rect 2710 1400 2711 1404
rect 2715 1400 2716 1404
rect 2710 1399 2716 1400
rect 2846 1404 2852 1405
rect 2846 1400 2847 1404
rect 2851 1400 2852 1404
rect 2846 1399 2852 1400
rect 2982 1404 2988 1405
rect 2982 1400 2983 1404
rect 2987 1400 2988 1404
rect 2982 1399 2988 1400
rect 3118 1404 3124 1405
rect 3118 1400 3119 1404
rect 3123 1400 3124 1404
rect 3118 1399 3124 1400
rect 3254 1404 3260 1405
rect 3254 1400 3255 1404
rect 3259 1400 3260 1404
rect 3798 1401 3799 1405
rect 3803 1401 3804 1405
rect 3798 1400 3804 1401
rect 3254 1399 3260 1400
rect 2138 1389 2144 1390
rect 1974 1388 1980 1389
rect 1974 1384 1975 1388
rect 1979 1384 1980 1388
rect 2138 1385 2139 1389
rect 2143 1385 2144 1389
rect 2138 1384 2144 1385
rect 2274 1389 2280 1390
rect 2274 1385 2275 1389
rect 2279 1385 2280 1389
rect 2274 1384 2280 1385
rect 2410 1389 2416 1390
rect 2410 1385 2411 1389
rect 2415 1385 2416 1389
rect 2410 1384 2416 1385
rect 2546 1389 2552 1390
rect 2546 1385 2547 1389
rect 2551 1385 2552 1389
rect 2546 1384 2552 1385
rect 2682 1389 2688 1390
rect 2682 1385 2683 1389
rect 2687 1385 2688 1389
rect 2682 1384 2688 1385
rect 2818 1389 2824 1390
rect 2818 1385 2819 1389
rect 2823 1385 2824 1389
rect 2818 1384 2824 1385
rect 2954 1389 2960 1390
rect 2954 1385 2955 1389
rect 2959 1385 2960 1389
rect 2954 1384 2960 1385
rect 3090 1389 3096 1390
rect 3090 1385 3091 1389
rect 3095 1385 3096 1389
rect 3090 1384 3096 1385
rect 3226 1389 3232 1390
rect 3226 1385 3227 1389
rect 3231 1385 3232 1389
rect 3226 1384 3232 1385
rect 3798 1388 3804 1389
rect 3798 1384 3799 1388
rect 3803 1384 3804 1388
rect 1974 1383 1980 1384
rect 3798 1383 3804 1384
rect 110 1368 116 1369
rect 1934 1368 1940 1369
rect 110 1364 111 1368
rect 115 1364 116 1368
rect 110 1363 116 1364
rect 130 1367 136 1368
rect 130 1363 131 1367
rect 135 1363 136 1367
rect 130 1362 136 1363
rect 394 1367 400 1368
rect 394 1363 395 1367
rect 399 1363 400 1367
rect 394 1362 400 1363
rect 682 1367 688 1368
rect 682 1363 683 1367
rect 687 1363 688 1367
rect 682 1362 688 1363
rect 970 1367 976 1368
rect 970 1363 971 1367
rect 975 1363 976 1367
rect 970 1362 976 1363
rect 1258 1367 1264 1368
rect 1258 1363 1259 1367
rect 1263 1363 1264 1367
rect 1934 1364 1935 1368
rect 1939 1364 1940 1368
rect 1934 1363 1940 1364
rect 1258 1362 1264 1363
rect 158 1352 164 1353
rect 110 1351 116 1352
rect 110 1347 111 1351
rect 115 1347 116 1351
rect 158 1348 159 1352
rect 163 1348 164 1352
rect 158 1347 164 1348
rect 422 1352 428 1353
rect 422 1348 423 1352
rect 427 1348 428 1352
rect 422 1347 428 1348
rect 710 1352 716 1353
rect 710 1348 711 1352
rect 715 1348 716 1352
rect 710 1347 716 1348
rect 998 1352 1004 1353
rect 998 1348 999 1352
rect 1003 1348 1004 1352
rect 998 1347 1004 1348
rect 1286 1352 1292 1353
rect 1286 1348 1287 1352
rect 1291 1348 1292 1352
rect 1286 1347 1292 1348
rect 1934 1351 1940 1352
rect 1934 1347 1935 1351
rect 1939 1347 1940 1351
rect 110 1346 116 1347
rect 1934 1346 1940 1347
rect 3838 1336 3844 1337
rect 5662 1336 5668 1337
rect 3838 1332 3839 1336
rect 3843 1332 3844 1336
rect 3838 1331 3844 1332
rect 4810 1335 4816 1336
rect 4810 1331 4811 1335
rect 4815 1331 4816 1335
rect 4810 1330 4816 1331
rect 4946 1335 4952 1336
rect 4946 1331 4947 1335
rect 4951 1331 4952 1335
rect 4946 1330 4952 1331
rect 5082 1335 5088 1336
rect 5082 1331 5083 1335
rect 5087 1331 5088 1335
rect 5082 1330 5088 1331
rect 5218 1335 5224 1336
rect 5218 1331 5219 1335
rect 5223 1331 5224 1335
rect 5218 1330 5224 1331
rect 5354 1335 5360 1336
rect 5354 1331 5355 1335
rect 5359 1331 5360 1335
rect 5354 1330 5360 1331
rect 5490 1335 5496 1336
rect 5490 1331 5491 1335
rect 5495 1331 5496 1335
rect 5662 1332 5663 1336
rect 5667 1332 5668 1336
rect 5662 1331 5668 1332
rect 5490 1330 5496 1331
rect 4838 1320 4844 1321
rect 3838 1319 3844 1320
rect 3838 1315 3839 1319
rect 3843 1315 3844 1319
rect 4838 1316 4839 1320
rect 4843 1316 4844 1320
rect 4838 1315 4844 1316
rect 4974 1320 4980 1321
rect 4974 1316 4975 1320
rect 4979 1316 4980 1320
rect 4974 1315 4980 1316
rect 5110 1320 5116 1321
rect 5110 1316 5111 1320
rect 5115 1316 5116 1320
rect 5110 1315 5116 1316
rect 5246 1320 5252 1321
rect 5246 1316 5247 1320
rect 5251 1316 5252 1320
rect 5246 1315 5252 1316
rect 5382 1320 5388 1321
rect 5382 1316 5383 1320
rect 5387 1316 5388 1320
rect 5382 1315 5388 1316
rect 5518 1320 5524 1321
rect 5518 1316 5519 1320
rect 5523 1316 5524 1320
rect 5518 1315 5524 1316
rect 5662 1319 5668 1320
rect 5662 1315 5663 1319
rect 5667 1315 5668 1319
rect 3838 1314 3844 1315
rect 5662 1314 5668 1315
rect 110 1293 116 1294
rect 1934 1293 1940 1294
rect 110 1289 111 1293
rect 115 1289 116 1293
rect 110 1288 116 1289
rect 158 1292 164 1293
rect 158 1288 159 1292
rect 163 1288 164 1292
rect 158 1287 164 1288
rect 454 1292 460 1293
rect 454 1288 455 1292
rect 459 1288 460 1292
rect 454 1287 460 1288
rect 774 1292 780 1293
rect 774 1288 775 1292
rect 779 1288 780 1292
rect 774 1287 780 1288
rect 1094 1292 1100 1293
rect 1094 1288 1095 1292
rect 1099 1288 1100 1292
rect 1094 1287 1100 1288
rect 1422 1292 1428 1293
rect 1422 1288 1423 1292
rect 1427 1288 1428 1292
rect 1934 1289 1935 1293
rect 1939 1289 1940 1293
rect 1934 1288 1940 1289
rect 1422 1287 1428 1288
rect 130 1277 136 1278
rect 110 1276 116 1277
rect 110 1272 111 1276
rect 115 1272 116 1276
rect 130 1273 131 1277
rect 135 1273 136 1277
rect 130 1272 136 1273
rect 426 1277 432 1278
rect 426 1273 427 1277
rect 431 1273 432 1277
rect 426 1272 432 1273
rect 746 1277 752 1278
rect 746 1273 747 1277
rect 751 1273 752 1277
rect 746 1272 752 1273
rect 1066 1277 1072 1278
rect 1066 1273 1067 1277
rect 1071 1273 1072 1277
rect 1066 1272 1072 1273
rect 1394 1277 1400 1278
rect 1394 1273 1395 1277
rect 1399 1273 1400 1277
rect 1394 1272 1400 1273
rect 1934 1276 1940 1277
rect 1934 1272 1935 1276
rect 1939 1272 1940 1276
rect 110 1271 116 1272
rect 1934 1271 1940 1272
rect 3838 1257 3844 1258
rect 5662 1257 5668 1258
rect 1974 1256 1980 1257
rect 3798 1256 3804 1257
rect 1974 1252 1975 1256
rect 1979 1252 1980 1256
rect 1974 1251 1980 1252
rect 2130 1255 2136 1256
rect 2130 1251 2131 1255
rect 2135 1251 2136 1255
rect 2130 1250 2136 1251
rect 2266 1255 2272 1256
rect 2266 1251 2267 1255
rect 2271 1251 2272 1255
rect 2266 1250 2272 1251
rect 2402 1255 2408 1256
rect 2402 1251 2403 1255
rect 2407 1251 2408 1255
rect 2402 1250 2408 1251
rect 2554 1255 2560 1256
rect 2554 1251 2555 1255
rect 2559 1251 2560 1255
rect 2554 1250 2560 1251
rect 2714 1255 2720 1256
rect 2714 1251 2715 1255
rect 2719 1251 2720 1255
rect 2714 1250 2720 1251
rect 2890 1255 2896 1256
rect 2890 1251 2891 1255
rect 2895 1251 2896 1255
rect 2890 1250 2896 1251
rect 3074 1255 3080 1256
rect 3074 1251 3075 1255
rect 3079 1251 3080 1255
rect 3074 1250 3080 1251
rect 3266 1255 3272 1256
rect 3266 1251 3267 1255
rect 3271 1251 3272 1255
rect 3266 1250 3272 1251
rect 3466 1255 3472 1256
rect 3466 1251 3467 1255
rect 3471 1251 3472 1255
rect 3466 1250 3472 1251
rect 3650 1255 3656 1256
rect 3650 1251 3651 1255
rect 3655 1251 3656 1255
rect 3798 1252 3799 1256
rect 3803 1252 3804 1256
rect 3838 1253 3839 1257
rect 3843 1253 3844 1257
rect 3838 1252 3844 1253
rect 4734 1256 4740 1257
rect 4734 1252 4735 1256
rect 4739 1252 4740 1256
rect 3798 1251 3804 1252
rect 4734 1251 4740 1252
rect 4878 1256 4884 1257
rect 4878 1252 4879 1256
rect 4883 1252 4884 1256
rect 4878 1251 4884 1252
rect 5030 1256 5036 1257
rect 5030 1252 5031 1256
rect 5035 1252 5036 1256
rect 5030 1251 5036 1252
rect 5190 1256 5196 1257
rect 5190 1252 5191 1256
rect 5195 1252 5196 1256
rect 5190 1251 5196 1252
rect 5358 1256 5364 1257
rect 5358 1252 5359 1256
rect 5363 1252 5364 1256
rect 5358 1251 5364 1252
rect 5526 1256 5532 1257
rect 5526 1252 5527 1256
rect 5531 1252 5532 1256
rect 5662 1253 5663 1257
rect 5667 1253 5668 1257
rect 5662 1252 5668 1253
rect 5526 1251 5532 1252
rect 3650 1250 3656 1251
rect 4706 1241 4712 1242
rect 2158 1240 2164 1241
rect 1974 1239 1980 1240
rect 1974 1235 1975 1239
rect 1979 1235 1980 1239
rect 2158 1236 2159 1240
rect 2163 1236 2164 1240
rect 2158 1235 2164 1236
rect 2294 1240 2300 1241
rect 2294 1236 2295 1240
rect 2299 1236 2300 1240
rect 2294 1235 2300 1236
rect 2430 1240 2436 1241
rect 2430 1236 2431 1240
rect 2435 1236 2436 1240
rect 2430 1235 2436 1236
rect 2582 1240 2588 1241
rect 2582 1236 2583 1240
rect 2587 1236 2588 1240
rect 2582 1235 2588 1236
rect 2742 1240 2748 1241
rect 2742 1236 2743 1240
rect 2747 1236 2748 1240
rect 2742 1235 2748 1236
rect 2918 1240 2924 1241
rect 2918 1236 2919 1240
rect 2923 1236 2924 1240
rect 2918 1235 2924 1236
rect 3102 1240 3108 1241
rect 3102 1236 3103 1240
rect 3107 1236 3108 1240
rect 3102 1235 3108 1236
rect 3294 1240 3300 1241
rect 3294 1236 3295 1240
rect 3299 1236 3300 1240
rect 3294 1235 3300 1236
rect 3494 1240 3500 1241
rect 3494 1236 3495 1240
rect 3499 1236 3500 1240
rect 3494 1235 3500 1236
rect 3678 1240 3684 1241
rect 3838 1240 3844 1241
rect 3678 1236 3679 1240
rect 3683 1236 3684 1240
rect 3678 1235 3684 1236
rect 3798 1239 3804 1240
rect 3798 1235 3799 1239
rect 3803 1235 3804 1239
rect 3838 1236 3839 1240
rect 3843 1236 3844 1240
rect 4706 1237 4707 1241
rect 4711 1237 4712 1241
rect 4706 1236 4712 1237
rect 4850 1241 4856 1242
rect 4850 1237 4851 1241
rect 4855 1237 4856 1241
rect 4850 1236 4856 1237
rect 5002 1241 5008 1242
rect 5002 1237 5003 1241
rect 5007 1237 5008 1241
rect 5002 1236 5008 1237
rect 5162 1241 5168 1242
rect 5162 1237 5163 1241
rect 5167 1237 5168 1241
rect 5162 1236 5168 1237
rect 5330 1241 5336 1242
rect 5330 1237 5331 1241
rect 5335 1237 5336 1241
rect 5330 1236 5336 1237
rect 5498 1241 5504 1242
rect 5498 1237 5499 1241
rect 5503 1237 5504 1241
rect 5498 1236 5504 1237
rect 5662 1240 5668 1241
rect 5662 1236 5663 1240
rect 5667 1236 5668 1240
rect 3838 1235 3844 1236
rect 5662 1235 5668 1236
rect 1974 1234 1980 1235
rect 3798 1234 3804 1235
rect 1974 1181 1980 1182
rect 3798 1181 3804 1182
rect 1974 1177 1975 1181
rect 1979 1177 1980 1181
rect 1974 1176 1980 1177
rect 2022 1180 2028 1181
rect 2022 1176 2023 1180
rect 2027 1176 2028 1180
rect 2022 1175 2028 1176
rect 2238 1180 2244 1181
rect 2238 1176 2239 1180
rect 2243 1176 2244 1180
rect 2238 1175 2244 1176
rect 2478 1180 2484 1181
rect 2478 1176 2479 1180
rect 2483 1176 2484 1180
rect 2478 1175 2484 1176
rect 2718 1180 2724 1181
rect 2718 1176 2719 1180
rect 2723 1176 2724 1180
rect 2718 1175 2724 1176
rect 2958 1180 2964 1181
rect 2958 1176 2959 1180
rect 2963 1176 2964 1180
rect 2958 1175 2964 1176
rect 3206 1180 3212 1181
rect 3206 1176 3207 1180
rect 3211 1176 3212 1180
rect 3206 1175 3212 1176
rect 3454 1180 3460 1181
rect 3454 1176 3455 1180
rect 3459 1176 3460 1180
rect 3454 1175 3460 1176
rect 3678 1180 3684 1181
rect 3678 1176 3679 1180
rect 3683 1176 3684 1180
rect 3798 1177 3799 1181
rect 3803 1177 3804 1181
rect 3798 1176 3804 1177
rect 3678 1175 3684 1176
rect 1994 1165 2000 1166
rect 1974 1164 1980 1165
rect 1974 1160 1975 1164
rect 1979 1160 1980 1164
rect 1994 1161 1995 1165
rect 1999 1161 2000 1165
rect 1994 1160 2000 1161
rect 2210 1165 2216 1166
rect 2210 1161 2211 1165
rect 2215 1161 2216 1165
rect 2210 1160 2216 1161
rect 2450 1165 2456 1166
rect 2450 1161 2451 1165
rect 2455 1161 2456 1165
rect 2450 1160 2456 1161
rect 2690 1165 2696 1166
rect 2690 1161 2691 1165
rect 2695 1161 2696 1165
rect 2690 1160 2696 1161
rect 2930 1165 2936 1166
rect 2930 1161 2931 1165
rect 2935 1161 2936 1165
rect 2930 1160 2936 1161
rect 3178 1165 3184 1166
rect 3178 1161 3179 1165
rect 3183 1161 3184 1165
rect 3178 1160 3184 1161
rect 3426 1165 3432 1166
rect 3426 1161 3427 1165
rect 3431 1161 3432 1165
rect 3426 1160 3432 1161
rect 3650 1165 3656 1166
rect 3650 1161 3651 1165
rect 3655 1161 3656 1165
rect 3650 1160 3656 1161
rect 3798 1164 3804 1165
rect 3798 1160 3799 1164
rect 3803 1160 3804 1164
rect 1974 1159 1980 1160
rect 3798 1159 3804 1160
rect 110 1120 116 1121
rect 1934 1120 1940 1121
rect 110 1116 111 1120
rect 115 1116 116 1120
rect 110 1115 116 1116
rect 130 1119 136 1120
rect 130 1115 131 1119
rect 135 1115 136 1119
rect 130 1114 136 1115
rect 330 1119 336 1120
rect 330 1115 331 1119
rect 335 1115 336 1119
rect 330 1114 336 1115
rect 562 1119 568 1120
rect 562 1115 563 1119
rect 567 1115 568 1119
rect 562 1114 568 1115
rect 802 1119 808 1120
rect 802 1115 803 1119
rect 807 1115 808 1119
rect 802 1114 808 1115
rect 1042 1119 1048 1120
rect 1042 1115 1043 1119
rect 1047 1115 1048 1119
rect 1042 1114 1048 1115
rect 1282 1119 1288 1120
rect 1282 1115 1283 1119
rect 1287 1115 1288 1119
rect 1282 1114 1288 1115
rect 1522 1119 1528 1120
rect 1522 1115 1523 1119
rect 1527 1115 1528 1119
rect 1522 1114 1528 1115
rect 1770 1119 1776 1120
rect 1770 1115 1771 1119
rect 1775 1115 1776 1119
rect 1934 1116 1935 1120
rect 1939 1116 1940 1120
rect 1934 1115 1940 1116
rect 1770 1114 1776 1115
rect 158 1104 164 1105
rect 110 1103 116 1104
rect 110 1099 111 1103
rect 115 1099 116 1103
rect 158 1100 159 1104
rect 163 1100 164 1104
rect 158 1099 164 1100
rect 358 1104 364 1105
rect 358 1100 359 1104
rect 363 1100 364 1104
rect 358 1099 364 1100
rect 590 1104 596 1105
rect 590 1100 591 1104
rect 595 1100 596 1104
rect 590 1099 596 1100
rect 830 1104 836 1105
rect 830 1100 831 1104
rect 835 1100 836 1104
rect 830 1099 836 1100
rect 1070 1104 1076 1105
rect 1070 1100 1071 1104
rect 1075 1100 1076 1104
rect 1070 1099 1076 1100
rect 1310 1104 1316 1105
rect 1310 1100 1311 1104
rect 1315 1100 1316 1104
rect 1310 1099 1316 1100
rect 1550 1104 1556 1105
rect 1550 1100 1551 1104
rect 1555 1100 1556 1104
rect 1550 1099 1556 1100
rect 1798 1104 1804 1105
rect 1798 1100 1799 1104
rect 1803 1100 1804 1104
rect 1798 1099 1804 1100
rect 1934 1103 1940 1104
rect 1934 1099 1935 1103
rect 1939 1099 1940 1103
rect 110 1098 116 1099
rect 1934 1098 1940 1099
rect 3838 1100 3844 1101
rect 5662 1100 5668 1101
rect 3838 1096 3839 1100
rect 3843 1096 3844 1100
rect 3838 1095 3844 1096
rect 3858 1099 3864 1100
rect 3858 1095 3859 1099
rect 3863 1095 3864 1099
rect 3858 1094 3864 1095
rect 4066 1099 4072 1100
rect 4066 1095 4067 1099
rect 4071 1095 4072 1099
rect 4066 1094 4072 1095
rect 4298 1099 4304 1100
rect 4298 1095 4299 1099
rect 4303 1095 4304 1099
rect 4298 1094 4304 1095
rect 4538 1099 4544 1100
rect 4538 1095 4539 1099
rect 4543 1095 4544 1099
rect 4538 1094 4544 1095
rect 4778 1099 4784 1100
rect 4778 1095 4779 1099
rect 4783 1095 4784 1099
rect 4778 1094 4784 1095
rect 5026 1099 5032 1100
rect 5026 1095 5027 1099
rect 5031 1095 5032 1099
rect 5026 1094 5032 1095
rect 5282 1099 5288 1100
rect 5282 1095 5283 1099
rect 5287 1095 5288 1099
rect 5282 1094 5288 1095
rect 5514 1099 5520 1100
rect 5514 1095 5515 1099
rect 5519 1095 5520 1099
rect 5662 1096 5663 1100
rect 5667 1096 5668 1100
rect 5662 1095 5668 1096
rect 5514 1094 5520 1095
rect 3886 1084 3892 1085
rect 3838 1083 3844 1084
rect 3838 1079 3839 1083
rect 3843 1079 3844 1083
rect 3886 1080 3887 1084
rect 3891 1080 3892 1084
rect 3886 1079 3892 1080
rect 4094 1084 4100 1085
rect 4094 1080 4095 1084
rect 4099 1080 4100 1084
rect 4094 1079 4100 1080
rect 4326 1084 4332 1085
rect 4326 1080 4327 1084
rect 4331 1080 4332 1084
rect 4326 1079 4332 1080
rect 4566 1084 4572 1085
rect 4566 1080 4567 1084
rect 4571 1080 4572 1084
rect 4566 1079 4572 1080
rect 4806 1084 4812 1085
rect 4806 1080 4807 1084
rect 4811 1080 4812 1084
rect 4806 1079 4812 1080
rect 5054 1084 5060 1085
rect 5054 1080 5055 1084
rect 5059 1080 5060 1084
rect 5054 1079 5060 1080
rect 5310 1084 5316 1085
rect 5310 1080 5311 1084
rect 5315 1080 5316 1084
rect 5310 1079 5316 1080
rect 5542 1084 5548 1085
rect 5542 1080 5543 1084
rect 5547 1080 5548 1084
rect 5542 1079 5548 1080
rect 5662 1083 5668 1084
rect 5662 1079 5663 1083
rect 5667 1079 5668 1083
rect 3838 1078 3844 1079
rect 5662 1078 5668 1079
rect 110 1045 116 1046
rect 1934 1045 1940 1046
rect 110 1041 111 1045
rect 115 1041 116 1045
rect 110 1040 116 1041
rect 262 1044 268 1045
rect 262 1040 263 1044
rect 267 1040 268 1044
rect 262 1039 268 1040
rect 438 1044 444 1045
rect 438 1040 439 1044
rect 443 1040 444 1044
rect 438 1039 444 1040
rect 614 1044 620 1045
rect 614 1040 615 1044
rect 619 1040 620 1044
rect 614 1039 620 1040
rect 782 1044 788 1045
rect 782 1040 783 1044
rect 787 1040 788 1044
rect 782 1039 788 1040
rect 950 1044 956 1045
rect 950 1040 951 1044
rect 955 1040 956 1044
rect 950 1039 956 1040
rect 1110 1044 1116 1045
rect 1110 1040 1111 1044
rect 1115 1040 1116 1044
rect 1110 1039 1116 1040
rect 1270 1044 1276 1045
rect 1270 1040 1271 1044
rect 1275 1040 1276 1044
rect 1270 1039 1276 1040
rect 1430 1044 1436 1045
rect 1430 1040 1431 1044
rect 1435 1040 1436 1044
rect 1430 1039 1436 1040
rect 1590 1044 1596 1045
rect 1590 1040 1591 1044
rect 1595 1040 1596 1044
rect 1590 1039 1596 1040
rect 1750 1044 1756 1045
rect 1750 1040 1751 1044
rect 1755 1040 1756 1044
rect 1934 1041 1935 1045
rect 1939 1041 1940 1045
rect 1934 1040 1940 1041
rect 1750 1039 1756 1040
rect 234 1029 240 1030
rect 110 1028 116 1029
rect 110 1024 111 1028
rect 115 1024 116 1028
rect 234 1025 235 1029
rect 239 1025 240 1029
rect 234 1024 240 1025
rect 410 1029 416 1030
rect 410 1025 411 1029
rect 415 1025 416 1029
rect 410 1024 416 1025
rect 586 1029 592 1030
rect 586 1025 587 1029
rect 591 1025 592 1029
rect 586 1024 592 1025
rect 754 1029 760 1030
rect 754 1025 755 1029
rect 759 1025 760 1029
rect 754 1024 760 1025
rect 922 1029 928 1030
rect 922 1025 923 1029
rect 927 1025 928 1029
rect 922 1024 928 1025
rect 1082 1029 1088 1030
rect 1082 1025 1083 1029
rect 1087 1025 1088 1029
rect 1082 1024 1088 1025
rect 1242 1029 1248 1030
rect 1242 1025 1243 1029
rect 1247 1025 1248 1029
rect 1242 1024 1248 1025
rect 1402 1029 1408 1030
rect 1402 1025 1403 1029
rect 1407 1025 1408 1029
rect 1402 1024 1408 1025
rect 1562 1029 1568 1030
rect 1562 1025 1563 1029
rect 1567 1025 1568 1029
rect 1562 1024 1568 1025
rect 1722 1029 1728 1030
rect 1722 1025 1723 1029
rect 1727 1025 1728 1029
rect 1722 1024 1728 1025
rect 1934 1028 1940 1029
rect 1934 1024 1935 1028
rect 1939 1024 1940 1028
rect 110 1023 116 1024
rect 1934 1023 1940 1024
rect 3838 1025 3844 1026
rect 5662 1025 5668 1026
rect 3838 1021 3839 1025
rect 3843 1021 3844 1025
rect 3838 1020 3844 1021
rect 3886 1024 3892 1025
rect 3886 1020 3887 1024
rect 3891 1020 3892 1024
rect 3886 1019 3892 1020
rect 4070 1024 4076 1025
rect 4070 1020 4071 1024
rect 4075 1020 4076 1024
rect 4070 1019 4076 1020
rect 4278 1024 4284 1025
rect 4278 1020 4279 1024
rect 4283 1020 4284 1024
rect 4278 1019 4284 1020
rect 4510 1024 4516 1025
rect 4510 1020 4511 1024
rect 4515 1020 4516 1024
rect 4510 1019 4516 1020
rect 4758 1024 4764 1025
rect 4758 1020 4759 1024
rect 4763 1020 4764 1024
rect 4758 1019 4764 1020
rect 5022 1024 5028 1025
rect 5022 1020 5023 1024
rect 5027 1020 5028 1024
rect 5022 1019 5028 1020
rect 5294 1024 5300 1025
rect 5294 1020 5295 1024
rect 5299 1020 5300 1024
rect 5294 1019 5300 1020
rect 5542 1024 5548 1025
rect 5542 1020 5543 1024
rect 5547 1020 5548 1024
rect 5662 1021 5663 1025
rect 5667 1021 5668 1025
rect 5662 1020 5668 1021
rect 5542 1019 5548 1020
rect 3858 1009 3864 1010
rect 1974 1008 1980 1009
rect 3798 1008 3804 1009
rect 1974 1004 1975 1008
rect 1979 1004 1980 1008
rect 1974 1003 1980 1004
rect 3090 1007 3096 1008
rect 3090 1003 3091 1007
rect 3095 1003 3096 1007
rect 3090 1002 3096 1003
rect 3242 1007 3248 1008
rect 3242 1003 3243 1007
rect 3247 1003 3248 1007
rect 3242 1002 3248 1003
rect 3394 1007 3400 1008
rect 3394 1003 3395 1007
rect 3399 1003 3400 1007
rect 3798 1004 3799 1008
rect 3803 1004 3804 1008
rect 3798 1003 3804 1004
rect 3838 1008 3844 1009
rect 3838 1004 3839 1008
rect 3843 1004 3844 1008
rect 3858 1005 3859 1009
rect 3863 1005 3864 1009
rect 3858 1004 3864 1005
rect 4042 1009 4048 1010
rect 4042 1005 4043 1009
rect 4047 1005 4048 1009
rect 4042 1004 4048 1005
rect 4250 1009 4256 1010
rect 4250 1005 4251 1009
rect 4255 1005 4256 1009
rect 4250 1004 4256 1005
rect 4482 1009 4488 1010
rect 4482 1005 4483 1009
rect 4487 1005 4488 1009
rect 4482 1004 4488 1005
rect 4730 1009 4736 1010
rect 4730 1005 4731 1009
rect 4735 1005 4736 1009
rect 4730 1004 4736 1005
rect 4994 1009 5000 1010
rect 4994 1005 4995 1009
rect 4999 1005 5000 1009
rect 4994 1004 5000 1005
rect 5266 1009 5272 1010
rect 5266 1005 5267 1009
rect 5271 1005 5272 1009
rect 5266 1004 5272 1005
rect 5514 1009 5520 1010
rect 5514 1005 5515 1009
rect 5519 1005 5520 1009
rect 5514 1004 5520 1005
rect 5662 1008 5668 1009
rect 5662 1004 5663 1008
rect 5667 1004 5668 1008
rect 3838 1003 3844 1004
rect 5662 1003 5668 1004
rect 3394 1002 3400 1003
rect 3118 992 3124 993
rect 1974 991 1980 992
rect 1974 987 1975 991
rect 1979 987 1980 991
rect 3118 988 3119 992
rect 3123 988 3124 992
rect 3118 987 3124 988
rect 3270 992 3276 993
rect 3270 988 3271 992
rect 3275 988 3276 992
rect 3270 987 3276 988
rect 3422 992 3428 993
rect 3422 988 3423 992
rect 3427 988 3428 992
rect 3422 987 3428 988
rect 3798 991 3804 992
rect 3798 987 3799 991
rect 3803 987 3804 991
rect 1974 986 1980 987
rect 3798 986 3804 987
rect 1974 905 1980 906
rect 3798 905 3804 906
rect 1974 901 1975 905
rect 1979 901 1980 905
rect 1974 900 1980 901
rect 2046 904 2052 905
rect 2046 900 2047 904
rect 2051 900 2052 904
rect 2046 899 2052 900
rect 2350 904 2356 905
rect 2350 900 2351 904
rect 2355 900 2356 904
rect 2350 899 2356 900
rect 2646 904 2652 905
rect 2646 900 2647 904
rect 2651 900 2652 904
rect 2646 899 2652 900
rect 2926 904 2932 905
rect 2926 900 2927 904
rect 2931 900 2932 904
rect 2926 899 2932 900
rect 3206 904 3212 905
rect 3206 900 3207 904
rect 3211 900 3212 904
rect 3206 899 3212 900
rect 3494 904 3500 905
rect 3494 900 3495 904
rect 3499 900 3500 904
rect 3798 901 3799 905
rect 3803 901 3804 905
rect 3798 900 3804 901
rect 3494 899 3500 900
rect 110 892 116 893
rect 1934 892 1940 893
rect 110 888 111 892
rect 115 888 116 892
rect 110 887 116 888
rect 226 891 232 892
rect 226 887 227 891
rect 231 887 232 891
rect 226 886 232 887
rect 378 891 384 892
rect 378 887 379 891
rect 383 887 384 891
rect 378 886 384 887
rect 538 891 544 892
rect 538 887 539 891
rect 543 887 544 891
rect 538 886 544 887
rect 714 891 720 892
rect 714 887 715 891
rect 719 887 720 891
rect 714 886 720 887
rect 890 891 896 892
rect 890 887 891 891
rect 895 887 896 891
rect 890 886 896 887
rect 1074 891 1080 892
rect 1074 887 1075 891
rect 1079 887 1080 891
rect 1074 886 1080 887
rect 1258 891 1264 892
rect 1258 887 1259 891
rect 1263 887 1264 891
rect 1258 886 1264 887
rect 1442 891 1448 892
rect 1442 887 1443 891
rect 1447 887 1448 891
rect 1442 886 1448 887
rect 1626 891 1632 892
rect 1626 887 1627 891
rect 1631 887 1632 891
rect 1626 886 1632 887
rect 1786 891 1792 892
rect 1786 887 1787 891
rect 1791 887 1792 891
rect 1934 888 1935 892
rect 1939 888 1940 892
rect 2018 889 2024 890
rect 1934 887 1940 888
rect 1974 888 1980 889
rect 1786 886 1792 887
rect 1974 884 1975 888
rect 1979 884 1980 888
rect 2018 885 2019 889
rect 2023 885 2024 889
rect 2018 884 2024 885
rect 2322 889 2328 890
rect 2322 885 2323 889
rect 2327 885 2328 889
rect 2322 884 2328 885
rect 2618 889 2624 890
rect 2618 885 2619 889
rect 2623 885 2624 889
rect 2618 884 2624 885
rect 2898 889 2904 890
rect 2898 885 2899 889
rect 2903 885 2904 889
rect 2898 884 2904 885
rect 3178 889 3184 890
rect 3178 885 3179 889
rect 3183 885 3184 889
rect 3178 884 3184 885
rect 3466 889 3472 890
rect 3466 885 3467 889
rect 3471 885 3472 889
rect 3466 884 3472 885
rect 3798 888 3804 889
rect 3798 884 3799 888
rect 3803 884 3804 888
rect 1974 883 1980 884
rect 3798 883 3804 884
rect 254 876 260 877
rect 110 875 116 876
rect 110 871 111 875
rect 115 871 116 875
rect 254 872 255 876
rect 259 872 260 876
rect 254 871 260 872
rect 406 876 412 877
rect 406 872 407 876
rect 411 872 412 876
rect 406 871 412 872
rect 566 876 572 877
rect 566 872 567 876
rect 571 872 572 876
rect 566 871 572 872
rect 742 876 748 877
rect 742 872 743 876
rect 747 872 748 876
rect 742 871 748 872
rect 918 876 924 877
rect 918 872 919 876
rect 923 872 924 876
rect 918 871 924 872
rect 1102 876 1108 877
rect 1102 872 1103 876
rect 1107 872 1108 876
rect 1102 871 1108 872
rect 1286 876 1292 877
rect 1286 872 1287 876
rect 1291 872 1292 876
rect 1286 871 1292 872
rect 1470 876 1476 877
rect 1470 872 1471 876
rect 1475 872 1476 876
rect 1470 871 1476 872
rect 1654 876 1660 877
rect 1654 872 1655 876
rect 1659 872 1660 876
rect 1654 871 1660 872
rect 1814 876 1820 877
rect 3838 876 3844 877
rect 5662 876 5668 877
rect 1814 872 1815 876
rect 1819 872 1820 876
rect 1814 871 1820 872
rect 1934 875 1940 876
rect 1934 871 1935 875
rect 1939 871 1940 875
rect 3838 872 3839 876
rect 3843 872 3844 876
rect 3838 871 3844 872
rect 3970 875 3976 876
rect 3970 871 3971 875
rect 3975 871 3976 875
rect 110 870 116 871
rect 1934 870 1940 871
rect 3970 870 3976 871
rect 4178 875 4184 876
rect 4178 871 4179 875
rect 4183 871 4184 875
rect 4178 870 4184 871
rect 4402 875 4408 876
rect 4402 871 4403 875
rect 4407 871 4408 875
rect 4402 870 4408 871
rect 4642 875 4648 876
rect 4642 871 4643 875
rect 4647 871 4648 875
rect 4642 870 4648 871
rect 4898 875 4904 876
rect 4898 871 4899 875
rect 4903 871 4904 875
rect 4898 870 4904 871
rect 5170 875 5176 876
rect 5170 871 5171 875
rect 5175 871 5176 875
rect 5170 870 5176 871
rect 5442 875 5448 876
rect 5442 871 5443 875
rect 5447 871 5448 875
rect 5662 872 5663 876
rect 5667 872 5668 876
rect 5662 871 5668 872
rect 5442 870 5448 871
rect 3998 860 4004 861
rect 3838 859 3844 860
rect 3838 855 3839 859
rect 3843 855 3844 859
rect 3998 856 3999 860
rect 4003 856 4004 860
rect 3998 855 4004 856
rect 4206 860 4212 861
rect 4206 856 4207 860
rect 4211 856 4212 860
rect 4206 855 4212 856
rect 4430 860 4436 861
rect 4430 856 4431 860
rect 4435 856 4436 860
rect 4430 855 4436 856
rect 4670 860 4676 861
rect 4670 856 4671 860
rect 4675 856 4676 860
rect 4670 855 4676 856
rect 4926 860 4932 861
rect 4926 856 4927 860
rect 4931 856 4932 860
rect 4926 855 4932 856
rect 5198 860 5204 861
rect 5198 856 5199 860
rect 5203 856 5204 860
rect 5198 855 5204 856
rect 5470 860 5476 861
rect 5470 856 5471 860
rect 5475 856 5476 860
rect 5470 855 5476 856
rect 5662 859 5668 860
rect 5662 855 5663 859
rect 5667 855 5668 859
rect 3838 854 3844 855
rect 5662 854 5668 855
rect 110 801 116 802
rect 1934 801 1940 802
rect 110 797 111 801
rect 115 797 116 801
rect 110 796 116 797
rect 374 800 380 801
rect 374 796 375 800
rect 379 796 380 800
rect 374 795 380 796
rect 654 800 660 801
rect 654 796 655 800
rect 659 796 660 800
rect 654 795 660 796
rect 942 800 948 801
rect 942 796 943 800
rect 947 796 948 800
rect 942 795 948 796
rect 1238 800 1244 801
rect 1238 796 1239 800
rect 1243 796 1244 800
rect 1238 795 1244 796
rect 1534 800 1540 801
rect 1534 796 1535 800
rect 1539 796 1540 800
rect 1534 795 1540 796
rect 1814 800 1820 801
rect 1814 796 1815 800
rect 1819 796 1820 800
rect 1934 797 1935 801
rect 1939 797 1940 801
rect 1934 796 1940 797
rect 3838 801 3844 802
rect 5662 801 5668 802
rect 3838 797 3839 801
rect 3843 797 3844 801
rect 3838 796 3844 797
rect 3886 800 3892 801
rect 3886 796 3887 800
rect 3891 796 3892 800
rect 1814 795 1820 796
rect 3886 795 3892 796
rect 4046 800 4052 801
rect 4046 796 4047 800
rect 4051 796 4052 800
rect 4046 795 4052 796
rect 4278 800 4284 801
rect 4278 796 4279 800
rect 4283 796 4284 800
rect 4278 795 4284 796
rect 4558 800 4564 801
rect 4558 796 4559 800
rect 4563 796 4564 800
rect 4558 795 4564 796
rect 4878 800 4884 801
rect 4878 796 4879 800
rect 4883 796 4884 800
rect 4878 795 4884 796
rect 5222 800 5228 801
rect 5222 796 5223 800
rect 5227 796 5228 800
rect 5222 795 5228 796
rect 5542 800 5548 801
rect 5542 796 5543 800
rect 5547 796 5548 800
rect 5662 797 5663 801
rect 5667 797 5668 801
rect 5662 796 5668 797
rect 5542 795 5548 796
rect 346 785 352 786
rect 110 784 116 785
rect 110 780 111 784
rect 115 780 116 784
rect 346 781 347 785
rect 351 781 352 785
rect 346 780 352 781
rect 626 785 632 786
rect 626 781 627 785
rect 631 781 632 785
rect 626 780 632 781
rect 914 785 920 786
rect 914 781 915 785
rect 919 781 920 785
rect 914 780 920 781
rect 1210 785 1216 786
rect 1210 781 1211 785
rect 1215 781 1216 785
rect 1210 780 1216 781
rect 1506 785 1512 786
rect 1506 781 1507 785
rect 1511 781 1512 785
rect 1506 780 1512 781
rect 1786 785 1792 786
rect 3858 785 3864 786
rect 1786 781 1787 785
rect 1791 781 1792 785
rect 1786 780 1792 781
rect 1934 784 1940 785
rect 1934 780 1935 784
rect 1939 780 1940 784
rect 110 779 116 780
rect 1934 779 1940 780
rect 3838 784 3844 785
rect 3838 780 3839 784
rect 3843 780 3844 784
rect 3858 781 3859 785
rect 3863 781 3864 785
rect 3858 780 3864 781
rect 4018 785 4024 786
rect 4018 781 4019 785
rect 4023 781 4024 785
rect 4018 780 4024 781
rect 4250 785 4256 786
rect 4250 781 4251 785
rect 4255 781 4256 785
rect 4250 780 4256 781
rect 4530 785 4536 786
rect 4530 781 4531 785
rect 4535 781 4536 785
rect 4530 780 4536 781
rect 4850 785 4856 786
rect 4850 781 4851 785
rect 4855 781 4856 785
rect 4850 780 4856 781
rect 5194 785 5200 786
rect 5194 781 5195 785
rect 5199 781 5200 785
rect 5194 780 5200 781
rect 5514 785 5520 786
rect 5514 781 5515 785
rect 5519 781 5520 785
rect 5514 780 5520 781
rect 5662 784 5668 785
rect 5662 780 5663 784
rect 5667 780 5668 784
rect 3838 779 3844 780
rect 5662 779 5668 780
rect 1974 756 1980 757
rect 3798 756 3804 757
rect 1974 752 1975 756
rect 1979 752 1980 756
rect 1974 751 1980 752
rect 1994 755 2000 756
rect 1994 751 1995 755
rect 1999 751 2000 755
rect 1994 750 2000 751
rect 2250 755 2256 756
rect 2250 751 2251 755
rect 2255 751 2256 755
rect 2250 750 2256 751
rect 2522 755 2528 756
rect 2522 751 2523 755
rect 2527 751 2528 755
rect 2522 750 2528 751
rect 2770 755 2776 756
rect 2770 751 2771 755
rect 2775 751 2776 755
rect 2770 750 2776 751
rect 3002 755 3008 756
rect 3002 751 3003 755
rect 3007 751 3008 755
rect 3002 750 3008 751
rect 3226 755 3232 756
rect 3226 751 3227 755
rect 3231 751 3232 755
rect 3226 750 3232 751
rect 3450 755 3456 756
rect 3450 751 3451 755
rect 3455 751 3456 755
rect 3450 750 3456 751
rect 3650 755 3656 756
rect 3650 751 3651 755
rect 3655 751 3656 755
rect 3798 752 3799 756
rect 3803 752 3804 756
rect 3798 751 3804 752
rect 3650 750 3656 751
rect 2022 740 2028 741
rect 1974 739 1980 740
rect 1974 735 1975 739
rect 1979 735 1980 739
rect 2022 736 2023 740
rect 2027 736 2028 740
rect 2022 735 2028 736
rect 2278 740 2284 741
rect 2278 736 2279 740
rect 2283 736 2284 740
rect 2278 735 2284 736
rect 2550 740 2556 741
rect 2550 736 2551 740
rect 2555 736 2556 740
rect 2550 735 2556 736
rect 2798 740 2804 741
rect 2798 736 2799 740
rect 2803 736 2804 740
rect 2798 735 2804 736
rect 3030 740 3036 741
rect 3030 736 3031 740
rect 3035 736 3036 740
rect 3030 735 3036 736
rect 3254 740 3260 741
rect 3254 736 3255 740
rect 3259 736 3260 740
rect 3254 735 3260 736
rect 3478 740 3484 741
rect 3478 736 3479 740
rect 3483 736 3484 740
rect 3478 735 3484 736
rect 3678 740 3684 741
rect 3678 736 3679 740
rect 3683 736 3684 740
rect 3678 735 3684 736
rect 3798 739 3804 740
rect 3798 735 3799 739
rect 3803 735 3804 739
rect 1974 734 1980 735
rect 3798 734 3804 735
rect 110 652 116 653
rect 1934 652 1940 653
rect 110 648 111 652
rect 115 648 116 652
rect 110 647 116 648
rect 130 651 136 652
rect 130 647 131 651
rect 135 647 136 651
rect 130 646 136 647
rect 306 651 312 652
rect 306 647 307 651
rect 311 647 312 651
rect 306 646 312 647
rect 498 651 504 652
rect 498 647 499 651
rect 503 647 504 651
rect 498 646 504 647
rect 682 651 688 652
rect 682 647 683 651
rect 687 647 688 651
rect 682 646 688 647
rect 858 651 864 652
rect 858 647 859 651
rect 863 647 864 651
rect 858 646 864 647
rect 1026 651 1032 652
rect 1026 647 1027 651
rect 1031 647 1032 651
rect 1026 646 1032 647
rect 1186 651 1192 652
rect 1186 647 1187 651
rect 1191 647 1192 651
rect 1186 646 1192 647
rect 1338 651 1344 652
rect 1338 647 1339 651
rect 1343 647 1344 651
rect 1338 646 1344 647
rect 1490 651 1496 652
rect 1490 647 1491 651
rect 1495 647 1496 651
rect 1490 646 1496 647
rect 1650 651 1656 652
rect 1650 647 1651 651
rect 1655 647 1656 651
rect 1650 646 1656 647
rect 1786 651 1792 652
rect 1786 647 1787 651
rect 1791 647 1792 651
rect 1934 648 1935 652
rect 1939 648 1940 652
rect 1934 647 1940 648
rect 1786 646 1792 647
rect 3838 644 3844 645
rect 5662 644 5668 645
rect 3838 640 3839 644
rect 3843 640 3844 644
rect 3838 639 3844 640
rect 3858 643 3864 644
rect 3858 639 3859 643
rect 3863 639 3864 643
rect 3858 638 3864 639
rect 3994 643 4000 644
rect 3994 639 3995 643
rect 3999 639 4000 643
rect 3994 638 4000 639
rect 4130 643 4136 644
rect 4130 639 4131 643
rect 4135 639 4136 643
rect 4130 638 4136 639
rect 4266 643 4272 644
rect 4266 639 4267 643
rect 4271 639 4272 643
rect 4266 638 4272 639
rect 4402 643 4408 644
rect 4402 639 4403 643
rect 4407 639 4408 643
rect 4402 638 4408 639
rect 4570 643 4576 644
rect 4570 639 4571 643
rect 4575 639 4576 643
rect 4570 638 4576 639
rect 4770 643 4776 644
rect 4770 639 4771 643
rect 4775 639 4776 643
rect 4770 638 4776 639
rect 4994 643 5000 644
rect 4994 639 4995 643
rect 4999 639 5000 643
rect 4994 638 5000 639
rect 5226 643 5232 644
rect 5226 639 5227 643
rect 5231 639 5232 643
rect 5226 638 5232 639
rect 5458 643 5464 644
rect 5458 639 5459 643
rect 5463 639 5464 643
rect 5662 640 5663 644
rect 5667 640 5668 644
rect 5662 639 5668 640
rect 5458 638 5464 639
rect 158 636 164 637
rect 110 635 116 636
rect 110 631 111 635
rect 115 631 116 635
rect 158 632 159 636
rect 163 632 164 636
rect 158 631 164 632
rect 334 636 340 637
rect 334 632 335 636
rect 339 632 340 636
rect 334 631 340 632
rect 526 636 532 637
rect 526 632 527 636
rect 531 632 532 636
rect 526 631 532 632
rect 710 636 716 637
rect 710 632 711 636
rect 715 632 716 636
rect 710 631 716 632
rect 886 636 892 637
rect 886 632 887 636
rect 891 632 892 636
rect 886 631 892 632
rect 1054 636 1060 637
rect 1054 632 1055 636
rect 1059 632 1060 636
rect 1054 631 1060 632
rect 1214 636 1220 637
rect 1214 632 1215 636
rect 1219 632 1220 636
rect 1214 631 1220 632
rect 1366 636 1372 637
rect 1366 632 1367 636
rect 1371 632 1372 636
rect 1366 631 1372 632
rect 1518 636 1524 637
rect 1518 632 1519 636
rect 1523 632 1524 636
rect 1518 631 1524 632
rect 1678 636 1684 637
rect 1678 632 1679 636
rect 1683 632 1684 636
rect 1678 631 1684 632
rect 1814 636 1820 637
rect 1814 632 1815 636
rect 1819 632 1820 636
rect 1814 631 1820 632
rect 1934 635 1940 636
rect 1934 631 1935 635
rect 1939 631 1940 635
rect 110 630 116 631
rect 1934 630 1940 631
rect 3886 628 3892 629
rect 3838 627 3844 628
rect 3838 623 3839 627
rect 3843 623 3844 627
rect 3886 624 3887 628
rect 3891 624 3892 628
rect 3886 623 3892 624
rect 4022 628 4028 629
rect 4022 624 4023 628
rect 4027 624 4028 628
rect 4022 623 4028 624
rect 4158 628 4164 629
rect 4158 624 4159 628
rect 4163 624 4164 628
rect 4158 623 4164 624
rect 4294 628 4300 629
rect 4294 624 4295 628
rect 4299 624 4300 628
rect 4294 623 4300 624
rect 4430 628 4436 629
rect 4430 624 4431 628
rect 4435 624 4436 628
rect 4430 623 4436 624
rect 4598 628 4604 629
rect 4598 624 4599 628
rect 4603 624 4604 628
rect 4598 623 4604 624
rect 4798 628 4804 629
rect 4798 624 4799 628
rect 4803 624 4804 628
rect 4798 623 4804 624
rect 5022 628 5028 629
rect 5022 624 5023 628
rect 5027 624 5028 628
rect 5022 623 5028 624
rect 5254 628 5260 629
rect 5254 624 5255 628
rect 5259 624 5260 628
rect 5254 623 5260 624
rect 5486 628 5492 629
rect 5486 624 5487 628
rect 5491 624 5492 628
rect 5486 623 5492 624
rect 5662 627 5668 628
rect 5662 623 5663 627
rect 5667 623 5668 627
rect 3838 622 3844 623
rect 5662 622 5668 623
rect 110 577 116 578
rect 1934 577 1940 578
rect 110 573 111 577
rect 115 573 116 577
rect 110 572 116 573
rect 158 576 164 577
rect 158 572 159 576
rect 163 572 164 576
rect 158 571 164 572
rect 374 576 380 577
rect 374 572 375 576
rect 379 572 380 576
rect 374 571 380 572
rect 598 576 604 577
rect 598 572 599 576
rect 603 572 604 576
rect 598 571 604 572
rect 806 576 812 577
rect 806 572 807 576
rect 811 572 812 576
rect 806 571 812 572
rect 998 576 1004 577
rect 998 572 999 576
rect 1003 572 1004 576
rect 998 571 1004 572
rect 1174 576 1180 577
rect 1174 572 1175 576
rect 1179 572 1180 576
rect 1174 571 1180 572
rect 1342 576 1348 577
rect 1342 572 1343 576
rect 1347 572 1348 576
rect 1342 571 1348 572
rect 1510 576 1516 577
rect 1510 572 1511 576
rect 1515 572 1516 576
rect 1510 571 1516 572
rect 1670 576 1676 577
rect 1670 572 1671 576
rect 1675 572 1676 576
rect 1670 571 1676 572
rect 1814 576 1820 577
rect 1814 572 1815 576
rect 1819 572 1820 576
rect 1934 573 1935 577
rect 1939 573 1940 577
rect 1934 572 1940 573
rect 1814 571 1820 572
rect 3838 569 3844 570
rect 5662 569 5668 570
rect 3838 565 3839 569
rect 3843 565 3844 569
rect 3838 564 3844 565
rect 3886 568 3892 569
rect 3886 564 3887 568
rect 3891 564 3892 568
rect 3886 563 3892 564
rect 4022 568 4028 569
rect 4022 564 4023 568
rect 4027 564 4028 568
rect 4022 563 4028 564
rect 4158 568 4164 569
rect 4158 564 4159 568
rect 4163 564 4164 568
rect 4158 563 4164 564
rect 4294 568 4300 569
rect 4294 564 4295 568
rect 4299 564 4300 568
rect 4294 563 4300 564
rect 4478 568 4484 569
rect 4478 564 4479 568
rect 4483 564 4484 568
rect 4478 563 4484 564
rect 4694 568 4700 569
rect 4694 564 4695 568
rect 4699 564 4700 568
rect 4694 563 4700 564
rect 4934 568 4940 569
rect 4934 564 4935 568
rect 4939 564 4940 568
rect 4934 563 4940 564
rect 5190 568 5196 569
rect 5190 564 5191 568
rect 5195 564 5196 568
rect 5190 563 5196 564
rect 5446 568 5452 569
rect 5446 564 5447 568
rect 5451 564 5452 568
rect 5662 565 5663 569
rect 5667 565 5668 569
rect 5662 564 5668 565
rect 5446 563 5452 564
rect 130 561 136 562
rect 110 560 116 561
rect 110 556 111 560
rect 115 556 116 560
rect 130 557 131 561
rect 135 557 136 561
rect 130 556 136 557
rect 346 561 352 562
rect 346 557 347 561
rect 351 557 352 561
rect 346 556 352 557
rect 570 561 576 562
rect 570 557 571 561
rect 575 557 576 561
rect 570 556 576 557
rect 778 561 784 562
rect 778 557 779 561
rect 783 557 784 561
rect 778 556 784 557
rect 970 561 976 562
rect 970 557 971 561
rect 975 557 976 561
rect 970 556 976 557
rect 1146 561 1152 562
rect 1146 557 1147 561
rect 1151 557 1152 561
rect 1146 556 1152 557
rect 1314 561 1320 562
rect 1314 557 1315 561
rect 1319 557 1320 561
rect 1314 556 1320 557
rect 1482 561 1488 562
rect 1482 557 1483 561
rect 1487 557 1488 561
rect 1482 556 1488 557
rect 1642 561 1648 562
rect 1642 557 1643 561
rect 1647 557 1648 561
rect 1642 556 1648 557
rect 1786 561 1792 562
rect 1786 557 1787 561
rect 1791 557 1792 561
rect 1786 556 1792 557
rect 1934 560 1940 561
rect 1934 556 1935 560
rect 1939 556 1940 560
rect 110 555 116 556
rect 1934 555 1940 556
rect 3858 553 3864 554
rect 3838 552 3844 553
rect 1974 549 1980 550
rect 3798 549 3804 550
rect 1974 545 1975 549
rect 1979 545 1980 549
rect 1974 544 1980 545
rect 3310 548 3316 549
rect 3310 544 3311 548
rect 3315 544 3316 548
rect 3310 543 3316 544
rect 3446 548 3452 549
rect 3446 544 3447 548
rect 3451 544 3452 548
rect 3446 543 3452 544
rect 3582 548 3588 549
rect 3582 544 3583 548
rect 3587 544 3588 548
rect 3798 545 3799 549
rect 3803 545 3804 549
rect 3838 548 3839 552
rect 3843 548 3844 552
rect 3858 549 3859 553
rect 3863 549 3864 553
rect 3858 548 3864 549
rect 3994 553 4000 554
rect 3994 549 3995 553
rect 3999 549 4000 553
rect 3994 548 4000 549
rect 4130 553 4136 554
rect 4130 549 4131 553
rect 4135 549 4136 553
rect 4130 548 4136 549
rect 4266 553 4272 554
rect 4266 549 4267 553
rect 4271 549 4272 553
rect 4266 548 4272 549
rect 4450 553 4456 554
rect 4450 549 4451 553
rect 4455 549 4456 553
rect 4450 548 4456 549
rect 4666 553 4672 554
rect 4666 549 4667 553
rect 4671 549 4672 553
rect 4666 548 4672 549
rect 4906 553 4912 554
rect 4906 549 4907 553
rect 4911 549 4912 553
rect 4906 548 4912 549
rect 5162 553 5168 554
rect 5162 549 5163 553
rect 5167 549 5168 553
rect 5162 548 5168 549
rect 5418 553 5424 554
rect 5418 549 5419 553
rect 5423 549 5424 553
rect 5418 548 5424 549
rect 5662 552 5668 553
rect 5662 548 5663 552
rect 5667 548 5668 552
rect 3838 547 3844 548
rect 5662 547 5668 548
rect 3798 544 3804 545
rect 3582 543 3588 544
rect 3282 533 3288 534
rect 1974 532 1980 533
rect 1974 528 1975 532
rect 1979 528 1980 532
rect 3282 529 3283 533
rect 3287 529 3288 533
rect 3282 528 3288 529
rect 3418 533 3424 534
rect 3418 529 3419 533
rect 3423 529 3424 533
rect 3418 528 3424 529
rect 3554 533 3560 534
rect 3554 529 3555 533
rect 3559 529 3560 533
rect 3554 528 3560 529
rect 3798 532 3804 533
rect 3798 528 3799 532
rect 3803 528 3804 532
rect 1974 527 1980 528
rect 3798 527 3804 528
rect 110 428 116 429
rect 1934 428 1940 429
rect 110 424 111 428
rect 115 424 116 428
rect 110 423 116 424
rect 130 427 136 428
rect 130 423 131 427
rect 135 423 136 427
rect 130 422 136 423
rect 426 427 432 428
rect 426 423 427 427
rect 431 423 432 427
rect 426 422 432 423
rect 762 427 768 428
rect 762 423 763 427
rect 767 423 768 427
rect 762 422 768 423
rect 1106 427 1112 428
rect 1106 423 1107 427
rect 1111 423 1112 427
rect 1106 422 1112 423
rect 1458 427 1464 428
rect 1458 423 1459 427
rect 1463 423 1464 427
rect 1458 422 1464 423
rect 1786 427 1792 428
rect 1786 423 1787 427
rect 1791 423 1792 427
rect 1934 424 1935 428
rect 1939 424 1940 428
rect 1934 423 1940 424
rect 1786 422 1792 423
rect 158 412 164 413
rect 110 411 116 412
rect 110 407 111 411
rect 115 407 116 411
rect 158 408 159 412
rect 163 408 164 412
rect 158 407 164 408
rect 454 412 460 413
rect 454 408 455 412
rect 459 408 460 412
rect 454 407 460 408
rect 790 412 796 413
rect 790 408 791 412
rect 795 408 796 412
rect 790 407 796 408
rect 1134 412 1140 413
rect 1134 408 1135 412
rect 1139 408 1140 412
rect 1134 407 1140 408
rect 1486 412 1492 413
rect 1486 408 1487 412
rect 1491 408 1492 412
rect 1486 407 1492 408
rect 1814 412 1820 413
rect 1814 408 1815 412
rect 1819 408 1820 412
rect 1814 407 1820 408
rect 1934 411 1940 412
rect 1934 407 1935 411
rect 1939 407 1940 411
rect 110 406 116 407
rect 1934 406 1940 407
rect 3838 408 3844 409
rect 5662 408 5668 409
rect 3838 404 3839 408
rect 3843 404 3844 408
rect 3838 403 3844 404
rect 4450 407 4456 408
rect 4450 403 4451 407
rect 4455 403 4456 407
rect 4450 402 4456 403
rect 4650 407 4656 408
rect 4650 403 4651 407
rect 4655 403 4656 407
rect 4650 402 4656 403
rect 4858 407 4864 408
rect 4858 403 4859 407
rect 4863 403 4864 407
rect 4858 402 4864 403
rect 5066 407 5072 408
rect 5066 403 5067 407
rect 5071 403 5072 407
rect 5066 402 5072 403
rect 5282 407 5288 408
rect 5282 403 5283 407
rect 5287 403 5288 407
rect 5282 402 5288 403
rect 5506 407 5512 408
rect 5506 403 5507 407
rect 5511 403 5512 407
rect 5662 404 5663 408
rect 5667 404 5668 408
rect 5662 403 5668 404
rect 5506 402 5512 403
rect 1974 400 1980 401
rect 3798 400 3804 401
rect 1974 396 1975 400
rect 1979 396 1980 400
rect 1974 395 1980 396
rect 1994 399 2000 400
rect 1994 395 1995 399
rect 1999 395 2000 399
rect 1994 394 2000 395
rect 2154 399 2160 400
rect 2154 395 2155 399
rect 2159 395 2160 399
rect 2154 394 2160 395
rect 2346 399 2352 400
rect 2346 395 2347 399
rect 2351 395 2352 399
rect 2346 394 2352 395
rect 2538 399 2544 400
rect 2538 395 2539 399
rect 2543 395 2544 399
rect 2538 394 2544 395
rect 2730 399 2736 400
rect 2730 395 2731 399
rect 2735 395 2736 399
rect 2730 394 2736 395
rect 2922 399 2928 400
rect 2922 395 2923 399
rect 2927 395 2928 399
rect 2922 394 2928 395
rect 3114 399 3120 400
rect 3114 395 3115 399
rect 3119 395 3120 399
rect 3114 394 3120 395
rect 3298 399 3304 400
rect 3298 395 3299 399
rect 3303 395 3304 399
rect 3298 394 3304 395
rect 3482 399 3488 400
rect 3482 395 3483 399
rect 3487 395 3488 399
rect 3482 394 3488 395
rect 3650 399 3656 400
rect 3650 395 3651 399
rect 3655 395 3656 399
rect 3798 396 3799 400
rect 3803 396 3804 400
rect 3798 395 3804 396
rect 3650 394 3656 395
rect 4478 392 4484 393
rect 3838 391 3844 392
rect 3838 387 3839 391
rect 3843 387 3844 391
rect 4478 388 4479 392
rect 4483 388 4484 392
rect 4478 387 4484 388
rect 4678 392 4684 393
rect 4678 388 4679 392
rect 4683 388 4684 392
rect 4678 387 4684 388
rect 4886 392 4892 393
rect 4886 388 4887 392
rect 4891 388 4892 392
rect 4886 387 4892 388
rect 5094 392 5100 393
rect 5094 388 5095 392
rect 5099 388 5100 392
rect 5094 387 5100 388
rect 5310 392 5316 393
rect 5310 388 5311 392
rect 5315 388 5316 392
rect 5310 387 5316 388
rect 5534 392 5540 393
rect 5534 388 5535 392
rect 5539 388 5540 392
rect 5534 387 5540 388
rect 5662 391 5668 392
rect 5662 387 5663 391
rect 5667 387 5668 391
rect 3838 386 3844 387
rect 5662 386 5668 387
rect 2022 384 2028 385
rect 1974 383 1980 384
rect 1974 379 1975 383
rect 1979 379 1980 383
rect 2022 380 2023 384
rect 2027 380 2028 384
rect 2022 379 2028 380
rect 2182 384 2188 385
rect 2182 380 2183 384
rect 2187 380 2188 384
rect 2182 379 2188 380
rect 2374 384 2380 385
rect 2374 380 2375 384
rect 2379 380 2380 384
rect 2374 379 2380 380
rect 2566 384 2572 385
rect 2566 380 2567 384
rect 2571 380 2572 384
rect 2566 379 2572 380
rect 2758 384 2764 385
rect 2758 380 2759 384
rect 2763 380 2764 384
rect 2758 379 2764 380
rect 2950 384 2956 385
rect 2950 380 2951 384
rect 2955 380 2956 384
rect 2950 379 2956 380
rect 3142 384 3148 385
rect 3142 380 3143 384
rect 3147 380 3148 384
rect 3142 379 3148 380
rect 3326 384 3332 385
rect 3326 380 3327 384
rect 3331 380 3332 384
rect 3326 379 3332 380
rect 3510 384 3516 385
rect 3510 380 3511 384
rect 3515 380 3516 384
rect 3510 379 3516 380
rect 3678 384 3684 385
rect 3678 380 3679 384
rect 3683 380 3684 384
rect 3678 379 3684 380
rect 3798 383 3804 384
rect 3798 379 3799 383
rect 3803 379 3804 383
rect 1974 378 1980 379
rect 3798 378 3804 379
rect 110 337 116 338
rect 1934 337 1940 338
rect 110 333 111 337
rect 115 333 116 337
rect 110 332 116 333
rect 238 336 244 337
rect 238 332 239 336
rect 243 332 244 336
rect 238 331 244 332
rect 390 336 396 337
rect 390 332 391 336
rect 395 332 396 336
rect 390 331 396 332
rect 550 336 556 337
rect 550 332 551 336
rect 555 332 556 336
rect 550 331 556 332
rect 710 336 716 337
rect 710 332 711 336
rect 715 332 716 336
rect 710 331 716 332
rect 870 336 876 337
rect 870 332 871 336
rect 875 332 876 336
rect 870 331 876 332
rect 1030 336 1036 337
rect 1030 332 1031 336
rect 1035 332 1036 336
rect 1934 333 1935 337
rect 1939 333 1940 337
rect 1934 332 1940 333
rect 1030 331 1036 332
rect 3838 329 3844 330
rect 5662 329 5668 330
rect 3838 325 3839 329
rect 3843 325 3844 329
rect 3838 324 3844 325
rect 4750 328 4756 329
rect 4750 324 4751 328
rect 4755 324 4756 328
rect 4750 323 4756 324
rect 4910 328 4916 329
rect 4910 324 4911 328
rect 4915 324 4916 328
rect 4910 323 4916 324
rect 5070 328 5076 329
rect 5070 324 5071 328
rect 5075 324 5076 328
rect 5070 323 5076 324
rect 5230 328 5236 329
rect 5230 324 5231 328
rect 5235 324 5236 328
rect 5230 323 5236 324
rect 5398 328 5404 329
rect 5398 324 5399 328
rect 5403 324 5404 328
rect 5398 323 5404 324
rect 5542 328 5548 329
rect 5542 324 5543 328
rect 5547 324 5548 328
rect 5662 325 5663 329
rect 5667 325 5668 329
rect 5662 324 5668 325
rect 5542 323 5548 324
rect 210 321 216 322
rect 110 320 116 321
rect 110 316 111 320
rect 115 316 116 320
rect 210 317 211 321
rect 215 317 216 321
rect 210 316 216 317
rect 362 321 368 322
rect 362 317 363 321
rect 367 317 368 321
rect 362 316 368 317
rect 522 321 528 322
rect 522 317 523 321
rect 527 317 528 321
rect 522 316 528 317
rect 682 321 688 322
rect 682 317 683 321
rect 687 317 688 321
rect 682 316 688 317
rect 842 321 848 322
rect 842 317 843 321
rect 847 317 848 321
rect 842 316 848 317
rect 1002 321 1008 322
rect 1002 317 1003 321
rect 1007 317 1008 321
rect 1002 316 1008 317
rect 1934 320 1940 321
rect 1934 316 1935 320
rect 1939 316 1940 320
rect 110 315 116 316
rect 1934 315 1940 316
rect 4722 313 4728 314
rect 3838 312 3844 313
rect 3838 308 3839 312
rect 3843 308 3844 312
rect 4722 309 4723 313
rect 4727 309 4728 313
rect 4722 308 4728 309
rect 4882 313 4888 314
rect 4882 309 4883 313
rect 4887 309 4888 313
rect 4882 308 4888 309
rect 5042 313 5048 314
rect 5042 309 5043 313
rect 5047 309 5048 313
rect 5042 308 5048 309
rect 5202 313 5208 314
rect 5202 309 5203 313
rect 5207 309 5208 313
rect 5202 308 5208 309
rect 5370 313 5376 314
rect 5370 309 5371 313
rect 5375 309 5376 313
rect 5370 308 5376 309
rect 5514 313 5520 314
rect 5514 309 5515 313
rect 5519 309 5520 313
rect 5514 308 5520 309
rect 5662 312 5668 313
rect 5662 308 5663 312
rect 5667 308 5668 312
rect 3838 307 3844 308
rect 5662 307 5668 308
rect 1974 301 1980 302
rect 3798 301 3804 302
rect 1974 297 1975 301
rect 1979 297 1980 301
rect 1974 296 1980 297
rect 2046 300 2052 301
rect 2046 296 2047 300
rect 2051 296 2052 300
rect 2046 295 2052 296
rect 2182 300 2188 301
rect 2182 296 2183 300
rect 2187 296 2188 300
rect 2182 295 2188 296
rect 2318 300 2324 301
rect 2318 296 2319 300
rect 2323 296 2324 300
rect 2318 295 2324 296
rect 2454 300 2460 301
rect 2454 296 2455 300
rect 2459 296 2460 300
rect 2454 295 2460 296
rect 2590 300 2596 301
rect 2590 296 2591 300
rect 2595 296 2596 300
rect 2590 295 2596 296
rect 2726 300 2732 301
rect 2726 296 2727 300
rect 2731 296 2732 300
rect 2726 295 2732 296
rect 2862 300 2868 301
rect 2862 296 2863 300
rect 2867 296 2868 300
rect 2862 295 2868 296
rect 2998 300 3004 301
rect 2998 296 2999 300
rect 3003 296 3004 300
rect 2998 295 3004 296
rect 3134 300 3140 301
rect 3134 296 3135 300
rect 3139 296 3140 300
rect 3134 295 3140 296
rect 3270 300 3276 301
rect 3270 296 3271 300
rect 3275 296 3276 300
rect 3270 295 3276 296
rect 3406 300 3412 301
rect 3406 296 3407 300
rect 3411 296 3412 300
rect 3406 295 3412 296
rect 3542 300 3548 301
rect 3542 296 3543 300
rect 3547 296 3548 300
rect 3542 295 3548 296
rect 3678 300 3684 301
rect 3678 296 3679 300
rect 3683 296 3684 300
rect 3798 297 3799 301
rect 3803 297 3804 301
rect 3798 296 3804 297
rect 3678 295 3684 296
rect 2018 285 2024 286
rect 1974 284 1980 285
rect 1974 280 1975 284
rect 1979 280 1980 284
rect 2018 281 2019 285
rect 2023 281 2024 285
rect 2018 280 2024 281
rect 2154 285 2160 286
rect 2154 281 2155 285
rect 2159 281 2160 285
rect 2154 280 2160 281
rect 2290 285 2296 286
rect 2290 281 2291 285
rect 2295 281 2296 285
rect 2290 280 2296 281
rect 2426 285 2432 286
rect 2426 281 2427 285
rect 2431 281 2432 285
rect 2426 280 2432 281
rect 2562 285 2568 286
rect 2562 281 2563 285
rect 2567 281 2568 285
rect 2562 280 2568 281
rect 2698 285 2704 286
rect 2698 281 2699 285
rect 2703 281 2704 285
rect 2698 280 2704 281
rect 2834 285 2840 286
rect 2834 281 2835 285
rect 2839 281 2840 285
rect 2834 280 2840 281
rect 2970 285 2976 286
rect 2970 281 2971 285
rect 2975 281 2976 285
rect 2970 280 2976 281
rect 3106 285 3112 286
rect 3106 281 3107 285
rect 3111 281 3112 285
rect 3106 280 3112 281
rect 3242 285 3248 286
rect 3242 281 3243 285
rect 3247 281 3248 285
rect 3242 280 3248 281
rect 3378 285 3384 286
rect 3378 281 3379 285
rect 3383 281 3384 285
rect 3378 280 3384 281
rect 3514 285 3520 286
rect 3514 281 3515 285
rect 3519 281 3520 285
rect 3514 280 3520 281
rect 3650 285 3656 286
rect 3650 281 3651 285
rect 3655 281 3656 285
rect 3650 280 3656 281
rect 3798 284 3804 285
rect 3798 280 3799 284
rect 3803 280 3804 284
rect 1974 279 1980 280
rect 3798 279 3804 280
rect 110 156 116 157
rect 1934 156 1940 157
rect 110 152 111 156
rect 115 152 116 156
rect 110 151 116 152
rect 146 155 152 156
rect 146 151 147 155
rect 151 151 152 155
rect 146 150 152 151
rect 282 155 288 156
rect 282 151 283 155
rect 287 151 288 155
rect 282 150 288 151
rect 418 155 424 156
rect 418 151 419 155
rect 423 151 424 155
rect 418 150 424 151
rect 554 155 560 156
rect 554 151 555 155
rect 559 151 560 155
rect 554 150 560 151
rect 690 155 696 156
rect 690 151 691 155
rect 695 151 696 155
rect 690 150 696 151
rect 826 155 832 156
rect 826 151 827 155
rect 831 151 832 155
rect 826 150 832 151
rect 962 155 968 156
rect 962 151 963 155
rect 967 151 968 155
rect 962 150 968 151
rect 1098 155 1104 156
rect 1098 151 1099 155
rect 1103 151 1104 155
rect 1934 152 1935 156
rect 1939 152 1940 156
rect 1934 151 1940 152
rect 1098 150 1104 151
rect 174 140 180 141
rect 110 139 116 140
rect 110 135 111 139
rect 115 135 116 139
rect 174 136 175 140
rect 179 136 180 140
rect 174 135 180 136
rect 310 140 316 141
rect 310 136 311 140
rect 315 136 316 140
rect 310 135 316 136
rect 446 140 452 141
rect 446 136 447 140
rect 451 136 452 140
rect 446 135 452 136
rect 582 140 588 141
rect 582 136 583 140
rect 587 136 588 140
rect 582 135 588 136
rect 718 140 724 141
rect 718 136 719 140
rect 723 136 724 140
rect 718 135 724 136
rect 854 140 860 141
rect 854 136 855 140
rect 859 136 860 140
rect 854 135 860 136
rect 990 140 996 141
rect 990 136 991 140
rect 995 136 996 140
rect 990 135 996 136
rect 1126 140 1132 141
rect 3838 140 3844 141
rect 5662 140 5668 141
rect 1126 136 1127 140
rect 1131 136 1132 140
rect 1126 135 1132 136
rect 1934 139 1940 140
rect 1934 135 1935 139
rect 1939 135 1940 139
rect 110 134 116 135
rect 1934 134 1940 135
rect 1974 136 1980 137
rect 3798 136 3804 137
rect 1974 132 1975 136
rect 1979 132 1980 136
rect 1974 131 1980 132
rect 1994 135 2000 136
rect 1994 131 1995 135
rect 1999 131 2000 135
rect 1994 130 2000 131
rect 2130 135 2136 136
rect 2130 131 2131 135
rect 2135 131 2136 135
rect 2130 130 2136 131
rect 2266 135 2272 136
rect 2266 131 2267 135
rect 2271 131 2272 135
rect 2266 130 2272 131
rect 2402 135 2408 136
rect 2402 131 2403 135
rect 2407 131 2408 135
rect 2402 130 2408 131
rect 2538 135 2544 136
rect 2538 131 2539 135
rect 2543 131 2544 135
rect 2538 130 2544 131
rect 2674 135 2680 136
rect 2674 131 2675 135
rect 2679 131 2680 135
rect 2674 130 2680 131
rect 2810 135 2816 136
rect 2810 131 2811 135
rect 2815 131 2816 135
rect 2810 130 2816 131
rect 2946 135 2952 136
rect 2946 131 2947 135
rect 2951 131 2952 135
rect 2946 130 2952 131
rect 3082 135 3088 136
rect 3082 131 3083 135
rect 3087 131 3088 135
rect 3082 130 3088 131
rect 3218 135 3224 136
rect 3218 131 3219 135
rect 3223 131 3224 135
rect 3218 130 3224 131
rect 3354 135 3360 136
rect 3354 131 3355 135
rect 3359 131 3360 135
rect 3354 130 3360 131
rect 3490 135 3496 136
rect 3490 131 3491 135
rect 3495 131 3496 135
rect 3490 130 3496 131
rect 3626 135 3632 136
rect 3626 131 3627 135
rect 3631 131 3632 135
rect 3798 132 3799 136
rect 3803 132 3804 136
rect 3838 136 3839 140
rect 3843 136 3844 140
rect 3838 135 3844 136
rect 4290 139 4296 140
rect 4290 135 4291 139
rect 4295 135 4296 139
rect 4290 134 4296 135
rect 4426 139 4432 140
rect 4426 135 4427 139
rect 4431 135 4432 139
rect 4426 134 4432 135
rect 4562 139 4568 140
rect 4562 135 4563 139
rect 4567 135 4568 139
rect 4562 134 4568 135
rect 4698 139 4704 140
rect 4698 135 4699 139
rect 4703 135 4704 139
rect 4698 134 4704 135
rect 4834 139 4840 140
rect 4834 135 4835 139
rect 4839 135 4840 139
rect 4834 134 4840 135
rect 4970 139 4976 140
rect 4970 135 4971 139
rect 4975 135 4976 139
rect 4970 134 4976 135
rect 5106 139 5112 140
rect 5106 135 5107 139
rect 5111 135 5112 139
rect 5106 134 5112 135
rect 5242 139 5248 140
rect 5242 135 5243 139
rect 5247 135 5248 139
rect 5242 134 5248 135
rect 5378 139 5384 140
rect 5378 135 5379 139
rect 5383 135 5384 139
rect 5378 134 5384 135
rect 5514 139 5520 140
rect 5514 135 5515 139
rect 5519 135 5520 139
rect 5662 136 5663 140
rect 5667 136 5668 140
rect 5662 135 5668 136
rect 5514 134 5520 135
rect 3798 131 3804 132
rect 3626 130 3632 131
rect 4318 124 4324 125
rect 3838 123 3844 124
rect 2022 120 2028 121
rect 1974 119 1980 120
rect 1974 115 1975 119
rect 1979 115 1980 119
rect 2022 116 2023 120
rect 2027 116 2028 120
rect 2022 115 2028 116
rect 2158 120 2164 121
rect 2158 116 2159 120
rect 2163 116 2164 120
rect 2158 115 2164 116
rect 2294 120 2300 121
rect 2294 116 2295 120
rect 2299 116 2300 120
rect 2294 115 2300 116
rect 2430 120 2436 121
rect 2430 116 2431 120
rect 2435 116 2436 120
rect 2430 115 2436 116
rect 2566 120 2572 121
rect 2566 116 2567 120
rect 2571 116 2572 120
rect 2566 115 2572 116
rect 2702 120 2708 121
rect 2702 116 2703 120
rect 2707 116 2708 120
rect 2702 115 2708 116
rect 2838 120 2844 121
rect 2838 116 2839 120
rect 2843 116 2844 120
rect 2838 115 2844 116
rect 2974 120 2980 121
rect 2974 116 2975 120
rect 2979 116 2980 120
rect 2974 115 2980 116
rect 3110 120 3116 121
rect 3110 116 3111 120
rect 3115 116 3116 120
rect 3110 115 3116 116
rect 3246 120 3252 121
rect 3246 116 3247 120
rect 3251 116 3252 120
rect 3246 115 3252 116
rect 3382 120 3388 121
rect 3382 116 3383 120
rect 3387 116 3388 120
rect 3382 115 3388 116
rect 3518 120 3524 121
rect 3518 116 3519 120
rect 3523 116 3524 120
rect 3518 115 3524 116
rect 3654 120 3660 121
rect 3654 116 3655 120
rect 3659 116 3660 120
rect 3654 115 3660 116
rect 3798 119 3804 120
rect 3798 115 3799 119
rect 3803 115 3804 119
rect 3838 119 3839 123
rect 3843 119 3844 123
rect 4318 120 4319 124
rect 4323 120 4324 124
rect 4318 119 4324 120
rect 4454 124 4460 125
rect 4454 120 4455 124
rect 4459 120 4460 124
rect 4454 119 4460 120
rect 4590 124 4596 125
rect 4590 120 4591 124
rect 4595 120 4596 124
rect 4590 119 4596 120
rect 4726 124 4732 125
rect 4726 120 4727 124
rect 4731 120 4732 124
rect 4726 119 4732 120
rect 4862 124 4868 125
rect 4862 120 4863 124
rect 4867 120 4868 124
rect 4862 119 4868 120
rect 4998 124 5004 125
rect 4998 120 4999 124
rect 5003 120 5004 124
rect 4998 119 5004 120
rect 5134 124 5140 125
rect 5134 120 5135 124
rect 5139 120 5140 124
rect 5134 119 5140 120
rect 5270 124 5276 125
rect 5270 120 5271 124
rect 5275 120 5276 124
rect 5270 119 5276 120
rect 5406 124 5412 125
rect 5406 120 5407 124
rect 5411 120 5412 124
rect 5406 119 5412 120
rect 5542 124 5548 125
rect 5542 120 5543 124
rect 5547 120 5548 124
rect 5542 119 5548 120
rect 5662 123 5668 124
rect 5662 119 5663 123
rect 5667 119 5668 123
rect 3838 118 3844 119
rect 5662 118 5668 119
rect 1974 114 1980 115
rect 3798 114 3804 115
<< m3c >>
rect 111 5688 115 5692
rect 131 5687 135 5691
rect 267 5687 271 5691
rect 403 5687 407 5691
rect 1935 5688 1939 5692
rect 111 5671 115 5675
rect 159 5672 163 5676
rect 295 5672 299 5676
rect 431 5672 435 5676
rect 1935 5671 1939 5675
rect 1975 5620 1979 5624
rect 1995 5619 1999 5623
rect 2171 5619 2175 5623
rect 2371 5619 2375 5623
rect 2563 5619 2567 5623
rect 2747 5619 2751 5623
rect 2931 5619 2935 5623
rect 3107 5619 3111 5623
rect 3275 5619 3279 5623
rect 3443 5619 3447 5623
rect 3619 5619 3623 5623
rect 3799 5620 3803 5624
rect 3839 5624 3843 5628
rect 4467 5623 4471 5627
rect 4603 5623 4607 5627
rect 4739 5623 4743 5627
rect 4875 5623 4879 5627
rect 5663 5624 5667 5628
rect 111 5613 115 5617
rect 343 5612 347 5616
rect 535 5612 539 5616
rect 735 5612 739 5616
rect 943 5612 947 5616
rect 1159 5612 1163 5616
rect 1383 5612 1387 5616
rect 1607 5612 1611 5616
rect 1815 5612 1819 5616
rect 1935 5613 1939 5617
rect 1975 5603 1979 5607
rect 2023 5604 2027 5608
rect 2199 5604 2203 5608
rect 2399 5604 2403 5608
rect 2591 5604 2595 5608
rect 2775 5604 2779 5608
rect 2959 5604 2963 5608
rect 3135 5604 3139 5608
rect 3303 5604 3307 5608
rect 3471 5604 3475 5608
rect 3647 5604 3651 5608
rect 3799 5603 3803 5607
rect 3839 5607 3843 5611
rect 4495 5608 4499 5612
rect 4631 5608 4635 5612
rect 4767 5608 4771 5612
rect 4903 5608 4907 5612
rect 5663 5607 5667 5611
rect 111 5596 115 5600
rect 315 5597 319 5601
rect 507 5597 511 5601
rect 707 5597 711 5601
rect 915 5597 919 5601
rect 1131 5597 1135 5601
rect 1355 5597 1359 5601
rect 1579 5597 1583 5601
rect 1787 5597 1791 5601
rect 1935 5596 1939 5600
rect 1975 5545 1979 5549
rect 2375 5544 2379 5548
rect 2607 5544 2611 5548
rect 2831 5544 2835 5548
rect 3047 5544 3051 5548
rect 3263 5544 3267 5548
rect 3479 5544 3483 5548
rect 3679 5544 3683 5548
rect 3799 5545 3803 5549
rect 3839 5549 3843 5553
rect 4431 5548 4435 5552
rect 4567 5548 4571 5552
rect 4703 5548 4707 5552
rect 4839 5548 4843 5552
rect 4975 5548 4979 5552
rect 5111 5548 5115 5552
rect 5663 5549 5667 5553
rect 1975 5528 1979 5532
rect 2347 5529 2351 5533
rect 2579 5529 2583 5533
rect 2803 5529 2807 5533
rect 3019 5529 3023 5533
rect 3235 5529 3239 5533
rect 3451 5529 3455 5533
rect 3651 5529 3655 5533
rect 3799 5528 3803 5532
rect 3839 5532 3843 5536
rect 4403 5533 4407 5537
rect 4539 5533 4543 5537
rect 4675 5533 4679 5537
rect 4811 5533 4815 5537
rect 4947 5533 4951 5537
rect 5083 5533 5087 5537
rect 5663 5532 5667 5536
rect 111 5464 115 5468
rect 875 5463 879 5467
rect 1011 5463 1015 5467
rect 1147 5463 1151 5467
rect 1291 5463 1295 5467
rect 1435 5463 1439 5467
rect 1579 5463 1583 5467
rect 1723 5463 1727 5467
rect 1935 5464 1939 5468
rect 111 5447 115 5451
rect 903 5448 907 5452
rect 1039 5448 1043 5452
rect 1175 5448 1179 5452
rect 1319 5448 1323 5452
rect 1463 5448 1467 5452
rect 1607 5448 1611 5452
rect 1751 5448 1755 5452
rect 1935 5447 1939 5451
rect 3839 5400 3843 5404
rect 4427 5399 4431 5403
rect 4587 5399 4591 5403
rect 4747 5399 4751 5403
rect 4907 5399 4911 5403
rect 5075 5399 5079 5403
rect 5663 5400 5667 5404
rect 111 5389 115 5393
rect 719 5388 723 5392
rect 855 5388 859 5392
rect 991 5388 995 5392
rect 1127 5388 1131 5392
rect 1263 5388 1267 5392
rect 1399 5388 1403 5392
rect 1535 5388 1539 5392
rect 1671 5388 1675 5392
rect 1807 5388 1811 5392
rect 1935 5389 1939 5393
rect 1975 5392 1979 5396
rect 2451 5391 2455 5395
rect 2699 5391 2703 5395
rect 2947 5391 2951 5395
rect 3187 5391 3191 5395
rect 3427 5391 3431 5395
rect 3651 5391 3655 5395
rect 3799 5392 3803 5396
rect 3839 5383 3843 5387
rect 4455 5384 4459 5388
rect 4615 5384 4619 5388
rect 4775 5384 4779 5388
rect 4935 5384 4939 5388
rect 5103 5384 5107 5388
rect 5663 5383 5667 5387
rect 111 5372 115 5376
rect 691 5373 695 5377
rect 827 5373 831 5377
rect 963 5373 967 5377
rect 1099 5373 1103 5377
rect 1235 5373 1239 5377
rect 1371 5373 1375 5377
rect 1507 5373 1511 5377
rect 1643 5373 1647 5377
rect 1779 5373 1783 5377
rect 1935 5372 1939 5376
rect 1975 5375 1979 5379
rect 2479 5376 2483 5380
rect 2727 5376 2731 5380
rect 2975 5376 2979 5380
rect 3215 5376 3219 5380
rect 3455 5376 3459 5380
rect 3679 5376 3683 5380
rect 3799 5375 3803 5379
rect 1975 5317 1979 5321
rect 2319 5316 2323 5320
rect 2519 5316 2523 5320
rect 2719 5316 2723 5320
rect 2919 5316 2923 5320
rect 3119 5316 3123 5320
rect 3327 5316 3331 5320
rect 3535 5316 3539 5320
rect 3799 5317 3803 5321
rect 3839 5317 3843 5321
rect 4431 5316 4435 5320
rect 4615 5316 4619 5320
rect 4799 5316 4803 5320
rect 4983 5316 4987 5320
rect 5175 5316 5179 5320
rect 5663 5317 5667 5321
rect 1975 5300 1979 5304
rect 2291 5301 2295 5305
rect 2491 5301 2495 5305
rect 2691 5301 2695 5305
rect 2891 5301 2895 5305
rect 3091 5301 3095 5305
rect 3299 5301 3303 5305
rect 3507 5301 3511 5305
rect 3799 5300 3803 5304
rect 3839 5300 3843 5304
rect 4403 5301 4407 5305
rect 4587 5301 4591 5305
rect 4771 5301 4775 5305
rect 4955 5301 4959 5305
rect 5147 5301 5151 5305
rect 5663 5300 5667 5304
rect 111 5240 115 5244
rect 723 5239 727 5243
rect 875 5239 879 5243
rect 1027 5239 1031 5243
rect 1187 5239 1191 5243
rect 1355 5239 1359 5243
rect 1523 5239 1527 5243
rect 1935 5240 1939 5244
rect 111 5223 115 5227
rect 751 5224 755 5228
rect 903 5224 907 5228
rect 1055 5224 1059 5228
rect 1215 5224 1219 5228
rect 1383 5224 1387 5228
rect 1551 5224 1555 5228
rect 1935 5223 1939 5227
rect 111 5165 115 5169
rect 447 5164 451 5168
rect 623 5164 627 5168
rect 807 5164 811 5168
rect 999 5164 1003 5168
rect 1199 5164 1203 5168
rect 1399 5164 1403 5168
rect 1607 5164 1611 5168
rect 1815 5164 1819 5168
rect 1935 5165 1939 5169
rect 1975 5164 1979 5168
rect 2275 5163 2279 5167
rect 2475 5163 2479 5167
rect 2683 5163 2687 5167
rect 2891 5163 2895 5167
rect 3099 5163 3103 5167
rect 3307 5163 3311 5167
rect 3799 5164 3803 5168
rect 111 5148 115 5152
rect 419 5149 423 5153
rect 595 5149 599 5153
rect 779 5149 783 5153
rect 971 5149 975 5153
rect 1171 5149 1175 5153
rect 1371 5149 1375 5153
rect 1579 5149 1583 5153
rect 1787 5149 1791 5153
rect 1935 5148 1939 5152
rect 1975 5147 1979 5151
rect 2303 5148 2307 5152
rect 2503 5148 2507 5152
rect 2711 5148 2715 5152
rect 2919 5148 2923 5152
rect 3127 5148 3131 5152
rect 3839 5152 3843 5156
rect 3335 5148 3339 5152
rect 4435 5151 4439 5155
rect 3799 5147 3803 5151
rect 4595 5151 4599 5155
rect 4755 5151 4759 5155
rect 4915 5151 4919 5155
rect 5067 5151 5071 5155
rect 5219 5151 5223 5155
rect 5379 5151 5383 5155
rect 5515 5151 5519 5155
rect 5663 5152 5667 5156
rect 3839 5135 3843 5139
rect 4463 5136 4467 5140
rect 4623 5136 4627 5140
rect 4783 5136 4787 5140
rect 4943 5136 4947 5140
rect 5095 5136 5099 5140
rect 5247 5136 5251 5140
rect 5407 5136 5411 5140
rect 5543 5136 5547 5140
rect 5663 5135 5667 5139
rect 1975 5073 1979 5077
rect 2119 5072 2123 5076
rect 2327 5072 2331 5076
rect 2535 5072 2539 5076
rect 2751 5072 2755 5076
rect 2975 5072 2979 5076
rect 3207 5072 3211 5076
rect 3799 5073 3803 5077
rect 3839 5069 3843 5073
rect 3887 5068 3891 5072
rect 4087 5068 4091 5072
rect 4327 5068 4331 5072
rect 4567 5068 4571 5072
rect 4815 5068 4819 5072
rect 5063 5068 5067 5072
rect 5311 5068 5315 5072
rect 5543 5068 5547 5072
rect 5663 5069 5667 5073
rect 1975 5056 1979 5060
rect 2091 5057 2095 5061
rect 2299 5057 2303 5061
rect 2507 5057 2511 5061
rect 2723 5057 2727 5061
rect 2947 5057 2951 5061
rect 3179 5057 3183 5061
rect 3799 5056 3803 5060
rect 3839 5052 3843 5056
rect 3859 5053 3863 5057
rect 4059 5053 4063 5057
rect 4299 5053 4303 5057
rect 4539 5053 4543 5057
rect 4787 5053 4791 5057
rect 5035 5053 5039 5057
rect 5283 5053 5287 5057
rect 5515 5053 5519 5057
rect 5663 5052 5667 5056
rect 111 5008 115 5012
rect 155 5007 159 5011
rect 379 5007 383 5011
rect 627 5007 631 5011
rect 899 5007 903 5011
rect 1195 5007 1199 5011
rect 1499 5007 1503 5011
rect 1787 5007 1791 5011
rect 1935 5008 1939 5012
rect 111 4991 115 4995
rect 183 4992 187 4996
rect 407 4992 411 4996
rect 655 4992 659 4996
rect 927 4992 931 4996
rect 1223 4992 1227 4996
rect 1527 4992 1531 4996
rect 1815 4992 1819 4996
rect 1935 4991 1939 4995
rect 1975 4916 1979 4920
rect 1995 4915 1999 4919
rect 2131 4915 2135 4919
rect 2267 4915 2271 4919
rect 2419 4915 2423 4919
rect 2619 4915 2623 4919
rect 2859 4915 2863 4919
rect 3123 4915 3127 4919
rect 3395 4915 3399 4919
rect 3651 4915 3655 4919
rect 3799 4916 3803 4920
rect 3839 4920 3843 4924
rect 3859 4919 3863 4923
rect 3995 4919 3999 4923
rect 4131 4919 4135 4923
rect 4267 4919 4271 4923
rect 4403 4919 4407 4923
rect 4539 4919 4543 4923
rect 4675 4919 4679 4923
rect 4811 4919 4815 4923
rect 4947 4919 4951 4923
rect 5083 4919 5087 4923
rect 5227 4919 5231 4923
rect 5379 4919 5383 4923
rect 5515 4919 5519 4923
rect 5663 4920 5667 4924
rect 111 4905 115 4909
rect 159 4904 163 4908
rect 295 4904 299 4908
rect 431 4904 435 4908
rect 567 4904 571 4908
rect 703 4904 707 4908
rect 1935 4905 1939 4909
rect 1975 4899 1979 4903
rect 2023 4900 2027 4904
rect 2159 4900 2163 4904
rect 2295 4900 2299 4904
rect 2447 4900 2451 4904
rect 2647 4900 2651 4904
rect 2887 4900 2891 4904
rect 3151 4900 3155 4904
rect 3423 4900 3427 4904
rect 3679 4900 3683 4904
rect 3799 4899 3803 4903
rect 3839 4903 3843 4907
rect 3887 4904 3891 4908
rect 4023 4904 4027 4908
rect 4159 4904 4163 4908
rect 4295 4904 4299 4908
rect 4431 4904 4435 4908
rect 4567 4904 4571 4908
rect 4703 4904 4707 4908
rect 4839 4904 4843 4908
rect 4975 4904 4979 4908
rect 5111 4904 5115 4908
rect 5255 4904 5259 4908
rect 5407 4904 5411 4908
rect 5543 4904 5547 4908
rect 5663 4903 5667 4907
rect 111 4888 115 4892
rect 131 4889 135 4893
rect 267 4889 271 4893
rect 403 4889 407 4893
rect 539 4889 543 4893
rect 675 4889 679 4893
rect 1935 4888 1939 4892
rect 1975 4833 1979 4837
rect 2327 4832 2331 4836
rect 2559 4832 2563 4836
rect 2823 4832 2827 4836
rect 3103 4832 3107 4836
rect 3399 4832 3403 4836
rect 3679 4832 3683 4836
rect 3799 4833 3803 4837
rect 1975 4816 1979 4820
rect 2299 4817 2303 4821
rect 2531 4817 2535 4821
rect 2795 4817 2799 4821
rect 3075 4817 3079 4821
rect 3371 4817 3375 4821
rect 3651 4817 3655 4821
rect 3799 4816 3803 4820
rect 3839 4769 3843 4773
rect 3887 4768 3891 4772
rect 4071 4768 4075 4772
rect 4295 4768 4299 4772
rect 4535 4768 4539 4772
rect 4783 4768 4787 4772
rect 5039 4768 5043 4772
rect 5303 4768 5307 4772
rect 5543 4768 5547 4772
rect 5663 4769 5667 4773
rect 3839 4752 3843 4756
rect 3859 4753 3863 4757
rect 4043 4753 4047 4757
rect 4267 4753 4271 4757
rect 4507 4753 4511 4757
rect 4755 4753 4759 4757
rect 5011 4753 5015 4757
rect 5275 4753 5279 4757
rect 5515 4753 5519 4757
rect 5663 4752 5667 4756
rect 111 4744 115 4748
rect 131 4743 135 4747
rect 267 4743 271 4747
rect 403 4743 407 4747
rect 539 4743 543 4747
rect 675 4743 679 4747
rect 1935 4744 1939 4748
rect 111 4727 115 4731
rect 159 4728 163 4732
rect 295 4728 299 4732
rect 431 4728 435 4732
rect 567 4728 571 4732
rect 703 4728 707 4732
rect 1935 4727 1939 4731
rect 1975 4672 1979 4676
rect 2019 4671 2023 4675
rect 2195 4671 2199 4675
rect 2371 4671 2375 4675
rect 2547 4671 2551 4675
rect 2723 4671 2727 4675
rect 3799 4672 3803 4676
rect 111 4665 115 4669
rect 159 4664 163 4668
rect 295 4664 299 4668
rect 431 4664 435 4668
rect 567 4664 571 4668
rect 703 4664 707 4668
rect 1935 4665 1939 4669
rect 1975 4655 1979 4659
rect 2047 4656 2051 4660
rect 2223 4656 2227 4660
rect 2399 4656 2403 4660
rect 2575 4656 2579 4660
rect 2751 4656 2755 4660
rect 3799 4655 3803 4659
rect 111 4648 115 4652
rect 131 4649 135 4653
rect 267 4649 271 4653
rect 403 4649 407 4653
rect 539 4649 543 4653
rect 675 4649 679 4653
rect 1935 4648 1939 4652
rect 3839 4620 3843 4624
rect 3859 4619 3863 4623
rect 3995 4619 3999 4623
rect 4131 4619 4135 4623
rect 4267 4619 4271 4623
rect 4403 4619 4407 4623
rect 4539 4619 4543 4623
rect 4675 4619 4679 4623
rect 4819 4619 4823 4623
rect 4963 4619 4967 4623
rect 5107 4619 5111 4623
rect 5243 4619 5247 4623
rect 5379 4619 5383 4623
rect 5515 4619 5519 4623
rect 5663 4620 5667 4624
rect 3839 4603 3843 4607
rect 3887 4604 3891 4608
rect 4023 4604 4027 4608
rect 4159 4604 4163 4608
rect 4295 4604 4299 4608
rect 4431 4604 4435 4608
rect 4567 4604 4571 4608
rect 4703 4604 4707 4608
rect 4847 4604 4851 4608
rect 4991 4604 4995 4608
rect 5135 4604 5139 4608
rect 5271 4604 5275 4608
rect 5407 4604 5411 4608
rect 5543 4604 5547 4608
rect 5663 4603 5667 4607
rect 1975 4593 1979 4597
rect 2023 4592 2027 4596
rect 2263 4592 2267 4596
rect 2527 4592 2531 4596
rect 2775 4592 2779 4596
rect 3015 4592 3019 4596
rect 3247 4592 3251 4596
rect 3471 4592 3475 4596
rect 3679 4592 3683 4596
rect 3799 4593 3803 4597
rect 1975 4576 1979 4580
rect 1995 4577 1999 4581
rect 2235 4577 2239 4581
rect 2499 4577 2503 4581
rect 2747 4577 2751 4581
rect 2987 4577 2991 4581
rect 3219 4577 3223 4581
rect 3443 4577 3447 4581
rect 3651 4577 3655 4581
rect 3799 4576 3803 4580
rect 3839 4545 3843 4549
rect 4671 4544 4675 4548
rect 4807 4544 4811 4548
rect 4943 4544 4947 4548
rect 5079 4544 5083 4548
rect 5663 4545 5667 4549
rect 3839 4528 3843 4532
rect 4643 4529 4647 4533
rect 4779 4529 4783 4533
rect 4915 4529 4919 4533
rect 5051 4529 5055 4533
rect 5663 4528 5667 4532
rect 111 4504 115 4508
rect 251 4503 255 4507
rect 443 4503 447 4507
rect 651 4503 655 4507
rect 875 4503 879 4507
rect 1099 4503 1103 4507
rect 1331 4503 1335 4507
rect 1571 4503 1575 4507
rect 1787 4503 1791 4507
rect 1935 4504 1939 4508
rect 111 4487 115 4491
rect 279 4488 283 4492
rect 471 4488 475 4492
rect 679 4488 683 4492
rect 903 4488 907 4492
rect 1127 4488 1131 4492
rect 1359 4488 1363 4492
rect 1599 4488 1603 4492
rect 1815 4488 1819 4492
rect 1935 4487 1939 4491
rect 111 4429 115 4433
rect 511 4428 515 4432
rect 687 4428 691 4432
rect 871 4428 875 4432
rect 1071 4428 1075 4432
rect 1279 4428 1283 4432
rect 1495 4428 1499 4432
rect 1719 4428 1723 4432
rect 1935 4429 1939 4433
rect 1975 4432 1979 4436
rect 2267 4431 2271 4435
rect 2515 4431 2519 4435
rect 2747 4431 2751 4435
rect 2971 4431 2975 4435
rect 3187 4431 3191 4435
rect 3395 4431 3399 4435
rect 3611 4431 3615 4435
rect 3799 4432 3803 4436
rect 111 4412 115 4416
rect 483 4413 487 4417
rect 659 4413 663 4417
rect 843 4413 847 4417
rect 1043 4413 1047 4417
rect 1251 4413 1255 4417
rect 1467 4413 1471 4417
rect 1691 4413 1695 4417
rect 1935 4412 1939 4416
rect 1975 4415 1979 4419
rect 2295 4416 2299 4420
rect 2543 4416 2547 4420
rect 2775 4416 2779 4420
rect 2999 4416 3003 4420
rect 3215 4416 3219 4420
rect 3423 4416 3427 4420
rect 3639 4416 3643 4420
rect 3799 4415 3803 4419
rect 3839 4392 3843 4396
rect 4347 4391 4351 4395
rect 4483 4391 4487 4395
rect 4619 4391 4623 4395
rect 4755 4391 4759 4395
rect 4891 4391 4895 4395
rect 5663 4392 5667 4396
rect 3839 4375 3843 4379
rect 4375 4376 4379 4380
rect 4511 4376 4515 4380
rect 4647 4376 4651 4380
rect 4783 4376 4787 4380
rect 4919 4376 4923 4380
rect 5663 4375 5667 4379
rect 1975 4345 1979 4349
rect 2023 4344 2027 4348
rect 2199 4344 2203 4348
rect 2399 4344 2403 4348
rect 2591 4344 2595 4348
rect 2775 4344 2779 4348
rect 2951 4344 2955 4348
rect 3135 4344 3139 4348
rect 3319 4344 3323 4348
rect 3799 4345 3803 4349
rect 1975 4328 1979 4332
rect 1995 4329 1999 4333
rect 2171 4329 2175 4333
rect 2371 4329 2375 4333
rect 2563 4329 2567 4333
rect 2747 4329 2751 4333
rect 2923 4329 2927 4333
rect 3107 4329 3111 4333
rect 3291 4329 3295 4333
rect 3799 4328 3803 4332
rect 3839 4301 3843 4305
rect 4135 4300 4139 4304
rect 4271 4300 4275 4304
rect 4407 4300 4411 4304
rect 4543 4300 4547 4304
rect 4679 4300 4683 4304
rect 5663 4301 5667 4305
rect 3839 4284 3843 4288
rect 4107 4285 4111 4289
rect 4243 4285 4247 4289
rect 4379 4285 4383 4289
rect 4515 4285 4519 4289
rect 4651 4285 4655 4289
rect 5663 4284 5667 4288
rect 111 4276 115 4280
rect 715 4275 719 4279
rect 851 4275 855 4279
rect 987 4275 991 4279
rect 1123 4275 1127 4279
rect 1259 4275 1263 4279
rect 1395 4275 1399 4279
rect 1531 4275 1535 4279
rect 1667 4275 1671 4279
rect 1935 4276 1939 4280
rect 111 4259 115 4263
rect 743 4260 747 4264
rect 879 4260 883 4264
rect 1015 4260 1019 4264
rect 1151 4260 1155 4264
rect 1287 4260 1291 4264
rect 1423 4260 1427 4264
rect 1559 4260 1563 4264
rect 1695 4260 1699 4264
rect 1935 4259 1939 4263
rect 111 4193 115 4197
rect 727 4192 731 4196
rect 863 4192 867 4196
rect 999 4192 1003 4196
rect 1135 4192 1139 4196
rect 1271 4192 1275 4196
rect 1407 4192 1411 4196
rect 1543 4192 1547 4196
rect 1679 4192 1683 4196
rect 1815 4192 1819 4196
rect 1935 4193 1939 4197
rect 1975 4192 1979 4196
rect 1995 4191 1999 4195
rect 2243 4191 2247 4195
rect 2507 4191 2511 4195
rect 2763 4191 2767 4195
rect 3019 4191 3023 4195
rect 3283 4191 3287 4195
rect 3799 4192 3803 4196
rect 111 4176 115 4180
rect 699 4177 703 4181
rect 835 4177 839 4181
rect 971 4177 975 4181
rect 1107 4177 1111 4181
rect 1243 4177 1247 4181
rect 1379 4177 1383 4181
rect 1515 4177 1519 4181
rect 1651 4177 1655 4181
rect 1787 4177 1791 4181
rect 1935 4176 1939 4180
rect 1975 4175 1979 4179
rect 2023 4176 2027 4180
rect 2271 4176 2275 4180
rect 2535 4176 2539 4180
rect 2791 4176 2795 4180
rect 3047 4176 3051 4180
rect 3311 4176 3315 4180
rect 3799 4175 3803 4179
rect 3839 4140 3843 4144
rect 3971 4139 3975 4143
rect 4107 4139 4111 4143
rect 4243 4139 4247 4143
rect 4379 4139 4383 4143
rect 4515 4139 4519 4143
rect 5663 4140 5667 4144
rect 3839 4123 3843 4127
rect 3999 4124 4003 4128
rect 4135 4124 4139 4128
rect 4271 4124 4275 4128
rect 4407 4124 4411 4128
rect 4543 4124 4547 4128
rect 5663 4123 5667 4127
rect 1975 4105 1979 4109
rect 3135 4104 3139 4108
rect 3271 4104 3275 4108
rect 3407 4104 3411 4108
rect 3543 4104 3547 4108
rect 3679 4104 3683 4108
rect 3799 4105 3803 4109
rect 1975 4088 1979 4092
rect 3107 4089 3111 4093
rect 3243 4089 3247 4093
rect 3379 4089 3383 4093
rect 3515 4089 3519 4093
rect 3651 4089 3655 4093
rect 3799 4088 3803 4092
rect 111 4044 115 4048
rect 563 4043 567 4047
rect 699 4043 703 4047
rect 835 4043 839 4047
rect 971 4043 975 4047
rect 1107 4043 1111 4047
rect 1243 4043 1247 4047
rect 1379 4043 1383 4047
rect 1515 4043 1519 4047
rect 1651 4043 1655 4047
rect 1787 4043 1791 4047
rect 1935 4044 1939 4048
rect 3839 4041 3843 4045
rect 3887 4040 3891 4044
rect 4023 4040 4027 4044
rect 4159 4040 4163 4044
rect 4295 4040 4299 4044
rect 4431 4040 4435 4044
rect 4567 4040 4571 4044
rect 4703 4040 4707 4044
rect 4839 4040 4843 4044
rect 5663 4041 5667 4045
rect 111 4027 115 4031
rect 591 4028 595 4032
rect 727 4028 731 4032
rect 863 4028 867 4032
rect 999 4028 1003 4032
rect 1135 4028 1139 4032
rect 1271 4028 1275 4032
rect 1407 4028 1411 4032
rect 1543 4028 1547 4032
rect 1679 4028 1683 4032
rect 1815 4028 1819 4032
rect 1935 4027 1939 4031
rect 3839 4024 3843 4028
rect 3859 4025 3863 4029
rect 3995 4025 3999 4029
rect 4131 4025 4135 4029
rect 4267 4025 4271 4029
rect 4403 4025 4407 4029
rect 4539 4025 4543 4029
rect 4675 4025 4679 4029
rect 4811 4025 4815 4029
rect 5663 4024 5667 4028
rect 111 3969 115 3973
rect 159 3968 163 3972
rect 327 3968 331 3972
rect 535 3968 539 3972
rect 751 3968 755 3972
rect 967 3968 971 3972
rect 1183 3968 1187 3972
rect 1399 3968 1403 3972
rect 1615 3968 1619 3972
rect 1815 3968 1819 3972
rect 1935 3969 1939 3973
rect 111 3952 115 3956
rect 131 3953 135 3957
rect 299 3953 303 3957
rect 507 3953 511 3957
rect 723 3953 727 3957
rect 939 3953 943 3957
rect 1155 3953 1159 3957
rect 1371 3953 1375 3957
rect 1587 3953 1591 3957
rect 1787 3953 1791 3957
rect 1935 3952 1939 3956
rect 3839 3892 3843 3896
rect 3859 3891 3863 3895
rect 3995 3891 3999 3895
rect 4147 3891 4151 3895
rect 4299 3891 4303 3895
rect 4459 3891 4463 3895
rect 4619 3891 4623 3895
rect 4779 3891 4783 3895
rect 5663 3892 5667 3896
rect 3839 3875 3843 3879
rect 3887 3876 3891 3880
rect 4023 3876 4027 3880
rect 4175 3876 4179 3880
rect 4327 3876 4331 3880
rect 4487 3876 4491 3880
rect 4647 3876 4651 3880
rect 4807 3876 4811 3880
rect 5663 3875 5667 3879
rect 1975 3864 1979 3868
rect 1995 3863 1999 3867
rect 2403 3863 2407 3867
rect 2827 3863 2831 3867
rect 3251 3863 3255 3867
rect 3651 3863 3655 3867
rect 3799 3864 3803 3868
rect 1975 3847 1979 3851
rect 2023 3848 2027 3852
rect 2431 3848 2435 3852
rect 2855 3848 2859 3852
rect 3279 3848 3283 3852
rect 3679 3848 3683 3852
rect 3799 3847 3803 3851
rect 111 3820 115 3824
rect 131 3819 135 3823
rect 355 3819 359 3823
rect 619 3819 623 3823
rect 899 3819 903 3823
rect 1195 3819 1199 3823
rect 1499 3819 1503 3823
rect 1787 3819 1791 3823
rect 1935 3820 1939 3824
rect 111 3803 115 3807
rect 159 3804 163 3808
rect 383 3804 387 3808
rect 647 3804 651 3808
rect 927 3804 931 3808
rect 1223 3804 1227 3808
rect 1527 3804 1531 3808
rect 1815 3804 1819 3808
rect 1935 3803 1939 3807
rect 1975 3789 1979 3793
rect 2023 3788 2027 3792
rect 2175 3788 2179 3792
rect 2351 3788 2355 3792
rect 2535 3788 2539 3792
rect 2719 3788 2723 3792
rect 2895 3788 2899 3792
rect 3071 3788 3075 3792
rect 3247 3788 3251 3792
rect 3423 3788 3427 3792
rect 3607 3788 3611 3792
rect 3799 3789 3803 3793
rect 3839 3789 3843 3793
rect 4503 3788 4507 3792
rect 4639 3788 4643 3792
rect 4775 3788 4779 3792
rect 4911 3788 4915 3792
rect 5047 3788 5051 3792
rect 5663 3789 5667 3793
rect 1975 3772 1979 3776
rect 1995 3773 1999 3777
rect 2147 3773 2151 3777
rect 2323 3773 2327 3777
rect 2507 3773 2511 3777
rect 2691 3773 2695 3777
rect 2867 3773 2871 3777
rect 3043 3773 3047 3777
rect 3219 3773 3223 3777
rect 3395 3773 3399 3777
rect 3579 3773 3583 3777
rect 3799 3772 3803 3776
rect 3839 3772 3843 3776
rect 4475 3773 4479 3777
rect 4611 3773 4615 3777
rect 4747 3773 4751 3777
rect 4883 3773 4887 3777
rect 5019 3773 5023 3777
rect 5663 3772 5667 3776
rect 111 3733 115 3737
rect 247 3732 251 3736
rect 519 3732 523 3736
rect 791 3732 795 3736
rect 1063 3732 1067 3736
rect 1343 3732 1347 3736
rect 1935 3733 1939 3737
rect 111 3716 115 3720
rect 219 3717 223 3721
rect 491 3717 495 3721
rect 763 3717 767 3721
rect 1035 3717 1039 3721
rect 1315 3717 1319 3721
rect 1935 3716 1939 3720
rect 1975 3632 1979 3636
rect 2011 3631 2015 3635
rect 2147 3631 2151 3635
rect 2291 3631 2295 3635
rect 2435 3631 2439 3635
rect 2579 3631 2583 3635
rect 2723 3631 2727 3635
rect 2867 3631 2871 3635
rect 3011 3631 3015 3635
rect 3155 3631 3159 3635
rect 3299 3631 3303 3635
rect 3799 3632 3803 3636
rect 1975 3615 1979 3619
rect 2039 3616 2043 3620
rect 2175 3616 2179 3620
rect 2319 3616 2323 3620
rect 2463 3616 2467 3620
rect 2607 3616 2611 3620
rect 2751 3616 2755 3620
rect 2895 3616 2899 3620
rect 3039 3616 3043 3620
rect 3183 3616 3187 3620
rect 3839 3620 3843 3624
rect 3327 3616 3331 3620
rect 4019 3619 4023 3623
rect 3799 3615 3803 3619
rect 4155 3619 4159 3623
rect 4291 3619 4295 3623
rect 4427 3619 4431 3623
rect 4563 3619 4567 3623
rect 4699 3619 4703 3623
rect 4835 3619 4839 3623
rect 4971 3619 4975 3623
rect 5107 3619 5111 3623
rect 5243 3619 5247 3623
rect 5379 3619 5383 3623
rect 5515 3619 5519 3623
rect 5663 3620 5667 3624
rect 3839 3603 3843 3607
rect 4047 3604 4051 3608
rect 4183 3604 4187 3608
rect 4319 3604 4323 3608
rect 4455 3604 4459 3608
rect 4591 3604 4595 3608
rect 4727 3604 4731 3608
rect 4863 3604 4867 3608
rect 4999 3604 5003 3608
rect 5135 3604 5139 3608
rect 5271 3604 5275 3608
rect 5407 3604 5411 3608
rect 5543 3604 5547 3608
rect 5663 3603 5667 3607
rect 111 3568 115 3572
rect 491 3567 495 3571
rect 635 3567 639 3571
rect 779 3567 783 3571
rect 923 3567 927 3571
rect 1067 3567 1071 3571
rect 1211 3567 1215 3571
rect 1935 3568 1939 3572
rect 111 3551 115 3555
rect 519 3552 523 3556
rect 663 3552 667 3556
rect 807 3552 811 3556
rect 951 3552 955 3556
rect 1095 3552 1099 3556
rect 1239 3552 1243 3556
rect 1935 3551 1939 3555
rect 1975 3549 1979 3553
rect 2239 3548 2243 3552
rect 2375 3548 2379 3552
rect 2511 3548 2515 3552
rect 2647 3548 2651 3552
rect 2783 3548 2787 3552
rect 2919 3548 2923 3552
rect 3055 3548 3059 3552
rect 3191 3548 3195 3552
rect 3327 3548 3331 3552
rect 3463 3548 3467 3552
rect 3799 3549 3803 3553
rect 1975 3532 1979 3536
rect 2211 3533 2215 3537
rect 2347 3533 2351 3537
rect 2483 3533 2487 3537
rect 2619 3533 2623 3537
rect 2755 3533 2759 3537
rect 2891 3533 2895 3537
rect 3027 3533 3031 3537
rect 3163 3533 3167 3537
rect 3299 3533 3303 3537
rect 3435 3533 3439 3537
rect 3799 3532 3803 3536
rect 3839 3497 3843 3501
rect 5407 3496 5411 3500
rect 5543 3496 5547 3500
rect 5663 3497 5667 3501
rect 3839 3480 3843 3484
rect 5379 3481 5383 3485
rect 5515 3481 5519 3485
rect 5663 3480 5667 3484
rect 111 3473 115 3477
rect 431 3472 435 3476
rect 567 3472 571 3476
rect 703 3472 707 3476
rect 839 3472 843 3476
rect 975 3472 979 3476
rect 1935 3473 1939 3477
rect 111 3456 115 3460
rect 403 3457 407 3461
rect 539 3457 543 3461
rect 675 3457 679 3461
rect 811 3457 815 3461
rect 947 3457 951 3461
rect 1935 3456 1939 3460
rect 1975 3396 1979 3400
rect 2171 3395 2175 3399
rect 2347 3395 2351 3399
rect 2531 3395 2535 3399
rect 2715 3395 2719 3399
rect 2907 3395 2911 3399
rect 3099 3395 3103 3399
rect 3291 3395 3295 3399
rect 3483 3395 3487 3399
rect 3651 3395 3655 3399
rect 3799 3396 3803 3400
rect 1975 3379 1979 3383
rect 2199 3380 2203 3384
rect 2375 3380 2379 3384
rect 2559 3380 2563 3384
rect 2743 3380 2747 3384
rect 2935 3380 2939 3384
rect 3127 3380 3131 3384
rect 3319 3380 3323 3384
rect 3511 3380 3515 3384
rect 3679 3380 3683 3384
rect 3799 3379 3803 3383
rect 3839 3340 3843 3344
rect 3859 3339 3863 3343
rect 4099 3339 4103 3343
rect 4347 3339 4351 3343
rect 4587 3339 4591 3343
rect 4811 3339 4815 3343
rect 5027 3339 5031 3343
rect 5235 3339 5239 3343
rect 5451 3339 5455 3343
rect 5663 3340 5667 3344
rect 3839 3323 3843 3327
rect 3887 3324 3891 3328
rect 4127 3324 4131 3328
rect 4375 3324 4379 3328
rect 4615 3324 4619 3328
rect 4839 3324 4843 3328
rect 5055 3324 5059 3328
rect 5263 3324 5267 3328
rect 5479 3324 5483 3328
rect 5663 3323 5667 3327
rect 111 3316 115 3320
rect 323 3315 327 3319
rect 459 3315 463 3319
rect 595 3315 599 3319
rect 731 3315 735 3319
rect 867 3315 871 3319
rect 1935 3316 1939 3320
rect 111 3299 115 3303
rect 351 3300 355 3304
rect 487 3300 491 3304
rect 623 3300 627 3304
rect 759 3300 763 3304
rect 895 3300 899 3304
rect 1935 3299 1939 3303
rect 1975 3297 1979 3301
rect 2151 3296 2155 3300
rect 2399 3296 2403 3300
rect 2687 3296 2691 3300
rect 3015 3296 3019 3300
rect 3359 3296 3363 3300
rect 3679 3296 3683 3300
rect 3799 3297 3803 3301
rect 1975 3280 1979 3284
rect 2123 3281 2127 3285
rect 2371 3281 2375 3285
rect 2659 3281 2663 3285
rect 2987 3281 2991 3285
rect 3331 3281 3335 3285
rect 3651 3281 3655 3285
rect 3799 3280 3803 3284
rect 3839 3265 3843 3269
rect 3887 3264 3891 3268
rect 4127 3264 4131 3268
rect 4375 3264 4379 3268
rect 4607 3264 4611 3268
rect 4815 3264 4819 3268
rect 5015 3264 5019 3268
rect 5199 3264 5203 3268
rect 5383 3264 5387 3268
rect 5543 3264 5547 3268
rect 5663 3265 5667 3269
rect 3839 3248 3843 3252
rect 3859 3249 3863 3253
rect 4099 3249 4103 3253
rect 4347 3249 4351 3253
rect 4579 3249 4583 3253
rect 4787 3249 4791 3253
rect 4987 3249 4991 3253
rect 5171 3249 5175 3253
rect 5355 3249 5359 3253
rect 5515 3249 5519 3253
rect 5663 3248 5667 3252
rect 111 3233 115 3237
rect 159 3232 163 3236
rect 335 3232 339 3236
rect 543 3232 547 3236
rect 751 3232 755 3236
rect 959 3232 963 3236
rect 1935 3233 1939 3237
rect 111 3216 115 3220
rect 131 3217 135 3221
rect 307 3217 311 3221
rect 515 3217 519 3221
rect 723 3217 727 3221
rect 931 3217 935 3221
rect 1935 3216 1939 3220
rect 1975 3148 1979 3152
rect 1995 3147 1999 3151
rect 2147 3147 2151 3151
rect 2347 3147 2351 3151
rect 2555 3147 2559 3151
rect 2771 3147 2775 3151
rect 2987 3147 2991 3151
rect 3211 3147 3215 3151
rect 3443 3147 3447 3151
rect 3651 3147 3655 3151
rect 3799 3148 3803 3152
rect 1975 3131 1979 3135
rect 2023 3132 2027 3136
rect 2175 3132 2179 3136
rect 2375 3132 2379 3136
rect 2583 3132 2587 3136
rect 2799 3132 2803 3136
rect 3015 3132 3019 3136
rect 3239 3132 3243 3136
rect 3471 3132 3475 3136
rect 3679 3132 3683 3136
rect 3799 3131 3803 3135
rect 3839 3100 3843 3104
rect 4467 3099 4471 3103
rect 4651 3099 4655 3103
rect 4859 3099 4863 3103
rect 5075 3099 5079 3103
rect 5307 3099 5311 3103
rect 5515 3099 5519 3103
rect 5663 3100 5667 3104
rect 3839 3083 3843 3087
rect 4495 3084 4499 3088
rect 4679 3084 4683 3088
rect 4887 3084 4891 3088
rect 5103 3084 5107 3088
rect 5335 3084 5339 3088
rect 5543 3084 5547 3088
rect 5663 3083 5667 3087
rect 1975 3073 1979 3077
rect 2647 3072 2651 3076
rect 111 3068 115 3072
rect 131 3067 135 3071
rect 371 3067 375 3071
rect 627 3067 631 3071
rect 875 3067 879 3071
rect 1115 3067 1119 3071
rect 1347 3067 1351 3071
rect 1579 3067 1583 3071
rect 1787 3067 1791 3071
rect 1935 3068 1939 3072
rect 2783 3072 2787 3076
rect 2927 3072 2931 3076
rect 3079 3072 3083 3076
rect 3239 3072 3243 3076
rect 3399 3072 3403 3076
rect 3567 3072 3571 3076
rect 3799 3073 3803 3077
rect 111 3051 115 3055
rect 159 3052 163 3056
rect 399 3052 403 3056
rect 655 3052 659 3056
rect 903 3052 907 3056
rect 1143 3052 1147 3056
rect 1375 3052 1379 3056
rect 1607 3052 1611 3056
rect 1975 3056 1979 3060
rect 2619 3057 2623 3061
rect 2755 3057 2759 3061
rect 2899 3057 2903 3061
rect 3051 3057 3055 3061
rect 3211 3057 3215 3061
rect 3371 3057 3375 3061
rect 3539 3057 3543 3061
rect 3799 3056 3803 3060
rect 1815 3052 1819 3056
rect 1935 3051 1939 3055
rect 3839 3025 3843 3029
rect 4255 3024 4259 3028
rect 4455 3024 4459 3028
rect 4671 3024 4675 3028
rect 4911 3024 4915 3028
rect 5167 3024 5171 3028
rect 5423 3024 5427 3028
rect 5663 3025 5667 3029
rect 3839 3008 3843 3012
rect 4227 3009 4231 3013
rect 4427 3009 4431 3013
rect 4643 3009 4647 3013
rect 4883 3009 4887 3013
rect 5139 3009 5143 3013
rect 5395 3009 5399 3013
rect 5663 3008 5667 3012
rect 111 2993 115 2997
rect 175 2992 179 2996
rect 407 2992 411 2996
rect 623 2992 627 2996
rect 823 2992 827 2996
rect 1007 2992 1011 2996
rect 1183 2992 1187 2996
rect 1351 2992 1355 2996
rect 1511 2992 1515 2996
rect 1671 2992 1675 2996
rect 1815 2992 1819 2996
rect 1935 2993 1939 2997
rect 111 2976 115 2980
rect 147 2977 151 2981
rect 379 2977 383 2981
rect 595 2977 599 2981
rect 795 2977 799 2981
rect 979 2977 983 2981
rect 1155 2977 1159 2981
rect 1323 2977 1327 2981
rect 1483 2977 1487 2981
rect 1643 2977 1647 2981
rect 1787 2977 1791 2981
rect 1935 2976 1939 2980
rect 1975 2924 1979 2928
rect 2803 2923 2807 2927
rect 2939 2923 2943 2927
rect 3075 2923 3079 2927
rect 3211 2923 3215 2927
rect 3347 2923 3351 2927
rect 3483 2923 3487 2927
rect 3799 2924 3803 2928
rect 1975 2907 1979 2911
rect 2831 2908 2835 2912
rect 2967 2908 2971 2912
rect 3103 2908 3107 2912
rect 3239 2908 3243 2912
rect 3375 2908 3379 2912
rect 3511 2908 3515 2912
rect 3799 2907 3803 2911
rect 3839 2852 3843 2856
rect 3995 2851 3999 2855
rect 4211 2851 4215 2855
rect 4443 2851 4447 2855
rect 4699 2851 4703 2855
rect 4971 2851 4975 2855
rect 5251 2851 5255 2855
rect 5515 2851 5519 2855
rect 5663 2852 5667 2856
rect 111 2840 115 2844
rect 395 2839 399 2843
rect 595 2839 599 2843
rect 787 2839 791 2843
rect 971 2839 975 2843
rect 1147 2839 1151 2843
rect 1315 2839 1319 2843
rect 1483 2839 1487 2843
rect 1643 2839 1647 2843
rect 1787 2839 1791 2843
rect 1935 2840 1939 2844
rect 3839 2835 3843 2839
rect 4023 2836 4027 2840
rect 4239 2836 4243 2840
rect 4471 2836 4475 2840
rect 4727 2836 4731 2840
rect 4999 2836 5003 2840
rect 5279 2836 5283 2840
rect 5543 2836 5547 2840
rect 5663 2835 5667 2839
rect 111 2823 115 2827
rect 423 2824 427 2828
rect 623 2824 627 2828
rect 815 2824 819 2828
rect 999 2824 1003 2828
rect 1175 2824 1179 2828
rect 1343 2824 1347 2828
rect 1511 2824 1515 2828
rect 1671 2824 1675 2828
rect 1815 2824 1819 2828
rect 1935 2823 1939 2827
rect 1975 2797 1979 2801
rect 2023 2796 2027 2800
rect 2167 2796 2171 2800
rect 2335 2796 2339 2800
rect 2495 2796 2499 2800
rect 2663 2796 2667 2800
rect 2831 2796 2835 2800
rect 2999 2796 3003 2800
rect 3167 2796 3171 2800
rect 3799 2797 3803 2801
rect 1975 2780 1979 2784
rect 1995 2781 1999 2785
rect 2139 2781 2143 2785
rect 2307 2781 2311 2785
rect 2467 2781 2471 2785
rect 2635 2781 2639 2785
rect 2803 2781 2807 2785
rect 2971 2781 2975 2785
rect 3139 2781 3143 2785
rect 3799 2780 3803 2784
rect 3839 2773 3843 2777
rect 3919 2772 3923 2776
rect 4055 2772 4059 2776
rect 4191 2772 4195 2776
rect 4327 2772 4331 2776
rect 4463 2772 4467 2776
rect 5663 2773 5667 2777
rect 111 2753 115 2757
rect 655 2752 659 2756
rect 815 2752 819 2756
rect 975 2752 979 2756
rect 1143 2752 1147 2756
rect 1311 2752 1315 2756
rect 1479 2752 1483 2756
rect 1935 2753 1939 2757
rect 3839 2756 3843 2760
rect 3891 2757 3895 2761
rect 4027 2757 4031 2761
rect 4163 2757 4167 2761
rect 4299 2757 4303 2761
rect 4435 2757 4439 2761
rect 5663 2756 5667 2760
rect 111 2736 115 2740
rect 627 2737 631 2741
rect 787 2737 791 2741
rect 947 2737 951 2741
rect 1115 2737 1119 2741
rect 1283 2737 1287 2741
rect 1451 2737 1455 2741
rect 1935 2736 1939 2740
rect 1975 2648 1979 2652
rect 2379 2647 2383 2651
rect 2515 2647 2519 2651
rect 2659 2647 2663 2651
rect 2803 2647 2807 2651
rect 2947 2647 2951 2651
rect 3091 2647 3095 2651
rect 3235 2647 3239 2651
rect 3799 2648 3803 2652
rect 1975 2631 1979 2635
rect 2407 2632 2411 2636
rect 2543 2632 2547 2636
rect 2687 2632 2691 2636
rect 2831 2632 2835 2636
rect 2975 2632 2979 2636
rect 3119 2632 3123 2636
rect 3263 2632 3267 2636
rect 3799 2631 3803 2635
rect 3839 2612 3843 2616
rect 4099 2611 4103 2615
rect 4299 2611 4303 2615
rect 4515 2611 4519 2615
rect 4755 2611 4759 2615
rect 5011 2611 5015 2615
rect 5275 2611 5279 2615
rect 5515 2611 5519 2615
rect 5663 2612 5667 2616
rect 111 2604 115 2608
rect 771 2603 775 2607
rect 907 2603 911 2607
rect 1043 2603 1047 2607
rect 1179 2603 1183 2607
rect 1315 2603 1319 2607
rect 1451 2603 1455 2607
rect 1587 2603 1591 2607
rect 1723 2603 1727 2607
rect 1935 2604 1939 2608
rect 3839 2595 3843 2599
rect 4127 2596 4131 2600
rect 4327 2596 4331 2600
rect 4543 2596 4547 2600
rect 4783 2596 4787 2600
rect 5039 2596 5043 2600
rect 5303 2596 5307 2600
rect 5543 2596 5547 2600
rect 5663 2595 5667 2599
rect 111 2587 115 2591
rect 799 2588 803 2592
rect 935 2588 939 2592
rect 1071 2588 1075 2592
rect 1207 2588 1211 2592
rect 1343 2588 1347 2592
rect 1479 2588 1483 2592
rect 1615 2588 1619 2592
rect 1751 2588 1755 2592
rect 1935 2587 1939 2591
rect 1975 2569 1979 2573
rect 2511 2568 2515 2572
rect 2647 2568 2651 2572
rect 2783 2568 2787 2572
rect 2919 2568 2923 2572
rect 3055 2568 3059 2572
rect 3191 2568 3195 2572
rect 3327 2568 3331 2572
rect 3463 2568 3467 2572
rect 3799 2569 3803 2573
rect 1975 2552 1979 2556
rect 2483 2553 2487 2557
rect 2619 2553 2623 2557
rect 2755 2553 2759 2557
rect 2891 2553 2895 2557
rect 3027 2553 3031 2557
rect 3163 2553 3167 2557
rect 3299 2553 3303 2557
rect 3435 2553 3439 2557
rect 3799 2552 3803 2556
rect 3839 2533 3843 2537
rect 4495 2532 4499 2536
rect 4631 2532 4635 2536
rect 4767 2532 4771 2536
rect 4903 2532 4907 2536
rect 5039 2532 5043 2536
rect 5663 2533 5667 2537
rect 111 2513 115 2517
rect 551 2512 555 2516
rect 687 2512 691 2516
rect 831 2512 835 2516
rect 983 2512 987 2516
rect 1135 2512 1139 2516
rect 1295 2512 1299 2516
rect 1455 2512 1459 2516
rect 1615 2512 1619 2516
rect 1783 2512 1787 2516
rect 1935 2513 1939 2517
rect 3839 2516 3843 2520
rect 4467 2517 4471 2521
rect 4603 2517 4607 2521
rect 4739 2517 4743 2521
rect 4875 2517 4879 2521
rect 5011 2517 5015 2521
rect 5663 2516 5667 2520
rect 111 2496 115 2500
rect 523 2497 527 2501
rect 659 2497 663 2501
rect 803 2497 807 2501
rect 955 2497 959 2501
rect 1107 2497 1111 2501
rect 1267 2497 1271 2501
rect 1427 2497 1431 2501
rect 1587 2497 1591 2501
rect 1755 2497 1759 2501
rect 1935 2496 1939 2500
rect 1975 2404 1979 2408
rect 2307 2403 2311 2407
rect 2515 2403 2519 2407
rect 2715 2403 2719 2407
rect 2907 2403 2911 2407
rect 3099 2403 3103 2407
rect 3283 2403 3287 2407
rect 3467 2403 3471 2407
rect 3651 2403 3655 2407
rect 3799 2404 3803 2408
rect 1975 2387 1979 2391
rect 2335 2388 2339 2392
rect 2543 2388 2547 2392
rect 2743 2388 2747 2392
rect 2935 2388 2939 2392
rect 3127 2388 3131 2392
rect 3311 2388 3315 2392
rect 3495 2388 3499 2392
rect 3679 2388 3683 2392
rect 3799 2387 3803 2391
rect 3839 2368 3843 2372
rect 4699 2367 4703 2371
rect 4835 2367 4839 2371
rect 4971 2367 4975 2371
rect 5107 2367 5111 2371
rect 5243 2367 5247 2371
rect 5379 2367 5383 2371
rect 5515 2367 5519 2371
rect 5663 2368 5667 2372
rect 111 2352 115 2356
rect 131 2351 135 2355
rect 339 2351 343 2355
rect 563 2351 567 2355
rect 803 2351 807 2355
rect 1043 2351 1047 2355
rect 1291 2351 1295 2355
rect 1547 2351 1551 2355
rect 1787 2351 1791 2355
rect 1935 2352 1939 2356
rect 3839 2351 3843 2355
rect 4727 2352 4731 2356
rect 4863 2352 4867 2356
rect 4999 2352 5003 2356
rect 5135 2352 5139 2356
rect 5271 2352 5275 2356
rect 5407 2352 5411 2356
rect 5543 2352 5547 2356
rect 5663 2351 5667 2355
rect 111 2335 115 2339
rect 159 2336 163 2340
rect 367 2336 371 2340
rect 591 2336 595 2340
rect 831 2336 835 2340
rect 1071 2336 1075 2340
rect 1319 2336 1323 2340
rect 1575 2336 1579 2340
rect 1815 2336 1819 2340
rect 1935 2335 1939 2339
rect 1975 2321 1979 2325
rect 2223 2320 2227 2324
rect 2503 2320 2507 2324
rect 2767 2320 2771 2324
rect 3007 2320 3011 2324
rect 3239 2320 3243 2324
rect 3471 2320 3475 2324
rect 3679 2320 3683 2324
rect 3799 2321 3803 2325
rect 1975 2304 1979 2308
rect 2195 2305 2199 2309
rect 2475 2305 2479 2309
rect 2739 2305 2743 2309
rect 2979 2305 2983 2309
rect 3211 2305 3215 2309
rect 3443 2305 3447 2309
rect 3651 2305 3655 2309
rect 3799 2304 3803 2308
rect 3839 2281 3843 2285
rect 3887 2280 3891 2284
rect 4183 2280 4187 2284
rect 4495 2280 4499 2284
rect 4791 2280 4795 2284
rect 5087 2280 5091 2284
rect 5383 2280 5387 2284
rect 5663 2281 5667 2285
rect 111 2273 115 2277
rect 159 2272 163 2276
rect 319 2272 323 2276
rect 551 2272 555 2276
rect 831 2272 835 2276
rect 1151 2272 1155 2276
rect 1495 2272 1499 2276
rect 1815 2272 1819 2276
rect 1935 2273 1939 2277
rect 3839 2264 3843 2268
rect 3859 2265 3863 2269
rect 4155 2265 4159 2269
rect 4467 2265 4471 2269
rect 4763 2265 4767 2269
rect 5059 2265 5063 2269
rect 5355 2265 5359 2269
rect 5663 2264 5667 2268
rect 111 2256 115 2260
rect 131 2257 135 2261
rect 291 2257 295 2261
rect 523 2257 527 2261
rect 803 2257 807 2261
rect 1123 2257 1127 2261
rect 1467 2257 1471 2261
rect 1787 2257 1791 2261
rect 1935 2256 1939 2260
rect 1975 2172 1979 2176
rect 1995 2171 1999 2175
rect 2155 2171 2159 2175
rect 2387 2171 2391 2175
rect 2667 2171 2671 2175
rect 2987 2171 2991 2175
rect 3331 2171 3335 2175
rect 3651 2171 3655 2175
rect 3799 2172 3803 2176
rect 1975 2155 1979 2159
rect 2023 2156 2027 2160
rect 2183 2156 2187 2160
rect 2415 2156 2419 2160
rect 2695 2156 2699 2160
rect 3015 2156 3019 2160
rect 3359 2156 3363 2160
rect 3679 2156 3683 2160
rect 3799 2155 3803 2159
rect 3839 2128 3843 2132
rect 3859 2127 3863 2131
rect 3995 2127 3999 2131
rect 4131 2127 4135 2131
rect 4267 2127 4271 2131
rect 4403 2127 4407 2131
rect 4539 2127 4543 2131
rect 4699 2127 4703 2131
rect 4891 2127 4895 2131
rect 5099 2127 5103 2131
rect 5315 2127 5319 2131
rect 5515 2127 5519 2131
rect 5663 2128 5667 2132
rect 3839 2111 3843 2115
rect 3887 2112 3891 2116
rect 4023 2112 4027 2116
rect 4159 2112 4163 2116
rect 4295 2112 4299 2116
rect 4431 2112 4435 2116
rect 4567 2112 4571 2116
rect 4727 2112 4731 2116
rect 4919 2112 4923 2116
rect 5127 2112 5131 2116
rect 5343 2112 5347 2116
rect 5543 2112 5547 2116
rect 5663 2111 5667 2115
rect 111 2100 115 2104
rect 291 2099 295 2103
rect 483 2099 487 2103
rect 691 2099 695 2103
rect 915 2099 919 2103
rect 1147 2099 1151 2103
rect 1387 2099 1391 2103
rect 1635 2099 1639 2103
rect 1935 2100 1939 2104
rect 111 2083 115 2087
rect 319 2084 323 2088
rect 511 2084 515 2088
rect 719 2084 723 2088
rect 943 2084 947 2088
rect 1175 2084 1179 2088
rect 1415 2084 1419 2088
rect 1663 2084 1667 2088
rect 1935 2083 1939 2087
rect 3839 2033 3843 2037
rect 3887 2032 3891 2036
rect 4023 2032 4027 2036
rect 4159 2032 4163 2036
rect 4295 2032 4299 2036
rect 4431 2032 4435 2036
rect 4567 2032 4571 2036
rect 4719 2032 4723 2036
rect 4895 2032 4899 2036
rect 5087 2032 5091 2036
rect 5279 2032 5283 2036
rect 5479 2032 5483 2036
rect 5663 2033 5667 2037
rect 111 2021 115 2025
rect 263 2020 267 2024
rect 399 2020 403 2024
rect 535 2020 539 2024
rect 679 2020 683 2024
rect 823 2020 827 2024
rect 967 2020 971 2024
rect 1111 2020 1115 2024
rect 1255 2020 1259 2024
rect 1399 2020 1403 2024
rect 1543 2020 1547 2024
rect 1679 2020 1683 2024
rect 1815 2020 1819 2024
rect 1935 2021 1939 2025
rect 3839 2016 3843 2020
rect 3859 2017 3863 2021
rect 3995 2017 3999 2021
rect 4131 2017 4135 2021
rect 4267 2017 4271 2021
rect 4403 2017 4407 2021
rect 4539 2017 4543 2021
rect 4691 2017 4695 2021
rect 4867 2017 4871 2021
rect 5059 2017 5063 2021
rect 5251 2017 5255 2021
rect 5451 2017 5455 2021
rect 5663 2016 5667 2020
rect 111 2004 115 2008
rect 235 2005 239 2009
rect 371 2005 375 2009
rect 507 2005 511 2009
rect 651 2005 655 2009
rect 795 2005 799 2009
rect 939 2005 943 2009
rect 1083 2005 1087 2009
rect 1227 2005 1231 2009
rect 1371 2005 1375 2009
rect 1515 2005 1519 2009
rect 1651 2005 1655 2009
rect 1787 2005 1791 2009
rect 1935 2004 1939 2008
rect 1975 1897 1979 1901
rect 3135 1896 3139 1900
rect 3271 1896 3275 1900
rect 3407 1896 3411 1900
rect 3543 1896 3547 1900
rect 3679 1896 3683 1900
rect 3799 1897 3803 1901
rect 1975 1880 1979 1884
rect 3107 1881 3111 1885
rect 3243 1881 3247 1885
rect 3379 1881 3383 1885
rect 3515 1881 3519 1885
rect 3651 1881 3655 1885
rect 3799 1880 3803 1884
rect 3839 1884 3843 1888
rect 3859 1883 3863 1887
rect 4043 1883 4047 1887
rect 4283 1883 4287 1887
rect 4563 1883 4567 1887
rect 4875 1883 4879 1887
rect 5203 1883 5207 1887
rect 5515 1883 5519 1887
rect 5663 1884 5667 1888
rect 3839 1867 3843 1871
rect 3887 1868 3891 1872
rect 4071 1868 4075 1872
rect 4311 1868 4315 1872
rect 4591 1868 4595 1872
rect 4903 1868 4907 1872
rect 5231 1868 5235 1872
rect 5543 1868 5547 1872
rect 5663 1867 5667 1871
rect 111 1860 115 1864
rect 235 1859 239 1863
rect 435 1859 439 1863
rect 627 1859 631 1863
rect 811 1859 815 1863
rect 987 1859 991 1863
rect 1155 1859 1159 1863
rect 1323 1859 1327 1863
rect 1483 1859 1487 1863
rect 1643 1859 1647 1863
rect 1787 1859 1791 1863
rect 1935 1860 1939 1864
rect 111 1843 115 1847
rect 263 1844 267 1848
rect 463 1844 467 1848
rect 655 1844 659 1848
rect 839 1844 843 1848
rect 1015 1844 1019 1848
rect 1183 1844 1187 1848
rect 1351 1844 1355 1848
rect 1511 1844 1515 1848
rect 1671 1844 1675 1848
rect 1815 1844 1819 1848
rect 1935 1843 1939 1847
rect 3839 1809 3843 1813
rect 4407 1808 4411 1812
rect 4543 1808 4547 1812
rect 4679 1808 4683 1812
rect 4815 1808 4819 1812
rect 4951 1808 4955 1812
rect 5663 1809 5667 1813
rect 3839 1792 3843 1796
rect 4379 1793 4383 1797
rect 4515 1793 4519 1797
rect 4651 1793 4655 1797
rect 4787 1793 4791 1797
rect 4923 1793 4927 1797
rect 5663 1792 5667 1796
rect 111 1773 115 1777
rect 223 1772 227 1776
rect 463 1772 467 1776
rect 695 1772 699 1776
rect 927 1772 931 1776
rect 1159 1772 1163 1776
rect 1391 1772 1395 1776
rect 1935 1773 1939 1777
rect 111 1756 115 1760
rect 195 1757 199 1761
rect 435 1757 439 1761
rect 667 1757 671 1761
rect 899 1757 903 1761
rect 1131 1757 1135 1761
rect 1363 1757 1367 1761
rect 1935 1756 1939 1760
rect 1975 1736 1979 1740
rect 1995 1735 1999 1739
rect 2131 1735 2135 1739
rect 2267 1735 2271 1739
rect 2419 1735 2423 1739
rect 2579 1735 2583 1739
rect 2739 1735 2743 1739
rect 2899 1735 2903 1739
rect 3051 1735 3055 1739
rect 3203 1735 3207 1739
rect 3355 1735 3359 1739
rect 3515 1735 3519 1739
rect 3651 1735 3655 1739
rect 3799 1736 3803 1740
rect 1975 1719 1979 1723
rect 2023 1720 2027 1724
rect 2159 1720 2163 1724
rect 2295 1720 2299 1724
rect 2447 1720 2451 1724
rect 2607 1720 2611 1724
rect 2767 1720 2771 1724
rect 2927 1720 2931 1724
rect 3079 1720 3083 1724
rect 3231 1720 3235 1724
rect 3383 1720 3387 1724
rect 3543 1720 3547 1724
rect 3679 1720 3683 1724
rect 3799 1719 3803 1723
rect 1975 1649 1979 1653
rect 2023 1648 2027 1652
rect 2167 1648 2171 1652
rect 2319 1648 2323 1652
rect 2479 1648 2483 1652
rect 2639 1648 2643 1652
rect 2791 1648 2795 1652
rect 2943 1648 2947 1652
rect 3103 1648 3107 1652
rect 3263 1648 3267 1652
rect 3423 1648 3427 1652
rect 3799 1649 3803 1653
rect 3839 1644 3843 1648
rect 4563 1643 4567 1647
rect 4699 1643 4703 1647
rect 4835 1643 4839 1647
rect 4971 1643 4975 1647
rect 5107 1643 5111 1647
rect 5243 1643 5247 1647
rect 5379 1643 5383 1647
rect 5515 1643 5519 1647
rect 5663 1644 5667 1648
rect 1975 1632 1979 1636
rect 1995 1633 1999 1637
rect 2139 1633 2143 1637
rect 2291 1633 2295 1637
rect 2451 1633 2455 1637
rect 2611 1633 2615 1637
rect 2763 1633 2767 1637
rect 2915 1633 2919 1637
rect 3075 1633 3079 1637
rect 3235 1633 3239 1637
rect 3395 1633 3399 1637
rect 3799 1632 3803 1636
rect 3839 1627 3843 1631
rect 4591 1628 4595 1632
rect 4727 1628 4731 1632
rect 4863 1628 4867 1632
rect 4999 1628 5003 1632
rect 5135 1628 5139 1632
rect 5271 1628 5275 1632
rect 5407 1628 5411 1632
rect 5543 1628 5547 1632
rect 5663 1627 5667 1631
rect 111 1612 115 1616
rect 131 1611 135 1615
rect 363 1611 367 1615
rect 619 1611 623 1615
rect 875 1611 879 1615
rect 1139 1611 1143 1615
rect 1935 1612 1939 1616
rect 111 1595 115 1599
rect 159 1596 163 1600
rect 391 1596 395 1600
rect 647 1596 651 1600
rect 903 1596 907 1600
rect 1167 1596 1171 1600
rect 1935 1595 1939 1599
rect 3839 1553 3843 1557
rect 4591 1552 4595 1556
rect 4727 1552 4731 1556
rect 4863 1552 4867 1556
rect 4999 1552 5003 1556
rect 5135 1552 5139 1556
rect 5271 1552 5275 1556
rect 5407 1552 5411 1556
rect 5543 1552 5547 1556
rect 5663 1553 5667 1557
rect 3839 1536 3843 1540
rect 4563 1537 4567 1541
rect 4699 1537 4703 1541
rect 4835 1537 4839 1541
rect 4971 1537 4975 1541
rect 5107 1537 5111 1541
rect 5243 1537 5247 1541
rect 5379 1537 5383 1541
rect 5515 1537 5519 1541
rect 5663 1536 5667 1540
rect 111 1525 115 1529
rect 159 1524 163 1528
rect 327 1524 331 1528
rect 511 1524 515 1528
rect 695 1524 699 1528
rect 887 1524 891 1528
rect 1079 1524 1083 1528
rect 1935 1525 1939 1529
rect 111 1508 115 1512
rect 131 1509 135 1513
rect 299 1509 303 1513
rect 483 1509 487 1513
rect 667 1509 671 1513
rect 859 1509 863 1513
rect 1051 1509 1055 1513
rect 1935 1508 1939 1512
rect 1975 1488 1979 1492
rect 1995 1487 1999 1491
rect 2131 1487 2135 1491
rect 2267 1487 2271 1491
rect 2403 1487 2407 1491
rect 2539 1487 2543 1491
rect 2675 1487 2679 1491
rect 2811 1487 2815 1491
rect 2947 1487 2951 1491
rect 3083 1487 3087 1491
rect 3219 1487 3223 1491
rect 3355 1487 3359 1491
rect 3491 1487 3495 1491
rect 3799 1488 3803 1492
rect 1975 1471 1979 1475
rect 2023 1472 2027 1476
rect 2159 1472 2163 1476
rect 2295 1472 2299 1476
rect 2431 1472 2435 1476
rect 2567 1472 2571 1476
rect 2703 1472 2707 1476
rect 2839 1472 2843 1476
rect 2975 1472 2979 1476
rect 3111 1472 3115 1476
rect 3247 1472 3251 1476
rect 3383 1472 3387 1476
rect 3519 1472 3523 1476
rect 3799 1471 3803 1475
rect 1975 1401 1979 1405
rect 2167 1400 2171 1404
rect 2303 1400 2307 1404
rect 2439 1400 2443 1404
rect 2575 1400 2579 1404
rect 2711 1400 2715 1404
rect 2847 1400 2851 1404
rect 2983 1400 2987 1404
rect 3119 1400 3123 1404
rect 3255 1400 3259 1404
rect 3799 1401 3803 1405
rect 1975 1384 1979 1388
rect 2139 1385 2143 1389
rect 2275 1385 2279 1389
rect 2411 1385 2415 1389
rect 2547 1385 2551 1389
rect 2683 1385 2687 1389
rect 2819 1385 2823 1389
rect 2955 1385 2959 1389
rect 3091 1385 3095 1389
rect 3227 1385 3231 1389
rect 3799 1384 3803 1388
rect 111 1364 115 1368
rect 131 1363 135 1367
rect 395 1363 399 1367
rect 683 1363 687 1367
rect 971 1363 975 1367
rect 1259 1363 1263 1367
rect 1935 1364 1939 1368
rect 111 1347 115 1351
rect 159 1348 163 1352
rect 423 1348 427 1352
rect 711 1348 715 1352
rect 999 1348 1003 1352
rect 1287 1348 1291 1352
rect 1935 1347 1939 1351
rect 3839 1332 3843 1336
rect 4811 1331 4815 1335
rect 4947 1331 4951 1335
rect 5083 1331 5087 1335
rect 5219 1331 5223 1335
rect 5355 1331 5359 1335
rect 5491 1331 5495 1335
rect 5663 1332 5667 1336
rect 3839 1315 3843 1319
rect 4839 1316 4843 1320
rect 4975 1316 4979 1320
rect 5111 1316 5115 1320
rect 5247 1316 5251 1320
rect 5383 1316 5387 1320
rect 5519 1316 5523 1320
rect 5663 1315 5667 1319
rect 111 1289 115 1293
rect 159 1288 163 1292
rect 455 1288 459 1292
rect 775 1288 779 1292
rect 1095 1288 1099 1292
rect 1423 1288 1427 1292
rect 1935 1289 1939 1293
rect 111 1272 115 1276
rect 131 1273 135 1277
rect 427 1273 431 1277
rect 747 1273 751 1277
rect 1067 1273 1071 1277
rect 1395 1273 1399 1277
rect 1935 1272 1939 1276
rect 1975 1252 1979 1256
rect 2131 1251 2135 1255
rect 2267 1251 2271 1255
rect 2403 1251 2407 1255
rect 2555 1251 2559 1255
rect 2715 1251 2719 1255
rect 2891 1251 2895 1255
rect 3075 1251 3079 1255
rect 3267 1251 3271 1255
rect 3467 1251 3471 1255
rect 3651 1251 3655 1255
rect 3799 1252 3803 1256
rect 3839 1253 3843 1257
rect 4735 1252 4739 1256
rect 4879 1252 4883 1256
rect 5031 1252 5035 1256
rect 5191 1252 5195 1256
rect 5359 1252 5363 1256
rect 5527 1252 5531 1256
rect 5663 1253 5667 1257
rect 1975 1235 1979 1239
rect 2159 1236 2163 1240
rect 2295 1236 2299 1240
rect 2431 1236 2435 1240
rect 2583 1236 2587 1240
rect 2743 1236 2747 1240
rect 2919 1236 2923 1240
rect 3103 1236 3107 1240
rect 3295 1236 3299 1240
rect 3495 1236 3499 1240
rect 3679 1236 3683 1240
rect 3799 1235 3803 1239
rect 3839 1236 3843 1240
rect 4707 1237 4711 1241
rect 4851 1237 4855 1241
rect 5003 1237 5007 1241
rect 5163 1237 5167 1241
rect 5331 1237 5335 1241
rect 5499 1237 5503 1241
rect 5663 1236 5667 1240
rect 1975 1177 1979 1181
rect 2023 1176 2027 1180
rect 2239 1176 2243 1180
rect 2479 1176 2483 1180
rect 2719 1176 2723 1180
rect 2959 1176 2963 1180
rect 3207 1176 3211 1180
rect 3455 1176 3459 1180
rect 3679 1176 3683 1180
rect 3799 1177 3803 1181
rect 1975 1160 1979 1164
rect 1995 1161 1999 1165
rect 2211 1161 2215 1165
rect 2451 1161 2455 1165
rect 2691 1161 2695 1165
rect 2931 1161 2935 1165
rect 3179 1161 3183 1165
rect 3427 1161 3431 1165
rect 3651 1161 3655 1165
rect 3799 1160 3803 1164
rect 111 1116 115 1120
rect 131 1115 135 1119
rect 331 1115 335 1119
rect 563 1115 567 1119
rect 803 1115 807 1119
rect 1043 1115 1047 1119
rect 1283 1115 1287 1119
rect 1523 1115 1527 1119
rect 1771 1115 1775 1119
rect 1935 1116 1939 1120
rect 111 1099 115 1103
rect 159 1100 163 1104
rect 359 1100 363 1104
rect 591 1100 595 1104
rect 831 1100 835 1104
rect 1071 1100 1075 1104
rect 1311 1100 1315 1104
rect 1551 1100 1555 1104
rect 1799 1100 1803 1104
rect 1935 1099 1939 1103
rect 3839 1096 3843 1100
rect 3859 1095 3863 1099
rect 4067 1095 4071 1099
rect 4299 1095 4303 1099
rect 4539 1095 4543 1099
rect 4779 1095 4783 1099
rect 5027 1095 5031 1099
rect 5283 1095 5287 1099
rect 5515 1095 5519 1099
rect 5663 1096 5667 1100
rect 3839 1079 3843 1083
rect 3887 1080 3891 1084
rect 4095 1080 4099 1084
rect 4327 1080 4331 1084
rect 4567 1080 4571 1084
rect 4807 1080 4811 1084
rect 5055 1080 5059 1084
rect 5311 1080 5315 1084
rect 5543 1080 5547 1084
rect 5663 1079 5667 1083
rect 111 1041 115 1045
rect 263 1040 267 1044
rect 439 1040 443 1044
rect 615 1040 619 1044
rect 783 1040 787 1044
rect 951 1040 955 1044
rect 1111 1040 1115 1044
rect 1271 1040 1275 1044
rect 1431 1040 1435 1044
rect 1591 1040 1595 1044
rect 1751 1040 1755 1044
rect 1935 1041 1939 1045
rect 111 1024 115 1028
rect 235 1025 239 1029
rect 411 1025 415 1029
rect 587 1025 591 1029
rect 755 1025 759 1029
rect 923 1025 927 1029
rect 1083 1025 1087 1029
rect 1243 1025 1247 1029
rect 1403 1025 1407 1029
rect 1563 1025 1567 1029
rect 1723 1025 1727 1029
rect 1935 1024 1939 1028
rect 3839 1021 3843 1025
rect 3887 1020 3891 1024
rect 4071 1020 4075 1024
rect 4279 1020 4283 1024
rect 4511 1020 4515 1024
rect 4759 1020 4763 1024
rect 5023 1020 5027 1024
rect 5295 1020 5299 1024
rect 5543 1020 5547 1024
rect 5663 1021 5667 1025
rect 1975 1004 1979 1008
rect 3091 1003 3095 1007
rect 3243 1003 3247 1007
rect 3395 1003 3399 1007
rect 3799 1004 3803 1008
rect 3839 1004 3843 1008
rect 3859 1005 3863 1009
rect 4043 1005 4047 1009
rect 4251 1005 4255 1009
rect 4483 1005 4487 1009
rect 4731 1005 4735 1009
rect 4995 1005 4999 1009
rect 5267 1005 5271 1009
rect 5515 1005 5519 1009
rect 5663 1004 5667 1008
rect 1975 987 1979 991
rect 3119 988 3123 992
rect 3271 988 3275 992
rect 3423 988 3427 992
rect 3799 987 3803 991
rect 1975 901 1979 905
rect 2047 900 2051 904
rect 2351 900 2355 904
rect 2647 900 2651 904
rect 2927 900 2931 904
rect 3207 900 3211 904
rect 3495 900 3499 904
rect 3799 901 3803 905
rect 111 888 115 892
rect 227 887 231 891
rect 379 887 383 891
rect 539 887 543 891
rect 715 887 719 891
rect 891 887 895 891
rect 1075 887 1079 891
rect 1259 887 1263 891
rect 1443 887 1447 891
rect 1627 887 1631 891
rect 1787 887 1791 891
rect 1935 888 1939 892
rect 1975 884 1979 888
rect 2019 885 2023 889
rect 2323 885 2327 889
rect 2619 885 2623 889
rect 2899 885 2903 889
rect 3179 885 3183 889
rect 3467 885 3471 889
rect 3799 884 3803 888
rect 111 871 115 875
rect 255 872 259 876
rect 407 872 411 876
rect 567 872 571 876
rect 743 872 747 876
rect 919 872 923 876
rect 1103 872 1107 876
rect 1287 872 1291 876
rect 1471 872 1475 876
rect 1655 872 1659 876
rect 1815 872 1819 876
rect 1935 871 1939 875
rect 3839 872 3843 876
rect 3971 871 3975 875
rect 4179 871 4183 875
rect 4403 871 4407 875
rect 4643 871 4647 875
rect 4899 871 4903 875
rect 5171 871 5175 875
rect 5443 871 5447 875
rect 5663 872 5667 876
rect 3839 855 3843 859
rect 3999 856 4003 860
rect 4207 856 4211 860
rect 4431 856 4435 860
rect 4671 856 4675 860
rect 4927 856 4931 860
rect 5199 856 5203 860
rect 5471 856 5475 860
rect 5663 855 5667 859
rect 111 797 115 801
rect 375 796 379 800
rect 655 796 659 800
rect 943 796 947 800
rect 1239 796 1243 800
rect 1535 796 1539 800
rect 1815 796 1819 800
rect 1935 797 1939 801
rect 3839 797 3843 801
rect 3887 796 3891 800
rect 4047 796 4051 800
rect 4279 796 4283 800
rect 4559 796 4563 800
rect 4879 796 4883 800
rect 5223 796 5227 800
rect 5543 796 5547 800
rect 5663 797 5667 801
rect 111 780 115 784
rect 347 781 351 785
rect 627 781 631 785
rect 915 781 919 785
rect 1211 781 1215 785
rect 1507 781 1511 785
rect 1787 781 1791 785
rect 1935 780 1939 784
rect 3839 780 3843 784
rect 3859 781 3863 785
rect 4019 781 4023 785
rect 4251 781 4255 785
rect 4531 781 4535 785
rect 4851 781 4855 785
rect 5195 781 5199 785
rect 5515 781 5519 785
rect 5663 780 5667 784
rect 1975 752 1979 756
rect 1995 751 1999 755
rect 2251 751 2255 755
rect 2523 751 2527 755
rect 2771 751 2775 755
rect 3003 751 3007 755
rect 3227 751 3231 755
rect 3451 751 3455 755
rect 3651 751 3655 755
rect 3799 752 3803 756
rect 1975 735 1979 739
rect 2023 736 2027 740
rect 2279 736 2283 740
rect 2551 736 2555 740
rect 2799 736 2803 740
rect 3031 736 3035 740
rect 3255 736 3259 740
rect 3479 736 3483 740
rect 3679 736 3683 740
rect 3799 735 3803 739
rect 111 648 115 652
rect 131 647 135 651
rect 307 647 311 651
rect 499 647 503 651
rect 683 647 687 651
rect 859 647 863 651
rect 1027 647 1031 651
rect 1187 647 1191 651
rect 1339 647 1343 651
rect 1491 647 1495 651
rect 1651 647 1655 651
rect 1787 647 1791 651
rect 1935 648 1939 652
rect 3839 640 3843 644
rect 3859 639 3863 643
rect 3995 639 3999 643
rect 4131 639 4135 643
rect 4267 639 4271 643
rect 4403 639 4407 643
rect 4571 639 4575 643
rect 4771 639 4775 643
rect 4995 639 4999 643
rect 5227 639 5231 643
rect 5459 639 5463 643
rect 5663 640 5667 644
rect 111 631 115 635
rect 159 632 163 636
rect 335 632 339 636
rect 527 632 531 636
rect 711 632 715 636
rect 887 632 891 636
rect 1055 632 1059 636
rect 1215 632 1219 636
rect 1367 632 1371 636
rect 1519 632 1523 636
rect 1679 632 1683 636
rect 1815 632 1819 636
rect 1935 631 1939 635
rect 3839 623 3843 627
rect 3887 624 3891 628
rect 4023 624 4027 628
rect 4159 624 4163 628
rect 4295 624 4299 628
rect 4431 624 4435 628
rect 4599 624 4603 628
rect 4799 624 4803 628
rect 5023 624 5027 628
rect 5255 624 5259 628
rect 5487 624 5491 628
rect 5663 623 5667 627
rect 111 573 115 577
rect 159 572 163 576
rect 375 572 379 576
rect 599 572 603 576
rect 807 572 811 576
rect 999 572 1003 576
rect 1175 572 1179 576
rect 1343 572 1347 576
rect 1511 572 1515 576
rect 1671 572 1675 576
rect 1815 572 1819 576
rect 1935 573 1939 577
rect 3839 565 3843 569
rect 3887 564 3891 568
rect 4023 564 4027 568
rect 4159 564 4163 568
rect 4295 564 4299 568
rect 4479 564 4483 568
rect 4695 564 4699 568
rect 4935 564 4939 568
rect 5191 564 5195 568
rect 5447 564 5451 568
rect 5663 565 5667 569
rect 111 556 115 560
rect 131 557 135 561
rect 347 557 351 561
rect 571 557 575 561
rect 779 557 783 561
rect 971 557 975 561
rect 1147 557 1151 561
rect 1315 557 1319 561
rect 1483 557 1487 561
rect 1643 557 1647 561
rect 1787 557 1791 561
rect 1935 556 1939 560
rect 1975 545 1979 549
rect 3311 544 3315 548
rect 3447 544 3451 548
rect 3583 544 3587 548
rect 3799 545 3803 549
rect 3839 548 3843 552
rect 3859 549 3863 553
rect 3995 549 3999 553
rect 4131 549 4135 553
rect 4267 549 4271 553
rect 4451 549 4455 553
rect 4667 549 4671 553
rect 4907 549 4911 553
rect 5163 549 5167 553
rect 5419 549 5423 553
rect 5663 548 5667 552
rect 1975 528 1979 532
rect 3283 529 3287 533
rect 3419 529 3423 533
rect 3555 529 3559 533
rect 3799 528 3803 532
rect 111 424 115 428
rect 131 423 135 427
rect 427 423 431 427
rect 763 423 767 427
rect 1107 423 1111 427
rect 1459 423 1463 427
rect 1787 423 1791 427
rect 1935 424 1939 428
rect 111 407 115 411
rect 159 408 163 412
rect 455 408 459 412
rect 791 408 795 412
rect 1135 408 1139 412
rect 1487 408 1491 412
rect 1815 408 1819 412
rect 1935 407 1939 411
rect 3839 404 3843 408
rect 4451 403 4455 407
rect 4651 403 4655 407
rect 4859 403 4863 407
rect 5067 403 5071 407
rect 5283 403 5287 407
rect 5507 403 5511 407
rect 5663 404 5667 408
rect 1975 396 1979 400
rect 1995 395 1999 399
rect 2155 395 2159 399
rect 2347 395 2351 399
rect 2539 395 2543 399
rect 2731 395 2735 399
rect 2923 395 2927 399
rect 3115 395 3119 399
rect 3299 395 3303 399
rect 3483 395 3487 399
rect 3651 395 3655 399
rect 3799 396 3803 400
rect 3839 387 3843 391
rect 4479 388 4483 392
rect 4679 388 4683 392
rect 4887 388 4891 392
rect 5095 388 5099 392
rect 5311 388 5315 392
rect 5535 388 5539 392
rect 5663 387 5667 391
rect 1975 379 1979 383
rect 2023 380 2027 384
rect 2183 380 2187 384
rect 2375 380 2379 384
rect 2567 380 2571 384
rect 2759 380 2763 384
rect 2951 380 2955 384
rect 3143 380 3147 384
rect 3327 380 3331 384
rect 3511 380 3515 384
rect 3679 380 3683 384
rect 3799 379 3803 383
rect 111 333 115 337
rect 239 332 243 336
rect 391 332 395 336
rect 551 332 555 336
rect 711 332 715 336
rect 871 332 875 336
rect 1031 332 1035 336
rect 1935 333 1939 337
rect 3839 325 3843 329
rect 4751 324 4755 328
rect 4911 324 4915 328
rect 5071 324 5075 328
rect 5231 324 5235 328
rect 5399 324 5403 328
rect 5543 324 5547 328
rect 5663 325 5667 329
rect 111 316 115 320
rect 211 317 215 321
rect 363 317 367 321
rect 523 317 527 321
rect 683 317 687 321
rect 843 317 847 321
rect 1003 317 1007 321
rect 1935 316 1939 320
rect 3839 308 3843 312
rect 4723 309 4727 313
rect 4883 309 4887 313
rect 5043 309 5047 313
rect 5203 309 5207 313
rect 5371 309 5375 313
rect 5515 309 5519 313
rect 5663 308 5667 312
rect 1975 297 1979 301
rect 2047 296 2051 300
rect 2183 296 2187 300
rect 2319 296 2323 300
rect 2455 296 2459 300
rect 2591 296 2595 300
rect 2727 296 2731 300
rect 2863 296 2867 300
rect 2999 296 3003 300
rect 3135 296 3139 300
rect 3271 296 3275 300
rect 3407 296 3411 300
rect 3543 296 3547 300
rect 3679 296 3683 300
rect 3799 297 3803 301
rect 1975 280 1979 284
rect 2019 281 2023 285
rect 2155 281 2159 285
rect 2291 281 2295 285
rect 2427 281 2431 285
rect 2563 281 2567 285
rect 2699 281 2703 285
rect 2835 281 2839 285
rect 2971 281 2975 285
rect 3107 281 3111 285
rect 3243 281 3247 285
rect 3379 281 3383 285
rect 3515 281 3519 285
rect 3651 281 3655 285
rect 3799 280 3803 284
rect 111 152 115 156
rect 147 151 151 155
rect 283 151 287 155
rect 419 151 423 155
rect 555 151 559 155
rect 691 151 695 155
rect 827 151 831 155
rect 963 151 967 155
rect 1099 151 1103 155
rect 1935 152 1939 156
rect 111 135 115 139
rect 175 136 179 140
rect 311 136 315 140
rect 447 136 451 140
rect 583 136 587 140
rect 719 136 723 140
rect 855 136 859 140
rect 991 136 995 140
rect 1127 136 1131 140
rect 1935 135 1939 139
rect 1975 132 1979 136
rect 1995 131 1999 135
rect 2131 131 2135 135
rect 2267 131 2271 135
rect 2403 131 2407 135
rect 2539 131 2543 135
rect 2675 131 2679 135
rect 2811 131 2815 135
rect 2947 131 2951 135
rect 3083 131 3087 135
rect 3219 131 3223 135
rect 3355 131 3359 135
rect 3491 131 3495 135
rect 3627 131 3631 135
rect 3799 132 3803 136
rect 3839 136 3843 140
rect 4291 135 4295 139
rect 4427 135 4431 139
rect 4563 135 4567 139
rect 4699 135 4703 139
rect 4835 135 4839 139
rect 4971 135 4975 139
rect 5107 135 5111 139
rect 5243 135 5247 139
rect 5379 135 5383 139
rect 5515 135 5519 139
rect 5663 136 5667 140
rect 1975 115 1979 119
rect 2023 116 2027 120
rect 2159 116 2163 120
rect 2295 116 2299 120
rect 2431 116 2435 120
rect 2567 116 2571 120
rect 2703 116 2707 120
rect 2839 116 2843 120
rect 2975 116 2979 120
rect 3111 116 3115 120
rect 3247 116 3251 120
rect 3383 116 3387 120
rect 3519 116 3523 120
rect 3655 116 3659 120
rect 3799 115 3803 119
rect 3839 119 3843 123
rect 4319 120 4323 124
rect 4455 120 4459 124
rect 4591 120 4595 124
rect 4727 120 4731 124
rect 4863 120 4867 124
rect 4999 120 5003 124
rect 5135 120 5139 124
rect 5271 120 5275 124
rect 5407 120 5411 124
rect 5543 120 5547 124
rect 5663 119 5667 123
<< m3 >>
rect 111 5758 115 5759
rect 111 5753 115 5754
rect 131 5758 135 5759
rect 131 5753 135 5754
rect 267 5758 271 5759
rect 267 5753 271 5754
rect 403 5758 407 5759
rect 403 5753 407 5754
rect 1935 5758 1939 5759
rect 1935 5753 1939 5754
rect 112 5693 114 5753
rect 110 5692 116 5693
rect 132 5692 134 5753
rect 268 5692 270 5753
rect 404 5692 406 5753
rect 1936 5693 1938 5753
rect 3839 5694 3843 5695
rect 1934 5692 1940 5693
rect 110 5688 111 5692
rect 115 5688 116 5692
rect 110 5687 116 5688
rect 130 5691 136 5692
rect 130 5687 131 5691
rect 135 5687 136 5691
rect 130 5686 136 5687
rect 266 5691 272 5692
rect 266 5687 267 5691
rect 271 5687 272 5691
rect 266 5686 272 5687
rect 402 5691 408 5692
rect 402 5687 403 5691
rect 407 5687 408 5691
rect 1934 5688 1935 5692
rect 1939 5688 1940 5692
rect 1934 5687 1940 5688
rect 1975 5690 1979 5691
rect 402 5686 408 5687
rect 1975 5685 1979 5686
rect 1995 5690 1999 5691
rect 1995 5685 1999 5686
rect 2171 5690 2175 5691
rect 2171 5685 2175 5686
rect 2371 5690 2375 5691
rect 2371 5685 2375 5686
rect 2563 5690 2567 5691
rect 2563 5685 2567 5686
rect 2747 5690 2751 5691
rect 2747 5685 2751 5686
rect 2931 5690 2935 5691
rect 2931 5685 2935 5686
rect 3107 5690 3111 5691
rect 3107 5685 3111 5686
rect 3275 5690 3279 5691
rect 3275 5685 3279 5686
rect 3443 5690 3447 5691
rect 3443 5685 3447 5686
rect 3619 5690 3623 5691
rect 3619 5685 3623 5686
rect 3799 5690 3803 5691
rect 3839 5689 3843 5690
rect 4467 5694 4471 5695
rect 4467 5689 4471 5690
rect 4603 5694 4607 5695
rect 4603 5689 4607 5690
rect 4739 5694 4743 5695
rect 4739 5689 4743 5690
rect 4875 5694 4879 5695
rect 4875 5689 4879 5690
rect 5663 5694 5667 5695
rect 5663 5689 5667 5690
rect 3799 5685 3803 5686
rect 158 5676 164 5677
rect 110 5675 116 5676
rect 110 5671 111 5675
rect 115 5671 116 5675
rect 158 5672 159 5676
rect 163 5672 164 5676
rect 158 5671 164 5672
rect 294 5676 300 5677
rect 294 5672 295 5676
rect 299 5672 300 5676
rect 294 5671 300 5672
rect 430 5676 436 5677
rect 430 5672 431 5676
rect 435 5672 436 5676
rect 430 5671 436 5672
rect 1934 5675 1940 5676
rect 1934 5671 1935 5675
rect 1939 5671 1940 5675
rect 110 5670 116 5671
rect 112 5647 114 5670
rect 160 5647 162 5671
rect 296 5647 298 5671
rect 432 5647 434 5671
rect 1934 5670 1940 5671
rect 1936 5647 1938 5670
rect 111 5646 115 5647
rect 111 5641 115 5642
rect 159 5646 163 5647
rect 159 5641 163 5642
rect 295 5646 299 5647
rect 295 5641 299 5642
rect 343 5646 347 5647
rect 343 5641 347 5642
rect 431 5646 435 5647
rect 431 5641 435 5642
rect 535 5646 539 5647
rect 535 5641 539 5642
rect 735 5646 739 5647
rect 735 5641 739 5642
rect 943 5646 947 5647
rect 943 5641 947 5642
rect 1159 5646 1163 5647
rect 1159 5641 1163 5642
rect 1383 5646 1387 5647
rect 1383 5641 1387 5642
rect 1607 5646 1611 5647
rect 1607 5641 1611 5642
rect 1815 5646 1819 5647
rect 1815 5641 1819 5642
rect 1935 5646 1939 5647
rect 1935 5641 1939 5642
rect 112 5618 114 5641
rect 110 5617 116 5618
rect 344 5617 346 5641
rect 536 5617 538 5641
rect 736 5617 738 5641
rect 944 5617 946 5641
rect 1160 5617 1162 5641
rect 1384 5617 1386 5641
rect 1608 5617 1610 5641
rect 1816 5617 1818 5641
rect 1936 5618 1938 5641
rect 1976 5625 1978 5685
rect 1974 5624 1980 5625
rect 1996 5624 1998 5685
rect 2172 5624 2174 5685
rect 2372 5624 2374 5685
rect 2564 5624 2566 5685
rect 2748 5624 2750 5685
rect 2932 5624 2934 5685
rect 3108 5624 3110 5685
rect 3276 5624 3278 5685
rect 3444 5624 3446 5685
rect 3620 5624 3622 5685
rect 3800 5625 3802 5685
rect 3840 5629 3842 5689
rect 3838 5628 3844 5629
rect 4468 5628 4470 5689
rect 4604 5628 4606 5689
rect 4740 5628 4742 5689
rect 4876 5628 4878 5689
rect 5664 5629 5666 5689
rect 5662 5628 5668 5629
rect 3798 5624 3804 5625
rect 1974 5620 1975 5624
rect 1979 5620 1980 5624
rect 1974 5619 1980 5620
rect 1994 5623 2000 5624
rect 1994 5619 1995 5623
rect 1999 5619 2000 5623
rect 1994 5618 2000 5619
rect 2170 5623 2176 5624
rect 2170 5619 2171 5623
rect 2175 5619 2176 5623
rect 2170 5618 2176 5619
rect 2370 5623 2376 5624
rect 2370 5619 2371 5623
rect 2375 5619 2376 5623
rect 2370 5618 2376 5619
rect 2562 5623 2568 5624
rect 2562 5619 2563 5623
rect 2567 5619 2568 5623
rect 2562 5618 2568 5619
rect 2746 5623 2752 5624
rect 2746 5619 2747 5623
rect 2751 5619 2752 5623
rect 2746 5618 2752 5619
rect 2930 5623 2936 5624
rect 2930 5619 2931 5623
rect 2935 5619 2936 5623
rect 2930 5618 2936 5619
rect 3106 5623 3112 5624
rect 3106 5619 3107 5623
rect 3111 5619 3112 5623
rect 3106 5618 3112 5619
rect 3274 5623 3280 5624
rect 3274 5619 3275 5623
rect 3279 5619 3280 5623
rect 3274 5618 3280 5619
rect 3442 5623 3448 5624
rect 3442 5619 3443 5623
rect 3447 5619 3448 5623
rect 3442 5618 3448 5619
rect 3618 5623 3624 5624
rect 3618 5619 3619 5623
rect 3623 5619 3624 5623
rect 3798 5620 3799 5624
rect 3803 5620 3804 5624
rect 3838 5624 3839 5628
rect 3843 5624 3844 5628
rect 3838 5623 3844 5624
rect 4466 5627 4472 5628
rect 4466 5623 4467 5627
rect 4471 5623 4472 5627
rect 4466 5622 4472 5623
rect 4602 5627 4608 5628
rect 4602 5623 4603 5627
rect 4607 5623 4608 5627
rect 4602 5622 4608 5623
rect 4738 5627 4744 5628
rect 4738 5623 4739 5627
rect 4743 5623 4744 5627
rect 4738 5622 4744 5623
rect 4874 5627 4880 5628
rect 4874 5623 4875 5627
rect 4879 5623 4880 5627
rect 5662 5624 5663 5628
rect 5667 5624 5668 5628
rect 5662 5623 5668 5624
rect 4874 5622 4880 5623
rect 3798 5619 3804 5620
rect 3618 5618 3624 5619
rect 1934 5617 1940 5618
rect 110 5613 111 5617
rect 115 5613 116 5617
rect 110 5612 116 5613
rect 342 5616 348 5617
rect 342 5612 343 5616
rect 347 5612 348 5616
rect 342 5611 348 5612
rect 534 5616 540 5617
rect 534 5612 535 5616
rect 539 5612 540 5616
rect 534 5611 540 5612
rect 734 5616 740 5617
rect 734 5612 735 5616
rect 739 5612 740 5616
rect 734 5611 740 5612
rect 942 5616 948 5617
rect 942 5612 943 5616
rect 947 5612 948 5616
rect 942 5611 948 5612
rect 1158 5616 1164 5617
rect 1158 5612 1159 5616
rect 1163 5612 1164 5616
rect 1158 5611 1164 5612
rect 1382 5616 1388 5617
rect 1382 5612 1383 5616
rect 1387 5612 1388 5616
rect 1382 5611 1388 5612
rect 1606 5616 1612 5617
rect 1606 5612 1607 5616
rect 1611 5612 1612 5616
rect 1606 5611 1612 5612
rect 1814 5616 1820 5617
rect 1814 5612 1815 5616
rect 1819 5612 1820 5616
rect 1934 5613 1935 5617
rect 1939 5613 1940 5617
rect 1934 5612 1940 5613
rect 4494 5612 4500 5613
rect 1814 5611 1820 5612
rect 3838 5611 3844 5612
rect 2022 5608 2028 5609
rect 1974 5607 1980 5608
rect 1974 5603 1975 5607
rect 1979 5603 1980 5607
rect 2022 5604 2023 5608
rect 2027 5604 2028 5608
rect 2022 5603 2028 5604
rect 2198 5608 2204 5609
rect 2198 5604 2199 5608
rect 2203 5604 2204 5608
rect 2198 5603 2204 5604
rect 2398 5608 2404 5609
rect 2398 5604 2399 5608
rect 2403 5604 2404 5608
rect 2398 5603 2404 5604
rect 2590 5608 2596 5609
rect 2590 5604 2591 5608
rect 2595 5604 2596 5608
rect 2590 5603 2596 5604
rect 2774 5608 2780 5609
rect 2774 5604 2775 5608
rect 2779 5604 2780 5608
rect 2774 5603 2780 5604
rect 2958 5608 2964 5609
rect 2958 5604 2959 5608
rect 2963 5604 2964 5608
rect 2958 5603 2964 5604
rect 3134 5608 3140 5609
rect 3134 5604 3135 5608
rect 3139 5604 3140 5608
rect 3134 5603 3140 5604
rect 3302 5608 3308 5609
rect 3302 5604 3303 5608
rect 3307 5604 3308 5608
rect 3302 5603 3308 5604
rect 3470 5608 3476 5609
rect 3470 5604 3471 5608
rect 3475 5604 3476 5608
rect 3470 5603 3476 5604
rect 3646 5608 3652 5609
rect 3646 5604 3647 5608
rect 3651 5604 3652 5608
rect 3646 5603 3652 5604
rect 3798 5607 3804 5608
rect 3798 5603 3799 5607
rect 3803 5603 3804 5607
rect 3838 5607 3839 5611
rect 3843 5607 3844 5611
rect 4494 5608 4495 5612
rect 4499 5608 4500 5612
rect 4494 5607 4500 5608
rect 4630 5612 4636 5613
rect 4630 5608 4631 5612
rect 4635 5608 4636 5612
rect 4630 5607 4636 5608
rect 4766 5612 4772 5613
rect 4766 5608 4767 5612
rect 4771 5608 4772 5612
rect 4766 5607 4772 5608
rect 4902 5612 4908 5613
rect 4902 5608 4903 5612
rect 4907 5608 4908 5612
rect 4902 5607 4908 5608
rect 5662 5611 5668 5612
rect 5662 5607 5663 5611
rect 5667 5607 5668 5611
rect 3838 5606 3844 5607
rect 1974 5602 1980 5603
rect 314 5601 320 5602
rect 110 5600 116 5601
rect 110 5596 111 5600
rect 115 5596 116 5600
rect 314 5597 315 5601
rect 319 5597 320 5601
rect 314 5596 320 5597
rect 506 5601 512 5602
rect 506 5597 507 5601
rect 511 5597 512 5601
rect 506 5596 512 5597
rect 706 5601 712 5602
rect 706 5597 707 5601
rect 711 5597 712 5601
rect 706 5596 712 5597
rect 914 5601 920 5602
rect 914 5597 915 5601
rect 919 5597 920 5601
rect 914 5596 920 5597
rect 1130 5601 1136 5602
rect 1130 5597 1131 5601
rect 1135 5597 1136 5601
rect 1130 5596 1136 5597
rect 1354 5601 1360 5602
rect 1354 5597 1355 5601
rect 1359 5597 1360 5601
rect 1354 5596 1360 5597
rect 1578 5601 1584 5602
rect 1578 5597 1579 5601
rect 1583 5597 1584 5601
rect 1578 5596 1584 5597
rect 1786 5601 1792 5602
rect 1786 5597 1787 5601
rect 1791 5597 1792 5601
rect 1786 5596 1792 5597
rect 1934 5600 1940 5601
rect 1934 5596 1935 5600
rect 1939 5596 1940 5600
rect 110 5595 116 5596
rect 112 5535 114 5595
rect 316 5535 318 5596
rect 508 5535 510 5596
rect 708 5535 710 5596
rect 916 5535 918 5596
rect 1132 5535 1134 5596
rect 1356 5535 1358 5596
rect 1580 5535 1582 5596
rect 1788 5535 1790 5596
rect 1934 5595 1940 5596
rect 1936 5535 1938 5595
rect 1976 5579 1978 5602
rect 2024 5579 2026 5603
rect 2200 5579 2202 5603
rect 2400 5579 2402 5603
rect 2592 5579 2594 5603
rect 2776 5579 2778 5603
rect 2960 5579 2962 5603
rect 3136 5579 3138 5603
rect 3304 5579 3306 5603
rect 3472 5579 3474 5603
rect 3648 5579 3650 5603
rect 3798 5602 3804 5603
rect 3800 5579 3802 5602
rect 3840 5583 3842 5606
rect 4496 5583 4498 5607
rect 4632 5583 4634 5607
rect 4768 5583 4770 5607
rect 4904 5583 4906 5607
rect 5662 5606 5668 5607
rect 5664 5583 5666 5606
rect 3839 5582 3843 5583
rect 1975 5578 1979 5579
rect 1975 5573 1979 5574
rect 2023 5578 2027 5579
rect 2023 5573 2027 5574
rect 2199 5578 2203 5579
rect 2199 5573 2203 5574
rect 2375 5578 2379 5579
rect 2375 5573 2379 5574
rect 2399 5578 2403 5579
rect 2399 5573 2403 5574
rect 2591 5578 2595 5579
rect 2591 5573 2595 5574
rect 2607 5578 2611 5579
rect 2607 5573 2611 5574
rect 2775 5578 2779 5579
rect 2775 5573 2779 5574
rect 2831 5578 2835 5579
rect 2831 5573 2835 5574
rect 2959 5578 2963 5579
rect 2959 5573 2963 5574
rect 3047 5578 3051 5579
rect 3047 5573 3051 5574
rect 3135 5578 3139 5579
rect 3135 5573 3139 5574
rect 3263 5578 3267 5579
rect 3263 5573 3267 5574
rect 3303 5578 3307 5579
rect 3303 5573 3307 5574
rect 3471 5578 3475 5579
rect 3471 5573 3475 5574
rect 3479 5578 3483 5579
rect 3479 5573 3483 5574
rect 3647 5578 3651 5579
rect 3647 5573 3651 5574
rect 3679 5578 3683 5579
rect 3679 5573 3683 5574
rect 3799 5578 3803 5579
rect 3839 5577 3843 5578
rect 4431 5582 4435 5583
rect 4431 5577 4435 5578
rect 4495 5582 4499 5583
rect 4495 5577 4499 5578
rect 4567 5582 4571 5583
rect 4567 5577 4571 5578
rect 4631 5582 4635 5583
rect 4631 5577 4635 5578
rect 4703 5582 4707 5583
rect 4703 5577 4707 5578
rect 4767 5582 4771 5583
rect 4767 5577 4771 5578
rect 4839 5582 4843 5583
rect 4839 5577 4843 5578
rect 4903 5582 4907 5583
rect 4903 5577 4907 5578
rect 4975 5582 4979 5583
rect 4975 5577 4979 5578
rect 5111 5582 5115 5583
rect 5111 5577 5115 5578
rect 5663 5582 5667 5583
rect 5663 5577 5667 5578
rect 3799 5573 3803 5574
rect 1976 5550 1978 5573
rect 1974 5549 1980 5550
rect 2376 5549 2378 5573
rect 2608 5549 2610 5573
rect 2832 5549 2834 5573
rect 3048 5549 3050 5573
rect 3264 5549 3266 5573
rect 3480 5549 3482 5573
rect 3680 5549 3682 5573
rect 3800 5550 3802 5573
rect 3840 5554 3842 5577
rect 3838 5553 3844 5554
rect 4432 5553 4434 5577
rect 4568 5553 4570 5577
rect 4704 5553 4706 5577
rect 4840 5553 4842 5577
rect 4976 5553 4978 5577
rect 5112 5553 5114 5577
rect 5664 5554 5666 5577
rect 5662 5553 5668 5554
rect 3798 5549 3804 5550
rect 1974 5545 1975 5549
rect 1979 5545 1980 5549
rect 1974 5544 1980 5545
rect 2374 5548 2380 5549
rect 2374 5544 2375 5548
rect 2379 5544 2380 5548
rect 2374 5543 2380 5544
rect 2606 5548 2612 5549
rect 2606 5544 2607 5548
rect 2611 5544 2612 5548
rect 2606 5543 2612 5544
rect 2830 5548 2836 5549
rect 2830 5544 2831 5548
rect 2835 5544 2836 5548
rect 2830 5543 2836 5544
rect 3046 5548 3052 5549
rect 3046 5544 3047 5548
rect 3051 5544 3052 5548
rect 3046 5543 3052 5544
rect 3262 5548 3268 5549
rect 3262 5544 3263 5548
rect 3267 5544 3268 5548
rect 3262 5543 3268 5544
rect 3478 5548 3484 5549
rect 3478 5544 3479 5548
rect 3483 5544 3484 5548
rect 3478 5543 3484 5544
rect 3678 5548 3684 5549
rect 3678 5544 3679 5548
rect 3683 5544 3684 5548
rect 3798 5545 3799 5549
rect 3803 5545 3804 5549
rect 3838 5549 3839 5553
rect 3843 5549 3844 5553
rect 3838 5548 3844 5549
rect 4430 5552 4436 5553
rect 4430 5548 4431 5552
rect 4435 5548 4436 5552
rect 4430 5547 4436 5548
rect 4566 5552 4572 5553
rect 4566 5548 4567 5552
rect 4571 5548 4572 5552
rect 4566 5547 4572 5548
rect 4702 5552 4708 5553
rect 4702 5548 4703 5552
rect 4707 5548 4708 5552
rect 4702 5547 4708 5548
rect 4838 5552 4844 5553
rect 4838 5548 4839 5552
rect 4843 5548 4844 5552
rect 4838 5547 4844 5548
rect 4974 5552 4980 5553
rect 4974 5548 4975 5552
rect 4979 5548 4980 5552
rect 4974 5547 4980 5548
rect 5110 5552 5116 5553
rect 5110 5548 5111 5552
rect 5115 5548 5116 5552
rect 5662 5549 5663 5553
rect 5667 5549 5668 5553
rect 5662 5548 5668 5549
rect 5110 5547 5116 5548
rect 3798 5544 3804 5545
rect 3678 5543 3684 5544
rect 4402 5537 4408 5538
rect 3838 5536 3844 5537
rect 111 5534 115 5535
rect 111 5529 115 5530
rect 315 5534 319 5535
rect 315 5529 319 5530
rect 507 5534 511 5535
rect 507 5529 511 5530
rect 707 5534 711 5535
rect 707 5529 711 5530
rect 875 5534 879 5535
rect 875 5529 879 5530
rect 915 5534 919 5535
rect 915 5529 919 5530
rect 1011 5534 1015 5535
rect 1011 5529 1015 5530
rect 1131 5534 1135 5535
rect 1131 5529 1135 5530
rect 1147 5534 1151 5535
rect 1147 5529 1151 5530
rect 1291 5534 1295 5535
rect 1291 5529 1295 5530
rect 1355 5534 1359 5535
rect 1355 5529 1359 5530
rect 1435 5534 1439 5535
rect 1435 5529 1439 5530
rect 1579 5534 1583 5535
rect 1579 5529 1583 5530
rect 1723 5534 1727 5535
rect 1723 5529 1727 5530
rect 1787 5534 1791 5535
rect 1787 5529 1791 5530
rect 1935 5534 1939 5535
rect 2346 5533 2352 5534
rect 1935 5529 1939 5530
rect 1974 5532 1980 5533
rect 112 5469 114 5529
rect 110 5468 116 5469
rect 876 5468 878 5529
rect 1012 5468 1014 5529
rect 1148 5468 1150 5529
rect 1292 5468 1294 5529
rect 1436 5468 1438 5529
rect 1580 5468 1582 5529
rect 1724 5468 1726 5529
rect 1936 5469 1938 5529
rect 1974 5528 1975 5532
rect 1979 5528 1980 5532
rect 2346 5529 2347 5533
rect 2351 5529 2352 5533
rect 2346 5528 2352 5529
rect 2578 5533 2584 5534
rect 2578 5529 2579 5533
rect 2583 5529 2584 5533
rect 2578 5528 2584 5529
rect 2802 5533 2808 5534
rect 2802 5529 2803 5533
rect 2807 5529 2808 5533
rect 2802 5528 2808 5529
rect 3018 5533 3024 5534
rect 3018 5529 3019 5533
rect 3023 5529 3024 5533
rect 3018 5528 3024 5529
rect 3234 5533 3240 5534
rect 3234 5529 3235 5533
rect 3239 5529 3240 5533
rect 3234 5528 3240 5529
rect 3450 5533 3456 5534
rect 3450 5529 3451 5533
rect 3455 5529 3456 5533
rect 3450 5528 3456 5529
rect 3650 5533 3656 5534
rect 3650 5529 3651 5533
rect 3655 5529 3656 5533
rect 3650 5528 3656 5529
rect 3798 5532 3804 5533
rect 3798 5528 3799 5532
rect 3803 5528 3804 5532
rect 3838 5532 3839 5536
rect 3843 5532 3844 5536
rect 4402 5533 4403 5537
rect 4407 5533 4408 5537
rect 4402 5532 4408 5533
rect 4538 5537 4544 5538
rect 4538 5533 4539 5537
rect 4543 5533 4544 5537
rect 4538 5532 4544 5533
rect 4674 5537 4680 5538
rect 4674 5533 4675 5537
rect 4679 5533 4680 5537
rect 4674 5532 4680 5533
rect 4810 5537 4816 5538
rect 4810 5533 4811 5537
rect 4815 5533 4816 5537
rect 4810 5532 4816 5533
rect 4946 5537 4952 5538
rect 4946 5533 4947 5537
rect 4951 5533 4952 5537
rect 4946 5532 4952 5533
rect 5082 5537 5088 5538
rect 5082 5533 5083 5537
rect 5087 5533 5088 5537
rect 5082 5532 5088 5533
rect 5662 5536 5668 5537
rect 5662 5532 5663 5536
rect 5667 5532 5668 5536
rect 3838 5531 3844 5532
rect 1974 5527 1980 5528
rect 1934 5468 1940 5469
rect 110 5464 111 5468
rect 115 5464 116 5468
rect 110 5463 116 5464
rect 874 5467 880 5468
rect 874 5463 875 5467
rect 879 5463 880 5467
rect 874 5462 880 5463
rect 1010 5467 1016 5468
rect 1010 5463 1011 5467
rect 1015 5463 1016 5467
rect 1010 5462 1016 5463
rect 1146 5467 1152 5468
rect 1146 5463 1147 5467
rect 1151 5463 1152 5467
rect 1146 5462 1152 5463
rect 1290 5467 1296 5468
rect 1290 5463 1291 5467
rect 1295 5463 1296 5467
rect 1290 5462 1296 5463
rect 1434 5467 1440 5468
rect 1434 5463 1435 5467
rect 1439 5463 1440 5467
rect 1434 5462 1440 5463
rect 1578 5467 1584 5468
rect 1578 5463 1579 5467
rect 1583 5463 1584 5467
rect 1578 5462 1584 5463
rect 1722 5467 1728 5468
rect 1722 5463 1723 5467
rect 1727 5463 1728 5467
rect 1934 5464 1935 5468
rect 1939 5464 1940 5468
rect 1934 5463 1940 5464
rect 1976 5463 1978 5527
rect 2348 5463 2350 5528
rect 2580 5463 2582 5528
rect 2804 5463 2806 5528
rect 3020 5463 3022 5528
rect 3236 5463 3238 5528
rect 3452 5463 3454 5528
rect 3652 5463 3654 5528
rect 3798 5527 3804 5528
rect 3800 5463 3802 5527
rect 3840 5471 3842 5531
rect 4404 5471 4406 5532
rect 4540 5471 4542 5532
rect 4676 5471 4678 5532
rect 4812 5471 4814 5532
rect 4948 5471 4950 5532
rect 5084 5471 5086 5532
rect 5662 5531 5668 5532
rect 5664 5471 5666 5531
rect 3839 5470 3843 5471
rect 3839 5465 3843 5466
rect 4403 5470 4407 5471
rect 4403 5465 4407 5466
rect 4427 5470 4431 5471
rect 4427 5465 4431 5466
rect 4539 5470 4543 5471
rect 4539 5465 4543 5466
rect 4587 5470 4591 5471
rect 4587 5465 4591 5466
rect 4675 5470 4679 5471
rect 4675 5465 4679 5466
rect 4747 5470 4751 5471
rect 4747 5465 4751 5466
rect 4811 5470 4815 5471
rect 4811 5465 4815 5466
rect 4907 5470 4911 5471
rect 4907 5465 4911 5466
rect 4947 5470 4951 5471
rect 4947 5465 4951 5466
rect 5075 5470 5079 5471
rect 5075 5465 5079 5466
rect 5083 5470 5087 5471
rect 5083 5465 5087 5466
rect 5663 5470 5667 5471
rect 5663 5465 5667 5466
rect 1722 5462 1728 5463
rect 1975 5462 1979 5463
rect 1975 5457 1979 5458
rect 2347 5462 2351 5463
rect 2347 5457 2351 5458
rect 2451 5462 2455 5463
rect 2451 5457 2455 5458
rect 2579 5462 2583 5463
rect 2579 5457 2583 5458
rect 2699 5462 2703 5463
rect 2699 5457 2703 5458
rect 2803 5462 2807 5463
rect 2803 5457 2807 5458
rect 2947 5462 2951 5463
rect 2947 5457 2951 5458
rect 3019 5462 3023 5463
rect 3019 5457 3023 5458
rect 3187 5462 3191 5463
rect 3187 5457 3191 5458
rect 3235 5462 3239 5463
rect 3235 5457 3239 5458
rect 3427 5462 3431 5463
rect 3427 5457 3431 5458
rect 3451 5462 3455 5463
rect 3451 5457 3455 5458
rect 3651 5462 3655 5463
rect 3651 5457 3655 5458
rect 3799 5462 3803 5463
rect 3799 5457 3803 5458
rect 902 5452 908 5453
rect 110 5451 116 5452
rect 110 5447 111 5451
rect 115 5447 116 5451
rect 902 5448 903 5452
rect 907 5448 908 5452
rect 902 5447 908 5448
rect 1038 5452 1044 5453
rect 1038 5448 1039 5452
rect 1043 5448 1044 5452
rect 1038 5447 1044 5448
rect 1174 5452 1180 5453
rect 1174 5448 1175 5452
rect 1179 5448 1180 5452
rect 1174 5447 1180 5448
rect 1318 5452 1324 5453
rect 1318 5448 1319 5452
rect 1323 5448 1324 5452
rect 1318 5447 1324 5448
rect 1462 5452 1468 5453
rect 1462 5448 1463 5452
rect 1467 5448 1468 5452
rect 1462 5447 1468 5448
rect 1606 5452 1612 5453
rect 1606 5448 1607 5452
rect 1611 5448 1612 5452
rect 1606 5447 1612 5448
rect 1750 5452 1756 5453
rect 1750 5448 1751 5452
rect 1755 5448 1756 5452
rect 1750 5447 1756 5448
rect 1934 5451 1940 5452
rect 1934 5447 1935 5451
rect 1939 5447 1940 5451
rect 110 5446 116 5447
rect 112 5423 114 5446
rect 904 5423 906 5447
rect 1040 5423 1042 5447
rect 1176 5423 1178 5447
rect 1320 5423 1322 5447
rect 1464 5423 1466 5447
rect 1608 5423 1610 5447
rect 1752 5423 1754 5447
rect 1934 5446 1940 5447
rect 1936 5423 1938 5446
rect 111 5422 115 5423
rect 111 5417 115 5418
rect 719 5422 723 5423
rect 719 5417 723 5418
rect 855 5422 859 5423
rect 855 5417 859 5418
rect 903 5422 907 5423
rect 903 5417 907 5418
rect 991 5422 995 5423
rect 991 5417 995 5418
rect 1039 5422 1043 5423
rect 1039 5417 1043 5418
rect 1127 5422 1131 5423
rect 1127 5417 1131 5418
rect 1175 5422 1179 5423
rect 1175 5417 1179 5418
rect 1263 5422 1267 5423
rect 1263 5417 1267 5418
rect 1319 5422 1323 5423
rect 1319 5417 1323 5418
rect 1399 5422 1403 5423
rect 1399 5417 1403 5418
rect 1463 5422 1467 5423
rect 1463 5417 1467 5418
rect 1535 5422 1539 5423
rect 1535 5417 1539 5418
rect 1607 5422 1611 5423
rect 1607 5417 1611 5418
rect 1671 5422 1675 5423
rect 1671 5417 1675 5418
rect 1751 5422 1755 5423
rect 1751 5417 1755 5418
rect 1807 5422 1811 5423
rect 1807 5417 1811 5418
rect 1935 5422 1939 5423
rect 1935 5417 1939 5418
rect 112 5394 114 5417
rect 110 5393 116 5394
rect 720 5393 722 5417
rect 856 5393 858 5417
rect 992 5393 994 5417
rect 1128 5393 1130 5417
rect 1264 5393 1266 5417
rect 1400 5393 1402 5417
rect 1536 5393 1538 5417
rect 1672 5393 1674 5417
rect 1808 5393 1810 5417
rect 1936 5394 1938 5417
rect 1976 5397 1978 5457
rect 1974 5396 1980 5397
rect 2452 5396 2454 5457
rect 2700 5396 2702 5457
rect 2948 5396 2950 5457
rect 3188 5396 3190 5457
rect 3428 5396 3430 5457
rect 3652 5396 3654 5457
rect 3800 5397 3802 5457
rect 3840 5405 3842 5465
rect 3838 5404 3844 5405
rect 4428 5404 4430 5465
rect 4588 5404 4590 5465
rect 4748 5404 4750 5465
rect 4908 5404 4910 5465
rect 5076 5404 5078 5465
rect 5664 5405 5666 5465
rect 5662 5404 5668 5405
rect 3838 5400 3839 5404
rect 3843 5400 3844 5404
rect 3838 5399 3844 5400
rect 4426 5403 4432 5404
rect 4426 5399 4427 5403
rect 4431 5399 4432 5403
rect 4426 5398 4432 5399
rect 4586 5403 4592 5404
rect 4586 5399 4587 5403
rect 4591 5399 4592 5403
rect 4586 5398 4592 5399
rect 4746 5403 4752 5404
rect 4746 5399 4747 5403
rect 4751 5399 4752 5403
rect 4746 5398 4752 5399
rect 4906 5403 4912 5404
rect 4906 5399 4907 5403
rect 4911 5399 4912 5403
rect 4906 5398 4912 5399
rect 5074 5403 5080 5404
rect 5074 5399 5075 5403
rect 5079 5399 5080 5403
rect 5662 5400 5663 5404
rect 5667 5400 5668 5404
rect 5662 5399 5668 5400
rect 5074 5398 5080 5399
rect 3798 5396 3804 5397
rect 1934 5393 1940 5394
rect 110 5389 111 5393
rect 115 5389 116 5393
rect 110 5388 116 5389
rect 718 5392 724 5393
rect 718 5388 719 5392
rect 723 5388 724 5392
rect 718 5387 724 5388
rect 854 5392 860 5393
rect 854 5388 855 5392
rect 859 5388 860 5392
rect 854 5387 860 5388
rect 990 5392 996 5393
rect 990 5388 991 5392
rect 995 5388 996 5392
rect 990 5387 996 5388
rect 1126 5392 1132 5393
rect 1126 5388 1127 5392
rect 1131 5388 1132 5392
rect 1126 5387 1132 5388
rect 1262 5392 1268 5393
rect 1262 5388 1263 5392
rect 1267 5388 1268 5392
rect 1262 5387 1268 5388
rect 1398 5392 1404 5393
rect 1398 5388 1399 5392
rect 1403 5388 1404 5392
rect 1398 5387 1404 5388
rect 1534 5392 1540 5393
rect 1534 5388 1535 5392
rect 1539 5388 1540 5392
rect 1534 5387 1540 5388
rect 1670 5392 1676 5393
rect 1670 5388 1671 5392
rect 1675 5388 1676 5392
rect 1670 5387 1676 5388
rect 1806 5392 1812 5393
rect 1806 5388 1807 5392
rect 1811 5388 1812 5392
rect 1934 5389 1935 5393
rect 1939 5389 1940 5393
rect 1974 5392 1975 5396
rect 1979 5392 1980 5396
rect 1974 5391 1980 5392
rect 2450 5395 2456 5396
rect 2450 5391 2451 5395
rect 2455 5391 2456 5395
rect 2450 5390 2456 5391
rect 2698 5395 2704 5396
rect 2698 5391 2699 5395
rect 2703 5391 2704 5395
rect 2698 5390 2704 5391
rect 2946 5395 2952 5396
rect 2946 5391 2947 5395
rect 2951 5391 2952 5395
rect 2946 5390 2952 5391
rect 3186 5395 3192 5396
rect 3186 5391 3187 5395
rect 3191 5391 3192 5395
rect 3186 5390 3192 5391
rect 3426 5395 3432 5396
rect 3426 5391 3427 5395
rect 3431 5391 3432 5395
rect 3426 5390 3432 5391
rect 3650 5395 3656 5396
rect 3650 5391 3651 5395
rect 3655 5391 3656 5395
rect 3798 5392 3799 5396
rect 3803 5392 3804 5396
rect 3798 5391 3804 5392
rect 3650 5390 3656 5391
rect 1934 5388 1940 5389
rect 4454 5388 4460 5389
rect 1806 5387 1812 5388
rect 3838 5387 3844 5388
rect 3838 5383 3839 5387
rect 3843 5383 3844 5387
rect 4454 5384 4455 5388
rect 4459 5384 4460 5388
rect 4454 5383 4460 5384
rect 4614 5388 4620 5389
rect 4614 5384 4615 5388
rect 4619 5384 4620 5388
rect 4614 5383 4620 5384
rect 4774 5388 4780 5389
rect 4774 5384 4775 5388
rect 4779 5384 4780 5388
rect 4774 5383 4780 5384
rect 4934 5388 4940 5389
rect 4934 5384 4935 5388
rect 4939 5384 4940 5388
rect 4934 5383 4940 5384
rect 5102 5388 5108 5389
rect 5102 5384 5103 5388
rect 5107 5384 5108 5388
rect 5102 5383 5108 5384
rect 5662 5387 5668 5388
rect 5662 5383 5663 5387
rect 5667 5383 5668 5387
rect 3838 5382 3844 5383
rect 2478 5380 2484 5381
rect 1974 5379 1980 5380
rect 690 5377 696 5378
rect 110 5376 116 5377
rect 110 5372 111 5376
rect 115 5372 116 5376
rect 690 5373 691 5377
rect 695 5373 696 5377
rect 690 5372 696 5373
rect 826 5377 832 5378
rect 826 5373 827 5377
rect 831 5373 832 5377
rect 826 5372 832 5373
rect 962 5377 968 5378
rect 962 5373 963 5377
rect 967 5373 968 5377
rect 962 5372 968 5373
rect 1098 5377 1104 5378
rect 1098 5373 1099 5377
rect 1103 5373 1104 5377
rect 1098 5372 1104 5373
rect 1234 5377 1240 5378
rect 1234 5373 1235 5377
rect 1239 5373 1240 5377
rect 1234 5372 1240 5373
rect 1370 5377 1376 5378
rect 1370 5373 1371 5377
rect 1375 5373 1376 5377
rect 1370 5372 1376 5373
rect 1506 5377 1512 5378
rect 1506 5373 1507 5377
rect 1511 5373 1512 5377
rect 1506 5372 1512 5373
rect 1642 5377 1648 5378
rect 1642 5373 1643 5377
rect 1647 5373 1648 5377
rect 1642 5372 1648 5373
rect 1778 5377 1784 5378
rect 1778 5373 1779 5377
rect 1783 5373 1784 5377
rect 1778 5372 1784 5373
rect 1934 5376 1940 5377
rect 1934 5372 1935 5376
rect 1939 5372 1940 5376
rect 1974 5375 1975 5379
rect 1979 5375 1980 5379
rect 2478 5376 2479 5380
rect 2483 5376 2484 5380
rect 2478 5375 2484 5376
rect 2726 5380 2732 5381
rect 2726 5376 2727 5380
rect 2731 5376 2732 5380
rect 2726 5375 2732 5376
rect 2974 5380 2980 5381
rect 2974 5376 2975 5380
rect 2979 5376 2980 5380
rect 2974 5375 2980 5376
rect 3214 5380 3220 5381
rect 3214 5376 3215 5380
rect 3219 5376 3220 5380
rect 3214 5375 3220 5376
rect 3454 5380 3460 5381
rect 3454 5376 3455 5380
rect 3459 5376 3460 5380
rect 3454 5375 3460 5376
rect 3678 5380 3684 5381
rect 3678 5376 3679 5380
rect 3683 5376 3684 5380
rect 3678 5375 3684 5376
rect 3798 5379 3804 5380
rect 3798 5375 3799 5379
rect 3803 5375 3804 5379
rect 1974 5374 1980 5375
rect 110 5371 116 5372
rect 112 5311 114 5371
rect 692 5311 694 5372
rect 828 5311 830 5372
rect 964 5311 966 5372
rect 1100 5311 1102 5372
rect 1236 5311 1238 5372
rect 1372 5311 1374 5372
rect 1508 5311 1510 5372
rect 1644 5311 1646 5372
rect 1780 5311 1782 5372
rect 1934 5371 1940 5372
rect 1936 5311 1938 5371
rect 1976 5351 1978 5374
rect 2480 5351 2482 5375
rect 2728 5351 2730 5375
rect 2976 5351 2978 5375
rect 3216 5351 3218 5375
rect 3456 5351 3458 5375
rect 3680 5351 3682 5375
rect 3798 5374 3804 5375
rect 3800 5351 3802 5374
rect 3840 5351 3842 5382
rect 4456 5351 4458 5383
rect 4616 5351 4618 5383
rect 4776 5351 4778 5383
rect 4936 5351 4938 5383
rect 5104 5351 5106 5383
rect 5662 5382 5668 5383
rect 5664 5351 5666 5382
rect 1975 5350 1979 5351
rect 1975 5345 1979 5346
rect 2319 5350 2323 5351
rect 2319 5345 2323 5346
rect 2479 5350 2483 5351
rect 2479 5345 2483 5346
rect 2519 5350 2523 5351
rect 2519 5345 2523 5346
rect 2719 5350 2723 5351
rect 2719 5345 2723 5346
rect 2727 5350 2731 5351
rect 2727 5345 2731 5346
rect 2919 5350 2923 5351
rect 2919 5345 2923 5346
rect 2975 5350 2979 5351
rect 2975 5345 2979 5346
rect 3119 5350 3123 5351
rect 3119 5345 3123 5346
rect 3215 5350 3219 5351
rect 3215 5345 3219 5346
rect 3327 5350 3331 5351
rect 3327 5345 3331 5346
rect 3455 5350 3459 5351
rect 3455 5345 3459 5346
rect 3535 5350 3539 5351
rect 3535 5345 3539 5346
rect 3679 5350 3683 5351
rect 3679 5345 3683 5346
rect 3799 5350 3803 5351
rect 3799 5345 3803 5346
rect 3839 5350 3843 5351
rect 3839 5345 3843 5346
rect 4431 5350 4435 5351
rect 4431 5345 4435 5346
rect 4455 5350 4459 5351
rect 4455 5345 4459 5346
rect 4615 5350 4619 5351
rect 4615 5345 4619 5346
rect 4775 5350 4779 5351
rect 4775 5345 4779 5346
rect 4799 5350 4803 5351
rect 4799 5345 4803 5346
rect 4935 5350 4939 5351
rect 4935 5345 4939 5346
rect 4983 5350 4987 5351
rect 4983 5345 4987 5346
rect 5103 5350 5107 5351
rect 5103 5345 5107 5346
rect 5175 5350 5179 5351
rect 5175 5345 5179 5346
rect 5663 5350 5667 5351
rect 5663 5345 5667 5346
rect 1976 5322 1978 5345
rect 1974 5321 1980 5322
rect 2320 5321 2322 5345
rect 2520 5321 2522 5345
rect 2720 5321 2722 5345
rect 2920 5321 2922 5345
rect 3120 5321 3122 5345
rect 3328 5321 3330 5345
rect 3536 5321 3538 5345
rect 3800 5322 3802 5345
rect 3840 5322 3842 5345
rect 3798 5321 3804 5322
rect 1974 5317 1975 5321
rect 1979 5317 1980 5321
rect 1974 5316 1980 5317
rect 2318 5320 2324 5321
rect 2318 5316 2319 5320
rect 2323 5316 2324 5320
rect 2318 5315 2324 5316
rect 2518 5320 2524 5321
rect 2518 5316 2519 5320
rect 2523 5316 2524 5320
rect 2518 5315 2524 5316
rect 2718 5320 2724 5321
rect 2718 5316 2719 5320
rect 2723 5316 2724 5320
rect 2718 5315 2724 5316
rect 2918 5320 2924 5321
rect 2918 5316 2919 5320
rect 2923 5316 2924 5320
rect 2918 5315 2924 5316
rect 3118 5320 3124 5321
rect 3118 5316 3119 5320
rect 3123 5316 3124 5320
rect 3118 5315 3124 5316
rect 3326 5320 3332 5321
rect 3326 5316 3327 5320
rect 3331 5316 3332 5320
rect 3326 5315 3332 5316
rect 3534 5320 3540 5321
rect 3534 5316 3535 5320
rect 3539 5316 3540 5320
rect 3798 5317 3799 5321
rect 3803 5317 3804 5321
rect 3798 5316 3804 5317
rect 3838 5321 3844 5322
rect 4432 5321 4434 5345
rect 4616 5321 4618 5345
rect 4800 5321 4802 5345
rect 4984 5321 4986 5345
rect 5176 5321 5178 5345
rect 5664 5322 5666 5345
rect 5662 5321 5668 5322
rect 3838 5317 3839 5321
rect 3843 5317 3844 5321
rect 3838 5316 3844 5317
rect 4430 5320 4436 5321
rect 4430 5316 4431 5320
rect 4435 5316 4436 5320
rect 3534 5315 3540 5316
rect 4430 5315 4436 5316
rect 4614 5320 4620 5321
rect 4614 5316 4615 5320
rect 4619 5316 4620 5320
rect 4614 5315 4620 5316
rect 4798 5320 4804 5321
rect 4798 5316 4799 5320
rect 4803 5316 4804 5320
rect 4798 5315 4804 5316
rect 4982 5320 4988 5321
rect 4982 5316 4983 5320
rect 4987 5316 4988 5320
rect 4982 5315 4988 5316
rect 5174 5320 5180 5321
rect 5174 5316 5175 5320
rect 5179 5316 5180 5320
rect 5662 5317 5663 5321
rect 5667 5317 5668 5321
rect 5662 5316 5668 5317
rect 5174 5315 5180 5316
rect 111 5310 115 5311
rect 111 5305 115 5306
rect 691 5310 695 5311
rect 691 5305 695 5306
rect 723 5310 727 5311
rect 723 5305 727 5306
rect 827 5310 831 5311
rect 827 5305 831 5306
rect 875 5310 879 5311
rect 875 5305 879 5306
rect 963 5310 967 5311
rect 963 5305 967 5306
rect 1027 5310 1031 5311
rect 1027 5305 1031 5306
rect 1099 5310 1103 5311
rect 1099 5305 1103 5306
rect 1187 5310 1191 5311
rect 1187 5305 1191 5306
rect 1235 5310 1239 5311
rect 1235 5305 1239 5306
rect 1355 5310 1359 5311
rect 1355 5305 1359 5306
rect 1371 5310 1375 5311
rect 1371 5305 1375 5306
rect 1507 5310 1511 5311
rect 1507 5305 1511 5306
rect 1523 5310 1527 5311
rect 1523 5305 1527 5306
rect 1643 5310 1647 5311
rect 1643 5305 1647 5306
rect 1779 5310 1783 5311
rect 1779 5305 1783 5306
rect 1935 5310 1939 5311
rect 1935 5305 1939 5306
rect 2290 5305 2296 5306
rect 112 5245 114 5305
rect 110 5244 116 5245
rect 724 5244 726 5305
rect 876 5244 878 5305
rect 1028 5244 1030 5305
rect 1188 5244 1190 5305
rect 1356 5244 1358 5305
rect 1524 5244 1526 5305
rect 1936 5245 1938 5305
rect 1974 5304 1980 5305
rect 1974 5300 1975 5304
rect 1979 5300 1980 5304
rect 2290 5301 2291 5305
rect 2295 5301 2296 5305
rect 2290 5300 2296 5301
rect 2490 5305 2496 5306
rect 2490 5301 2491 5305
rect 2495 5301 2496 5305
rect 2490 5300 2496 5301
rect 2690 5305 2696 5306
rect 2690 5301 2691 5305
rect 2695 5301 2696 5305
rect 2690 5300 2696 5301
rect 2890 5305 2896 5306
rect 2890 5301 2891 5305
rect 2895 5301 2896 5305
rect 2890 5300 2896 5301
rect 3090 5305 3096 5306
rect 3090 5301 3091 5305
rect 3095 5301 3096 5305
rect 3090 5300 3096 5301
rect 3298 5305 3304 5306
rect 3298 5301 3299 5305
rect 3303 5301 3304 5305
rect 3298 5300 3304 5301
rect 3506 5305 3512 5306
rect 4402 5305 4408 5306
rect 3506 5301 3507 5305
rect 3511 5301 3512 5305
rect 3506 5300 3512 5301
rect 3798 5304 3804 5305
rect 3798 5300 3799 5304
rect 3803 5300 3804 5304
rect 1974 5299 1980 5300
rect 1934 5244 1940 5245
rect 110 5240 111 5244
rect 115 5240 116 5244
rect 110 5239 116 5240
rect 722 5243 728 5244
rect 722 5239 723 5243
rect 727 5239 728 5243
rect 722 5238 728 5239
rect 874 5243 880 5244
rect 874 5239 875 5243
rect 879 5239 880 5243
rect 874 5238 880 5239
rect 1026 5243 1032 5244
rect 1026 5239 1027 5243
rect 1031 5239 1032 5243
rect 1026 5238 1032 5239
rect 1186 5243 1192 5244
rect 1186 5239 1187 5243
rect 1191 5239 1192 5243
rect 1186 5238 1192 5239
rect 1354 5243 1360 5244
rect 1354 5239 1355 5243
rect 1359 5239 1360 5243
rect 1354 5238 1360 5239
rect 1522 5243 1528 5244
rect 1522 5239 1523 5243
rect 1527 5239 1528 5243
rect 1934 5240 1935 5244
rect 1939 5240 1940 5244
rect 1934 5239 1940 5240
rect 1522 5238 1528 5239
rect 1976 5235 1978 5299
rect 2292 5235 2294 5300
rect 2492 5235 2494 5300
rect 2692 5235 2694 5300
rect 2892 5235 2894 5300
rect 3092 5235 3094 5300
rect 3300 5235 3302 5300
rect 3508 5235 3510 5300
rect 3798 5299 3804 5300
rect 3838 5304 3844 5305
rect 3838 5300 3839 5304
rect 3843 5300 3844 5304
rect 4402 5301 4403 5305
rect 4407 5301 4408 5305
rect 4402 5300 4408 5301
rect 4586 5305 4592 5306
rect 4586 5301 4587 5305
rect 4591 5301 4592 5305
rect 4586 5300 4592 5301
rect 4770 5305 4776 5306
rect 4770 5301 4771 5305
rect 4775 5301 4776 5305
rect 4770 5300 4776 5301
rect 4954 5305 4960 5306
rect 4954 5301 4955 5305
rect 4959 5301 4960 5305
rect 4954 5300 4960 5301
rect 5146 5305 5152 5306
rect 5146 5301 5147 5305
rect 5151 5301 5152 5305
rect 5146 5300 5152 5301
rect 5662 5304 5668 5305
rect 5662 5300 5663 5304
rect 5667 5300 5668 5304
rect 3838 5299 3844 5300
rect 3800 5235 3802 5299
rect 1975 5234 1979 5235
rect 1975 5229 1979 5230
rect 2275 5234 2279 5235
rect 2275 5229 2279 5230
rect 2291 5234 2295 5235
rect 2291 5229 2295 5230
rect 2475 5234 2479 5235
rect 2475 5229 2479 5230
rect 2491 5234 2495 5235
rect 2491 5229 2495 5230
rect 2683 5234 2687 5235
rect 2683 5229 2687 5230
rect 2691 5234 2695 5235
rect 2691 5229 2695 5230
rect 2891 5234 2895 5235
rect 2891 5229 2895 5230
rect 3091 5234 3095 5235
rect 3091 5229 3095 5230
rect 3099 5234 3103 5235
rect 3099 5229 3103 5230
rect 3299 5234 3303 5235
rect 3299 5229 3303 5230
rect 3307 5234 3311 5235
rect 3307 5229 3311 5230
rect 3507 5234 3511 5235
rect 3507 5229 3511 5230
rect 3799 5234 3803 5235
rect 3799 5229 3803 5230
rect 750 5228 756 5229
rect 110 5227 116 5228
rect 110 5223 111 5227
rect 115 5223 116 5227
rect 750 5224 751 5228
rect 755 5224 756 5228
rect 750 5223 756 5224
rect 902 5228 908 5229
rect 902 5224 903 5228
rect 907 5224 908 5228
rect 902 5223 908 5224
rect 1054 5228 1060 5229
rect 1054 5224 1055 5228
rect 1059 5224 1060 5228
rect 1054 5223 1060 5224
rect 1214 5228 1220 5229
rect 1214 5224 1215 5228
rect 1219 5224 1220 5228
rect 1214 5223 1220 5224
rect 1382 5228 1388 5229
rect 1382 5224 1383 5228
rect 1387 5224 1388 5228
rect 1382 5223 1388 5224
rect 1550 5228 1556 5229
rect 1550 5224 1551 5228
rect 1555 5224 1556 5228
rect 1550 5223 1556 5224
rect 1934 5227 1940 5228
rect 1934 5223 1935 5227
rect 1939 5223 1940 5227
rect 110 5222 116 5223
rect 112 5199 114 5222
rect 752 5199 754 5223
rect 904 5199 906 5223
rect 1056 5199 1058 5223
rect 1216 5199 1218 5223
rect 1384 5199 1386 5223
rect 1552 5199 1554 5223
rect 1934 5222 1940 5223
rect 1936 5199 1938 5222
rect 111 5198 115 5199
rect 111 5193 115 5194
rect 447 5198 451 5199
rect 447 5193 451 5194
rect 623 5198 627 5199
rect 623 5193 627 5194
rect 751 5198 755 5199
rect 751 5193 755 5194
rect 807 5198 811 5199
rect 807 5193 811 5194
rect 903 5198 907 5199
rect 903 5193 907 5194
rect 999 5198 1003 5199
rect 999 5193 1003 5194
rect 1055 5198 1059 5199
rect 1055 5193 1059 5194
rect 1199 5198 1203 5199
rect 1199 5193 1203 5194
rect 1215 5198 1219 5199
rect 1215 5193 1219 5194
rect 1383 5198 1387 5199
rect 1383 5193 1387 5194
rect 1399 5198 1403 5199
rect 1399 5193 1403 5194
rect 1551 5198 1555 5199
rect 1551 5193 1555 5194
rect 1607 5198 1611 5199
rect 1607 5193 1611 5194
rect 1815 5198 1819 5199
rect 1815 5193 1819 5194
rect 1935 5198 1939 5199
rect 1935 5193 1939 5194
rect 112 5170 114 5193
rect 110 5169 116 5170
rect 448 5169 450 5193
rect 624 5169 626 5193
rect 808 5169 810 5193
rect 1000 5169 1002 5193
rect 1200 5169 1202 5193
rect 1400 5169 1402 5193
rect 1608 5169 1610 5193
rect 1816 5169 1818 5193
rect 1936 5170 1938 5193
rect 1934 5169 1940 5170
rect 1976 5169 1978 5229
rect 110 5165 111 5169
rect 115 5165 116 5169
rect 110 5164 116 5165
rect 446 5168 452 5169
rect 446 5164 447 5168
rect 451 5164 452 5168
rect 446 5163 452 5164
rect 622 5168 628 5169
rect 622 5164 623 5168
rect 627 5164 628 5168
rect 622 5163 628 5164
rect 806 5168 812 5169
rect 806 5164 807 5168
rect 811 5164 812 5168
rect 806 5163 812 5164
rect 998 5168 1004 5169
rect 998 5164 999 5168
rect 1003 5164 1004 5168
rect 998 5163 1004 5164
rect 1198 5168 1204 5169
rect 1198 5164 1199 5168
rect 1203 5164 1204 5168
rect 1198 5163 1204 5164
rect 1398 5168 1404 5169
rect 1398 5164 1399 5168
rect 1403 5164 1404 5168
rect 1398 5163 1404 5164
rect 1606 5168 1612 5169
rect 1606 5164 1607 5168
rect 1611 5164 1612 5168
rect 1606 5163 1612 5164
rect 1814 5168 1820 5169
rect 1814 5164 1815 5168
rect 1819 5164 1820 5168
rect 1934 5165 1935 5169
rect 1939 5165 1940 5169
rect 1934 5164 1940 5165
rect 1974 5168 1980 5169
rect 2276 5168 2278 5229
rect 2476 5168 2478 5229
rect 2684 5168 2686 5229
rect 2892 5168 2894 5229
rect 3100 5168 3102 5229
rect 3308 5168 3310 5229
rect 3800 5169 3802 5229
rect 3840 5223 3842 5299
rect 4404 5223 4406 5300
rect 4588 5223 4590 5300
rect 4772 5223 4774 5300
rect 4956 5223 4958 5300
rect 5148 5223 5150 5300
rect 5662 5299 5668 5300
rect 5664 5223 5666 5299
rect 3839 5222 3843 5223
rect 3839 5217 3843 5218
rect 4403 5222 4407 5223
rect 4403 5217 4407 5218
rect 4435 5222 4439 5223
rect 4435 5217 4439 5218
rect 4587 5222 4591 5223
rect 4587 5217 4591 5218
rect 4595 5222 4599 5223
rect 4595 5217 4599 5218
rect 4755 5222 4759 5223
rect 4755 5217 4759 5218
rect 4771 5222 4775 5223
rect 4771 5217 4775 5218
rect 4915 5222 4919 5223
rect 4915 5217 4919 5218
rect 4955 5222 4959 5223
rect 4955 5217 4959 5218
rect 5067 5222 5071 5223
rect 5067 5217 5071 5218
rect 5147 5222 5151 5223
rect 5147 5217 5151 5218
rect 5219 5222 5223 5223
rect 5219 5217 5223 5218
rect 5379 5222 5383 5223
rect 5379 5217 5383 5218
rect 5515 5222 5519 5223
rect 5515 5217 5519 5218
rect 5663 5222 5667 5223
rect 5663 5217 5667 5218
rect 3798 5168 3804 5169
rect 1974 5164 1975 5168
rect 1979 5164 1980 5168
rect 1814 5163 1820 5164
rect 1974 5163 1980 5164
rect 2274 5167 2280 5168
rect 2274 5163 2275 5167
rect 2279 5163 2280 5167
rect 2274 5162 2280 5163
rect 2474 5167 2480 5168
rect 2474 5163 2475 5167
rect 2479 5163 2480 5167
rect 2474 5162 2480 5163
rect 2682 5167 2688 5168
rect 2682 5163 2683 5167
rect 2687 5163 2688 5167
rect 2682 5162 2688 5163
rect 2890 5167 2896 5168
rect 2890 5163 2891 5167
rect 2895 5163 2896 5167
rect 2890 5162 2896 5163
rect 3098 5167 3104 5168
rect 3098 5163 3099 5167
rect 3103 5163 3104 5167
rect 3098 5162 3104 5163
rect 3306 5167 3312 5168
rect 3306 5163 3307 5167
rect 3311 5163 3312 5167
rect 3798 5164 3799 5168
rect 3803 5164 3804 5168
rect 3798 5163 3804 5164
rect 3306 5162 3312 5163
rect 3840 5157 3842 5217
rect 3838 5156 3844 5157
rect 4436 5156 4438 5217
rect 4596 5156 4598 5217
rect 4756 5156 4758 5217
rect 4916 5156 4918 5217
rect 5068 5156 5070 5217
rect 5220 5156 5222 5217
rect 5380 5156 5382 5217
rect 5516 5156 5518 5217
rect 5664 5157 5666 5217
rect 5662 5156 5668 5157
rect 418 5153 424 5154
rect 110 5152 116 5153
rect 110 5148 111 5152
rect 115 5148 116 5152
rect 418 5149 419 5153
rect 423 5149 424 5153
rect 418 5148 424 5149
rect 594 5153 600 5154
rect 594 5149 595 5153
rect 599 5149 600 5153
rect 594 5148 600 5149
rect 778 5153 784 5154
rect 778 5149 779 5153
rect 783 5149 784 5153
rect 778 5148 784 5149
rect 970 5153 976 5154
rect 970 5149 971 5153
rect 975 5149 976 5153
rect 970 5148 976 5149
rect 1170 5153 1176 5154
rect 1170 5149 1171 5153
rect 1175 5149 1176 5153
rect 1170 5148 1176 5149
rect 1370 5153 1376 5154
rect 1370 5149 1371 5153
rect 1375 5149 1376 5153
rect 1370 5148 1376 5149
rect 1578 5153 1584 5154
rect 1578 5149 1579 5153
rect 1583 5149 1584 5153
rect 1578 5148 1584 5149
rect 1786 5153 1792 5154
rect 1786 5149 1787 5153
rect 1791 5149 1792 5153
rect 1786 5148 1792 5149
rect 1934 5152 1940 5153
rect 2302 5152 2308 5153
rect 1934 5148 1935 5152
rect 1939 5148 1940 5152
rect 110 5147 116 5148
rect 112 5079 114 5147
rect 420 5079 422 5148
rect 596 5079 598 5148
rect 780 5079 782 5148
rect 972 5079 974 5148
rect 1172 5079 1174 5148
rect 1372 5079 1374 5148
rect 1580 5079 1582 5148
rect 1788 5079 1790 5148
rect 1934 5147 1940 5148
rect 1974 5151 1980 5152
rect 1974 5147 1975 5151
rect 1979 5147 1980 5151
rect 2302 5148 2303 5152
rect 2307 5148 2308 5152
rect 2302 5147 2308 5148
rect 2502 5152 2508 5153
rect 2502 5148 2503 5152
rect 2507 5148 2508 5152
rect 2502 5147 2508 5148
rect 2710 5152 2716 5153
rect 2710 5148 2711 5152
rect 2715 5148 2716 5152
rect 2710 5147 2716 5148
rect 2918 5152 2924 5153
rect 2918 5148 2919 5152
rect 2923 5148 2924 5152
rect 2918 5147 2924 5148
rect 3126 5152 3132 5153
rect 3126 5148 3127 5152
rect 3131 5148 3132 5152
rect 3126 5147 3132 5148
rect 3334 5152 3340 5153
rect 3838 5152 3839 5156
rect 3843 5152 3844 5156
rect 3334 5148 3335 5152
rect 3339 5148 3340 5152
rect 3334 5147 3340 5148
rect 3798 5151 3804 5152
rect 3838 5151 3844 5152
rect 4434 5155 4440 5156
rect 4434 5151 4435 5155
rect 4439 5151 4440 5155
rect 3798 5147 3799 5151
rect 3803 5147 3804 5151
rect 4434 5150 4440 5151
rect 4594 5155 4600 5156
rect 4594 5151 4595 5155
rect 4599 5151 4600 5155
rect 4594 5150 4600 5151
rect 4754 5155 4760 5156
rect 4754 5151 4755 5155
rect 4759 5151 4760 5155
rect 4754 5150 4760 5151
rect 4914 5155 4920 5156
rect 4914 5151 4915 5155
rect 4919 5151 4920 5155
rect 4914 5150 4920 5151
rect 5066 5155 5072 5156
rect 5066 5151 5067 5155
rect 5071 5151 5072 5155
rect 5066 5150 5072 5151
rect 5218 5155 5224 5156
rect 5218 5151 5219 5155
rect 5223 5151 5224 5155
rect 5218 5150 5224 5151
rect 5378 5155 5384 5156
rect 5378 5151 5379 5155
rect 5383 5151 5384 5155
rect 5378 5150 5384 5151
rect 5514 5155 5520 5156
rect 5514 5151 5515 5155
rect 5519 5151 5520 5155
rect 5662 5152 5663 5156
rect 5667 5152 5668 5156
rect 5662 5151 5668 5152
rect 5514 5150 5520 5151
rect 1936 5079 1938 5147
rect 1974 5146 1980 5147
rect 1976 5107 1978 5146
rect 2304 5107 2306 5147
rect 2504 5107 2506 5147
rect 2712 5107 2714 5147
rect 2920 5107 2922 5147
rect 3128 5107 3130 5147
rect 3336 5107 3338 5147
rect 3798 5146 3804 5147
rect 3800 5107 3802 5146
rect 4462 5140 4468 5141
rect 3838 5139 3844 5140
rect 3838 5135 3839 5139
rect 3843 5135 3844 5139
rect 4462 5136 4463 5140
rect 4467 5136 4468 5140
rect 4462 5135 4468 5136
rect 4622 5140 4628 5141
rect 4622 5136 4623 5140
rect 4627 5136 4628 5140
rect 4622 5135 4628 5136
rect 4782 5140 4788 5141
rect 4782 5136 4783 5140
rect 4787 5136 4788 5140
rect 4782 5135 4788 5136
rect 4942 5140 4948 5141
rect 4942 5136 4943 5140
rect 4947 5136 4948 5140
rect 4942 5135 4948 5136
rect 5094 5140 5100 5141
rect 5094 5136 5095 5140
rect 5099 5136 5100 5140
rect 5094 5135 5100 5136
rect 5246 5140 5252 5141
rect 5246 5136 5247 5140
rect 5251 5136 5252 5140
rect 5246 5135 5252 5136
rect 5406 5140 5412 5141
rect 5406 5136 5407 5140
rect 5411 5136 5412 5140
rect 5406 5135 5412 5136
rect 5542 5140 5548 5141
rect 5542 5136 5543 5140
rect 5547 5136 5548 5140
rect 5542 5135 5548 5136
rect 5662 5139 5668 5140
rect 5662 5135 5663 5139
rect 5667 5135 5668 5139
rect 3838 5134 3844 5135
rect 1975 5106 1979 5107
rect 1975 5101 1979 5102
rect 2119 5106 2123 5107
rect 2119 5101 2123 5102
rect 2303 5106 2307 5107
rect 2303 5101 2307 5102
rect 2327 5106 2331 5107
rect 2327 5101 2331 5102
rect 2503 5106 2507 5107
rect 2503 5101 2507 5102
rect 2535 5106 2539 5107
rect 2535 5101 2539 5102
rect 2711 5106 2715 5107
rect 2711 5101 2715 5102
rect 2751 5106 2755 5107
rect 2751 5101 2755 5102
rect 2919 5106 2923 5107
rect 2919 5101 2923 5102
rect 2975 5106 2979 5107
rect 2975 5101 2979 5102
rect 3127 5106 3131 5107
rect 3127 5101 3131 5102
rect 3207 5106 3211 5107
rect 3207 5101 3211 5102
rect 3335 5106 3339 5107
rect 3335 5101 3339 5102
rect 3799 5106 3803 5107
rect 3840 5103 3842 5134
rect 4464 5103 4466 5135
rect 4624 5103 4626 5135
rect 4784 5103 4786 5135
rect 4944 5103 4946 5135
rect 5096 5103 5098 5135
rect 5248 5103 5250 5135
rect 5408 5103 5410 5135
rect 5544 5103 5546 5135
rect 5662 5134 5668 5135
rect 5664 5103 5666 5134
rect 3799 5101 3803 5102
rect 3839 5102 3843 5103
rect 111 5078 115 5079
rect 111 5073 115 5074
rect 155 5078 159 5079
rect 155 5073 159 5074
rect 379 5078 383 5079
rect 379 5073 383 5074
rect 419 5078 423 5079
rect 419 5073 423 5074
rect 595 5078 599 5079
rect 595 5073 599 5074
rect 627 5078 631 5079
rect 627 5073 631 5074
rect 779 5078 783 5079
rect 779 5073 783 5074
rect 899 5078 903 5079
rect 899 5073 903 5074
rect 971 5078 975 5079
rect 971 5073 975 5074
rect 1171 5078 1175 5079
rect 1171 5073 1175 5074
rect 1195 5078 1199 5079
rect 1195 5073 1199 5074
rect 1371 5078 1375 5079
rect 1371 5073 1375 5074
rect 1499 5078 1503 5079
rect 1499 5073 1503 5074
rect 1579 5078 1583 5079
rect 1579 5073 1583 5074
rect 1787 5078 1791 5079
rect 1787 5073 1791 5074
rect 1935 5078 1939 5079
rect 1976 5078 1978 5101
rect 1935 5073 1939 5074
rect 1974 5077 1980 5078
rect 2120 5077 2122 5101
rect 2328 5077 2330 5101
rect 2536 5077 2538 5101
rect 2752 5077 2754 5101
rect 2976 5077 2978 5101
rect 3208 5077 3210 5101
rect 3800 5078 3802 5101
rect 3839 5097 3843 5098
rect 3887 5102 3891 5103
rect 3887 5097 3891 5098
rect 4087 5102 4091 5103
rect 4087 5097 4091 5098
rect 4327 5102 4331 5103
rect 4327 5097 4331 5098
rect 4463 5102 4467 5103
rect 4463 5097 4467 5098
rect 4567 5102 4571 5103
rect 4567 5097 4571 5098
rect 4623 5102 4627 5103
rect 4623 5097 4627 5098
rect 4783 5102 4787 5103
rect 4783 5097 4787 5098
rect 4815 5102 4819 5103
rect 4815 5097 4819 5098
rect 4943 5102 4947 5103
rect 4943 5097 4947 5098
rect 5063 5102 5067 5103
rect 5063 5097 5067 5098
rect 5095 5102 5099 5103
rect 5095 5097 5099 5098
rect 5247 5102 5251 5103
rect 5247 5097 5251 5098
rect 5311 5102 5315 5103
rect 5311 5097 5315 5098
rect 5407 5102 5411 5103
rect 5407 5097 5411 5098
rect 5543 5102 5547 5103
rect 5543 5097 5547 5098
rect 5663 5102 5667 5103
rect 5663 5097 5667 5098
rect 3798 5077 3804 5078
rect 1974 5073 1975 5077
rect 1979 5073 1980 5077
rect 112 5013 114 5073
rect 110 5012 116 5013
rect 156 5012 158 5073
rect 380 5012 382 5073
rect 628 5012 630 5073
rect 900 5012 902 5073
rect 1196 5012 1198 5073
rect 1500 5012 1502 5073
rect 1788 5012 1790 5073
rect 1936 5013 1938 5073
rect 1974 5072 1980 5073
rect 2118 5076 2124 5077
rect 2118 5072 2119 5076
rect 2123 5072 2124 5076
rect 2118 5071 2124 5072
rect 2326 5076 2332 5077
rect 2326 5072 2327 5076
rect 2331 5072 2332 5076
rect 2326 5071 2332 5072
rect 2534 5076 2540 5077
rect 2534 5072 2535 5076
rect 2539 5072 2540 5076
rect 2534 5071 2540 5072
rect 2750 5076 2756 5077
rect 2750 5072 2751 5076
rect 2755 5072 2756 5076
rect 2750 5071 2756 5072
rect 2974 5076 2980 5077
rect 2974 5072 2975 5076
rect 2979 5072 2980 5076
rect 2974 5071 2980 5072
rect 3206 5076 3212 5077
rect 3206 5072 3207 5076
rect 3211 5072 3212 5076
rect 3798 5073 3799 5077
rect 3803 5073 3804 5077
rect 3840 5074 3842 5097
rect 3798 5072 3804 5073
rect 3838 5073 3844 5074
rect 3888 5073 3890 5097
rect 4088 5073 4090 5097
rect 4328 5073 4330 5097
rect 4568 5073 4570 5097
rect 4816 5073 4818 5097
rect 5064 5073 5066 5097
rect 5312 5073 5314 5097
rect 5544 5073 5546 5097
rect 5664 5074 5666 5097
rect 5662 5073 5668 5074
rect 3206 5071 3212 5072
rect 3838 5069 3839 5073
rect 3843 5069 3844 5073
rect 3838 5068 3844 5069
rect 3886 5072 3892 5073
rect 3886 5068 3887 5072
rect 3891 5068 3892 5072
rect 3886 5067 3892 5068
rect 4086 5072 4092 5073
rect 4086 5068 4087 5072
rect 4091 5068 4092 5072
rect 4086 5067 4092 5068
rect 4326 5072 4332 5073
rect 4326 5068 4327 5072
rect 4331 5068 4332 5072
rect 4326 5067 4332 5068
rect 4566 5072 4572 5073
rect 4566 5068 4567 5072
rect 4571 5068 4572 5072
rect 4566 5067 4572 5068
rect 4814 5072 4820 5073
rect 4814 5068 4815 5072
rect 4819 5068 4820 5072
rect 4814 5067 4820 5068
rect 5062 5072 5068 5073
rect 5062 5068 5063 5072
rect 5067 5068 5068 5072
rect 5062 5067 5068 5068
rect 5310 5072 5316 5073
rect 5310 5068 5311 5072
rect 5315 5068 5316 5072
rect 5310 5067 5316 5068
rect 5542 5072 5548 5073
rect 5542 5068 5543 5072
rect 5547 5068 5548 5072
rect 5662 5069 5663 5073
rect 5667 5069 5668 5073
rect 5662 5068 5668 5069
rect 5542 5067 5548 5068
rect 2090 5061 2096 5062
rect 1974 5060 1980 5061
rect 1974 5056 1975 5060
rect 1979 5056 1980 5060
rect 2090 5057 2091 5061
rect 2095 5057 2096 5061
rect 2090 5056 2096 5057
rect 2298 5061 2304 5062
rect 2298 5057 2299 5061
rect 2303 5057 2304 5061
rect 2298 5056 2304 5057
rect 2506 5061 2512 5062
rect 2506 5057 2507 5061
rect 2511 5057 2512 5061
rect 2506 5056 2512 5057
rect 2722 5061 2728 5062
rect 2722 5057 2723 5061
rect 2727 5057 2728 5061
rect 2722 5056 2728 5057
rect 2946 5061 2952 5062
rect 2946 5057 2947 5061
rect 2951 5057 2952 5061
rect 2946 5056 2952 5057
rect 3178 5061 3184 5062
rect 3178 5057 3179 5061
rect 3183 5057 3184 5061
rect 3178 5056 3184 5057
rect 3798 5060 3804 5061
rect 3798 5056 3799 5060
rect 3803 5056 3804 5060
rect 3858 5057 3864 5058
rect 1974 5055 1980 5056
rect 1934 5012 1940 5013
rect 110 5008 111 5012
rect 115 5008 116 5012
rect 110 5007 116 5008
rect 154 5011 160 5012
rect 154 5007 155 5011
rect 159 5007 160 5011
rect 154 5006 160 5007
rect 378 5011 384 5012
rect 378 5007 379 5011
rect 383 5007 384 5011
rect 378 5006 384 5007
rect 626 5011 632 5012
rect 626 5007 627 5011
rect 631 5007 632 5011
rect 626 5006 632 5007
rect 898 5011 904 5012
rect 898 5007 899 5011
rect 903 5007 904 5011
rect 898 5006 904 5007
rect 1194 5011 1200 5012
rect 1194 5007 1195 5011
rect 1199 5007 1200 5011
rect 1194 5006 1200 5007
rect 1498 5011 1504 5012
rect 1498 5007 1499 5011
rect 1503 5007 1504 5011
rect 1498 5006 1504 5007
rect 1786 5011 1792 5012
rect 1786 5007 1787 5011
rect 1791 5007 1792 5011
rect 1934 5008 1935 5012
rect 1939 5008 1940 5012
rect 1934 5007 1940 5008
rect 1786 5006 1792 5007
rect 182 4996 188 4997
rect 110 4995 116 4996
rect 110 4991 111 4995
rect 115 4991 116 4995
rect 182 4992 183 4996
rect 187 4992 188 4996
rect 182 4991 188 4992
rect 406 4996 412 4997
rect 406 4992 407 4996
rect 411 4992 412 4996
rect 406 4991 412 4992
rect 654 4996 660 4997
rect 654 4992 655 4996
rect 659 4992 660 4996
rect 654 4991 660 4992
rect 926 4996 932 4997
rect 926 4992 927 4996
rect 931 4992 932 4996
rect 926 4991 932 4992
rect 1222 4996 1228 4997
rect 1222 4992 1223 4996
rect 1227 4992 1228 4996
rect 1222 4991 1228 4992
rect 1526 4996 1532 4997
rect 1526 4992 1527 4996
rect 1531 4992 1532 4996
rect 1526 4991 1532 4992
rect 1814 4996 1820 4997
rect 1814 4992 1815 4996
rect 1819 4992 1820 4996
rect 1814 4991 1820 4992
rect 1934 4995 1940 4996
rect 1934 4991 1935 4995
rect 1939 4991 1940 4995
rect 110 4990 116 4991
rect 112 4939 114 4990
rect 184 4939 186 4991
rect 408 4939 410 4991
rect 656 4939 658 4991
rect 928 4939 930 4991
rect 1224 4939 1226 4991
rect 1528 4939 1530 4991
rect 1816 4939 1818 4991
rect 1934 4990 1940 4991
rect 1936 4939 1938 4990
rect 1976 4987 1978 5055
rect 2092 4987 2094 5056
rect 2300 4987 2302 5056
rect 2508 4987 2510 5056
rect 2724 4987 2726 5056
rect 2948 4987 2950 5056
rect 3180 4987 3182 5056
rect 3798 5055 3804 5056
rect 3838 5056 3844 5057
rect 3800 4987 3802 5055
rect 3838 5052 3839 5056
rect 3843 5052 3844 5056
rect 3858 5053 3859 5057
rect 3863 5053 3864 5057
rect 3858 5052 3864 5053
rect 4058 5057 4064 5058
rect 4058 5053 4059 5057
rect 4063 5053 4064 5057
rect 4058 5052 4064 5053
rect 4298 5057 4304 5058
rect 4298 5053 4299 5057
rect 4303 5053 4304 5057
rect 4298 5052 4304 5053
rect 4538 5057 4544 5058
rect 4538 5053 4539 5057
rect 4543 5053 4544 5057
rect 4538 5052 4544 5053
rect 4786 5057 4792 5058
rect 4786 5053 4787 5057
rect 4791 5053 4792 5057
rect 4786 5052 4792 5053
rect 5034 5057 5040 5058
rect 5034 5053 5035 5057
rect 5039 5053 5040 5057
rect 5034 5052 5040 5053
rect 5282 5057 5288 5058
rect 5282 5053 5283 5057
rect 5287 5053 5288 5057
rect 5282 5052 5288 5053
rect 5514 5057 5520 5058
rect 5514 5053 5515 5057
rect 5519 5053 5520 5057
rect 5514 5052 5520 5053
rect 5662 5056 5668 5057
rect 5662 5052 5663 5056
rect 5667 5052 5668 5056
rect 3838 5051 3844 5052
rect 3840 4991 3842 5051
rect 3860 4991 3862 5052
rect 4060 4991 4062 5052
rect 4300 4991 4302 5052
rect 4540 4991 4542 5052
rect 4788 4991 4790 5052
rect 5036 4991 5038 5052
rect 5284 4991 5286 5052
rect 5516 4991 5518 5052
rect 5662 5051 5668 5052
rect 5664 4991 5666 5051
rect 3839 4990 3843 4991
rect 1975 4986 1979 4987
rect 1975 4981 1979 4982
rect 1995 4986 1999 4987
rect 1995 4981 1999 4982
rect 2091 4986 2095 4987
rect 2091 4981 2095 4982
rect 2131 4986 2135 4987
rect 2131 4981 2135 4982
rect 2267 4986 2271 4987
rect 2267 4981 2271 4982
rect 2299 4986 2303 4987
rect 2299 4981 2303 4982
rect 2419 4986 2423 4987
rect 2419 4981 2423 4982
rect 2507 4986 2511 4987
rect 2507 4981 2511 4982
rect 2619 4986 2623 4987
rect 2619 4981 2623 4982
rect 2723 4986 2727 4987
rect 2723 4981 2727 4982
rect 2859 4986 2863 4987
rect 2859 4981 2863 4982
rect 2947 4986 2951 4987
rect 2947 4981 2951 4982
rect 3123 4986 3127 4987
rect 3123 4981 3127 4982
rect 3179 4986 3183 4987
rect 3179 4981 3183 4982
rect 3395 4986 3399 4987
rect 3395 4981 3399 4982
rect 3651 4986 3655 4987
rect 3651 4981 3655 4982
rect 3799 4986 3803 4987
rect 3839 4985 3843 4986
rect 3859 4990 3863 4991
rect 3859 4985 3863 4986
rect 3995 4990 3999 4991
rect 3995 4985 3999 4986
rect 4059 4990 4063 4991
rect 4059 4985 4063 4986
rect 4131 4990 4135 4991
rect 4131 4985 4135 4986
rect 4267 4990 4271 4991
rect 4267 4985 4271 4986
rect 4299 4990 4303 4991
rect 4299 4985 4303 4986
rect 4403 4990 4407 4991
rect 4403 4985 4407 4986
rect 4539 4990 4543 4991
rect 4539 4985 4543 4986
rect 4675 4990 4679 4991
rect 4675 4985 4679 4986
rect 4787 4990 4791 4991
rect 4787 4985 4791 4986
rect 4811 4990 4815 4991
rect 4811 4985 4815 4986
rect 4947 4990 4951 4991
rect 4947 4985 4951 4986
rect 5035 4990 5039 4991
rect 5035 4985 5039 4986
rect 5083 4990 5087 4991
rect 5083 4985 5087 4986
rect 5227 4990 5231 4991
rect 5227 4985 5231 4986
rect 5283 4990 5287 4991
rect 5283 4985 5287 4986
rect 5379 4990 5383 4991
rect 5379 4985 5383 4986
rect 5515 4990 5519 4991
rect 5515 4985 5519 4986
rect 5663 4990 5667 4991
rect 5663 4985 5667 4986
rect 3799 4981 3803 4982
rect 111 4938 115 4939
rect 111 4933 115 4934
rect 159 4938 163 4939
rect 159 4933 163 4934
rect 183 4938 187 4939
rect 183 4933 187 4934
rect 295 4938 299 4939
rect 295 4933 299 4934
rect 407 4938 411 4939
rect 407 4933 411 4934
rect 431 4938 435 4939
rect 431 4933 435 4934
rect 567 4938 571 4939
rect 567 4933 571 4934
rect 655 4938 659 4939
rect 655 4933 659 4934
rect 703 4938 707 4939
rect 703 4933 707 4934
rect 927 4938 931 4939
rect 927 4933 931 4934
rect 1223 4938 1227 4939
rect 1223 4933 1227 4934
rect 1527 4938 1531 4939
rect 1527 4933 1531 4934
rect 1815 4938 1819 4939
rect 1815 4933 1819 4934
rect 1935 4938 1939 4939
rect 1935 4933 1939 4934
rect 112 4910 114 4933
rect 110 4909 116 4910
rect 160 4909 162 4933
rect 296 4909 298 4933
rect 432 4909 434 4933
rect 568 4909 570 4933
rect 704 4909 706 4933
rect 1936 4910 1938 4933
rect 1976 4921 1978 4981
rect 1974 4920 1980 4921
rect 1996 4920 1998 4981
rect 2132 4920 2134 4981
rect 2268 4920 2270 4981
rect 2420 4920 2422 4981
rect 2620 4920 2622 4981
rect 2860 4920 2862 4981
rect 3124 4920 3126 4981
rect 3396 4920 3398 4981
rect 3652 4920 3654 4981
rect 3800 4921 3802 4981
rect 3840 4925 3842 4985
rect 3838 4924 3844 4925
rect 3860 4924 3862 4985
rect 3996 4924 3998 4985
rect 4132 4924 4134 4985
rect 4268 4924 4270 4985
rect 4404 4924 4406 4985
rect 4540 4924 4542 4985
rect 4676 4924 4678 4985
rect 4812 4924 4814 4985
rect 4948 4924 4950 4985
rect 5084 4924 5086 4985
rect 5228 4924 5230 4985
rect 5380 4924 5382 4985
rect 5516 4924 5518 4985
rect 5664 4925 5666 4985
rect 5662 4924 5668 4925
rect 3798 4920 3804 4921
rect 1974 4916 1975 4920
rect 1979 4916 1980 4920
rect 1974 4915 1980 4916
rect 1994 4919 2000 4920
rect 1994 4915 1995 4919
rect 1999 4915 2000 4919
rect 1994 4914 2000 4915
rect 2130 4919 2136 4920
rect 2130 4915 2131 4919
rect 2135 4915 2136 4919
rect 2130 4914 2136 4915
rect 2266 4919 2272 4920
rect 2266 4915 2267 4919
rect 2271 4915 2272 4919
rect 2266 4914 2272 4915
rect 2418 4919 2424 4920
rect 2418 4915 2419 4919
rect 2423 4915 2424 4919
rect 2418 4914 2424 4915
rect 2618 4919 2624 4920
rect 2618 4915 2619 4919
rect 2623 4915 2624 4919
rect 2618 4914 2624 4915
rect 2858 4919 2864 4920
rect 2858 4915 2859 4919
rect 2863 4915 2864 4919
rect 2858 4914 2864 4915
rect 3122 4919 3128 4920
rect 3122 4915 3123 4919
rect 3127 4915 3128 4919
rect 3122 4914 3128 4915
rect 3394 4919 3400 4920
rect 3394 4915 3395 4919
rect 3399 4915 3400 4919
rect 3394 4914 3400 4915
rect 3650 4919 3656 4920
rect 3650 4915 3651 4919
rect 3655 4915 3656 4919
rect 3798 4916 3799 4920
rect 3803 4916 3804 4920
rect 3838 4920 3839 4924
rect 3843 4920 3844 4924
rect 3838 4919 3844 4920
rect 3858 4923 3864 4924
rect 3858 4919 3859 4923
rect 3863 4919 3864 4923
rect 3858 4918 3864 4919
rect 3994 4923 4000 4924
rect 3994 4919 3995 4923
rect 3999 4919 4000 4923
rect 3994 4918 4000 4919
rect 4130 4923 4136 4924
rect 4130 4919 4131 4923
rect 4135 4919 4136 4923
rect 4130 4918 4136 4919
rect 4266 4923 4272 4924
rect 4266 4919 4267 4923
rect 4271 4919 4272 4923
rect 4266 4918 4272 4919
rect 4402 4923 4408 4924
rect 4402 4919 4403 4923
rect 4407 4919 4408 4923
rect 4402 4918 4408 4919
rect 4538 4923 4544 4924
rect 4538 4919 4539 4923
rect 4543 4919 4544 4923
rect 4538 4918 4544 4919
rect 4674 4923 4680 4924
rect 4674 4919 4675 4923
rect 4679 4919 4680 4923
rect 4674 4918 4680 4919
rect 4810 4923 4816 4924
rect 4810 4919 4811 4923
rect 4815 4919 4816 4923
rect 4810 4918 4816 4919
rect 4946 4923 4952 4924
rect 4946 4919 4947 4923
rect 4951 4919 4952 4923
rect 4946 4918 4952 4919
rect 5082 4923 5088 4924
rect 5082 4919 5083 4923
rect 5087 4919 5088 4923
rect 5082 4918 5088 4919
rect 5226 4923 5232 4924
rect 5226 4919 5227 4923
rect 5231 4919 5232 4923
rect 5226 4918 5232 4919
rect 5378 4923 5384 4924
rect 5378 4919 5379 4923
rect 5383 4919 5384 4923
rect 5378 4918 5384 4919
rect 5514 4923 5520 4924
rect 5514 4919 5515 4923
rect 5519 4919 5520 4923
rect 5662 4920 5663 4924
rect 5667 4920 5668 4924
rect 5662 4919 5668 4920
rect 5514 4918 5520 4919
rect 3798 4915 3804 4916
rect 3650 4914 3656 4915
rect 1934 4909 1940 4910
rect 110 4905 111 4909
rect 115 4905 116 4909
rect 110 4904 116 4905
rect 158 4908 164 4909
rect 158 4904 159 4908
rect 163 4904 164 4908
rect 158 4903 164 4904
rect 294 4908 300 4909
rect 294 4904 295 4908
rect 299 4904 300 4908
rect 294 4903 300 4904
rect 430 4908 436 4909
rect 430 4904 431 4908
rect 435 4904 436 4908
rect 430 4903 436 4904
rect 566 4908 572 4909
rect 566 4904 567 4908
rect 571 4904 572 4908
rect 566 4903 572 4904
rect 702 4908 708 4909
rect 702 4904 703 4908
rect 707 4904 708 4908
rect 1934 4905 1935 4909
rect 1939 4905 1940 4909
rect 3886 4908 3892 4909
rect 3838 4907 3844 4908
rect 1934 4904 1940 4905
rect 2022 4904 2028 4905
rect 702 4903 708 4904
rect 1974 4903 1980 4904
rect 1974 4899 1975 4903
rect 1979 4899 1980 4903
rect 2022 4900 2023 4904
rect 2027 4900 2028 4904
rect 2022 4899 2028 4900
rect 2158 4904 2164 4905
rect 2158 4900 2159 4904
rect 2163 4900 2164 4904
rect 2158 4899 2164 4900
rect 2294 4904 2300 4905
rect 2294 4900 2295 4904
rect 2299 4900 2300 4904
rect 2294 4899 2300 4900
rect 2446 4904 2452 4905
rect 2446 4900 2447 4904
rect 2451 4900 2452 4904
rect 2446 4899 2452 4900
rect 2646 4904 2652 4905
rect 2646 4900 2647 4904
rect 2651 4900 2652 4904
rect 2646 4899 2652 4900
rect 2886 4904 2892 4905
rect 2886 4900 2887 4904
rect 2891 4900 2892 4904
rect 2886 4899 2892 4900
rect 3150 4904 3156 4905
rect 3150 4900 3151 4904
rect 3155 4900 3156 4904
rect 3150 4899 3156 4900
rect 3422 4904 3428 4905
rect 3422 4900 3423 4904
rect 3427 4900 3428 4904
rect 3422 4899 3428 4900
rect 3678 4904 3684 4905
rect 3678 4900 3679 4904
rect 3683 4900 3684 4904
rect 3678 4899 3684 4900
rect 3798 4903 3804 4904
rect 3798 4899 3799 4903
rect 3803 4899 3804 4903
rect 3838 4903 3839 4907
rect 3843 4903 3844 4907
rect 3886 4904 3887 4908
rect 3891 4904 3892 4908
rect 3886 4903 3892 4904
rect 4022 4908 4028 4909
rect 4022 4904 4023 4908
rect 4027 4904 4028 4908
rect 4022 4903 4028 4904
rect 4158 4908 4164 4909
rect 4158 4904 4159 4908
rect 4163 4904 4164 4908
rect 4158 4903 4164 4904
rect 4294 4908 4300 4909
rect 4294 4904 4295 4908
rect 4299 4904 4300 4908
rect 4294 4903 4300 4904
rect 4430 4908 4436 4909
rect 4430 4904 4431 4908
rect 4435 4904 4436 4908
rect 4430 4903 4436 4904
rect 4566 4908 4572 4909
rect 4566 4904 4567 4908
rect 4571 4904 4572 4908
rect 4566 4903 4572 4904
rect 4702 4908 4708 4909
rect 4702 4904 4703 4908
rect 4707 4904 4708 4908
rect 4702 4903 4708 4904
rect 4838 4908 4844 4909
rect 4838 4904 4839 4908
rect 4843 4904 4844 4908
rect 4838 4903 4844 4904
rect 4974 4908 4980 4909
rect 4974 4904 4975 4908
rect 4979 4904 4980 4908
rect 4974 4903 4980 4904
rect 5110 4908 5116 4909
rect 5110 4904 5111 4908
rect 5115 4904 5116 4908
rect 5110 4903 5116 4904
rect 5254 4908 5260 4909
rect 5254 4904 5255 4908
rect 5259 4904 5260 4908
rect 5254 4903 5260 4904
rect 5406 4908 5412 4909
rect 5406 4904 5407 4908
rect 5411 4904 5412 4908
rect 5406 4903 5412 4904
rect 5542 4908 5548 4909
rect 5542 4904 5543 4908
rect 5547 4904 5548 4908
rect 5542 4903 5548 4904
rect 5662 4907 5668 4908
rect 5662 4903 5663 4907
rect 5667 4903 5668 4907
rect 3838 4902 3844 4903
rect 1974 4898 1980 4899
rect 130 4893 136 4894
rect 110 4892 116 4893
rect 110 4888 111 4892
rect 115 4888 116 4892
rect 130 4889 131 4893
rect 135 4889 136 4893
rect 130 4888 136 4889
rect 266 4893 272 4894
rect 266 4889 267 4893
rect 271 4889 272 4893
rect 266 4888 272 4889
rect 402 4893 408 4894
rect 402 4889 403 4893
rect 407 4889 408 4893
rect 402 4888 408 4889
rect 538 4893 544 4894
rect 538 4889 539 4893
rect 543 4889 544 4893
rect 538 4888 544 4889
rect 674 4893 680 4894
rect 674 4889 675 4893
rect 679 4889 680 4893
rect 674 4888 680 4889
rect 1934 4892 1940 4893
rect 1934 4888 1935 4892
rect 1939 4888 1940 4892
rect 110 4887 116 4888
rect 112 4815 114 4887
rect 132 4815 134 4888
rect 268 4815 270 4888
rect 404 4815 406 4888
rect 540 4815 542 4888
rect 676 4815 678 4888
rect 1934 4887 1940 4888
rect 1936 4815 1938 4887
rect 1976 4867 1978 4898
rect 2024 4867 2026 4899
rect 2160 4867 2162 4899
rect 2296 4867 2298 4899
rect 2448 4867 2450 4899
rect 2648 4867 2650 4899
rect 2888 4867 2890 4899
rect 3152 4867 3154 4899
rect 3424 4867 3426 4899
rect 3680 4867 3682 4899
rect 3798 4898 3804 4899
rect 3800 4867 3802 4898
rect 1975 4866 1979 4867
rect 1975 4861 1979 4862
rect 2023 4866 2027 4867
rect 2023 4861 2027 4862
rect 2159 4866 2163 4867
rect 2159 4861 2163 4862
rect 2295 4866 2299 4867
rect 2295 4861 2299 4862
rect 2327 4866 2331 4867
rect 2327 4861 2331 4862
rect 2447 4866 2451 4867
rect 2447 4861 2451 4862
rect 2559 4866 2563 4867
rect 2559 4861 2563 4862
rect 2647 4866 2651 4867
rect 2647 4861 2651 4862
rect 2823 4866 2827 4867
rect 2823 4861 2827 4862
rect 2887 4866 2891 4867
rect 2887 4861 2891 4862
rect 3103 4866 3107 4867
rect 3103 4861 3107 4862
rect 3151 4866 3155 4867
rect 3151 4861 3155 4862
rect 3399 4866 3403 4867
rect 3399 4861 3403 4862
rect 3423 4866 3427 4867
rect 3423 4861 3427 4862
rect 3679 4866 3683 4867
rect 3679 4861 3683 4862
rect 3799 4866 3803 4867
rect 3799 4861 3803 4862
rect 1976 4838 1978 4861
rect 1974 4837 1980 4838
rect 2328 4837 2330 4861
rect 2560 4837 2562 4861
rect 2824 4837 2826 4861
rect 3104 4837 3106 4861
rect 3400 4837 3402 4861
rect 3680 4837 3682 4861
rect 3800 4838 3802 4861
rect 3798 4837 3804 4838
rect 1974 4833 1975 4837
rect 1979 4833 1980 4837
rect 1974 4832 1980 4833
rect 2326 4836 2332 4837
rect 2326 4832 2327 4836
rect 2331 4832 2332 4836
rect 2326 4831 2332 4832
rect 2558 4836 2564 4837
rect 2558 4832 2559 4836
rect 2563 4832 2564 4836
rect 2558 4831 2564 4832
rect 2822 4836 2828 4837
rect 2822 4832 2823 4836
rect 2827 4832 2828 4836
rect 2822 4831 2828 4832
rect 3102 4836 3108 4837
rect 3102 4832 3103 4836
rect 3107 4832 3108 4836
rect 3102 4831 3108 4832
rect 3398 4836 3404 4837
rect 3398 4832 3399 4836
rect 3403 4832 3404 4836
rect 3398 4831 3404 4832
rect 3678 4836 3684 4837
rect 3678 4832 3679 4836
rect 3683 4832 3684 4836
rect 3798 4833 3799 4837
rect 3803 4833 3804 4837
rect 3798 4832 3804 4833
rect 3678 4831 3684 4832
rect 2298 4821 2304 4822
rect 1974 4820 1980 4821
rect 1974 4816 1975 4820
rect 1979 4816 1980 4820
rect 2298 4817 2299 4821
rect 2303 4817 2304 4821
rect 2298 4816 2304 4817
rect 2530 4821 2536 4822
rect 2530 4817 2531 4821
rect 2535 4817 2536 4821
rect 2530 4816 2536 4817
rect 2794 4821 2800 4822
rect 2794 4817 2795 4821
rect 2799 4817 2800 4821
rect 2794 4816 2800 4817
rect 3074 4821 3080 4822
rect 3074 4817 3075 4821
rect 3079 4817 3080 4821
rect 3074 4816 3080 4817
rect 3370 4821 3376 4822
rect 3370 4817 3371 4821
rect 3375 4817 3376 4821
rect 3370 4816 3376 4817
rect 3650 4821 3656 4822
rect 3650 4817 3651 4821
rect 3655 4817 3656 4821
rect 3650 4816 3656 4817
rect 3798 4820 3804 4821
rect 3798 4816 3799 4820
rect 3803 4816 3804 4820
rect 1974 4815 1980 4816
rect 111 4814 115 4815
rect 111 4809 115 4810
rect 131 4814 135 4815
rect 131 4809 135 4810
rect 267 4814 271 4815
rect 267 4809 271 4810
rect 403 4814 407 4815
rect 403 4809 407 4810
rect 539 4814 543 4815
rect 539 4809 543 4810
rect 675 4814 679 4815
rect 675 4809 679 4810
rect 1935 4814 1939 4815
rect 1935 4809 1939 4810
rect 112 4749 114 4809
rect 110 4748 116 4749
rect 132 4748 134 4809
rect 268 4748 270 4809
rect 404 4748 406 4809
rect 540 4748 542 4809
rect 676 4748 678 4809
rect 1936 4749 1938 4809
rect 1934 4748 1940 4749
rect 110 4744 111 4748
rect 115 4744 116 4748
rect 110 4743 116 4744
rect 130 4747 136 4748
rect 130 4743 131 4747
rect 135 4743 136 4747
rect 130 4742 136 4743
rect 266 4747 272 4748
rect 266 4743 267 4747
rect 271 4743 272 4747
rect 266 4742 272 4743
rect 402 4747 408 4748
rect 402 4743 403 4747
rect 407 4743 408 4747
rect 402 4742 408 4743
rect 538 4747 544 4748
rect 538 4743 539 4747
rect 543 4743 544 4747
rect 538 4742 544 4743
rect 674 4747 680 4748
rect 674 4743 675 4747
rect 679 4743 680 4747
rect 1934 4744 1935 4748
rect 1939 4744 1940 4748
rect 1934 4743 1940 4744
rect 1976 4743 1978 4815
rect 2300 4743 2302 4816
rect 2532 4743 2534 4816
rect 2796 4743 2798 4816
rect 3076 4743 3078 4816
rect 3372 4743 3374 4816
rect 3652 4743 3654 4816
rect 3798 4815 3804 4816
rect 3800 4743 3802 4815
rect 3840 4803 3842 4902
rect 3888 4803 3890 4903
rect 4024 4803 4026 4903
rect 4160 4803 4162 4903
rect 4296 4803 4298 4903
rect 4432 4803 4434 4903
rect 4568 4803 4570 4903
rect 4704 4803 4706 4903
rect 4840 4803 4842 4903
rect 4976 4803 4978 4903
rect 5112 4803 5114 4903
rect 5256 4803 5258 4903
rect 5408 4803 5410 4903
rect 5544 4803 5546 4903
rect 5662 4902 5668 4903
rect 5664 4803 5666 4902
rect 3839 4802 3843 4803
rect 3839 4797 3843 4798
rect 3887 4802 3891 4803
rect 3887 4797 3891 4798
rect 4023 4802 4027 4803
rect 4023 4797 4027 4798
rect 4071 4802 4075 4803
rect 4071 4797 4075 4798
rect 4159 4802 4163 4803
rect 4159 4797 4163 4798
rect 4295 4802 4299 4803
rect 4295 4797 4299 4798
rect 4431 4802 4435 4803
rect 4431 4797 4435 4798
rect 4535 4802 4539 4803
rect 4535 4797 4539 4798
rect 4567 4802 4571 4803
rect 4567 4797 4571 4798
rect 4703 4802 4707 4803
rect 4703 4797 4707 4798
rect 4783 4802 4787 4803
rect 4783 4797 4787 4798
rect 4839 4802 4843 4803
rect 4839 4797 4843 4798
rect 4975 4802 4979 4803
rect 4975 4797 4979 4798
rect 5039 4802 5043 4803
rect 5039 4797 5043 4798
rect 5111 4802 5115 4803
rect 5111 4797 5115 4798
rect 5255 4802 5259 4803
rect 5255 4797 5259 4798
rect 5303 4802 5307 4803
rect 5303 4797 5307 4798
rect 5407 4802 5411 4803
rect 5407 4797 5411 4798
rect 5543 4802 5547 4803
rect 5543 4797 5547 4798
rect 5663 4802 5667 4803
rect 5663 4797 5667 4798
rect 3840 4774 3842 4797
rect 3838 4773 3844 4774
rect 3888 4773 3890 4797
rect 4072 4773 4074 4797
rect 4296 4773 4298 4797
rect 4536 4773 4538 4797
rect 4784 4773 4786 4797
rect 5040 4773 5042 4797
rect 5304 4773 5306 4797
rect 5544 4773 5546 4797
rect 5664 4774 5666 4797
rect 5662 4773 5668 4774
rect 3838 4769 3839 4773
rect 3843 4769 3844 4773
rect 3838 4768 3844 4769
rect 3886 4772 3892 4773
rect 3886 4768 3887 4772
rect 3891 4768 3892 4772
rect 3886 4767 3892 4768
rect 4070 4772 4076 4773
rect 4070 4768 4071 4772
rect 4075 4768 4076 4772
rect 4070 4767 4076 4768
rect 4294 4772 4300 4773
rect 4294 4768 4295 4772
rect 4299 4768 4300 4772
rect 4294 4767 4300 4768
rect 4534 4772 4540 4773
rect 4534 4768 4535 4772
rect 4539 4768 4540 4772
rect 4534 4767 4540 4768
rect 4782 4772 4788 4773
rect 4782 4768 4783 4772
rect 4787 4768 4788 4772
rect 4782 4767 4788 4768
rect 5038 4772 5044 4773
rect 5038 4768 5039 4772
rect 5043 4768 5044 4772
rect 5038 4767 5044 4768
rect 5302 4772 5308 4773
rect 5302 4768 5303 4772
rect 5307 4768 5308 4772
rect 5302 4767 5308 4768
rect 5542 4772 5548 4773
rect 5542 4768 5543 4772
rect 5547 4768 5548 4772
rect 5662 4769 5663 4773
rect 5667 4769 5668 4773
rect 5662 4768 5668 4769
rect 5542 4767 5548 4768
rect 3858 4757 3864 4758
rect 3838 4756 3844 4757
rect 3838 4752 3839 4756
rect 3843 4752 3844 4756
rect 3858 4753 3859 4757
rect 3863 4753 3864 4757
rect 3858 4752 3864 4753
rect 4042 4757 4048 4758
rect 4042 4753 4043 4757
rect 4047 4753 4048 4757
rect 4042 4752 4048 4753
rect 4266 4757 4272 4758
rect 4266 4753 4267 4757
rect 4271 4753 4272 4757
rect 4266 4752 4272 4753
rect 4506 4757 4512 4758
rect 4506 4753 4507 4757
rect 4511 4753 4512 4757
rect 4506 4752 4512 4753
rect 4754 4757 4760 4758
rect 4754 4753 4755 4757
rect 4759 4753 4760 4757
rect 4754 4752 4760 4753
rect 5010 4757 5016 4758
rect 5010 4753 5011 4757
rect 5015 4753 5016 4757
rect 5010 4752 5016 4753
rect 5274 4757 5280 4758
rect 5274 4753 5275 4757
rect 5279 4753 5280 4757
rect 5274 4752 5280 4753
rect 5514 4757 5520 4758
rect 5514 4753 5515 4757
rect 5519 4753 5520 4757
rect 5514 4752 5520 4753
rect 5662 4756 5668 4757
rect 5662 4752 5663 4756
rect 5667 4752 5668 4756
rect 3838 4751 3844 4752
rect 674 4742 680 4743
rect 1975 4742 1979 4743
rect 1975 4737 1979 4738
rect 2019 4742 2023 4743
rect 2019 4737 2023 4738
rect 2195 4742 2199 4743
rect 2195 4737 2199 4738
rect 2299 4742 2303 4743
rect 2299 4737 2303 4738
rect 2371 4742 2375 4743
rect 2371 4737 2375 4738
rect 2531 4742 2535 4743
rect 2531 4737 2535 4738
rect 2547 4742 2551 4743
rect 2547 4737 2551 4738
rect 2723 4742 2727 4743
rect 2723 4737 2727 4738
rect 2795 4742 2799 4743
rect 2795 4737 2799 4738
rect 3075 4742 3079 4743
rect 3075 4737 3079 4738
rect 3371 4742 3375 4743
rect 3371 4737 3375 4738
rect 3651 4742 3655 4743
rect 3651 4737 3655 4738
rect 3799 4742 3803 4743
rect 3799 4737 3803 4738
rect 158 4732 164 4733
rect 110 4731 116 4732
rect 110 4727 111 4731
rect 115 4727 116 4731
rect 158 4728 159 4732
rect 163 4728 164 4732
rect 158 4727 164 4728
rect 294 4732 300 4733
rect 294 4728 295 4732
rect 299 4728 300 4732
rect 294 4727 300 4728
rect 430 4732 436 4733
rect 430 4728 431 4732
rect 435 4728 436 4732
rect 430 4727 436 4728
rect 566 4732 572 4733
rect 566 4728 567 4732
rect 571 4728 572 4732
rect 566 4727 572 4728
rect 702 4732 708 4733
rect 702 4728 703 4732
rect 707 4728 708 4732
rect 702 4727 708 4728
rect 1934 4731 1940 4732
rect 1934 4727 1935 4731
rect 1939 4727 1940 4731
rect 110 4726 116 4727
rect 112 4699 114 4726
rect 160 4699 162 4727
rect 296 4699 298 4727
rect 432 4699 434 4727
rect 568 4699 570 4727
rect 704 4699 706 4727
rect 1934 4726 1940 4727
rect 1936 4699 1938 4726
rect 111 4698 115 4699
rect 111 4693 115 4694
rect 159 4698 163 4699
rect 159 4693 163 4694
rect 295 4698 299 4699
rect 295 4693 299 4694
rect 431 4698 435 4699
rect 431 4693 435 4694
rect 567 4698 571 4699
rect 567 4693 571 4694
rect 703 4698 707 4699
rect 703 4693 707 4694
rect 1935 4698 1939 4699
rect 1935 4693 1939 4694
rect 112 4670 114 4693
rect 110 4669 116 4670
rect 160 4669 162 4693
rect 296 4669 298 4693
rect 432 4669 434 4693
rect 568 4669 570 4693
rect 704 4669 706 4693
rect 1936 4670 1938 4693
rect 1976 4677 1978 4737
rect 1974 4676 1980 4677
rect 2020 4676 2022 4737
rect 2196 4676 2198 4737
rect 2372 4676 2374 4737
rect 2548 4676 2550 4737
rect 2724 4676 2726 4737
rect 3800 4677 3802 4737
rect 3840 4691 3842 4751
rect 3860 4691 3862 4752
rect 4044 4691 4046 4752
rect 4268 4691 4270 4752
rect 4508 4691 4510 4752
rect 4756 4691 4758 4752
rect 5012 4691 5014 4752
rect 5276 4691 5278 4752
rect 5516 4691 5518 4752
rect 5662 4751 5668 4752
rect 5664 4691 5666 4751
rect 3839 4690 3843 4691
rect 3839 4685 3843 4686
rect 3859 4690 3863 4691
rect 3859 4685 3863 4686
rect 3995 4690 3999 4691
rect 3995 4685 3999 4686
rect 4043 4690 4047 4691
rect 4043 4685 4047 4686
rect 4131 4690 4135 4691
rect 4131 4685 4135 4686
rect 4267 4690 4271 4691
rect 4267 4685 4271 4686
rect 4403 4690 4407 4691
rect 4403 4685 4407 4686
rect 4507 4690 4511 4691
rect 4507 4685 4511 4686
rect 4539 4690 4543 4691
rect 4539 4685 4543 4686
rect 4675 4690 4679 4691
rect 4675 4685 4679 4686
rect 4755 4690 4759 4691
rect 4755 4685 4759 4686
rect 4819 4690 4823 4691
rect 4819 4685 4823 4686
rect 4963 4690 4967 4691
rect 4963 4685 4967 4686
rect 5011 4690 5015 4691
rect 5011 4685 5015 4686
rect 5107 4690 5111 4691
rect 5107 4685 5111 4686
rect 5243 4690 5247 4691
rect 5243 4685 5247 4686
rect 5275 4690 5279 4691
rect 5275 4685 5279 4686
rect 5379 4690 5383 4691
rect 5379 4685 5383 4686
rect 5515 4690 5519 4691
rect 5515 4685 5519 4686
rect 5663 4690 5667 4691
rect 5663 4685 5667 4686
rect 3798 4676 3804 4677
rect 1974 4672 1975 4676
rect 1979 4672 1980 4676
rect 1974 4671 1980 4672
rect 2018 4675 2024 4676
rect 2018 4671 2019 4675
rect 2023 4671 2024 4675
rect 2018 4670 2024 4671
rect 2194 4675 2200 4676
rect 2194 4671 2195 4675
rect 2199 4671 2200 4675
rect 2194 4670 2200 4671
rect 2370 4675 2376 4676
rect 2370 4671 2371 4675
rect 2375 4671 2376 4675
rect 2370 4670 2376 4671
rect 2546 4675 2552 4676
rect 2546 4671 2547 4675
rect 2551 4671 2552 4675
rect 2546 4670 2552 4671
rect 2722 4675 2728 4676
rect 2722 4671 2723 4675
rect 2727 4671 2728 4675
rect 3798 4672 3799 4676
rect 3803 4672 3804 4676
rect 3798 4671 3804 4672
rect 2722 4670 2728 4671
rect 1934 4669 1940 4670
rect 110 4665 111 4669
rect 115 4665 116 4669
rect 110 4664 116 4665
rect 158 4668 164 4669
rect 158 4664 159 4668
rect 163 4664 164 4668
rect 158 4663 164 4664
rect 294 4668 300 4669
rect 294 4664 295 4668
rect 299 4664 300 4668
rect 294 4663 300 4664
rect 430 4668 436 4669
rect 430 4664 431 4668
rect 435 4664 436 4668
rect 430 4663 436 4664
rect 566 4668 572 4669
rect 566 4664 567 4668
rect 571 4664 572 4668
rect 566 4663 572 4664
rect 702 4668 708 4669
rect 702 4664 703 4668
rect 707 4664 708 4668
rect 1934 4665 1935 4669
rect 1939 4665 1940 4669
rect 1934 4664 1940 4665
rect 702 4663 708 4664
rect 2046 4660 2052 4661
rect 1974 4659 1980 4660
rect 1974 4655 1975 4659
rect 1979 4655 1980 4659
rect 2046 4656 2047 4660
rect 2051 4656 2052 4660
rect 2046 4655 2052 4656
rect 2222 4660 2228 4661
rect 2222 4656 2223 4660
rect 2227 4656 2228 4660
rect 2222 4655 2228 4656
rect 2398 4660 2404 4661
rect 2398 4656 2399 4660
rect 2403 4656 2404 4660
rect 2398 4655 2404 4656
rect 2574 4660 2580 4661
rect 2574 4656 2575 4660
rect 2579 4656 2580 4660
rect 2574 4655 2580 4656
rect 2750 4660 2756 4661
rect 2750 4656 2751 4660
rect 2755 4656 2756 4660
rect 2750 4655 2756 4656
rect 3798 4659 3804 4660
rect 3798 4655 3799 4659
rect 3803 4655 3804 4659
rect 1974 4654 1980 4655
rect 130 4653 136 4654
rect 110 4652 116 4653
rect 110 4648 111 4652
rect 115 4648 116 4652
rect 130 4649 131 4653
rect 135 4649 136 4653
rect 130 4648 136 4649
rect 266 4653 272 4654
rect 266 4649 267 4653
rect 271 4649 272 4653
rect 266 4648 272 4649
rect 402 4653 408 4654
rect 402 4649 403 4653
rect 407 4649 408 4653
rect 402 4648 408 4649
rect 538 4653 544 4654
rect 538 4649 539 4653
rect 543 4649 544 4653
rect 538 4648 544 4649
rect 674 4653 680 4654
rect 674 4649 675 4653
rect 679 4649 680 4653
rect 674 4648 680 4649
rect 1934 4652 1940 4653
rect 1934 4648 1935 4652
rect 1939 4648 1940 4652
rect 110 4647 116 4648
rect 112 4575 114 4647
rect 132 4575 134 4648
rect 268 4575 270 4648
rect 404 4575 406 4648
rect 540 4575 542 4648
rect 676 4575 678 4648
rect 1934 4647 1940 4648
rect 1936 4575 1938 4647
rect 1976 4627 1978 4654
rect 2048 4627 2050 4655
rect 2224 4627 2226 4655
rect 2400 4627 2402 4655
rect 2576 4627 2578 4655
rect 2752 4627 2754 4655
rect 3798 4654 3804 4655
rect 3800 4627 3802 4654
rect 1975 4626 1979 4627
rect 1975 4621 1979 4622
rect 2023 4626 2027 4627
rect 2023 4621 2027 4622
rect 2047 4626 2051 4627
rect 2047 4621 2051 4622
rect 2223 4626 2227 4627
rect 2223 4621 2227 4622
rect 2263 4626 2267 4627
rect 2263 4621 2267 4622
rect 2399 4626 2403 4627
rect 2399 4621 2403 4622
rect 2527 4626 2531 4627
rect 2527 4621 2531 4622
rect 2575 4626 2579 4627
rect 2575 4621 2579 4622
rect 2751 4626 2755 4627
rect 2751 4621 2755 4622
rect 2775 4626 2779 4627
rect 2775 4621 2779 4622
rect 3015 4626 3019 4627
rect 3015 4621 3019 4622
rect 3247 4626 3251 4627
rect 3247 4621 3251 4622
rect 3471 4626 3475 4627
rect 3471 4621 3475 4622
rect 3679 4626 3683 4627
rect 3679 4621 3683 4622
rect 3799 4626 3803 4627
rect 3840 4625 3842 4685
rect 3799 4621 3803 4622
rect 3838 4624 3844 4625
rect 3860 4624 3862 4685
rect 3996 4624 3998 4685
rect 4132 4624 4134 4685
rect 4268 4624 4270 4685
rect 4404 4624 4406 4685
rect 4540 4624 4542 4685
rect 4676 4624 4678 4685
rect 4820 4624 4822 4685
rect 4964 4624 4966 4685
rect 5108 4624 5110 4685
rect 5244 4624 5246 4685
rect 5380 4624 5382 4685
rect 5516 4624 5518 4685
rect 5664 4625 5666 4685
rect 5662 4624 5668 4625
rect 1976 4598 1978 4621
rect 1974 4597 1980 4598
rect 2024 4597 2026 4621
rect 2264 4597 2266 4621
rect 2528 4597 2530 4621
rect 2776 4597 2778 4621
rect 3016 4597 3018 4621
rect 3248 4597 3250 4621
rect 3472 4597 3474 4621
rect 3680 4597 3682 4621
rect 3800 4598 3802 4621
rect 3838 4620 3839 4624
rect 3843 4620 3844 4624
rect 3838 4619 3844 4620
rect 3858 4623 3864 4624
rect 3858 4619 3859 4623
rect 3863 4619 3864 4623
rect 3858 4618 3864 4619
rect 3994 4623 4000 4624
rect 3994 4619 3995 4623
rect 3999 4619 4000 4623
rect 3994 4618 4000 4619
rect 4130 4623 4136 4624
rect 4130 4619 4131 4623
rect 4135 4619 4136 4623
rect 4130 4618 4136 4619
rect 4266 4623 4272 4624
rect 4266 4619 4267 4623
rect 4271 4619 4272 4623
rect 4266 4618 4272 4619
rect 4402 4623 4408 4624
rect 4402 4619 4403 4623
rect 4407 4619 4408 4623
rect 4402 4618 4408 4619
rect 4538 4623 4544 4624
rect 4538 4619 4539 4623
rect 4543 4619 4544 4623
rect 4538 4618 4544 4619
rect 4674 4623 4680 4624
rect 4674 4619 4675 4623
rect 4679 4619 4680 4623
rect 4674 4618 4680 4619
rect 4818 4623 4824 4624
rect 4818 4619 4819 4623
rect 4823 4619 4824 4623
rect 4818 4618 4824 4619
rect 4962 4623 4968 4624
rect 4962 4619 4963 4623
rect 4967 4619 4968 4623
rect 4962 4618 4968 4619
rect 5106 4623 5112 4624
rect 5106 4619 5107 4623
rect 5111 4619 5112 4623
rect 5106 4618 5112 4619
rect 5242 4623 5248 4624
rect 5242 4619 5243 4623
rect 5247 4619 5248 4623
rect 5242 4618 5248 4619
rect 5378 4623 5384 4624
rect 5378 4619 5379 4623
rect 5383 4619 5384 4623
rect 5378 4618 5384 4619
rect 5514 4623 5520 4624
rect 5514 4619 5515 4623
rect 5519 4619 5520 4623
rect 5662 4620 5663 4624
rect 5667 4620 5668 4624
rect 5662 4619 5668 4620
rect 5514 4618 5520 4619
rect 3886 4608 3892 4609
rect 3838 4607 3844 4608
rect 3838 4603 3839 4607
rect 3843 4603 3844 4607
rect 3886 4604 3887 4608
rect 3891 4604 3892 4608
rect 3886 4603 3892 4604
rect 4022 4608 4028 4609
rect 4022 4604 4023 4608
rect 4027 4604 4028 4608
rect 4022 4603 4028 4604
rect 4158 4608 4164 4609
rect 4158 4604 4159 4608
rect 4163 4604 4164 4608
rect 4158 4603 4164 4604
rect 4294 4608 4300 4609
rect 4294 4604 4295 4608
rect 4299 4604 4300 4608
rect 4294 4603 4300 4604
rect 4430 4608 4436 4609
rect 4430 4604 4431 4608
rect 4435 4604 4436 4608
rect 4430 4603 4436 4604
rect 4566 4608 4572 4609
rect 4566 4604 4567 4608
rect 4571 4604 4572 4608
rect 4566 4603 4572 4604
rect 4702 4608 4708 4609
rect 4702 4604 4703 4608
rect 4707 4604 4708 4608
rect 4702 4603 4708 4604
rect 4846 4608 4852 4609
rect 4846 4604 4847 4608
rect 4851 4604 4852 4608
rect 4846 4603 4852 4604
rect 4990 4608 4996 4609
rect 4990 4604 4991 4608
rect 4995 4604 4996 4608
rect 4990 4603 4996 4604
rect 5134 4608 5140 4609
rect 5134 4604 5135 4608
rect 5139 4604 5140 4608
rect 5134 4603 5140 4604
rect 5270 4608 5276 4609
rect 5270 4604 5271 4608
rect 5275 4604 5276 4608
rect 5270 4603 5276 4604
rect 5406 4608 5412 4609
rect 5406 4604 5407 4608
rect 5411 4604 5412 4608
rect 5406 4603 5412 4604
rect 5542 4608 5548 4609
rect 5542 4604 5543 4608
rect 5547 4604 5548 4608
rect 5542 4603 5548 4604
rect 5662 4607 5668 4608
rect 5662 4603 5663 4607
rect 5667 4603 5668 4607
rect 3838 4602 3844 4603
rect 3798 4597 3804 4598
rect 1974 4593 1975 4597
rect 1979 4593 1980 4597
rect 1974 4592 1980 4593
rect 2022 4596 2028 4597
rect 2022 4592 2023 4596
rect 2027 4592 2028 4596
rect 2022 4591 2028 4592
rect 2262 4596 2268 4597
rect 2262 4592 2263 4596
rect 2267 4592 2268 4596
rect 2262 4591 2268 4592
rect 2526 4596 2532 4597
rect 2526 4592 2527 4596
rect 2531 4592 2532 4596
rect 2526 4591 2532 4592
rect 2774 4596 2780 4597
rect 2774 4592 2775 4596
rect 2779 4592 2780 4596
rect 2774 4591 2780 4592
rect 3014 4596 3020 4597
rect 3014 4592 3015 4596
rect 3019 4592 3020 4596
rect 3014 4591 3020 4592
rect 3246 4596 3252 4597
rect 3246 4592 3247 4596
rect 3251 4592 3252 4596
rect 3246 4591 3252 4592
rect 3470 4596 3476 4597
rect 3470 4592 3471 4596
rect 3475 4592 3476 4596
rect 3470 4591 3476 4592
rect 3678 4596 3684 4597
rect 3678 4592 3679 4596
rect 3683 4592 3684 4596
rect 3798 4593 3799 4597
rect 3803 4593 3804 4597
rect 3798 4592 3804 4593
rect 3678 4591 3684 4592
rect 1994 4581 2000 4582
rect 1974 4580 1980 4581
rect 1974 4576 1975 4580
rect 1979 4576 1980 4580
rect 1994 4577 1995 4581
rect 1999 4577 2000 4581
rect 1994 4576 2000 4577
rect 2234 4581 2240 4582
rect 2234 4577 2235 4581
rect 2239 4577 2240 4581
rect 2234 4576 2240 4577
rect 2498 4581 2504 4582
rect 2498 4577 2499 4581
rect 2503 4577 2504 4581
rect 2498 4576 2504 4577
rect 2746 4581 2752 4582
rect 2746 4577 2747 4581
rect 2751 4577 2752 4581
rect 2746 4576 2752 4577
rect 2986 4581 2992 4582
rect 2986 4577 2987 4581
rect 2991 4577 2992 4581
rect 2986 4576 2992 4577
rect 3218 4581 3224 4582
rect 3218 4577 3219 4581
rect 3223 4577 3224 4581
rect 3218 4576 3224 4577
rect 3442 4581 3448 4582
rect 3442 4577 3443 4581
rect 3447 4577 3448 4581
rect 3442 4576 3448 4577
rect 3650 4581 3656 4582
rect 3650 4577 3651 4581
rect 3655 4577 3656 4581
rect 3650 4576 3656 4577
rect 3798 4580 3804 4581
rect 3798 4576 3799 4580
rect 3803 4576 3804 4580
rect 3840 4579 3842 4602
rect 3888 4579 3890 4603
rect 4024 4579 4026 4603
rect 4160 4579 4162 4603
rect 4296 4579 4298 4603
rect 4432 4579 4434 4603
rect 4568 4579 4570 4603
rect 4704 4579 4706 4603
rect 4848 4579 4850 4603
rect 4992 4579 4994 4603
rect 5136 4579 5138 4603
rect 5272 4579 5274 4603
rect 5408 4579 5410 4603
rect 5544 4579 5546 4603
rect 5662 4602 5668 4603
rect 5664 4579 5666 4602
rect 1974 4575 1980 4576
rect 111 4574 115 4575
rect 111 4569 115 4570
rect 131 4574 135 4575
rect 131 4569 135 4570
rect 251 4574 255 4575
rect 251 4569 255 4570
rect 267 4574 271 4575
rect 267 4569 271 4570
rect 403 4574 407 4575
rect 403 4569 407 4570
rect 443 4574 447 4575
rect 443 4569 447 4570
rect 539 4574 543 4575
rect 539 4569 543 4570
rect 651 4574 655 4575
rect 651 4569 655 4570
rect 675 4574 679 4575
rect 675 4569 679 4570
rect 875 4574 879 4575
rect 875 4569 879 4570
rect 1099 4574 1103 4575
rect 1099 4569 1103 4570
rect 1331 4574 1335 4575
rect 1331 4569 1335 4570
rect 1571 4574 1575 4575
rect 1571 4569 1575 4570
rect 1787 4574 1791 4575
rect 1787 4569 1791 4570
rect 1935 4574 1939 4575
rect 1935 4569 1939 4570
rect 112 4509 114 4569
rect 110 4508 116 4509
rect 252 4508 254 4569
rect 444 4508 446 4569
rect 652 4508 654 4569
rect 876 4508 878 4569
rect 1100 4508 1102 4569
rect 1332 4508 1334 4569
rect 1572 4508 1574 4569
rect 1788 4508 1790 4569
rect 1936 4509 1938 4569
rect 1934 4508 1940 4509
rect 110 4504 111 4508
rect 115 4504 116 4508
rect 110 4503 116 4504
rect 250 4507 256 4508
rect 250 4503 251 4507
rect 255 4503 256 4507
rect 250 4502 256 4503
rect 442 4507 448 4508
rect 442 4503 443 4507
rect 447 4503 448 4507
rect 442 4502 448 4503
rect 650 4507 656 4508
rect 650 4503 651 4507
rect 655 4503 656 4507
rect 650 4502 656 4503
rect 874 4507 880 4508
rect 874 4503 875 4507
rect 879 4503 880 4507
rect 874 4502 880 4503
rect 1098 4507 1104 4508
rect 1098 4503 1099 4507
rect 1103 4503 1104 4507
rect 1098 4502 1104 4503
rect 1330 4507 1336 4508
rect 1330 4503 1331 4507
rect 1335 4503 1336 4507
rect 1330 4502 1336 4503
rect 1570 4507 1576 4508
rect 1570 4503 1571 4507
rect 1575 4503 1576 4507
rect 1570 4502 1576 4503
rect 1786 4507 1792 4508
rect 1786 4503 1787 4507
rect 1791 4503 1792 4507
rect 1934 4504 1935 4508
rect 1939 4504 1940 4508
rect 1934 4503 1940 4504
rect 1976 4503 1978 4575
rect 1996 4503 1998 4576
rect 2236 4503 2238 4576
rect 2500 4503 2502 4576
rect 2748 4503 2750 4576
rect 2988 4503 2990 4576
rect 3220 4503 3222 4576
rect 3444 4503 3446 4576
rect 3652 4503 3654 4576
rect 3798 4575 3804 4576
rect 3839 4578 3843 4579
rect 3800 4503 3802 4575
rect 3839 4573 3843 4574
rect 3887 4578 3891 4579
rect 3887 4573 3891 4574
rect 4023 4578 4027 4579
rect 4023 4573 4027 4574
rect 4159 4578 4163 4579
rect 4159 4573 4163 4574
rect 4295 4578 4299 4579
rect 4295 4573 4299 4574
rect 4431 4578 4435 4579
rect 4431 4573 4435 4574
rect 4567 4578 4571 4579
rect 4567 4573 4571 4574
rect 4671 4578 4675 4579
rect 4671 4573 4675 4574
rect 4703 4578 4707 4579
rect 4703 4573 4707 4574
rect 4807 4578 4811 4579
rect 4807 4573 4811 4574
rect 4847 4578 4851 4579
rect 4847 4573 4851 4574
rect 4943 4578 4947 4579
rect 4943 4573 4947 4574
rect 4991 4578 4995 4579
rect 4991 4573 4995 4574
rect 5079 4578 5083 4579
rect 5079 4573 5083 4574
rect 5135 4578 5139 4579
rect 5135 4573 5139 4574
rect 5271 4578 5275 4579
rect 5271 4573 5275 4574
rect 5407 4578 5411 4579
rect 5407 4573 5411 4574
rect 5543 4578 5547 4579
rect 5543 4573 5547 4574
rect 5663 4578 5667 4579
rect 5663 4573 5667 4574
rect 3840 4550 3842 4573
rect 3838 4549 3844 4550
rect 4672 4549 4674 4573
rect 4808 4549 4810 4573
rect 4944 4549 4946 4573
rect 5080 4549 5082 4573
rect 5664 4550 5666 4573
rect 5662 4549 5668 4550
rect 3838 4545 3839 4549
rect 3843 4545 3844 4549
rect 3838 4544 3844 4545
rect 4670 4548 4676 4549
rect 4670 4544 4671 4548
rect 4675 4544 4676 4548
rect 4670 4543 4676 4544
rect 4806 4548 4812 4549
rect 4806 4544 4807 4548
rect 4811 4544 4812 4548
rect 4806 4543 4812 4544
rect 4942 4548 4948 4549
rect 4942 4544 4943 4548
rect 4947 4544 4948 4548
rect 4942 4543 4948 4544
rect 5078 4548 5084 4549
rect 5078 4544 5079 4548
rect 5083 4544 5084 4548
rect 5662 4545 5663 4549
rect 5667 4545 5668 4549
rect 5662 4544 5668 4545
rect 5078 4543 5084 4544
rect 4642 4533 4648 4534
rect 3838 4532 3844 4533
rect 3838 4528 3839 4532
rect 3843 4528 3844 4532
rect 4642 4529 4643 4533
rect 4647 4529 4648 4533
rect 4642 4528 4648 4529
rect 4778 4533 4784 4534
rect 4778 4529 4779 4533
rect 4783 4529 4784 4533
rect 4778 4528 4784 4529
rect 4914 4533 4920 4534
rect 4914 4529 4915 4533
rect 4919 4529 4920 4533
rect 4914 4528 4920 4529
rect 5050 4533 5056 4534
rect 5050 4529 5051 4533
rect 5055 4529 5056 4533
rect 5050 4528 5056 4529
rect 5662 4532 5668 4533
rect 5662 4528 5663 4532
rect 5667 4528 5668 4532
rect 3838 4527 3844 4528
rect 1786 4502 1792 4503
rect 1975 4502 1979 4503
rect 1975 4497 1979 4498
rect 1995 4502 1999 4503
rect 1995 4497 1999 4498
rect 2235 4502 2239 4503
rect 2235 4497 2239 4498
rect 2267 4502 2271 4503
rect 2267 4497 2271 4498
rect 2499 4502 2503 4503
rect 2499 4497 2503 4498
rect 2515 4502 2519 4503
rect 2515 4497 2519 4498
rect 2747 4502 2751 4503
rect 2747 4497 2751 4498
rect 2971 4502 2975 4503
rect 2971 4497 2975 4498
rect 2987 4502 2991 4503
rect 2987 4497 2991 4498
rect 3187 4502 3191 4503
rect 3187 4497 3191 4498
rect 3219 4502 3223 4503
rect 3219 4497 3223 4498
rect 3395 4502 3399 4503
rect 3395 4497 3399 4498
rect 3443 4502 3447 4503
rect 3443 4497 3447 4498
rect 3611 4502 3615 4503
rect 3611 4497 3615 4498
rect 3651 4502 3655 4503
rect 3651 4497 3655 4498
rect 3799 4502 3803 4503
rect 3799 4497 3803 4498
rect 278 4492 284 4493
rect 110 4491 116 4492
rect 110 4487 111 4491
rect 115 4487 116 4491
rect 278 4488 279 4492
rect 283 4488 284 4492
rect 278 4487 284 4488
rect 470 4492 476 4493
rect 470 4488 471 4492
rect 475 4488 476 4492
rect 470 4487 476 4488
rect 678 4492 684 4493
rect 678 4488 679 4492
rect 683 4488 684 4492
rect 678 4487 684 4488
rect 902 4492 908 4493
rect 902 4488 903 4492
rect 907 4488 908 4492
rect 902 4487 908 4488
rect 1126 4492 1132 4493
rect 1126 4488 1127 4492
rect 1131 4488 1132 4492
rect 1126 4487 1132 4488
rect 1358 4492 1364 4493
rect 1358 4488 1359 4492
rect 1363 4488 1364 4492
rect 1358 4487 1364 4488
rect 1598 4492 1604 4493
rect 1598 4488 1599 4492
rect 1603 4488 1604 4492
rect 1598 4487 1604 4488
rect 1814 4492 1820 4493
rect 1814 4488 1815 4492
rect 1819 4488 1820 4492
rect 1814 4487 1820 4488
rect 1934 4491 1940 4492
rect 1934 4487 1935 4491
rect 1939 4487 1940 4491
rect 110 4486 116 4487
rect 112 4463 114 4486
rect 280 4463 282 4487
rect 472 4463 474 4487
rect 680 4463 682 4487
rect 904 4463 906 4487
rect 1128 4463 1130 4487
rect 1360 4463 1362 4487
rect 1600 4463 1602 4487
rect 1816 4463 1818 4487
rect 1934 4486 1940 4487
rect 1936 4463 1938 4486
rect 111 4462 115 4463
rect 111 4457 115 4458
rect 279 4462 283 4463
rect 279 4457 283 4458
rect 471 4462 475 4463
rect 471 4457 475 4458
rect 511 4462 515 4463
rect 511 4457 515 4458
rect 679 4462 683 4463
rect 679 4457 683 4458
rect 687 4462 691 4463
rect 687 4457 691 4458
rect 871 4462 875 4463
rect 871 4457 875 4458
rect 903 4462 907 4463
rect 903 4457 907 4458
rect 1071 4462 1075 4463
rect 1071 4457 1075 4458
rect 1127 4462 1131 4463
rect 1127 4457 1131 4458
rect 1279 4462 1283 4463
rect 1279 4457 1283 4458
rect 1359 4462 1363 4463
rect 1359 4457 1363 4458
rect 1495 4462 1499 4463
rect 1495 4457 1499 4458
rect 1599 4462 1603 4463
rect 1599 4457 1603 4458
rect 1719 4462 1723 4463
rect 1719 4457 1723 4458
rect 1815 4462 1819 4463
rect 1815 4457 1819 4458
rect 1935 4462 1939 4463
rect 1935 4457 1939 4458
rect 112 4434 114 4457
rect 110 4433 116 4434
rect 512 4433 514 4457
rect 688 4433 690 4457
rect 872 4433 874 4457
rect 1072 4433 1074 4457
rect 1280 4433 1282 4457
rect 1496 4433 1498 4457
rect 1720 4433 1722 4457
rect 1936 4434 1938 4457
rect 1976 4437 1978 4497
rect 1974 4436 1980 4437
rect 2268 4436 2270 4497
rect 2516 4436 2518 4497
rect 2748 4436 2750 4497
rect 2972 4436 2974 4497
rect 3188 4436 3190 4497
rect 3396 4436 3398 4497
rect 3612 4436 3614 4497
rect 3800 4437 3802 4497
rect 3840 4463 3842 4527
rect 4644 4463 4646 4528
rect 4780 4463 4782 4528
rect 4916 4463 4918 4528
rect 5052 4463 5054 4528
rect 5662 4527 5668 4528
rect 5664 4463 5666 4527
rect 3839 4462 3843 4463
rect 3839 4457 3843 4458
rect 4347 4462 4351 4463
rect 4347 4457 4351 4458
rect 4483 4462 4487 4463
rect 4483 4457 4487 4458
rect 4619 4462 4623 4463
rect 4619 4457 4623 4458
rect 4643 4462 4647 4463
rect 4643 4457 4647 4458
rect 4755 4462 4759 4463
rect 4755 4457 4759 4458
rect 4779 4462 4783 4463
rect 4779 4457 4783 4458
rect 4891 4462 4895 4463
rect 4891 4457 4895 4458
rect 4915 4462 4919 4463
rect 4915 4457 4919 4458
rect 5051 4462 5055 4463
rect 5051 4457 5055 4458
rect 5663 4462 5667 4463
rect 5663 4457 5667 4458
rect 3798 4436 3804 4437
rect 1934 4433 1940 4434
rect 110 4429 111 4433
rect 115 4429 116 4433
rect 110 4428 116 4429
rect 510 4432 516 4433
rect 510 4428 511 4432
rect 515 4428 516 4432
rect 510 4427 516 4428
rect 686 4432 692 4433
rect 686 4428 687 4432
rect 691 4428 692 4432
rect 686 4427 692 4428
rect 870 4432 876 4433
rect 870 4428 871 4432
rect 875 4428 876 4432
rect 870 4427 876 4428
rect 1070 4432 1076 4433
rect 1070 4428 1071 4432
rect 1075 4428 1076 4432
rect 1070 4427 1076 4428
rect 1278 4432 1284 4433
rect 1278 4428 1279 4432
rect 1283 4428 1284 4432
rect 1278 4427 1284 4428
rect 1494 4432 1500 4433
rect 1494 4428 1495 4432
rect 1499 4428 1500 4432
rect 1494 4427 1500 4428
rect 1718 4432 1724 4433
rect 1718 4428 1719 4432
rect 1723 4428 1724 4432
rect 1934 4429 1935 4433
rect 1939 4429 1940 4433
rect 1974 4432 1975 4436
rect 1979 4432 1980 4436
rect 1974 4431 1980 4432
rect 2266 4435 2272 4436
rect 2266 4431 2267 4435
rect 2271 4431 2272 4435
rect 2266 4430 2272 4431
rect 2514 4435 2520 4436
rect 2514 4431 2515 4435
rect 2519 4431 2520 4435
rect 2514 4430 2520 4431
rect 2746 4435 2752 4436
rect 2746 4431 2747 4435
rect 2751 4431 2752 4435
rect 2746 4430 2752 4431
rect 2970 4435 2976 4436
rect 2970 4431 2971 4435
rect 2975 4431 2976 4435
rect 2970 4430 2976 4431
rect 3186 4435 3192 4436
rect 3186 4431 3187 4435
rect 3191 4431 3192 4435
rect 3186 4430 3192 4431
rect 3394 4435 3400 4436
rect 3394 4431 3395 4435
rect 3399 4431 3400 4435
rect 3394 4430 3400 4431
rect 3610 4435 3616 4436
rect 3610 4431 3611 4435
rect 3615 4431 3616 4435
rect 3798 4432 3799 4436
rect 3803 4432 3804 4436
rect 3798 4431 3804 4432
rect 3610 4430 3616 4431
rect 1934 4428 1940 4429
rect 1718 4427 1724 4428
rect 2294 4420 2300 4421
rect 1974 4419 1980 4420
rect 482 4417 488 4418
rect 110 4416 116 4417
rect 110 4412 111 4416
rect 115 4412 116 4416
rect 482 4413 483 4417
rect 487 4413 488 4417
rect 482 4412 488 4413
rect 658 4417 664 4418
rect 658 4413 659 4417
rect 663 4413 664 4417
rect 658 4412 664 4413
rect 842 4417 848 4418
rect 842 4413 843 4417
rect 847 4413 848 4417
rect 842 4412 848 4413
rect 1042 4417 1048 4418
rect 1042 4413 1043 4417
rect 1047 4413 1048 4417
rect 1042 4412 1048 4413
rect 1250 4417 1256 4418
rect 1250 4413 1251 4417
rect 1255 4413 1256 4417
rect 1250 4412 1256 4413
rect 1466 4417 1472 4418
rect 1466 4413 1467 4417
rect 1471 4413 1472 4417
rect 1466 4412 1472 4413
rect 1690 4417 1696 4418
rect 1690 4413 1691 4417
rect 1695 4413 1696 4417
rect 1690 4412 1696 4413
rect 1934 4416 1940 4417
rect 1934 4412 1935 4416
rect 1939 4412 1940 4416
rect 1974 4415 1975 4419
rect 1979 4415 1980 4419
rect 2294 4416 2295 4420
rect 2299 4416 2300 4420
rect 2294 4415 2300 4416
rect 2542 4420 2548 4421
rect 2542 4416 2543 4420
rect 2547 4416 2548 4420
rect 2542 4415 2548 4416
rect 2774 4420 2780 4421
rect 2774 4416 2775 4420
rect 2779 4416 2780 4420
rect 2774 4415 2780 4416
rect 2998 4420 3004 4421
rect 2998 4416 2999 4420
rect 3003 4416 3004 4420
rect 2998 4415 3004 4416
rect 3214 4420 3220 4421
rect 3214 4416 3215 4420
rect 3219 4416 3220 4420
rect 3214 4415 3220 4416
rect 3422 4420 3428 4421
rect 3422 4416 3423 4420
rect 3427 4416 3428 4420
rect 3422 4415 3428 4416
rect 3638 4420 3644 4421
rect 3638 4416 3639 4420
rect 3643 4416 3644 4420
rect 3638 4415 3644 4416
rect 3798 4419 3804 4420
rect 3798 4415 3799 4419
rect 3803 4415 3804 4419
rect 1974 4414 1980 4415
rect 110 4411 116 4412
rect 112 4347 114 4411
rect 484 4347 486 4412
rect 660 4347 662 4412
rect 844 4347 846 4412
rect 1044 4347 1046 4412
rect 1252 4347 1254 4412
rect 1468 4347 1470 4412
rect 1692 4347 1694 4412
rect 1934 4411 1940 4412
rect 1936 4347 1938 4411
rect 1976 4379 1978 4414
rect 2296 4379 2298 4415
rect 2544 4379 2546 4415
rect 2776 4379 2778 4415
rect 3000 4379 3002 4415
rect 3216 4379 3218 4415
rect 3424 4379 3426 4415
rect 3640 4379 3642 4415
rect 3798 4414 3804 4415
rect 3800 4379 3802 4414
rect 3840 4397 3842 4457
rect 3838 4396 3844 4397
rect 4348 4396 4350 4457
rect 4484 4396 4486 4457
rect 4620 4396 4622 4457
rect 4756 4396 4758 4457
rect 4892 4396 4894 4457
rect 5664 4397 5666 4457
rect 5662 4396 5668 4397
rect 3838 4392 3839 4396
rect 3843 4392 3844 4396
rect 3838 4391 3844 4392
rect 4346 4395 4352 4396
rect 4346 4391 4347 4395
rect 4351 4391 4352 4395
rect 4346 4390 4352 4391
rect 4482 4395 4488 4396
rect 4482 4391 4483 4395
rect 4487 4391 4488 4395
rect 4482 4390 4488 4391
rect 4618 4395 4624 4396
rect 4618 4391 4619 4395
rect 4623 4391 4624 4395
rect 4618 4390 4624 4391
rect 4754 4395 4760 4396
rect 4754 4391 4755 4395
rect 4759 4391 4760 4395
rect 4754 4390 4760 4391
rect 4890 4395 4896 4396
rect 4890 4391 4891 4395
rect 4895 4391 4896 4395
rect 5662 4392 5663 4396
rect 5667 4392 5668 4396
rect 5662 4391 5668 4392
rect 4890 4390 4896 4391
rect 4374 4380 4380 4381
rect 3838 4379 3844 4380
rect 1975 4378 1979 4379
rect 1975 4373 1979 4374
rect 2023 4378 2027 4379
rect 2023 4373 2027 4374
rect 2199 4378 2203 4379
rect 2199 4373 2203 4374
rect 2295 4378 2299 4379
rect 2295 4373 2299 4374
rect 2399 4378 2403 4379
rect 2399 4373 2403 4374
rect 2543 4378 2547 4379
rect 2543 4373 2547 4374
rect 2591 4378 2595 4379
rect 2591 4373 2595 4374
rect 2775 4378 2779 4379
rect 2775 4373 2779 4374
rect 2951 4378 2955 4379
rect 2951 4373 2955 4374
rect 2999 4378 3003 4379
rect 2999 4373 3003 4374
rect 3135 4378 3139 4379
rect 3135 4373 3139 4374
rect 3215 4378 3219 4379
rect 3215 4373 3219 4374
rect 3319 4378 3323 4379
rect 3319 4373 3323 4374
rect 3423 4378 3427 4379
rect 3423 4373 3427 4374
rect 3639 4378 3643 4379
rect 3639 4373 3643 4374
rect 3799 4378 3803 4379
rect 3838 4375 3839 4379
rect 3843 4375 3844 4379
rect 4374 4376 4375 4380
rect 4379 4376 4380 4380
rect 4374 4375 4380 4376
rect 4510 4380 4516 4381
rect 4510 4376 4511 4380
rect 4515 4376 4516 4380
rect 4510 4375 4516 4376
rect 4646 4380 4652 4381
rect 4646 4376 4647 4380
rect 4651 4376 4652 4380
rect 4646 4375 4652 4376
rect 4782 4380 4788 4381
rect 4782 4376 4783 4380
rect 4787 4376 4788 4380
rect 4782 4375 4788 4376
rect 4918 4380 4924 4381
rect 4918 4376 4919 4380
rect 4923 4376 4924 4380
rect 4918 4375 4924 4376
rect 5662 4379 5668 4380
rect 5662 4375 5663 4379
rect 5667 4375 5668 4379
rect 3838 4374 3844 4375
rect 3799 4373 3803 4374
rect 1976 4350 1978 4373
rect 1974 4349 1980 4350
rect 2024 4349 2026 4373
rect 2200 4349 2202 4373
rect 2400 4349 2402 4373
rect 2592 4349 2594 4373
rect 2776 4349 2778 4373
rect 2952 4349 2954 4373
rect 3136 4349 3138 4373
rect 3320 4349 3322 4373
rect 3800 4350 3802 4373
rect 3798 4349 3804 4350
rect 111 4346 115 4347
rect 111 4341 115 4342
rect 483 4346 487 4347
rect 483 4341 487 4342
rect 659 4346 663 4347
rect 659 4341 663 4342
rect 715 4346 719 4347
rect 715 4341 719 4342
rect 843 4346 847 4347
rect 843 4341 847 4342
rect 851 4346 855 4347
rect 851 4341 855 4342
rect 987 4346 991 4347
rect 987 4341 991 4342
rect 1043 4346 1047 4347
rect 1043 4341 1047 4342
rect 1123 4346 1127 4347
rect 1123 4341 1127 4342
rect 1251 4346 1255 4347
rect 1251 4341 1255 4342
rect 1259 4346 1263 4347
rect 1259 4341 1263 4342
rect 1395 4346 1399 4347
rect 1395 4341 1399 4342
rect 1467 4346 1471 4347
rect 1467 4341 1471 4342
rect 1531 4346 1535 4347
rect 1531 4341 1535 4342
rect 1667 4346 1671 4347
rect 1667 4341 1671 4342
rect 1691 4346 1695 4347
rect 1691 4341 1695 4342
rect 1935 4346 1939 4347
rect 1974 4345 1975 4349
rect 1979 4345 1980 4349
rect 1974 4344 1980 4345
rect 2022 4348 2028 4349
rect 2022 4344 2023 4348
rect 2027 4344 2028 4348
rect 2022 4343 2028 4344
rect 2198 4348 2204 4349
rect 2198 4344 2199 4348
rect 2203 4344 2204 4348
rect 2198 4343 2204 4344
rect 2398 4348 2404 4349
rect 2398 4344 2399 4348
rect 2403 4344 2404 4348
rect 2398 4343 2404 4344
rect 2590 4348 2596 4349
rect 2590 4344 2591 4348
rect 2595 4344 2596 4348
rect 2590 4343 2596 4344
rect 2774 4348 2780 4349
rect 2774 4344 2775 4348
rect 2779 4344 2780 4348
rect 2774 4343 2780 4344
rect 2950 4348 2956 4349
rect 2950 4344 2951 4348
rect 2955 4344 2956 4348
rect 2950 4343 2956 4344
rect 3134 4348 3140 4349
rect 3134 4344 3135 4348
rect 3139 4344 3140 4348
rect 3134 4343 3140 4344
rect 3318 4348 3324 4349
rect 3318 4344 3319 4348
rect 3323 4344 3324 4348
rect 3798 4345 3799 4349
rect 3803 4345 3804 4349
rect 3798 4344 3804 4345
rect 3318 4343 3324 4344
rect 1935 4341 1939 4342
rect 112 4281 114 4341
rect 110 4280 116 4281
rect 716 4280 718 4341
rect 852 4280 854 4341
rect 988 4280 990 4341
rect 1124 4280 1126 4341
rect 1260 4280 1262 4341
rect 1396 4280 1398 4341
rect 1532 4280 1534 4341
rect 1668 4280 1670 4341
rect 1936 4281 1938 4341
rect 3840 4335 3842 4374
rect 4376 4335 4378 4375
rect 4512 4335 4514 4375
rect 4648 4335 4650 4375
rect 4784 4335 4786 4375
rect 4920 4335 4922 4375
rect 5662 4374 5668 4375
rect 5664 4335 5666 4374
rect 3839 4334 3843 4335
rect 1994 4333 2000 4334
rect 1974 4332 1980 4333
rect 1974 4328 1975 4332
rect 1979 4328 1980 4332
rect 1994 4329 1995 4333
rect 1999 4329 2000 4333
rect 1994 4328 2000 4329
rect 2170 4333 2176 4334
rect 2170 4329 2171 4333
rect 2175 4329 2176 4333
rect 2170 4328 2176 4329
rect 2370 4333 2376 4334
rect 2370 4329 2371 4333
rect 2375 4329 2376 4333
rect 2370 4328 2376 4329
rect 2562 4333 2568 4334
rect 2562 4329 2563 4333
rect 2567 4329 2568 4333
rect 2562 4328 2568 4329
rect 2746 4333 2752 4334
rect 2746 4329 2747 4333
rect 2751 4329 2752 4333
rect 2746 4328 2752 4329
rect 2922 4333 2928 4334
rect 2922 4329 2923 4333
rect 2927 4329 2928 4333
rect 2922 4328 2928 4329
rect 3106 4333 3112 4334
rect 3106 4329 3107 4333
rect 3111 4329 3112 4333
rect 3106 4328 3112 4329
rect 3290 4333 3296 4334
rect 3290 4329 3291 4333
rect 3295 4329 3296 4333
rect 3290 4328 3296 4329
rect 3798 4332 3804 4333
rect 3798 4328 3799 4332
rect 3803 4328 3804 4332
rect 3839 4329 3843 4330
rect 4135 4334 4139 4335
rect 4135 4329 4139 4330
rect 4271 4334 4275 4335
rect 4271 4329 4275 4330
rect 4375 4334 4379 4335
rect 4375 4329 4379 4330
rect 4407 4334 4411 4335
rect 4407 4329 4411 4330
rect 4511 4334 4515 4335
rect 4511 4329 4515 4330
rect 4543 4334 4547 4335
rect 4543 4329 4547 4330
rect 4647 4334 4651 4335
rect 4647 4329 4651 4330
rect 4679 4334 4683 4335
rect 4679 4329 4683 4330
rect 4783 4334 4787 4335
rect 4783 4329 4787 4330
rect 4919 4334 4923 4335
rect 4919 4329 4923 4330
rect 5663 4334 5667 4335
rect 5663 4329 5667 4330
rect 1974 4327 1980 4328
rect 1934 4280 1940 4281
rect 110 4276 111 4280
rect 115 4276 116 4280
rect 110 4275 116 4276
rect 714 4279 720 4280
rect 714 4275 715 4279
rect 719 4275 720 4279
rect 714 4274 720 4275
rect 850 4279 856 4280
rect 850 4275 851 4279
rect 855 4275 856 4279
rect 850 4274 856 4275
rect 986 4279 992 4280
rect 986 4275 987 4279
rect 991 4275 992 4279
rect 986 4274 992 4275
rect 1122 4279 1128 4280
rect 1122 4275 1123 4279
rect 1127 4275 1128 4279
rect 1122 4274 1128 4275
rect 1258 4279 1264 4280
rect 1258 4275 1259 4279
rect 1263 4275 1264 4279
rect 1258 4274 1264 4275
rect 1394 4279 1400 4280
rect 1394 4275 1395 4279
rect 1399 4275 1400 4279
rect 1394 4274 1400 4275
rect 1530 4279 1536 4280
rect 1530 4275 1531 4279
rect 1535 4275 1536 4279
rect 1530 4274 1536 4275
rect 1666 4279 1672 4280
rect 1666 4275 1667 4279
rect 1671 4275 1672 4279
rect 1934 4276 1935 4280
rect 1939 4276 1940 4280
rect 1934 4275 1940 4276
rect 1666 4274 1672 4275
rect 742 4264 748 4265
rect 110 4263 116 4264
rect 110 4259 111 4263
rect 115 4259 116 4263
rect 742 4260 743 4264
rect 747 4260 748 4264
rect 742 4259 748 4260
rect 878 4264 884 4265
rect 878 4260 879 4264
rect 883 4260 884 4264
rect 878 4259 884 4260
rect 1014 4264 1020 4265
rect 1014 4260 1015 4264
rect 1019 4260 1020 4264
rect 1014 4259 1020 4260
rect 1150 4264 1156 4265
rect 1150 4260 1151 4264
rect 1155 4260 1156 4264
rect 1150 4259 1156 4260
rect 1286 4264 1292 4265
rect 1286 4260 1287 4264
rect 1291 4260 1292 4264
rect 1286 4259 1292 4260
rect 1422 4264 1428 4265
rect 1422 4260 1423 4264
rect 1427 4260 1428 4264
rect 1422 4259 1428 4260
rect 1558 4264 1564 4265
rect 1558 4260 1559 4264
rect 1563 4260 1564 4264
rect 1558 4259 1564 4260
rect 1694 4264 1700 4265
rect 1694 4260 1695 4264
rect 1699 4260 1700 4264
rect 1694 4259 1700 4260
rect 1934 4263 1940 4264
rect 1976 4263 1978 4327
rect 1996 4263 1998 4328
rect 2172 4263 2174 4328
rect 2372 4263 2374 4328
rect 2564 4263 2566 4328
rect 2748 4263 2750 4328
rect 2924 4263 2926 4328
rect 3108 4263 3110 4328
rect 3292 4263 3294 4328
rect 3798 4327 3804 4328
rect 3800 4263 3802 4327
rect 3840 4306 3842 4329
rect 3838 4305 3844 4306
rect 4136 4305 4138 4329
rect 4272 4305 4274 4329
rect 4408 4305 4410 4329
rect 4544 4305 4546 4329
rect 4680 4305 4682 4329
rect 5664 4306 5666 4329
rect 5662 4305 5668 4306
rect 3838 4301 3839 4305
rect 3843 4301 3844 4305
rect 3838 4300 3844 4301
rect 4134 4304 4140 4305
rect 4134 4300 4135 4304
rect 4139 4300 4140 4304
rect 4134 4299 4140 4300
rect 4270 4304 4276 4305
rect 4270 4300 4271 4304
rect 4275 4300 4276 4304
rect 4270 4299 4276 4300
rect 4406 4304 4412 4305
rect 4406 4300 4407 4304
rect 4411 4300 4412 4304
rect 4406 4299 4412 4300
rect 4542 4304 4548 4305
rect 4542 4300 4543 4304
rect 4547 4300 4548 4304
rect 4542 4299 4548 4300
rect 4678 4304 4684 4305
rect 4678 4300 4679 4304
rect 4683 4300 4684 4304
rect 5662 4301 5663 4305
rect 5667 4301 5668 4305
rect 5662 4300 5668 4301
rect 4678 4299 4684 4300
rect 4106 4289 4112 4290
rect 3838 4288 3844 4289
rect 3838 4284 3839 4288
rect 3843 4284 3844 4288
rect 4106 4285 4107 4289
rect 4111 4285 4112 4289
rect 4106 4284 4112 4285
rect 4242 4289 4248 4290
rect 4242 4285 4243 4289
rect 4247 4285 4248 4289
rect 4242 4284 4248 4285
rect 4378 4289 4384 4290
rect 4378 4285 4379 4289
rect 4383 4285 4384 4289
rect 4378 4284 4384 4285
rect 4514 4289 4520 4290
rect 4514 4285 4515 4289
rect 4519 4285 4520 4289
rect 4514 4284 4520 4285
rect 4650 4289 4656 4290
rect 4650 4285 4651 4289
rect 4655 4285 4656 4289
rect 4650 4284 4656 4285
rect 5662 4288 5668 4289
rect 5662 4284 5663 4288
rect 5667 4284 5668 4288
rect 3838 4283 3844 4284
rect 1934 4259 1935 4263
rect 1939 4259 1940 4263
rect 110 4258 116 4259
rect 112 4227 114 4258
rect 744 4227 746 4259
rect 880 4227 882 4259
rect 1016 4227 1018 4259
rect 1152 4227 1154 4259
rect 1288 4227 1290 4259
rect 1424 4227 1426 4259
rect 1560 4227 1562 4259
rect 1696 4227 1698 4259
rect 1934 4258 1940 4259
rect 1975 4262 1979 4263
rect 1936 4227 1938 4258
rect 1975 4257 1979 4258
rect 1995 4262 1999 4263
rect 1995 4257 1999 4258
rect 2171 4262 2175 4263
rect 2171 4257 2175 4258
rect 2243 4262 2247 4263
rect 2243 4257 2247 4258
rect 2371 4262 2375 4263
rect 2371 4257 2375 4258
rect 2507 4262 2511 4263
rect 2507 4257 2511 4258
rect 2563 4262 2567 4263
rect 2563 4257 2567 4258
rect 2747 4262 2751 4263
rect 2747 4257 2751 4258
rect 2763 4262 2767 4263
rect 2763 4257 2767 4258
rect 2923 4262 2927 4263
rect 2923 4257 2927 4258
rect 3019 4262 3023 4263
rect 3019 4257 3023 4258
rect 3107 4262 3111 4263
rect 3107 4257 3111 4258
rect 3283 4262 3287 4263
rect 3283 4257 3287 4258
rect 3291 4262 3295 4263
rect 3291 4257 3295 4258
rect 3799 4262 3803 4263
rect 3799 4257 3803 4258
rect 111 4226 115 4227
rect 111 4221 115 4222
rect 727 4226 731 4227
rect 727 4221 731 4222
rect 743 4226 747 4227
rect 743 4221 747 4222
rect 863 4226 867 4227
rect 863 4221 867 4222
rect 879 4226 883 4227
rect 879 4221 883 4222
rect 999 4226 1003 4227
rect 999 4221 1003 4222
rect 1015 4226 1019 4227
rect 1015 4221 1019 4222
rect 1135 4226 1139 4227
rect 1135 4221 1139 4222
rect 1151 4226 1155 4227
rect 1151 4221 1155 4222
rect 1271 4226 1275 4227
rect 1271 4221 1275 4222
rect 1287 4226 1291 4227
rect 1287 4221 1291 4222
rect 1407 4226 1411 4227
rect 1407 4221 1411 4222
rect 1423 4226 1427 4227
rect 1423 4221 1427 4222
rect 1543 4226 1547 4227
rect 1543 4221 1547 4222
rect 1559 4226 1563 4227
rect 1559 4221 1563 4222
rect 1679 4226 1683 4227
rect 1679 4221 1683 4222
rect 1695 4226 1699 4227
rect 1695 4221 1699 4222
rect 1815 4226 1819 4227
rect 1815 4221 1819 4222
rect 1935 4226 1939 4227
rect 1935 4221 1939 4222
rect 112 4198 114 4221
rect 110 4197 116 4198
rect 728 4197 730 4221
rect 864 4197 866 4221
rect 1000 4197 1002 4221
rect 1136 4197 1138 4221
rect 1272 4197 1274 4221
rect 1408 4197 1410 4221
rect 1544 4197 1546 4221
rect 1680 4197 1682 4221
rect 1816 4197 1818 4221
rect 1936 4198 1938 4221
rect 1934 4197 1940 4198
rect 1976 4197 1978 4257
rect 110 4193 111 4197
rect 115 4193 116 4197
rect 110 4192 116 4193
rect 726 4196 732 4197
rect 726 4192 727 4196
rect 731 4192 732 4196
rect 726 4191 732 4192
rect 862 4196 868 4197
rect 862 4192 863 4196
rect 867 4192 868 4196
rect 862 4191 868 4192
rect 998 4196 1004 4197
rect 998 4192 999 4196
rect 1003 4192 1004 4196
rect 998 4191 1004 4192
rect 1134 4196 1140 4197
rect 1134 4192 1135 4196
rect 1139 4192 1140 4196
rect 1134 4191 1140 4192
rect 1270 4196 1276 4197
rect 1270 4192 1271 4196
rect 1275 4192 1276 4196
rect 1270 4191 1276 4192
rect 1406 4196 1412 4197
rect 1406 4192 1407 4196
rect 1411 4192 1412 4196
rect 1406 4191 1412 4192
rect 1542 4196 1548 4197
rect 1542 4192 1543 4196
rect 1547 4192 1548 4196
rect 1542 4191 1548 4192
rect 1678 4196 1684 4197
rect 1678 4192 1679 4196
rect 1683 4192 1684 4196
rect 1678 4191 1684 4192
rect 1814 4196 1820 4197
rect 1814 4192 1815 4196
rect 1819 4192 1820 4196
rect 1934 4193 1935 4197
rect 1939 4193 1940 4197
rect 1934 4192 1940 4193
rect 1974 4196 1980 4197
rect 1996 4196 1998 4257
rect 2244 4196 2246 4257
rect 2508 4196 2510 4257
rect 2764 4196 2766 4257
rect 3020 4196 3022 4257
rect 3284 4196 3286 4257
rect 3800 4197 3802 4257
rect 3840 4211 3842 4283
rect 4108 4211 4110 4284
rect 4244 4211 4246 4284
rect 4380 4211 4382 4284
rect 4516 4211 4518 4284
rect 4652 4211 4654 4284
rect 5662 4283 5668 4284
rect 5664 4211 5666 4283
rect 3839 4210 3843 4211
rect 3839 4205 3843 4206
rect 3971 4210 3975 4211
rect 3971 4205 3975 4206
rect 4107 4210 4111 4211
rect 4107 4205 4111 4206
rect 4243 4210 4247 4211
rect 4243 4205 4247 4206
rect 4379 4210 4383 4211
rect 4379 4205 4383 4206
rect 4515 4210 4519 4211
rect 4515 4205 4519 4206
rect 4651 4210 4655 4211
rect 4651 4205 4655 4206
rect 5663 4210 5667 4211
rect 5663 4205 5667 4206
rect 3798 4196 3804 4197
rect 1974 4192 1975 4196
rect 1979 4192 1980 4196
rect 1814 4191 1820 4192
rect 1974 4191 1980 4192
rect 1994 4195 2000 4196
rect 1994 4191 1995 4195
rect 1999 4191 2000 4195
rect 1994 4190 2000 4191
rect 2242 4195 2248 4196
rect 2242 4191 2243 4195
rect 2247 4191 2248 4195
rect 2242 4190 2248 4191
rect 2506 4195 2512 4196
rect 2506 4191 2507 4195
rect 2511 4191 2512 4195
rect 2506 4190 2512 4191
rect 2762 4195 2768 4196
rect 2762 4191 2763 4195
rect 2767 4191 2768 4195
rect 2762 4190 2768 4191
rect 3018 4195 3024 4196
rect 3018 4191 3019 4195
rect 3023 4191 3024 4195
rect 3018 4190 3024 4191
rect 3282 4195 3288 4196
rect 3282 4191 3283 4195
rect 3287 4191 3288 4195
rect 3798 4192 3799 4196
rect 3803 4192 3804 4196
rect 3798 4191 3804 4192
rect 3282 4190 3288 4191
rect 698 4181 704 4182
rect 110 4180 116 4181
rect 110 4176 111 4180
rect 115 4176 116 4180
rect 698 4177 699 4181
rect 703 4177 704 4181
rect 698 4176 704 4177
rect 834 4181 840 4182
rect 834 4177 835 4181
rect 839 4177 840 4181
rect 834 4176 840 4177
rect 970 4181 976 4182
rect 970 4177 971 4181
rect 975 4177 976 4181
rect 970 4176 976 4177
rect 1106 4181 1112 4182
rect 1106 4177 1107 4181
rect 1111 4177 1112 4181
rect 1106 4176 1112 4177
rect 1242 4181 1248 4182
rect 1242 4177 1243 4181
rect 1247 4177 1248 4181
rect 1242 4176 1248 4177
rect 1378 4181 1384 4182
rect 1378 4177 1379 4181
rect 1383 4177 1384 4181
rect 1378 4176 1384 4177
rect 1514 4181 1520 4182
rect 1514 4177 1515 4181
rect 1519 4177 1520 4181
rect 1514 4176 1520 4177
rect 1650 4181 1656 4182
rect 1650 4177 1651 4181
rect 1655 4177 1656 4181
rect 1650 4176 1656 4177
rect 1786 4181 1792 4182
rect 1786 4177 1787 4181
rect 1791 4177 1792 4181
rect 1786 4176 1792 4177
rect 1934 4180 1940 4181
rect 2022 4180 2028 4181
rect 1934 4176 1935 4180
rect 1939 4176 1940 4180
rect 110 4175 116 4176
rect 112 4115 114 4175
rect 700 4115 702 4176
rect 836 4115 838 4176
rect 972 4115 974 4176
rect 1108 4115 1110 4176
rect 1244 4115 1246 4176
rect 1380 4115 1382 4176
rect 1516 4115 1518 4176
rect 1652 4115 1654 4176
rect 1788 4115 1790 4176
rect 1934 4175 1940 4176
rect 1974 4179 1980 4180
rect 1974 4175 1975 4179
rect 1979 4175 1980 4179
rect 2022 4176 2023 4180
rect 2027 4176 2028 4180
rect 2022 4175 2028 4176
rect 2270 4180 2276 4181
rect 2270 4176 2271 4180
rect 2275 4176 2276 4180
rect 2270 4175 2276 4176
rect 2534 4180 2540 4181
rect 2534 4176 2535 4180
rect 2539 4176 2540 4180
rect 2534 4175 2540 4176
rect 2790 4180 2796 4181
rect 2790 4176 2791 4180
rect 2795 4176 2796 4180
rect 2790 4175 2796 4176
rect 3046 4180 3052 4181
rect 3046 4176 3047 4180
rect 3051 4176 3052 4180
rect 3046 4175 3052 4176
rect 3310 4180 3316 4181
rect 3310 4176 3311 4180
rect 3315 4176 3316 4180
rect 3310 4175 3316 4176
rect 3798 4179 3804 4180
rect 3798 4175 3799 4179
rect 3803 4175 3804 4179
rect 1936 4115 1938 4175
rect 1974 4174 1980 4175
rect 1976 4139 1978 4174
rect 2024 4139 2026 4175
rect 2272 4139 2274 4175
rect 2536 4139 2538 4175
rect 2792 4139 2794 4175
rect 3048 4139 3050 4175
rect 3312 4139 3314 4175
rect 3798 4174 3804 4175
rect 3800 4139 3802 4174
rect 3840 4145 3842 4205
rect 3838 4144 3844 4145
rect 3972 4144 3974 4205
rect 4108 4144 4110 4205
rect 4244 4144 4246 4205
rect 4380 4144 4382 4205
rect 4516 4144 4518 4205
rect 5664 4145 5666 4205
rect 5662 4144 5668 4145
rect 3838 4140 3839 4144
rect 3843 4140 3844 4144
rect 3838 4139 3844 4140
rect 3970 4143 3976 4144
rect 3970 4139 3971 4143
rect 3975 4139 3976 4143
rect 1975 4138 1979 4139
rect 1975 4133 1979 4134
rect 2023 4138 2027 4139
rect 2023 4133 2027 4134
rect 2271 4138 2275 4139
rect 2271 4133 2275 4134
rect 2535 4138 2539 4139
rect 2535 4133 2539 4134
rect 2791 4138 2795 4139
rect 2791 4133 2795 4134
rect 3047 4138 3051 4139
rect 3047 4133 3051 4134
rect 3135 4138 3139 4139
rect 3135 4133 3139 4134
rect 3271 4138 3275 4139
rect 3271 4133 3275 4134
rect 3311 4138 3315 4139
rect 3311 4133 3315 4134
rect 3407 4138 3411 4139
rect 3407 4133 3411 4134
rect 3543 4138 3547 4139
rect 3543 4133 3547 4134
rect 3679 4138 3683 4139
rect 3679 4133 3683 4134
rect 3799 4138 3803 4139
rect 3970 4138 3976 4139
rect 4106 4143 4112 4144
rect 4106 4139 4107 4143
rect 4111 4139 4112 4143
rect 4106 4138 4112 4139
rect 4242 4143 4248 4144
rect 4242 4139 4243 4143
rect 4247 4139 4248 4143
rect 4242 4138 4248 4139
rect 4378 4143 4384 4144
rect 4378 4139 4379 4143
rect 4383 4139 4384 4143
rect 4378 4138 4384 4139
rect 4514 4143 4520 4144
rect 4514 4139 4515 4143
rect 4519 4139 4520 4143
rect 5662 4140 5663 4144
rect 5667 4140 5668 4144
rect 5662 4139 5668 4140
rect 4514 4138 4520 4139
rect 3799 4133 3803 4134
rect 111 4114 115 4115
rect 111 4109 115 4110
rect 563 4114 567 4115
rect 563 4109 567 4110
rect 699 4114 703 4115
rect 699 4109 703 4110
rect 835 4114 839 4115
rect 835 4109 839 4110
rect 971 4114 975 4115
rect 971 4109 975 4110
rect 1107 4114 1111 4115
rect 1107 4109 1111 4110
rect 1243 4114 1247 4115
rect 1243 4109 1247 4110
rect 1379 4114 1383 4115
rect 1379 4109 1383 4110
rect 1515 4114 1519 4115
rect 1515 4109 1519 4110
rect 1651 4114 1655 4115
rect 1651 4109 1655 4110
rect 1787 4114 1791 4115
rect 1787 4109 1791 4110
rect 1935 4114 1939 4115
rect 1976 4110 1978 4133
rect 1935 4109 1939 4110
rect 1974 4109 1980 4110
rect 3136 4109 3138 4133
rect 3272 4109 3274 4133
rect 3408 4109 3410 4133
rect 3544 4109 3546 4133
rect 3680 4109 3682 4133
rect 3800 4110 3802 4133
rect 3998 4128 4004 4129
rect 3838 4127 3844 4128
rect 3838 4123 3839 4127
rect 3843 4123 3844 4127
rect 3998 4124 3999 4128
rect 4003 4124 4004 4128
rect 3998 4123 4004 4124
rect 4134 4128 4140 4129
rect 4134 4124 4135 4128
rect 4139 4124 4140 4128
rect 4134 4123 4140 4124
rect 4270 4128 4276 4129
rect 4270 4124 4271 4128
rect 4275 4124 4276 4128
rect 4270 4123 4276 4124
rect 4406 4128 4412 4129
rect 4406 4124 4407 4128
rect 4411 4124 4412 4128
rect 4406 4123 4412 4124
rect 4542 4128 4548 4129
rect 4542 4124 4543 4128
rect 4547 4124 4548 4128
rect 4542 4123 4548 4124
rect 5662 4127 5668 4128
rect 5662 4123 5663 4127
rect 5667 4123 5668 4127
rect 3838 4122 3844 4123
rect 3798 4109 3804 4110
rect 112 4049 114 4109
rect 110 4048 116 4049
rect 564 4048 566 4109
rect 700 4048 702 4109
rect 836 4048 838 4109
rect 972 4048 974 4109
rect 1108 4048 1110 4109
rect 1244 4048 1246 4109
rect 1380 4048 1382 4109
rect 1516 4048 1518 4109
rect 1652 4048 1654 4109
rect 1788 4048 1790 4109
rect 1936 4049 1938 4109
rect 1974 4105 1975 4109
rect 1979 4105 1980 4109
rect 1974 4104 1980 4105
rect 3134 4108 3140 4109
rect 3134 4104 3135 4108
rect 3139 4104 3140 4108
rect 3134 4103 3140 4104
rect 3270 4108 3276 4109
rect 3270 4104 3271 4108
rect 3275 4104 3276 4108
rect 3270 4103 3276 4104
rect 3406 4108 3412 4109
rect 3406 4104 3407 4108
rect 3411 4104 3412 4108
rect 3406 4103 3412 4104
rect 3542 4108 3548 4109
rect 3542 4104 3543 4108
rect 3547 4104 3548 4108
rect 3542 4103 3548 4104
rect 3678 4108 3684 4109
rect 3678 4104 3679 4108
rect 3683 4104 3684 4108
rect 3798 4105 3799 4109
rect 3803 4105 3804 4109
rect 3798 4104 3804 4105
rect 3678 4103 3684 4104
rect 3106 4093 3112 4094
rect 1974 4092 1980 4093
rect 1974 4088 1975 4092
rect 1979 4088 1980 4092
rect 3106 4089 3107 4093
rect 3111 4089 3112 4093
rect 3106 4088 3112 4089
rect 3242 4093 3248 4094
rect 3242 4089 3243 4093
rect 3247 4089 3248 4093
rect 3242 4088 3248 4089
rect 3378 4093 3384 4094
rect 3378 4089 3379 4093
rect 3383 4089 3384 4093
rect 3378 4088 3384 4089
rect 3514 4093 3520 4094
rect 3514 4089 3515 4093
rect 3519 4089 3520 4093
rect 3514 4088 3520 4089
rect 3650 4093 3656 4094
rect 3650 4089 3651 4093
rect 3655 4089 3656 4093
rect 3650 4088 3656 4089
rect 3798 4092 3804 4093
rect 3798 4088 3799 4092
rect 3803 4088 3804 4092
rect 1974 4087 1980 4088
rect 1934 4048 1940 4049
rect 110 4044 111 4048
rect 115 4044 116 4048
rect 110 4043 116 4044
rect 562 4047 568 4048
rect 562 4043 563 4047
rect 567 4043 568 4047
rect 562 4042 568 4043
rect 698 4047 704 4048
rect 698 4043 699 4047
rect 703 4043 704 4047
rect 698 4042 704 4043
rect 834 4047 840 4048
rect 834 4043 835 4047
rect 839 4043 840 4047
rect 834 4042 840 4043
rect 970 4047 976 4048
rect 970 4043 971 4047
rect 975 4043 976 4047
rect 970 4042 976 4043
rect 1106 4047 1112 4048
rect 1106 4043 1107 4047
rect 1111 4043 1112 4047
rect 1106 4042 1112 4043
rect 1242 4047 1248 4048
rect 1242 4043 1243 4047
rect 1247 4043 1248 4047
rect 1242 4042 1248 4043
rect 1378 4047 1384 4048
rect 1378 4043 1379 4047
rect 1383 4043 1384 4047
rect 1378 4042 1384 4043
rect 1514 4047 1520 4048
rect 1514 4043 1515 4047
rect 1519 4043 1520 4047
rect 1514 4042 1520 4043
rect 1650 4047 1656 4048
rect 1650 4043 1651 4047
rect 1655 4043 1656 4047
rect 1650 4042 1656 4043
rect 1786 4047 1792 4048
rect 1786 4043 1787 4047
rect 1791 4043 1792 4047
rect 1934 4044 1935 4048
rect 1939 4044 1940 4048
rect 1934 4043 1940 4044
rect 1786 4042 1792 4043
rect 590 4032 596 4033
rect 110 4031 116 4032
rect 110 4027 111 4031
rect 115 4027 116 4031
rect 590 4028 591 4032
rect 595 4028 596 4032
rect 590 4027 596 4028
rect 726 4032 732 4033
rect 726 4028 727 4032
rect 731 4028 732 4032
rect 726 4027 732 4028
rect 862 4032 868 4033
rect 862 4028 863 4032
rect 867 4028 868 4032
rect 862 4027 868 4028
rect 998 4032 1004 4033
rect 998 4028 999 4032
rect 1003 4028 1004 4032
rect 998 4027 1004 4028
rect 1134 4032 1140 4033
rect 1134 4028 1135 4032
rect 1139 4028 1140 4032
rect 1134 4027 1140 4028
rect 1270 4032 1276 4033
rect 1270 4028 1271 4032
rect 1275 4028 1276 4032
rect 1270 4027 1276 4028
rect 1406 4032 1412 4033
rect 1406 4028 1407 4032
rect 1411 4028 1412 4032
rect 1406 4027 1412 4028
rect 1542 4032 1548 4033
rect 1542 4028 1543 4032
rect 1547 4028 1548 4032
rect 1542 4027 1548 4028
rect 1678 4032 1684 4033
rect 1678 4028 1679 4032
rect 1683 4028 1684 4032
rect 1678 4027 1684 4028
rect 1814 4032 1820 4033
rect 1814 4028 1815 4032
rect 1819 4028 1820 4032
rect 1814 4027 1820 4028
rect 1934 4031 1940 4032
rect 1934 4027 1935 4031
rect 1939 4027 1940 4031
rect 110 4026 116 4027
rect 112 4003 114 4026
rect 592 4003 594 4027
rect 728 4003 730 4027
rect 864 4003 866 4027
rect 1000 4003 1002 4027
rect 1136 4003 1138 4027
rect 1272 4003 1274 4027
rect 1408 4003 1410 4027
rect 1544 4003 1546 4027
rect 1680 4003 1682 4027
rect 1816 4003 1818 4027
rect 1934 4026 1940 4027
rect 1936 4003 1938 4026
rect 111 4002 115 4003
rect 111 3997 115 3998
rect 159 4002 163 4003
rect 159 3997 163 3998
rect 327 4002 331 4003
rect 327 3997 331 3998
rect 535 4002 539 4003
rect 535 3997 539 3998
rect 591 4002 595 4003
rect 591 3997 595 3998
rect 727 4002 731 4003
rect 727 3997 731 3998
rect 751 4002 755 4003
rect 751 3997 755 3998
rect 863 4002 867 4003
rect 863 3997 867 3998
rect 967 4002 971 4003
rect 967 3997 971 3998
rect 999 4002 1003 4003
rect 999 3997 1003 3998
rect 1135 4002 1139 4003
rect 1135 3997 1139 3998
rect 1183 4002 1187 4003
rect 1183 3997 1187 3998
rect 1271 4002 1275 4003
rect 1271 3997 1275 3998
rect 1399 4002 1403 4003
rect 1399 3997 1403 3998
rect 1407 4002 1411 4003
rect 1407 3997 1411 3998
rect 1543 4002 1547 4003
rect 1543 3997 1547 3998
rect 1615 4002 1619 4003
rect 1615 3997 1619 3998
rect 1679 4002 1683 4003
rect 1679 3997 1683 3998
rect 1815 4002 1819 4003
rect 1815 3997 1819 3998
rect 1935 4002 1939 4003
rect 1935 3997 1939 3998
rect 112 3974 114 3997
rect 110 3973 116 3974
rect 160 3973 162 3997
rect 328 3973 330 3997
rect 536 3973 538 3997
rect 752 3973 754 3997
rect 968 3973 970 3997
rect 1184 3973 1186 3997
rect 1400 3973 1402 3997
rect 1616 3973 1618 3997
rect 1816 3973 1818 3997
rect 1936 3974 1938 3997
rect 1934 3973 1940 3974
rect 110 3969 111 3973
rect 115 3969 116 3973
rect 110 3968 116 3969
rect 158 3972 164 3973
rect 158 3968 159 3972
rect 163 3968 164 3972
rect 158 3967 164 3968
rect 326 3972 332 3973
rect 326 3968 327 3972
rect 331 3968 332 3972
rect 326 3967 332 3968
rect 534 3972 540 3973
rect 534 3968 535 3972
rect 539 3968 540 3972
rect 534 3967 540 3968
rect 750 3972 756 3973
rect 750 3968 751 3972
rect 755 3968 756 3972
rect 750 3967 756 3968
rect 966 3972 972 3973
rect 966 3968 967 3972
rect 971 3968 972 3972
rect 966 3967 972 3968
rect 1182 3972 1188 3973
rect 1182 3968 1183 3972
rect 1187 3968 1188 3972
rect 1182 3967 1188 3968
rect 1398 3972 1404 3973
rect 1398 3968 1399 3972
rect 1403 3968 1404 3972
rect 1398 3967 1404 3968
rect 1614 3972 1620 3973
rect 1614 3968 1615 3972
rect 1619 3968 1620 3972
rect 1614 3967 1620 3968
rect 1814 3972 1820 3973
rect 1814 3968 1815 3972
rect 1819 3968 1820 3972
rect 1934 3969 1935 3973
rect 1939 3969 1940 3973
rect 1934 3968 1940 3969
rect 1814 3967 1820 3968
rect 130 3957 136 3958
rect 110 3956 116 3957
rect 110 3952 111 3956
rect 115 3952 116 3956
rect 130 3953 131 3957
rect 135 3953 136 3957
rect 130 3952 136 3953
rect 298 3957 304 3958
rect 298 3953 299 3957
rect 303 3953 304 3957
rect 298 3952 304 3953
rect 506 3957 512 3958
rect 506 3953 507 3957
rect 511 3953 512 3957
rect 506 3952 512 3953
rect 722 3957 728 3958
rect 722 3953 723 3957
rect 727 3953 728 3957
rect 722 3952 728 3953
rect 938 3957 944 3958
rect 938 3953 939 3957
rect 943 3953 944 3957
rect 938 3952 944 3953
rect 1154 3957 1160 3958
rect 1154 3953 1155 3957
rect 1159 3953 1160 3957
rect 1154 3952 1160 3953
rect 1370 3957 1376 3958
rect 1370 3953 1371 3957
rect 1375 3953 1376 3957
rect 1370 3952 1376 3953
rect 1586 3957 1592 3958
rect 1586 3953 1587 3957
rect 1591 3953 1592 3957
rect 1586 3952 1592 3953
rect 1786 3957 1792 3958
rect 1786 3953 1787 3957
rect 1791 3953 1792 3957
rect 1786 3952 1792 3953
rect 1934 3956 1940 3957
rect 1934 3952 1935 3956
rect 1939 3952 1940 3956
rect 110 3951 116 3952
rect 112 3891 114 3951
rect 132 3891 134 3952
rect 300 3891 302 3952
rect 508 3891 510 3952
rect 724 3891 726 3952
rect 940 3891 942 3952
rect 1156 3891 1158 3952
rect 1372 3891 1374 3952
rect 1588 3891 1590 3952
rect 1788 3891 1790 3952
rect 1934 3951 1940 3952
rect 1936 3891 1938 3951
rect 1976 3935 1978 4087
rect 3108 3935 3110 4088
rect 3244 3935 3246 4088
rect 3380 3935 3382 4088
rect 3516 3935 3518 4088
rect 3652 3935 3654 4088
rect 3798 4087 3804 4088
rect 3800 3935 3802 4087
rect 3840 4075 3842 4122
rect 4000 4075 4002 4123
rect 4136 4075 4138 4123
rect 4272 4075 4274 4123
rect 4408 4075 4410 4123
rect 4544 4075 4546 4123
rect 5662 4122 5668 4123
rect 5664 4075 5666 4122
rect 3839 4074 3843 4075
rect 3839 4069 3843 4070
rect 3887 4074 3891 4075
rect 3887 4069 3891 4070
rect 3999 4074 4003 4075
rect 3999 4069 4003 4070
rect 4023 4074 4027 4075
rect 4023 4069 4027 4070
rect 4135 4074 4139 4075
rect 4135 4069 4139 4070
rect 4159 4074 4163 4075
rect 4159 4069 4163 4070
rect 4271 4074 4275 4075
rect 4271 4069 4275 4070
rect 4295 4074 4299 4075
rect 4295 4069 4299 4070
rect 4407 4074 4411 4075
rect 4407 4069 4411 4070
rect 4431 4074 4435 4075
rect 4431 4069 4435 4070
rect 4543 4074 4547 4075
rect 4543 4069 4547 4070
rect 4567 4074 4571 4075
rect 4567 4069 4571 4070
rect 4703 4074 4707 4075
rect 4703 4069 4707 4070
rect 4839 4074 4843 4075
rect 4839 4069 4843 4070
rect 5663 4074 5667 4075
rect 5663 4069 5667 4070
rect 3840 4046 3842 4069
rect 3838 4045 3844 4046
rect 3888 4045 3890 4069
rect 4024 4045 4026 4069
rect 4160 4045 4162 4069
rect 4296 4045 4298 4069
rect 4432 4045 4434 4069
rect 4568 4045 4570 4069
rect 4704 4045 4706 4069
rect 4840 4045 4842 4069
rect 5664 4046 5666 4069
rect 5662 4045 5668 4046
rect 3838 4041 3839 4045
rect 3843 4041 3844 4045
rect 3838 4040 3844 4041
rect 3886 4044 3892 4045
rect 3886 4040 3887 4044
rect 3891 4040 3892 4044
rect 3886 4039 3892 4040
rect 4022 4044 4028 4045
rect 4022 4040 4023 4044
rect 4027 4040 4028 4044
rect 4022 4039 4028 4040
rect 4158 4044 4164 4045
rect 4158 4040 4159 4044
rect 4163 4040 4164 4044
rect 4158 4039 4164 4040
rect 4294 4044 4300 4045
rect 4294 4040 4295 4044
rect 4299 4040 4300 4044
rect 4294 4039 4300 4040
rect 4430 4044 4436 4045
rect 4430 4040 4431 4044
rect 4435 4040 4436 4044
rect 4430 4039 4436 4040
rect 4566 4044 4572 4045
rect 4566 4040 4567 4044
rect 4571 4040 4572 4044
rect 4566 4039 4572 4040
rect 4702 4044 4708 4045
rect 4702 4040 4703 4044
rect 4707 4040 4708 4044
rect 4702 4039 4708 4040
rect 4838 4044 4844 4045
rect 4838 4040 4839 4044
rect 4843 4040 4844 4044
rect 5662 4041 5663 4045
rect 5667 4041 5668 4045
rect 5662 4040 5668 4041
rect 4838 4039 4844 4040
rect 3858 4029 3864 4030
rect 3838 4028 3844 4029
rect 3838 4024 3839 4028
rect 3843 4024 3844 4028
rect 3858 4025 3859 4029
rect 3863 4025 3864 4029
rect 3858 4024 3864 4025
rect 3994 4029 4000 4030
rect 3994 4025 3995 4029
rect 3999 4025 4000 4029
rect 3994 4024 4000 4025
rect 4130 4029 4136 4030
rect 4130 4025 4131 4029
rect 4135 4025 4136 4029
rect 4130 4024 4136 4025
rect 4266 4029 4272 4030
rect 4266 4025 4267 4029
rect 4271 4025 4272 4029
rect 4266 4024 4272 4025
rect 4402 4029 4408 4030
rect 4402 4025 4403 4029
rect 4407 4025 4408 4029
rect 4402 4024 4408 4025
rect 4538 4029 4544 4030
rect 4538 4025 4539 4029
rect 4543 4025 4544 4029
rect 4538 4024 4544 4025
rect 4674 4029 4680 4030
rect 4674 4025 4675 4029
rect 4679 4025 4680 4029
rect 4674 4024 4680 4025
rect 4810 4029 4816 4030
rect 4810 4025 4811 4029
rect 4815 4025 4816 4029
rect 4810 4024 4816 4025
rect 5662 4028 5668 4029
rect 5662 4024 5663 4028
rect 5667 4024 5668 4028
rect 3838 4023 3844 4024
rect 3840 3963 3842 4023
rect 3860 3963 3862 4024
rect 3996 3963 3998 4024
rect 4132 3963 4134 4024
rect 4268 3963 4270 4024
rect 4404 3963 4406 4024
rect 4540 3963 4542 4024
rect 4676 3963 4678 4024
rect 4812 3963 4814 4024
rect 5662 4023 5668 4024
rect 5664 3963 5666 4023
rect 3839 3962 3843 3963
rect 3839 3957 3843 3958
rect 3859 3962 3863 3963
rect 3859 3957 3863 3958
rect 3995 3962 3999 3963
rect 3995 3957 3999 3958
rect 4131 3962 4135 3963
rect 4131 3957 4135 3958
rect 4147 3962 4151 3963
rect 4147 3957 4151 3958
rect 4267 3962 4271 3963
rect 4267 3957 4271 3958
rect 4299 3962 4303 3963
rect 4299 3957 4303 3958
rect 4403 3962 4407 3963
rect 4403 3957 4407 3958
rect 4459 3962 4463 3963
rect 4459 3957 4463 3958
rect 4539 3962 4543 3963
rect 4539 3957 4543 3958
rect 4619 3962 4623 3963
rect 4619 3957 4623 3958
rect 4675 3962 4679 3963
rect 4675 3957 4679 3958
rect 4779 3962 4783 3963
rect 4779 3957 4783 3958
rect 4811 3962 4815 3963
rect 4811 3957 4815 3958
rect 5663 3962 5667 3963
rect 5663 3957 5667 3958
rect 1975 3934 1979 3935
rect 1975 3929 1979 3930
rect 1995 3934 1999 3935
rect 1995 3929 1999 3930
rect 2403 3934 2407 3935
rect 2403 3929 2407 3930
rect 2827 3934 2831 3935
rect 2827 3929 2831 3930
rect 3107 3934 3111 3935
rect 3107 3929 3111 3930
rect 3243 3934 3247 3935
rect 3243 3929 3247 3930
rect 3251 3934 3255 3935
rect 3251 3929 3255 3930
rect 3379 3934 3383 3935
rect 3379 3929 3383 3930
rect 3515 3934 3519 3935
rect 3515 3929 3519 3930
rect 3651 3934 3655 3935
rect 3651 3929 3655 3930
rect 3799 3934 3803 3935
rect 3799 3929 3803 3930
rect 111 3890 115 3891
rect 111 3885 115 3886
rect 131 3890 135 3891
rect 131 3885 135 3886
rect 299 3890 303 3891
rect 299 3885 303 3886
rect 355 3890 359 3891
rect 355 3885 359 3886
rect 507 3890 511 3891
rect 507 3885 511 3886
rect 619 3890 623 3891
rect 619 3885 623 3886
rect 723 3890 727 3891
rect 723 3885 727 3886
rect 899 3890 903 3891
rect 899 3885 903 3886
rect 939 3890 943 3891
rect 939 3885 943 3886
rect 1155 3890 1159 3891
rect 1155 3885 1159 3886
rect 1195 3890 1199 3891
rect 1195 3885 1199 3886
rect 1371 3890 1375 3891
rect 1371 3885 1375 3886
rect 1499 3890 1503 3891
rect 1499 3885 1503 3886
rect 1587 3890 1591 3891
rect 1587 3885 1591 3886
rect 1787 3890 1791 3891
rect 1787 3885 1791 3886
rect 1935 3890 1939 3891
rect 1935 3885 1939 3886
rect 112 3825 114 3885
rect 110 3824 116 3825
rect 132 3824 134 3885
rect 356 3824 358 3885
rect 620 3824 622 3885
rect 900 3824 902 3885
rect 1196 3824 1198 3885
rect 1500 3824 1502 3885
rect 1788 3824 1790 3885
rect 1936 3825 1938 3885
rect 1976 3869 1978 3929
rect 1974 3868 1980 3869
rect 1996 3868 1998 3929
rect 2404 3868 2406 3929
rect 2828 3868 2830 3929
rect 3252 3868 3254 3929
rect 3652 3868 3654 3929
rect 3800 3869 3802 3929
rect 3840 3897 3842 3957
rect 3838 3896 3844 3897
rect 3860 3896 3862 3957
rect 3996 3896 3998 3957
rect 4148 3896 4150 3957
rect 4300 3896 4302 3957
rect 4460 3896 4462 3957
rect 4620 3896 4622 3957
rect 4780 3896 4782 3957
rect 5664 3897 5666 3957
rect 5662 3896 5668 3897
rect 3838 3892 3839 3896
rect 3843 3892 3844 3896
rect 3838 3891 3844 3892
rect 3858 3895 3864 3896
rect 3858 3891 3859 3895
rect 3863 3891 3864 3895
rect 3858 3890 3864 3891
rect 3994 3895 4000 3896
rect 3994 3891 3995 3895
rect 3999 3891 4000 3895
rect 3994 3890 4000 3891
rect 4146 3895 4152 3896
rect 4146 3891 4147 3895
rect 4151 3891 4152 3895
rect 4146 3890 4152 3891
rect 4298 3895 4304 3896
rect 4298 3891 4299 3895
rect 4303 3891 4304 3895
rect 4298 3890 4304 3891
rect 4458 3895 4464 3896
rect 4458 3891 4459 3895
rect 4463 3891 4464 3895
rect 4458 3890 4464 3891
rect 4618 3895 4624 3896
rect 4618 3891 4619 3895
rect 4623 3891 4624 3895
rect 4618 3890 4624 3891
rect 4778 3895 4784 3896
rect 4778 3891 4779 3895
rect 4783 3891 4784 3895
rect 5662 3892 5663 3896
rect 5667 3892 5668 3896
rect 5662 3891 5668 3892
rect 4778 3890 4784 3891
rect 3886 3880 3892 3881
rect 3838 3879 3844 3880
rect 3838 3875 3839 3879
rect 3843 3875 3844 3879
rect 3886 3876 3887 3880
rect 3891 3876 3892 3880
rect 3886 3875 3892 3876
rect 4022 3880 4028 3881
rect 4022 3876 4023 3880
rect 4027 3876 4028 3880
rect 4022 3875 4028 3876
rect 4174 3880 4180 3881
rect 4174 3876 4175 3880
rect 4179 3876 4180 3880
rect 4174 3875 4180 3876
rect 4326 3880 4332 3881
rect 4326 3876 4327 3880
rect 4331 3876 4332 3880
rect 4326 3875 4332 3876
rect 4486 3880 4492 3881
rect 4486 3876 4487 3880
rect 4491 3876 4492 3880
rect 4486 3875 4492 3876
rect 4646 3880 4652 3881
rect 4646 3876 4647 3880
rect 4651 3876 4652 3880
rect 4646 3875 4652 3876
rect 4806 3880 4812 3881
rect 4806 3876 4807 3880
rect 4811 3876 4812 3880
rect 4806 3875 4812 3876
rect 5662 3879 5668 3880
rect 5662 3875 5663 3879
rect 5667 3875 5668 3879
rect 3838 3874 3844 3875
rect 3798 3868 3804 3869
rect 1974 3864 1975 3868
rect 1979 3864 1980 3868
rect 1974 3863 1980 3864
rect 1994 3867 2000 3868
rect 1994 3863 1995 3867
rect 1999 3863 2000 3867
rect 1994 3862 2000 3863
rect 2402 3867 2408 3868
rect 2402 3863 2403 3867
rect 2407 3863 2408 3867
rect 2402 3862 2408 3863
rect 2826 3867 2832 3868
rect 2826 3863 2827 3867
rect 2831 3863 2832 3867
rect 2826 3862 2832 3863
rect 3250 3867 3256 3868
rect 3250 3863 3251 3867
rect 3255 3863 3256 3867
rect 3250 3862 3256 3863
rect 3650 3867 3656 3868
rect 3650 3863 3651 3867
rect 3655 3863 3656 3867
rect 3798 3864 3799 3868
rect 3803 3864 3804 3868
rect 3798 3863 3804 3864
rect 3650 3862 3656 3863
rect 2022 3852 2028 3853
rect 1974 3851 1980 3852
rect 1974 3847 1975 3851
rect 1979 3847 1980 3851
rect 2022 3848 2023 3852
rect 2027 3848 2028 3852
rect 2022 3847 2028 3848
rect 2430 3852 2436 3853
rect 2430 3848 2431 3852
rect 2435 3848 2436 3852
rect 2430 3847 2436 3848
rect 2854 3852 2860 3853
rect 2854 3848 2855 3852
rect 2859 3848 2860 3852
rect 2854 3847 2860 3848
rect 3278 3852 3284 3853
rect 3278 3848 3279 3852
rect 3283 3848 3284 3852
rect 3278 3847 3284 3848
rect 3678 3852 3684 3853
rect 3678 3848 3679 3852
rect 3683 3848 3684 3852
rect 3678 3847 3684 3848
rect 3798 3851 3804 3852
rect 3798 3847 3799 3851
rect 3803 3847 3804 3851
rect 1974 3846 1980 3847
rect 1934 3824 1940 3825
rect 110 3820 111 3824
rect 115 3820 116 3824
rect 110 3819 116 3820
rect 130 3823 136 3824
rect 130 3819 131 3823
rect 135 3819 136 3823
rect 130 3818 136 3819
rect 354 3823 360 3824
rect 354 3819 355 3823
rect 359 3819 360 3823
rect 354 3818 360 3819
rect 618 3823 624 3824
rect 618 3819 619 3823
rect 623 3819 624 3823
rect 618 3818 624 3819
rect 898 3823 904 3824
rect 898 3819 899 3823
rect 903 3819 904 3823
rect 898 3818 904 3819
rect 1194 3823 1200 3824
rect 1194 3819 1195 3823
rect 1199 3819 1200 3823
rect 1194 3818 1200 3819
rect 1498 3823 1504 3824
rect 1498 3819 1499 3823
rect 1503 3819 1504 3823
rect 1498 3818 1504 3819
rect 1786 3823 1792 3824
rect 1786 3819 1787 3823
rect 1791 3819 1792 3823
rect 1934 3820 1935 3824
rect 1939 3820 1940 3824
rect 1976 3823 1978 3846
rect 2024 3823 2026 3847
rect 2432 3823 2434 3847
rect 2856 3823 2858 3847
rect 3280 3823 3282 3847
rect 3680 3823 3682 3847
rect 3798 3846 3804 3847
rect 3800 3823 3802 3846
rect 3840 3823 3842 3874
rect 3888 3823 3890 3875
rect 4024 3823 4026 3875
rect 4176 3823 4178 3875
rect 4328 3823 4330 3875
rect 4488 3823 4490 3875
rect 4648 3823 4650 3875
rect 4808 3823 4810 3875
rect 5662 3874 5668 3875
rect 5664 3823 5666 3874
rect 1934 3819 1940 3820
rect 1975 3822 1979 3823
rect 1786 3818 1792 3819
rect 1975 3817 1979 3818
rect 2023 3822 2027 3823
rect 2023 3817 2027 3818
rect 2175 3822 2179 3823
rect 2175 3817 2179 3818
rect 2351 3822 2355 3823
rect 2351 3817 2355 3818
rect 2431 3822 2435 3823
rect 2431 3817 2435 3818
rect 2535 3822 2539 3823
rect 2535 3817 2539 3818
rect 2719 3822 2723 3823
rect 2719 3817 2723 3818
rect 2855 3822 2859 3823
rect 2855 3817 2859 3818
rect 2895 3822 2899 3823
rect 2895 3817 2899 3818
rect 3071 3822 3075 3823
rect 3071 3817 3075 3818
rect 3247 3822 3251 3823
rect 3247 3817 3251 3818
rect 3279 3822 3283 3823
rect 3279 3817 3283 3818
rect 3423 3822 3427 3823
rect 3423 3817 3427 3818
rect 3607 3822 3611 3823
rect 3607 3817 3611 3818
rect 3679 3822 3683 3823
rect 3679 3817 3683 3818
rect 3799 3822 3803 3823
rect 3799 3817 3803 3818
rect 3839 3822 3843 3823
rect 3839 3817 3843 3818
rect 3887 3822 3891 3823
rect 3887 3817 3891 3818
rect 4023 3822 4027 3823
rect 4023 3817 4027 3818
rect 4175 3822 4179 3823
rect 4175 3817 4179 3818
rect 4327 3822 4331 3823
rect 4327 3817 4331 3818
rect 4487 3822 4491 3823
rect 4487 3817 4491 3818
rect 4503 3822 4507 3823
rect 4503 3817 4507 3818
rect 4639 3822 4643 3823
rect 4639 3817 4643 3818
rect 4647 3822 4651 3823
rect 4647 3817 4651 3818
rect 4775 3822 4779 3823
rect 4775 3817 4779 3818
rect 4807 3822 4811 3823
rect 4807 3817 4811 3818
rect 4911 3822 4915 3823
rect 4911 3817 4915 3818
rect 5047 3822 5051 3823
rect 5047 3817 5051 3818
rect 5663 3822 5667 3823
rect 5663 3817 5667 3818
rect 158 3808 164 3809
rect 110 3807 116 3808
rect 110 3803 111 3807
rect 115 3803 116 3807
rect 158 3804 159 3808
rect 163 3804 164 3808
rect 158 3803 164 3804
rect 382 3808 388 3809
rect 382 3804 383 3808
rect 387 3804 388 3808
rect 382 3803 388 3804
rect 646 3808 652 3809
rect 646 3804 647 3808
rect 651 3804 652 3808
rect 646 3803 652 3804
rect 926 3808 932 3809
rect 926 3804 927 3808
rect 931 3804 932 3808
rect 926 3803 932 3804
rect 1222 3808 1228 3809
rect 1222 3804 1223 3808
rect 1227 3804 1228 3808
rect 1222 3803 1228 3804
rect 1526 3808 1532 3809
rect 1526 3804 1527 3808
rect 1531 3804 1532 3808
rect 1526 3803 1532 3804
rect 1814 3808 1820 3809
rect 1814 3804 1815 3808
rect 1819 3804 1820 3808
rect 1814 3803 1820 3804
rect 1934 3807 1940 3808
rect 1934 3803 1935 3807
rect 1939 3803 1940 3807
rect 110 3802 116 3803
rect 112 3767 114 3802
rect 160 3767 162 3803
rect 384 3767 386 3803
rect 648 3767 650 3803
rect 928 3767 930 3803
rect 1224 3767 1226 3803
rect 1528 3767 1530 3803
rect 1816 3767 1818 3803
rect 1934 3802 1940 3803
rect 1936 3767 1938 3802
rect 1976 3794 1978 3817
rect 1974 3793 1980 3794
rect 2024 3793 2026 3817
rect 2176 3793 2178 3817
rect 2352 3793 2354 3817
rect 2536 3793 2538 3817
rect 2720 3793 2722 3817
rect 2896 3793 2898 3817
rect 3072 3793 3074 3817
rect 3248 3793 3250 3817
rect 3424 3793 3426 3817
rect 3608 3793 3610 3817
rect 3800 3794 3802 3817
rect 3840 3794 3842 3817
rect 3798 3793 3804 3794
rect 1974 3789 1975 3793
rect 1979 3789 1980 3793
rect 1974 3788 1980 3789
rect 2022 3792 2028 3793
rect 2022 3788 2023 3792
rect 2027 3788 2028 3792
rect 2022 3787 2028 3788
rect 2174 3792 2180 3793
rect 2174 3788 2175 3792
rect 2179 3788 2180 3792
rect 2174 3787 2180 3788
rect 2350 3792 2356 3793
rect 2350 3788 2351 3792
rect 2355 3788 2356 3792
rect 2350 3787 2356 3788
rect 2534 3792 2540 3793
rect 2534 3788 2535 3792
rect 2539 3788 2540 3792
rect 2534 3787 2540 3788
rect 2718 3792 2724 3793
rect 2718 3788 2719 3792
rect 2723 3788 2724 3792
rect 2718 3787 2724 3788
rect 2894 3792 2900 3793
rect 2894 3788 2895 3792
rect 2899 3788 2900 3792
rect 2894 3787 2900 3788
rect 3070 3792 3076 3793
rect 3070 3788 3071 3792
rect 3075 3788 3076 3792
rect 3070 3787 3076 3788
rect 3246 3792 3252 3793
rect 3246 3788 3247 3792
rect 3251 3788 3252 3792
rect 3246 3787 3252 3788
rect 3422 3792 3428 3793
rect 3422 3788 3423 3792
rect 3427 3788 3428 3792
rect 3422 3787 3428 3788
rect 3606 3792 3612 3793
rect 3606 3788 3607 3792
rect 3611 3788 3612 3792
rect 3798 3789 3799 3793
rect 3803 3789 3804 3793
rect 3798 3788 3804 3789
rect 3838 3793 3844 3794
rect 4504 3793 4506 3817
rect 4640 3793 4642 3817
rect 4776 3793 4778 3817
rect 4912 3793 4914 3817
rect 5048 3793 5050 3817
rect 5664 3794 5666 3817
rect 5662 3793 5668 3794
rect 3838 3789 3839 3793
rect 3843 3789 3844 3793
rect 3838 3788 3844 3789
rect 4502 3792 4508 3793
rect 4502 3788 4503 3792
rect 4507 3788 4508 3792
rect 3606 3787 3612 3788
rect 4502 3787 4508 3788
rect 4638 3792 4644 3793
rect 4638 3788 4639 3792
rect 4643 3788 4644 3792
rect 4638 3787 4644 3788
rect 4774 3792 4780 3793
rect 4774 3788 4775 3792
rect 4779 3788 4780 3792
rect 4774 3787 4780 3788
rect 4910 3792 4916 3793
rect 4910 3788 4911 3792
rect 4915 3788 4916 3792
rect 4910 3787 4916 3788
rect 5046 3792 5052 3793
rect 5046 3788 5047 3792
rect 5051 3788 5052 3792
rect 5662 3789 5663 3793
rect 5667 3789 5668 3793
rect 5662 3788 5668 3789
rect 5046 3787 5052 3788
rect 1994 3777 2000 3778
rect 1974 3776 1980 3777
rect 1974 3772 1975 3776
rect 1979 3772 1980 3776
rect 1994 3773 1995 3777
rect 1999 3773 2000 3777
rect 1994 3772 2000 3773
rect 2146 3777 2152 3778
rect 2146 3773 2147 3777
rect 2151 3773 2152 3777
rect 2146 3772 2152 3773
rect 2322 3777 2328 3778
rect 2322 3773 2323 3777
rect 2327 3773 2328 3777
rect 2322 3772 2328 3773
rect 2506 3777 2512 3778
rect 2506 3773 2507 3777
rect 2511 3773 2512 3777
rect 2506 3772 2512 3773
rect 2690 3777 2696 3778
rect 2690 3773 2691 3777
rect 2695 3773 2696 3777
rect 2690 3772 2696 3773
rect 2866 3777 2872 3778
rect 2866 3773 2867 3777
rect 2871 3773 2872 3777
rect 2866 3772 2872 3773
rect 3042 3777 3048 3778
rect 3042 3773 3043 3777
rect 3047 3773 3048 3777
rect 3042 3772 3048 3773
rect 3218 3777 3224 3778
rect 3218 3773 3219 3777
rect 3223 3773 3224 3777
rect 3218 3772 3224 3773
rect 3394 3777 3400 3778
rect 3394 3773 3395 3777
rect 3399 3773 3400 3777
rect 3394 3772 3400 3773
rect 3578 3777 3584 3778
rect 4474 3777 4480 3778
rect 3578 3773 3579 3777
rect 3583 3773 3584 3777
rect 3578 3772 3584 3773
rect 3798 3776 3804 3777
rect 3798 3772 3799 3776
rect 3803 3772 3804 3776
rect 1974 3771 1980 3772
rect 111 3766 115 3767
rect 111 3761 115 3762
rect 159 3766 163 3767
rect 159 3761 163 3762
rect 247 3766 251 3767
rect 247 3761 251 3762
rect 383 3766 387 3767
rect 383 3761 387 3762
rect 519 3766 523 3767
rect 519 3761 523 3762
rect 647 3766 651 3767
rect 647 3761 651 3762
rect 791 3766 795 3767
rect 791 3761 795 3762
rect 927 3766 931 3767
rect 927 3761 931 3762
rect 1063 3766 1067 3767
rect 1063 3761 1067 3762
rect 1223 3766 1227 3767
rect 1223 3761 1227 3762
rect 1343 3766 1347 3767
rect 1343 3761 1347 3762
rect 1527 3766 1531 3767
rect 1527 3761 1531 3762
rect 1815 3766 1819 3767
rect 1815 3761 1819 3762
rect 1935 3766 1939 3767
rect 1935 3761 1939 3762
rect 112 3738 114 3761
rect 110 3737 116 3738
rect 248 3737 250 3761
rect 520 3737 522 3761
rect 792 3737 794 3761
rect 1064 3737 1066 3761
rect 1344 3737 1346 3761
rect 1936 3738 1938 3761
rect 1934 3737 1940 3738
rect 110 3733 111 3737
rect 115 3733 116 3737
rect 110 3732 116 3733
rect 246 3736 252 3737
rect 246 3732 247 3736
rect 251 3732 252 3736
rect 246 3731 252 3732
rect 518 3736 524 3737
rect 518 3732 519 3736
rect 523 3732 524 3736
rect 518 3731 524 3732
rect 790 3736 796 3737
rect 790 3732 791 3736
rect 795 3732 796 3736
rect 790 3731 796 3732
rect 1062 3736 1068 3737
rect 1062 3732 1063 3736
rect 1067 3732 1068 3736
rect 1062 3731 1068 3732
rect 1342 3736 1348 3737
rect 1342 3732 1343 3736
rect 1347 3732 1348 3736
rect 1934 3733 1935 3737
rect 1939 3733 1940 3737
rect 1934 3732 1940 3733
rect 1342 3731 1348 3732
rect 218 3721 224 3722
rect 110 3720 116 3721
rect 110 3716 111 3720
rect 115 3716 116 3720
rect 218 3717 219 3721
rect 223 3717 224 3721
rect 218 3716 224 3717
rect 490 3721 496 3722
rect 490 3717 491 3721
rect 495 3717 496 3721
rect 490 3716 496 3717
rect 762 3721 768 3722
rect 762 3717 763 3721
rect 767 3717 768 3721
rect 762 3716 768 3717
rect 1034 3721 1040 3722
rect 1034 3717 1035 3721
rect 1039 3717 1040 3721
rect 1034 3716 1040 3717
rect 1314 3721 1320 3722
rect 1314 3717 1315 3721
rect 1319 3717 1320 3721
rect 1314 3716 1320 3717
rect 1934 3720 1940 3721
rect 1934 3716 1935 3720
rect 1939 3716 1940 3720
rect 110 3715 116 3716
rect 112 3639 114 3715
rect 220 3639 222 3716
rect 492 3639 494 3716
rect 764 3639 766 3716
rect 1036 3639 1038 3716
rect 1316 3639 1318 3716
rect 1934 3715 1940 3716
rect 1936 3639 1938 3715
rect 1976 3703 1978 3771
rect 1996 3703 1998 3772
rect 2148 3703 2150 3772
rect 2324 3703 2326 3772
rect 2508 3703 2510 3772
rect 2692 3703 2694 3772
rect 2868 3703 2870 3772
rect 3044 3703 3046 3772
rect 3220 3703 3222 3772
rect 3396 3703 3398 3772
rect 3580 3703 3582 3772
rect 3798 3771 3804 3772
rect 3838 3776 3844 3777
rect 3838 3772 3839 3776
rect 3843 3772 3844 3776
rect 4474 3773 4475 3777
rect 4479 3773 4480 3777
rect 4474 3772 4480 3773
rect 4610 3777 4616 3778
rect 4610 3773 4611 3777
rect 4615 3773 4616 3777
rect 4610 3772 4616 3773
rect 4746 3777 4752 3778
rect 4746 3773 4747 3777
rect 4751 3773 4752 3777
rect 4746 3772 4752 3773
rect 4882 3777 4888 3778
rect 4882 3773 4883 3777
rect 4887 3773 4888 3777
rect 4882 3772 4888 3773
rect 5018 3777 5024 3778
rect 5018 3773 5019 3777
rect 5023 3773 5024 3777
rect 5018 3772 5024 3773
rect 5662 3776 5668 3777
rect 5662 3772 5663 3776
rect 5667 3772 5668 3776
rect 3838 3771 3844 3772
rect 3800 3703 3802 3771
rect 1975 3702 1979 3703
rect 1975 3697 1979 3698
rect 1995 3702 1999 3703
rect 1995 3697 1999 3698
rect 2011 3702 2015 3703
rect 2011 3697 2015 3698
rect 2147 3702 2151 3703
rect 2147 3697 2151 3698
rect 2291 3702 2295 3703
rect 2291 3697 2295 3698
rect 2323 3702 2327 3703
rect 2323 3697 2327 3698
rect 2435 3702 2439 3703
rect 2435 3697 2439 3698
rect 2507 3702 2511 3703
rect 2507 3697 2511 3698
rect 2579 3702 2583 3703
rect 2579 3697 2583 3698
rect 2691 3702 2695 3703
rect 2691 3697 2695 3698
rect 2723 3702 2727 3703
rect 2723 3697 2727 3698
rect 2867 3702 2871 3703
rect 2867 3697 2871 3698
rect 3011 3702 3015 3703
rect 3011 3697 3015 3698
rect 3043 3702 3047 3703
rect 3043 3697 3047 3698
rect 3155 3702 3159 3703
rect 3155 3697 3159 3698
rect 3219 3702 3223 3703
rect 3219 3697 3223 3698
rect 3299 3702 3303 3703
rect 3299 3697 3303 3698
rect 3395 3702 3399 3703
rect 3395 3697 3399 3698
rect 3579 3702 3583 3703
rect 3579 3697 3583 3698
rect 3799 3702 3803 3703
rect 3799 3697 3803 3698
rect 111 3638 115 3639
rect 111 3633 115 3634
rect 219 3638 223 3639
rect 219 3633 223 3634
rect 491 3638 495 3639
rect 491 3633 495 3634
rect 635 3638 639 3639
rect 635 3633 639 3634
rect 763 3638 767 3639
rect 763 3633 767 3634
rect 779 3638 783 3639
rect 779 3633 783 3634
rect 923 3638 927 3639
rect 923 3633 927 3634
rect 1035 3638 1039 3639
rect 1035 3633 1039 3634
rect 1067 3638 1071 3639
rect 1067 3633 1071 3634
rect 1211 3638 1215 3639
rect 1211 3633 1215 3634
rect 1315 3638 1319 3639
rect 1315 3633 1319 3634
rect 1935 3638 1939 3639
rect 1976 3637 1978 3697
rect 1935 3633 1939 3634
rect 1974 3636 1980 3637
rect 2012 3636 2014 3697
rect 2148 3636 2150 3697
rect 2292 3636 2294 3697
rect 2436 3636 2438 3697
rect 2580 3636 2582 3697
rect 2724 3636 2726 3697
rect 2868 3636 2870 3697
rect 3012 3636 3014 3697
rect 3156 3636 3158 3697
rect 3300 3636 3302 3697
rect 3800 3637 3802 3697
rect 3840 3691 3842 3771
rect 4476 3691 4478 3772
rect 4612 3691 4614 3772
rect 4748 3691 4750 3772
rect 4884 3691 4886 3772
rect 5020 3691 5022 3772
rect 5662 3771 5668 3772
rect 5664 3691 5666 3771
rect 3839 3690 3843 3691
rect 3839 3685 3843 3686
rect 4019 3690 4023 3691
rect 4019 3685 4023 3686
rect 4155 3690 4159 3691
rect 4155 3685 4159 3686
rect 4291 3690 4295 3691
rect 4291 3685 4295 3686
rect 4427 3690 4431 3691
rect 4427 3685 4431 3686
rect 4475 3690 4479 3691
rect 4475 3685 4479 3686
rect 4563 3690 4567 3691
rect 4563 3685 4567 3686
rect 4611 3690 4615 3691
rect 4611 3685 4615 3686
rect 4699 3690 4703 3691
rect 4699 3685 4703 3686
rect 4747 3690 4751 3691
rect 4747 3685 4751 3686
rect 4835 3690 4839 3691
rect 4835 3685 4839 3686
rect 4883 3690 4887 3691
rect 4883 3685 4887 3686
rect 4971 3690 4975 3691
rect 4971 3685 4975 3686
rect 5019 3690 5023 3691
rect 5019 3685 5023 3686
rect 5107 3690 5111 3691
rect 5107 3685 5111 3686
rect 5243 3690 5247 3691
rect 5243 3685 5247 3686
rect 5379 3690 5383 3691
rect 5379 3685 5383 3686
rect 5515 3690 5519 3691
rect 5515 3685 5519 3686
rect 5663 3690 5667 3691
rect 5663 3685 5667 3686
rect 3798 3636 3804 3637
rect 112 3573 114 3633
rect 110 3572 116 3573
rect 492 3572 494 3633
rect 636 3572 638 3633
rect 780 3572 782 3633
rect 924 3572 926 3633
rect 1068 3572 1070 3633
rect 1212 3572 1214 3633
rect 1936 3573 1938 3633
rect 1974 3632 1975 3636
rect 1979 3632 1980 3636
rect 1974 3631 1980 3632
rect 2010 3635 2016 3636
rect 2010 3631 2011 3635
rect 2015 3631 2016 3635
rect 2010 3630 2016 3631
rect 2146 3635 2152 3636
rect 2146 3631 2147 3635
rect 2151 3631 2152 3635
rect 2146 3630 2152 3631
rect 2290 3635 2296 3636
rect 2290 3631 2291 3635
rect 2295 3631 2296 3635
rect 2290 3630 2296 3631
rect 2434 3635 2440 3636
rect 2434 3631 2435 3635
rect 2439 3631 2440 3635
rect 2434 3630 2440 3631
rect 2578 3635 2584 3636
rect 2578 3631 2579 3635
rect 2583 3631 2584 3635
rect 2578 3630 2584 3631
rect 2722 3635 2728 3636
rect 2722 3631 2723 3635
rect 2727 3631 2728 3635
rect 2722 3630 2728 3631
rect 2866 3635 2872 3636
rect 2866 3631 2867 3635
rect 2871 3631 2872 3635
rect 2866 3630 2872 3631
rect 3010 3635 3016 3636
rect 3010 3631 3011 3635
rect 3015 3631 3016 3635
rect 3010 3630 3016 3631
rect 3154 3635 3160 3636
rect 3154 3631 3155 3635
rect 3159 3631 3160 3635
rect 3154 3630 3160 3631
rect 3298 3635 3304 3636
rect 3298 3631 3299 3635
rect 3303 3631 3304 3635
rect 3798 3632 3799 3636
rect 3803 3632 3804 3636
rect 3798 3631 3804 3632
rect 3298 3630 3304 3631
rect 3840 3625 3842 3685
rect 3838 3624 3844 3625
rect 4020 3624 4022 3685
rect 4156 3624 4158 3685
rect 4292 3624 4294 3685
rect 4428 3624 4430 3685
rect 4564 3624 4566 3685
rect 4700 3624 4702 3685
rect 4836 3624 4838 3685
rect 4972 3624 4974 3685
rect 5108 3624 5110 3685
rect 5244 3624 5246 3685
rect 5380 3624 5382 3685
rect 5516 3624 5518 3685
rect 5664 3625 5666 3685
rect 5662 3624 5668 3625
rect 2038 3620 2044 3621
rect 1974 3619 1980 3620
rect 1974 3615 1975 3619
rect 1979 3615 1980 3619
rect 2038 3616 2039 3620
rect 2043 3616 2044 3620
rect 2038 3615 2044 3616
rect 2174 3620 2180 3621
rect 2174 3616 2175 3620
rect 2179 3616 2180 3620
rect 2174 3615 2180 3616
rect 2318 3620 2324 3621
rect 2318 3616 2319 3620
rect 2323 3616 2324 3620
rect 2318 3615 2324 3616
rect 2462 3620 2468 3621
rect 2462 3616 2463 3620
rect 2467 3616 2468 3620
rect 2462 3615 2468 3616
rect 2606 3620 2612 3621
rect 2606 3616 2607 3620
rect 2611 3616 2612 3620
rect 2606 3615 2612 3616
rect 2750 3620 2756 3621
rect 2750 3616 2751 3620
rect 2755 3616 2756 3620
rect 2750 3615 2756 3616
rect 2894 3620 2900 3621
rect 2894 3616 2895 3620
rect 2899 3616 2900 3620
rect 2894 3615 2900 3616
rect 3038 3620 3044 3621
rect 3038 3616 3039 3620
rect 3043 3616 3044 3620
rect 3038 3615 3044 3616
rect 3182 3620 3188 3621
rect 3182 3616 3183 3620
rect 3187 3616 3188 3620
rect 3182 3615 3188 3616
rect 3326 3620 3332 3621
rect 3838 3620 3839 3624
rect 3843 3620 3844 3624
rect 3326 3616 3327 3620
rect 3331 3616 3332 3620
rect 3326 3615 3332 3616
rect 3798 3619 3804 3620
rect 3838 3619 3844 3620
rect 4018 3623 4024 3624
rect 4018 3619 4019 3623
rect 4023 3619 4024 3623
rect 3798 3615 3799 3619
rect 3803 3615 3804 3619
rect 4018 3618 4024 3619
rect 4154 3623 4160 3624
rect 4154 3619 4155 3623
rect 4159 3619 4160 3623
rect 4154 3618 4160 3619
rect 4290 3623 4296 3624
rect 4290 3619 4291 3623
rect 4295 3619 4296 3623
rect 4290 3618 4296 3619
rect 4426 3623 4432 3624
rect 4426 3619 4427 3623
rect 4431 3619 4432 3623
rect 4426 3618 4432 3619
rect 4562 3623 4568 3624
rect 4562 3619 4563 3623
rect 4567 3619 4568 3623
rect 4562 3618 4568 3619
rect 4698 3623 4704 3624
rect 4698 3619 4699 3623
rect 4703 3619 4704 3623
rect 4698 3618 4704 3619
rect 4834 3623 4840 3624
rect 4834 3619 4835 3623
rect 4839 3619 4840 3623
rect 4834 3618 4840 3619
rect 4970 3623 4976 3624
rect 4970 3619 4971 3623
rect 4975 3619 4976 3623
rect 4970 3618 4976 3619
rect 5106 3623 5112 3624
rect 5106 3619 5107 3623
rect 5111 3619 5112 3623
rect 5106 3618 5112 3619
rect 5242 3623 5248 3624
rect 5242 3619 5243 3623
rect 5247 3619 5248 3623
rect 5242 3618 5248 3619
rect 5378 3623 5384 3624
rect 5378 3619 5379 3623
rect 5383 3619 5384 3623
rect 5378 3618 5384 3619
rect 5514 3623 5520 3624
rect 5514 3619 5515 3623
rect 5519 3619 5520 3623
rect 5662 3620 5663 3624
rect 5667 3620 5668 3624
rect 5662 3619 5668 3620
rect 5514 3618 5520 3619
rect 1974 3614 1980 3615
rect 1976 3583 1978 3614
rect 2040 3583 2042 3615
rect 2176 3583 2178 3615
rect 2320 3583 2322 3615
rect 2464 3583 2466 3615
rect 2608 3583 2610 3615
rect 2752 3583 2754 3615
rect 2896 3583 2898 3615
rect 3040 3583 3042 3615
rect 3184 3583 3186 3615
rect 3328 3583 3330 3615
rect 3798 3614 3804 3615
rect 3800 3583 3802 3614
rect 4046 3608 4052 3609
rect 3838 3607 3844 3608
rect 3838 3603 3839 3607
rect 3843 3603 3844 3607
rect 4046 3604 4047 3608
rect 4051 3604 4052 3608
rect 4046 3603 4052 3604
rect 4182 3608 4188 3609
rect 4182 3604 4183 3608
rect 4187 3604 4188 3608
rect 4182 3603 4188 3604
rect 4318 3608 4324 3609
rect 4318 3604 4319 3608
rect 4323 3604 4324 3608
rect 4318 3603 4324 3604
rect 4454 3608 4460 3609
rect 4454 3604 4455 3608
rect 4459 3604 4460 3608
rect 4454 3603 4460 3604
rect 4590 3608 4596 3609
rect 4590 3604 4591 3608
rect 4595 3604 4596 3608
rect 4590 3603 4596 3604
rect 4726 3608 4732 3609
rect 4726 3604 4727 3608
rect 4731 3604 4732 3608
rect 4726 3603 4732 3604
rect 4862 3608 4868 3609
rect 4862 3604 4863 3608
rect 4867 3604 4868 3608
rect 4862 3603 4868 3604
rect 4998 3608 5004 3609
rect 4998 3604 4999 3608
rect 5003 3604 5004 3608
rect 4998 3603 5004 3604
rect 5134 3608 5140 3609
rect 5134 3604 5135 3608
rect 5139 3604 5140 3608
rect 5134 3603 5140 3604
rect 5270 3608 5276 3609
rect 5270 3604 5271 3608
rect 5275 3604 5276 3608
rect 5270 3603 5276 3604
rect 5406 3608 5412 3609
rect 5406 3604 5407 3608
rect 5411 3604 5412 3608
rect 5406 3603 5412 3604
rect 5542 3608 5548 3609
rect 5542 3604 5543 3608
rect 5547 3604 5548 3608
rect 5542 3603 5548 3604
rect 5662 3607 5668 3608
rect 5662 3603 5663 3607
rect 5667 3603 5668 3607
rect 3838 3602 3844 3603
rect 1975 3582 1979 3583
rect 1975 3577 1979 3578
rect 2039 3582 2043 3583
rect 2039 3577 2043 3578
rect 2175 3582 2179 3583
rect 2175 3577 2179 3578
rect 2239 3582 2243 3583
rect 2239 3577 2243 3578
rect 2319 3582 2323 3583
rect 2319 3577 2323 3578
rect 2375 3582 2379 3583
rect 2375 3577 2379 3578
rect 2463 3582 2467 3583
rect 2463 3577 2467 3578
rect 2511 3582 2515 3583
rect 2511 3577 2515 3578
rect 2607 3582 2611 3583
rect 2607 3577 2611 3578
rect 2647 3582 2651 3583
rect 2647 3577 2651 3578
rect 2751 3582 2755 3583
rect 2751 3577 2755 3578
rect 2783 3582 2787 3583
rect 2783 3577 2787 3578
rect 2895 3582 2899 3583
rect 2895 3577 2899 3578
rect 2919 3582 2923 3583
rect 2919 3577 2923 3578
rect 3039 3582 3043 3583
rect 3039 3577 3043 3578
rect 3055 3582 3059 3583
rect 3055 3577 3059 3578
rect 3183 3582 3187 3583
rect 3183 3577 3187 3578
rect 3191 3582 3195 3583
rect 3191 3577 3195 3578
rect 3327 3582 3331 3583
rect 3327 3577 3331 3578
rect 3463 3582 3467 3583
rect 3463 3577 3467 3578
rect 3799 3582 3803 3583
rect 3799 3577 3803 3578
rect 1934 3572 1940 3573
rect 110 3568 111 3572
rect 115 3568 116 3572
rect 110 3567 116 3568
rect 490 3571 496 3572
rect 490 3567 491 3571
rect 495 3567 496 3571
rect 490 3566 496 3567
rect 634 3571 640 3572
rect 634 3567 635 3571
rect 639 3567 640 3571
rect 634 3566 640 3567
rect 778 3571 784 3572
rect 778 3567 779 3571
rect 783 3567 784 3571
rect 778 3566 784 3567
rect 922 3571 928 3572
rect 922 3567 923 3571
rect 927 3567 928 3571
rect 922 3566 928 3567
rect 1066 3571 1072 3572
rect 1066 3567 1067 3571
rect 1071 3567 1072 3571
rect 1066 3566 1072 3567
rect 1210 3571 1216 3572
rect 1210 3567 1211 3571
rect 1215 3567 1216 3571
rect 1934 3568 1935 3572
rect 1939 3568 1940 3572
rect 1934 3567 1940 3568
rect 1210 3566 1216 3567
rect 518 3556 524 3557
rect 110 3555 116 3556
rect 110 3551 111 3555
rect 115 3551 116 3555
rect 518 3552 519 3556
rect 523 3552 524 3556
rect 518 3551 524 3552
rect 662 3556 668 3557
rect 662 3552 663 3556
rect 667 3552 668 3556
rect 662 3551 668 3552
rect 806 3556 812 3557
rect 806 3552 807 3556
rect 811 3552 812 3556
rect 806 3551 812 3552
rect 950 3556 956 3557
rect 950 3552 951 3556
rect 955 3552 956 3556
rect 950 3551 956 3552
rect 1094 3556 1100 3557
rect 1094 3552 1095 3556
rect 1099 3552 1100 3556
rect 1094 3551 1100 3552
rect 1238 3556 1244 3557
rect 1238 3552 1239 3556
rect 1243 3552 1244 3556
rect 1238 3551 1244 3552
rect 1934 3555 1940 3556
rect 1934 3551 1935 3555
rect 1939 3551 1940 3555
rect 1976 3554 1978 3577
rect 110 3550 116 3551
rect 112 3507 114 3550
rect 520 3507 522 3551
rect 664 3507 666 3551
rect 808 3507 810 3551
rect 952 3507 954 3551
rect 1096 3507 1098 3551
rect 1240 3507 1242 3551
rect 1934 3550 1940 3551
rect 1974 3553 1980 3554
rect 2240 3553 2242 3577
rect 2376 3553 2378 3577
rect 2512 3553 2514 3577
rect 2648 3553 2650 3577
rect 2784 3553 2786 3577
rect 2920 3553 2922 3577
rect 3056 3553 3058 3577
rect 3192 3553 3194 3577
rect 3328 3553 3330 3577
rect 3464 3553 3466 3577
rect 3800 3554 3802 3577
rect 3798 3553 3804 3554
rect 1936 3507 1938 3550
rect 1974 3549 1975 3553
rect 1979 3549 1980 3553
rect 1974 3548 1980 3549
rect 2238 3552 2244 3553
rect 2238 3548 2239 3552
rect 2243 3548 2244 3552
rect 2238 3547 2244 3548
rect 2374 3552 2380 3553
rect 2374 3548 2375 3552
rect 2379 3548 2380 3552
rect 2374 3547 2380 3548
rect 2510 3552 2516 3553
rect 2510 3548 2511 3552
rect 2515 3548 2516 3552
rect 2510 3547 2516 3548
rect 2646 3552 2652 3553
rect 2646 3548 2647 3552
rect 2651 3548 2652 3552
rect 2646 3547 2652 3548
rect 2782 3552 2788 3553
rect 2782 3548 2783 3552
rect 2787 3548 2788 3552
rect 2782 3547 2788 3548
rect 2918 3552 2924 3553
rect 2918 3548 2919 3552
rect 2923 3548 2924 3552
rect 2918 3547 2924 3548
rect 3054 3552 3060 3553
rect 3054 3548 3055 3552
rect 3059 3548 3060 3552
rect 3054 3547 3060 3548
rect 3190 3552 3196 3553
rect 3190 3548 3191 3552
rect 3195 3548 3196 3552
rect 3190 3547 3196 3548
rect 3326 3552 3332 3553
rect 3326 3548 3327 3552
rect 3331 3548 3332 3552
rect 3326 3547 3332 3548
rect 3462 3552 3468 3553
rect 3462 3548 3463 3552
rect 3467 3548 3468 3552
rect 3798 3549 3799 3553
rect 3803 3549 3804 3553
rect 3798 3548 3804 3549
rect 3462 3547 3468 3548
rect 2210 3537 2216 3538
rect 1974 3536 1980 3537
rect 1974 3532 1975 3536
rect 1979 3532 1980 3536
rect 2210 3533 2211 3537
rect 2215 3533 2216 3537
rect 2210 3532 2216 3533
rect 2346 3537 2352 3538
rect 2346 3533 2347 3537
rect 2351 3533 2352 3537
rect 2346 3532 2352 3533
rect 2482 3537 2488 3538
rect 2482 3533 2483 3537
rect 2487 3533 2488 3537
rect 2482 3532 2488 3533
rect 2618 3537 2624 3538
rect 2618 3533 2619 3537
rect 2623 3533 2624 3537
rect 2618 3532 2624 3533
rect 2754 3537 2760 3538
rect 2754 3533 2755 3537
rect 2759 3533 2760 3537
rect 2754 3532 2760 3533
rect 2890 3537 2896 3538
rect 2890 3533 2891 3537
rect 2895 3533 2896 3537
rect 2890 3532 2896 3533
rect 3026 3537 3032 3538
rect 3026 3533 3027 3537
rect 3031 3533 3032 3537
rect 3026 3532 3032 3533
rect 3162 3537 3168 3538
rect 3162 3533 3163 3537
rect 3167 3533 3168 3537
rect 3162 3532 3168 3533
rect 3298 3537 3304 3538
rect 3298 3533 3299 3537
rect 3303 3533 3304 3537
rect 3298 3532 3304 3533
rect 3434 3537 3440 3538
rect 3434 3533 3435 3537
rect 3439 3533 3440 3537
rect 3434 3532 3440 3533
rect 3798 3536 3804 3537
rect 3798 3532 3799 3536
rect 3803 3532 3804 3536
rect 1974 3531 1980 3532
rect 111 3506 115 3507
rect 111 3501 115 3502
rect 431 3506 435 3507
rect 431 3501 435 3502
rect 519 3506 523 3507
rect 519 3501 523 3502
rect 567 3506 571 3507
rect 567 3501 571 3502
rect 663 3506 667 3507
rect 663 3501 667 3502
rect 703 3506 707 3507
rect 703 3501 707 3502
rect 807 3506 811 3507
rect 807 3501 811 3502
rect 839 3506 843 3507
rect 839 3501 843 3502
rect 951 3506 955 3507
rect 951 3501 955 3502
rect 975 3506 979 3507
rect 975 3501 979 3502
rect 1095 3506 1099 3507
rect 1095 3501 1099 3502
rect 1239 3506 1243 3507
rect 1239 3501 1243 3502
rect 1935 3506 1939 3507
rect 1935 3501 1939 3502
rect 112 3478 114 3501
rect 110 3477 116 3478
rect 432 3477 434 3501
rect 568 3477 570 3501
rect 704 3477 706 3501
rect 840 3477 842 3501
rect 976 3477 978 3501
rect 1936 3478 1938 3501
rect 1934 3477 1940 3478
rect 110 3473 111 3477
rect 115 3473 116 3477
rect 110 3472 116 3473
rect 430 3476 436 3477
rect 430 3472 431 3476
rect 435 3472 436 3476
rect 430 3471 436 3472
rect 566 3476 572 3477
rect 566 3472 567 3476
rect 571 3472 572 3476
rect 566 3471 572 3472
rect 702 3476 708 3477
rect 702 3472 703 3476
rect 707 3472 708 3476
rect 702 3471 708 3472
rect 838 3476 844 3477
rect 838 3472 839 3476
rect 843 3472 844 3476
rect 838 3471 844 3472
rect 974 3476 980 3477
rect 974 3472 975 3476
rect 979 3472 980 3476
rect 1934 3473 1935 3477
rect 1939 3473 1940 3477
rect 1934 3472 1940 3473
rect 974 3471 980 3472
rect 1976 3467 1978 3531
rect 2212 3467 2214 3532
rect 2348 3467 2350 3532
rect 2484 3467 2486 3532
rect 2620 3467 2622 3532
rect 2756 3467 2758 3532
rect 2892 3467 2894 3532
rect 3028 3467 3030 3532
rect 3164 3467 3166 3532
rect 3300 3467 3302 3532
rect 3436 3467 3438 3532
rect 3798 3531 3804 3532
rect 3840 3531 3842 3602
rect 4048 3531 4050 3603
rect 4184 3531 4186 3603
rect 4320 3531 4322 3603
rect 4456 3531 4458 3603
rect 4592 3531 4594 3603
rect 4728 3531 4730 3603
rect 4864 3531 4866 3603
rect 5000 3531 5002 3603
rect 5136 3531 5138 3603
rect 5272 3531 5274 3603
rect 5408 3531 5410 3603
rect 5544 3531 5546 3603
rect 5662 3602 5668 3603
rect 5664 3531 5666 3602
rect 3800 3467 3802 3531
rect 3839 3530 3843 3531
rect 3839 3525 3843 3526
rect 4047 3530 4051 3531
rect 4047 3525 4051 3526
rect 4183 3530 4187 3531
rect 4183 3525 4187 3526
rect 4319 3530 4323 3531
rect 4319 3525 4323 3526
rect 4455 3530 4459 3531
rect 4455 3525 4459 3526
rect 4591 3530 4595 3531
rect 4591 3525 4595 3526
rect 4727 3530 4731 3531
rect 4727 3525 4731 3526
rect 4863 3530 4867 3531
rect 4863 3525 4867 3526
rect 4999 3530 5003 3531
rect 4999 3525 5003 3526
rect 5135 3530 5139 3531
rect 5135 3525 5139 3526
rect 5271 3530 5275 3531
rect 5271 3525 5275 3526
rect 5407 3530 5411 3531
rect 5407 3525 5411 3526
rect 5543 3530 5547 3531
rect 5543 3525 5547 3526
rect 5663 3530 5667 3531
rect 5663 3525 5667 3526
rect 3840 3502 3842 3525
rect 3838 3501 3844 3502
rect 5408 3501 5410 3525
rect 5544 3501 5546 3525
rect 5664 3502 5666 3525
rect 5662 3501 5668 3502
rect 3838 3497 3839 3501
rect 3843 3497 3844 3501
rect 3838 3496 3844 3497
rect 5406 3500 5412 3501
rect 5406 3496 5407 3500
rect 5411 3496 5412 3500
rect 5406 3495 5412 3496
rect 5542 3500 5548 3501
rect 5542 3496 5543 3500
rect 5547 3496 5548 3500
rect 5662 3497 5663 3501
rect 5667 3497 5668 3501
rect 5662 3496 5668 3497
rect 5542 3495 5548 3496
rect 5378 3485 5384 3486
rect 3838 3484 3844 3485
rect 3838 3480 3839 3484
rect 3843 3480 3844 3484
rect 5378 3481 5379 3485
rect 5383 3481 5384 3485
rect 5378 3480 5384 3481
rect 5514 3485 5520 3486
rect 5514 3481 5515 3485
rect 5519 3481 5520 3485
rect 5514 3480 5520 3481
rect 5662 3484 5668 3485
rect 5662 3480 5663 3484
rect 5667 3480 5668 3484
rect 3838 3479 3844 3480
rect 1975 3466 1979 3467
rect 402 3461 408 3462
rect 110 3460 116 3461
rect 110 3456 111 3460
rect 115 3456 116 3460
rect 402 3457 403 3461
rect 407 3457 408 3461
rect 402 3456 408 3457
rect 538 3461 544 3462
rect 538 3457 539 3461
rect 543 3457 544 3461
rect 538 3456 544 3457
rect 674 3461 680 3462
rect 674 3457 675 3461
rect 679 3457 680 3461
rect 674 3456 680 3457
rect 810 3461 816 3462
rect 810 3457 811 3461
rect 815 3457 816 3461
rect 810 3456 816 3457
rect 946 3461 952 3462
rect 1975 3461 1979 3462
rect 2171 3466 2175 3467
rect 2171 3461 2175 3462
rect 2211 3466 2215 3467
rect 2211 3461 2215 3462
rect 2347 3466 2351 3467
rect 2347 3461 2351 3462
rect 2483 3466 2487 3467
rect 2483 3461 2487 3462
rect 2531 3466 2535 3467
rect 2531 3461 2535 3462
rect 2619 3466 2623 3467
rect 2619 3461 2623 3462
rect 2715 3466 2719 3467
rect 2715 3461 2719 3462
rect 2755 3466 2759 3467
rect 2755 3461 2759 3462
rect 2891 3466 2895 3467
rect 2891 3461 2895 3462
rect 2907 3466 2911 3467
rect 2907 3461 2911 3462
rect 3027 3466 3031 3467
rect 3027 3461 3031 3462
rect 3099 3466 3103 3467
rect 3099 3461 3103 3462
rect 3163 3466 3167 3467
rect 3163 3461 3167 3462
rect 3291 3466 3295 3467
rect 3291 3461 3295 3462
rect 3299 3466 3303 3467
rect 3299 3461 3303 3462
rect 3435 3466 3439 3467
rect 3435 3461 3439 3462
rect 3483 3466 3487 3467
rect 3483 3461 3487 3462
rect 3651 3466 3655 3467
rect 3651 3461 3655 3462
rect 3799 3466 3803 3467
rect 3799 3461 3803 3462
rect 946 3457 947 3461
rect 951 3457 952 3461
rect 946 3456 952 3457
rect 1934 3460 1940 3461
rect 1934 3456 1935 3460
rect 1939 3456 1940 3460
rect 110 3455 116 3456
rect 112 3387 114 3455
rect 404 3387 406 3456
rect 540 3387 542 3456
rect 676 3387 678 3456
rect 812 3387 814 3456
rect 948 3387 950 3456
rect 1934 3455 1940 3456
rect 1936 3387 1938 3455
rect 1976 3401 1978 3461
rect 1974 3400 1980 3401
rect 2172 3400 2174 3461
rect 2348 3400 2350 3461
rect 2532 3400 2534 3461
rect 2716 3400 2718 3461
rect 2908 3400 2910 3461
rect 3100 3400 3102 3461
rect 3292 3400 3294 3461
rect 3484 3400 3486 3461
rect 3652 3400 3654 3461
rect 3800 3401 3802 3461
rect 3840 3411 3842 3479
rect 5380 3411 5382 3480
rect 5516 3411 5518 3480
rect 5662 3479 5668 3480
rect 5664 3411 5666 3479
rect 3839 3410 3843 3411
rect 3839 3405 3843 3406
rect 3859 3410 3863 3411
rect 3859 3405 3863 3406
rect 4099 3410 4103 3411
rect 4099 3405 4103 3406
rect 4347 3410 4351 3411
rect 4347 3405 4351 3406
rect 4587 3410 4591 3411
rect 4587 3405 4591 3406
rect 4811 3410 4815 3411
rect 4811 3405 4815 3406
rect 5027 3410 5031 3411
rect 5027 3405 5031 3406
rect 5235 3410 5239 3411
rect 5235 3405 5239 3406
rect 5379 3410 5383 3411
rect 5379 3405 5383 3406
rect 5451 3410 5455 3411
rect 5451 3405 5455 3406
rect 5515 3410 5519 3411
rect 5515 3405 5519 3406
rect 5663 3410 5667 3411
rect 5663 3405 5667 3406
rect 3798 3400 3804 3401
rect 1974 3396 1975 3400
rect 1979 3396 1980 3400
rect 1974 3395 1980 3396
rect 2170 3399 2176 3400
rect 2170 3395 2171 3399
rect 2175 3395 2176 3399
rect 2170 3394 2176 3395
rect 2346 3399 2352 3400
rect 2346 3395 2347 3399
rect 2351 3395 2352 3399
rect 2346 3394 2352 3395
rect 2530 3399 2536 3400
rect 2530 3395 2531 3399
rect 2535 3395 2536 3399
rect 2530 3394 2536 3395
rect 2714 3399 2720 3400
rect 2714 3395 2715 3399
rect 2719 3395 2720 3399
rect 2714 3394 2720 3395
rect 2906 3399 2912 3400
rect 2906 3395 2907 3399
rect 2911 3395 2912 3399
rect 2906 3394 2912 3395
rect 3098 3399 3104 3400
rect 3098 3395 3099 3399
rect 3103 3395 3104 3399
rect 3098 3394 3104 3395
rect 3290 3399 3296 3400
rect 3290 3395 3291 3399
rect 3295 3395 3296 3399
rect 3290 3394 3296 3395
rect 3482 3399 3488 3400
rect 3482 3395 3483 3399
rect 3487 3395 3488 3399
rect 3482 3394 3488 3395
rect 3650 3399 3656 3400
rect 3650 3395 3651 3399
rect 3655 3395 3656 3399
rect 3798 3396 3799 3400
rect 3803 3396 3804 3400
rect 3798 3395 3804 3396
rect 3650 3394 3656 3395
rect 111 3386 115 3387
rect 111 3381 115 3382
rect 323 3386 327 3387
rect 323 3381 327 3382
rect 403 3386 407 3387
rect 403 3381 407 3382
rect 459 3386 463 3387
rect 459 3381 463 3382
rect 539 3386 543 3387
rect 539 3381 543 3382
rect 595 3386 599 3387
rect 595 3381 599 3382
rect 675 3386 679 3387
rect 675 3381 679 3382
rect 731 3386 735 3387
rect 731 3381 735 3382
rect 811 3386 815 3387
rect 811 3381 815 3382
rect 867 3386 871 3387
rect 867 3381 871 3382
rect 947 3386 951 3387
rect 947 3381 951 3382
rect 1935 3386 1939 3387
rect 2198 3384 2204 3385
rect 1935 3381 1939 3382
rect 1974 3383 1980 3384
rect 112 3321 114 3381
rect 110 3320 116 3321
rect 324 3320 326 3381
rect 460 3320 462 3381
rect 596 3320 598 3381
rect 732 3320 734 3381
rect 868 3320 870 3381
rect 1936 3321 1938 3381
rect 1974 3379 1975 3383
rect 1979 3379 1980 3383
rect 2198 3380 2199 3384
rect 2203 3380 2204 3384
rect 2198 3379 2204 3380
rect 2374 3384 2380 3385
rect 2374 3380 2375 3384
rect 2379 3380 2380 3384
rect 2374 3379 2380 3380
rect 2558 3384 2564 3385
rect 2558 3380 2559 3384
rect 2563 3380 2564 3384
rect 2558 3379 2564 3380
rect 2742 3384 2748 3385
rect 2742 3380 2743 3384
rect 2747 3380 2748 3384
rect 2742 3379 2748 3380
rect 2934 3384 2940 3385
rect 2934 3380 2935 3384
rect 2939 3380 2940 3384
rect 2934 3379 2940 3380
rect 3126 3384 3132 3385
rect 3126 3380 3127 3384
rect 3131 3380 3132 3384
rect 3126 3379 3132 3380
rect 3318 3384 3324 3385
rect 3318 3380 3319 3384
rect 3323 3380 3324 3384
rect 3318 3379 3324 3380
rect 3510 3384 3516 3385
rect 3510 3380 3511 3384
rect 3515 3380 3516 3384
rect 3510 3379 3516 3380
rect 3678 3384 3684 3385
rect 3678 3380 3679 3384
rect 3683 3380 3684 3384
rect 3678 3379 3684 3380
rect 3798 3383 3804 3384
rect 3798 3379 3799 3383
rect 3803 3379 3804 3383
rect 1974 3378 1980 3379
rect 1976 3331 1978 3378
rect 2200 3331 2202 3379
rect 2376 3331 2378 3379
rect 2560 3331 2562 3379
rect 2744 3331 2746 3379
rect 2936 3331 2938 3379
rect 3128 3331 3130 3379
rect 3320 3331 3322 3379
rect 3512 3331 3514 3379
rect 3680 3331 3682 3379
rect 3798 3378 3804 3379
rect 3800 3331 3802 3378
rect 3840 3345 3842 3405
rect 3838 3344 3844 3345
rect 3860 3344 3862 3405
rect 4100 3344 4102 3405
rect 4348 3344 4350 3405
rect 4588 3344 4590 3405
rect 4812 3344 4814 3405
rect 5028 3344 5030 3405
rect 5236 3344 5238 3405
rect 5452 3344 5454 3405
rect 5664 3345 5666 3405
rect 5662 3344 5668 3345
rect 3838 3340 3839 3344
rect 3843 3340 3844 3344
rect 3838 3339 3844 3340
rect 3858 3343 3864 3344
rect 3858 3339 3859 3343
rect 3863 3339 3864 3343
rect 3858 3338 3864 3339
rect 4098 3343 4104 3344
rect 4098 3339 4099 3343
rect 4103 3339 4104 3343
rect 4098 3338 4104 3339
rect 4346 3343 4352 3344
rect 4346 3339 4347 3343
rect 4351 3339 4352 3343
rect 4346 3338 4352 3339
rect 4586 3343 4592 3344
rect 4586 3339 4587 3343
rect 4591 3339 4592 3343
rect 4586 3338 4592 3339
rect 4810 3343 4816 3344
rect 4810 3339 4811 3343
rect 4815 3339 4816 3343
rect 4810 3338 4816 3339
rect 5026 3343 5032 3344
rect 5026 3339 5027 3343
rect 5031 3339 5032 3343
rect 5026 3338 5032 3339
rect 5234 3343 5240 3344
rect 5234 3339 5235 3343
rect 5239 3339 5240 3343
rect 5234 3338 5240 3339
rect 5450 3343 5456 3344
rect 5450 3339 5451 3343
rect 5455 3339 5456 3343
rect 5662 3340 5663 3344
rect 5667 3340 5668 3344
rect 5662 3339 5668 3340
rect 5450 3338 5456 3339
rect 1975 3330 1979 3331
rect 1975 3325 1979 3326
rect 2151 3330 2155 3331
rect 2151 3325 2155 3326
rect 2199 3330 2203 3331
rect 2199 3325 2203 3326
rect 2375 3330 2379 3331
rect 2375 3325 2379 3326
rect 2399 3330 2403 3331
rect 2399 3325 2403 3326
rect 2559 3330 2563 3331
rect 2559 3325 2563 3326
rect 2687 3330 2691 3331
rect 2687 3325 2691 3326
rect 2743 3330 2747 3331
rect 2743 3325 2747 3326
rect 2935 3330 2939 3331
rect 2935 3325 2939 3326
rect 3015 3330 3019 3331
rect 3015 3325 3019 3326
rect 3127 3330 3131 3331
rect 3127 3325 3131 3326
rect 3319 3330 3323 3331
rect 3319 3325 3323 3326
rect 3359 3330 3363 3331
rect 3359 3325 3363 3326
rect 3511 3330 3515 3331
rect 3511 3325 3515 3326
rect 3679 3330 3683 3331
rect 3679 3325 3683 3326
rect 3799 3330 3803 3331
rect 3886 3328 3892 3329
rect 3799 3325 3803 3326
rect 3838 3327 3844 3328
rect 1934 3320 1940 3321
rect 110 3316 111 3320
rect 115 3316 116 3320
rect 110 3315 116 3316
rect 322 3319 328 3320
rect 322 3315 323 3319
rect 327 3315 328 3319
rect 322 3314 328 3315
rect 458 3319 464 3320
rect 458 3315 459 3319
rect 463 3315 464 3319
rect 458 3314 464 3315
rect 594 3319 600 3320
rect 594 3315 595 3319
rect 599 3315 600 3319
rect 594 3314 600 3315
rect 730 3319 736 3320
rect 730 3315 731 3319
rect 735 3315 736 3319
rect 730 3314 736 3315
rect 866 3319 872 3320
rect 866 3315 867 3319
rect 871 3315 872 3319
rect 1934 3316 1935 3320
rect 1939 3316 1940 3320
rect 1934 3315 1940 3316
rect 866 3314 872 3315
rect 350 3304 356 3305
rect 110 3303 116 3304
rect 110 3299 111 3303
rect 115 3299 116 3303
rect 350 3300 351 3304
rect 355 3300 356 3304
rect 350 3299 356 3300
rect 486 3304 492 3305
rect 486 3300 487 3304
rect 491 3300 492 3304
rect 486 3299 492 3300
rect 622 3304 628 3305
rect 622 3300 623 3304
rect 627 3300 628 3304
rect 622 3299 628 3300
rect 758 3304 764 3305
rect 758 3300 759 3304
rect 763 3300 764 3304
rect 758 3299 764 3300
rect 894 3304 900 3305
rect 894 3300 895 3304
rect 899 3300 900 3304
rect 894 3299 900 3300
rect 1934 3303 1940 3304
rect 1934 3299 1935 3303
rect 1939 3299 1940 3303
rect 1976 3302 1978 3325
rect 110 3298 116 3299
rect 112 3267 114 3298
rect 352 3267 354 3299
rect 488 3267 490 3299
rect 624 3267 626 3299
rect 760 3267 762 3299
rect 896 3267 898 3299
rect 1934 3298 1940 3299
rect 1974 3301 1980 3302
rect 2152 3301 2154 3325
rect 2400 3301 2402 3325
rect 2688 3301 2690 3325
rect 3016 3301 3018 3325
rect 3360 3301 3362 3325
rect 3680 3301 3682 3325
rect 3800 3302 3802 3325
rect 3838 3323 3839 3327
rect 3843 3323 3844 3327
rect 3886 3324 3887 3328
rect 3891 3324 3892 3328
rect 3886 3323 3892 3324
rect 4126 3328 4132 3329
rect 4126 3324 4127 3328
rect 4131 3324 4132 3328
rect 4126 3323 4132 3324
rect 4374 3328 4380 3329
rect 4374 3324 4375 3328
rect 4379 3324 4380 3328
rect 4374 3323 4380 3324
rect 4614 3328 4620 3329
rect 4614 3324 4615 3328
rect 4619 3324 4620 3328
rect 4614 3323 4620 3324
rect 4838 3328 4844 3329
rect 4838 3324 4839 3328
rect 4843 3324 4844 3328
rect 4838 3323 4844 3324
rect 5054 3328 5060 3329
rect 5054 3324 5055 3328
rect 5059 3324 5060 3328
rect 5054 3323 5060 3324
rect 5262 3328 5268 3329
rect 5262 3324 5263 3328
rect 5267 3324 5268 3328
rect 5262 3323 5268 3324
rect 5478 3328 5484 3329
rect 5478 3324 5479 3328
rect 5483 3324 5484 3328
rect 5478 3323 5484 3324
rect 5662 3327 5668 3328
rect 5662 3323 5663 3327
rect 5667 3323 5668 3327
rect 3838 3322 3844 3323
rect 3798 3301 3804 3302
rect 1936 3267 1938 3298
rect 1974 3297 1975 3301
rect 1979 3297 1980 3301
rect 1974 3296 1980 3297
rect 2150 3300 2156 3301
rect 2150 3296 2151 3300
rect 2155 3296 2156 3300
rect 2150 3295 2156 3296
rect 2398 3300 2404 3301
rect 2398 3296 2399 3300
rect 2403 3296 2404 3300
rect 2398 3295 2404 3296
rect 2686 3300 2692 3301
rect 2686 3296 2687 3300
rect 2691 3296 2692 3300
rect 2686 3295 2692 3296
rect 3014 3300 3020 3301
rect 3014 3296 3015 3300
rect 3019 3296 3020 3300
rect 3014 3295 3020 3296
rect 3358 3300 3364 3301
rect 3358 3296 3359 3300
rect 3363 3296 3364 3300
rect 3358 3295 3364 3296
rect 3678 3300 3684 3301
rect 3678 3296 3679 3300
rect 3683 3296 3684 3300
rect 3798 3297 3799 3301
rect 3803 3297 3804 3301
rect 3840 3299 3842 3322
rect 3888 3299 3890 3323
rect 4128 3299 4130 3323
rect 4376 3299 4378 3323
rect 4616 3299 4618 3323
rect 4840 3299 4842 3323
rect 5056 3299 5058 3323
rect 5264 3299 5266 3323
rect 5480 3299 5482 3323
rect 5662 3322 5668 3323
rect 5664 3299 5666 3322
rect 3798 3296 3804 3297
rect 3839 3298 3843 3299
rect 3678 3295 3684 3296
rect 3839 3293 3843 3294
rect 3887 3298 3891 3299
rect 3887 3293 3891 3294
rect 4127 3298 4131 3299
rect 4127 3293 4131 3294
rect 4375 3298 4379 3299
rect 4375 3293 4379 3294
rect 4607 3298 4611 3299
rect 4607 3293 4611 3294
rect 4615 3298 4619 3299
rect 4615 3293 4619 3294
rect 4815 3298 4819 3299
rect 4815 3293 4819 3294
rect 4839 3298 4843 3299
rect 4839 3293 4843 3294
rect 5015 3298 5019 3299
rect 5015 3293 5019 3294
rect 5055 3298 5059 3299
rect 5055 3293 5059 3294
rect 5199 3298 5203 3299
rect 5199 3293 5203 3294
rect 5263 3298 5267 3299
rect 5263 3293 5267 3294
rect 5383 3298 5387 3299
rect 5383 3293 5387 3294
rect 5479 3298 5483 3299
rect 5479 3293 5483 3294
rect 5543 3298 5547 3299
rect 5543 3293 5547 3294
rect 5663 3298 5667 3299
rect 5663 3293 5667 3294
rect 2122 3285 2128 3286
rect 1974 3284 1980 3285
rect 1974 3280 1975 3284
rect 1979 3280 1980 3284
rect 2122 3281 2123 3285
rect 2127 3281 2128 3285
rect 2122 3280 2128 3281
rect 2370 3285 2376 3286
rect 2370 3281 2371 3285
rect 2375 3281 2376 3285
rect 2370 3280 2376 3281
rect 2658 3285 2664 3286
rect 2658 3281 2659 3285
rect 2663 3281 2664 3285
rect 2658 3280 2664 3281
rect 2986 3285 2992 3286
rect 2986 3281 2987 3285
rect 2991 3281 2992 3285
rect 2986 3280 2992 3281
rect 3330 3285 3336 3286
rect 3330 3281 3331 3285
rect 3335 3281 3336 3285
rect 3330 3280 3336 3281
rect 3650 3285 3656 3286
rect 3650 3281 3651 3285
rect 3655 3281 3656 3285
rect 3650 3280 3656 3281
rect 3798 3284 3804 3285
rect 3798 3280 3799 3284
rect 3803 3280 3804 3284
rect 1974 3279 1980 3280
rect 111 3266 115 3267
rect 111 3261 115 3262
rect 159 3266 163 3267
rect 159 3261 163 3262
rect 335 3266 339 3267
rect 335 3261 339 3262
rect 351 3266 355 3267
rect 351 3261 355 3262
rect 487 3266 491 3267
rect 487 3261 491 3262
rect 543 3266 547 3267
rect 543 3261 547 3262
rect 623 3266 627 3267
rect 623 3261 627 3262
rect 751 3266 755 3267
rect 751 3261 755 3262
rect 759 3266 763 3267
rect 759 3261 763 3262
rect 895 3266 899 3267
rect 895 3261 899 3262
rect 959 3266 963 3267
rect 959 3261 963 3262
rect 1935 3266 1939 3267
rect 1935 3261 1939 3262
rect 112 3238 114 3261
rect 110 3237 116 3238
rect 160 3237 162 3261
rect 336 3237 338 3261
rect 544 3237 546 3261
rect 752 3237 754 3261
rect 960 3237 962 3261
rect 1936 3238 1938 3261
rect 1934 3237 1940 3238
rect 110 3233 111 3237
rect 115 3233 116 3237
rect 110 3232 116 3233
rect 158 3236 164 3237
rect 158 3232 159 3236
rect 163 3232 164 3236
rect 158 3231 164 3232
rect 334 3236 340 3237
rect 334 3232 335 3236
rect 339 3232 340 3236
rect 334 3231 340 3232
rect 542 3236 548 3237
rect 542 3232 543 3236
rect 547 3232 548 3236
rect 542 3231 548 3232
rect 750 3236 756 3237
rect 750 3232 751 3236
rect 755 3232 756 3236
rect 750 3231 756 3232
rect 958 3236 964 3237
rect 958 3232 959 3236
rect 963 3232 964 3236
rect 1934 3233 1935 3237
rect 1939 3233 1940 3237
rect 1934 3232 1940 3233
rect 958 3231 964 3232
rect 130 3221 136 3222
rect 110 3220 116 3221
rect 110 3216 111 3220
rect 115 3216 116 3220
rect 130 3217 131 3221
rect 135 3217 136 3221
rect 130 3216 136 3217
rect 306 3221 312 3222
rect 306 3217 307 3221
rect 311 3217 312 3221
rect 306 3216 312 3217
rect 514 3221 520 3222
rect 514 3217 515 3221
rect 519 3217 520 3221
rect 514 3216 520 3217
rect 722 3221 728 3222
rect 722 3217 723 3221
rect 727 3217 728 3221
rect 722 3216 728 3217
rect 930 3221 936 3222
rect 930 3217 931 3221
rect 935 3217 936 3221
rect 930 3216 936 3217
rect 1934 3220 1940 3221
rect 1934 3216 1935 3220
rect 1939 3216 1940 3220
rect 1976 3219 1978 3279
rect 2124 3219 2126 3280
rect 2372 3219 2374 3280
rect 2660 3219 2662 3280
rect 2988 3219 2990 3280
rect 3332 3219 3334 3280
rect 3652 3219 3654 3280
rect 3798 3279 3804 3280
rect 3800 3219 3802 3279
rect 3840 3270 3842 3293
rect 3838 3269 3844 3270
rect 3888 3269 3890 3293
rect 4128 3269 4130 3293
rect 4376 3269 4378 3293
rect 4608 3269 4610 3293
rect 4816 3269 4818 3293
rect 5016 3269 5018 3293
rect 5200 3269 5202 3293
rect 5384 3269 5386 3293
rect 5544 3269 5546 3293
rect 5664 3270 5666 3293
rect 5662 3269 5668 3270
rect 3838 3265 3839 3269
rect 3843 3265 3844 3269
rect 3838 3264 3844 3265
rect 3886 3268 3892 3269
rect 3886 3264 3887 3268
rect 3891 3264 3892 3268
rect 3886 3263 3892 3264
rect 4126 3268 4132 3269
rect 4126 3264 4127 3268
rect 4131 3264 4132 3268
rect 4126 3263 4132 3264
rect 4374 3268 4380 3269
rect 4374 3264 4375 3268
rect 4379 3264 4380 3268
rect 4374 3263 4380 3264
rect 4606 3268 4612 3269
rect 4606 3264 4607 3268
rect 4611 3264 4612 3268
rect 4606 3263 4612 3264
rect 4814 3268 4820 3269
rect 4814 3264 4815 3268
rect 4819 3264 4820 3268
rect 4814 3263 4820 3264
rect 5014 3268 5020 3269
rect 5014 3264 5015 3268
rect 5019 3264 5020 3268
rect 5014 3263 5020 3264
rect 5198 3268 5204 3269
rect 5198 3264 5199 3268
rect 5203 3264 5204 3268
rect 5198 3263 5204 3264
rect 5382 3268 5388 3269
rect 5382 3264 5383 3268
rect 5387 3264 5388 3268
rect 5382 3263 5388 3264
rect 5542 3268 5548 3269
rect 5542 3264 5543 3268
rect 5547 3264 5548 3268
rect 5662 3265 5663 3269
rect 5667 3265 5668 3269
rect 5662 3264 5668 3265
rect 5542 3263 5548 3264
rect 3858 3253 3864 3254
rect 3838 3252 3844 3253
rect 3838 3248 3839 3252
rect 3843 3248 3844 3252
rect 3858 3249 3859 3253
rect 3863 3249 3864 3253
rect 3858 3248 3864 3249
rect 4098 3253 4104 3254
rect 4098 3249 4099 3253
rect 4103 3249 4104 3253
rect 4098 3248 4104 3249
rect 4346 3253 4352 3254
rect 4346 3249 4347 3253
rect 4351 3249 4352 3253
rect 4346 3248 4352 3249
rect 4578 3253 4584 3254
rect 4578 3249 4579 3253
rect 4583 3249 4584 3253
rect 4578 3248 4584 3249
rect 4786 3253 4792 3254
rect 4786 3249 4787 3253
rect 4791 3249 4792 3253
rect 4786 3248 4792 3249
rect 4986 3253 4992 3254
rect 4986 3249 4987 3253
rect 4991 3249 4992 3253
rect 4986 3248 4992 3249
rect 5170 3253 5176 3254
rect 5170 3249 5171 3253
rect 5175 3249 5176 3253
rect 5170 3248 5176 3249
rect 5354 3253 5360 3254
rect 5354 3249 5355 3253
rect 5359 3249 5360 3253
rect 5354 3248 5360 3249
rect 5514 3253 5520 3254
rect 5514 3249 5515 3253
rect 5519 3249 5520 3253
rect 5514 3248 5520 3249
rect 5662 3252 5668 3253
rect 5662 3248 5663 3252
rect 5667 3248 5668 3252
rect 3838 3247 3844 3248
rect 110 3215 116 3216
rect 112 3139 114 3215
rect 132 3139 134 3216
rect 308 3139 310 3216
rect 516 3139 518 3216
rect 724 3139 726 3216
rect 932 3139 934 3216
rect 1934 3215 1940 3216
rect 1975 3218 1979 3219
rect 1936 3139 1938 3215
rect 1975 3213 1979 3214
rect 1995 3218 1999 3219
rect 1995 3213 1999 3214
rect 2123 3218 2127 3219
rect 2123 3213 2127 3214
rect 2147 3218 2151 3219
rect 2147 3213 2151 3214
rect 2347 3218 2351 3219
rect 2347 3213 2351 3214
rect 2371 3218 2375 3219
rect 2371 3213 2375 3214
rect 2555 3218 2559 3219
rect 2555 3213 2559 3214
rect 2659 3218 2663 3219
rect 2659 3213 2663 3214
rect 2771 3218 2775 3219
rect 2771 3213 2775 3214
rect 2987 3218 2991 3219
rect 2987 3213 2991 3214
rect 3211 3218 3215 3219
rect 3211 3213 3215 3214
rect 3331 3218 3335 3219
rect 3331 3213 3335 3214
rect 3443 3218 3447 3219
rect 3443 3213 3447 3214
rect 3651 3218 3655 3219
rect 3651 3213 3655 3214
rect 3799 3218 3803 3219
rect 3799 3213 3803 3214
rect 1976 3153 1978 3213
rect 1974 3152 1980 3153
rect 1996 3152 1998 3213
rect 2148 3152 2150 3213
rect 2348 3152 2350 3213
rect 2556 3152 2558 3213
rect 2772 3152 2774 3213
rect 2988 3152 2990 3213
rect 3212 3152 3214 3213
rect 3444 3152 3446 3213
rect 3652 3152 3654 3213
rect 3800 3153 3802 3213
rect 3840 3171 3842 3247
rect 3860 3171 3862 3248
rect 4100 3171 4102 3248
rect 4348 3171 4350 3248
rect 4580 3171 4582 3248
rect 4788 3171 4790 3248
rect 4988 3171 4990 3248
rect 5172 3171 5174 3248
rect 5356 3171 5358 3248
rect 5516 3171 5518 3248
rect 5662 3247 5668 3248
rect 5664 3171 5666 3247
rect 3839 3170 3843 3171
rect 3839 3165 3843 3166
rect 3859 3170 3863 3171
rect 3859 3165 3863 3166
rect 4099 3170 4103 3171
rect 4099 3165 4103 3166
rect 4347 3170 4351 3171
rect 4347 3165 4351 3166
rect 4467 3170 4471 3171
rect 4467 3165 4471 3166
rect 4579 3170 4583 3171
rect 4579 3165 4583 3166
rect 4651 3170 4655 3171
rect 4651 3165 4655 3166
rect 4787 3170 4791 3171
rect 4787 3165 4791 3166
rect 4859 3170 4863 3171
rect 4859 3165 4863 3166
rect 4987 3170 4991 3171
rect 4987 3165 4991 3166
rect 5075 3170 5079 3171
rect 5075 3165 5079 3166
rect 5171 3170 5175 3171
rect 5171 3165 5175 3166
rect 5307 3170 5311 3171
rect 5307 3165 5311 3166
rect 5355 3170 5359 3171
rect 5355 3165 5359 3166
rect 5515 3170 5519 3171
rect 5515 3165 5519 3166
rect 5663 3170 5667 3171
rect 5663 3165 5667 3166
rect 3798 3152 3804 3153
rect 1974 3148 1975 3152
rect 1979 3148 1980 3152
rect 1974 3147 1980 3148
rect 1994 3151 2000 3152
rect 1994 3147 1995 3151
rect 1999 3147 2000 3151
rect 1994 3146 2000 3147
rect 2146 3151 2152 3152
rect 2146 3147 2147 3151
rect 2151 3147 2152 3151
rect 2146 3146 2152 3147
rect 2346 3151 2352 3152
rect 2346 3147 2347 3151
rect 2351 3147 2352 3151
rect 2346 3146 2352 3147
rect 2554 3151 2560 3152
rect 2554 3147 2555 3151
rect 2559 3147 2560 3151
rect 2554 3146 2560 3147
rect 2770 3151 2776 3152
rect 2770 3147 2771 3151
rect 2775 3147 2776 3151
rect 2770 3146 2776 3147
rect 2986 3151 2992 3152
rect 2986 3147 2987 3151
rect 2991 3147 2992 3151
rect 2986 3146 2992 3147
rect 3210 3151 3216 3152
rect 3210 3147 3211 3151
rect 3215 3147 3216 3151
rect 3210 3146 3216 3147
rect 3442 3151 3448 3152
rect 3442 3147 3443 3151
rect 3447 3147 3448 3151
rect 3442 3146 3448 3147
rect 3650 3151 3656 3152
rect 3650 3147 3651 3151
rect 3655 3147 3656 3151
rect 3798 3148 3799 3152
rect 3803 3148 3804 3152
rect 3798 3147 3804 3148
rect 3650 3146 3656 3147
rect 111 3138 115 3139
rect 111 3133 115 3134
rect 131 3138 135 3139
rect 131 3133 135 3134
rect 307 3138 311 3139
rect 307 3133 311 3134
rect 371 3138 375 3139
rect 371 3133 375 3134
rect 515 3138 519 3139
rect 515 3133 519 3134
rect 627 3138 631 3139
rect 627 3133 631 3134
rect 723 3138 727 3139
rect 723 3133 727 3134
rect 875 3138 879 3139
rect 875 3133 879 3134
rect 931 3138 935 3139
rect 931 3133 935 3134
rect 1115 3138 1119 3139
rect 1115 3133 1119 3134
rect 1347 3138 1351 3139
rect 1347 3133 1351 3134
rect 1579 3138 1583 3139
rect 1579 3133 1583 3134
rect 1787 3138 1791 3139
rect 1787 3133 1791 3134
rect 1935 3138 1939 3139
rect 2022 3136 2028 3137
rect 1935 3133 1939 3134
rect 1974 3135 1980 3136
rect 112 3073 114 3133
rect 110 3072 116 3073
rect 132 3072 134 3133
rect 372 3072 374 3133
rect 628 3072 630 3133
rect 876 3072 878 3133
rect 1116 3072 1118 3133
rect 1348 3072 1350 3133
rect 1580 3072 1582 3133
rect 1788 3072 1790 3133
rect 1936 3073 1938 3133
rect 1974 3131 1975 3135
rect 1979 3131 1980 3135
rect 2022 3132 2023 3136
rect 2027 3132 2028 3136
rect 2022 3131 2028 3132
rect 2174 3136 2180 3137
rect 2174 3132 2175 3136
rect 2179 3132 2180 3136
rect 2174 3131 2180 3132
rect 2374 3136 2380 3137
rect 2374 3132 2375 3136
rect 2379 3132 2380 3136
rect 2374 3131 2380 3132
rect 2582 3136 2588 3137
rect 2582 3132 2583 3136
rect 2587 3132 2588 3136
rect 2582 3131 2588 3132
rect 2798 3136 2804 3137
rect 2798 3132 2799 3136
rect 2803 3132 2804 3136
rect 2798 3131 2804 3132
rect 3014 3136 3020 3137
rect 3014 3132 3015 3136
rect 3019 3132 3020 3136
rect 3014 3131 3020 3132
rect 3238 3136 3244 3137
rect 3238 3132 3239 3136
rect 3243 3132 3244 3136
rect 3238 3131 3244 3132
rect 3470 3136 3476 3137
rect 3470 3132 3471 3136
rect 3475 3132 3476 3136
rect 3470 3131 3476 3132
rect 3678 3136 3684 3137
rect 3678 3132 3679 3136
rect 3683 3132 3684 3136
rect 3678 3131 3684 3132
rect 3798 3135 3804 3136
rect 3798 3131 3799 3135
rect 3803 3131 3804 3135
rect 1974 3130 1980 3131
rect 1976 3107 1978 3130
rect 2024 3107 2026 3131
rect 2176 3107 2178 3131
rect 2376 3107 2378 3131
rect 2584 3107 2586 3131
rect 2800 3107 2802 3131
rect 3016 3107 3018 3131
rect 3240 3107 3242 3131
rect 3472 3107 3474 3131
rect 3680 3107 3682 3131
rect 3798 3130 3804 3131
rect 3800 3107 3802 3130
rect 1975 3106 1979 3107
rect 1975 3101 1979 3102
rect 2023 3106 2027 3107
rect 2023 3101 2027 3102
rect 2175 3106 2179 3107
rect 2175 3101 2179 3102
rect 2375 3106 2379 3107
rect 2375 3101 2379 3102
rect 2583 3106 2587 3107
rect 2583 3101 2587 3102
rect 2647 3106 2651 3107
rect 2647 3101 2651 3102
rect 2783 3106 2787 3107
rect 2783 3101 2787 3102
rect 2799 3106 2803 3107
rect 2799 3101 2803 3102
rect 2927 3106 2931 3107
rect 2927 3101 2931 3102
rect 3015 3106 3019 3107
rect 3015 3101 3019 3102
rect 3079 3106 3083 3107
rect 3079 3101 3083 3102
rect 3239 3106 3243 3107
rect 3239 3101 3243 3102
rect 3399 3106 3403 3107
rect 3399 3101 3403 3102
rect 3471 3106 3475 3107
rect 3471 3101 3475 3102
rect 3567 3106 3571 3107
rect 3567 3101 3571 3102
rect 3679 3106 3683 3107
rect 3679 3101 3683 3102
rect 3799 3106 3803 3107
rect 3840 3105 3842 3165
rect 3799 3101 3803 3102
rect 3838 3104 3844 3105
rect 4468 3104 4470 3165
rect 4652 3104 4654 3165
rect 4860 3104 4862 3165
rect 5076 3104 5078 3165
rect 5308 3104 5310 3165
rect 5516 3104 5518 3165
rect 5664 3105 5666 3165
rect 5662 3104 5668 3105
rect 1976 3078 1978 3101
rect 1974 3077 1980 3078
rect 2648 3077 2650 3101
rect 2784 3077 2786 3101
rect 2928 3077 2930 3101
rect 3080 3077 3082 3101
rect 3240 3077 3242 3101
rect 3400 3077 3402 3101
rect 3568 3077 3570 3101
rect 3800 3078 3802 3101
rect 3838 3100 3839 3104
rect 3843 3100 3844 3104
rect 3838 3099 3844 3100
rect 4466 3103 4472 3104
rect 4466 3099 4467 3103
rect 4471 3099 4472 3103
rect 4466 3098 4472 3099
rect 4650 3103 4656 3104
rect 4650 3099 4651 3103
rect 4655 3099 4656 3103
rect 4650 3098 4656 3099
rect 4858 3103 4864 3104
rect 4858 3099 4859 3103
rect 4863 3099 4864 3103
rect 4858 3098 4864 3099
rect 5074 3103 5080 3104
rect 5074 3099 5075 3103
rect 5079 3099 5080 3103
rect 5074 3098 5080 3099
rect 5306 3103 5312 3104
rect 5306 3099 5307 3103
rect 5311 3099 5312 3103
rect 5306 3098 5312 3099
rect 5514 3103 5520 3104
rect 5514 3099 5515 3103
rect 5519 3099 5520 3103
rect 5662 3100 5663 3104
rect 5667 3100 5668 3104
rect 5662 3099 5668 3100
rect 5514 3098 5520 3099
rect 4494 3088 4500 3089
rect 3838 3087 3844 3088
rect 3838 3083 3839 3087
rect 3843 3083 3844 3087
rect 4494 3084 4495 3088
rect 4499 3084 4500 3088
rect 4494 3083 4500 3084
rect 4678 3088 4684 3089
rect 4678 3084 4679 3088
rect 4683 3084 4684 3088
rect 4678 3083 4684 3084
rect 4886 3088 4892 3089
rect 4886 3084 4887 3088
rect 4891 3084 4892 3088
rect 4886 3083 4892 3084
rect 5102 3088 5108 3089
rect 5102 3084 5103 3088
rect 5107 3084 5108 3088
rect 5102 3083 5108 3084
rect 5334 3088 5340 3089
rect 5334 3084 5335 3088
rect 5339 3084 5340 3088
rect 5334 3083 5340 3084
rect 5542 3088 5548 3089
rect 5542 3084 5543 3088
rect 5547 3084 5548 3088
rect 5542 3083 5548 3084
rect 5662 3087 5668 3088
rect 5662 3083 5663 3087
rect 5667 3083 5668 3087
rect 3838 3082 3844 3083
rect 3798 3077 3804 3078
rect 1974 3073 1975 3077
rect 1979 3073 1980 3077
rect 1934 3072 1940 3073
rect 1974 3072 1980 3073
rect 2646 3076 2652 3077
rect 2646 3072 2647 3076
rect 2651 3072 2652 3076
rect 110 3068 111 3072
rect 115 3068 116 3072
rect 110 3067 116 3068
rect 130 3071 136 3072
rect 130 3067 131 3071
rect 135 3067 136 3071
rect 130 3066 136 3067
rect 370 3071 376 3072
rect 370 3067 371 3071
rect 375 3067 376 3071
rect 370 3066 376 3067
rect 626 3071 632 3072
rect 626 3067 627 3071
rect 631 3067 632 3071
rect 626 3066 632 3067
rect 874 3071 880 3072
rect 874 3067 875 3071
rect 879 3067 880 3071
rect 874 3066 880 3067
rect 1114 3071 1120 3072
rect 1114 3067 1115 3071
rect 1119 3067 1120 3071
rect 1114 3066 1120 3067
rect 1346 3071 1352 3072
rect 1346 3067 1347 3071
rect 1351 3067 1352 3071
rect 1346 3066 1352 3067
rect 1578 3071 1584 3072
rect 1578 3067 1579 3071
rect 1583 3067 1584 3071
rect 1578 3066 1584 3067
rect 1786 3071 1792 3072
rect 1786 3067 1787 3071
rect 1791 3067 1792 3071
rect 1934 3068 1935 3072
rect 1939 3068 1940 3072
rect 2646 3071 2652 3072
rect 2782 3076 2788 3077
rect 2782 3072 2783 3076
rect 2787 3072 2788 3076
rect 2782 3071 2788 3072
rect 2926 3076 2932 3077
rect 2926 3072 2927 3076
rect 2931 3072 2932 3076
rect 2926 3071 2932 3072
rect 3078 3076 3084 3077
rect 3078 3072 3079 3076
rect 3083 3072 3084 3076
rect 3078 3071 3084 3072
rect 3238 3076 3244 3077
rect 3238 3072 3239 3076
rect 3243 3072 3244 3076
rect 3238 3071 3244 3072
rect 3398 3076 3404 3077
rect 3398 3072 3399 3076
rect 3403 3072 3404 3076
rect 3398 3071 3404 3072
rect 3566 3076 3572 3077
rect 3566 3072 3567 3076
rect 3571 3072 3572 3076
rect 3798 3073 3799 3077
rect 3803 3073 3804 3077
rect 3798 3072 3804 3073
rect 3566 3071 3572 3072
rect 1934 3067 1940 3068
rect 1786 3066 1792 3067
rect 2618 3061 2624 3062
rect 1974 3060 1980 3061
rect 158 3056 164 3057
rect 110 3055 116 3056
rect 110 3051 111 3055
rect 115 3051 116 3055
rect 158 3052 159 3056
rect 163 3052 164 3056
rect 158 3051 164 3052
rect 398 3056 404 3057
rect 398 3052 399 3056
rect 403 3052 404 3056
rect 398 3051 404 3052
rect 654 3056 660 3057
rect 654 3052 655 3056
rect 659 3052 660 3056
rect 654 3051 660 3052
rect 902 3056 908 3057
rect 902 3052 903 3056
rect 907 3052 908 3056
rect 902 3051 908 3052
rect 1142 3056 1148 3057
rect 1142 3052 1143 3056
rect 1147 3052 1148 3056
rect 1142 3051 1148 3052
rect 1374 3056 1380 3057
rect 1374 3052 1375 3056
rect 1379 3052 1380 3056
rect 1374 3051 1380 3052
rect 1606 3056 1612 3057
rect 1606 3052 1607 3056
rect 1611 3052 1612 3056
rect 1606 3051 1612 3052
rect 1814 3056 1820 3057
rect 1974 3056 1975 3060
rect 1979 3056 1980 3060
rect 2618 3057 2619 3061
rect 2623 3057 2624 3061
rect 2618 3056 2624 3057
rect 2754 3061 2760 3062
rect 2754 3057 2755 3061
rect 2759 3057 2760 3061
rect 2754 3056 2760 3057
rect 2898 3061 2904 3062
rect 2898 3057 2899 3061
rect 2903 3057 2904 3061
rect 2898 3056 2904 3057
rect 3050 3061 3056 3062
rect 3050 3057 3051 3061
rect 3055 3057 3056 3061
rect 3050 3056 3056 3057
rect 3210 3061 3216 3062
rect 3210 3057 3211 3061
rect 3215 3057 3216 3061
rect 3210 3056 3216 3057
rect 3370 3061 3376 3062
rect 3370 3057 3371 3061
rect 3375 3057 3376 3061
rect 3370 3056 3376 3057
rect 3538 3061 3544 3062
rect 3538 3057 3539 3061
rect 3543 3057 3544 3061
rect 3538 3056 3544 3057
rect 3798 3060 3804 3061
rect 3798 3056 3799 3060
rect 3803 3056 3804 3060
rect 3840 3059 3842 3082
rect 4496 3059 4498 3083
rect 4680 3059 4682 3083
rect 4888 3059 4890 3083
rect 5104 3059 5106 3083
rect 5336 3059 5338 3083
rect 5544 3059 5546 3083
rect 5662 3082 5668 3083
rect 5664 3059 5666 3082
rect 1814 3052 1815 3056
rect 1819 3052 1820 3056
rect 1814 3051 1820 3052
rect 1934 3055 1940 3056
rect 1974 3055 1980 3056
rect 1934 3051 1935 3055
rect 1939 3051 1940 3055
rect 110 3050 116 3051
rect 112 3027 114 3050
rect 160 3027 162 3051
rect 400 3027 402 3051
rect 656 3027 658 3051
rect 904 3027 906 3051
rect 1144 3027 1146 3051
rect 1376 3027 1378 3051
rect 1608 3027 1610 3051
rect 1816 3027 1818 3051
rect 1934 3050 1940 3051
rect 1936 3027 1938 3050
rect 111 3026 115 3027
rect 111 3021 115 3022
rect 159 3026 163 3027
rect 159 3021 163 3022
rect 175 3026 179 3027
rect 175 3021 179 3022
rect 399 3026 403 3027
rect 399 3021 403 3022
rect 407 3026 411 3027
rect 407 3021 411 3022
rect 623 3026 627 3027
rect 623 3021 627 3022
rect 655 3026 659 3027
rect 655 3021 659 3022
rect 823 3026 827 3027
rect 823 3021 827 3022
rect 903 3026 907 3027
rect 903 3021 907 3022
rect 1007 3026 1011 3027
rect 1007 3021 1011 3022
rect 1143 3026 1147 3027
rect 1143 3021 1147 3022
rect 1183 3026 1187 3027
rect 1183 3021 1187 3022
rect 1351 3026 1355 3027
rect 1351 3021 1355 3022
rect 1375 3026 1379 3027
rect 1375 3021 1379 3022
rect 1511 3026 1515 3027
rect 1511 3021 1515 3022
rect 1607 3026 1611 3027
rect 1607 3021 1611 3022
rect 1671 3026 1675 3027
rect 1671 3021 1675 3022
rect 1815 3026 1819 3027
rect 1815 3021 1819 3022
rect 1935 3026 1939 3027
rect 1935 3021 1939 3022
rect 112 2998 114 3021
rect 110 2997 116 2998
rect 176 2997 178 3021
rect 408 2997 410 3021
rect 624 2997 626 3021
rect 824 2997 826 3021
rect 1008 2997 1010 3021
rect 1184 2997 1186 3021
rect 1352 2997 1354 3021
rect 1512 2997 1514 3021
rect 1672 2997 1674 3021
rect 1816 2997 1818 3021
rect 1936 2998 1938 3021
rect 1934 2997 1940 2998
rect 110 2993 111 2997
rect 115 2993 116 2997
rect 110 2992 116 2993
rect 174 2996 180 2997
rect 174 2992 175 2996
rect 179 2992 180 2996
rect 174 2991 180 2992
rect 406 2996 412 2997
rect 406 2992 407 2996
rect 411 2992 412 2996
rect 406 2991 412 2992
rect 622 2996 628 2997
rect 622 2992 623 2996
rect 627 2992 628 2996
rect 622 2991 628 2992
rect 822 2996 828 2997
rect 822 2992 823 2996
rect 827 2992 828 2996
rect 822 2991 828 2992
rect 1006 2996 1012 2997
rect 1006 2992 1007 2996
rect 1011 2992 1012 2996
rect 1006 2991 1012 2992
rect 1182 2996 1188 2997
rect 1182 2992 1183 2996
rect 1187 2992 1188 2996
rect 1182 2991 1188 2992
rect 1350 2996 1356 2997
rect 1350 2992 1351 2996
rect 1355 2992 1356 2996
rect 1350 2991 1356 2992
rect 1510 2996 1516 2997
rect 1510 2992 1511 2996
rect 1515 2992 1516 2996
rect 1510 2991 1516 2992
rect 1670 2996 1676 2997
rect 1670 2992 1671 2996
rect 1675 2992 1676 2996
rect 1670 2991 1676 2992
rect 1814 2996 1820 2997
rect 1814 2992 1815 2996
rect 1819 2992 1820 2996
rect 1934 2993 1935 2997
rect 1939 2993 1940 2997
rect 1976 2995 1978 3055
rect 2620 2995 2622 3056
rect 2756 2995 2758 3056
rect 2900 2995 2902 3056
rect 3052 2995 3054 3056
rect 3212 2995 3214 3056
rect 3372 2995 3374 3056
rect 3540 2995 3542 3056
rect 3798 3055 3804 3056
rect 3839 3058 3843 3059
rect 3800 2995 3802 3055
rect 3839 3053 3843 3054
rect 4255 3058 4259 3059
rect 4255 3053 4259 3054
rect 4455 3058 4459 3059
rect 4455 3053 4459 3054
rect 4495 3058 4499 3059
rect 4495 3053 4499 3054
rect 4671 3058 4675 3059
rect 4671 3053 4675 3054
rect 4679 3058 4683 3059
rect 4679 3053 4683 3054
rect 4887 3058 4891 3059
rect 4887 3053 4891 3054
rect 4911 3058 4915 3059
rect 4911 3053 4915 3054
rect 5103 3058 5107 3059
rect 5103 3053 5107 3054
rect 5167 3058 5171 3059
rect 5167 3053 5171 3054
rect 5335 3058 5339 3059
rect 5335 3053 5339 3054
rect 5423 3058 5427 3059
rect 5423 3053 5427 3054
rect 5543 3058 5547 3059
rect 5543 3053 5547 3054
rect 5663 3058 5667 3059
rect 5663 3053 5667 3054
rect 3840 3030 3842 3053
rect 3838 3029 3844 3030
rect 4256 3029 4258 3053
rect 4456 3029 4458 3053
rect 4672 3029 4674 3053
rect 4912 3029 4914 3053
rect 5168 3029 5170 3053
rect 5424 3029 5426 3053
rect 5664 3030 5666 3053
rect 5662 3029 5668 3030
rect 3838 3025 3839 3029
rect 3843 3025 3844 3029
rect 3838 3024 3844 3025
rect 4254 3028 4260 3029
rect 4254 3024 4255 3028
rect 4259 3024 4260 3028
rect 4254 3023 4260 3024
rect 4454 3028 4460 3029
rect 4454 3024 4455 3028
rect 4459 3024 4460 3028
rect 4454 3023 4460 3024
rect 4670 3028 4676 3029
rect 4670 3024 4671 3028
rect 4675 3024 4676 3028
rect 4670 3023 4676 3024
rect 4910 3028 4916 3029
rect 4910 3024 4911 3028
rect 4915 3024 4916 3028
rect 4910 3023 4916 3024
rect 5166 3028 5172 3029
rect 5166 3024 5167 3028
rect 5171 3024 5172 3028
rect 5166 3023 5172 3024
rect 5422 3028 5428 3029
rect 5422 3024 5423 3028
rect 5427 3024 5428 3028
rect 5662 3025 5663 3029
rect 5667 3025 5668 3029
rect 5662 3024 5668 3025
rect 5422 3023 5428 3024
rect 4226 3013 4232 3014
rect 3838 3012 3844 3013
rect 3838 3008 3839 3012
rect 3843 3008 3844 3012
rect 4226 3009 4227 3013
rect 4231 3009 4232 3013
rect 4226 3008 4232 3009
rect 4426 3013 4432 3014
rect 4426 3009 4427 3013
rect 4431 3009 4432 3013
rect 4426 3008 4432 3009
rect 4642 3013 4648 3014
rect 4642 3009 4643 3013
rect 4647 3009 4648 3013
rect 4642 3008 4648 3009
rect 4882 3013 4888 3014
rect 4882 3009 4883 3013
rect 4887 3009 4888 3013
rect 4882 3008 4888 3009
rect 5138 3013 5144 3014
rect 5138 3009 5139 3013
rect 5143 3009 5144 3013
rect 5138 3008 5144 3009
rect 5394 3013 5400 3014
rect 5394 3009 5395 3013
rect 5399 3009 5400 3013
rect 5394 3008 5400 3009
rect 5662 3012 5668 3013
rect 5662 3008 5663 3012
rect 5667 3008 5668 3012
rect 3838 3007 3844 3008
rect 1934 2992 1940 2993
rect 1975 2994 1979 2995
rect 1814 2991 1820 2992
rect 1975 2989 1979 2990
rect 2619 2994 2623 2995
rect 2619 2989 2623 2990
rect 2755 2994 2759 2995
rect 2755 2989 2759 2990
rect 2803 2994 2807 2995
rect 2803 2989 2807 2990
rect 2899 2994 2903 2995
rect 2899 2989 2903 2990
rect 2939 2994 2943 2995
rect 2939 2989 2943 2990
rect 3051 2994 3055 2995
rect 3051 2989 3055 2990
rect 3075 2994 3079 2995
rect 3075 2989 3079 2990
rect 3211 2994 3215 2995
rect 3211 2989 3215 2990
rect 3347 2994 3351 2995
rect 3347 2989 3351 2990
rect 3371 2994 3375 2995
rect 3371 2989 3375 2990
rect 3483 2994 3487 2995
rect 3483 2989 3487 2990
rect 3539 2994 3543 2995
rect 3539 2989 3543 2990
rect 3799 2994 3803 2995
rect 3799 2989 3803 2990
rect 146 2981 152 2982
rect 110 2980 116 2981
rect 110 2976 111 2980
rect 115 2976 116 2980
rect 146 2977 147 2981
rect 151 2977 152 2981
rect 146 2976 152 2977
rect 378 2981 384 2982
rect 378 2977 379 2981
rect 383 2977 384 2981
rect 378 2976 384 2977
rect 594 2981 600 2982
rect 594 2977 595 2981
rect 599 2977 600 2981
rect 594 2976 600 2977
rect 794 2981 800 2982
rect 794 2977 795 2981
rect 799 2977 800 2981
rect 794 2976 800 2977
rect 978 2981 984 2982
rect 978 2977 979 2981
rect 983 2977 984 2981
rect 978 2976 984 2977
rect 1154 2981 1160 2982
rect 1154 2977 1155 2981
rect 1159 2977 1160 2981
rect 1154 2976 1160 2977
rect 1322 2981 1328 2982
rect 1322 2977 1323 2981
rect 1327 2977 1328 2981
rect 1322 2976 1328 2977
rect 1482 2981 1488 2982
rect 1482 2977 1483 2981
rect 1487 2977 1488 2981
rect 1482 2976 1488 2977
rect 1642 2981 1648 2982
rect 1642 2977 1643 2981
rect 1647 2977 1648 2981
rect 1642 2976 1648 2977
rect 1786 2981 1792 2982
rect 1786 2977 1787 2981
rect 1791 2977 1792 2981
rect 1786 2976 1792 2977
rect 1934 2980 1940 2981
rect 1934 2976 1935 2980
rect 1939 2976 1940 2980
rect 110 2975 116 2976
rect 112 2911 114 2975
rect 148 2911 150 2976
rect 380 2911 382 2976
rect 596 2911 598 2976
rect 796 2911 798 2976
rect 980 2911 982 2976
rect 1156 2911 1158 2976
rect 1324 2911 1326 2976
rect 1484 2911 1486 2976
rect 1644 2911 1646 2976
rect 1788 2911 1790 2976
rect 1934 2975 1940 2976
rect 1936 2911 1938 2975
rect 1976 2929 1978 2989
rect 1974 2928 1980 2929
rect 2804 2928 2806 2989
rect 2940 2928 2942 2989
rect 3076 2928 3078 2989
rect 3212 2928 3214 2989
rect 3348 2928 3350 2989
rect 3484 2928 3486 2989
rect 3800 2929 3802 2989
rect 3798 2928 3804 2929
rect 1974 2924 1975 2928
rect 1979 2924 1980 2928
rect 1974 2923 1980 2924
rect 2802 2927 2808 2928
rect 2802 2923 2803 2927
rect 2807 2923 2808 2927
rect 2802 2922 2808 2923
rect 2938 2927 2944 2928
rect 2938 2923 2939 2927
rect 2943 2923 2944 2927
rect 2938 2922 2944 2923
rect 3074 2927 3080 2928
rect 3074 2923 3075 2927
rect 3079 2923 3080 2927
rect 3074 2922 3080 2923
rect 3210 2927 3216 2928
rect 3210 2923 3211 2927
rect 3215 2923 3216 2927
rect 3210 2922 3216 2923
rect 3346 2927 3352 2928
rect 3346 2923 3347 2927
rect 3351 2923 3352 2927
rect 3346 2922 3352 2923
rect 3482 2927 3488 2928
rect 3482 2923 3483 2927
rect 3487 2923 3488 2927
rect 3798 2924 3799 2928
rect 3803 2924 3804 2928
rect 3798 2923 3804 2924
rect 3840 2923 3842 3007
rect 4228 2923 4230 3008
rect 4428 2923 4430 3008
rect 4644 2923 4646 3008
rect 4884 2923 4886 3008
rect 5140 2923 5142 3008
rect 5396 2923 5398 3008
rect 5662 3007 5668 3008
rect 5664 2923 5666 3007
rect 3482 2922 3488 2923
rect 3839 2922 3843 2923
rect 3839 2917 3843 2918
rect 3995 2922 3999 2923
rect 3995 2917 3999 2918
rect 4211 2922 4215 2923
rect 4211 2917 4215 2918
rect 4227 2922 4231 2923
rect 4227 2917 4231 2918
rect 4427 2922 4431 2923
rect 4427 2917 4431 2918
rect 4443 2922 4447 2923
rect 4443 2917 4447 2918
rect 4643 2922 4647 2923
rect 4643 2917 4647 2918
rect 4699 2922 4703 2923
rect 4699 2917 4703 2918
rect 4883 2922 4887 2923
rect 4883 2917 4887 2918
rect 4971 2922 4975 2923
rect 4971 2917 4975 2918
rect 5139 2922 5143 2923
rect 5139 2917 5143 2918
rect 5251 2922 5255 2923
rect 5251 2917 5255 2918
rect 5395 2922 5399 2923
rect 5395 2917 5399 2918
rect 5515 2922 5519 2923
rect 5515 2917 5519 2918
rect 5663 2922 5667 2923
rect 5663 2917 5667 2918
rect 2830 2912 2836 2913
rect 1974 2911 1980 2912
rect 111 2910 115 2911
rect 111 2905 115 2906
rect 147 2910 151 2911
rect 147 2905 151 2906
rect 379 2910 383 2911
rect 379 2905 383 2906
rect 395 2910 399 2911
rect 395 2905 399 2906
rect 595 2910 599 2911
rect 595 2905 599 2906
rect 787 2910 791 2911
rect 787 2905 791 2906
rect 795 2910 799 2911
rect 795 2905 799 2906
rect 971 2910 975 2911
rect 971 2905 975 2906
rect 979 2910 983 2911
rect 979 2905 983 2906
rect 1147 2910 1151 2911
rect 1147 2905 1151 2906
rect 1155 2910 1159 2911
rect 1155 2905 1159 2906
rect 1315 2910 1319 2911
rect 1315 2905 1319 2906
rect 1323 2910 1327 2911
rect 1323 2905 1327 2906
rect 1483 2910 1487 2911
rect 1483 2905 1487 2906
rect 1643 2910 1647 2911
rect 1643 2905 1647 2906
rect 1787 2910 1791 2911
rect 1787 2905 1791 2906
rect 1935 2910 1939 2911
rect 1974 2907 1975 2911
rect 1979 2907 1980 2911
rect 2830 2908 2831 2912
rect 2835 2908 2836 2912
rect 2830 2907 2836 2908
rect 2966 2912 2972 2913
rect 2966 2908 2967 2912
rect 2971 2908 2972 2912
rect 2966 2907 2972 2908
rect 3102 2912 3108 2913
rect 3102 2908 3103 2912
rect 3107 2908 3108 2912
rect 3102 2907 3108 2908
rect 3238 2912 3244 2913
rect 3238 2908 3239 2912
rect 3243 2908 3244 2912
rect 3238 2907 3244 2908
rect 3374 2912 3380 2913
rect 3374 2908 3375 2912
rect 3379 2908 3380 2912
rect 3374 2907 3380 2908
rect 3510 2912 3516 2913
rect 3510 2908 3511 2912
rect 3515 2908 3516 2912
rect 3510 2907 3516 2908
rect 3798 2911 3804 2912
rect 3798 2907 3799 2911
rect 3803 2907 3804 2911
rect 1974 2906 1980 2907
rect 1935 2905 1939 2906
rect 112 2845 114 2905
rect 110 2844 116 2845
rect 396 2844 398 2905
rect 596 2844 598 2905
rect 788 2844 790 2905
rect 972 2844 974 2905
rect 1148 2844 1150 2905
rect 1316 2844 1318 2905
rect 1484 2844 1486 2905
rect 1644 2844 1646 2905
rect 1788 2844 1790 2905
rect 1936 2845 1938 2905
rect 1934 2844 1940 2845
rect 110 2840 111 2844
rect 115 2840 116 2844
rect 110 2839 116 2840
rect 394 2843 400 2844
rect 394 2839 395 2843
rect 399 2839 400 2843
rect 394 2838 400 2839
rect 594 2843 600 2844
rect 594 2839 595 2843
rect 599 2839 600 2843
rect 594 2838 600 2839
rect 786 2843 792 2844
rect 786 2839 787 2843
rect 791 2839 792 2843
rect 786 2838 792 2839
rect 970 2843 976 2844
rect 970 2839 971 2843
rect 975 2839 976 2843
rect 970 2838 976 2839
rect 1146 2843 1152 2844
rect 1146 2839 1147 2843
rect 1151 2839 1152 2843
rect 1146 2838 1152 2839
rect 1314 2843 1320 2844
rect 1314 2839 1315 2843
rect 1319 2839 1320 2843
rect 1314 2838 1320 2839
rect 1482 2843 1488 2844
rect 1482 2839 1483 2843
rect 1487 2839 1488 2843
rect 1482 2838 1488 2839
rect 1642 2843 1648 2844
rect 1642 2839 1643 2843
rect 1647 2839 1648 2843
rect 1642 2838 1648 2839
rect 1786 2843 1792 2844
rect 1786 2839 1787 2843
rect 1791 2839 1792 2843
rect 1934 2840 1935 2844
rect 1939 2840 1940 2844
rect 1934 2839 1940 2840
rect 1786 2838 1792 2839
rect 1976 2831 1978 2906
rect 2832 2831 2834 2907
rect 2968 2831 2970 2907
rect 3104 2831 3106 2907
rect 3240 2831 3242 2907
rect 3376 2831 3378 2907
rect 3512 2831 3514 2907
rect 3798 2906 3804 2907
rect 3800 2831 3802 2906
rect 3840 2857 3842 2917
rect 3838 2856 3844 2857
rect 3996 2856 3998 2917
rect 4212 2856 4214 2917
rect 4444 2856 4446 2917
rect 4700 2856 4702 2917
rect 4972 2856 4974 2917
rect 5252 2856 5254 2917
rect 5516 2856 5518 2917
rect 5664 2857 5666 2917
rect 5662 2856 5668 2857
rect 3838 2852 3839 2856
rect 3843 2852 3844 2856
rect 3838 2851 3844 2852
rect 3994 2855 4000 2856
rect 3994 2851 3995 2855
rect 3999 2851 4000 2855
rect 3994 2850 4000 2851
rect 4210 2855 4216 2856
rect 4210 2851 4211 2855
rect 4215 2851 4216 2855
rect 4210 2850 4216 2851
rect 4442 2855 4448 2856
rect 4442 2851 4443 2855
rect 4447 2851 4448 2855
rect 4442 2850 4448 2851
rect 4698 2855 4704 2856
rect 4698 2851 4699 2855
rect 4703 2851 4704 2855
rect 4698 2850 4704 2851
rect 4970 2855 4976 2856
rect 4970 2851 4971 2855
rect 4975 2851 4976 2855
rect 4970 2850 4976 2851
rect 5250 2855 5256 2856
rect 5250 2851 5251 2855
rect 5255 2851 5256 2855
rect 5250 2850 5256 2851
rect 5514 2855 5520 2856
rect 5514 2851 5515 2855
rect 5519 2851 5520 2855
rect 5662 2852 5663 2856
rect 5667 2852 5668 2856
rect 5662 2851 5668 2852
rect 5514 2850 5520 2851
rect 4022 2840 4028 2841
rect 3838 2839 3844 2840
rect 3838 2835 3839 2839
rect 3843 2835 3844 2839
rect 4022 2836 4023 2840
rect 4027 2836 4028 2840
rect 4022 2835 4028 2836
rect 4238 2840 4244 2841
rect 4238 2836 4239 2840
rect 4243 2836 4244 2840
rect 4238 2835 4244 2836
rect 4470 2840 4476 2841
rect 4470 2836 4471 2840
rect 4475 2836 4476 2840
rect 4470 2835 4476 2836
rect 4726 2840 4732 2841
rect 4726 2836 4727 2840
rect 4731 2836 4732 2840
rect 4726 2835 4732 2836
rect 4998 2840 5004 2841
rect 4998 2836 4999 2840
rect 5003 2836 5004 2840
rect 4998 2835 5004 2836
rect 5278 2840 5284 2841
rect 5278 2836 5279 2840
rect 5283 2836 5284 2840
rect 5278 2835 5284 2836
rect 5542 2840 5548 2841
rect 5542 2836 5543 2840
rect 5547 2836 5548 2840
rect 5542 2835 5548 2836
rect 5662 2839 5668 2840
rect 5662 2835 5663 2839
rect 5667 2835 5668 2839
rect 3838 2834 3844 2835
rect 1975 2830 1979 2831
rect 422 2828 428 2829
rect 110 2827 116 2828
rect 110 2823 111 2827
rect 115 2823 116 2827
rect 422 2824 423 2828
rect 427 2824 428 2828
rect 422 2823 428 2824
rect 622 2828 628 2829
rect 622 2824 623 2828
rect 627 2824 628 2828
rect 622 2823 628 2824
rect 814 2828 820 2829
rect 814 2824 815 2828
rect 819 2824 820 2828
rect 814 2823 820 2824
rect 998 2828 1004 2829
rect 998 2824 999 2828
rect 1003 2824 1004 2828
rect 998 2823 1004 2824
rect 1174 2828 1180 2829
rect 1174 2824 1175 2828
rect 1179 2824 1180 2828
rect 1174 2823 1180 2824
rect 1342 2828 1348 2829
rect 1342 2824 1343 2828
rect 1347 2824 1348 2828
rect 1342 2823 1348 2824
rect 1510 2828 1516 2829
rect 1510 2824 1511 2828
rect 1515 2824 1516 2828
rect 1510 2823 1516 2824
rect 1670 2828 1676 2829
rect 1670 2824 1671 2828
rect 1675 2824 1676 2828
rect 1670 2823 1676 2824
rect 1814 2828 1820 2829
rect 1814 2824 1815 2828
rect 1819 2824 1820 2828
rect 1814 2823 1820 2824
rect 1934 2827 1940 2828
rect 1934 2823 1935 2827
rect 1939 2823 1940 2827
rect 1975 2825 1979 2826
rect 2023 2830 2027 2831
rect 2023 2825 2027 2826
rect 2167 2830 2171 2831
rect 2167 2825 2171 2826
rect 2335 2830 2339 2831
rect 2335 2825 2339 2826
rect 2495 2830 2499 2831
rect 2495 2825 2499 2826
rect 2663 2830 2667 2831
rect 2663 2825 2667 2826
rect 2831 2830 2835 2831
rect 2831 2825 2835 2826
rect 2967 2830 2971 2831
rect 2967 2825 2971 2826
rect 2999 2830 3003 2831
rect 2999 2825 3003 2826
rect 3103 2830 3107 2831
rect 3103 2825 3107 2826
rect 3167 2830 3171 2831
rect 3167 2825 3171 2826
rect 3239 2830 3243 2831
rect 3239 2825 3243 2826
rect 3375 2830 3379 2831
rect 3375 2825 3379 2826
rect 3511 2830 3515 2831
rect 3511 2825 3515 2826
rect 3799 2830 3803 2831
rect 3799 2825 3803 2826
rect 110 2822 116 2823
rect 112 2787 114 2822
rect 424 2787 426 2823
rect 624 2787 626 2823
rect 816 2787 818 2823
rect 1000 2787 1002 2823
rect 1176 2787 1178 2823
rect 1344 2787 1346 2823
rect 1512 2787 1514 2823
rect 1672 2787 1674 2823
rect 1816 2787 1818 2823
rect 1934 2822 1940 2823
rect 1936 2787 1938 2822
rect 1976 2802 1978 2825
rect 1974 2801 1980 2802
rect 2024 2801 2026 2825
rect 2168 2801 2170 2825
rect 2336 2801 2338 2825
rect 2496 2801 2498 2825
rect 2664 2801 2666 2825
rect 2832 2801 2834 2825
rect 3000 2801 3002 2825
rect 3168 2801 3170 2825
rect 3800 2802 3802 2825
rect 3840 2807 3842 2834
rect 4024 2807 4026 2835
rect 4240 2807 4242 2835
rect 4472 2807 4474 2835
rect 4728 2807 4730 2835
rect 5000 2807 5002 2835
rect 5280 2807 5282 2835
rect 5544 2807 5546 2835
rect 5662 2834 5668 2835
rect 5664 2807 5666 2834
rect 3839 2806 3843 2807
rect 3798 2801 3804 2802
rect 3839 2801 3843 2802
rect 3919 2806 3923 2807
rect 3919 2801 3923 2802
rect 4023 2806 4027 2807
rect 4023 2801 4027 2802
rect 4055 2806 4059 2807
rect 4055 2801 4059 2802
rect 4191 2806 4195 2807
rect 4191 2801 4195 2802
rect 4239 2806 4243 2807
rect 4239 2801 4243 2802
rect 4327 2806 4331 2807
rect 4327 2801 4331 2802
rect 4463 2806 4467 2807
rect 4463 2801 4467 2802
rect 4471 2806 4475 2807
rect 4471 2801 4475 2802
rect 4727 2806 4731 2807
rect 4727 2801 4731 2802
rect 4999 2806 5003 2807
rect 4999 2801 5003 2802
rect 5279 2806 5283 2807
rect 5279 2801 5283 2802
rect 5543 2806 5547 2807
rect 5543 2801 5547 2802
rect 5663 2806 5667 2807
rect 5663 2801 5667 2802
rect 1974 2797 1975 2801
rect 1979 2797 1980 2801
rect 1974 2796 1980 2797
rect 2022 2800 2028 2801
rect 2022 2796 2023 2800
rect 2027 2796 2028 2800
rect 2022 2795 2028 2796
rect 2166 2800 2172 2801
rect 2166 2796 2167 2800
rect 2171 2796 2172 2800
rect 2166 2795 2172 2796
rect 2334 2800 2340 2801
rect 2334 2796 2335 2800
rect 2339 2796 2340 2800
rect 2334 2795 2340 2796
rect 2494 2800 2500 2801
rect 2494 2796 2495 2800
rect 2499 2796 2500 2800
rect 2494 2795 2500 2796
rect 2662 2800 2668 2801
rect 2662 2796 2663 2800
rect 2667 2796 2668 2800
rect 2662 2795 2668 2796
rect 2830 2800 2836 2801
rect 2830 2796 2831 2800
rect 2835 2796 2836 2800
rect 2830 2795 2836 2796
rect 2998 2800 3004 2801
rect 2998 2796 2999 2800
rect 3003 2796 3004 2800
rect 2998 2795 3004 2796
rect 3166 2800 3172 2801
rect 3166 2796 3167 2800
rect 3171 2796 3172 2800
rect 3798 2797 3799 2801
rect 3803 2797 3804 2801
rect 3798 2796 3804 2797
rect 3166 2795 3172 2796
rect 111 2786 115 2787
rect 111 2781 115 2782
rect 423 2786 427 2787
rect 423 2781 427 2782
rect 623 2786 627 2787
rect 623 2781 627 2782
rect 655 2786 659 2787
rect 655 2781 659 2782
rect 815 2786 819 2787
rect 815 2781 819 2782
rect 975 2786 979 2787
rect 975 2781 979 2782
rect 999 2786 1003 2787
rect 999 2781 1003 2782
rect 1143 2786 1147 2787
rect 1143 2781 1147 2782
rect 1175 2786 1179 2787
rect 1175 2781 1179 2782
rect 1311 2786 1315 2787
rect 1311 2781 1315 2782
rect 1343 2786 1347 2787
rect 1343 2781 1347 2782
rect 1479 2786 1483 2787
rect 1479 2781 1483 2782
rect 1511 2786 1515 2787
rect 1511 2781 1515 2782
rect 1671 2786 1675 2787
rect 1671 2781 1675 2782
rect 1815 2786 1819 2787
rect 1815 2781 1819 2782
rect 1935 2786 1939 2787
rect 1994 2785 2000 2786
rect 1935 2781 1939 2782
rect 1974 2784 1980 2785
rect 112 2758 114 2781
rect 110 2757 116 2758
rect 656 2757 658 2781
rect 816 2757 818 2781
rect 976 2757 978 2781
rect 1144 2757 1146 2781
rect 1312 2757 1314 2781
rect 1480 2757 1482 2781
rect 1936 2758 1938 2781
rect 1974 2780 1975 2784
rect 1979 2780 1980 2784
rect 1994 2781 1995 2785
rect 1999 2781 2000 2785
rect 1994 2780 2000 2781
rect 2138 2785 2144 2786
rect 2138 2781 2139 2785
rect 2143 2781 2144 2785
rect 2138 2780 2144 2781
rect 2306 2785 2312 2786
rect 2306 2781 2307 2785
rect 2311 2781 2312 2785
rect 2306 2780 2312 2781
rect 2466 2785 2472 2786
rect 2466 2781 2467 2785
rect 2471 2781 2472 2785
rect 2466 2780 2472 2781
rect 2634 2785 2640 2786
rect 2634 2781 2635 2785
rect 2639 2781 2640 2785
rect 2634 2780 2640 2781
rect 2802 2785 2808 2786
rect 2802 2781 2803 2785
rect 2807 2781 2808 2785
rect 2802 2780 2808 2781
rect 2970 2785 2976 2786
rect 2970 2781 2971 2785
rect 2975 2781 2976 2785
rect 2970 2780 2976 2781
rect 3138 2785 3144 2786
rect 3138 2781 3139 2785
rect 3143 2781 3144 2785
rect 3138 2780 3144 2781
rect 3798 2784 3804 2785
rect 3798 2780 3799 2784
rect 3803 2780 3804 2784
rect 1974 2779 1980 2780
rect 1934 2757 1940 2758
rect 110 2753 111 2757
rect 115 2753 116 2757
rect 110 2752 116 2753
rect 654 2756 660 2757
rect 654 2752 655 2756
rect 659 2752 660 2756
rect 654 2751 660 2752
rect 814 2756 820 2757
rect 814 2752 815 2756
rect 819 2752 820 2756
rect 814 2751 820 2752
rect 974 2756 980 2757
rect 974 2752 975 2756
rect 979 2752 980 2756
rect 974 2751 980 2752
rect 1142 2756 1148 2757
rect 1142 2752 1143 2756
rect 1147 2752 1148 2756
rect 1142 2751 1148 2752
rect 1310 2756 1316 2757
rect 1310 2752 1311 2756
rect 1315 2752 1316 2756
rect 1310 2751 1316 2752
rect 1478 2756 1484 2757
rect 1478 2752 1479 2756
rect 1483 2752 1484 2756
rect 1934 2753 1935 2757
rect 1939 2753 1940 2757
rect 1934 2752 1940 2753
rect 1478 2751 1484 2752
rect 626 2741 632 2742
rect 110 2740 116 2741
rect 110 2736 111 2740
rect 115 2736 116 2740
rect 626 2737 627 2741
rect 631 2737 632 2741
rect 626 2736 632 2737
rect 786 2741 792 2742
rect 786 2737 787 2741
rect 791 2737 792 2741
rect 786 2736 792 2737
rect 946 2741 952 2742
rect 946 2737 947 2741
rect 951 2737 952 2741
rect 946 2736 952 2737
rect 1114 2741 1120 2742
rect 1114 2737 1115 2741
rect 1119 2737 1120 2741
rect 1114 2736 1120 2737
rect 1282 2741 1288 2742
rect 1282 2737 1283 2741
rect 1287 2737 1288 2741
rect 1282 2736 1288 2737
rect 1450 2741 1456 2742
rect 1450 2737 1451 2741
rect 1455 2737 1456 2741
rect 1450 2736 1456 2737
rect 1934 2740 1940 2741
rect 1934 2736 1935 2740
rect 1939 2736 1940 2740
rect 110 2735 116 2736
rect 112 2675 114 2735
rect 628 2675 630 2736
rect 788 2675 790 2736
rect 948 2675 950 2736
rect 1116 2675 1118 2736
rect 1284 2675 1286 2736
rect 1452 2675 1454 2736
rect 1934 2735 1940 2736
rect 1936 2675 1938 2735
rect 1976 2719 1978 2779
rect 1996 2719 1998 2780
rect 2140 2719 2142 2780
rect 2308 2719 2310 2780
rect 2468 2719 2470 2780
rect 2636 2719 2638 2780
rect 2804 2719 2806 2780
rect 2972 2719 2974 2780
rect 3140 2719 3142 2780
rect 3798 2779 3804 2780
rect 3800 2719 3802 2779
rect 3840 2778 3842 2801
rect 3838 2777 3844 2778
rect 3920 2777 3922 2801
rect 4056 2777 4058 2801
rect 4192 2777 4194 2801
rect 4328 2777 4330 2801
rect 4464 2777 4466 2801
rect 5664 2778 5666 2801
rect 5662 2777 5668 2778
rect 3838 2773 3839 2777
rect 3843 2773 3844 2777
rect 3838 2772 3844 2773
rect 3918 2776 3924 2777
rect 3918 2772 3919 2776
rect 3923 2772 3924 2776
rect 3918 2771 3924 2772
rect 4054 2776 4060 2777
rect 4054 2772 4055 2776
rect 4059 2772 4060 2776
rect 4054 2771 4060 2772
rect 4190 2776 4196 2777
rect 4190 2772 4191 2776
rect 4195 2772 4196 2776
rect 4190 2771 4196 2772
rect 4326 2776 4332 2777
rect 4326 2772 4327 2776
rect 4331 2772 4332 2776
rect 4326 2771 4332 2772
rect 4462 2776 4468 2777
rect 4462 2772 4463 2776
rect 4467 2772 4468 2776
rect 5662 2773 5663 2777
rect 5667 2773 5668 2777
rect 5662 2772 5668 2773
rect 4462 2771 4468 2772
rect 3890 2761 3896 2762
rect 3838 2760 3844 2761
rect 3838 2756 3839 2760
rect 3843 2756 3844 2760
rect 3890 2757 3891 2761
rect 3895 2757 3896 2761
rect 3890 2756 3896 2757
rect 4026 2761 4032 2762
rect 4026 2757 4027 2761
rect 4031 2757 4032 2761
rect 4026 2756 4032 2757
rect 4162 2761 4168 2762
rect 4162 2757 4163 2761
rect 4167 2757 4168 2761
rect 4162 2756 4168 2757
rect 4298 2761 4304 2762
rect 4298 2757 4299 2761
rect 4303 2757 4304 2761
rect 4298 2756 4304 2757
rect 4434 2761 4440 2762
rect 4434 2757 4435 2761
rect 4439 2757 4440 2761
rect 4434 2756 4440 2757
rect 5662 2760 5668 2761
rect 5662 2756 5663 2760
rect 5667 2756 5668 2760
rect 3838 2755 3844 2756
rect 1975 2718 1979 2719
rect 1975 2713 1979 2714
rect 1995 2718 1999 2719
rect 1995 2713 1999 2714
rect 2139 2718 2143 2719
rect 2139 2713 2143 2714
rect 2307 2718 2311 2719
rect 2307 2713 2311 2714
rect 2379 2718 2383 2719
rect 2379 2713 2383 2714
rect 2467 2718 2471 2719
rect 2467 2713 2471 2714
rect 2515 2718 2519 2719
rect 2515 2713 2519 2714
rect 2635 2718 2639 2719
rect 2635 2713 2639 2714
rect 2659 2718 2663 2719
rect 2659 2713 2663 2714
rect 2803 2718 2807 2719
rect 2803 2713 2807 2714
rect 2947 2718 2951 2719
rect 2947 2713 2951 2714
rect 2971 2718 2975 2719
rect 2971 2713 2975 2714
rect 3091 2718 3095 2719
rect 3091 2713 3095 2714
rect 3139 2718 3143 2719
rect 3139 2713 3143 2714
rect 3235 2718 3239 2719
rect 3235 2713 3239 2714
rect 3799 2718 3803 2719
rect 3799 2713 3803 2714
rect 111 2674 115 2675
rect 111 2669 115 2670
rect 627 2674 631 2675
rect 627 2669 631 2670
rect 771 2674 775 2675
rect 771 2669 775 2670
rect 787 2674 791 2675
rect 787 2669 791 2670
rect 907 2674 911 2675
rect 907 2669 911 2670
rect 947 2674 951 2675
rect 947 2669 951 2670
rect 1043 2674 1047 2675
rect 1043 2669 1047 2670
rect 1115 2674 1119 2675
rect 1115 2669 1119 2670
rect 1179 2674 1183 2675
rect 1179 2669 1183 2670
rect 1283 2674 1287 2675
rect 1283 2669 1287 2670
rect 1315 2674 1319 2675
rect 1315 2669 1319 2670
rect 1451 2674 1455 2675
rect 1451 2669 1455 2670
rect 1587 2674 1591 2675
rect 1587 2669 1591 2670
rect 1723 2674 1727 2675
rect 1723 2669 1727 2670
rect 1935 2674 1939 2675
rect 1935 2669 1939 2670
rect 112 2609 114 2669
rect 110 2608 116 2609
rect 772 2608 774 2669
rect 908 2608 910 2669
rect 1044 2608 1046 2669
rect 1180 2608 1182 2669
rect 1316 2608 1318 2669
rect 1452 2608 1454 2669
rect 1588 2608 1590 2669
rect 1724 2608 1726 2669
rect 1936 2609 1938 2669
rect 1976 2653 1978 2713
rect 1974 2652 1980 2653
rect 2380 2652 2382 2713
rect 2516 2652 2518 2713
rect 2660 2652 2662 2713
rect 2804 2652 2806 2713
rect 2948 2652 2950 2713
rect 3092 2652 3094 2713
rect 3236 2652 3238 2713
rect 3800 2653 3802 2713
rect 3840 2683 3842 2755
rect 3892 2683 3894 2756
rect 4028 2683 4030 2756
rect 4164 2683 4166 2756
rect 4300 2683 4302 2756
rect 4436 2683 4438 2756
rect 5662 2755 5668 2756
rect 5664 2683 5666 2755
rect 3839 2682 3843 2683
rect 3839 2677 3843 2678
rect 3891 2682 3895 2683
rect 3891 2677 3895 2678
rect 4027 2682 4031 2683
rect 4027 2677 4031 2678
rect 4099 2682 4103 2683
rect 4099 2677 4103 2678
rect 4163 2682 4167 2683
rect 4163 2677 4167 2678
rect 4299 2682 4303 2683
rect 4299 2677 4303 2678
rect 4435 2682 4439 2683
rect 4435 2677 4439 2678
rect 4515 2682 4519 2683
rect 4515 2677 4519 2678
rect 4755 2682 4759 2683
rect 4755 2677 4759 2678
rect 5011 2682 5015 2683
rect 5011 2677 5015 2678
rect 5275 2682 5279 2683
rect 5275 2677 5279 2678
rect 5515 2682 5519 2683
rect 5515 2677 5519 2678
rect 5663 2682 5667 2683
rect 5663 2677 5667 2678
rect 3798 2652 3804 2653
rect 1974 2648 1975 2652
rect 1979 2648 1980 2652
rect 1974 2647 1980 2648
rect 2378 2651 2384 2652
rect 2378 2647 2379 2651
rect 2383 2647 2384 2651
rect 2378 2646 2384 2647
rect 2514 2651 2520 2652
rect 2514 2647 2515 2651
rect 2519 2647 2520 2651
rect 2514 2646 2520 2647
rect 2658 2651 2664 2652
rect 2658 2647 2659 2651
rect 2663 2647 2664 2651
rect 2658 2646 2664 2647
rect 2802 2651 2808 2652
rect 2802 2647 2803 2651
rect 2807 2647 2808 2651
rect 2802 2646 2808 2647
rect 2946 2651 2952 2652
rect 2946 2647 2947 2651
rect 2951 2647 2952 2651
rect 2946 2646 2952 2647
rect 3090 2651 3096 2652
rect 3090 2647 3091 2651
rect 3095 2647 3096 2651
rect 3090 2646 3096 2647
rect 3234 2651 3240 2652
rect 3234 2647 3235 2651
rect 3239 2647 3240 2651
rect 3798 2648 3799 2652
rect 3803 2648 3804 2652
rect 3798 2647 3804 2648
rect 3234 2646 3240 2647
rect 2406 2636 2412 2637
rect 1974 2635 1980 2636
rect 1974 2631 1975 2635
rect 1979 2631 1980 2635
rect 2406 2632 2407 2636
rect 2411 2632 2412 2636
rect 2406 2631 2412 2632
rect 2542 2636 2548 2637
rect 2542 2632 2543 2636
rect 2547 2632 2548 2636
rect 2542 2631 2548 2632
rect 2686 2636 2692 2637
rect 2686 2632 2687 2636
rect 2691 2632 2692 2636
rect 2686 2631 2692 2632
rect 2830 2636 2836 2637
rect 2830 2632 2831 2636
rect 2835 2632 2836 2636
rect 2830 2631 2836 2632
rect 2974 2636 2980 2637
rect 2974 2632 2975 2636
rect 2979 2632 2980 2636
rect 2974 2631 2980 2632
rect 3118 2636 3124 2637
rect 3118 2632 3119 2636
rect 3123 2632 3124 2636
rect 3118 2631 3124 2632
rect 3262 2636 3268 2637
rect 3262 2632 3263 2636
rect 3267 2632 3268 2636
rect 3262 2631 3268 2632
rect 3798 2635 3804 2636
rect 3798 2631 3799 2635
rect 3803 2631 3804 2635
rect 1974 2630 1980 2631
rect 1934 2608 1940 2609
rect 110 2604 111 2608
rect 115 2604 116 2608
rect 110 2603 116 2604
rect 770 2607 776 2608
rect 770 2603 771 2607
rect 775 2603 776 2607
rect 770 2602 776 2603
rect 906 2607 912 2608
rect 906 2603 907 2607
rect 911 2603 912 2607
rect 906 2602 912 2603
rect 1042 2607 1048 2608
rect 1042 2603 1043 2607
rect 1047 2603 1048 2607
rect 1042 2602 1048 2603
rect 1178 2607 1184 2608
rect 1178 2603 1179 2607
rect 1183 2603 1184 2607
rect 1178 2602 1184 2603
rect 1314 2607 1320 2608
rect 1314 2603 1315 2607
rect 1319 2603 1320 2607
rect 1314 2602 1320 2603
rect 1450 2607 1456 2608
rect 1450 2603 1451 2607
rect 1455 2603 1456 2607
rect 1450 2602 1456 2603
rect 1586 2607 1592 2608
rect 1586 2603 1587 2607
rect 1591 2603 1592 2607
rect 1586 2602 1592 2603
rect 1722 2607 1728 2608
rect 1722 2603 1723 2607
rect 1727 2603 1728 2607
rect 1934 2604 1935 2608
rect 1939 2604 1940 2608
rect 1934 2603 1940 2604
rect 1976 2603 1978 2630
rect 2408 2603 2410 2631
rect 2544 2603 2546 2631
rect 2688 2603 2690 2631
rect 2832 2603 2834 2631
rect 2976 2603 2978 2631
rect 3120 2603 3122 2631
rect 3264 2603 3266 2631
rect 3798 2630 3804 2631
rect 3800 2603 3802 2630
rect 3840 2617 3842 2677
rect 3838 2616 3844 2617
rect 4100 2616 4102 2677
rect 4300 2616 4302 2677
rect 4516 2616 4518 2677
rect 4756 2616 4758 2677
rect 5012 2616 5014 2677
rect 5276 2616 5278 2677
rect 5516 2616 5518 2677
rect 5664 2617 5666 2677
rect 5662 2616 5668 2617
rect 3838 2612 3839 2616
rect 3843 2612 3844 2616
rect 3838 2611 3844 2612
rect 4098 2615 4104 2616
rect 4098 2611 4099 2615
rect 4103 2611 4104 2615
rect 4098 2610 4104 2611
rect 4298 2615 4304 2616
rect 4298 2611 4299 2615
rect 4303 2611 4304 2615
rect 4298 2610 4304 2611
rect 4514 2615 4520 2616
rect 4514 2611 4515 2615
rect 4519 2611 4520 2615
rect 4514 2610 4520 2611
rect 4754 2615 4760 2616
rect 4754 2611 4755 2615
rect 4759 2611 4760 2615
rect 4754 2610 4760 2611
rect 5010 2615 5016 2616
rect 5010 2611 5011 2615
rect 5015 2611 5016 2615
rect 5010 2610 5016 2611
rect 5274 2615 5280 2616
rect 5274 2611 5275 2615
rect 5279 2611 5280 2615
rect 5274 2610 5280 2611
rect 5514 2615 5520 2616
rect 5514 2611 5515 2615
rect 5519 2611 5520 2615
rect 5662 2612 5663 2616
rect 5667 2612 5668 2616
rect 5662 2611 5668 2612
rect 5514 2610 5520 2611
rect 1722 2602 1728 2603
rect 1975 2602 1979 2603
rect 1975 2597 1979 2598
rect 2407 2602 2411 2603
rect 2407 2597 2411 2598
rect 2511 2602 2515 2603
rect 2511 2597 2515 2598
rect 2543 2602 2547 2603
rect 2543 2597 2547 2598
rect 2647 2602 2651 2603
rect 2647 2597 2651 2598
rect 2687 2602 2691 2603
rect 2687 2597 2691 2598
rect 2783 2602 2787 2603
rect 2783 2597 2787 2598
rect 2831 2602 2835 2603
rect 2831 2597 2835 2598
rect 2919 2602 2923 2603
rect 2919 2597 2923 2598
rect 2975 2602 2979 2603
rect 2975 2597 2979 2598
rect 3055 2602 3059 2603
rect 3055 2597 3059 2598
rect 3119 2602 3123 2603
rect 3119 2597 3123 2598
rect 3191 2602 3195 2603
rect 3191 2597 3195 2598
rect 3263 2602 3267 2603
rect 3263 2597 3267 2598
rect 3327 2602 3331 2603
rect 3327 2597 3331 2598
rect 3463 2602 3467 2603
rect 3463 2597 3467 2598
rect 3799 2602 3803 2603
rect 4126 2600 4132 2601
rect 3799 2597 3803 2598
rect 3838 2599 3844 2600
rect 798 2592 804 2593
rect 110 2591 116 2592
rect 110 2587 111 2591
rect 115 2587 116 2591
rect 798 2588 799 2592
rect 803 2588 804 2592
rect 798 2587 804 2588
rect 934 2592 940 2593
rect 934 2588 935 2592
rect 939 2588 940 2592
rect 934 2587 940 2588
rect 1070 2592 1076 2593
rect 1070 2588 1071 2592
rect 1075 2588 1076 2592
rect 1070 2587 1076 2588
rect 1206 2592 1212 2593
rect 1206 2588 1207 2592
rect 1211 2588 1212 2592
rect 1206 2587 1212 2588
rect 1342 2592 1348 2593
rect 1342 2588 1343 2592
rect 1347 2588 1348 2592
rect 1342 2587 1348 2588
rect 1478 2592 1484 2593
rect 1478 2588 1479 2592
rect 1483 2588 1484 2592
rect 1478 2587 1484 2588
rect 1614 2592 1620 2593
rect 1614 2588 1615 2592
rect 1619 2588 1620 2592
rect 1614 2587 1620 2588
rect 1750 2592 1756 2593
rect 1750 2588 1751 2592
rect 1755 2588 1756 2592
rect 1750 2587 1756 2588
rect 1934 2591 1940 2592
rect 1934 2587 1935 2591
rect 1939 2587 1940 2591
rect 110 2586 116 2587
rect 112 2547 114 2586
rect 800 2547 802 2587
rect 936 2547 938 2587
rect 1072 2547 1074 2587
rect 1208 2547 1210 2587
rect 1344 2547 1346 2587
rect 1480 2547 1482 2587
rect 1616 2547 1618 2587
rect 1752 2547 1754 2587
rect 1934 2586 1940 2587
rect 1936 2547 1938 2586
rect 1976 2574 1978 2597
rect 1974 2573 1980 2574
rect 2512 2573 2514 2597
rect 2648 2573 2650 2597
rect 2784 2573 2786 2597
rect 2920 2573 2922 2597
rect 3056 2573 3058 2597
rect 3192 2573 3194 2597
rect 3328 2573 3330 2597
rect 3464 2573 3466 2597
rect 3800 2574 3802 2597
rect 3838 2595 3839 2599
rect 3843 2595 3844 2599
rect 4126 2596 4127 2600
rect 4131 2596 4132 2600
rect 4126 2595 4132 2596
rect 4326 2600 4332 2601
rect 4326 2596 4327 2600
rect 4331 2596 4332 2600
rect 4326 2595 4332 2596
rect 4542 2600 4548 2601
rect 4542 2596 4543 2600
rect 4547 2596 4548 2600
rect 4542 2595 4548 2596
rect 4782 2600 4788 2601
rect 4782 2596 4783 2600
rect 4787 2596 4788 2600
rect 4782 2595 4788 2596
rect 5038 2600 5044 2601
rect 5038 2596 5039 2600
rect 5043 2596 5044 2600
rect 5038 2595 5044 2596
rect 5302 2600 5308 2601
rect 5302 2596 5303 2600
rect 5307 2596 5308 2600
rect 5302 2595 5308 2596
rect 5542 2600 5548 2601
rect 5542 2596 5543 2600
rect 5547 2596 5548 2600
rect 5542 2595 5548 2596
rect 5662 2599 5668 2600
rect 5662 2595 5663 2599
rect 5667 2595 5668 2599
rect 3838 2594 3844 2595
rect 3798 2573 3804 2574
rect 1974 2569 1975 2573
rect 1979 2569 1980 2573
rect 1974 2568 1980 2569
rect 2510 2572 2516 2573
rect 2510 2568 2511 2572
rect 2515 2568 2516 2572
rect 2510 2567 2516 2568
rect 2646 2572 2652 2573
rect 2646 2568 2647 2572
rect 2651 2568 2652 2572
rect 2646 2567 2652 2568
rect 2782 2572 2788 2573
rect 2782 2568 2783 2572
rect 2787 2568 2788 2572
rect 2782 2567 2788 2568
rect 2918 2572 2924 2573
rect 2918 2568 2919 2572
rect 2923 2568 2924 2572
rect 2918 2567 2924 2568
rect 3054 2572 3060 2573
rect 3054 2568 3055 2572
rect 3059 2568 3060 2572
rect 3054 2567 3060 2568
rect 3190 2572 3196 2573
rect 3190 2568 3191 2572
rect 3195 2568 3196 2572
rect 3190 2567 3196 2568
rect 3326 2572 3332 2573
rect 3326 2568 3327 2572
rect 3331 2568 3332 2572
rect 3326 2567 3332 2568
rect 3462 2572 3468 2573
rect 3462 2568 3463 2572
rect 3467 2568 3468 2572
rect 3798 2569 3799 2573
rect 3803 2569 3804 2573
rect 3798 2568 3804 2569
rect 3462 2567 3468 2568
rect 3840 2567 3842 2594
rect 4128 2567 4130 2595
rect 4328 2567 4330 2595
rect 4544 2567 4546 2595
rect 4784 2567 4786 2595
rect 5040 2567 5042 2595
rect 5304 2567 5306 2595
rect 5544 2567 5546 2595
rect 5662 2594 5668 2595
rect 5664 2567 5666 2594
rect 3839 2566 3843 2567
rect 3839 2561 3843 2562
rect 4127 2566 4131 2567
rect 4127 2561 4131 2562
rect 4327 2566 4331 2567
rect 4327 2561 4331 2562
rect 4495 2566 4499 2567
rect 4495 2561 4499 2562
rect 4543 2566 4547 2567
rect 4543 2561 4547 2562
rect 4631 2566 4635 2567
rect 4631 2561 4635 2562
rect 4767 2566 4771 2567
rect 4767 2561 4771 2562
rect 4783 2566 4787 2567
rect 4783 2561 4787 2562
rect 4903 2566 4907 2567
rect 4903 2561 4907 2562
rect 5039 2566 5043 2567
rect 5039 2561 5043 2562
rect 5303 2566 5307 2567
rect 5303 2561 5307 2562
rect 5543 2566 5547 2567
rect 5543 2561 5547 2562
rect 5663 2566 5667 2567
rect 5663 2561 5667 2562
rect 2482 2557 2488 2558
rect 1974 2556 1980 2557
rect 1974 2552 1975 2556
rect 1979 2552 1980 2556
rect 2482 2553 2483 2557
rect 2487 2553 2488 2557
rect 2482 2552 2488 2553
rect 2618 2557 2624 2558
rect 2618 2553 2619 2557
rect 2623 2553 2624 2557
rect 2618 2552 2624 2553
rect 2754 2557 2760 2558
rect 2754 2553 2755 2557
rect 2759 2553 2760 2557
rect 2754 2552 2760 2553
rect 2890 2557 2896 2558
rect 2890 2553 2891 2557
rect 2895 2553 2896 2557
rect 2890 2552 2896 2553
rect 3026 2557 3032 2558
rect 3026 2553 3027 2557
rect 3031 2553 3032 2557
rect 3026 2552 3032 2553
rect 3162 2557 3168 2558
rect 3162 2553 3163 2557
rect 3167 2553 3168 2557
rect 3162 2552 3168 2553
rect 3298 2557 3304 2558
rect 3298 2553 3299 2557
rect 3303 2553 3304 2557
rect 3298 2552 3304 2553
rect 3434 2557 3440 2558
rect 3434 2553 3435 2557
rect 3439 2553 3440 2557
rect 3434 2552 3440 2553
rect 3798 2556 3804 2557
rect 3798 2552 3799 2556
rect 3803 2552 3804 2556
rect 1974 2551 1980 2552
rect 111 2546 115 2547
rect 111 2541 115 2542
rect 551 2546 555 2547
rect 551 2541 555 2542
rect 687 2546 691 2547
rect 687 2541 691 2542
rect 799 2546 803 2547
rect 799 2541 803 2542
rect 831 2546 835 2547
rect 831 2541 835 2542
rect 935 2546 939 2547
rect 935 2541 939 2542
rect 983 2546 987 2547
rect 983 2541 987 2542
rect 1071 2546 1075 2547
rect 1071 2541 1075 2542
rect 1135 2546 1139 2547
rect 1135 2541 1139 2542
rect 1207 2546 1211 2547
rect 1207 2541 1211 2542
rect 1295 2546 1299 2547
rect 1295 2541 1299 2542
rect 1343 2546 1347 2547
rect 1343 2541 1347 2542
rect 1455 2546 1459 2547
rect 1455 2541 1459 2542
rect 1479 2546 1483 2547
rect 1479 2541 1483 2542
rect 1615 2546 1619 2547
rect 1615 2541 1619 2542
rect 1751 2546 1755 2547
rect 1751 2541 1755 2542
rect 1783 2546 1787 2547
rect 1783 2541 1787 2542
rect 1935 2546 1939 2547
rect 1935 2541 1939 2542
rect 112 2518 114 2541
rect 110 2517 116 2518
rect 552 2517 554 2541
rect 688 2517 690 2541
rect 832 2517 834 2541
rect 984 2517 986 2541
rect 1136 2517 1138 2541
rect 1296 2517 1298 2541
rect 1456 2517 1458 2541
rect 1616 2517 1618 2541
rect 1784 2517 1786 2541
rect 1936 2518 1938 2541
rect 1934 2517 1940 2518
rect 110 2513 111 2517
rect 115 2513 116 2517
rect 110 2512 116 2513
rect 550 2516 556 2517
rect 550 2512 551 2516
rect 555 2512 556 2516
rect 550 2511 556 2512
rect 686 2516 692 2517
rect 686 2512 687 2516
rect 691 2512 692 2516
rect 686 2511 692 2512
rect 830 2516 836 2517
rect 830 2512 831 2516
rect 835 2512 836 2516
rect 830 2511 836 2512
rect 982 2516 988 2517
rect 982 2512 983 2516
rect 987 2512 988 2516
rect 982 2511 988 2512
rect 1134 2516 1140 2517
rect 1134 2512 1135 2516
rect 1139 2512 1140 2516
rect 1134 2511 1140 2512
rect 1294 2516 1300 2517
rect 1294 2512 1295 2516
rect 1299 2512 1300 2516
rect 1294 2511 1300 2512
rect 1454 2516 1460 2517
rect 1454 2512 1455 2516
rect 1459 2512 1460 2516
rect 1454 2511 1460 2512
rect 1614 2516 1620 2517
rect 1614 2512 1615 2516
rect 1619 2512 1620 2516
rect 1614 2511 1620 2512
rect 1782 2516 1788 2517
rect 1782 2512 1783 2516
rect 1787 2512 1788 2516
rect 1934 2513 1935 2517
rect 1939 2513 1940 2517
rect 1934 2512 1940 2513
rect 1782 2511 1788 2512
rect 522 2501 528 2502
rect 110 2500 116 2501
rect 110 2496 111 2500
rect 115 2496 116 2500
rect 522 2497 523 2501
rect 527 2497 528 2501
rect 522 2496 528 2497
rect 658 2501 664 2502
rect 658 2497 659 2501
rect 663 2497 664 2501
rect 658 2496 664 2497
rect 802 2501 808 2502
rect 802 2497 803 2501
rect 807 2497 808 2501
rect 802 2496 808 2497
rect 954 2501 960 2502
rect 954 2497 955 2501
rect 959 2497 960 2501
rect 954 2496 960 2497
rect 1106 2501 1112 2502
rect 1106 2497 1107 2501
rect 1111 2497 1112 2501
rect 1106 2496 1112 2497
rect 1266 2501 1272 2502
rect 1266 2497 1267 2501
rect 1271 2497 1272 2501
rect 1266 2496 1272 2497
rect 1426 2501 1432 2502
rect 1426 2497 1427 2501
rect 1431 2497 1432 2501
rect 1426 2496 1432 2497
rect 1586 2501 1592 2502
rect 1586 2497 1587 2501
rect 1591 2497 1592 2501
rect 1586 2496 1592 2497
rect 1754 2501 1760 2502
rect 1754 2497 1755 2501
rect 1759 2497 1760 2501
rect 1754 2496 1760 2497
rect 1934 2500 1940 2501
rect 1934 2496 1935 2500
rect 1939 2496 1940 2500
rect 110 2495 116 2496
rect 112 2423 114 2495
rect 524 2423 526 2496
rect 660 2423 662 2496
rect 804 2423 806 2496
rect 956 2423 958 2496
rect 1108 2423 1110 2496
rect 1268 2423 1270 2496
rect 1428 2423 1430 2496
rect 1588 2423 1590 2496
rect 1756 2423 1758 2496
rect 1934 2495 1940 2496
rect 1936 2423 1938 2495
rect 1976 2475 1978 2551
rect 2484 2475 2486 2552
rect 2620 2475 2622 2552
rect 2756 2475 2758 2552
rect 2892 2475 2894 2552
rect 3028 2475 3030 2552
rect 3164 2475 3166 2552
rect 3300 2475 3302 2552
rect 3436 2475 3438 2552
rect 3798 2551 3804 2552
rect 3800 2475 3802 2551
rect 3840 2538 3842 2561
rect 3838 2537 3844 2538
rect 4496 2537 4498 2561
rect 4632 2537 4634 2561
rect 4768 2537 4770 2561
rect 4904 2537 4906 2561
rect 5040 2537 5042 2561
rect 5664 2538 5666 2561
rect 5662 2537 5668 2538
rect 3838 2533 3839 2537
rect 3843 2533 3844 2537
rect 3838 2532 3844 2533
rect 4494 2536 4500 2537
rect 4494 2532 4495 2536
rect 4499 2532 4500 2536
rect 4494 2531 4500 2532
rect 4630 2536 4636 2537
rect 4630 2532 4631 2536
rect 4635 2532 4636 2536
rect 4630 2531 4636 2532
rect 4766 2536 4772 2537
rect 4766 2532 4767 2536
rect 4771 2532 4772 2536
rect 4766 2531 4772 2532
rect 4902 2536 4908 2537
rect 4902 2532 4903 2536
rect 4907 2532 4908 2536
rect 4902 2531 4908 2532
rect 5038 2536 5044 2537
rect 5038 2532 5039 2536
rect 5043 2532 5044 2536
rect 5662 2533 5663 2537
rect 5667 2533 5668 2537
rect 5662 2532 5668 2533
rect 5038 2531 5044 2532
rect 4466 2521 4472 2522
rect 3838 2520 3844 2521
rect 3838 2516 3839 2520
rect 3843 2516 3844 2520
rect 4466 2517 4467 2521
rect 4471 2517 4472 2521
rect 4466 2516 4472 2517
rect 4602 2521 4608 2522
rect 4602 2517 4603 2521
rect 4607 2517 4608 2521
rect 4602 2516 4608 2517
rect 4738 2521 4744 2522
rect 4738 2517 4739 2521
rect 4743 2517 4744 2521
rect 4738 2516 4744 2517
rect 4874 2521 4880 2522
rect 4874 2517 4875 2521
rect 4879 2517 4880 2521
rect 4874 2516 4880 2517
rect 5010 2521 5016 2522
rect 5010 2517 5011 2521
rect 5015 2517 5016 2521
rect 5010 2516 5016 2517
rect 5662 2520 5668 2521
rect 5662 2516 5663 2520
rect 5667 2516 5668 2520
rect 3838 2515 3844 2516
rect 1975 2474 1979 2475
rect 1975 2469 1979 2470
rect 2307 2474 2311 2475
rect 2307 2469 2311 2470
rect 2483 2474 2487 2475
rect 2483 2469 2487 2470
rect 2515 2474 2519 2475
rect 2515 2469 2519 2470
rect 2619 2474 2623 2475
rect 2619 2469 2623 2470
rect 2715 2474 2719 2475
rect 2715 2469 2719 2470
rect 2755 2474 2759 2475
rect 2755 2469 2759 2470
rect 2891 2474 2895 2475
rect 2891 2469 2895 2470
rect 2907 2474 2911 2475
rect 2907 2469 2911 2470
rect 3027 2474 3031 2475
rect 3027 2469 3031 2470
rect 3099 2474 3103 2475
rect 3099 2469 3103 2470
rect 3163 2474 3167 2475
rect 3163 2469 3167 2470
rect 3283 2474 3287 2475
rect 3283 2469 3287 2470
rect 3299 2474 3303 2475
rect 3299 2469 3303 2470
rect 3435 2474 3439 2475
rect 3435 2469 3439 2470
rect 3467 2474 3471 2475
rect 3467 2469 3471 2470
rect 3651 2474 3655 2475
rect 3651 2469 3655 2470
rect 3799 2474 3803 2475
rect 3799 2469 3803 2470
rect 111 2422 115 2423
rect 111 2417 115 2418
rect 131 2422 135 2423
rect 131 2417 135 2418
rect 339 2422 343 2423
rect 339 2417 343 2418
rect 523 2422 527 2423
rect 523 2417 527 2418
rect 563 2422 567 2423
rect 563 2417 567 2418
rect 659 2422 663 2423
rect 659 2417 663 2418
rect 803 2422 807 2423
rect 803 2417 807 2418
rect 955 2422 959 2423
rect 955 2417 959 2418
rect 1043 2422 1047 2423
rect 1043 2417 1047 2418
rect 1107 2422 1111 2423
rect 1107 2417 1111 2418
rect 1267 2422 1271 2423
rect 1267 2417 1271 2418
rect 1291 2422 1295 2423
rect 1291 2417 1295 2418
rect 1427 2422 1431 2423
rect 1427 2417 1431 2418
rect 1547 2422 1551 2423
rect 1547 2417 1551 2418
rect 1587 2422 1591 2423
rect 1587 2417 1591 2418
rect 1755 2422 1759 2423
rect 1755 2417 1759 2418
rect 1787 2422 1791 2423
rect 1787 2417 1791 2418
rect 1935 2422 1939 2423
rect 1935 2417 1939 2418
rect 112 2357 114 2417
rect 110 2356 116 2357
rect 132 2356 134 2417
rect 340 2356 342 2417
rect 564 2356 566 2417
rect 804 2356 806 2417
rect 1044 2356 1046 2417
rect 1292 2356 1294 2417
rect 1548 2356 1550 2417
rect 1788 2356 1790 2417
rect 1936 2357 1938 2417
rect 1976 2409 1978 2469
rect 1974 2408 1980 2409
rect 2308 2408 2310 2469
rect 2516 2408 2518 2469
rect 2716 2408 2718 2469
rect 2908 2408 2910 2469
rect 3100 2408 3102 2469
rect 3284 2408 3286 2469
rect 3468 2408 3470 2469
rect 3652 2408 3654 2469
rect 3800 2409 3802 2469
rect 3840 2439 3842 2515
rect 4468 2439 4470 2516
rect 4604 2439 4606 2516
rect 4740 2439 4742 2516
rect 4876 2439 4878 2516
rect 5012 2439 5014 2516
rect 5662 2515 5668 2516
rect 5664 2439 5666 2515
rect 3839 2438 3843 2439
rect 3839 2433 3843 2434
rect 4467 2438 4471 2439
rect 4467 2433 4471 2434
rect 4603 2438 4607 2439
rect 4603 2433 4607 2434
rect 4699 2438 4703 2439
rect 4699 2433 4703 2434
rect 4739 2438 4743 2439
rect 4739 2433 4743 2434
rect 4835 2438 4839 2439
rect 4835 2433 4839 2434
rect 4875 2438 4879 2439
rect 4875 2433 4879 2434
rect 4971 2438 4975 2439
rect 4971 2433 4975 2434
rect 5011 2438 5015 2439
rect 5011 2433 5015 2434
rect 5107 2438 5111 2439
rect 5107 2433 5111 2434
rect 5243 2438 5247 2439
rect 5243 2433 5247 2434
rect 5379 2438 5383 2439
rect 5379 2433 5383 2434
rect 5515 2438 5519 2439
rect 5515 2433 5519 2434
rect 5663 2438 5667 2439
rect 5663 2433 5667 2434
rect 3798 2408 3804 2409
rect 1974 2404 1975 2408
rect 1979 2404 1980 2408
rect 1974 2403 1980 2404
rect 2306 2407 2312 2408
rect 2306 2403 2307 2407
rect 2311 2403 2312 2407
rect 2306 2402 2312 2403
rect 2514 2407 2520 2408
rect 2514 2403 2515 2407
rect 2519 2403 2520 2407
rect 2514 2402 2520 2403
rect 2714 2407 2720 2408
rect 2714 2403 2715 2407
rect 2719 2403 2720 2407
rect 2714 2402 2720 2403
rect 2906 2407 2912 2408
rect 2906 2403 2907 2407
rect 2911 2403 2912 2407
rect 2906 2402 2912 2403
rect 3098 2407 3104 2408
rect 3098 2403 3099 2407
rect 3103 2403 3104 2407
rect 3098 2402 3104 2403
rect 3282 2407 3288 2408
rect 3282 2403 3283 2407
rect 3287 2403 3288 2407
rect 3282 2402 3288 2403
rect 3466 2407 3472 2408
rect 3466 2403 3467 2407
rect 3471 2403 3472 2407
rect 3466 2402 3472 2403
rect 3650 2407 3656 2408
rect 3650 2403 3651 2407
rect 3655 2403 3656 2407
rect 3798 2404 3799 2408
rect 3803 2404 3804 2408
rect 3798 2403 3804 2404
rect 3650 2402 3656 2403
rect 2334 2392 2340 2393
rect 1974 2391 1980 2392
rect 1974 2387 1975 2391
rect 1979 2387 1980 2391
rect 2334 2388 2335 2392
rect 2339 2388 2340 2392
rect 2334 2387 2340 2388
rect 2542 2392 2548 2393
rect 2542 2388 2543 2392
rect 2547 2388 2548 2392
rect 2542 2387 2548 2388
rect 2742 2392 2748 2393
rect 2742 2388 2743 2392
rect 2747 2388 2748 2392
rect 2742 2387 2748 2388
rect 2934 2392 2940 2393
rect 2934 2388 2935 2392
rect 2939 2388 2940 2392
rect 2934 2387 2940 2388
rect 3126 2392 3132 2393
rect 3126 2388 3127 2392
rect 3131 2388 3132 2392
rect 3126 2387 3132 2388
rect 3310 2392 3316 2393
rect 3310 2388 3311 2392
rect 3315 2388 3316 2392
rect 3310 2387 3316 2388
rect 3494 2392 3500 2393
rect 3494 2388 3495 2392
rect 3499 2388 3500 2392
rect 3494 2387 3500 2388
rect 3678 2392 3684 2393
rect 3678 2388 3679 2392
rect 3683 2388 3684 2392
rect 3678 2387 3684 2388
rect 3798 2391 3804 2392
rect 3798 2387 3799 2391
rect 3803 2387 3804 2391
rect 1974 2386 1980 2387
rect 1934 2356 1940 2357
rect 110 2352 111 2356
rect 115 2352 116 2356
rect 110 2351 116 2352
rect 130 2355 136 2356
rect 130 2351 131 2355
rect 135 2351 136 2355
rect 130 2350 136 2351
rect 338 2355 344 2356
rect 338 2351 339 2355
rect 343 2351 344 2355
rect 338 2350 344 2351
rect 562 2355 568 2356
rect 562 2351 563 2355
rect 567 2351 568 2355
rect 562 2350 568 2351
rect 802 2355 808 2356
rect 802 2351 803 2355
rect 807 2351 808 2355
rect 802 2350 808 2351
rect 1042 2355 1048 2356
rect 1042 2351 1043 2355
rect 1047 2351 1048 2355
rect 1042 2350 1048 2351
rect 1290 2355 1296 2356
rect 1290 2351 1291 2355
rect 1295 2351 1296 2355
rect 1290 2350 1296 2351
rect 1546 2355 1552 2356
rect 1546 2351 1547 2355
rect 1551 2351 1552 2355
rect 1546 2350 1552 2351
rect 1786 2355 1792 2356
rect 1786 2351 1787 2355
rect 1791 2351 1792 2355
rect 1934 2352 1935 2356
rect 1939 2352 1940 2356
rect 1976 2355 1978 2386
rect 2336 2355 2338 2387
rect 2544 2355 2546 2387
rect 2744 2355 2746 2387
rect 2936 2355 2938 2387
rect 3128 2355 3130 2387
rect 3312 2355 3314 2387
rect 3496 2355 3498 2387
rect 3680 2355 3682 2387
rect 3798 2386 3804 2387
rect 3800 2355 3802 2386
rect 3840 2373 3842 2433
rect 3838 2372 3844 2373
rect 4700 2372 4702 2433
rect 4836 2372 4838 2433
rect 4972 2372 4974 2433
rect 5108 2372 5110 2433
rect 5244 2372 5246 2433
rect 5380 2372 5382 2433
rect 5516 2372 5518 2433
rect 5664 2373 5666 2433
rect 5662 2372 5668 2373
rect 3838 2368 3839 2372
rect 3843 2368 3844 2372
rect 3838 2367 3844 2368
rect 4698 2371 4704 2372
rect 4698 2367 4699 2371
rect 4703 2367 4704 2371
rect 4698 2366 4704 2367
rect 4834 2371 4840 2372
rect 4834 2367 4835 2371
rect 4839 2367 4840 2371
rect 4834 2366 4840 2367
rect 4970 2371 4976 2372
rect 4970 2367 4971 2371
rect 4975 2367 4976 2371
rect 4970 2366 4976 2367
rect 5106 2371 5112 2372
rect 5106 2367 5107 2371
rect 5111 2367 5112 2371
rect 5106 2366 5112 2367
rect 5242 2371 5248 2372
rect 5242 2367 5243 2371
rect 5247 2367 5248 2371
rect 5242 2366 5248 2367
rect 5378 2371 5384 2372
rect 5378 2367 5379 2371
rect 5383 2367 5384 2371
rect 5378 2366 5384 2367
rect 5514 2371 5520 2372
rect 5514 2367 5515 2371
rect 5519 2367 5520 2371
rect 5662 2368 5663 2372
rect 5667 2368 5668 2372
rect 5662 2367 5668 2368
rect 5514 2366 5520 2367
rect 4726 2356 4732 2357
rect 3838 2355 3844 2356
rect 1934 2351 1940 2352
rect 1975 2354 1979 2355
rect 1786 2350 1792 2351
rect 1975 2349 1979 2350
rect 2223 2354 2227 2355
rect 2223 2349 2227 2350
rect 2335 2354 2339 2355
rect 2335 2349 2339 2350
rect 2503 2354 2507 2355
rect 2503 2349 2507 2350
rect 2543 2354 2547 2355
rect 2543 2349 2547 2350
rect 2743 2354 2747 2355
rect 2743 2349 2747 2350
rect 2767 2354 2771 2355
rect 2767 2349 2771 2350
rect 2935 2354 2939 2355
rect 2935 2349 2939 2350
rect 3007 2354 3011 2355
rect 3007 2349 3011 2350
rect 3127 2354 3131 2355
rect 3127 2349 3131 2350
rect 3239 2354 3243 2355
rect 3239 2349 3243 2350
rect 3311 2354 3315 2355
rect 3311 2349 3315 2350
rect 3471 2354 3475 2355
rect 3471 2349 3475 2350
rect 3495 2354 3499 2355
rect 3495 2349 3499 2350
rect 3679 2354 3683 2355
rect 3679 2349 3683 2350
rect 3799 2354 3803 2355
rect 3838 2351 3839 2355
rect 3843 2351 3844 2355
rect 4726 2352 4727 2356
rect 4731 2352 4732 2356
rect 4726 2351 4732 2352
rect 4862 2356 4868 2357
rect 4862 2352 4863 2356
rect 4867 2352 4868 2356
rect 4862 2351 4868 2352
rect 4998 2356 5004 2357
rect 4998 2352 4999 2356
rect 5003 2352 5004 2356
rect 4998 2351 5004 2352
rect 5134 2356 5140 2357
rect 5134 2352 5135 2356
rect 5139 2352 5140 2356
rect 5134 2351 5140 2352
rect 5270 2356 5276 2357
rect 5270 2352 5271 2356
rect 5275 2352 5276 2356
rect 5270 2351 5276 2352
rect 5406 2356 5412 2357
rect 5406 2352 5407 2356
rect 5411 2352 5412 2356
rect 5406 2351 5412 2352
rect 5542 2356 5548 2357
rect 5542 2352 5543 2356
rect 5547 2352 5548 2356
rect 5542 2351 5548 2352
rect 5662 2355 5668 2356
rect 5662 2351 5663 2355
rect 5667 2351 5668 2355
rect 3838 2350 3844 2351
rect 3799 2349 3803 2350
rect 158 2340 164 2341
rect 110 2339 116 2340
rect 110 2335 111 2339
rect 115 2335 116 2339
rect 158 2336 159 2340
rect 163 2336 164 2340
rect 158 2335 164 2336
rect 366 2340 372 2341
rect 366 2336 367 2340
rect 371 2336 372 2340
rect 366 2335 372 2336
rect 590 2340 596 2341
rect 590 2336 591 2340
rect 595 2336 596 2340
rect 590 2335 596 2336
rect 830 2340 836 2341
rect 830 2336 831 2340
rect 835 2336 836 2340
rect 830 2335 836 2336
rect 1070 2340 1076 2341
rect 1070 2336 1071 2340
rect 1075 2336 1076 2340
rect 1070 2335 1076 2336
rect 1318 2340 1324 2341
rect 1318 2336 1319 2340
rect 1323 2336 1324 2340
rect 1318 2335 1324 2336
rect 1574 2340 1580 2341
rect 1574 2336 1575 2340
rect 1579 2336 1580 2340
rect 1574 2335 1580 2336
rect 1814 2340 1820 2341
rect 1814 2336 1815 2340
rect 1819 2336 1820 2340
rect 1814 2335 1820 2336
rect 1934 2339 1940 2340
rect 1934 2335 1935 2339
rect 1939 2335 1940 2339
rect 110 2334 116 2335
rect 112 2307 114 2334
rect 160 2307 162 2335
rect 368 2307 370 2335
rect 592 2307 594 2335
rect 832 2307 834 2335
rect 1072 2307 1074 2335
rect 1320 2307 1322 2335
rect 1576 2307 1578 2335
rect 1816 2307 1818 2335
rect 1934 2334 1940 2335
rect 1936 2307 1938 2334
rect 1976 2326 1978 2349
rect 1974 2325 1980 2326
rect 2224 2325 2226 2349
rect 2504 2325 2506 2349
rect 2768 2325 2770 2349
rect 3008 2325 3010 2349
rect 3240 2325 3242 2349
rect 3472 2325 3474 2349
rect 3680 2325 3682 2349
rect 3800 2326 3802 2349
rect 3798 2325 3804 2326
rect 1974 2321 1975 2325
rect 1979 2321 1980 2325
rect 1974 2320 1980 2321
rect 2222 2324 2228 2325
rect 2222 2320 2223 2324
rect 2227 2320 2228 2324
rect 2222 2319 2228 2320
rect 2502 2324 2508 2325
rect 2502 2320 2503 2324
rect 2507 2320 2508 2324
rect 2502 2319 2508 2320
rect 2766 2324 2772 2325
rect 2766 2320 2767 2324
rect 2771 2320 2772 2324
rect 2766 2319 2772 2320
rect 3006 2324 3012 2325
rect 3006 2320 3007 2324
rect 3011 2320 3012 2324
rect 3006 2319 3012 2320
rect 3238 2324 3244 2325
rect 3238 2320 3239 2324
rect 3243 2320 3244 2324
rect 3238 2319 3244 2320
rect 3470 2324 3476 2325
rect 3470 2320 3471 2324
rect 3475 2320 3476 2324
rect 3470 2319 3476 2320
rect 3678 2324 3684 2325
rect 3678 2320 3679 2324
rect 3683 2320 3684 2324
rect 3798 2321 3799 2325
rect 3803 2321 3804 2325
rect 3798 2320 3804 2321
rect 3678 2319 3684 2320
rect 3840 2315 3842 2350
rect 4728 2315 4730 2351
rect 4864 2315 4866 2351
rect 5000 2315 5002 2351
rect 5136 2315 5138 2351
rect 5272 2315 5274 2351
rect 5408 2315 5410 2351
rect 5544 2315 5546 2351
rect 5662 2350 5668 2351
rect 5664 2315 5666 2350
rect 3839 2314 3843 2315
rect 2194 2309 2200 2310
rect 1974 2308 1980 2309
rect 111 2306 115 2307
rect 111 2301 115 2302
rect 159 2306 163 2307
rect 159 2301 163 2302
rect 319 2306 323 2307
rect 319 2301 323 2302
rect 367 2306 371 2307
rect 367 2301 371 2302
rect 551 2306 555 2307
rect 551 2301 555 2302
rect 591 2306 595 2307
rect 591 2301 595 2302
rect 831 2306 835 2307
rect 831 2301 835 2302
rect 1071 2306 1075 2307
rect 1071 2301 1075 2302
rect 1151 2306 1155 2307
rect 1151 2301 1155 2302
rect 1319 2306 1323 2307
rect 1319 2301 1323 2302
rect 1495 2306 1499 2307
rect 1495 2301 1499 2302
rect 1575 2306 1579 2307
rect 1575 2301 1579 2302
rect 1815 2306 1819 2307
rect 1815 2301 1819 2302
rect 1935 2306 1939 2307
rect 1974 2304 1975 2308
rect 1979 2304 1980 2308
rect 2194 2305 2195 2309
rect 2199 2305 2200 2309
rect 2194 2304 2200 2305
rect 2474 2309 2480 2310
rect 2474 2305 2475 2309
rect 2479 2305 2480 2309
rect 2474 2304 2480 2305
rect 2738 2309 2744 2310
rect 2738 2305 2739 2309
rect 2743 2305 2744 2309
rect 2738 2304 2744 2305
rect 2978 2309 2984 2310
rect 2978 2305 2979 2309
rect 2983 2305 2984 2309
rect 2978 2304 2984 2305
rect 3210 2309 3216 2310
rect 3210 2305 3211 2309
rect 3215 2305 3216 2309
rect 3210 2304 3216 2305
rect 3442 2309 3448 2310
rect 3442 2305 3443 2309
rect 3447 2305 3448 2309
rect 3442 2304 3448 2305
rect 3650 2309 3656 2310
rect 3839 2309 3843 2310
rect 3887 2314 3891 2315
rect 3887 2309 3891 2310
rect 4183 2314 4187 2315
rect 4183 2309 4187 2310
rect 4495 2314 4499 2315
rect 4495 2309 4499 2310
rect 4727 2314 4731 2315
rect 4727 2309 4731 2310
rect 4791 2314 4795 2315
rect 4791 2309 4795 2310
rect 4863 2314 4867 2315
rect 4863 2309 4867 2310
rect 4999 2314 5003 2315
rect 4999 2309 5003 2310
rect 5087 2314 5091 2315
rect 5087 2309 5091 2310
rect 5135 2314 5139 2315
rect 5135 2309 5139 2310
rect 5271 2314 5275 2315
rect 5271 2309 5275 2310
rect 5383 2314 5387 2315
rect 5383 2309 5387 2310
rect 5407 2314 5411 2315
rect 5407 2309 5411 2310
rect 5543 2314 5547 2315
rect 5543 2309 5547 2310
rect 5663 2314 5667 2315
rect 5663 2309 5667 2310
rect 3650 2305 3651 2309
rect 3655 2305 3656 2309
rect 3650 2304 3656 2305
rect 3798 2308 3804 2309
rect 3798 2304 3799 2308
rect 3803 2304 3804 2308
rect 1974 2303 1980 2304
rect 1935 2301 1939 2302
rect 112 2278 114 2301
rect 110 2277 116 2278
rect 160 2277 162 2301
rect 320 2277 322 2301
rect 552 2277 554 2301
rect 832 2277 834 2301
rect 1152 2277 1154 2301
rect 1496 2277 1498 2301
rect 1816 2277 1818 2301
rect 1936 2278 1938 2301
rect 1934 2277 1940 2278
rect 110 2273 111 2277
rect 115 2273 116 2277
rect 110 2272 116 2273
rect 158 2276 164 2277
rect 158 2272 159 2276
rect 163 2272 164 2276
rect 158 2271 164 2272
rect 318 2276 324 2277
rect 318 2272 319 2276
rect 323 2272 324 2276
rect 318 2271 324 2272
rect 550 2276 556 2277
rect 550 2272 551 2276
rect 555 2272 556 2276
rect 550 2271 556 2272
rect 830 2276 836 2277
rect 830 2272 831 2276
rect 835 2272 836 2276
rect 830 2271 836 2272
rect 1150 2276 1156 2277
rect 1150 2272 1151 2276
rect 1155 2272 1156 2276
rect 1150 2271 1156 2272
rect 1494 2276 1500 2277
rect 1494 2272 1495 2276
rect 1499 2272 1500 2276
rect 1494 2271 1500 2272
rect 1814 2276 1820 2277
rect 1814 2272 1815 2276
rect 1819 2272 1820 2276
rect 1934 2273 1935 2277
rect 1939 2273 1940 2277
rect 1934 2272 1940 2273
rect 1814 2271 1820 2272
rect 130 2261 136 2262
rect 110 2260 116 2261
rect 110 2256 111 2260
rect 115 2256 116 2260
rect 130 2257 131 2261
rect 135 2257 136 2261
rect 130 2256 136 2257
rect 290 2261 296 2262
rect 290 2257 291 2261
rect 295 2257 296 2261
rect 290 2256 296 2257
rect 522 2261 528 2262
rect 522 2257 523 2261
rect 527 2257 528 2261
rect 522 2256 528 2257
rect 802 2261 808 2262
rect 802 2257 803 2261
rect 807 2257 808 2261
rect 802 2256 808 2257
rect 1122 2261 1128 2262
rect 1122 2257 1123 2261
rect 1127 2257 1128 2261
rect 1122 2256 1128 2257
rect 1466 2261 1472 2262
rect 1466 2257 1467 2261
rect 1471 2257 1472 2261
rect 1466 2256 1472 2257
rect 1786 2261 1792 2262
rect 1786 2257 1787 2261
rect 1791 2257 1792 2261
rect 1786 2256 1792 2257
rect 1934 2260 1940 2261
rect 1934 2256 1935 2260
rect 1939 2256 1940 2260
rect 110 2255 116 2256
rect 112 2171 114 2255
rect 132 2171 134 2256
rect 292 2171 294 2256
rect 524 2171 526 2256
rect 804 2171 806 2256
rect 1124 2171 1126 2256
rect 1468 2171 1470 2256
rect 1788 2171 1790 2256
rect 1934 2255 1940 2256
rect 1936 2171 1938 2255
rect 1976 2243 1978 2303
rect 2196 2243 2198 2304
rect 2476 2243 2478 2304
rect 2740 2243 2742 2304
rect 2980 2243 2982 2304
rect 3212 2243 3214 2304
rect 3444 2243 3446 2304
rect 3652 2243 3654 2304
rect 3798 2303 3804 2304
rect 3800 2243 3802 2303
rect 3840 2286 3842 2309
rect 3838 2285 3844 2286
rect 3888 2285 3890 2309
rect 4184 2285 4186 2309
rect 4496 2285 4498 2309
rect 4792 2285 4794 2309
rect 5088 2285 5090 2309
rect 5384 2285 5386 2309
rect 5664 2286 5666 2309
rect 5662 2285 5668 2286
rect 3838 2281 3839 2285
rect 3843 2281 3844 2285
rect 3838 2280 3844 2281
rect 3886 2284 3892 2285
rect 3886 2280 3887 2284
rect 3891 2280 3892 2284
rect 3886 2279 3892 2280
rect 4182 2284 4188 2285
rect 4182 2280 4183 2284
rect 4187 2280 4188 2284
rect 4182 2279 4188 2280
rect 4494 2284 4500 2285
rect 4494 2280 4495 2284
rect 4499 2280 4500 2284
rect 4494 2279 4500 2280
rect 4790 2284 4796 2285
rect 4790 2280 4791 2284
rect 4795 2280 4796 2284
rect 4790 2279 4796 2280
rect 5086 2284 5092 2285
rect 5086 2280 5087 2284
rect 5091 2280 5092 2284
rect 5086 2279 5092 2280
rect 5382 2284 5388 2285
rect 5382 2280 5383 2284
rect 5387 2280 5388 2284
rect 5662 2281 5663 2285
rect 5667 2281 5668 2285
rect 5662 2280 5668 2281
rect 5382 2279 5388 2280
rect 3858 2269 3864 2270
rect 3838 2268 3844 2269
rect 3838 2264 3839 2268
rect 3843 2264 3844 2268
rect 3858 2265 3859 2269
rect 3863 2265 3864 2269
rect 3858 2264 3864 2265
rect 4154 2269 4160 2270
rect 4154 2265 4155 2269
rect 4159 2265 4160 2269
rect 4154 2264 4160 2265
rect 4466 2269 4472 2270
rect 4466 2265 4467 2269
rect 4471 2265 4472 2269
rect 4466 2264 4472 2265
rect 4762 2269 4768 2270
rect 4762 2265 4763 2269
rect 4767 2265 4768 2269
rect 4762 2264 4768 2265
rect 5058 2269 5064 2270
rect 5058 2265 5059 2269
rect 5063 2265 5064 2269
rect 5058 2264 5064 2265
rect 5354 2269 5360 2270
rect 5354 2265 5355 2269
rect 5359 2265 5360 2269
rect 5354 2264 5360 2265
rect 5662 2268 5668 2269
rect 5662 2264 5663 2268
rect 5667 2264 5668 2268
rect 3838 2263 3844 2264
rect 1975 2242 1979 2243
rect 1975 2237 1979 2238
rect 1995 2242 1999 2243
rect 1995 2237 1999 2238
rect 2155 2242 2159 2243
rect 2155 2237 2159 2238
rect 2195 2242 2199 2243
rect 2195 2237 2199 2238
rect 2387 2242 2391 2243
rect 2387 2237 2391 2238
rect 2475 2242 2479 2243
rect 2475 2237 2479 2238
rect 2667 2242 2671 2243
rect 2667 2237 2671 2238
rect 2739 2242 2743 2243
rect 2739 2237 2743 2238
rect 2979 2242 2983 2243
rect 2979 2237 2983 2238
rect 2987 2242 2991 2243
rect 2987 2237 2991 2238
rect 3211 2242 3215 2243
rect 3211 2237 3215 2238
rect 3331 2242 3335 2243
rect 3331 2237 3335 2238
rect 3443 2242 3447 2243
rect 3443 2237 3447 2238
rect 3651 2242 3655 2243
rect 3651 2237 3655 2238
rect 3799 2242 3803 2243
rect 3799 2237 3803 2238
rect 1976 2177 1978 2237
rect 1974 2176 1980 2177
rect 1996 2176 1998 2237
rect 2156 2176 2158 2237
rect 2388 2176 2390 2237
rect 2668 2176 2670 2237
rect 2988 2176 2990 2237
rect 3332 2176 3334 2237
rect 3652 2176 3654 2237
rect 3800 2177 3802 2237
rect 3840 2199 3842 2263
rect 3860 2199 3862 2264
rect 4156 2199 4158 2264
rect 4468 2199 4470 2264
rect 4764 2199 4766 2264
rect 5060 2199 5062 2264
rect 5356 2199 5358 2264
rect 5662 2263 5668 2264
rect 5664 2199 5666 2263
rect 3839 2198 3843 2199
rect 3839 2193 3843 2194
rect 3859 2198 3863 2199
rect 3859 2193 3863 2194
rect 3995 2198 3999 2199
rect 3995 2193 3999 2194
rect 4131 2198 4135 2199
rect 4131 2193 4135 2194
rect 4155 2198 4159 2199
rect 4155 2193 4159 2194
rect 4267 2198 4271 2199
rect 4267 2193 4271 2194
rect 4403 2198 4407 2199
rect 4403 2193 4407 2194
rect 4467 2198 4471 2199
rect 4467 2193 4471 2194
rect 4539 2198 4543 2199
rect 4539 2193 4543 2194
rect 4699 2198 4703 2199
rect 4699 2193 4703 2194
rect 4763 2198 4767 2199
rect 4763 2193 4767 2194
rect 4891 2198 4895 2199
rect 4891 2193 4895 2194
rect 5059 2198 5063 2199
rect 5059 2193 5063 2194
rect 5099 2198 5103 2199
rect 5099 2193 5103 2194
rect 5315 2198 5319 2199
rect 5315 2193 5319 2194
rect 5355 2198 5359 2199
rect 5355 2193 5359 2194
rect 5515 2198 5519 2199
rect 5515 2193 5519 2194
rect 5663 2198 5667 2199
rect 5663 2193 5667 2194
rect 3798 2176 3804 2177
rect 1974 2172 1975 2176
rect 1979 2172 1980 2176
rect 1974 2171 1980 2172
rect 1994 2175 2000 2176
rect 1994 2171 1995 2175
rect 1999 2171 2000 2175
rect 111 2170 115 2171
rect 111 2165 115 2166
rect 131 2170 135 2171
rect 131 2165 135 2166
rect 291 2170 295 2171
rect 291 2165 295 2166
rect 483 2170 487 2171
rect 483 2165 487 2166
rect 523 2170 527 2171
rect 523 2165 527 2166
rect 691 2170 695 2171
rect 691 2165 695 2166
rect 803 2170 807 2171
rect 803 2165 807 2166
rect 915 2170 919 2171
rect 915 2165 919 2166
rect 1123 2170 1127 2171
rect 1123 2165 1127 2166
rect 1147 2170 1151 2171
rect 1147 2165 1151 2166
rect 1387 2170 1391 2171
rect 1387 2165 1391 2166
rect 1467 2170 1471 2171
rect 1467 2165 1471 2166
rect 1635 2170 1639 2171
rect 1635 2165 1639 2166
rect 1787 2170 1791 2171
rect 1787 2165 1791 2166
rect 1935 2170 1939 2171
rect 1994 2170 2000 2171
rect 2154 2175 2160 2176
rect 2154 2171 2155 2175
rect 2159 2171 2160 2175
rect 2154 2170 2160 2171
rect 2386 2175 2392 2176
rect 2386 2171 2387 2175
rect 2391 2171 2392 2175
rect 2386 2170 2392 2171
rect 2666 2175 2672 2176
rect 2666 2171 2667 2175
rect 2671 2171 2672 2175
rect 2666 2170 2672 2171
rect 2986 2175 2992 2176
rect 2986 2171 2987 2175
rect 2991 2171 2992 2175
rect 2986 2170 2992 2171
rect 3330 2175 3336 2176
rect 3330 2171 3331 2175
rect 3335 2171 3336 2175
rect 3330 2170 3336 2171
rect 3650 2175 3656 2176
rect 3650 2171 3651 2175
rect 3655 2171 3656 2175
rect 3798 2172 3799 2176
rect 3803 2172 3804 2176
rect 3798 2171 3804 2172
rect 3650 2170 3656 2171
rect 1935 2165 1939 2166
rect 112 2105 114 2165
rect 110 2104 116 2105
rect 292 2104 294 2165
rect 484 2104 486 2165
rect 692 2104 694 2165
rect 916 2104 918 2165
rect 1148 2104 1150 2165
rect 1388 2104 1390 2165
rect 1636 2104 1638 2165
rect 1936 2105 1938 2165
rect 2022 2160 2028 2161
rect 1974 2159 1980 2160
rect 1974 2155 1975 2159
rect 1979 2155 1980 2159
rect 2022 2156 2023 2160
rect 2027 2156 2028 2160
rect 2022 2155 2028 2156
rect 2182 2160 2188 2161
rect 2182 2156 2183 2160
rect 2187 2156 2188 2160
rect 2182 2155 2188 2156
rect 2414 2160 2420 2161
rect 2414 2156 2415 2160
rect 2419 2156 2420 2160
rect 2414 2155 2420 2156
rect 2694 2160 2700 2161
rect 2694 2156 2695 2160
rect 2699 2156 2700 2160
rect 2694 2155 2700 2156
rect 3014 2160 3020 2161
rect 3014 2156 3015 2160
rect 3019 2156 3020 2160
rect 3014 2155 3020 2156
rect 3358 2160 3364 2161
rect 3358 2156 3359 2160
rect 3363 2156 3364 2160
rect 3358 2155 3364 2156
rect 3678 2160 3684 2161
rect 3678 2156 3679 2160
rect 3683 2156 3684 2160
rect 3678 2155 3684 2156
rect 3798 2159 3804 2160
rect 3798 2155 3799 2159
rect 3803 2155 3804 2159
rect 1974 2154 1980 2155
rect 1934 2104 1940 2105
rect 110 2100 111 2104
rect 115 2100 116 2104
rect 110 2099 116 2100
rect 290 2103 296 2104
rect 290 2099 291 2103
rect 295 2099 296 2103
rect 290 2098 296 2099
rect 482 2103 488 2104
rect 482 2099 483 2103
rect 487 2099 488 2103
rect 482 2098 488 2099
rect 690 2103 696 2104
rect 690 2099 691 2103
rect 695 2099 696 2103
rect 690 2098 696 2099
rect 914 2103 920 2104
rect 914 2099 915 2103
rect 919 2099 920 2103
rect 914 2098 920 2099
rect 1146 2103 1152 2104
rect 1146 2099 1147 2103
rect 1151 2099 1152 2103
rect 1146 2098 1152 2099
rect 1386 2103 1392 2104
rect 1386 2099 1387 2103
rect 1391 2099 1392 2103
rect 1386 2098 1392 2099
rect 1634 2103 1640 2104
rect 1634 2099 1635 2103
rect 1639 2099 1640 2103
rect 1934 2100 1935 2104
rect 1939 2100 1940 2104
rect 1934 2099 1940 2100
rect 1634 2098 1640 2099
rect 318 2088 324 2089
rect 110 2087 116 2088
rect 110 2083 111 2087
rect 115 2083 116 2087
rect 318 2084 319 2088
rect 323 2084 324 2088
rect 318 2083 324 2084
rect 510 2088 516 2089
rect 510 2084 511 2088
rect 515 2084 516 2088
rect 510 2083 516 2084
rect 718 2088 724 2089
rect 718 2084 719 2088
rect 723 2084 724 2088
rect 718 2083 724 2084
rect 942 2088 948 2089
rect 942 2084 943 2088
rect 947 2084 948 2088
rect 942 2083 948 2084
rect 1174 2088 1180 2089
rect 1174 2084 1175 2088
rect 1179 2084 1180 2088
rect 1174 2083 1180 2084
rect 1414 2088 1420 2089
rect 1414 2084 1415 2088
rect 1419 2084 1420 2088
rect 1414 2083 1420 2084
rect 1662 2088 1668 2089
rect 1662 2084 1663 2088
rect 1667 2084 1668 2088
rect 1662 2083 1668 2084
rect 1934 2087 1940 2088
rect 1934 2083 1935 2087
rect 1939 2083 1940 2087
rect 110 2082 116 2083
rect 112 2055 114 2082
rect 320 2055 322 2083
rect 512 2055 514 2083
rect 720 2055 722 2083
rect 944 2055 946 2083
rect 1176 2055 1178 2083
rect 1416 2055 1418 2083
rect 1664 2055 1666 2083
rect 1934 2082 1940 2083
rect 1936 2055 1938 2082
rect 111 2054 115 2055
rect 111 2049 115 2050
rect 263 2054 267 2055
rect 263 2049 267 2050
rect 319 2054 323 2055
rect 319 2049 323 2050
rect 399 2054 403 2055
rect 399 2049 403 2050
rect 511 2054 515 2055
rect 511 2049 515 2050
rect 535 2054 539 2055
rect 535 2049 539 2050
rect 679 2054 683 2055
rect 679 2049 683 2050
rect 719 2054 723 2055
rect 719 2049 723 2050
rect 823 2054 827 2055
rect 823 2049 827 2050
rect 943 2054 947 2055
rect 943 2049 947 2050
rect 967 2054 971 2055
rect 967 2049 971 2050
rect 1111 2054 1115 2055
rect 1111 2049 1115 2050
rect 1175 2054 1179 2055
rect 1175 2049 1179 2050
rect 1255 2054 1259 2055
rect 1255 2049 1259 2050
rect 1399 2054 1403 2055
rect 1399 2049 1403 2050
rect 1415 2054 1419 2055
rect 1415 2049 1419 2050
rect 1543 2054 1547 2055
rect 1543 2049 1547 2050
rect 1663 2054 1667 2055
rect 1663 2049 1667 2050
rect 1679 2054 1683 2055
rect 1679 2049 1683 2050
rect 1815 2054 1819 2055
rect 1815 2049 1819 2050
rect 1935 2054 1939 2055
rect 1935 2049 1939 2050
rect 112 2026 114 2049
rect 110 2025 116 2026
rect 264 2025 266 2049
rect 400 2025 402 2049
rect 536 2025 538 2049
rect 680 2025 682 2049
rect 824 2025 826 2049
rect 968 2025 970 2049
rect 1112 2025 1114 2049
rect 1256 2025 1258 2049
rect 1400 2025 1402 2049
rect 1544 2025 1546 2049
rect 1680 2025 1682 2049
rect 1816 2025 1818 2049
rect 1936 2026 1938 2049
rect 1934 2025 1940 2026
rect 110 2021 111 2025
rect 115 2021 116 2025
rect 110 2020 116 2021
rect 262 2024 268 2025
rect 262 2020 263 2024
rect 267 2020 268 2024
rect 262 2019 268 2020
rect 398 2024 404 2025
rect 398 2020 399 2024
rect 403 2020 404 2024
rect 398 2019 404 2020
rect 534 2024 540 2025
rect 534 2020 535 2024
rect 539 2020 540 2024
rect 534 2019 540 2020
rect 678 2024 684 2025
rect 678 2020 679 2024
rect 683 2020 684 2024
rect 678 2019 684 2020
rect 822 2024 828 2025
rect 822 2020 823 2024
rect 827 2020 828 2024
rect 822 2019 828 2020
rect 966 2024 972 2025
rect 966 2020 967 2024
rect 971 2020 972 2024
rect 966 2019 972 2020
rect 1110 2024 1116 2025
rect 1110 2020 1111 2024
rect 1115 2020 1116 2024
rect 1110 2019 1116 2020
rect 1254 2024 1260 2025
rect 1254 2020 1255 2024
rect 1259 2020 1260 2024
rect 1254 2019 1260 2020
rect 1398 2024 1404 2025
rect 1398 2020 1399 2024
rect 1403 2020 1404 2024
rect 1398 2019 1404 2020
rect 1542 2024 1548 2025
rect 1542 2020 1543 2024
rect 1547 2020 1548 2024
rect 1542 2019 1548 2020
rect 1678 2024 1684 2025
rect 1678 2020 1679 2024
rect 1683 2020 1684 2024
rect 1678 2019 1684 2020
rect 1814 2024 1820 2025
rect 1814 2020 1815 2024
rect 1819 2020 1820 2024
rect 1934 2021 1935 2025
rect 1939 2021 1940 2025
rect 1934 2020 1940 2021
rect 1814 2019 1820 2020
rect 234 2009 240 2010
rect 110 2008 116 2009
rect 110 2004 111 2008
rect 115 2004 116 2008
rect 234 2005 235 2009
rect 239 2005 240 2009
rect 234 2004 240 2005
rect 370 2009 376 2010
rect 370 2005 371 2009
rect 375 2005 376 2009
rect 370 2004 376 2005
rect 506 2009 512 2010
rect 506 2005 507 2009
rect 511 2005 512 2009
rect 506 2004 512 2005
rect 650 2009 656 2010
rect 650 2005 651 2009
rect 655 2005 656 2009
rect 650 2004 656 2005
rect 794 2009 800 2010
rect 794 2005 795 2009
rect 799 2005 800 2009
rect 794 2004 800 2005
rect 938 2009 944 2010
rect 938 2005 939 2009
rect 943 2005 944 2009
rect 938 2004 944 2005
rect 1082 2009 1088 2010
rect 1082 2005 1083 2009
rect 1087 2005 1088 2009
rect 1082 2004 1088 2005
rect 1226 2009 1232 2010
rect 1226 2005 1227 2009
rect 1231 2005 1232 2009
rect 1226 2004 1232 2005
rect 1370 2009 1376 2010
rect 1370 2005 1371 2009
rect 1375 2005 1376 2009
rect 1370 2004 1376 2005
rect 1514 2009 1520 2010
rect 1514 2005 1515 2009
rect 1519 2005 1520 2009
rect 1514 2004 1520 2005
rect 1650 2009 1656 2010
rect 1650 2005 1651 2009
rect 1655 2005 1656 2009
rect 1650 2004 1656 2005
rect 1786 2009 1792 2010
rect 1786 2005 1787 2009
rect 1791 2005 1792 2009
rect 1786 2004 1792 2005
rect 1934 2008 1940 2009
rect 1934 2004 1935 2008
rect 1939 2004 1940 2008
rect 110 2003 116 2004
rect 112 1931 114 2003
rect 236 1931 238 2004
rect 372 1931 374 2004
rect 508 1931 510 2004
rect 652 1931 654 2004
rect 796 1931 798 2004
rect 940 1931 942 2004
rect 1084 1931 1086 2004
rect 1228 1931 1230 2004
rect 1372 1931 1374 2004
rect 1516 1931 1518 2004
rect 1652 1931 1654 2004
rect 1788 1931 1790 2004
rect 1934 2003 1940 2004
rect 1936 1931 1938 2003
rect 1976 1931 1978 2154
rect 2024 1931 2026 2155
rect 2184 1931 2186 2155
rect 2416 1931 2418 2155
rect 2696 1931 2698 2155
rect 3016 1931 3018 2155
rect 3360 1931 3362 2155
rect 3680 1931 3682 2155
rect 3798 2154 3804 2155
rect 3800 1931 3802 2154
rect 3840 2133 3842 2193
rect 3838 2132 3844 2133
rect 3860 2132 3862 2193
rect 3996 2132 3998 2193
rect 4132 2132 4134 2193
rect 4268 2132 4270 2193
rect 4404 2132 4406 2193
rect 4540 2132 4542 2193
rect 4700 2132 4702 2193
rect 4892 2132 4894 2193
rect 5100 2132 5102 2193
rect 5316 2132 5318 2193
rect 5516 2132 5518 2193
rect 5664 2133 5666 2193
rect 5662 2132 5668 2133
rect 3838 2128 3839 2132
rect 3843 2128 3844 2132
rect 3838 2127 3844 2128
rect 3858 2131 3864 2132
rect 3858 2127 3859 2131
rect 3863 2127 3864 2131
rect 3858 2126 3864 2127
rect 3994 2131 4000 2132
rect 3994 2127 3995 2131
rect 3999 2127 4000 2131
rect 3994 2126 4000 2127
rect 4130 2131 4136 2132
rect 4130 2127 4131 2131
rect 4135 2127 4136 2131
rect 4130 2126 4136 2127
rect 4266 2131 4272 2132
rect 4266 2127 4267 2131
rect 4271 2127 4272 2131
rect 4266 2126 4272 2127
rect 4402 2131 4408 2132
rect 4402 2127 4403 2131
rect 4407 2127 4408 2131
rect 4402 2126 4408 2127
rect 4538 2131 4544 2132
rect 4538 2127 4539 2131
rect 4543 2127 4544 2131
rect 4538 2126 4544 2127
rect 4698 2131 4704 2132
rect 4698 2127 4699 2131
rect 4703 2127 4704 2131
rect 4698 2126 4704 2127
rect 4890 2131 4896 2132
rect 4890 2127 4891 2131
rect 4895 2127 4896 2131
rect 4890 2126 4896 2127
rect 5098 2131 5104 2132
rect 5098 2127 5099 2131
rect 5103 2127 5104 2131
rect 5098 2126 5104 2127
rect 5314 2131 5320 2132
rect 5314 2127 5315 2131
rect 5319 2127 5320 2131
rect 5314 2126 5320 2127
rect 5514 2131 5520 2132
rect 5514 2127 5515 2131
rect 5519 2127 5520 2131
rect 5662 2128 5663 2132
rect 5667 2128 5668 2132
rect 5662 2127 5668 2128
rect 5514 2126 5520 2127
rect 3886 2116 3892 2117
rect 3838 2115 3844 2116
rect 3838 2111 3839 2115
rect 3843 2111 3844 2115
rect 3886 2112 3887 2116
rect 3891 2112 3892 2116
rect 3886 2111 3892 2112
rect 4022 2116 4028 2117
rect 4022 2112 4023 2116
rect 4027 2112 4028 2116
rect 4022 2111 4028 2112
rect 4158 2116 4164 2117
rect 4158 2112 4159 2116
rect 4163 2112 4164 2116
rect 4158 2111 4164 2112
rect 4294 2116 4300 2117
rect 4294 2112 4295 2116
rect 4299 2112 4300 2116
rect 4294 2111 4300 2112
rect 4430 2116 4436 2117
rect 4430 2112 4431 2116
rect 4435 2112 4436 2116
rect 4430 2111 4436 2112
rect 4566 2116 4572 2117
rect 4566 2112 4567 2116
rect 4571 2112 4572 2116
rect 4566 2111 4572 2112
rect 4726 2116 4732 2117
rect 4726 2112 4727 2116
rect 4731 2112 4732 2116
rect 4726 2111 4732 2112
rect 4918 2116 4924 2117
rect 4918 2112 4919 2116
rect 4923 2112 4924 2116
rect 4918 2111 4924 2112
rect 5126 2116 5132 2117
rect 5126 2112 5127 2116
rect 5131 2112 5132 2116
rect 5126 2111 5132 2112
rect 5342 2116 5348 2117
rect 5342 2112 5343 2116
rect 5347 2112 5348 2116
rect 5342 2111 5348 2112
rect 5542 2116 5548 2117
rect 5542 2112 5543 2116
rect 5547 2112 5548 2116
rect 5542 2111 5548 2112
rect 5662 2115 5668 2116
rect 5662 2111 5663 2115
rect 5667 2111 5668 2115
rect 3838 2110 3844 2111
rect 3840 2067 3842 2110
rect 3888 2067 3890 2111
rect 4024 2067 4026 2111
rect 4160 2067 4162 2111
rect 4296 2067 4298 2111
rect 4432 2067 4434 2111
rect 4568 2067 4570 2111
rect 4728 2067 4730 2111
rect 4920 2067 4922 2111
rect 5128 2067 5130 2111
rect 5344 2067 5346 2111
rect 5544 2067 5546 2111
rect 5662 2110 5668 2111
rect 5664 2067 5666 2110
rect 3839 2066 3843 2067
rect 3839 2061 3843 2062
rect 3887 2066 3891 2067
rect 3887 2061 3891 2062
rect 4023 2066 4027 2067
rect 4023 2061 4027 2062
rect 4159 2066 4163 2067
rect 4159 2061 4163 2062
rect 4295 2066 4299 2067
rect 4295 2061 4299 2062
rect 4431 2066 4435 2067
rect 4431 2061 4435 2062
rect 4567 2066 4571 2067
rect 4567 2061 4571 2062
rect 4719 2066 4723 2067
rect 4719 2061 4723 2062
rect 4727 2066 4731 2067
rect 4727 2061 4731 2062
rect 4895 2066 4899 2067
rect 4895 2061 4899 2062
rect 4919 2066 4923 2067
rect 4919 2061 4923 2062
rect 5087 2066 5091 2067
rect 5087 2061 5091 2062
rect 5127 2066 5131 2067
rect 5127 2061 5131 2062
rect 5279 2066 5283 2067
rect 5279 2061 5283 2062
rect 5343 2066 5347 2067
rect 5343 2061 5347 2062
rect 5479 2066 5483 2067
rect 5479 2061 5483 2062
rect 5543 2066 5547 2067
rect 5543 2061 5547 2062
rect 5663 2066 5667 2067
rect 5663 2061 5667 2062
rect 3840 2038 3842 2061
rect 3838 2037 3844 2038
rect 3888 2037 3890 2061
rect 4024 2037 4026 2061
rect 4160 2037 4162 2061
rect 4296 2037 4298 2061
rect 4432 2037 4434 2061
rect 4568 2037 4570 2061
rect 4720 2037 4722 2061
rect 4896 2037 4898 2061
rect 5088 2037 5090 2061
rect 5280 2037 5282 2061
rect 5480 2037 5482 2061
rect 5664 2038 5666 2061
rect 5662 2037 5668 2038
rect 3838 2033 3839 2037
rect 3843 2033 3844 2037
rect 3838 2032 3844 2033
rect 3886 2036 3892 2037
rect 3886 2032 3887 2036
rect 3891 2032 3892 2036
rect 3886 2031 3892 2032
rect 4022 2036 4028 2037
rect 4022 2032 4023 2036
rect 4027 2032 4028 2036
rect 4022 2031 4028 2032
rect 4158 2036 4164 2037
rect 4158 2032 4159 2036
rect 4163 2032 4164 2036
rect 4158 2031 4164 2032
rect 4294 2036 4300 2037
rect 4294 2032 4295 2036
rect 4299 2032 4300 2036
rect 4294 2031 4300 2032
rect 4430 2036 4436 2037
rect 4430 2032 4431 2036
rect 4435 2032 4436 2036
rect 4430 2031 4436 2032
rect 4566 2036 4572 2037
rect 4566 2032 4567 2036
rect 4571 2032 4572 2036
rect 4566 2031 4572 2032
rect 4718 2036 4724 2037
rect 4718 2032 4719 2036
rect 4723 2032 4724 2036
rect 4718 2031 4724 2032
rect 4894 2036 4900 2037
rect 4894 2032 4895 2036
rect 4899 2032 4900 2036
rect 4894 2031 4900 2032
rect 5086 2036 5092 2037
rect 5086 2032 5087 2036
rect 5091 2032 5092 2036
rect 5086 2031 5092 2032
rect 5278 2036 5284 2037
rect 5278 2032 5279 2036
rect 5283 2032 5284 2036
rect 5278 2031 5284 2032
rect 5478 2036 5484 2037
rect 5478 2032 5479 2036
rect 5483 2032 5484 2036
rect 5662 2033 5663 2037
rect 5667 2033 5668 2037
rect 5662 2032 5668 2033
rect 5478 2031 5484 2032
rect 3858 2021 3864 2022
rect 3838 2020 3844 2021
rect 3838 2016 3839 2020
rect 3843 2016 3844 2020
rect 3858 2017 3859 2021
rect 3863 2017 3864 2021
rect 3858 2016 3864 2017
rect 3994 2021 4000 2022
rect 3994 2017 3995 2021
rect 3999 2017 4000 2021
rect 3994 2016 4000 2017
rect 4130 2021 4136 2022
rect 4130 2017 4131 2021
rect 4135 2017 4136 2021
rect 4130 2016 4136 2017
rect 4266 2021 4272 2022
rect 4266 2017 4267 2021
rect 4271 2017 4272 2021
rect 4266 2016 4272 2017
rect 4402 2021 4408 2022
rect 4402 2017 4403 2021
rect 4407 2017 4408 2021
rect 4402 2016 4408 2017
rect 4538 2021 4544 2022
rect 4538 2017 4539 2021
rect 4543 2017 4544 2021
rect 4538 2016 4544 2017
rect 4690 2021 4696 2022
rect 4690 2017 4691 2021
rect 4695 2017 4696 2021
rect 4690 2016 4696 2017
rect 4866 2021 4872 2022
rect 4866 2017 4867 2021
rect 4871 2017 4872 2021
rect 4866 2016 4872 2017
rect 5058 2021 5064 2022
rect 5058 2017 5059 2021
rect 5063 2017 5064 2021
rect 5058 2016 5064 2017
rect 5250 2021 5256 2022
rect 5250 2017 5251 2021
rect 5255 2017 5256 2021
rect 5250 2016 5256 2017
rect 5450 2021 5456 2022
rect 5450 2017 5451 2021
rect 5455 2017 5456 2021
rect 5450 2016 5456 2017
rect 5662 2020 5668 2021
rect 5662 2016 5663 2020
rect 5667 2016 5668 2020
rect 3838 2015 3844 2016
rect 3840 1955 3842 2015
rect 3860 1955 3862 2016
rect 3996 1955 3998 2016
rect 4132 1955 4134 2016
rect 4268 1955 4270 2016
rect 4404 1955 4406 2016
rect 4540 1955 4542 2016
rect 4692 1955 4694 2016
rect 4868 1955 4870 2016
rect 5060 1955 5062 2016
rect 5252 1955 5254 2016
rect 5452 1955 5454 2016
rect 5662 2015 5668 2016
rect 5664 1955 5666 2015
rect 3839 1954 3843 1955
rect 3839 1949 3843 1950
rect 3859 1954 3863 1955
rect 3859 1949 3863 1950
rect 3995 1954 3999 1955
rect 3995 1949 3999 1950
rect 4043 1954 4047 1955
rect 4043 1949 4047 1950
rect 4131 1954 4135 1955
rect 4131 1949 4135 1950
rect 4267 1954 4271 1955
rect 4267 1949 4271 1950
rect 4283 1954 4287 1955
rect 4283 1949 4287 1950
rect 4403 1954 4407 1955
rect 4403 1949 4407 1950
rect 4539 1954 4543 1955
rect 4539 1949 4543 1950
rect 4563 1954 4567 1955
rect 4563 1949 4567 1950
rect 4691 1954 4695 1955
rect 4691 1949 4695 1950
rect 4867 1954 4871 1955
rect 4867 1949 4871 1950
rect 4875 1954 4879 1955
rect 4875 1949 4879 1950
rect 5059 1954 5063 1955
rect 5059 1949 5063 1950
rect 5203 1954 5207 1955
rect 5203 1949 5207 1950
rect 5251 1954 5255 1955
rect 5251 1949 5255 1950
rect 5451 1954 5455 1955
rect 5451 1949 5455 1950
rect 5515 1954 5519 1955
rect 5515 1949 5519 1950
rect 5663 1954 5667 1955
rect 5663 1949 5667 1950
rect 111 1930 115 1931
rect 111 1925 115 1926
rect 235 1930 239 1931
rect 235 1925 239 1926
rect 371 1930 375 1931
rect 371 1925 375 1926
rect 435 1930 439 1931
rect 435 1925 439 1926
rect 507 1930 511 1931
rect 507 1925 511 1926
rect 627 1930 631 1931
rect 627 1925 631 1926
rect 651 1930 655 1931
rect 651 1925 655 1926
rect 795 1930 799 1931
rect 795 1925 799 1926
rect 811 1930 815 1931
rect 811 1925 815 1926
rect 939 1930 943 1931
rect 939 1925 943 1926
rect 987 1930 991 1931
rect 987 1925 991 1926
rect 1083 1930 1087 1931
rect 1083 1925 1087 1926
rect 1155 1930 1159 1931
rect 1155 1925 1159 1926
rect 1227 1930 1231 1931
rect 1227 1925 1231 1926
rect 1323 1930 1327 1931
rect 1323 1925 1327 1926
rect 1371 1930 1375 1931
rect 1371 1925 1375 1926
rect 1483 1930 1487 1931
rect 1483 1925 1487 1926
rect 1515 1930 1519 1931
rect 1515 1925 1519 1926
rect 1643 1930 1647 1931
rect 1643 1925 1647 1926
rect 1651 1930 1655 1931
rect 1651 1925 1655 1926
rect 1787 1930 1791 1931
rect 1787 1925 1791 1926
rect 1935 1930 1939 1931
rect 1935 1925 1939 1926
rect 1975 1930 1979 1931
rect 1975 1925 1979 1926
rect 2023 1930 2027 1931
rect 2023 1925 2027 1926
rect 2183 1930 2187 1931
rect 2183 1925 2187 1926
rect 2415 1930 2419 1931
rect 2415 1925 2419 1926
rect 2695 1930 2699 1931
rect 2695 1925 2699 1926
rect 3015 1930 3019 1931
rect 3015 1925 3019 1926
rect 3135 1930 3139 1931
rect 3135 1925 3139 1926
rect 3271 1930 3275 1931
rect 3271 1925 3275 1926
rect 3359 1930 3363 1931
rect 3359 1925 3363 1926
rect 3407 1930 3411 1931
rect 3407 1925 3411 1926
rect 3543 1930 3547 1931
rect 3543 1925 3547 1926
rect 3679 1930 3683 1931
rect 3679 1925 3683 1926
rect 3799 1930 3803 1931
rect 3799 1925 3803 1926
rect 112 1865 114 1925
rect 110 1864 116 1865
rect 236 1864 238 1925
rect 436 1864 438 1925
rect 628 1864 630 1925
rect 812 1864 814 1925
rect 988 1864 990 1925
rect 1156 1864 1158 1925
rect 1324 1864 1326 1925
rect 1484 1864 1486 1925
rect 1644 1864 1646 1925
rect 1788 1864 1790 1925
rect 1936 1865 1938 1925
rect 1976 1902 1978 1925
rect 1974 1901 1980 1902
rect 3136 1901 3138 1925
rect 3272 1901 3274 1925
rect 3408 1901 3410 1925
rect 3544 1901 3546 1925
rect 3680 1901 3682 1925
rect 3800 1902 3802 1925
rect 3798 1901 3804 1902
rect 1974 1897 1975 1901
rect 1979 1897 1980 1901
rect 1974 1896 1980 1897
rect 3134 1900 3140 1901
rect 3134 1896 3135 1900
rect 3139 1896 3140 1900
rect 3134 1895 3140 1896
rect 3270 1900 3276 1901
rect 3270 1896 3271 1900
rect 3275 1896 3276 1900
rect 3270 1895 3276 1896
rect 3406 1900 3412 1901
rect 3406 1896 3407 1900
rect 3411 1896 3412 1900
rect 3406 1895 3412 1896
rect 3542 1900 3548 1901
rect 3542 1896 3543 1900
rect 3547 1896 3548 1900
rect 3542 1895 3548 1896
rect 3678 1900 3684 1901
rect 3678 1896 3679 1900
rect 3683 1896 3684 1900
rect 3798 1897 3799 1901
rect 3803 1897 3804 1901
rect 3798 1896 3804 1897
rect 3678 1895 3684 1896
rect 3840 1889 3842 1949
rect 3838 1888 3844 1889
rect 3860 1888 3862 1949
rect 4044 1888 4046 1949
rect 4284 1888 4286 1949
rect 4564 1888 4566 1949
rect 4876 1888 4878 1949
rect 5204 1888 5206 1949
rect 5516 1888 5518 1949
rect 5664 1889 5666 1949
rect 5662 1888 5668 1889
rect 3106 1885 3112 1886
rect 1974 1884 1980 1885
rect 1974 1880 1975 1884
rect 1979 1880 1980 1884
rect 3106 1881 3107 1885
rect 3111 1881 3112 1885
rect 3106 1880 3112 1881
rect 3242 1885 3248 1886
rect 3242 1881 3243 1885
rect 3247 1881 3248 1885
rect 3242 1880 3248 1881
rect 3378 1885 3384 1886
rect 3378 1881 3379 1885
rect 3383 1881 3384 1885
rect 3378 1880 3384 1881
rect 3514 1885 3520 1886
rect 3514 1881 3515 1885
rect 3519 1881 3520 1885
rect 3514 1880 3520 1881
rect 3650 1885 3656 1886
rect 3650 1881 3651 1885
rect 3655 1881 3656 1885
rect 3650 1880 3656 1881
rect 3798 1884 3804 1885
rect 3798 1880 3799 1884
rect 3803 1880 3804 1884
rect 3838 1884 3839 1888
rect 3843 1884 3844 1888
rect 3838 1883 3844 1884
rect 3858 1887 3864 1888
rect 3858 1883 3859 1887
rect 3863 1883 3864 1887
rect 3858 1882 3864 1883
rect 4042 1887 4048 1888
rect 4042 1883 4043 1887
rect 4047 1883 4048 1887
rect 4042 1882 4048 1883
rect 4282 1887 4288 1888
rect 4282 1883 4283 1887
rect 4287 1883 4288 1887
rect 4282 1882 4288 1883
rect 4562 1887 4568 1888
rect 4562 1883 4563 1887
rect 4567 1883 4568 1887
rect 4562 1882 4568 1883
rect 4874 1887 4880 1888
rect 4874 1883 4875 1887
rect 4879 1883 4880 1887
rect 4874 1882 4880 1883
rect 5202 1887 5208 1888
rect 5202 1883 5203 1887
rect 5207 1883 5208 1887
rect 5202 1882 5208 1883
rect 5514 1887 5520 1888
rect 5514 1883 5515 1887
rect 5519 1883 5520 1887
rect 5662 1884 5663 1888
rect 5667 1884 5668 1888
rect 5662 1883 5668 1884
rect 5514 1882 5520 1883
rect 1974 1879 1980 1880
rect 1934 1864 1940 1865
rect 110 1860 111 1864
rect 115 1860 116 1864
rect 110 1859 116 1860
rect 234 1863 240 1864
rect 234 1859 235 1863
rect 239 1859 240 1863
rect 234 1858 240 1859
rect 434 1863 440 1864
rect 434 1859 435 1863
rect 439 1859 440 1863
rect 434 1858 440 1859
rect 626 1863 632 1864
rect 626 1859 627 1863
rect 631 1859 632 1863
rect 626 1858 632 1859
rect 810 1863 816 1864
rect 810 1859 811 1863
rect 815 1859 816 1863
rect 810 1858 816 1859
rect 986 1863 992 1864
rect 986 1859 987 1863
rect 991 1859 992 1863
rect 986 1858 992 1859
rect 1154 1863 1160 1864
rect 1154 1859 1155 1863
rect 1159 1859 1160 1863
rect 1154 1858 1160 1859
rect 1322 1863 1328 1864
rect 1322 1859 1323 1863
rect 1327 1859 1328 1863
rect 1322 1858 1328 1859
rect 1482 1863 1488 1864
rect 1482 1859 1483 1863
rect 1487 1859 1488 1863
rect 1482 1858 1488 1859
rect 1642 1863 1648 1864
rect 1642 1859 1643 1863
rect 1647 1859 1648 1863
rect 1642 1858 1648 1859
rect 1786 1863 1792 1864
rect 1786 1859 1787 1863
rect 1791 1859 1792 1863
rect 1934 1860 1935 1864
rect 1939 1860 1940 1864
rect 1934 1859 1940 1860
rect 1786 1858 1792 1859
rect 262 1848 268 1849
rect 110 1847 116 1848
rect 110 1843 111 1847
rect 115 1843 116 1847
rect 262 1844 263 1848
rect 267 1844 268 1848
rect 262 1843 268 1844
rect 462 1848 468 1849
rect 462 1844 463 1848
rect 467 1844 468 1848
rect 462 1843 468 1844
rect 654 1848 660 1849
rect 654 1844 655 1848
rect 659 1844 660 1848
rect 654 1843 660 1844
rect 838 1848 844 1849
rect 838 1844 839 1848
rect 843 1844 844 1848
rect 838 1843 844 1844
rect 1014 1848 1020 1849
rect 1014 1844 1015 1848
rect 1019 1844 1020 1848
rect 1014 1843 1020 1844
rect 1182 1848 1188 1849
rect 1182 1844 1183 1848
rect 1187 1844 1188 1848
rect 1182 1843 1188 1844
rect 1350 1848 1356 1849
rect 1350 1844 1351 1848
rect 1355 1844 1356 1848
rect 1350 1843 1356 1844
rect 1510 1848 1516 1849
rect 1510 1844 1511 1848
rect 1515 1844 1516 1848
rect 1510 1843 1516 1844
rect 1670 1848 1676 1849
rect 1670 1844 1671 1848
rect 1675 1844 1676 1848
rect 1670 1843 1676 1844
rect 1814 1848 1820 1849
rect 1814 1844 1815 1848
rect 1819 1844 1820 1848
rect 1814 1843 1820 1844
rect 1934 1847 1940 1848
rect 1934 1843 1935 1847
rect 1939 1843 1940 1847
rect 110 1842 116 1843
rect 112 1807 114 1842
rect 264 1807 266 1843
rect 464 1807 466 1843
rect 656 1807 658 1843
rect 840 1807 842 1843
rect 1016 1807 1018 1843
rect 1184 1807 1186 1843
rect 1352 1807 1354 1843
rect 1512 1807 1514 1843
rect 1672 1807 1674 1843
rect 1816 1807 1818 1843
rect 1934 1842 1940 1843
rect 1936 1807 1938 1842
rect 1976 1807 1978 1879
rect 3108 1807 3110 1880
rect 3244 1807 3246 1880
rect 3380 1807 3382 1880
rect 3516 1807 3518 1880
rect 3652 1807 3654 1880
rect 3798 1879 3804 1880
rect 3800 1807 3802 1879
rect 3886 1872 3892 1873
rect 3838 1871 3844 1872
rect 3838 1867 3839 1871
rect 3843 1867 3844 1871
rect 3886 1868 3887 1872
rect 3891 1868 3892 1872
rect 3886 1867 3892 1868
rect 4070 1872 4076 1873
rect 4070 1868 4071 1872
rect 4075 1868 4076 1872
rect 4070 1867 4076 1868
rect 4310 1872 4316 1873
rect 4310 1868 4311 1872
rect 4315 1868 4316 1872
rect 4310 1867 4316 1868
rect 4590 1872 4596 1873
rect 4590 1868 4591 1872
rect 4595 1868 4596 1872
rect 4590 1867 4596 1868
rect 4902 1872 4908 1873
rect 4902 1868 4903 1872
rect 4907 1868 4908 1872
rect 4902 1867 4908 1868
rect 5230 1872 5236 1873
rect 5230 1868 5231 1872
rect 5235 1868 5236 1872
rect 5230 1867 5236 1868
rect 5542 1872 5548 1873
rect 5542 1868 5543 1872
rect 5547 1868 5548 1872
rect 5542 1867 5548 1868
rect 5662 1871 5668 1872
rect 5662 1867 5663 1871
rect 5667 1867 5668 1871
rect 3838 1866 3844 1867
rect 3840 1843 3842 1866
rect 3888 1843 3890 1867
rect 4072 1843 4074 1867
rect 4312 1843 4314 1867
rect 4592 1843 4594 1867
rect 4904 1843 4906 1867
rect 5232 1843 5234 1867
rect 5544 1843 5546 1867
rect 5662 1866 5668 1867
rect 5664 1843 5666 1866
rect 3839 1842 3843 1843
rect 3839 1837 3843 1838
rect 3887 1842 3891 1843
rect 3887 1837 3891 1838
rect 4071 1842 4075 1843
rect 4071 1837 4075 1838
rect 4311 1842 4315 1843
rect 4311 1837 4315 1838
rect 4407 1842 4411 1843
rect 4407 1837 4411 1838
rect 4543 1842 4547 1843
rect 4543 1837 4547 1838
rect 4591 1842 4595 1843
rect 4591 1837 4595 1838
rect 4679 1842 4683 1843
rect 4679 1837 4683 1838
rect 4815 1842 4819 1843
rect 4815 1837 4819 1838
rect 4903 1842 4907 1843
rect 4903 1837 4907 1838
rect 4951 1842 4955 1843
rect 4951 1837 4955 1838
rect 5231 1842 5235 1843
rect 5231 1837 5235 1838
rect 5543 1842 5547 1843
rect 5543 1837 5547 1838
rect 5663 1842 5667 1843
rect 5663 1837 5667 1838
rect 3840 1814 3842 1837
rect 3838 1813 3844 1814
rect 4408 1813 4410 1837
rect 4544 1813 4546 1837
rect 4680 1813 4682 1837
rect 4816 1813 4818 1837
rect 4952 1813 4954 1837
rect 5664 1814 5666 1837
rect 5662 1813 5668 1814
rect 3838 1809 3839 1813
rect 3843 1809 3844 1813
rect 3838 1808 3844 1809
rect 4406 1812 4412 1813
rect 4406 1808 4407 1812
rect 4411 1808 4412 1812
rect 4406 1807 4412 1808
rect 4542 1812 4548 1813
rect 4542 1808 4543 1812
rect 4547 1808 4548 1812
rect 4542 1807 4548 1808
rect 4678 1812 4684 1813
rect 4678 1808 4679 1812
rect 4683 1808 4684 1812
rect 4678 1807 4684 1808
rect 4814 1812 4820 1813
rect 4814 1808 4815 1812
rect 4819 1808 4820 1812
rect 4814 1807 4820 1808
rect 4950 1812 4956 1813
rect 4950 1808 4951 1812
rect 4955 1808 4956 1812
rect 5662 1809 5663 1813
rect 5667 1809 5668 1813
rect 5662 1808 5668 1809
rect 4950 1807 4956 1808
rect 111 1806 115 1807
rect 111 1801 115 1802
rect 223 1806 227 1807
rect 223 1801 227 1802
rect 263 1806 267 1807
rect 263 1801 267 1802
rect 463 1806 467 1807
rect 463 1801 467 1802
rect 655 1806 659 1807
rect 655 1801 659 1802
rect 695 1806 699 1807
rect 695 1801 699 1802
rect 839 1806 843 1807
rect 839 1801 843 1802
rect 927 1806 931 1807
rect 927 1801 931 1802
rect 1015 1806 1019 1807
rect 1015 1801 1019 1802
rect 1159 1806 1163 1807
rect 1159 1801 1163 1802
rect 1183 1806 1187 1807
rect 1183 1801 1187 1802
rect 1351 1806 1355 1807
rect 1351 1801 1355 1802
rect 1391 1806 1395 1807
rect 1391 1801 1395 1802
rect 1511 1806 1515 1807
rect 1511 1801 1515 1802
rect 1671 1806 1675 1807
rect 1671 1801 1675 1802
rect 1815 1806 1819 1807
rect 1815 1801 1819 1802
rect 1935 1806 1939 1807
rect 1935 1801 1939 1802
rect 1975 1806 1979 1807
rect 1975 1801 1979 1802
rect 1995 1806 1999 1807
rect 1995 1801 1999 1802
rect 2131 1806 2135 1807
rect 2131 1801 2135 1802
rect 2267 1806 2271 1807
rect 2267 1801 2271 1802
rect 2419 1806 2423 1807
rect 2419 1801 2423 1802
rect 2579 1806 2583 1807
rect 2579 1801 2583 1802
rect 2739 1806 2743 1807
rect 2739 1801 2743 1802
rect 2899 1806 2903 1807
rect 2899 1801 2903 1802
rect 3051 1806 3055 1807
rect 3051 1801 3055 1802
rect 3107 1806 3111 1807
rect 3107 1801 3111 1802
rect 3203 1806 3207 1807
rect 3203 1801 3207 1802
rect 3243 1806 3247 1807
rect 3243 1801 3247 1802
rect 3355 1806 3359 1807
rect 3355 1801 3359 1802
rect 3379 1806 3383 1807
rect 3379 1801 3383 1802
rect 3515 1806 3519 1807
rect 3515 1801 3519 1802
rect 3651 1806 3655 1807
rect 3651 1801 3655 1802
rect 3799 1806 3803 1807
rect 3799 1801 3803 1802
rect 112 1778 114 1801
rect 110 1777 116 1778
rect 224 1777 226 1801
rect 464 1777 466 1801
rect 696 1777 698 1801
rect 928 1777 930 1801
rect 1160 1777 1162 1801
rect 1392 1777 1394 1801
rect 1936 1778 1938 1801
rect 1934 1777 1940 1778
rect 110 1773 111 1777
rect 115 1773 116 1777
rect 110 1772 116 1773
rect 222 1776 228 1777
rect 222 1772 223 1776
rect 227 1772 228 1776
rect 222 1771 228 1772
rect 462 1776 468 1777
rect 462 1772 463 1776
rect 467 1772 468 1776
rect 462 1771 468 1772
rect 694 1776 700 1777
rect 694 1772 695 1776
rect 699 1772 700 1776
rect 694 1771 700 1772
rect 926 1776 932 1777
rect 926 1772 927 1776
rect 931 1772 932 1776
rect 926 1771 932 1772
rect 1158 1776 1164 1777
rect 1158 1772 1159 1776
rect 1163 1772 1164 1776
rect 1158 1771 1164 1772
rect 1390 1776 1396 1777
rect 1390 1772 1391 1776
rect 1395 1772 1396 1776
rect 1934 1773 1935 1777
rect 1939 1773 1940 1777
rect 1934 1772 1940 1773
rect 1390 1771 1396 1772
rect 194 1761 200 1762
rect 110 1760 116 1761
rect 110 1756 111 1760
rect 115 1756 116 1760
rect 194 1757 195 1761
rect 199 1757 200 1761
rect 194 1756 200 1757
rect 434 1761 440 1762
rect 434 1757 435 1761
rect 439 1757 440 1761
rect 434 1756 440 1757
rect 666 1761 672 1762
rect 666 1757 667 1761
rect 671 1757 672 1761
rect 666 1756 672 1757
rect 898 1761 904 1762
rect 898 1757 899 1761
rect 903 1757 904 1761
rect 898 1756 904 1757
rect 1130 1761 1136 1762
rect 1130 1757 1131 1761
rect 1135 1757 1136 1761
rect 1130 1756 1136 1757
rect 1362 1761 1368 1762
rect 1362 1757 1363 1761
rect 1367 1757 1368 1761
rect 1362 1756 1368 1757
rect 1934 1760 1940 1761
rect 1934 1756 1935 1760
rect 1939 1756 1940 1760
rect 110 1755 116 1756
rect 112 1683 114 1755
rect 196 1683 198 1756
rect 436 1683 438 1756
rect 668 1683 670 1756
rect 900 1683 902 1756
rect 1132 1683 1134 1756
rect 1364 1683 1366 1756
rect 1934 1755 1940 1756
rect 1936 1683 1938 1755
rect 1976 1741 1978 1801
rect 1974 1740 1980 1741
rect 1996 1740 1998 1801
rect 2132 1740 2134 1801
rect 2268 1740 2270 1801
rect 2420 1740 2422 1801
rect 2580 1740 2582 1801
rect 2740 1740 2742 1801
rect 2900 1740 2902 1801
rect 3052 1740 3054 1801
rect 3204 1740 3206 1801
rect 3356 1740 3358 1801
rect 3516 1740 3518 1801
rect 3652 1740 3654 1801
rect 3800 1741 3802 1801
rect 4378 1797 4384 1798
rect 3838 1796 3844 1797
rect 3838 1792 3839 1796
rect 3843 1792 3844 1796
rect 4378 1793 4379 1797
rect 4383 1793 4384 1797
rect 4378 1792 4384 1793
rect 4514 1797 4520 1798
rect 4514 1793 4515 1797
rect 4519 1793 4520 1797
rect 4514 1792 4520 1793
rect 4650 1797 4656 1798
rect 4650 1793 4651 1797
rect 4655 1793 4656 1797
rect 4650 1792 4656 1793
rect 4786 1797 4792 1798
rect 4786 1793 4787 1797
rect 4791 1793 4792 1797
rect 4786 1792 4792 1793
rect 4922 1797 4928 1798
rect 4922 1793 4923 1797
rect 4927 1793 4928 1797
rect 4922 1792 4928 1793
rect 5662 1796 5668 1797
rect 5662 1792 5663 1796
rect 5667 1792 5668 1796
rect 3838 1791 3844 1792
rect 3798 1740 3804 1741
rect 1974 1736 1975 1740
rect 1979 1736 1980 1740
rect 1974 1735 1980 1736
rect 1994 1739 2000 1740
rect 1994 1735 1995 1739
rect 1999 1735 2000 1739
rect 1994 1734 2000 1735
rect 2130 1739 2136 1740
rect 2130 1735 2131 1739
rect 2135 1735 2136 1739
rect 2130 1734 2136 1735
rect 2266 1739 2272 1740
rect 2266 1735 2267 1739
rect 2271 1735 2272 1739
rect 2266 1734 2272 1735
rect 2418 1739 2424 1740
rect 2418 1735 2419 1739
rect 2423 1735 2424 1739
rect 2418 1734 2424 1735
rect 2578 1739 2584 1740
rect 2578 1735 2579 1739
rect 2583 1735 2584 1739
rect 2578 1734 2584 1735
rect 2738 1739 2744 1740
rect 2738 1735 2739 1739
rect 2743 1735 2744 1739
rect 2738 1734 2744 1735
rect 2898 1739 2904 1740
rect 2898 1735 2899 1739
rect 2903 1735 2904 1739
rect 2898 1734 2904 1735
rect 3050 1739 3056 1740
rect 3050 1735 3051 1739
rect 3055 1735 3056 1739
rect 3050 1734 3056 1735
rect 3202 1739 3208 1740
rect 3202 1735 3203 1739
rect 3207 1735 3208 1739
rect 3202 1734 3208 1735
rect 3354 1739 3360 1740
rect 3354 1735 3355 1739
rect 3359 1735 3360 1739
rect 3354 1734 3360 1735
rect 3514 1739 3520 1740
rect 3514 1735 3515 1739
rect 3519 1735 3520 1739
rect 3514 1734 3520 1735
rect 3650 1739 3656 1740
rect 3650 1735 3651 1739
rect 3655 1735 3656 1739
rect 3798 1736 3799 1740
rect 3803 1736 3804 1740
rect 3798 1735 3804 1736
rect 3650 1734 3656 1735
rect 2022 1724 2028 1725
rect 1974 1723 1980 1724
rect 1974 1719 1975 1723
rect 1979 1719 1980 1723
rect 2022 1720 2023 1724
rect 2027 1720 2028 1724
rect 2022 1719 2028 1720
rect 2158 1724 2164 1725
rect 2158 1720 2159 1724
rect 2163 1720 2164 1724
rect 2158 1719 2164 1720
rect 2294 1724 2300 1725
rect 2294 1720 2295 1724
rect 2299 1720 2300 1724
rect 2294 1719 2300 1720
rect 2446 1724 2452 1725
rect 2446 1720 2447 1724
rect 2451 1720 2452 1724
rect 2446 1719 2452 1720
rect 2606 1724 2612 1725
rect 2606 1720 2607 1724
rect 2611 1720 2612 1724
rect 2606 1719 2612 1720
rect 2766 1724 2772 1725
rect 2766 1720 2767 1724
rect 2771 1720 2772 1724
rect 2766 1719 2772 1720
rect 2926 1724 2932 1725
rect 2926 1720 2927 1724
rect 2931 1720 2932 1724
rect 2926 1719 2932 1720
rect 3078 1724 3084 1725
rect 3078 1720 3079 1724
rect 3083 1720 3084 1724
rect 3078 1719 3084 1720
rect 3230 1724 3236 1725
rect 3230 1720 3231 1724
rect 3235 1720 3236 1724
rect 3230 1719 3236 1720
rect 3382 1724 3388 1725
rect 3382 1720 3383 1724
rect 3387 1720 3388 1724
rect 3382 1719 3388 1720
rect 3542 1724 3548 1725
rect 3542 1720 3543 1724
rect 3547 1720 3548 1724
rect 3542 1719 3548 1720
rect 3678 1724 3684 1725
rect 3678 1720 3679 1724
rect 3683 1720 3684 1724
rect 3678 1719 3684 1720
rect 3798 1723 3804 1724
rect 3798 1719 3799 1723
rect 3803 1719 3804 1723
rect 1974 1718 1980 1719
rect 1976 1683 1978 1718
rect 2024 1683 2026 1719
rect 2160 1683 2162 1719
rect 2296 1683 2298 1719
rect 2448 1683 2450 1719
rect 2608 1683 2610 1719
rect 2768 1683 2770 1719
rect 2928 1683 2930 1719
rect 3080 1683 3082 1719
rect 3232 1683 3234 1719
rect 3384 1683 3386 1719
rect 3544 1683 3546 1719
rect 3680 1683 3682 1719
rect 3798 1718 3804 1719
rect 3800 1683 3802 1718
rect 3840 1715 3842 1791
rect 4380 1715 4382 1792
rect 4516 1715 4518 1792
rect 4652 1715 4654 1792
rect 4788 1715 4790 1792
rect 4924 1715 4926 1792
rect 5662 1791 5668 1792
rect 5664 1715 5666 1791
rect 3839 1714 3843 1715
rect 3839 1709 3843 1710
rect 4379 1714 4383 1715
rect 4379 1709 4383 1710
rect 4515 1714 4519 1715
rect 4515 1709 4519 1710
rect 4563 1714 4567 1715
rect 4563 1709 4567 1710
rect 4651 1714 4655 1715
rect 4651 1709 4655 1710
rect 4699 1714 4703 1715
rect 4699 1709 4703 1710
rect 4787 1714 4791 1715
rect 4787 1709 4791 1710
rect 4835 1714 4839 1715
rect 4835 1709 4839 1710
rect 4923 1714 4927 1715
rect 4923 1709 4927 1710
rect 4971 1714 4975 1715
rect 4971 1709 4975 1710
rect 5107 1714 5111 1715
rect 5107 1709 5111 1710
rect 5243 1714 5247 1715
rect 5243 1709 5247 1710
rect 5379 1714 5383 1715
rect 5379 1709 5383 1710
rect 5515 1714 5519 1715
rect 5515 1709 5519 1710
rect 5663 1714 5667 1715
rect 5663 1709 5667 1710
rect 111 1682 115 1683
rect 111 1677 115 1678
rect 131 1682 135 1683
rect 131 1677 135 1678
rect 195 1682 199 1683
rect 195 1677 199 1678
rect 363 1682 367 1683
rect 363 1677 367 1678
rect 435 1682 439 1683
rect 435 1677 439 1678
rect 619 1682 623 1683
rect 619 1677 623 1678
rect 667 1682 671 1683
rect 667 1677 671 1678
rect 875 1682 879 1683
rect 875 1677 879 1678
rect 899 1682 903 1683
rect 899 1677 903 1678
rect 1131 1682 1135 1683
rect 1131 1677 1135 1678
rect 1139 1682 1143 1683
rect 1139 1677 1143 1678
rect 1363 1682 1367 1683
rect 1363 1677 1367 1678
rect 1935 1682 1939 1683
rect 1935 1677 1939 1678
rect 1975 1682 1979 1683
rect 1975 1677 1979 1678
rect 2023 1682 2027 1683
rect 2023 1677 2027 1678
rect 2159 1682 2163 1683
rect 2159 1677 2163 1678
rect 2167 1682 2171 1683
rect 2167 1677 2171 1678
rect 2295 1682 2299 1683
rect 2295 1677 2299 1678
rect 2319 1682 2323 1683
rect 2319 1677 2323 1678
rect 2447 1682 2451 1683
rect 2447 1677 2451 1678
rect 2479 1682 2483 1683
rect 2479 1677 2483 1678
rect 2607 1682 2611 1683
rect 2607 1677 2611 1678
rect 2639 1682 2643 1683
rect 2639 1677 2643 1678
rect 2767 1682 2771 1683
rect 2767 1677 2771 1678
rect 2791 1682 2795 1683
rect 2791 1677 2795 1678
rect 2927 1682 2931 1683
rect 2927 1677 2931 1678
rect 2943 1682 2947 1683
rect 2943 1677 2947 1678
rect 3079 1682 3083 1683
rect 3079 1677 3083 1678
rect 3103 1682 3107 1683
rect 3103 1677 3107 1678
rect 3231 1682 3235 1683
rect 3231 1677 3235 1678
rect 3263 1682 3267 1683
rect 3263 1677 3267 1678
rect 3383 1682 3387 1683
rect 3383 1677 3387 1678
rect 3423 1682 3427 1683
rect 3423 1677 3427 1678
rect 3543 1682 3547 1683
rect 3543 1677 3547 1678
rect 3679 1682 3683 1683
rect 3679 1677 3683 1678
rect 3799 1682 3803 1683
rect 3799 1677 3803 1678
rect 112 1617 114 1677
rect 110 1616 116 1617
rect 132 1616 134 1677
rect 364 1616 366 1677
rect 620 1616 622 1677
rect 876 1616 878 1677
rect 1140 1616 1142 1677
rect 1936 1617 1938 1677
rect 1976 1654 1978 1677
rect 1974 1653 1980 1654
rect 2024 1653 2026 1677
rect 2168 1653 2170 1677
rect 2320 1653 2322 1677
rect 2480 1653 2482 1677
rect 2640 1653 2642 1677
rect 2792 1653 2794 1677
rect 2944 1653 2946 1677
rect 3104 1653 3106 1677
rect 3264 1653 3266 1677
rect 3424 1653 3426 1677
rect 3800 1654 3802 1677
rect 3798 1653 3804 1654
rect 1974 1649 1975 1653
rect 1979 1649 1980 1653
rect 1974 1648 1980 1649
rect 2022 1652 2028 1653
rect 2022 1648 2023 1652
rect 2027 1648 2028 1652
rect 2022 1647 2028 1648
rect 2166 1652 2172 1653
rect 2166 1648 2167 1652
rect 2171 1648 2172 1652
rect 2166 1647 2172 1648
rect 2318 1652 2324 1653
rect 2318 1648 2319 1652
rect 2323 1648 2324 1652
rect 2318 1647 2324 1648
rect 2478 1652 2484 1653
rect 2478 1648 2479 1652
rect 2483 1648 2484 1652
rect 2478 1647 2484 1648
rect 2638 1652 2644 1653
rect 2638 1648 2639 1652
rect 2643 1648 2644 1652
rect 2638 1647 2644 1648
rect 2790 1652 2796 1653
rect 2790 1648 2791 1652
rect 2795 1648 2796 1652
rect 2790 1647 2796 1648
rect 2942 1652 2948 1653
rect 2942 1648 2943 1652
rect 2947 1648 2948 1652
rect 2942 1647 2948 1648
rect 3102 1652 3108 1653
rect 3102 1648 3103 1652
rect 3107 1648 3108 1652
rect 3102 1647 3108 1648
rect 3262 1652 3268 1653
rect 3262 1648 3263 1652
rect 3267 1648 3268 1652
rect 3262 1647 3268 1648
rect 3422 1652 3428 1653
rect 3422 1648 3423 1652
rect 3427 1648 3428 1652
rect 3798 1649 3799 1653
rect 3803 1649 3804 1653
rect 3840 1649 3842 1709
rect 3798 1648 3804 1649
rect 3838 1648 3844 1649
rect 4564 1648 4566 1709
rect 4700 1648 4702 1709
rect 4836 1648 4838 1709
rect 4972 1648 4974 1709
rect 5108 1648 5110 1709
rect 5244 1648 5246 1709
rect 5380 1648 5382 1709
rect 5516 1648 5518 1709
rect 5664 1649 5666 1709
rect 5662 1648 5668 1649
rect 3422 1647 3428 1648
rect 3838 1644 3839 1648
rect 3843 1644 3844 1648
rect 3838 1643 3844 1644
rect 4562 1647 4568 1648
rect 4562 1643 4563 1647
rect 4567 1643 4568 1647
rect 4562 1642 4568 1643
rect 4698 1647 4704 1648
rect 4698 1643 4699 1647
rect 4703 1643 4704 1647
rect 4698 1642 4704 1643
rect 4834 1647 4840 1648
rect 4834 1643 4835 1647
rect 4839 1643 4840 1647
rect 4834 1642 4840 1643
rect 4970 1647 4976 1648
rect 4970 1643 4971 1647
rect 4975 1643 4976 1647
rect 4970 1642 4976 1643
rect 5106 1647 5112 1648
rect 5106 1643 5107 1647
rect 5111 1643 5112 1647
rect 5106 1642 5112 1643
rect 5242 1647 5248 1648
rect 5242 1643 5243 1647
rect 5247 1643 5248 1647
rect 5242 1642 5248 1643
rect 5378 1647 5384 1648
rect 5378 1643 5379 1647
rect 5383 1643 5384 1647
rect 5378 1642 5384 1643
rect 5514 1647 5520 1648
rect 5514 1643 5515 1647
rect 5519 1643 5520 1647
rect 5662 1644 5663 1648
rect 5667 1644 5668 1648
rect 5662 1643 5668 1644
rect 5514 1642 5520 1643
rect 1994 1637 2000 1638
rect 1974 1636 1980 1637
rect 1974 1632 1975 1636
rect 1979 1632 1980 1636
rect 1994 1633 1995 1637
rect 1999 1633 2000 1637
rect 1994 1632 2000 1633
rect 2138 1637 2144 1638
rect 2138 1633 2139 1637
rect 2143 1633 2144 1637
rect 2138 1632 2144 1633
rect 2290 1637 2296 1638
rect 2290 1633 2291 1637
rect 2295 1633 2296 1637
rect 2290 1632 2296 1633
rect 2450 1637 2456 1638
rect 2450 1633 2451 1637
rect 2455 1633 2456 1637
rect 2450 1632 2456 1633
rect 2610 1637 2616 1638
rect 2610 1633 2611 1637
rect 2615 1633 2616 1637
rect 2610 1632 2616 1633
rect 2762 1637 2768 1638
rect 2762 1633 2763 1637
rect 2767 1633 2768 1637
rect 2762 1632 2768 1633
rect 2914 1637 2920 1638
rect 2914 1633 2915 1637
rect 2919 1633 2920 1637
rect 2914 1632 2920 1633
rect 3074 1637 3080 1638
rect 3074 1633 3075 1637
rect 3079 1633 3080 1637
rect 3074 1632 3080 1633
rect 3234 1637 3240 1638
rect 3234 1633 3235 1637
rect 3239 1633 3240 1637
rect 3234 1632 3240 1633
rect 3394 1637 3400 1638
rect 3394 1633 3395 1637
rect 3399 1633 3400 1637
rect 3394 1632 3400 1633
rect 3798 1636 3804 1637
rect 3798 1632 3799 1636
rect 3803 1632 3804 1636
rect 4590 1632 4596 1633
rect 1974 1631 1980 1632
rect 1934 1616 1940 1617
rect 110 1612 111 1616
rect 115 1612 116 1616
rect 110 1611 116 1612
rect 130 1615 136 1616
rect 130 1611 131 1615
rect 135 1611 136 1615
rect 130 1610 136 1611
rect 362 1615 368 1616
rect 362 1611 363 1615
rect 367 1611 368 1615
rect 362 1610 368 1611
rect 618 1615 624 1616
rect 618 1611 619 1615
rect 623 1611 624 1615
rect 618 1610 624 1611
rect 874 1615 880 1616
rect 874 1611 875 1615
rect 879 1611 880 1615
rect 874 1610 880 1611
rect 1138 1615 1144 1616
rect 1138 1611 1139 1615
rect 1143 1611 1144 1615
rect 1934 1612 1935 1616
rect 1939 1612 1940 1616
rect 1934 1611 1940 1612
rect 1138 1610 1144 1611
rect 158 1600 164 1601
rect 110 1599 116 1600
rect 110 1595 111 1599
rect 115 1595 116 1599
rect 158 1596 159 1600
rect 163 1596 164 1600
rect 158 1595 164 1596
rect 390 1600 396 1601
rect 390 1596 391 1600
rect 395 1596 396 1600
rect 390 1595 396 1596
rect 646 1600 652 1601
rect 646 1596 647 1600
rect 651 1596 652 1600
rect 646 1595 652 1596
rect 902 1600 908 1601
rect 902 1596 903 1600
rect 907 1596 908 1600
rect 902 1595 908 1596
rect 1166 1600 1172 1601
rect 1166 1596 1167 1600
rect 1171 1596 1172 1600
rect 1166 1595 1172 1596
rect 1934 1599 1940 1600
rect 1934 1595 1935 1599
rect 1939 1595 1940 1599
rect 110 1594 116 1595
rect 112 1559 114 1594
rect 160 1559 162 1595
rect 392 1559 394 1595
rect 648 1559 650 1595
rect 904 1559 906 1595
rect 1168 1559 1170 1595
rect 1934 1594 1940 1595
rect 1936 1559 1938 1594
rect 1976 1559 1978 1631
rect 1996 1559 1998 1632
rect 2140 1559 2142 1632
rect 2292 1559 2294 1632
rect 2452 1559 2454 1632
rect 2612 1559 2614 1632
rect 2764 1559 2766 1632
rect 2916 1559 2918 1632
rect 3076 1559 3078 1632
rect 3236 1559 3238 1632
rect 3396 1559 3398 1632
rect 3798 1631 3804 1632
rect 3838 1631 3844 1632
rect 3800 1559 3802 1631
rect 3838 1627 3839 1631
rect 3843 1627 3844 1631
rect 4590 1628 4591 1632
rect 4595 1628 4596 1632
rect 4590 1627 4596 1628
rect 4726 1632 4732 1633
rect 4726 1628 4727 1632
rect 4731 1628 4732 1632
rect 4726 1627 4732 1628
rect 4862 1632 4868 1633
rect 4862 1628 4863 1632
rect 4867 1628 4868 1632
rect 4862 1627 4868 1628
rect 4998 1632 5004 1633
rect 4998 1628 4999 1632
rect 5003 1628 5004 1632
rect 4998 1627 5004 1628
rect 5134 1632 5140 1633
rect 5134 1628 5135 1632
rect 5139 1628 5140 1632
rect 5134 1627 5140 1628
rect 5270 1632 5276 1633
rect 5270 1628 5271 1632
rect 5275 1628 5276 1632
rect 5270 1627 5276 1628
rect 5406 1632 5412 1633
rect 5406 1628 5407 1632
rect 5411 1628 5412 1632
rect 5406 1627 5412 1628
rect 5542 1632 5548 1633
rect 5542 1628 5543 1632
rect 5547 1628 5548 1632
rect 5542 1627 5548 1628
rect 5662 1631 5668 1632
rect 5662 1627 5663 1631
rect 5667 1627 5668 1631
rect 3838 1626 3844 1627
rect 3840 1587 3842 1626
rect 4592 1587 4594 1627
rect 4728 1587 4730 1627
rect 4864 1587 4866 1627
rect 5000 1587 5002 1627
rect 5136 1587 5138 1627
rect 5272 1587 5274 1627
rect 5408 1587 5410 1627
rect 5544 1587 5546 1627
rect 5662 1626 5668 1627
rect 5664 1587 5666 1626
rect 3839 1586 3843 1587
rect 3839 1581 3843 1582
rect 4591 1586 4595 1587
rect 4591 1581 4595 1582
rect 4727 1586 4731 1587
rect 4727 1581 4731 1582
rect 4863 1586 4867 1587
rect 4863 1581 4867 1582
rect 4999 1586 5003 1587
rect 4999 1581 5003 1582
rect 5135 1586 5139 1587
rect 5135 1581 5139 1582
rect 5271 1586 5275 1587
rect 5271 1581 5275 1582
rect 5407 1586 5411 1587
rect 5407 1581 5411 1582
rect 5543 1586 5547 1587
rect 5543 1581 5547 1582
rect 5663 1586 5667 1587
rect 5663 1581 5667 1582
rect 111 1558 115 1559
rect 111 1553 115 1554
rect 159 1558 163 1559
rect 159 1553 163 1554
rect 327 1558 331 1559
rect 327 1553 331 1554
rect 391 1558 395 1559
rect 391 1553 395 1554
rect 511 1558 515 1559
rect 511 1553 515 1554
rect 647 1558 651 1559
rect 647 1553 651 1554
rect 695 1558 699 1559
rect 695 1553 699 1554
rect 887 1558 891 1559
rect 887 1553 891 1554
rect 903 1558 907 1559
rect 903 1553 907 1554
rect 1079 1558 1083 1559
rect 1079 1553 1083 1554
rect 1167 1558 1171 1559
rect 1167 1553 1171 1554
rect 1935 1558 1939 1559
rect 1935 1553 1939 1554
rect 1975 1558 1979 1559
rect 1975 1553 1979 1554
rect 1995 1558 1999 1559
rect 1995 1553 1999 1554
rect 2131 1558 2135 1559
rect 2131 1553 2135 1554
rect 2139 1558 2143 1559
rect 2139 1553 2143 1554
rect 2267 1558 2271 1559
rect 2267 1553 2271 1554
rect 2291 1558 2295 1559
rect 2291 1553 2295 1554
rect 2403 1558 2407 1559
rect 2403 1553 2407 1554
rect 2451 1558 2455 1559
rect 2451 1553 2455 1554
rect 2539 1558 2543 1559
rect 2539 1553 2543 1554
rect 2611 1558 2615 1559
rect 2611 1553 2615 1554
rect 2675 1558 2679 1559
rect 2675 1553 2679 1554
rect 2763 1558 2767 1559
rect 2763 1553 2767 1554
rect 2811 1558 2815 1559
rect 2811 1553 2815 1554
rect 2915 1558 2919 1559
rect 2915 1553 2919 1554
rect 2947 1558 2951 1559
rect 2947 1553 2951 1554
rect 3075 1558 3079 1559
rect 3075 1553 3079 1554
rect 3083 1558 3087 1559
rect 3083 1553 3087 1554
rect 3219 1558 3223 1559
rect 3219 1553 3223 1554
rect 3235 1558 3239 1559
rect 3235 1553 3239 1554
rect 3355 1558 3359 1559
rect 3355 1553 3359 1554
rect 3395 1558 3399 1559
rect 3395 1553 3399 1554
rect 3491 1558 3495 1559
rect 3491 1553 3495 1554
rect 3799 1558 3803 1559
rect 3840 1558 3842 1581
rect 3799 1553 3803 1554
rect 3838 1557 3844 1558
rect 4592 1557 4594 1581
rect 4728 1557 4730 1581
rect 4864 1557 4866 1581
rect 5000 1557 5002 1581
rect 5136 1557 5138 1581
rect 5272 1557 5274 1581
rect 5408 1557 5410 1581
rect 5544 1557 5546 1581
rect 5664 1558 5666 1581
rect 5662 1557 5668 1558
rect 3838 1553 3839 1557
rect 3843 1553 3844 1557
rect 112 1530 114 1553
rect 110 1529 116 1530
rect 160 1529 162 1553
rect 328 1529 330 1553
rect 512 1529 514 1553
rect 696 1529 698 1553
rect 888 1529 890 1553
rect 1080 1529 1082 1553
rect 1936 1530 1938 1553
rect 1934 1529 1940 1530
rect 110 1525 111 1529
rect 115 1525 116 1529
rect 110 1524 116 1525
rect 158 1528 164 1529
rect 158 1524 159 1528
rect 163 1524 164 1528
rect 158 1523 164 1524
rect 326 1528 332 1529
rect 326 1524 327 1528
rect 331 1524 332 1528
rect 326 1523 332 1524
rect 510 1528 516 1529
rect 510 1524 511 1528
rect 515 1524 516 1528
rect 510 1523 516 1524
rect 694 1528 700 1529
rect 694 1524 695 1528
rect 699 1524 700 1528
rect 694 1523 700 1524
rect 886 1528 892 1529
rect 886 1524 887 1528
rect 891 1524 892 1528
rect 886 1523 892 1524
rect 1078 1528 1084 1529
rect 1078 1524 1079 1528
rect 1083 1524 1084 1528
rect 1934 1525 1935 1529
rect 1939 1525 1940 1529
rect 1934 1524 1940 1525
rect 1078 1523 1084 1524
rect 130 1513 136 1514
rect 110 1512 116 1513
rect 110 1508 111 1512
rect 115 1508 116 1512
rect 130 1509 131 1513
rect 135 1509 136 1513
rect 130 1508 136 1509
rect 298 1513 304 1514
rect 298 1509 299 1513
rect 303 1509 304 1513
rect 298 1508 304 1509
rect 482 1513 488 1514
rect 482 1509 483 1513
rect 487 1509 488 1513
rect 482 1508 488 1509
rect 666 1513 672 1514
rect 666 1509 667 1513
rect 671 1509 672 1513
rect 666 1508 672 1509
rect 858 1513 864 1514
rect 858 1509 859 1513
rect 863 1509 864 1513
rect 858 1508 864 1509
rect 1050 1513 1056 1514
rect 1050 1509 1051 1513
rect 1055 1509 1056 1513
rect 1050 1508 1056 1509
rect 1934 1512 1940 1513
rect 1934 1508 1935 1512
rect 1939 1508 1940 1512
rect 110 1507 116 1508
rect 112 1435 114 1507
rect 132 1435 134 1508
rect 300 1435 302 1508
rect 484 1435 486 1508
rect 668 1435 670 1508
rect 860 1435 862 1508
rect 1052 1435 1054 1508
rect 1934 1507 1940 1508
rect 1936 1435 1938 1507
rect 1976 1493 1978 1553
rect 1974 1492 1980 1493
rect 1996 1492 1998 1553
rect 2132 1492 2134 1553
rect 2268 1492 2270 1553
rect 2404 1492 2406 1553
rect 2540 1492 2542 1553
rect 2676 1492 2678 1553
rect 2812 1492 2814 1553
rect 2948 1492 2950 1553
rect 3084 1492 3086 1553
rect 3220 1492 3222 1553
rect 3356 1492 3358 1553
rect 3492 1492 3494 1553
rect 3800 1493 3802 1553
rect 3838 1552 3844 1553
rect 4590 1556 4596 1557
rect 4590 1552 4591 1556
rect 4595 1552 4596 1556
rect 4590 1551 4596 1552
rect 4726 1556 4732 1557
rect 4726 1552 4727 1556
rect 4731 1552 4732 1556
rect 4726 1551 4732 1552
rect 4862 1556 4868 1557
rect 4862 1552 4863 1556
rect 4867 1552 4868 1556
rect 4862 1551 4868 1552
rect 4998 1556 5004 1557
rect 4998 1552 4999 1556
rect 5003 1552 5004 1556
rect 4998 1551 5004 1552
rect 5134 1556 5140 1557
rect 5134 1552 5135 1556
rect 5139 1552 5140 1556
rect 5134 1551 5140 1552
rect 5270 1556 5276 1557
rect 5270 1552 5271 1556
rect 5275 1552 5276 1556
rect 5270 1551 5276 1552
rect 5406 1556 5412 1557
rect 5406 1552 5407 1556
rect 5411 1552 5412 1556
rect 5406 1551 5412 1552
rect 5542 1556 5548 1557
rect 5542 1552 5543 1556
rect 5547 1552 5548 1556
rect 5662 1553 5663 1557
rect 5667 1553 5668 1557
rect 5662 1552 5668 1553
rect 5542 1551 5548 1552
rect 4562 1541 4568 1542
rect 3838 1540 3844 1541
rect 3838 1536 3839 1540
rect 3843 1536 3844 1540
rect 4562 1537 4563 1541
rect 4567 1537 4568 1541
rect 4562 1536 4568 1537
rect 4698 1541 4704 1542
rect 4698 1537 4699 1541
rect 4703 1537 4704 1541
rect 4698 1536 4704 1537
rect 4834 1541 4840 1542
rect 4834 1537 4835 1541
rect 4839 1537 4840 1541
rect 4834 1536 4840 1537
rect 4970 1541 4976 1542
rect 4970 1537 4971 1541
rect 4975 1537 4976 1541
rect 4970 1536 4976 1537
rect 5106 1541 5112 1542
rect 5106 1537 5107 1541
rect 5111 1537 5112 1541
rect 5106 1536 5112 1537
rect 5242 1541 5248 1542
rect 5242 1537 5243 1541
rect 5247 1537 5248 1541
rect 5242 1536 5248 1537
rect 5378 1541 5384 1542
rect 5378 1537 5379 1541
rect 5383 1537 5384 1541
rect 5378 1536 5384 1537
rect 5514 1541 5520 1542
rect 5514 1537 5515 1541
rect 5519 1537 5520 1541
rect 5514 1536 5520 1537
rect 5662 1540 5668 1541
rect 5662 1536 5663 1540
rect 5667 1536 5668 1540
rect 3838 1535 3844 1536
rect 3798 1492 3804 1493
rect 1974 1488 1975 1492
rect 1979 1488 1980 1492
rect 1974 1487 1980 1488
rect 1994 1491 2000 1492
rect 1994 1487 1995 1491
rect 1999 1487 2000 1491
rect 1994 1486 2000 1487
rect 2130 1491 2136 1492
rect 2130 1487 2131 1491
rect 2135 1487 2136 1491
rect 2130 1486 2136 1487
rect 2266 1491 2272 1492
rect 2266 1487 2267 1491
rect 2271 1487 2272 1491
rect 2266 1486 2272 1487
rect 2402 1491 2408 1492
rect 2402 1487 2403 1491
rect 2407 1487 2408 1491
rect 2402 1486 2408 1487
rect 2538 1491 2544 1492
rect 2538 1487 2539 1491
rect 2543 1487 2544 1491
rect 2538 1486 2544 1487
rect 2674 1491 2680 1492
rect 2674 1487 2675 1491
rect 2679 1487 2680 1491
rect 2674 1486 2680 1487
rect 2810 1491 2816 1492
rect 2810 1487 2811 1491
rect 2815 1487 2816 1491
rect 2810 1486 2816 1487
rect 2946 1491 2952 1492
rect 2946 1487 2947 1491
rect 2951 1487 2952 1491
rect 2946 1486 2952 1487
rect 3082 1491 3088 1492
rect 3082 1487 3083 1491
rect 3087 1487 3088 1491
rect 3082 1486 3088 1487
rect 3218 1491 3224 1492
rect 3218 1487 3219 1491
rect 3223 1487 3224 1491
rect 3218 1486 3224 1487
rect 3354 1491 3360 1492
rect 3354 1487 3355 1491
rect 3359 1487 3360 1491
rect 3354 1486 3360 1487
rect 3490 1491 3496 1492
rect 3490 1487 3491 1491
rect 3495 1487 3496 1491
rect 3798 1488 3799 1492
rect 3803 1488 3804 1492
rect 3798 1487 3804 1488
rect 3490 1486 3496 1487
rect 2022 1476 2028 1477
rect 1974 1475 1980 1476
rect 1974 1471 1975 1475
rect 1979 1471 1980 1475
rect 2022 1472 2023 1476
rect 2027 1472 2028 1476
rect 2022 1471 2028 1472
rect 2158 1476 2164 1477
rect 2158 1472 2159 1476
rect 2163 1472 2164 1476
rect 2158 1471 2164 1472
rect 2294 1476 2300 1477
rect 2294 1472 2295 1476
rect 2299 1472 2300 1476
rect 2294 1471 2300 1472
rect 2430 1476 2436 1477
rect 2430 1472 2431 1476
rect 2435 1472 2436 1476
rect 2430 1471 2436 1472
rect 2566 1476 2572 1477
rect 2566 1472 2567 1476
rect 2571 1472 2572 1476
rect 2566 1471 2572 1472
rect 2702 1476 2708 1477
rect 2702 1472 2703 1476
rect 2707 1472 2708 1476
rect 2702 1471 2708 1472
rect 2838 1476 2844 1477
rect 2838 1472 2839 1476
rect 2843 1472 2844 1476
rect 2838 1471 2844 1472
rect 2974 1476 2980 1477
rect 2974 1472 2975 1476
rect 2979 1472 2980 1476
rect 2974 1471 2980 1472
rect 3110 1476 3116 1477
rect 3110 1472 3111 1476
rect 3115 1472 3116 1476
rect 3110 1471 3116 1472
rect 3246 1476 3252 1477
rect 3246 1472 3247 1476
rect 3251 1472 3252 1476
rect 3246 1471 3252 1472
rect 3382 1476 3388 1477
rect 3382 1472 3383 1476
rect 3387 1472 3388 1476
rect 3382 1471 3388 1472
rect 3518 1476 3524 1477
rect 3518 1472 3519 1476
rect 3523 1472 3524 1476
rect 3518 1471 3524 1472
rect 3798 1475 3804 1476
rect 3798 1471 3799 1475
rect 3803 1471 3804 1475
rect 1974 1470 1980 1471
rect 1976 1435 1978 1470
rect 2024 1435 2026 1471
rect 2160 1435 2162 1471
rect 2296 1435 2298 1471
rect 2432 1435 2434 1471
rect 2568 1435 2570 1471
rect 2704 1435 2706 1471
rect 2840 1435 2842 1471
rect 2976 1435 2978 1471
rect 3112 1435 3114 1471
rect 3248 1435 3250 1471
rect 3384 1435 3386 1471
rect 3520 1435 3522 1471
rect 3798 1470 3804 1471
rect 3800 1435 3802 1470
rect 111 1434 115 1435
rect 111 1429 115 1430
rect 131 1434 135 1435
rect 131 1429 135 1430
rect 299 1434 303 1435
rect 299 1429 303 1430
rect 395 1434 399 1435
rect 395 1429 399 1430
rect 483 1434 487 1435
rect 483 1429 487 1430
rect 667 1434 671 1435
rect 667 1429 671 1430
rect 683 1434 687 1435
rect 683 1429 687 1430
rect 859 1434 863 1435
rect 859 1429 863 1430
rect 971 1434 975 1435
rect 971 1429 975 1430
rect 1051 1434 1055 1435
rect 1051 1429 1055 1430
rect 1259 1434 1263 1435
rect 1259 1429 1263 1430
rect 1935 1434 1939 1435
rect 1935 1429 1939 1430
rect 1975 1434 1979 1435
rect 1975 1429 1979 1430
rect 2023 1434 2027 1435
rect 2023 1429 2027 1430
rect 2159 1434 2163 1435
rect 2159 1429 2163 1430
rect 2167 1434 2171 1435
rect 2167 1429 2171 1430
rect 2295 1434 2299 1435
rect 2295 1429 2299 1430
rect 2303 1434 2307 1435
rect 2303 1429 2307 1430
rect 2431 1434 2435 1435
rect 2431 1429 2435 1430
rect 2439 1434 2443 1435
rect 2439 1429 2443 1430
rect 2567 1434 2571 1435
rect 2567 1429 2571 1430
rect 2575 1434 2579 1435
rect 2575 1429 2579 1430
rect 2703 1434 2707 1435
rect 2703 1429 2707 1430
rect 2711 1434 2715 1435
rect 2711 1429 2715 1430
rect 2839 1434 2843 1435
rect 2839 1429 2843 1430
rect 2847 1434 2851 1435
rect 2847 1429 2851 1430
rect 2975 1434 2979 1435
rect 2975 1429 2979 1430
rect 2983 1434 2987 1435
rect 2983 1429 2987 1430
rect 3111 1434 3115 1435
rect 3111 1429 3115 1430
rect 3119 1434 3123 1435
rect 3119 1429 3123 1430
rect 3247 1434 3251 1435
rect 3247 1429 3251 1430
rect 3255 1434 3259 1435
rect 3255 1429 3259 1430
rect 3383 1434 3387 1435
rect 3383 1429 3387 1430
rect 3519 1434 3523 1435
rect 3519 1429 3523 1430
rect 3799 1434 3803 1435
rect 3799 1429 3803 1430
rect 112 1369 114 1429
rect 110 1368 116 1369
rect 132 1368 134 1429
rect 396 1368 398 1429
rect 684 1368 686 1429
rect 972 1368 974 1429
rect 1260 1368 1262 1429
rect 1936 1369 1938 1429
rect 1976 1406 1978 1429
rect 1974 1405 1980 1406
rect 2168 1405 2170 1429
rect 2304 1405 2306 1429
rect 2440 1405 2442 1429
rect 2576 1405 2578 1429
rect 2712 1405 2714 1429
rect 2848 1405 2850 1429
rect 2984 1405 2986 1429
rect 3120 1405 3122 1429
rect 3256 1405 3258 1429
rect 3800 1406 3802 1429
rect 3798 1405 3804 1406
rect 1974 1401 1975 1405
rect 1979 1401 1980 1405
rect 1974 1400 1980 1401
rect 2166 1404 2172 1405
rect 2166 1400 2167 1404
rect 2171 1400 2172 1404
rect 2166 1399 2172 1400
rect 2302 1404 2308 1405
rect 2302 1400 2303 1404
rect 2307 1400 2308 1404
rect 2302 1399 2308 1400
rect 2438 1404 2444 1405
rect 2438 1400 2439 1404
rect 2443 1400 2444 1404
rect 2438 1399 2444 1400
rect 2574 1404 2580 1405
rect 2574 1400 2575 1404
rect 2579 1400 2580 1404
rect 2574 1399 2580 1400
rect 2710 1404 2716 1405
rect 2710 1400 2711 1404
rect 2715 1400 2716 1404
rect 2710 1399 2716 1400
rect 2846 1404 2852 1405
rect 2846 1400 2847 1404
rect 2851 1400 2852 1404
rect 2846 1399 2852 1400
rect 2982 1404 2988 1405
rect 2982 1400 2983 1404
rect 2987 1400 2988 1404
rect 2982 1399 2988 1400
rect 3118 1404 3124 1405
rect 3118 1400 3119 1404
rect 3123 1400 3124 1404
rect 3118 1399 3124 1400
rect 3254 1404 3260 1405
rect 3254 1400 3255 1404
rect 3259 1400 3260 1404
rect 3798 1401 3799 1405
rect 3803 1401 3804 1405
rect 3840 1403 3842 1535
rect 4564 1403 4566 1536
rect 4700 1403 4702 1536
rect 4836 1403 4838 1536
rect 4972 1403 4974 1536
rect 5108 1403 5110 1536
rect 5244 1403 5246 1536
rect 5380 1403 5382 1536
rect 5516 1403 5518 1536
rect 5662 1535 5668 1536
rect 5664 1403 5666 1535
rect 3798 1400 3804 1401
rect 3839 1402 3843 1403
rect 3254 1399 3260 1400
rect 3839 1397 3843 1398
rect 4563 1402 4567 1403
rect 4563 1397 4567 1398
rect 4699 1402 4703 1403
rect 4699 1397 4703 1398
rect 4811 1402 4815 1403
rect 4811 1397 4815 1398
rect 4835 1402 4839 1403
rect 4835 1397 4839 1398
rect 4947 1402 4951 1403
rect 4947 1397 4951 1398
rect 4971 1402 4975 1403
rect 4971 1397 4975 1398
rect 5083 1402 5087 1403
rect 5083 1397 5087 1398
rect 5107 1402 5111 1403
rect 5107 1397 5111 1398
rect 5219 1402 5223 1403
rect 5219 1397 5223 1398
rect 5243 1402 5247 1403
rect 5243 1397 5247 1398
rect 5355 1402 5359 1403
rect 5355 1397 5359 1398
rect 5379 1402 5383 1403
rect 5379 1397 5383 1398
rect 5491 1402 5495 1403
rect 5491 1397 5495 1398
rect 5515 1402 5519 1403
rect 5515 1397 5519 1398
rect 5663 1402 5667 1403
rect 5663 1397 5667 1398
rect 2138 1389 2144 1390
rect 1974 1388 1980 1389
rect 1974 1384 1975 1388
rect 1979 1384 1980 1388
rect 2138 1385 2139 1389
rect 2143 1385 2144 1389
rect 2138 1384 2144 1385
rect 2274 1389 2280 1390
rect 2274 1385 2275 1389
rect 2279 1385 2280 1389
rect 2274 1384 2280 1385
rect 2410 1389 2416 1390
rect 2410 1385 2411 1389
rect 2415 1385 2416 1389
rect 2410 1384 2416 1385
rect 2546 1389 2552 1390
rect 2546 1385 2547 1389
rect 2551 1385 2552 1389
rect 2546 1384 2552 1385
rect 2682 1389 2688 1390
rect 2682 1385 2683 1389
rect 2687 1385 2688 1389
rect 2682 1384 2688 1385
rect 2818 1389 2824 1390
rect 2818 1385 2819 1389
rect 2823 1385 2824 1389
rect 2818 1384 2824 1385
rect 2954 1389 2960 1390
rect 2954 1385 2955 1389
rect 2959 1385 2960 1389
rect 2954 1384 2960 1385
rect 3090 1389 3096 1390
rect 3090 1385 3091 1389
rect 3095 1385 3096 1389
rect 3090 1384 3096 1385
rect 3226 1389 3232 1390
rect 3226 1385 3227 1389
rect 3231 1385 3232 1389
rect 3226 1384 3232 1385
rect 3798 1388 3804 1389
rect 3798 1384 3799 1388
rect 3803 1384 3804 1388
rect 1974 1383 1980 1384
rect 1934 1368 1940 1369
rect 110 1364 111 1368
rect 115 1364 116 1368
rect 110 1363 116 1364
rect 130 1367 136 1368
rect 130 1363 131 1367
rect 135 1363 136 1367
rect 130 1362 136 1363
rect 394 1367 400 1368
rect 394 1363 395 1367
rect 399 1363 400 1367
rect 394 1362 400 1363
rect 682 1367 688 1368
rect 682 1363 683 1367
rect 687 1363 688 1367
rect 682 1362 688 1363
rect 970 1367 976 1368
rect 970 1363 971 1367
rect 975 1363 976 1367
rect 970 1362 976 1363
rect 1258 1367 1264 1368
rect 1258 1363 1259 1367
rect 1263 1363 1264 1367
rect 1934 1364 1935 1368
rect 1939 1364 1940 1368
rect 1934 1363 1940 1364
rect 1258 1362 1264 1363
rect 158 1352 164 1353
rect 110 1351 116 1352
rect 110 1347 111 1351
rect 115 1347 116 1351
rect 158 1348 159 1352
rect 163 1348 164 1352
rect 158 1347 164 1348
rect 422 1352 428 1353
rect 422 1348 423 1352
rect 427 1348 428 1352
rect 422 1347 428 1348
rect 710 1352 716 1353
rect 710 1348 711 1352
rect 715 1348 716 1352
rect 710 1347 716 1348
rect 998 1352 1004 1353
rect 998 1348 999 1352
rect 1003 1348 1004 1352
rect 998 1347 1004 1348
rect 1286 1352 1292 1353
rect 1286 1348 1287 1352
rect 1291 1348 1292 1352
rect 1286 1347 1292 1348
rect 1934 1351 1940 1352
rect 1934 1347 1935 1351
rect 1939 1347 1940 1351
rect 110 1346 116 1347
rect 112 1323 114 1346
rect 160 1323 162 1347
rect 424 1323 426 1347
rect 712 1323 714 1347
rect 1000 1323 1002 1347
rect 1288 1323 1290 1347
rect 1934 1346 1940 1347
rect 1936 1323 1938 1346
rect 1976 1323 1978 1383
rect 2140 1323 2142 1384
rect 2276 1323 2278 1384
rect 2412 1323 2414 1384
rect 2548 1323 2550 1384
rect 2684 1323 2686 1384
rect 2820 1323 2822 1384
rect 2956 1323 2958 1384
rect 3092 1323 3094 1384
rect 3228 1323 3230 1384
rect 3798 1383 3804 1384
rect 3800 1323 3802 1383
rect 3840 1337 3842 1397
rect 3838 1336 3844 1337
rect 4812 1336 4814 1397
rect 4948 1336 4950 1397
rect 5084 1336 5086 1397
rect 5220 1336 5222 1397
rect 5356 1336 5358 1397
rect 5492 1336 5494 1397
rect 5664 1337 5666 1397
rect 5662 1336 5668 1337
rect 3838 1332 3839 1336
rect 3843 1332 3844 1336
rect 3838 1331 3844 1332
rect 4810 1335 4816 1336
rect 4810 1331 4811 1335
rect 4815 1331 4816 1335
rect 4810 1330 4816 1331
rect 4946 1335 4952 1336
rect 4946 1331 4947 1335
rect 4951 1331 4952 1335
rect 4946 1330 4952 1331
rect 5082 1335 5088 1336
rect 5082 1331 5083 1335
rect 5087 1331 5088 1335
rect 5082 1330 5088 1331
rect 5218 1335 5224 1336
rect 5218 1331 5219 1335
rect 5223 1331 5224 1335
rect 5218 1330 5224 1331
rect 5354 1335 5360 1336
rect 5354 1331 5355 1335
rect 5359 1331 5360 1335
rect 5354 1330 5360 1331
rect 5490 1335 5496 1336
rect 5490 1331 5491 1335
rect 5495 1331 5496 1335
rect 5662 1332 5663 1336
rect 5667 1332 5668 1336
rect 5662 1331 5668 1332
rect 5490 1330 5496 1331
rect 111 1322 115 1323
rect 111 1317 115 1318
rect 159 1322 163 1323
rect 159 1317 163 1318
rect 423 1322 427 1323
rect 423 1317 427 1318
rect 455 1322 459 1323
rect 455 1317 459 1318
rect 711 1322 715 1323
rect 711 1317 715 1318
rect 775 1322 779 1323
rect 775 1317 779 1318
rect 999 1322 1003 1323
rect 999 1317 1003 1318
rect 1095 1322 1099 1323
rect 1095 1317 1099 1318
rect 1287 1322 1291 1323
rect 1287 1317 1291 1318
rect 1423 1322 1427 1323
rect 1423 1317 1427 1318
rect 1935 1322 1939 1323
rect 1935 1317 1939 1318
rect 1975 1322 1979 1323
rect 1975 1317 1979 1318
rect 2131 1322 2135 1323
rect 2131 1317 2135 1318
rect 2139 1322 2143 1323
rect 2139 1317 2143 1318
rect 2267 1322 2271 1323
rect 2267 1317 2271 1318
rect 2275 1322 2279 1323
rect 2275 1317 2279 1318
rect 2403 1322 2407 1323
rect 2403 1317 2407 1318
rect 2411 1322 2415 1323
rect 2411 1317 2415 1318
rect 2547 1322 2551 1323
rect 2547 1317 2551 1318
rect 2555 1322 2559 1323
rect 2555 1317 2559 1318
rect 2683 1322 2687 1323
rect 2683 1317 2687 1318
rect 2715 1322 2719 1323
rect 2715 1317 2719 1318
rect 2819 1322 2823 1323
rect 2819 1317 2823 1318
rect 2891 1322 2895 1323
rect 2891 1317 2895 1318
rect 2955 1322 2959 1323
rect 2955 1317 2959 1318
rect 3075 1322 3079 1323
rect 3075 1317 3079 1318
rect 3091 1322 3095 1323
rect 3091 1317 3095 1318
rect 3227 1322 3231 1323
rect 3227 1317 3231 1318
rect 3267 1322 3271 1323
rect 3267 1317 3271 1318
rect 3467 1322 3471 1323
rect 3467 1317 3471 1318
rect 3651 1322 3655 1323
rect 3651 1317 3655 1318
rect 3799 1322 3803 1323
rect 4838 1320 4844 1321
rect 3799 1317 3803 1318
rect 3838 1319 3844 1320
rect 112 1294 114 1317
rect 110 1293 116 1294
rect 160 1293 162 1317
rect 456 1293 458 1317
rect 776 1293 778 1317
rect 1096 1293 1098 1317
rect 1424 1293 1426 1317
rect 1936 1294 1938 1317
rect 1934 1293 1940 1294
rect 110 1289 111 1293
rect 115 1289 116 1293
rect 110 1288 116 1289
rect 158 1292 164 1293
rect 158 1288 159 1292
rect 163 1288 164 1292
rect 158 1287 164 1288
rect 454 1292 460 1293
rect 454 1288 455 1292
rect 459 1288 460 1292
rect 454 1287 460 1288
rect 774 1292 780 1293
rect 774 1288 775 1292
rect 779 1288 780 1292
rect 774 1287 780 1288
rect 1094 1292 1100 1293
rect 1094 1288 1095 1292
rect 1099 1288 1100 1292
rect 1094 1287 1100 1288
rect 1422 1292 1428 1293
rect 1422 1288 1423 1292
rect 1427 1288 1428 1292
rect 1934 1289 1935 1293
rect 1939 1289 1940 1293
rect 1934 1288 1940 1289
rect 1422 1287 1428 1288
rect 130 1277 136 1278
rect 110 1276 116 1277
rect 110 1272 111 1276
rect 115 1272 116 1276
rect 130 1273 131 1277
rect 135 1273 136 1277
rect 130 1272 136 1273
rect 426 1277 432 1278
rect 426 1273 427 1277
rect 431 1273 432 1277
rect 426 1272 432 1273
rect 746 1277 752 1278
rect 746 1273 747 1277
rect 751 1273 752 1277
rect 746 1272 752 1273
rect 1066 1277 1072 1278
rect 1066 1273 1067 1277
rect 1071 1273 1072 1277
rect 1066 1272 1072 1273
rect 1394 1277 1400 1278
rect 1394 1273 1395 1277
rect 1399 1273 1400 1277
rect 1394 1272 1400 1273
rect 1934 1276 1940 1277
rect 1934 1272 1935 1276
rect 1939 1272 1940 1276
rect 110 1271 116 1272
rect 112 1187 114 1271
rect 132 1187 134 1272
rect 428 1187 430 1272
rect 748 1187 750 1272
rect 1068 1187 1070 1272
rect 1396 1187 1398 1272
rect 1934 1271 1940 1272
rect 1936 1187 1938 1271
rect 1976 1257 1978 1317
rect 1974 1256 1980 1257
rect 2132 1256 2134 1317
rect 2268 1256 2270 1317
rect 2404 1256 2406 1317
rect 2556 1256 2558 1317
rect 2716 1256 2718 1317
rect 2892 1256 2894 1317
rect 3076 1256 3078 1317
rect 3268 1256 3270 1317
rect 3468 1256 3470 1317
rect 3652 1256 3654 1317
rect 3800 1257 3802 1317
rect 3838 1315 3839 1319
rect 3843 1315 3844 1319
rect 4838 1316 4839 1320
rect 4843 1316 4844 1320
rect 4838 1315 4844 1316
rect 4974 1320 4980 1321
rect 4974 1316 4975 1320
rect 4979 1316 4980 1320
rect 4974 1315 4980 1316
rect 5110 1320 5116 1321
rect 5110 1316 5111 1320
rect 5115 1316 5116 1320
rect 5110 1315 5116 1316
rect 5246 1320 5252 1321
rect 5246 1316 5247 1320
rect 5251 1316 5252 1320
rect 5246 1315 5252 1316
rect 5382 1320 5388 1321
rect 5382 1316 5383 1320
rect 5387 1316 5388 1320
rect 5382 1315 5388 1316
rect 5518 1320 5524 1321
rect 5518 1316 5519 1320
rect 5523 1316 5524 1320
rect 5518 1315 5524 1316
rect 5662 1319 5668 1320
rect 5662 1315 5663 1319
rect 5667 1315 5668 1319
rect 3838 1314 3844 1315
rect 3840 1287 3842 1314
rect 4840 1287 4842 1315
rect 4976 1287 4978 1315
rect 5112 1287 5114 1315
rect 5248 1287 5250 1315
rect 5384 1287 5386 1315
rect 5520 1287 5522 1315
rect 5662 1314 5668 1315
rect 5664 1287 5666 1314
rect 3839 1286 3843 1287
rect 3839 1281 3843 1282
rect 4735 1286 4739 1287
rect 4735 1281 4739 1282
rect 4839 1286 4843 1287
rect 4839 1281 4843 1282
rect 4879 1286 4883 1287
rect 4879 1281 4883 1282
rect 4975 1286 4979 1287
rect 4975 1281 4979 1282
rect 5031 1286 5035 1287
rect 5031 1281 5035 1282
rect 5111 1286 5115 1287
rect 5111 1281 5115 1282
rect 5191 1286 5195 1287
rect 5191 1281 5195 1282
rect 5247 1286 5251 1287
rect 5247 1281 5251 1282
rect 5359 1286 5363 1287
rect 5359 1281 5363 1282
rect 5383 1286 5387 1287
rect 5383 1281 5387 1282
rect 5519 1286 5523 1287
rect 5519 1281 5523 1282
rect 5527 1286 5531 1287
rect 5527 1281 5531 1282
rect 5663 1286 5667 1287
rect 5663 1281 5667 1282
rect 3840 1258 3842 1281
rect 3838 1257 3844 1258
rect 4736 1257 4738 1281
rect 4880 1257 4882 1281
rect 5032 1257 5034 1281
rect 5192 1257 5194 1281
rect 5360 1257 5362 1281
rect 5528 1257 5530 1281
rect 5664 1258 5666 1281
rect 5662 1257 5668 1258
rect 3798 1256 3804 1257
rect 1974 1252 1975 1256
rect 1979 1252 1980 1256
rect 1974 1251 1980 1252
rect 2130 1255 2136 1256
rect 2130 1251 2131 1255
rect 2135 1251 2136 1255
rect 2130 1250 2136 1251
rect 2266 1255 2272 1256
rect 2266 1251 2267 1255
rect 2271 1251 2272 1255
rect 2266 1250 2272 1251
rect 2402 1255 2408 1256
rect 2402 1251 2403 1255
rect 2407 1251 2408 1255
rect 2402 1250 2408 1251
rect 2554 1255 2560 1256
rect 2554 1251 2555 1255
rect 2559 1251 2560 1255
rect 2554 1250 2560 1251
rect 2714 1255 2720 1256
rect 2714 1251 2715 1255
rect 2719 1251 2720 1255
rect 2714 1250 2720 1251
rect 2890 1255 2896 1256
rect 2890 1251 2891 1255
rect 2895 1251 2896 1255
rect 2890 1250 2896 1251
rect 3074 1255 3080 1256
rect 3074 1251 3075 1255
rect 3079 1251 3080 1255
rect 3074 1250 3080 1251
rect 3266 1255 3272 1256
rect 3266 1251 3267 1255
rect 3271 1251 3272 1255
rect 3266 1250 3272 1251
rect 3466 1255 3472 1256
rect 3466 1251 3467 1255
rect 3471 1251 3472 1255
rect 3466 1250 3472 1251
rect 3650 1255 3656 1256
rect 3650 1251 3651 1255
rect 3655 1251 3656 1255
rect 3798 1252 3799 1256
rect 3803 1252 3804 1256
rect 3838 1253 3839 1257
rect 3843 1253 3844 1257
rect 3838 1252 3844 1253
rect 4734 1256 4740 1257
rect 4734 1252 4735 1256
rect 4739 1252 4740 1256
rect 3798 1251 3804 1252
rect 4734 1251 4740 1252
rect 4878 1256 4884 1257
rect 4878 1252 4879 1256
rect 4883 1252 4884 1256
rect 4878 1251 4884 1252
rect 5030 1256 5036 1257
rect 5030 1252 5031 1256
rect 5035 1252 5036 1256
rect 5030 1251 5036 1252
rect 5190 1256 5196 1257
rect 5190 1252 5191 1256
rect 5195 1252 5196 1256
rect 5190 1251 5196 1252
rect 5358 1256 5364 1257
rect 5358 1252 5359 1256
rect 5363 1252 5364 1256
rect 5358 1251 5364 1252
rect 5526 1256 5532 1257
rect 5526 1252 5527 1256
rect 5531 1252 5532 1256
rect 5662 1253 5663 1257
rect 5667 1253 5668 1257
rect 5662 1252 5668 1253
rect 5526 1251 5532 1252
rect 3650 1250 3656 1251
rect 4706 1241 4712 1242
rect 2158 1240 2164 1241
rect 1974 1239 1980 1240
rect 1974 1235 1975 1239
rect 1979 1235 1980 1239
rect 2158 1236 2159 1240
rect 2163 1236 2164 1240
rect 2158 1235 2164 1236
rect 2294 1240 2300 1241
rect 2294 1236 2295 1240
rect 2299 1236 2300 1240
rect 2294 1235 2300 1236
rect 2430 1240 2436 1241
rect 2430 1236 2431 1240
rect 2435 1236 2436 1240
rect 2430 1235 2436 1236
rect 2582 1240 2588 1241
rect 2582 1236 2583 1240
rect 2587 1236 2588 1240
rect 2582 1235 2588 1236
rect 2742 1240 2748 1241
rect 2742 1236 2743 1240
rect 2747 1236 2748 1240
rect 2742 1235 2748 1236
rect 2918 1240 2924 1241
rect 2918 1236 2919 1240
rect 2923 1236 2924 1240
rect 2918 1235 2924 1236
rect 3102 1240 3108 1241
rect 3102 1236 3103 1240
rect 3107 1236 3108 1240
rect 3102 1235 3108 1236
rect 3294 1240 3300 1241
rect 3294 1236 3295 1240
rect 3299 1236 3300 1240
rect 3294 1235 3300 1236
rect 3494 1240 3500 1241
rect 3494 1236 3495 1240
rect 3499 1236 3500 1240
rect 3494 1235 3500 1236
rect 3678 1240 3684 1241
rect 3838 1240 3844 1241
rect 3678 1236 3679 1240
rect 3683 1236 3684 1240
rect 3678 1235 3684 1236
rect 3798 1239 3804 1240
rect 3798 1235 3799 1239
rect 3803 1235 3804 1239
rect 3838 1236 3839 1240
rect 3843 1236 3844 1240
rect 4706 1237 4707 1241
rect 4711 1237 4712 1241
rect 4706 1236 4712 1237
rect 4850 1241 4856 1242
rect 4850 1237 4851 1241
rect 4855 1237 4856 1241
rect 4850 1236 4856 1237
rect 5002 1241 5008 1242
rect 5002 1237 5003 1241
rect 5007 1237 5008 1241
rect 5002 1236 5008 1237
rect 5162 1241 5168 1242
rect 5162 1237 5163 1241
rect 5167 1237 5168 1241
rect 5162 1236 5168 1237
rect 5330 1241 5336 1242
rect 5330 1237 5331 1241
rect 5335 1237 5336 1241
rect 5330 1236 5336 1237
rect 5498 1241 5504 1242
rect 5498 1237 5499 1241
rect 5503 1237 5504 1241
rect 5498 1236 5504 1237
rect 5662 1240 5668 1241
rect 5662 1236 5663 1240
rect 5667 1236 5668 1240
rect 3838 1235 3844 1236
rect 1974 1234 1980 1235
rect 1976 1211 1978 1234
rect 2160 1211 2162 1235
rect 2296 1211 2298 1235
rect 2432 1211 2434 1235
rect 2584 1211 2586 1235
rect 2744 1211 2746 1235
rect 2920 1211 2922 1235
rect 3104 1211 3106 1235
rect 3296 1211 3298 1235
rect 3496 1211 3498 1235
rect 3680 1211 3682 1235
rect 3798 1234 3804 1235
rect 3800 1211 3802 1234
rect 1975 1210 1979 1211
rect 1975 1205 1979 1206
rect 2023 1210 2027 1211
rect 2023 1205 2027 1206
rect 2159 1210 2163 1211
rect 2159 1205 2163 1206
rect 2239 1210 2243 1211
rect 2239 1205 2243 1206
rect 2295 1210 2299 1211
rect 2295 1205 2299 1206
rect 2431 1210 2435 1211
rect 2431 1205 2435 1206
rect 2479 1210 2483 1211
rect 2479 1205 2483 1206
rect 2583 1210 2587 1211
rect 2583 1205 2587 1206
rect 2719 1210 2723 1211
rect 2719 1205 2723 1206
rect 2743 1210 2747 1211
rect 2743 1205 2747 1206
rect 2919 1210 2923 1211
rect 2919 1205 2923 1206
rect 2959 1210 2963 1211
rect 2959 1205 2963 1206
rect 3103 1210 3107 1211
rect 3103 1205 3107 1206
rect 3207 1210 3211 1211
rect 3207 1205 3211 1206
rect 3295 1210 3299 1211
rect 3295 1205 3299 1206
rect 3455 1210 3459 1211
rect 3455 1205 3459 1206
rect 3495 1210 3499 1211
rect 3495 1205 3499 1206
rect 3679 1210 3683 1211
rect 3679 1205 3683 1206
rect 3799 1210 3803 1211
rect 3799 1205 3803 1206
rect 111 1186 115 1187
rect 111 1181 115 1182
rect 131 1186 135 1187
rect 131 1181 135 1182
rect 331 1186 335 1187
rect 331 1181 335 1182
rect 427 1186 431 1187
rect 427 1181 431 1182
rect 563 1186 567 1187
rect 563 1181 567 1182
rect 747 1186 751 1187
rect 747 1181 751 1182
rect 803 1186 807 1187
rect 803 1181 807 1182
rect 1043 1186 1047 1187
rect 1043 1181 1047 1182
rect 1067 1186 1071 1187
rect 1067 1181 1071 1182
rect 1283 1186 1287 1187
rect 1283 1181 1287 1182
rect 1395 1186 1399 1187
rect 1395 1181 1399 1182
rect 1523 1186 1527 1187
rect 1523 1181 1527 1182
rect 1771 1186 1775 1187
rect 1771 1181 1775 1182
rect 1935 1186 1939 1187
rect 1976 1182 1978 1205
rect 1935 1181 1939 1182
rect 1974 1181 1980 1182
rect 2024 1181 2026 1205
rect 2240 1181 2242 1205
rect 2480 1181 2482 1205
rect 2720 1181 2722 1205
rect 2960 1181 2962 1205
rect 3208 1181 3210 1205
rect 3456 1181 3458 1205
rect 3680 1181 3682 1205
rect 3800 1182 3802 1205
rect 3798 1181 3804 1182
rect 112 1121 114 1181
rect 110 1120 116 1121
rect 132 1120 134 1181
rect 332 1120 334 1181
rect 564 1120 566 1181
rect 804 1120 806 1181
rect 1044 1120 1046 1181
rect 1284 1120 1286 1181
rect 1524 1120 1526 1181
rect 1772 1120 1774 1181
rect 1936 1121 1938 1181
rect 1974 1177 1975 1181
rect 1979 1177 1980 1181
rect 1974 1176 1980 1177
rect 2022 1180 2028 1181
rect 2022 1176 2023 1180
rect 2027 1176 2028 1180
rect 2022 1175 2028 1176
rect 2238 1180 2244 1181
rect 2238 1176 2239 1180
rect 2243 1176 2244 1180
rect 2238 1175 2244 1176
rect 2478 1180 2484 1181
rect 2478 1176 2479 1180
rect 2483 1176 2484 1180
rect 2478 1175 2484 1176
rect 2718 1180 2724 1181
rect 2718 1176 2719 1180
rect 2723 1176 2724 1180
rect 2718 1175 2724 1176
rect 2958 1180 2964 1181
rect 2958 1176 2959 1180
rect 2963 1176 2964 1180
rect 2958 1175 2964 1176
rect 3206 1180 3212 1181
rect 3206 1176 3207 1180
rect 3211 1176 3212 1180
rect 3206 1175 3212 1176
rect 3454 1180 3460 1181
rect 3454 1176 3455 1180
rect 3459 1176 3460 1180
rect 3454 1175 3460 1176
rect 3678 1180 3684 1181
rect 3678 1176 3679 1180
rect 3683 1176 3684 1180
rect 3798 1177 3799 1181
rect 3803 1177 3804 1181
rect 3798 1176 3804 1177
rect 3678 1175 3684 1176
rect 3840 1167 3842 1235
rect 4708 1167 4710 1236
rect 4852 1167 4854 1236
rect 5004 1167 5006 1236
rect 5164 1167 5166 1236
rect 5332 1167 5334 1236
rect 5500 1167 5502 1236
rect 5662 1235 5668 1236
rect 5664 1167 5666 1235
rect 3839 1166 3843 1167
rect 1994 1165 2000 1166
rect 1974 1164 1980 1165
rect 1974 1160 1975 1164
rect 1979 1160 1980 1164
rect 1994 1161 1995 1165
rect 1999 1161 2000 1165
rect 1994 1160 2000 1161
rect 2210 1165 2216 1166
rect 2210 1161 2211 1165
rect 2215 1161 2216 1165
rect 2210 1160 2216 1161
rect 2450 1165 2456 1166
rect 2450 1161 2451 1165
rect 2455 1161 2456 1165
rect 2450 1160 2456 1161
rect 2690 1165 2696 1166
rect 2690 1161 2691 1165
rect 2695 1161 2696 1165
rect 2690 1160 2696 1161
rect 2930 1165 2936 1166
rect 2930 1161 2931 1165
rect 2935 1161 2936 1165
rect 2930 1160 2936 1161
rect 3178 1165 3184 1166
rect 3178 1161 3179 1165
rect 3183 1161 3184 1165
rect 3178 1160 3184 1161
rect 3426 1165 3432 1166
rect 3426 1161 3427 1165
rect 3431 1161 3432 1165
rect 3426 1160 3432 1161
rect 3650 1165 3656 1166
rect 3650 1161 3651 1165
rect 3655 1161 3656 1165
rect 3650 1160 3656 1161
rect 3798 1164 3804 1165
rect 3798 1160 3799 1164
rect 3803 1160 3804 1164
rect 3839 1161 3843 1162
rect 3859 1166 3863 1167
rect 3859 1161 3863 1162
rect 4067 1166 4071 1167
rect 4067 1161 4071 1162
rect 4299 1166 4303 1167
rect 4299 1161 4303 1162
rect 4539 1166 4543 1167
rect 4539 1161 4543 1162
rect 4707 1166 4711 1167
rect 4707 1161 4711 1162
rect 4779 1166 4783 1167
rect 4779 1161 4783 1162
rect 4851 1166 4855 1167
rect 4851 1161 4855 1162
rect 5003 1166 5007 1167
rect 5003 1161 5007 1162
rect 5027 1166 5031 1167
rect 5027 1161 5031 1162
rect 5163 1166 5167 1167
rect 5163 1161 5167 1162
rect 5283 1166 5287 1167
rect 5283 1161 5287 1162
rect 5331 1166 5335 1167
rect 5331 1161 5335 1162
rect 5499 1166 5503 1167
rect 5499 1161 5503 1162
rect 5515 1166 5519 1167
rect 5515 1161 5519 1162
rect 5663 1166 5667 1167
rect 5663 1161 5667 1162
rect 1974 1159 1980 1160
rect 1934 1120 1940 1121
rect 110 1116 111 1120
rect 115 1116 116 1120
rect 110 1115 116 1116
rect 130 1119 136 1120
rect 130 1115 131 1119
rect 135 1115 136 1119
rect 130 1114 136 1115
rect 330 1119 336 1120
rect 330 1115 331 1119
rect 335 1115 336 1119
rect 330 1114 336 1115
rect 562 1119 568 1120
rect 562 1115 563 1119
rect 567 1115 568 1119
rect 562 1114 568 1115
rect 802 1119 808 1120
rect 802 1115 803 1119
rect 807 1115 808 1119
rect 802 1114 808 1115
rect 1042 1119 1048 1120
rect 1042 1115 1043 1119
rect 1047 1115 1048 1119
rect 1042 1114 1048 1115
rect 1282 1119 1288 1120
rect 1282 1115 1283 1119
rect 1287 1115 1288 1119
rect 1282 1114 1288 1115
rect 1522 1119 1528 1120
rect 1522 1115 1523 1119
rect 1527 1115 1528 1119
rect 1522 1114 1528 1115
rect 1770 1119 1776 1120
rect 1770 1115 1771 1119
rect 1775 1115 1776 1119
rect 1934 1116 1935 1120
rect 1939 1116 1940 1120
rect 1934 1115 1940 1116
rect 1770 1114 1776 1115
rect 158 1104 164 1105
rect 110 1103 116 1104
rect 110 1099 111 1103
rect 115 1099 116 1103
rect 158 1100 159 1104
rect 163 1100 164 1104
rect 158 1099 164 1100
rect 358 1104 364 1105
rect 358 1100 359 1104
rect 363 1100 364 1104
rect 358 1099 364 1100
rect 590 1104 596 1105
rect 590 1100 591 1104
rect 595 1100 596 1104
rect 590 1099 596 1100
rect 830 1104 836 1105
rect 830 1100 831 1104
rect 835 1100 836 1104
rect 830 1099 836 1100
rect 1070 1104 1076 1105
rect 1070 1100 1071 1104
rect 1075 1100 1076 1104
rect 1070 1099 1076 1100
rect 1310 1104 1316 1105
rect 1310 1100 1311 1104
rect 1315 1100 1316 1104
rect 1310 1099 1316 1100
rect 1550 1104 1556 1105
rect 1550 1100 1551 1104
rect 1555 1100 1556 1104
rect 1550 1099 1556 1100
rect 1798 1104 1804 1105
rect 1798 1100 1799 1104
rect 1803 1100 1804 1104
rect 1798 1099 1804 1100
rect 1934 1103 1940 1104
rect 1934 1099 1935 1103
rect 1939 1099 1940 1103
rect 110 1098 116 1099
rect 112 1075 114 1098
rect 160 1075 162 1099
rect 360 1075 362 1099
rect 592 1075 594 1099
rect 832 1075 834 1099
rect 1072 1075 1074 1099
rect 1312 1075 1314 1099
rect 1552 1075 1554 1099
rect 1800 1075 1802 1099
rect 1934 1098 1940 1099
rect 1936 1075 1938 1098
rect 1976 1075 1978 1159
rect 1996 1075 1998 1160
rect 2212 1075 2214 1160
rect 2452 1075 2454 1160
rect 2692 1075 2694 1160
rect 2932 1075 2934 1160
rect 3180 1075 3182 1160
rect 3428 1075 3430 1160
rect 3652 1075 3654 1160
rect 3798 1159 3804 1160
rect 3800 1075 3802 1159
rect 3840 1101 3842 1161
rect 3838 1100 3844 1101
rect 3860 1100 3862 1161
rect 4068 1100 4070 1161
rect 4300 1100 4302 1161
rect 4540 1100 4542 1161
rect 4780 1100 4782 1161
rect 5028 1100 5030 1161
rect 5284 1100 5286 1161
rect 5516 1100 5518 1161
rect 5664 1101 5666 1161
rect 5662 1100 5668 1101
rect 3838 1096 3839 1100
rect 3843 1096 3844 1100
rect 3838 1095 3844 1096
rect 3858 1099 3864 1100
rect 3858 1095 3859 1099
rect 3863 1095 3864 1099
rect 3858 1094 3864 1095
rect 4066 1099 4072 1100
rect 4066 1095 4067 1099
rect 4071 1095 4072 1099
rect 4066 1094 4072 1095
rect 4298 1099 4304 1100
rect 4298 1095 4299 1099
rect 4303 1095 4304 1099
rect 4298 1094 4304 1095
rect 4538 1099 4544 1100
rect 4538 1095 4539 1099
rect 4543 1095 4544 1099
rect 4538 1094 4544 1095
rect 4778 1099 4784 1100
rect 4778 1095 4779 1099
rect 4783 1095 4784 1099
rect 4778 1094 4784 1095
rect 5026 1099 5032 1100
rect 5026 1095 5027 1099
rect 5031 1095 5032 1099
rect 5026 1094 5032 1095
rect 5282 1099 5288 1100
rect 5282 1095 5283 1099
rect 5287 1095 5288 1099
rect 5282 1094 5288 1095
rect 5514 1099 5520 1100
rect 5514 1095 5515 1099
rect 5519 1095 5520 1099
rect 5662 1096 5663 1100
rect 5667 1096 5668 1100
rect 5662 1095 5668 1096
rect 5514 1094 5520 1095
rect 3886 1084 3892 1085
rect 3838 1083 3844 1084
rect 3838 1079 3839 1083
rect 3843 1079 3844 1083
rect 3886 1080 3887 1084
rect 3891 1080 3892 1084
rect 3886 1079 3892 1080
rect 4094 1084 4100 1085
rect 4094 1080 4095 1084
rect 4099 1080 4100 1084
rect 4094 1079 4100 1080
rect 4326 1084 4332 1085
rect 4326 1080 4327 1084
rect 4331 1080 4332 1084
rect 4326 1079 4332 1080
rect 4566 1084 4572 1085
rect 4566 1080 4567 1084
rect 4571 1080 4572 1084
rect 4566 1079 4572 1080
rect 4806 1084 4812 1085
rect 4806 1080 4807 1084
rect 4811 1080 4812 1084
rect 4806 1079 4812 1080
rect 5054 1084 5060 1085
rect 5054 1080 5055 1084
rect 5059 1080 5060 1084
rect 5054 1079 5060 1080
rect 5310 1084 5316 1085
rect 5310 1080 5311 1084
rect 5315 1080 5316 1084
rect 5310 1079 5316 1080
rect 5542 1084 5548 1085
rect 5542 1080 5543 1084
rect 5547 1080 5548 1084
rect 5542 1079 5548 1080
rect 5662 1083 5668 1084
rect 5662 1079 5663 1083
rect 5667 1079 5668 1083
rect 3838 1078 3844 1079
rect 111 1074 115 1075
rect 111 1069 115 1070
rect 159 1074 163 1075
rect 159 1069 163 1070
rect 263 1074 267 1075
rect 263 1069 267 1070
rect 359 1074 363 1075
rect 359 1069 363 1070
rect 439 1074 443 1075
rect 439 1069 443 1070
rect 591 1074 595 1075
rect 591 1069 595 1070
rect 615 1074 619 1075
rect 615 1069 619 1070
rect 783 1074 787 1075
rect 783 1069 787 1070
rect 831 1074 835 1075
rect 831 1069 835 1070
rect 951 1074 955 1075
rect 951 1069 955 1070
rect 1071 1074 1075 1075
rect 1071 1069 1075 1070
rect 1111 1074 1115 1075
rect 1111 1069 1115 1070
rect 1271 1074 1275 1075
rect 1271 1069 1275 1070
rect 1311 1074 1315 1075
rect 1311 1069 1315 1070
rect 1431 1074 1435 1075
rect 1431 1069 1435 1070
rect 1551 1074 1555 1075
rect 1551 1069 1555 1070
rect 1591 1074 1595 1075
rect 1591 1069 1595 1070
rect 1751 1074 1755 1075
rect 1751 1069 1755 1070
rect 1799 1074 1803 1075
rect 1799 1069 1803 1070
rect 1935 1074 1939 1075
rect 1935 1069 1939 1070
rect 1975 1074 1979 1075
rect 1975 1069 1979 1070
rect 1995 1074 1999 1075
rect 1995 1069 1999 1070
rect 2211 1074 2215 1075
rect 2211 1069 2215 1070
rect 2451 1074 2455 1075
rect 2451 1069 2455 1070
rect 2691 1074 2695 1075
rect 2691 1069 2695 1070
rect 2931 1074 2935 1075
rect 2931 1069 2935 1070
rect 3091 1074 3095 1075
rect 3091 1069 3095 1070
rect 3179 1074 3183 1075
rect 3179 1069 3183 1070
rect 3243 1074 3247 1075
rect 3243 1069 3247 1070
rect 3395 1074 3399 1075
rect 3395 1069 3399 1070
rect 3427 1074 3431 1075
rect 3427 1069 3431 1070
rect 3651 1074 3655 1075
rect 3651 1069 3655 1070
rect 3799 1074 3803 1075
rect 3799 1069 3803 1070
rect 112 1046 114 1069
rect 110 1045 116 1046
rect 264 1045 266 1069
rect 440 1045 442 1069
rect 616 1045 618 1069
rect 784 1045 786 1069
rect 952 1045 954 1069
rect 1112 1045 1114 1069
rect 1272 1045 1274 1069
rect 1432 1045 1434 1069
rect 1592 1045 1594 1069
rect 1752 1045 1754 1069
rect 1936 1046 1938 1069
rect 1934 1045 1940 1046
rect 110 1041 111 1045
rect 115 1041 116 1045
rect 110 1040 116 1041
rect 262 1044 268 1045
rect 262 1040 263 1044
rect 267 1040 268 1044
rect 262 1039 268 1040
rect 438 1044 444 1045
rect 438 1040 439 1044
rect 443 1040 444 1044
rect 438 1039 444 1040
rect 614 1044 620 1045
rect 614 1040 615 1044
rect 619 1040 620 1044
rect 614 1039 620 1040
rect 782 1044 788 1045
rect 782 1040 783 1044
rect 787 1040 788 1044
rect 782 1039 788 1040
rect 950 1044 956 1045
rect 950 1040 951 1044
rect 955 1040 956 1044
rect 950 1039 956 1040
rect 1110 1044 1116 1045
rect 1110 1040 1111 1044
rect 1115 1040 1116 1044
rect 1110 1039 1116 1040
rect 1270 1044 1276 1045
rect 1270 1040 1271 1044
rect 1275 1040 1276 1044
rect 1270 1039 1276 1040
rect 1430 1044 1436 1045
rect 1430 1040 1431 1044
rect 1435 1040 1436 1044
rect 1430 1039 1436 1040
rect 1590 1044 1596 1045
rect 1590 1040 1591 1044
rect 1595 1040 1596 1044
rect 1590 1039 1596 1040
rect 1750 1044 1756 1045
rect 1750 1040 1751 1044
rect 1755 1040 1756 1044
rect 1934 1041 1935 1045
rect 1939 1041 1940 1045
rect 1934 1040 1940 1041
rect 1750 1039 1756 1040
rect 234 1029 240 1030
rect 110 1028 116 1029
rect 110 1024 111 1028
rect 115 1024 116 1028
rect 234 1025 235 1029
rect 239 1025 240 1029
rect 234 1024 240 1025
rect 410 1029 416 1030
rect 410 1025 411 1029
rect 415 1025 416 1029
rect 410 1024 416 1025
rect 586 1029 592 1030
rect 586 1025 587 1029
rect 591 1025 592 1029
rect 586 1024 592 1025
rect 754 1029 760 1030
rect 754 1025 755 1029
rect 759 1025 760 1029
rect 754 1024 760 1025
rect 922 1029 928 1030
rect 922 1025 923 1029
rect 927 1025 928 1029
rect 922 1024 928 1025
rect 1082 1029 1088 1030
rect 1082 1025 1083 1029
rect 1087 1025 1088 1029
rect 1082 1024 1088 1025
rect 1242 1029 1248 1030
rect 1242 1025 1243 1029
rect 1247 1025 1248 1029
rect 1242 1024 1248 1025
rect 1402 1029 1408 1030
rect 1402 1025 1403 1029
rect 1407 1025 1408 1029
rect 1402 1024 1408 1025
rect 1562 1029 1568 1030
rect 1562 1025 1563 1029
rect 1567 1025 1568 1029
rect 1562 1024 1568 1025
rect 1722 1029 1728 1030
rect 1722 1025 1723 1029
rect 1727 1025 1728 1029
rect 1722 1024 1728 1025
rect 1934 1028 1940 1029
rect 1934 1024 1935 1028
rect 1939 1024 1940 1028
rect 110 1023 116 1024
rect 112 959 114 1023
rect 236 959 238 1024
rect 412 959 414 1024
rect 588 959 590 1024
rect 756 959 758 1024
rect 924 959 926 1024
rect 1084 959 1086 1024
rect 1244 959 1246 1024
rect 1404 959 1406 1024
rect 1564 959 1566 1024
rect 1724 959 1726 1024
rect 1934 1023 1940 1024
rect 1936 959 1938 1023
rect 1976 1009 1978 1069
rect 1974 1008 1980 1009
rect 3092 1008 3094 1069
rect 3244 1008 3246 1069
rect 3396 1008 3398 1069
rect 3800 1009 3802 1069
rect 3840 1055 3842 1078
rect 3888 1055 3890 1079
rect 4096 1055 4098 1079
rect 4328 1055 4330 1079
rect 4568 1055 4570 1079
rect 4808 1055 4810 1079
rect 5056 1055 5058 1079
rect 5312 1055 5314 1079
rect 5544 1055 5546 1079
rect 5662 1078 5668 1079
rect 5664 1055 5666 1078
rect 3839 1054 3843 1055
rect 3839 1049 3843 1050
rect 3887 1054 3891 1055
rect 3887 1049 3891 1050
rect 4071 1054 4075 1055
rect 4071 1049 4075 1050
rect 4095 1054 4099 1055
rect 4095 1049 4099 1050
rect 4279 1054 4283 1055
rect 4279 1049 4283 1050
rect 4327 1054 4331 1055
rect 4327 1049 4331 1050
rect 4511 1054 4515 1055
rect 4511 1049 4515 1050
rect 4567 1054 4571 1055
rect 4567 1049 4571 1050
rect 4759 1054 4763 1055
rect 4759 1049 4763 1050
rect 4807 1054 4811 1055
rect 4807 1049 4811 1050
rect 5023 1054 5027 1055
rect 5023 1049 5027 1050
rect 5055 1054 5059 1055
rect 5055 1049 5059 1050
rect 5295 1054 5299 1055
rect 5295 1049 5299 1050
rect 5311 1054 5315 1055
rect 5311 1049 5315 1050
rect 5543 1054 5547 1055
rect 5543 1049 5547 1050
rect 5663 1054 5667 1055
rect 5663 1049 5667 1050
rect 3840 1026 3842 1049
rect 3838 1025 3844 1026
rect 3888 1025 3890 1049
rect 4072 1025 4074 1049
rect 4280 1025 4282 1049
rect 4512 1025 4514 1049
rect 4760 1025 4762 1049
rect 5024 1025 5026 1049
rect 5296 1025 5298 1049
rect 5544 1025 5546 1049
rect 5664 1026 5666 1049
rect 5662 1025 5668 1026
rect 3838 1021 3839 1025
rect 3843 1021 3844 1025
rect 3838 1020 3844 1021
rect 3886 1024 3892 1025
rect 3886 1020 3887 1024
rect 3891 1020 3892 1024
rect 3886 1019 3892 1020
rect 4070 1024 4076 1025
rect 4070 1020 4071 1024
rect 4075 1020 4076 1024
rect 4070 1019 4076 1020
rect 4278 1024 4284 1025
rect 4278 1020 4279 1024
rect 4283 1020 4284 1024
rect 4278 1019 4284 1020
rect 4510 1024 4516 1025
rect 4510 1020 4511 1024
rect 4515 1020 4516 1024
rect 4510 1019 4516 1020
rect 4758 1024 4764 1025
rect 4758 1020 4759 1024
rect 4763 1020 4764 1024
rect 4758 1019 4764 1020
rect 5022 1024 5028 1025
rect 5022 1020 5023 1024
rect 5027 1020 5028 1024
rect 5022 1019 5028 1020
rect 5294 1024 5300 1025
rect 5294 1020 5295 1024
rect 5299 1020 5300 1024
rect 5294 1019 5300 1020
rect 5542 1024 5548 1025
rect 5542 1020 5543 1024
rect 5547 1020 5548 1024
rect 5662 1021 5663 1025
rect 5667 1021 5668 1025
rect 5662 1020 5668 1021
rect 5542 1019 5548 1020
rect 3858 1009 3864 1010
rect 3798 1008 3804 1009
rect 1974 1004 1975 1008
rect 1979 1004 1980 1008
rect 1974 1003 1980 1004
rect 3090 1007 3096 1008
rect 3090 1003 3091 1007
rect 3095 1003 3096 1007
rect 3090 1002 3096 1003
rect 3242 1007 3248 1008
rect 3242 1003 3243 1007
rect 3247 1003 3248 1007
rect 3242 1002 3248 1003
rect 3394 1007 3400 1008
rect 3394 1003 3395 1007
rect 3399 1003 3400 1007
rect 3798 1004 3799 1008
rect 3803 1004 3804 1008
rect 3798 1003 3804 1004
rect 3838 1008 3844 1009
rect 3838 1004 3839 1008
rect 3843 1004 3844 1008
rect 3858 1005 3859 1009
rect 3863 1005 3864 1009
rect 3858 1004 3864 1005
rect 4042 1009 4048 1010
rect 4042 1005 4043 1009
rect 4047 1005 4048 1009
rect 4042 1004 4048 1005
rect 4250 1009 4256 1010
rect 4250 1005 4251 1009
rect 4255 1005 4256 1009
rect 4250 1004 4256 1005
rect 4482 1009 4488 1010
rect 4482 1005 4483 1009
rect 4487 1005 4488 1009
rect 4482 1004 4488 1005
rect 4730 1009 4736 1010
rect 4730 1005 4731 1009
rect 4735 1005 4736 1009
rect 4730 1004 4736 1005
rect 4994 1009 5000 1010
rect 4994 1005 4995 1009
rect 4999 1005 5000 1009
rect 4994 1004 5000 1005
rect 5266 1009 5272 1010
rect 5266 1005 5267 1009
rect 5271 1005 5272 1009
rect 5266 1004 5272 1005
rect 5514 1009 5520 1010
rect 5514 1005 5515 1009
rect 5519 1005 5520 1009
rect 5514 1004 5520 1005
rect 5662 1008 5668 1009
rect 5662 1004 5663 1008
rect 5667 1004 5668 1008
rect 3838 1003 3844 1004
rect 3394 1002 3400 1003
rect 3118 992 3124 993
rect 1974 991 1980 992
rect 1974 987 1975 991
rect 1979 987 1980 991
rect 3118 988 3119 992
rect 3123 988 3124 992
rect 3118 987 3124 988
rect 3270 992 3276 993
rect 3270 988 3271 992
rect 3275 988 3276 992
rect 3270 987 3276 988
rect 3422 992 3428 993
rect 3422 988 3423 992
rect 3427 988 3428 992
rect 3422 987 3428 988
rect 3798 991 3804 992
rect 3798 987 3799 991
rect 3803 987 3804 991
rect 1974 986 1980 987
rect 111 958 115 959
rect 111 953 115 954
rect 227 958 231 959
rect 227 953 231 954
rect 235 958 239 959
rect 235 953 239 954
rect 379 958 383 959
rect 379 953 383 954
rect 411 958 415 959
rect 411 953 415 954
rect 539 958 543 959
rect 539 953 543 954
rect 587 958 591 959
rect 587 953 591 954
rect 715 958 719 959
rect 715 953 719 954
rect 755 958 759 959
rect 755 953 759 954
rect 891 958 895 959
rect 891 953 895 954
rect 923 958 927 959
rect 923 953 927 954
rect 1075 958 1079 959
rect 1075 953 1079 954
rect 1083 958 1087 959
rect 1083 953 1087 954
rect 1243 958 1247 959
rect 1243 953 1247 954
rect 1259 958 1263 959
rect 1259 953 1263 954
rect 1403 958 1407 959
rect 1403 953 1407 954
rect 1443 958 1447 959
rect 1443 953 1447 954
rect 1563 958 1567 959
rect 1563 953 1567 954
rect 1627 958 1631 959
rect 1627 953 1631 954
rect 1723 958 1727 959
rect 1723 953 1727 954
rect 1787 958 1791 959
rect 1787 953 1791 954
rect 1935 958 1939 959
rect 1935 953 1939 954
rect 112 893 114 953
rect 110 892 116 893
rect 228 892 230 953
rect 380 892 382 953
rect 540 892 542 953
rect 716 892 718 953
rect 892 892 894 953
rect 1076 892 1078 953
rect 1260 892 1262 953
rect 1444 892 1446 953
rect 1628 892 1630 953
rect 1788 892 1790 953
rect 1936 893 1938 953
rect 1976 935 1978 986
rect 3120 935 3122 987
rect 3272 935 3274 987
rect 3424 935 3426 987
rect 3798 986 3804 987
rect 3800 935 3802 986
rect 3840 943 3842 1003
rect 3860 943 3862 1004
rect 4044 943 4046 1004
rect 4252 943 4254 1004
rect 4484 943 4486 1004
rect 4732 943 4734 1004
rect 4996 943 4998 1004
rect 5268 943 5270 1004
rect 5516 943 5518 1004
rect 5662 1003 5668 1004
rect 5664 943 5666 1003
rect 3839 942 3843 943
rect 3839 937 3843 938
rect 3859 942 3863 943
rect 3859 937 3863 938
rect 3971 942 3975 943
rect 3971 937 3975 938
rect 4043 942 4047 943
rect 4043 937 4047 938
rect 4179 942 4183 943
rect 4179 937 4183 938
rect 4251 942 4255 943
rect 4251 937 4255 938
rect 4403 942 4407 943
rect 4403 937 4407 938
rect 4483 942 4487 943
rect 4483 937 4487 938
rect 4643 942 4647 943
rect 4643 937 4647 938
rect 4731 942 4735 943
rect 4731 937 4735 938
rect 4899 942 4903 943
rect 4899 937 4903 938
rect 4995 942 4999 943
rect 4995 937 4999 938
rect 5171 942 5175 943
rect 5171 937 5175 938
rect 5267 942 5271 943
rect 5267 937 5271 938
rect 5443 942 5447 943
rect 5443 937 5447 938
rect 5515 942 5519 943
rect 5515 937 5519 938
rect 5663 942 5667 943
rect 5663 937 5667 938
rect 1975 934 1979 935
rect 1975 929 1979 930
rect 2047 934 2051 935
rect 2047 929 2051 930
rect 2351 934 2355 935
rect 2351 929 2355 930
rect 2647 934 2651 935
rect 2647 929 2651 930
rect 2927 934 2931 935
rect 2927 929 2931 930
rect 3119 934 3123 935
rect 3119 929 3123 930
rect 3207 934 3211 935
rect 3207 929 3211 930
rect 3271 934 3275 935
rect 3271 929 3275 930
rect 3423 934 3427 935
rect 3423 929 3427 930
rect 3495 934 3499 935
rect 3495 929 3499 930
rect 3799 934 3803 935
rect 3799 929 3803 930
rect 1976 906 1978 929
rect 1974 905 1980 906
rect 2048 905 2050 929
rect 2352 905 2354 929
rect 2648 905 2650 929
rect 2928 905 2930 929
rect 3208 905 3210 929
rect 3496 905 3498 929
rect 3800 906 3802 929
rect 3798 905 3804 906
rect 1974 901 1975 905
rect 1979 901 1980 905
rect 1974 900 1980 901
rect 2046 904 2052 905
rect 2046 900 2047 904
rect 2051 900 2052 904
rect 2046 899 2052 900
rect 2350 904 2356 905
rect 2350 900 2351 904
rect 2355 900 2356 904
rect 2350 899 2356 900
rect 2646 904 2652 905
rect 2646 900 2647 904
rect 2651 900 2652 904
rect 2646 899 2652 900
rect 2926 904 2932 905
rect 2926 900 2927 904
rect 2931 900 2932 904
rect 2926 899 2932 900
rect 3206 904 3212 905
rect 3206 900 3207 904
rect 3211 900 3212 904
rect 3206 899 3212 900
rect 3494 904 3500 905
rect 3494 900 3495 904
rect 3499 900 3500 904
rect 3798 901 3799 905
rect 3803 901 3804 905
rect 3798 900 3804 901
rect 3494 899 3500 900
rect 1934 892 1940 893
rect 110 888 111 892
rect 115 888 116 892
rect 110 887 116 888
rect 226 891 232 892
rect 226 887 227 891
rect 231 887 232 891
rect 226 886 232 887
rect 378 891 384 892
rect 378 887 379 891
rect 383 887 384 891
rect 378 886 384 887
rect 538 891 544 892
rect 538 887 539 891
rect 543 887 544 891
rect 538 886 544 887
rect 714 891 720 892
rect 714 887 715 891
rect 719 887 720 891
rect 714 886 720 887
rect 890 891 896 892
rect 890 887 891 891
rect 895 887 896 891
rect 890 886 896 887
rect 1074 891 1080 892
rect 1074 887 1075 891
rect 1079 887 1080 891
rect 1074 886 1080 887
rect 1258 891 1264 892
rect 1258 887 1259 891
rect 1263 887 1264 891
rect 1258 886 1264 887
rect 1442 891 1448 892
rect 1442 887 1443 891
rect 1447 887 1448 891
rect 1442 886 1448 887
rect 1626 891 1632 892
rect 1626 887 1627 891
rect 1631 887 1632 891
rect 1626 886 1632 887
rect 1786 891 1792 892
rect 1786 887 1787 891
rect 1791 887 1792 891
rect 1934 888 1935 892
rect 1939 888 1940 892
rect 2018 889 2024 890
rect 1934 887 1940 888
rect 1974 888 1980 889
rect 1786 886 1792 887
rect 1974 884 1975 888
rect 1979 884 1980 888
rect 2018 885 2019 889
rect 2023 885 2024 889
rect 2018 884 2024 885
rect 2322 889 2328 890
rect 2322 885 2323 889
rect 2327 885 2328 889
rect 2322 884 2328 885
rect 2618 889 2624 890
rect 2618 885 2619 889
rect 2623 885 2624 889
rect 2618 884 2624 885
rect 2898 889 2904 890
rect 2898 885 2899 889
rect 2903 885 2904 889
rect 2898 884 2904 885
rect 3178 889 3184 890
rect 3178 885 3179 889
rect 3183 885 3184 889
rect 3178 884 3184 885
rect 3466 889 3472 890
rect 3466 885 3467 889
rect 3471 885 3472 889
rect 3466 884 3472 885
rect 3798 888 3804 889
rect 3798 884 3799 888
rect 3803 884 3804 888
rect 1974 883 1980 884
rect 254 876 260 877
rect 110 875 116 876
rect 110 871 111 875
rect 115 871 116 875
rect 254 872 255 876
rect 259 872 260 876
rect 254 871 260 872
rect 406 876 412 877
rect 406 872 407 876
rect 411 872 412 876
rect 406 871 412 872
rect 566 876 572 877
rect 566 872 567 876
rect 571 872 572 876
rect 566 871 572 872
rect 742 876 748 877
rect 742 872 743 876
rect 747 872 748 876
rect 742 871 748 872
rect 918 876 924 877
rect 918 872 919 876
rect 923 872 924 876
rect 918 871 924 872
rect 1102 876 1108 877
rect 1102 872 1103 876
rect 1107 872 1108 876
rect 1102 871 1108 872
rect 1286 876 1292 877
rect 1286 872 1287 876
rect 1291 872 1292 876
rect 1286 871 1292 872
rect 1470 876 1476 877
rect 1470 872 1471 876
rect 1475 872 1476 876
rect 1470 871 1476 872
rect 1654 876 1660 877
rect 1654 872 1655 876
rect 1659 872 1660 876
rect 1654 871 1660 872
rect 1814 876 1820 877
rect 1814 872 1815 876
rect 1819 872 1820 876
rect 1814 871 1820 872
rect 1934 875 1940 876
rect 1934 871 1935 875
rect 1939 871 1940 875
rect 110 870 116 871
rect 112 831 114 870
rect 256 831 258 871
rect 408 831 410 871
rect 568 831 570 871
rect 744 831 746 871
rect 920 831 922 871
rect 1104 831 1106 871
rect 1288 831 1290 871
rect 1472 831 1474 871
rect 1656 831 1658 871
rect 1816 831 1818 871
rect 1934 870 1940 871
rect 1936 831 1938 870
rect 111 830 115 831
rect 111 825 115 826
rect 255 830 259 831
rect 255 825 259 826
rect 375 830 379 831
rect 375 825 379 826
rect 407 830 411 831
rect 407 825 411 826
rect 567 830 571 831
rect 567 825 571 826
rect 655 830 659 831
rect 655 825 659 826
rect 743 830 747 831
rect 743 825 747 826
rect 919 830 923 831
rect 919 825 923 826
rect 943 830 947 831
rect 943 825 947 826
rect 1103 830 1107 831
rect 1103 825 1107 826
rect 1239 830 1243 831
rect 1239 825 1243 826
rect 1287 830 1291 831
rect 1287 825 1291 826
rect 1471 830 1475 831
rect 1471 825 1475 826
rect 1535 830 1539 831
rect 1535 825 1539 826
rect 1655 830 1659 831
rect 1655 825 1659 826
rect 1815 830 1819 831
rect 1815 825 1819 826
rect 1935 830 1939 831
rect 1935 825 1939 826
rect 112 802 114 825
rect 110 801 116 802
rect 376 801 378 825
rect 656 801 658 825
rect 944 801 946 825
rect 1240 801 1242 825
rect 1536 801 1538 825
rect 1816 801 1818 825
rect 1936 802 1938 825
rect 1976 823 1978 883
rect 2020 823 2022 884
rect 2324 823 2326 884
rect 2620 823 2622 884
rect 2900 823 2902 884
rect 3180 823 3182 884
rect 3468 823 3470 884
rect 3798 883 3804 884
rect 3800 823 3802 883
rect 3840 877 3842 937
rect 3838 876 3844 877
rect 3972 876 3974 937
rect 4180 876 4182 937
rect 4404 876 4406 937
rect 4644 876 4646 937
rect 4900 876 4902 937
rect 5172 876 5174 937
rect 5444 876 5446 937
rect 5664 877 5666 937
rect 5662 876 5668 877
rect 3838 872 3839 876
rect 3843 872 3844 876
rect 3838 871 3844 872
rect 3970 875 3976 876
rect 3970 871 3971 875
rect 3975 871 3976 875
rect 3970 870 3976 871
rect 4178 875 4184 876
rect 4178 871 4179 875
rect 4183 871 4184 875
rect 4178 870 4184 871
rect 4402 875 4408 876
rect 4402 871 4403 875
rect 4407 871 4408 875
rect 4402 870 4408 871
rect 4642 875 4648 876
rect 4642 871 4643 875
rect 4647 871 4648 875
rect 4642 870 4648 871
rect 4898 875 4904 876
rect 4898 871 4899 875
rect 4903 871 4904 875
rect 4898 870 4904 871
rect 5170 875 5176 876
rect 5170 871 5171 875
rect 5175 871 5176 875
rect 5170 870 5176 871
rect 5442 875 5448 876
rect 5442 871 5443 875
rect 5447 871 5448 875
rect 5662 872 5663 876
rect 5667 872 5668 876
rect 5662 871 5668 872
rect 5442 870 5448 871
rect 3998 860 4004 861
rect 3838 859 3844 860
rect 3838 855 3839 859
rect 3843 855 3844 859
rect 3998 856 3999 860
rect 4003 856 4004 860
rect 3998 855 4004 856
rect 4206 860 4212 861
rect 4206 856 4207 860
rect 4211 856 4212 860
rect 4206 855 4212 856
rect 4430 860 4436 861
rect 4430 856 4431 860
rect 4435 856 4436 860
rect 4430 855 4436 856
rect 4670 860 4676 861
rect 4670 856 4671 860
rect 4675 856 4676 860
rect 4670 855 4676 856
rect 4926 860 4932 861
rect 4926 856 4927 860
rect 4931 856 4932 860
rect 4926 855 4932 856
rect 5198 860 5204 861
rect 5198 856 5199 860
rect 5203 856 5204 860
rect 5198 855 5204 856
rect 5470 860 5476 861
rect 5470 856 5471 860
rect 5475 856 5476 860
rect 5470 855 5476 856
rect 5662 859 5668 860
rect 5662 855 5663 859
rect 5667 855 5668 859
rect 3838 854 3844 855
rect 3840 831 3842 854
rect 4000 831 4002 855
rect 4208 831 4210 855
rect 4432 831 4434 855
rect 4672 831 4674 855
rect 4928 831 4930 855
rect 5200 831 5202 855
rect 5472 831 5474 855
rect 5662 854 5668 855
rect 5664 831 5666 854
rect 3839 830 3843 831
rect 3839 825 3843 826
rect 3887 830 3891 831
rect 3887 825 3891 826
rect 3999 830 4003 831
rect 3999 825 4003 826
rect 4047 830 4051 831
rect 4047 825 4051 826
rect 4207 830 4211 831
rect 4207 825 4211 826
rect 4279 830 4283 831
rect 4279 825 4283 826
rect 4431 830 4435 831
rect 4431 825 4435 826
rect 4559 830 4563 831
rect 4559 825 4563 826
rect 4671 830 4675 831
rect 4671 825 4675 826
rect 4879 830 4883 831
rect 4879 825 4883 826
rect 4927 830 4931 831
rect 4927 825 4931 826
rect 5199 830 5203 831
rect 5199 825 5203 826
rect 5223 830 5227 831
rect 5223 825 5227 826
rect 5471 830 5475 831
rect 5471 825 5475 826
rect 5543 830 5547 831
rect 5543 825 5547 826
rect 5663 830 5667 831
rect 5663 825 5667 826
rect 1975 822 1979 823
rect 1975 817 1979 818
rect 1995 822 1999 823
rect 1995 817 1999 818
rect 2019 822 2023 823
rect 2019 817 2023 818
rect 2251 822 2255 823
rect 2251 817 2255 818
rect 2323 822 2327 823
rect 2323 817 2327 818
rect 2523 822 2527 823
rect 2523 817 2527 818
rect 2619 822 2623 823
rect 2619 817 2623 818
rect 2771 822 2775 823
rect 2771 817 2775 818
rect 2899 822 2903 823
rect 2899 817 2903 818
rect 3003 822 3007 823
rect 3003 817 3007 818
rect 3179 822 3183 823
rect 3179 817 3183 818
rect 3227 822 3231 823
rect 3227 817 3231 818
rect 3451 822 3455 823
rect 3451 817 3455 818
rect 3467 822 3471 823
rect 3467 817 3471 818
rect 3651 822 3655 823
rect 3651 817 3655 818
rect 3799 822 3803 823
rect 3799 817 3803 818
rect 1934 801 1940 802
rect 110 797 111 801
rect 115 797 116 801
rect 110 796 116 797
rect 374 800 380 801
rect 374 796 375 800
rect 379 796 380 800
rect 374 795 380 796
rect 654 800 660 801
rect 654 796 655 800
rect 659 796 660 800
rect 654 795 660 796
rect 942 800 948 801
rect 942 796 943 800
rect 947 796 948 800
rect 942 795 948 796
rect 1238 800 1244 801
rect 1238 796 1239 800
rect 1243 796 1244 800
rect 1238 795 1244 796
rect 1534 800 1540 801
rect 1534 796 1535 800
rect 1539 796 1540 800
rect 1534 795 1540 796
rect 1814 800 1820 801
rect 1814 796 1815 800
rect 1819 796 1820 800
rect 1934 797 1935 801
rect 1939 797 1940 801
rect 1934 796 1940 797
rect 1814 795 1820 796
rect 346 785 352 786
rect 110 784 116 785
rect 110 780 111 784
rect 115 780 116 784
rect 346 781 347 785
rect 351 781 352 785
rect 346 780 352 781
rect 626 785 632 786
rect 626 781 627 785
rect 631 781 632 785
rect 626 780 632 781
rect 914 785 920 786
rect 914 781 915 785
rect 919 781 920 785
rect 914 780 920 781
rect 1210 785 1216 786
rect 1210 781 1211 785
rect 1215 781 1216 785
rect 1210 780 1216 781
rect 1506 785 1512 786
rect 1506 781 1507 785
rect 1511 781 1512 785
rect 1506 780 1512 781
rect 1786 785 1792 786
rect 1786 781 1787 785
rect 1791 781 1792 785
rect 1786 780 1792 781
rect 1934 784 1940 785
rect 1934 780 1935 784
rect 1939 780 1940 784
rect 110 779 116 780
rect 112 719 114 779
rect 348 719 350 780
rect 628 719 630 780
rect 916 719 918 780
rect 1212 719 1214 780
rect 1508 719 1510 780
rect 1788 719 1790 780
rect 1934 779 1940 780
rect 1936 719 1938 779
rect 1976 757 1978 817
rect 1974 756 1980 757
rect 1996 756 1998 817
rect 2252 756 2254 817
rect 2524 756 2526 817
rect 2772 756 2774 817
rect 3004 756 3006 817
rect 3228 756 3230 817
rect 3452 756 3454 817
rect 3652 756 3654 817
rect 3800 757 3802 817
rect 3840 802 3842 825
rect 3838 801 3844 802
rect 3888 801 3890 825
rect 4048 801 4050 825
rect 4280 801 4282 825
rect 4560 801 4562 825
rect 4880 801 4882 825
rect 5224 801 5226 825
rect 5544 801 5546 825
rect 5664 802 5666 825
rect 5662 801 5668 802
rect 3838 797 3839 801
rect 3843 797 3844 801
rect 3838 796 3844 797
rect 3886 800 3892 801
rect 3886 796 3887 800
rect 3891 796 3892 800
rect 3886 795 3892 796
rect 4046 800 4052 801
rect 4046 796 4047 800
rect 4051 796 4052 800
rect 4046 795 4052 796
rect 4278 800 4284 801
rect 4278 796 4279 800
rect 4283 796 4284 800
rect 4278 795 4284 796
rect 4558 800 4564 801
rect 4558 796 4559 800
rect 4563 796 4564 800
rect 4558 795 4564 796
rect 4878 800 4884 801
rect 4878 796 4879 800
rect 4883 796 4884 800
rect 4878 795 4884 796
rect 5222 800 5228 801
rect 5222 796 5223 800
rect 5227 796 5228 800
rect 5222 795 5228 796
rect 5542 800 5548 801
rect 5542 796 5543 800
rect 5547 796 5548 800
rect 5662 797 5663 801
rect 5667 797 5668 801
rect 5662 796 5668 797
rect 5542 795 5548 796
rect 3858 785 3864 786
rect 3838 784 3844 785
rect 3838 780 3839 784
rect 3843 780 3844 784
rect 3858 781 3859 785
rect 3863 781 3864 785
rect 3858 780 3864 781
rect 4018 785 4024 786
rect 4018 781 4019 785
rect 4023 781 4024 785
rect 4018 780 4024 781
rect 4250 785 4256 786
rect 4250 781 4251 785
rect 4255 781 4256 785
rect 4250 780 4256 781
rect 4530 785 4536 786
rect 4530 781 4531 785
rect 4535 781 4536 785
rect 4530 780 4536 781
rect 4850 785 4856 786
rect 4850 781 4851 785
rect 4855 781 4856 785
rect 4850 780 4856 781
rect 5194 785 5200 786
rect 5194 781 5195 785
rect 5199 781 5200 785
rect 5194 780 5200 781
rect 5514 785 5520 786
rect 5514 781 5515 785
rect 5519 781 5520 785
rect 5514 780 5520 781
rect 5662 784 5668 785
rect 5662 780 5663 784
rect 5667 780 5668 784
rect 3838 779 3844 780
rect 3798 756 3804 757
rect 1974 752 1975 756
rect 1979 752 1980 756
rect 1974 751 1980 752
rect 1994 755 2000 756
rect 1994 751 1995 755
rect 1999 751 2000 755
rect 1994 750 2000 751
rect 2250 755 2256 756
rect 2250 751 2251 755
rect 2255 751 2256 755
rect 2250 750 2256 751
rect 2522 755 2528 756
rect 2522 751 2523 755
rect 2527 751 2528 755
rect 2522 750 2528 751
rect 2770 755 2776 756
rect 2770 751 2771 755
rect 2775 751 2776 755
rect 2770 750 2776 751
rect 3002 755 3008 756
rect 3002 751 3003 755
rect 3007 751 3008 755
rect 3002 750 3008 751
rect 3226 755 3232 756
rect 3226 751 3227 755
rect 3231 751 3232 755
rect 3226 750 3232 751
rect 3450 755 3456 756
rect 3450 751 3451 755
rect 3455 751 3456 755
rect 3450 750 3456 751
rect 3650 755 3656 756
rect 3650 751 3651 755
rect 3655 751 3656 755
rect 3798 752 3799 756
rect 3803 752 3804 756
rect 3798 751 3804 752
rect 3650 750 3656 751
rect 2022 740 2028 741
rect 1974 739 1980 740
rect 1974 735 1975 739
rect 1979 735 1980 739
rect 2022 736 2023 740
rect 2027 736 2028 740
rect 2022 735 2028 736
rect 2278 740 2284 741
rect 2278 736 2279 740
rect 2283 736 2284 740
rect 2278 735 2284 736
rect 2550 740 2556 741
rect 2550 736 2551 740
rect 2555 736 2556 740
rect 2550 735 2556 736
rect 2798 740 2804 741
rect 2798 736 2799 740
rect 2803 736 2804 740
rect 2798 735 2804 736
rect 3030 740 3036 741
rect 3030 736 3031 740
rect 3035 736 3036 740
rect 3030 735 3036 736
rect 3254 740 3260 741
rect 3254 736 3255 740
rect 3259 736 3260 740
rect 3254 735 3260 736
rect 3478 740 3484 741
rect 3478 736 3479 740
rect 3483 736 3484 740
rect 3478 735 3484 736
rect 3678 740 3684 741
rect 3678 736 3679 740
rect 3683 736 3684 740
rect 3678 735 3684 736
rect 3798 739 3804 740
rect 3798 735 3799 739
rect 3803 735 3804 739
rect 1974 734 1980 735
rect 111 718 115 719
rect 111 713 115 714
rect 131 718 135 719
rect 131 713 135 714
rect 307 718 311 719
rect 307 713 311 714
rect 347 718 351 719
rect 347 713 351 714
rect 499 718 503 719
rect 499 713 503 714
rect 627 718 631 719
rect 627 713 631 714
rect 683 718 687 719
rect 683 713 687 714
rect 859 718 863 719
rect 859 713 863 714
rect 915 718 919 719
rect 915 713 919 714
rect 1027 718 1031 719
rect 1027 713 1031 714
rect 1187 718 1191 719
rect 1187 713 1191 714
rect 1211 718 1215 719
rect 1211 713 1215 714
rect 1339 718 1343 719
rect 1339 713 1343 714
rect 1491 718 1495 719
rect 1491 713 1495 714
rect 1507 718 1511 719
rect 1507 713 1511 714
rect 1651 718 1655 719
rect 1651 713 1655 714
rect 1787 718 1791 719
rect 1787 713 1791 714
rect 1935 718 1939 719
rect 1935 713 1939 714
rect 112 653 114 713
rect 110 652 116 653
rect 132 652 134 713
rect 308 652 310 713
rect 500 652 502 713
rect 684 652 686 713
rect 860 652 862 713
rect 1028 652 1030 713
rect 1188 652 1190 713
rect 1340 652 1342 713
rect 1492 652 1494 713
rect 1652 652 1654 713
rect 1788 652 1790 713
rect 1936 653 1938 713
rect 1934 652 1940 653
rect 110 648 111 652
rect 115 648 116 652
rect 110 647 116 648
rect 130 651 136 652
rect 130 647 131 651
rect 135 647 136 651
rect 130 646 136 647
rect 306 651 312 652
rect 306 647 307 651
rect 311 647 312 651
rect 306 646 312 647
rect 498 651 504 652
rect 498 647 499 651
rect 503 647 504 651
rect 498 646 504 647
rect 682 651 688 652
rect 682 647 683 651
rect 687 647 688 651
rect 682 646 688 647
rect 858 651 864 652
rect 858 647 859 651
rect 863 647 864 651
rect 858 646 864 647
rect 1026 651 1032 652
rect 1026 647 1027 651
rect 1031 647 1032 651
rect 1026 646 1032 647
rect 1186 651 1192 652
rect 1186 647 1187 651
rect 1191 647 1192 651
rect 1186 646 1192 647
rect 1338 651 1344 652
rect 1338 647 1339 651
rect 1343 647 1344 651
rect 1338 646 1344 647
rect 1490 651 1496 652
rect 1490 647 1491 651
rect 1495 647 1496 651
rect 1490 646 1496 647
rect 1650 651 1656 652
rect 1650 647 1651 651
rect 1655 647 1656 651
rect 1650 646 1656 647
rect 1786 651 1792 652
rect 1786 647 1787 651
rect 1791 647 1792 651
rect 1934 648 1935 652
rect 1939 648 1940 652
rect 1934 647 1940 648
rect 1786 646 1792 647
rect 158 636 164 637
rect 110 635 116 636
rect 110 631 111 635
rect 115 631 116 635
rect 158 632 159 636
rect 163 632 164 636
rect 158 631 164 632
rect 334 636 340 637
rect 334 632 335 636
rect 339 632 340 636
rect 334 631 340 632
rect 526 636 532 637
rect 526 632 527 636
rect 531 632 532 636
rect 526 631 532 632
rect 710 636 716 637
rect 710 632 711 636
rect 715 632 716 636
rect 710 631 716 632
rect 886 636 892 637
rect 886 632 887 636
rect 891 632 892 636
rect 886 631 892 632
rect 1054 636 1060 637
rect 1054 632 1055 636
rect 1059 632 1060 636
rect 1054 631 1060 632
rect 1214 636 1220 637
rect 1214 632 1215 636
rect 1219 632 1220 636
rect 1214 631 1220 632
rect 1366 636 1372 637
rect 1366 632 1367 636
rect 1371 632 1372 636
rect 1366 631 1372 632
rect 1518 636 1524 637
rect 1518 632 1519 636
rect 1523 632 1524 636
rect 1518 631 1524 632
rect 1678 636 1684 637
rect 1678 632 1679 636
rect 1683 632 1684 636
rect 1678 631 1684 632
rect 1814 636 1820 637
rect 1814 632 1815 636
rect 1819 632 1820 636
rect 1814 631 1820 632
rect 1934 635 1940 636
rect 1934 631 1935 635
rect 1939 631 1940 635
rect 110 630 116 631
rect 112 607 114 630
rect 160 607 162 631
rect 336 607 338 631
rect 528 607 530 631
rect 712 607 714 631
rect 888 607 890 631
rect 1056 607 1058 631
rect 1216 607 1218 631
rect 1368 607 1370 631
rect 1520 607 1522 631
rect 1680 607 1682 631
rect 1816 607 1818 631
rect 1934 630 1940 631
rect 1936 607 1938 630
rect 111 606 115 607
rect 111 601 115 602
rect 159 606 163 607
rect 159 601 163 602
rect 335 606 339 607
rect 335 601 339 602
rect 375 606 379 607
rect 375 601 379 602
rect 527 606 531 607
rect 527 601 531 602
rect 599 606 603 607
rect 599 601 603 602
rect 711 606 715 607
rect 711 601 715 602
rect 807 606 811 607
rect 807 601 811 602
rect 887 606 891 607
rect 887 601 891 602
rect 999 606 1003 607
rect 999 601 1003 602
rect 1055 606 1059 607
rect 1055 601 1059 602
rect 1175 606 1179 607
rect 1175 601 1179 602
rect 1215 606 1219 607
rect 1215 601 1219 602
rect 1343 606 1347 607
rect 1343 601 1347 602
rect 1367 606 1371 607
rect 1367 601 1371 602
rect 1511 606 1515 607
rect 1511 601 1515 602
rect 1519 606 1523 607
rect 1519 601 1523 602
rect 1671 606 1675 607
rect 1671 601 1675 602
rect 1679 606 1683 607
rect 1679 601 1683 602
rect 1815 606 1819 607
rect 1815 601 1819 602
rect 1935 606 1939 607
rect 1935 601 1939 602
rect 112 578 114 601
rect 110 577 116 578
rect 160 577 162 601
rect 376 577 378 601
rect 600 577 602 601
rect 808 577 810 601
rect 1000 577 1002 601
rect 1176 577 1178 601
rect 1344 577 1346 601
rect 1512 577 1514 601
rect 1672 577 1674 601
rect 1816 577 1818 601
rect 1936 578 1938 601
rect 1976 579 1978 734
rect 2024 579 2026 735
rect 2280 579 2282 735
rect 2552 579 2554 735
rect 2800 579 2802 735
rect 3032 579 3034 735
rect 3256 579 3258 735
rect 3480 579 3482 735
rect 3680 579 3682 735
rect 3798 734 3804 735
rect 3800 579 3802 734
rect 3840 711 3842 779
rect 3860 711 3862 780
rect 4020 711 4022 780
rect 4252 711 4254 780
rect 4532 711 4534 780
rect 4852 711 4854 780
rect 5196 711 5198 780
rect 5516 711 5518 780
rect 5662 779 5668 780
rect 5664 711 5666 779
rect 3839 710 3843 711
rect 3839 705 3843 706
rect 3859 710 3863 711
rect 3859 705 3863 706
rect 3995 710 3999 711
rect 3995 705 3999 706
rect 4019 710 4023 711
rect 4019 705 4023 706
rect 4131 710 4135 711
rect 4131 705 4135 706
rect 4251 710 4255 711
rect 4251 705 4255 706
rect 4267 710 4271 711
rect 4267 705 4271 706
rect 4403 710 4407 711
rect 4403 705 4407 706
rect 4531 710 4535 711
rect 4531 705 4535 706
rect 4571 710 4575 711
rect 4571 705 4575 706
rect 4771 710 4775 711
rect 4771 705 4775 706
rect 4851 710 4855 711
rect 4851 705 4855 706
rect 4995 710 4999 711
rect 4995 705 4999 706
rect 5195 710 5199 711
rect 5195 705 5199 706
rect 5227 710 5231 711
rect 5227 705 5231 706
rect 5459 710 5463 711
rect 5459 705 5463 706
rect 5515 710 5519 711
rect 5515 705 5519 706
rect 5663 710 5667 711
rect 5663 705 5667 706
rect 3840 645 3842 705
rect 3838 644 3844 645
rect 3860 644 3862 705
rect 3996 644 3998 705
rect 4132 644 4134 705
rect 4268 644 4270 705
rect 4404 644 4406 705
rect 4572 644 4574 705
rect 4772 644 4774 705
rect 4996 644 4998 705
rect 5228 644 5230 705
rect 5460 644 5462 705
rect 5664 645 5666 705
rect 5662 644 5668 645
rect 3838 640 3839 644
rect 3843 640 3844 644
rect 3838 639 3844 640
rect 3858 643 3864 644
rect 3858 639 3859 643
rect 3863 639 3864 643
rect 3858 638 3864 639
rect 3994 643 4000 644
rect 3994 639 3995 643
rect 3999 639 4000 643
rect 3994 638 4000 639
rect 4130 643 4136 644
rect 4130 639 4131 643
rect 4135 639 4136 643
rect 4130 638 4136 639
rect 4266 643 4272 644
rect 4266 639 4267 643
rect 4271 639 4272 643
rect 4266 638 4272 639
rect 4402 643 4408 644
rect 4402 639 4403 643
rect 4407 639 4408 643
rect 4402 638 4408 639
rect 4570 643 4576 644
rect 4570 639 4571 643
rect 4575 639 4576 643
rect 4570 638 4576 639
rect 4770 643 4776 644
rect 4770 639 4771 643
rect 4775 639 4776 643
rect 4770 638 4776 639
rect 4994 643 5000 644
rect 4994 639 4995 643
rect 4999 639 5000 643
rect 4994 638 5000 639
rect 5226 643 5232 644
rect 5226 639 5227 643
rect 5231 639 5232 643
rect 5226 638 5232 639
rect 5458 643 5464 644
rect 5458 639 5459 643
rect 5463 639 5464 643
rect 5662 640 5663 644
rect 5667 640 5668 644
rect 5662 639 5668 640
rect 5458 638 5464 639
rect 3886 628 3892 629
rect 3838 627 3844 628
rect 3838 623 3839 627
rect 3843 623 3844 627
rect 3886 624 3887 628
rect 3891 624 3892 628
rect 3886 623 3892 624
rect 4022 628 4028 629
rect 4022 624 4023 628
rect 4027 624 4028 628
rect 4022 623 4028 624
rect 4158 628 4164 629
rect 4158 624 4159 628
rect 4163 624 4164 628
rect 4158 623 4164 624
rect 4294 628 4300 629
rect 4294 624 4295 628
rect 4299 624 4300 628
rect 4294 623 4300 624
rect 4430 628 4436 629
rect 4430 624 4431 628
rect 4435 624 4436 628
rect 4430 623 4436 624
rect 4598 628 4604 629
rect 4598 624 4599 628
rect 4603 624 4604 628
rect 4598 623 4604 624
rect 4798 628 4804 629
rect 4798 624 4799 628
rect 4803 624 4804 628
rect 4798 623 4804 624
rect 5022 628 5028 629
rect 5022 624 5023 628
rect 5027 624 5028 628
rect 5022 623 5028 624
rect 5254 628 5260 629
rect 5254 624 5255 628
rect 5259 624 5260 628
rect 5254 623 5260 624
rect 5486 628 5492 629
rect 5486 624 5487 628
rect 5491 624 5492 628
rect 5486 623 5492 624
rect 5662 627 5668 628
rect 5662 623 5663 627
rect 5667 623 5668 627
rect 3838 622 3844 623
rect 3840 599 3842 622
rect 3888 599 3890 623
rect 4024 599 4026 623
rect 4160 599 4162 623
rect 4296 599 4298 623
rect 4432 599 4434 623
rect 4600 599 4602 623
rect 4800 599 4802 623
rect 5024 599 5026 623
rect 5256 599 5258 623
rect 5488 599 5490 623
rect 5662 622 5668 623
rect 5664 599 5666 622
rect 3839 598 3843 599
rect 3839 593 3843 594
rect 3887 598 3891 599
rect 3887 593 3891 594
rect 4023 598 4027 599
rect 4023 593 4027 594
rect 4159 598 4163 599
rect 4159 593 4163 594
rect 4295 598 4299 599
rect 4295 593 4299 594
rect 4431 598 4435 599
rect 4431 593 4435 594
rect 4479 598 4483 599
rect 4479 593 4483 594
rect 4599 598 4603 599
rect 4599 593 4603 594
rect 4695 598 4699 599
rect 4695 593 4699 594
rect 4799 598 4803 599
rect 4799 593 4803 594
rect 4935 598 4939 599
rect 4935 593 4939 594
rect 5023 598 5027 599
rect 5023 593 5027 594
rect 5191 598 5195 599
rect 5191 593 5195 594
rect 5255 598 5259 599
rect 5255 593 5259 594
rect 5447 598 5451 599
rect 5447 593 5451 594
rect 5487 598 5491 599
rect 5487 593 5491 594
rect 5663 598 5667 599
rect 5663 593 5667 594
rect 1975 578 1979 579
rect 1934 577 1940 578
rect 110 573 111 577
rect 115 573 116 577
rect 110 572 116 573
rect 158 576 164 577
rect 158 572 159 576
rect 163 572 164 576
rect 158 571 164 572
rect 374 576 380 577
rect 374 572 375 576
rect 379 572 380 576
rect 374 571 380 572
rect 598 576 604 577
rect 598 572 599 576
rect 603 572 604 576
rect 598 571 604 572
rect 806 576 812 577
rect 806 572 807 576
rect 811 572 812 576
rect 806 571 812 572
rect 998 576 1004 577
rect 998 572 999 576
rect 1003 572 1004 576
rect 998 571 1004 572
rect 1174 576 1180 577
rect 1174 572 1175 576
rect 1179 572 1180 576
rect 1174 571 1180 572
rect 1342 576 1348 577
rect 1342 572 1343 576
rect 1347 572 1348 576
rect 1342 571 1348 572
rect 1510 576 1516 577
rect 1510 572 1511 576
rect 1515 572 1516 576
rect 1510 571 1516 572
rect 1670 576 1676 577
rect 1670 572 1671 576
rect 1675 572 1676 576
rect 1670 571 1676 572
rect 1814 576 1820 577
rect 1814 572 1815 576
rect 1819 572 1820 576
rect 1934 573 1935 577
rect 1939 573 1940 577
rect 1975 573 1979 574
rect 2023 578 2027 579
rect 2023 573 2027 574
rect 2279 578 2283 579
rect 2279 573 2283 574
rect 2551 578 2555 579
rect 2551 573 2555 574
rect 2799 578 2803 579
rect 2799 573 2803 574
rect 3031 578 3035 579
rect 3031 573 3035 574
rect 3255 578 3259 579
rect 3255 573 3259 574
rect 3311 578 3315 579
rect 3311 573 3315 574
rect 3447 578 3451 579
rect 3447 573 3451 574
rect 3479 578 3483 579
rect 3479 573 3483 574
rect 3583 578 3587 579
rect 3583 573 3587 574
rect 3679 578 3683 579
rect 3679 573 3683 574
rect 3799 578 3803 579
rect 3799 573 3803 574
rect 1934 572 1940 573
rect 1814 571 1820 572
rect 130 561 136 562
rect 110 560 116 561
rect 110 556 111 560
rect 115 556 116 560
rect 130 557 131 561
rect 135 557 136 561
rect 130 556 136 557
rect 346 561 352 562
rect 346 557 347 561
rect 351 557 352 561
rect 346 556 352 557
rect 570 561 576 562
rect 570 557 571 561
rect 575 557 576 561
rect 570 556 576 557
rect 778 561 784 562
rect 778 557 779 561
rect 783 557 784 561
rect 778 556 784 557
rect 970 561 976 562
rect 970 557 971 561
rect 975 557 976 561
rect 970 556 976 557
rect 1146 561 1152 562
rect 1146 557 1147 561
rect 1151 557 1152 561
rect 1146 556 1152 557
rect 1314 561 1320 562
rect 1314 557 1315 561
rect 1319 557 1320 561
rect 1314 556 1320 557
rect 1482 561 1488 562
rect 1482 557 1483 561
rect 1487 557 1488 561
rect 1482 556 1488 557
rect 1642 561 1648 562
rect 1642 557 1643 561
rect 1647 557 1648 561
rect 1642 556 1648 557
rect 1786 561 1792 562
rect 1786 557 1787 561
rect 1791 557 1792 561
rect 1786 556 1792 557
rect 1934 560 1940 561
rect 1934 556 1935 560
rect 1939 556 1940 560
rect 110 555 116 556
rect 112 495 114 555
rect 132 495 134 556
rect 348 495 350 556
rect 572 495 574 556
rect 780 495 782 556
rect 972 495 974 556
rect 1148 495 1150 556
rect 1316 495 1318 556
rect 1484 495 1486 556
rect 1644 495 1646 556
rect 1788 495 1790 556
rect 1934 555 1940 556
rect 1936 495 1938 555
rect 1976 550 1978 573
rect 1974 549 1980 550
rect 3312 549 3314 573
rect 3448 549 3450 573
rect 3584 549 3586 573
rect 3800 550 3802 573
rect 3840 570 3842 593
rect 3838 569 3844 570
rect 3888 569 3890 593
rect 4024 569 4026 593
rect 4160 569 4162 593
rect 4296 569 4298 593
rect 4480 569 4482 593
rect 4696 569 4698 593
rect 4936 569 4938 593
rect 5192 569 5194 593
rect 5448 569 5450 593
rect 5664 570 5666 593
rect 5662 569 5668 570
rect 3838 565 3839 569
rect 3843 565 3844 569
rect 3838 564 3844 565
rect 3886 568 3892 569
rect 3886 564 3887 568
rect 3891 564 3892 568
rect 3886 563 3892 564
rect 4022 568 4028 569
rect 4022 564 4023 568
rect 4027 564 4028 568
rect 4022 563 4028 564
rect 4158 568 4164 569
rect 4158 564 4159 568
rect 4163 564 4164 568
rect 4158 563 4164 564
rect 4294 568 4300 569
rect 4294 564 4295 568
rect 4299 564 4300 568
rect 4294 563 4300 564
rect 4478 568 4484 569
rect 4478 564 4479 568
rect 4483 564 4484 568
rect 4478 563 4484 564
rect 4694 568 4700 569
rect 4694 564 4695 568
rect 4699 564 4700 568
rect 4694 563 4700 564
rect 4934 568 4940 569
rect 4934 564 4935 568
rect 4939 564 4940 568
rect 4934 563 4940 564
rect 5190 568 5196 569
rect 5190 564 5191 568
rect 5195 564 5196 568
rect 5190 563 5196 564
rect 5446 568 5452 569
rect 5446 564 5447 568
rect 5451 564 5452 568
rect 5662 565 5663 569
rect 5667 565 5668 569
rect 5662 564 5668 565
rect 5446 563 5452 564
rect 3858 553 3864 554
rect 3838 552 3844 553
rect 3798 549 3804 550
rect 1974 545 1975 549
rect 1979 545 1980 549
rect 1974 544 1980 545
rect 3310 548 3316 549
rect 3310 544 3311 548
rect 3315 544 3316 548
rect 3310 543 3316 544
rect 3446 548 3452 549
rect 3446 544 3447 548
rect 3451 544 3452 548
rect 3446 543 3452 544
rect 3582 548 3588 549
rect 3582 544 3583 548
rect 3587 544 3588 548
rect 3798 545 3799 549
rect 3803 545 3804 549
rect 3838 548 3839 552
rect 3843 548 3844 552
rect 3858 549 3859 553
rect 3863 549 3864 553
rect 3858 548 3864 549
rect 3994 553 4000 554
rect 3994 549 3995 553
rect 3999 549 4000 553
rect 3994 548 4000 549
rect 4130 553 4136 554
rect 4130 549 4131 553
rect 4135 549 4136 553
rect 4130 548 4136 549
rect 4266 553 4272 554
rect 4266 549 4267 553
rect 4271 549 4272 553
rect 4266 548 4272 549
rect 4450 553 4456 554
rect 4450 549 4451 553
rect 4455 549 4456 553
rect 4450 548 4456 549
rect 4666 553 4672 554
rect 4666 549 4667 553
rect 4671 549 4672 553
rect 4666 548 4672 549
rect 4906 553 4912 554
rect 4906 549 4907 553
rect 4911 549 4912 553
rect 4906 548 4912 549
rect 5162 553 5168 554
rect 5162 549 5163 553
rect 5167 549 5168 553
rect 5162 548 5168 549
rect 5418 553 5424 554
rect 5418 549 5419 553
rect 5423 549 5424 553
rect 5418 548 5424 549
rect 5662 552 5668 553
rect 5662 548 5663 552
rect 5667 548 5668 552
rect 3838 547 3844 548
rect 3798 544 3804 545
rect 3582 543 3588 544
rect 3282 533 3288 534
rect 1974 532 1980 533
rect 1974 528 1975 532
rect 1979 528 1980 532
rect 3282 529 3283 533
rect 3287 529 3288 533
rect 3282 528 3288 529
rect 3418 533 3424 534
rect 3418 529 3419 533
rect 3423 529 3424 533
rect 3418 528 3424 529
rect 3554 533 3560 534
rect 3554 529 3555 533
rect 3559 529 3560 533
rect 3554 528 3560 529
rect 3798 532 3804 533
rect 3798 528 3799 532
rect 3803 528 3804 532
rect 1974 527 1980 528
rect 111 494 115 495
rect 111 489 115 490
rect 131 494 135 495
rect 131 489 135 490
rect 347 494 351 495
rect 347 489 351 490
rect 427 494 431 495
rect 427 489 431 490
rect 571 494 575 495
rect 571 489 575 490
rect 763 494 767 495
rect 763 489 767 490
rect 779 494 783 495
rect 779 489 783 490
rect 971 494 975 495
rect 971 489 975 490
rect 1107 494 1111 495
rect 1107 489 1111 490
rect 1147 494 1151 495
rect 1147 489 1151 490
rect 1315 494 1319 495
rect 1315 489 1319 490
rect 1459 494 1463 495
rect 1459 489 1463 490
rect 1483 494 1487 495
rect 1483 489 1487 490
rect 1643 494 1647 495
rect 1643 489 1647 490
rect 1787 494 1791 495
rect 1787 489 1791 490
rect 1935 494 1939 495
rect 1935 489 1939 490
rect 112 429 114 489
rect 110 428 116 429
rect 132 428 134 489
rect 428 428 430 489
rect 764 428 766 489
rect 1108 428 1110 489
rect 1460 428 1462 489
rect 1788 428 1790 489
rect 1936 429 1938 489
rect 1976 467 1978 527
rect 3284 467 3286 528
rect 3420 467 3422 528
rect 3556 467 3558 528
rect 3798 527 3804 528
rect 3800 467 3802 527
rect 3840 475 3842 547
rect 3860 475 3862 548
rect 3996 475 3998 548
rect 4132 475 4134 548
rect 4268 475 4270 548
rect 4452 475 4454 548
rect 4668 475 4670 548
rect 4908 475 4910 548
rect 5164 475 5166 548
rect 5420 475 5422 548
rect 5662 547 5668 548
rect 5664 475 5666 547
rect 3839 474 3843 475
rect 3839 469 3843 470
rect 3859 474 3863 475
rect 3859 469 3863 470
rect 3995 474 3999 475
rect 3995 469 3999 470
rect 4131 474 4135 475
rect 4131 469 4135 470
rect 4267 474 4271 475
rect 4267 469 4271 470
rect 4451 474 4455 475
rect 4451 469 4455 470
rect 4651 474 4655 475
rect 4651 469 4655 470
rect 4667 474 4671 475
rect 4667 469 4671 470
rect 4859 474 4863 475
rect 4859 469 4863 470
rect 4907 474 4911 475
rect 4907 469 4911 470
rect 5067 474 5071 475
rect 5067 469 5071 470
rect 5163 474 5167 475
rect 5163 469 5167 470
rect 5283 474 5287 475
rect 5283 469 5287 470
rect 5419 474 5423 475
rect 5419 469 5423 470
rect 5507 474 5511 475
rect 5507 469 5511 470
rect 5663 474 5667 475
rect 5663 469 5667 470
rect 1975 466 1979 467
rect 1975 461 1979 462
rect 1995 466 1999 467
rect 1995 461 1999 462
rect 2155 466 2159 467
rect 2155 461 2159 462
rect 2347 466 2351 467
rect 2347 461 2351 462
rect 2539 466 2543 467
rect 2539 461 2543 462
rect 2731 466 2735 467
rect 2731 461 2735 462
rect 2923 466 2927 467
rect 2923 461 2927 462
rect 3115 466 3119 467
rect 3115 461 3119 462
rect 3283 466 3287 467
rect 3283 461 3287 462
rect 3299 466 3303 467
rect 3299 461 3303 462
rect 3419 466 3423 467
rect 3419 461 3423 462
rect 3483 466 3487 467
rect 3483 461 3487 462
rect 3555 466 3559 467
rect 3555 461 3559 462
rect 3651 466 3655 467
rect 3651 461 3655 462
rect 3799 466 3803 467
rect 3799 461 3803 462
rect 1934 428 1940 429
rect 110 424 111 428
rect 115 424 116 428
rect 110 423 116 424
rect 130 427 136 428
rect 130 423 131 427
rect 135 423 136 427
rect 130 422 136 423
rect 426 427 432 428
rect 426 423 427 427
rect 431 423 432 427
rect 426 422 432 423
rect 762 427 768 428
rect 762 423 763 427
rect 767 423 768 427
rect 762 422 768 423
rect 1106 427 1112 428
rect 1106 423 1107 427
rect 1111 423 1112 427
rect 1106 422 1112 423
rect 1458 427 1464 428
rect 1458 423 1459 427
rect 1463 423 1464 427
rect 1458 422 1464 423
rect 1786 427 1792 428
rect 1786 423 1787 427
rect 1791 423 1792 427
rect 1934 424 1935 428
rect 1939 424 1940 428
rect 1934 423 1940 424
rect 1786 422 1792 423
rect 158 412 164 413
rect 110 411 116 412
rect 110 407 111 411
rect 115 407 116 411
rect 158 408 159 412
rect 163 408 164 412
rect 158 407 164 408
rect 454 412 460 413
rect 454 408 455 412
rect 459 408 460 412
rect 454 407 460 408
rect 790 412 796 413
rect 790 408 791 412
rect 795 408 796 412
rect 790 407 796 408
rect 1134 412 1140 413
rect 1134 408 1135 412
rect 1139 408 1140 412
rect 1134 407 1140 408
rect 1486 412 1492 413
rect 1486 408 1487 412
rect 1491 408 1492 412
rect 1486 407 1492 408
rect 1814 412 1820 413
rect 1814 408 1815 412
rect 1819 408 1820 412
rect 1814 407 1820 408
rect 1934 411 1940 412
rect 1934 407 1935 411
rect 1939 407 1940 411
rect 110 406 116 407
rect 112 367 114 406
rect 160 367 162 407
rect 456 367 458 407
rect 792 367 794 407
rect 1136 367 1138 407
rect 1488 367 1490 407
rect 1816 367 1818 407
rect 1934 406 1940 407
rect 1936 367 1938 406
rect 1976 401 1978 461
rect 1974 400 1980 401
rect 1996 400 1998 461
rect 2156 400 2158 461
rect 2348 400 2350 461
rect 2540 400 2542 461
rect 2732 400 2734 461
rect 2924 400 2926 461
rect 3116 400 3118 461
rect 3300 400 3302 461
rect 3484 400 3486 461
rect 3652 400 3654 461
rect 3800 401 3802 461
rect 3840 409 3842 469
rect 3838 408 3844 409
rect 4452 408 4454 469
rect 4652 408 4654 469
rect 4860 408 4862 469
rect 5068 408 5070 469
rect 5284 408 5286 469
rect 5508 408 5510 469
rect 5664 409 5666 469
rect 5662 408 5668 409
rect 3838 404 3839 408
rect 3843 404 3844 408
rect 3838 403 3844 404
rect 4450 407 4456 408
rect 4450 403 4451 407
rect 4455 403 4456 407
rect 4450 402 4456 403
rect 4650 407 4656 408
rect 4650 403 4651 407
rect 4655 403 4656 407
rect 4650 402 4656 403
rect 4858 407 4864 408
rect 4858 403 4859 407
rect 4863 403 4864 407
rect 4858 402 4864 403
rect 5066 407 5072 408
rect 5066 403 5067 407
rect 5071 403 5072 407
rect 5066 402 5072 403
rect 5282 407 5288 408
rect 5282 403 5283 407
rect 5287 403 5288 407
rect 5282 402 5288 403
rect 5506 407 5512 408
rect 5506 403 5507 407
rect 5511 403 5512 407
rect 5662 404 5663 408
rect 5667 404 5668 408
rect 5662 403 5668 404
rect 5506 402 5512 403
rect 3798 400 3804 401
rect 1974 396 1975 400
rect 1979 396 1980 400
rect 1974 395 1980 396
rect 1994 399 2000 400
rect 1994 395 1995 399
rect 1999 395 2000 399
rect 1994 394 2000 395
rect 2154 399 2160 400
rect 2154 395 2155 399
rect 2159 395 2160 399
rect 2154 394 2160 395
rect 2346 399 2352 400
rect 2346 395 2347 399
rect 2351 395 2352 399
rect 2346 394 2352 395
rect 2538 399 2544 400
rect 2538 395 2539 399
rect 2543 395 2544 399
rect 2538 394 2544 395
rect 2730 399 2736 400
rect 2730 395 2731 399
rect 2735 395 2736 399
rect 2730 394 2736 395
rect 2922 399 2928 400
rect 2922 395 2923 399
rect 2927 395 2928 399
rect 2922 394 2928 395
rect 3114 399 3120 400
rect 3114 395 3115 399
rect 3119 395 3120 399
rect 3114 394 3120 395
rect 3298 399 3304 400
rect 3298 395 3299 399
rect 3303 395 3304 399
rect 3298 394 3304 395
rect 3482 399 3488 400
rect 3482 395 3483 399
rect 3487 395 3488 399
rect 3482 394 3488 395
rect 3650 399 3656 400
rect 3650 395 3651 399
rect 3655 395 3656 399
rect 3798 396 3799 400
rect 3803 396 3804 400
rect 3798 395 3804 396
rect 3650 394 3656 395
rect 4478 392 4484 393
rect 3838 391 3844 392
rect 3838 387 3839 391
rect 3843 387 3844 391
rect 4478 388 4479 392
rect 4483 388 4484 392
rect 4478 387 4484 388
rect 4678 392 4684 393
rect 4678 388 4679 392
rect 4683 388 4684 392
rect 4678 387 4684 388
rect 4886 392 4892 393
rect 4886 388 4887 392
rect 4891 388 4892 392
rect 4886 387 4892 388
rect 5094 392 5100 393
rect 5094 388 5095 392
rect 5099 388 5100 392
rect 5094 387 5100 388
rect 5310 392 5316 393
rect 5310 388 5311 392
rect 5315 388 5316 392
rect 5310 387 5316 388
rect 5534 392 5540 393
rect 5534 388 5535 392
rect 5539 388 5540 392
rect 5534 387 5540 388
rect 5662 391 5668 392
rect 5662 387 5663 391
rect 5667 387 5668 391
rect 3838 386 3844 387
rect 2022 384 2028 385
rect 1974 383 1980 384
rect 1974 379 1975 383
rect 1979 379 1980 383
rect 2022 380 2023 384
rect 2027 380 2028 384
rect 2022 379 2028 380
rect 2182 384 2188 385
rect 2182 380 2183 384
rect 2187 380 2188 384
rect 2182 379 2188 380
rect 2374 384 2380 385
rect 2374 380 2375 384
rect 2379 380 2380 384
rect 2374 379 2380 380
rect 2566 384 2572 385
rect 2566 380 2567 384
rect 2571 380 2572 384
rect 2566 379 2572 380
rect 2758 384 2764 385
rect 2758 380 2759 384
rect 2763 380 2764 384
rect 2758 379 2764 380
rect 2950 384 2956 385
rect 2950 380 2951 384
rect 2955 380 2956 384
rect 2950 379 2956 380
rect 3142 384 3148 385
rect 3142 380 3143 384
rect 3147 380 3148 384
rect 3142 379 3148 380
rect 3326 384 3332 385
rect 3326 380 3327 384
rect 3331 380 3332 384
rect 3326 379 3332 380
rect 3510 384 3516 385
rect 3510 380 3511 384
rect 3515 380 3516 384
rect 3510 379 3516 380
rect 3678 384 3684 385
rect 3678 380 3679 384
rect 3683 380 3684 384
rect 3678 379 3684 380
rect 3798 383 3804 384
rect 3798 379 3799 383
rect 3803 379 3804 383
rect 1974 378 1980 379
rect 111 366 115 367
rect 111 361 115 362
rect 159 366 163 367
rect 159 361 163 362
rect 239 366 243 367
rect 239 361 243 362
rect 391 366 395 367
rect 391 361 395 362
rect 455 366 459 367
rect 455 361 459 362
rect 551 366 555 367
rect 551 361 555 362
rect 711 366 715 367
rect 711 361 715 362
rect 791 366 795 367
rect 791 361 795 362
rect 871 366 875 367
rect 871 361 875 362
rect 1031 366 1035 367
rect 1031 361 1035 362
rect 1135 366 1139 367
rect 1135 361 1139 362
rect 1487 366 1491 367
rect 1487 361 1491 362
rect 1815 366 1819 367
rect 1815 361 1819 362
rect 1935 366 1939 367
rect 1935 361 1939 362
rect 112 338 114 361
rect 110 337 116 338
rect 240 337 242 361
rect 392 337 394 361
rect 552 337 554 361
rect 712 337 714 361
rect 872 337 874 361
rect 1032 337 1034 361
rect 1936 338 1938 361
rect 1934 337 1940 338
rect 110 333 111 337
rect 115 333 116 337
rect 110 332 116 333
rect 238 336 244 337
rect 238 332 239 336
rect 243 332 244 336
rect 238 331 244 332
rect 390 336 396 337
rect 390 332 391 336
rect 395 332 396 336
rect 390 331 396 332
rect 550 336 556 337
rect 550 332 551 336
rect 555 332 556 336
rect 550 331 556 332
rect 710 336 716 337
rect 710 332 711 336
rect 715 332 716 336
rect 710 331 716 332
rect 870 336 876 337
rect 870 332 871 336
rect 875 332 876 336
rect 870 331 876 332
rect 1030 336 1036 337
rect 1030 332 1031 336
rect 1035 332 1036 336
rect 1934 333 1935 337
rect 1939 333 1940 337
rect 1934 332 1940 333
rect 1030 331 1036 332
rect 1976 331 1978 378
rect 2024 331 2026 379
rect 2184 331 2186 379
rect 2376 331 2378 379
rect 2568 331 2570 379
rect 2760 331 2762 379
rect 2952 331 2954 379
rect 3144 331 3146 379
rect 3328 331 3330 379
rect 3512 331 3514 379
rect 3680 331 3682 379
rect 3798 378 3804 379
rect 3800 331 3802 378
rect 3840 359 3842 386
rect 4480 359 4482 387
rect 4680 359 4682 387
rect 4888 359 4890 387
rect 5096 359 5098 387
rect 5312 359 5314 387
rect 5536 359 5538 387
rect 5662 386 5668 387
rect 5664 359 5666 386
rect 3839 358 3843 359
rect 3839 353 3843 354
rect 4479 358 4483 359
rect 4479 353 4483 354
rect 4679 358 4683 359
rect 4679 353 4683 354
rect 4751 358 4755 359
rect 4751 353 4755 354
rect 4887 358 4891 359
rect 4887 353 4891 354
rect 4911 358 4915 359
rect 4911 353 4915 354
rect 5071 358 5075 359
rect 5071 353 5075 354
rect 5095 358 5099 359
rect 5095 353 5099 354
rect 5231 358 5235 359
rect 5231 353 5235 354
rect 5311 358 5315 359
rect 5311 353 5315 354
rect 5399 358 5403 359
rect 5399 353 5403 354
rect 5535 358 5539 359
rect 5535 353 5539 354
rect 5543 358 5547 359
rect 5543 353 5547 354
rect 5663 358 5667 359
rect 5663 353 5667 354
rect 1975 330 1979 331
rect 1975 325 1979 326
rect 2023 330 2027 331
rect 2023 325 2027 326
rect 2047 330 2051 331
rect 2047 325 2051 326
rect 2183 330 2187 331
rect 2183 325 2187 326
rect 2319 330 2323 331
rect 2319 325 2323 326
rect 2375 330 2379 331
rect 2375 325 2379 326
rect 2455 330 2459 331
rect 2455 325 2459 326
rect 2567 330 2571 331
rect 2567 325 2571 326
rect 2591 330 2595 331
rect 2591 325 2595 326
rect 2727 330 2731 331
rect 2727 325 2731 326
rect 2759 330 2763 331
rect 2759 325 2763 326
rect 2863 330 2867 331
rect 2863 325 2867 326
rect 2951 330 2955 331
rect 2951 325 2955 326
rect 2999 330 3003 331
rect 2999 325 3003 326
rect 3135 330 3139 331
rect 3135 325 3139 326
rect 3143 330 3147 331
rect 3143 325 3147 326
rect 3271 330 3275 331
rect 3271 325 3275 326
rect 3327 330 3331 331
rect 3327 325 3331 326
rect 3407 330 3411 331
rect 3407 325 3411 326
rect 3511 330 3515 331
rect 3511 325 3515 326
rect 3543 330 3547 331
rect 3543 325 3547 326
rect 3679 330 3683 331
rect 3679 325 3683 326
rect 3799 330 3803 331
rect 3840 330 3842 353
rect 3799 325 3803 326
rect 3838 329 3844 330
rect 4752 329 4754 353
rect 4912 329 4914 353
rect 5072 329 5074 353
rect 5232 329 5234 353
rect 5400 329 5402 353
rect 5544 329 5546 353
rect 5664 330 5666 353
rect 5662 329 5668 330
rect 3838 325 3839 329
rect 3843 325 3844 329
rect 210 321 216 322
rect 110 320 116 321
rect 110 316 111 320
rect 115 316 116 320
rect 210 317 211 321
rect 215 317 216 321
rect 210 316 216 317
rect 362 321 368 322
rect 362 317 363 321
rect 367 317 368 321
rect 362 316 368 317
rect 522 321 528 322
rect 522 317 523 321
rect 527 317 528 321
rect 522 316 528 317
rect 682 321 688 322
rect 682 317 683 321
rect 687 317 688 321
rect 682 316 688 317
rect 842 321 848 322
rect 842 317 843 321
rect 847 317 848 321
rect 842 316 848 317
rect 1002 321 1008 322
rect 1002 317 1003 321
rect 1007 317 1008 321
rect 1002 316 1008 317
rect 1934 320 1940 321
rect 1934 316 1935 320
rect 1939 316 1940 320
rect 110 315 116 316
rect 112 223 114 315
rect 212 223 214 316
rect 364 223 366 316
rect 524 223 526 316
rect 684 223 686 316
rect 844 223 846 316
rect 1004 223 1006 316
rect 1934 315 1940 316
rect 1936 223 1938 315
rect 1976 302 1978 325
rect 1974 301 1980 302
rect 2048 301 2050 325
rect 2184 301 2186 325
rect 2320 301 2322 325
rect 2456 301 2458 325
rect 2592 301 2594 325
rect 2728 301 2730 325
rect 2864 301 2866 325
rect 3000 301 3002 325
rect 3136 301 3138 325
rect 3272 301 3274 325
rect 3408 301 3410 325
rect 3544 301 3546 325
rect 3680 301 3682 325
rect 3800 302 3802 325
rect 3838 324 3844 325
rect 4750 328 4756 329
rect 4750 324 4751 328
rect 4755 324 4756 328
rect 4750 323 4756 324
rect 4910 328 4916 329
rect 4910 324 4911 328
rect 4915 324 4916 328
rect 4910 323 4916 324
rect 5070 328 5076 329
rect 5070 324 5071 328
rect 5075 324 5076 328
rect 5070 323 5076 324
rect 5230 328 5236 329
rect 5230 324 5231 328
rect 5235 324 5236 328
rect 5230 323 5236 324
rect 5398 328 5404 329
rect 5398 324 5399 328
rect 5403 324 5404 328
rect 5398 323 5404 324
rect 5542 328 5548 329
rect 5542 324 5543 328
rect 5547 324 5548 328
rect 5662 325 5663 329
rect 5667 325 5668 329
rect 5662 324 5668 325
rect 5542 323 5548 324
rect 4722 313 4728 314
rect 3838 312 3844 313
rect 3838 308 3839 312
rect 3843 308 3844 312
rect 4722 309 4723 313
rect 4727 309 4728 313
rect 4722 308 4728 309
rect 4882 313 4888 314
rect 4882 309 4883 313
rect 4887 309 4888 313
rect 4882 308 4888 309
rect 5042 313 5048 314
rect 5042 309 5043 313
rect 5047 309 5048 313
rect 5042 308 5048 309
rect 5202 313 5208 314
rect 5202 309 5203 313
rect 5207 309 5208 313
rect 5202 308 5208 309
rect 5370 313 5376 314
rect 5370 309 5371 313
rect 5375 309 5376 313
rect 5370 308 5376 309
rect 5514 313 5520 314
rect 5514 309 5515 313
rect 5519 309 5520 313
rect 5514 308 5520 309
rect 5662 312 5668 313
rect 5662 308 5663 312
rect 5667 308 5668 312
rect 3838 307 3844 308
rect 3798 301 3804 302
rect 1974 297 1975 301
rect 1979 297 1980 301
rect 1974 296 1980 297
rect 2046 300 2052 301
rect 2046 296 2047 300
rect 2051 296 2052 300
rect 2046 295 2052 296
rect 2182 300 2188 301
rect 2182 296 2183 300
rect 2187 296 2188 300
rect 2182 295 2188 296
rect 2318 300 2324 301
rect 2318 296 2319 300
rect 2323 296 2324 300
rect 2318 295 2324 296
rect 2454 300 2460 301
rect 2454 296 2455 300
rect 2459 296 2460 300
rect 2454 295 2460 296
rect 2590 300 2596 301
rect 2590 296 2591 300
rect 2595 296 2596 300
rect 2590 295 2596 296
rect 2726 300 2732 301
rect 2726 296 2727 300
rect 2731 296 2732 300
rect 2726 295 2732 296
rect 2862 300 2868 301
rect 2862 296 2863 300
rect 2867 296 2868 300
rect 2862 295 2868 296
rect 2998 300 3004 301
rect 2998 296 2999 300
rect 3003 296 3004 300
rect 2998 295 3004 296
rect 3134 300 3140 301
rect 3134 296 3135 300
rect 3139 296 3140 300
rect 3134 295 3140 296
rect 3270 300 3276 301
rect 3270 296 3271 300
rect 3275 296 3276 300
rect 3270 295 3276 296
rect 3406 300 3412 301
rect 3406 296 3407 300
rect 3411 296 3412 300
rect 3406 295 3412 296
rect 3542 300 3548 301
rect 3542 296 3543 300
rect 3547 296 3548 300
rect 3542 295 3548 296
rect 3678 300 3684 301
rect 3678 296 3679 300
rect 3683 296 3684 300
rect 3798 297 3799 301
rect 3803 297 3804 301
rect 3798 296 3804 297
rect 3678 295 3684 296
rect 2018 285 2024 286
rect 1974 284 1980 285
rect 1974 280 1975 284
rect 1979 280 1980 284
rect 2018 281 2019 285
rect 2023 281 2024 285
rect 2018 280 2024 281
rect 2154 285 2160 286
rect 2154 281 2155 285
rect 2159 281 2160 285
rect 2154 280 2160 281
rect 2290 285 2296 286
rect 2290 281 2291 285
rect 2295 281 2296 285
rect 2290 280 2296 281
rect 2426 285 2432 286
rect 2426 281 2427 285
rect 2431 281 2432 285
rect 2426 280 2432 281
rect 2562 285 2568 286
rect 2562 281 2563 285
rect 2567 281 2568 285
rect 2562 280 2568 281
rect 2698 285 2704 286
rect 2698 281 2699 285
rect 2703 281 2704 285
rect 2698 280 2704 281
rect 2834 285 2840 286
rect 2834 281 2835 285
rect 2839 281 2840 285
rect 2834 280 2840 281
rect 2970 285 2976 286
rect 2970 281 2971 285
rect 2975 281 2976 285
rect 2970 280 2976 281
rect 3106 285 3112 286
rect 3106 281 3107 285
rect 3111 281 3112 285
rect 3106 280 3112 281
rect 3242 285 3248 286
rect 3242 281 3243 285
rect 3247 281 3248 285
rect 3242 280 3248 281
rect 3378 285 3384 286
rect 3378 281 3379 285
rect 3383 281 3384 285
rect 3378 280 3384 281
rect 3514 285 3520 286
rect 3514 281 3515 285
rect 3519 281 3520 285
rect 3514 280 3520 281
rect 3650 285 3656 286
rect 3650 281 3651 285
rect 3655 281 3656 285
rect 3650 280 3656 281
rect 3798 284 3804 285
rect 3798 280 3799 284
rect 3803 280 3804 284
rect 1974 279 1980 280
rect 111 222 115 223
rect 111 217 115 218
rect 147 222 151 223
rect 147 217 151 218
rect 211 222 215 223
rect 211 217 215 218
rect 283 222 287 223
rect 283 217 287 218
rect 363 222 367 223
rect 363 217 367 218
rect 419 222 423 223
rect 419 217 423 218
rect 523 222 527 223
rect 523 217 527 218
rect 555 222 559 223
rect 555 217 559 218
rect 683 222 687 223
rect 683 217 687 218
rect 691 222 695 223
rect 691 217 695 218
rect 827 222 831 223
rect 827 217 831 218
rect 843 222 847 223
rect 843 217 847 218
rect 963 222 967 223
rect 963 217 967 218
rect 1003 222 1007 223
rect 1003 217 1007 218
rect 1099 222 1103 223
rect 1099 217 1103 218
rect 1935 222 1939 223
rect 1935 217 1939 218
rect 112 157 114 217
rect 110 156 116 157
rect 148 156 150 217
rect 284 156 286 217
rect 420 156 422 217
rect 556 156 558 217
rect 692 156 694 217
rect 828 156 830 217
rect 964 156 966 217
rect 1100 156 1102 217
rect 1936 157 1938 217
rect 1976 203 1978 279
rect 2020 203 2022 280
rect 2156 203 2158 280
rect 2292 203 2294 280
rect 2428 203 2430 280
rect 2564 203 2566 280
rect 2700 203 2702 280
rect 2836 203 2838 280
rect 2972 203 2974 280
rect 3108 203 3110 280
rect 3244 203 3246 280
rect 3380 203 3382 280
rect 3516 203 3518 280
rect 3652 203 3654 280
rect 3798 279 3804 280
rect 3800 203 3802 279
rect 3840 207 3842 307
rect 4724 207 4726 308
rect 4884 207 4886 308
rect 5044 207 5046 308
rect 5204 207 5206 308
rect 5372 207 5374 308
rect 5516 207 5518 308
rect 5662 307 5668 308
rect 5664 207 5666 307
rect 3839 206 3843 207
rect 1975 202 1979 203
rect 1975 197 1979 198
rect 1995 202 1999 203
rect 1995 197 1999 198
rect 2019 202 2023 203
rect 2019 197 2023 198
rect 2131 202 2135 203
rect 2131 197 2135 198
rect 2155 202 2159 203
rect 2155 197 2159 198
rect 2267 202 2271 203
rect 2267 197 2271 198
rect 2291 202 2295 203
rect 2291 197 2295 198
rect 2403 202 2407 203
rect 2403 197 2407 198
rect 2427 202 2431 203
rect 2427 197 2431 198
rect 2539 202 2543 203
rect 2539 197 2543 198
rect 2563 202 2567 203
rect 2563 197 2567 198
rect 2675 202 2679 203
rect 2675 197 2679 198
rect 2699 202 2703 203
rect 2699 197 2703 198
rect 2811 202 2815 203
rect 2811 197 2815 198
rect 2835 202 2839 203
rect 2835 197 2839 198
rect 2947 202 2951 203
rect 2947 197 2951 198
rect 2971 202 2975 203
rect 2971 197 2975 198
rect 3083 202 3087 203
rect 3083 197 3087 198
rect 3107 202 3111 203
rect 3107 197 3111 198
rect 3219 202 3223 203
rect 3219 197 3223 198
rect 3243 202 3247 203
rect 3243 197 3247 198
rect 3355 202 3359 203
rect 3355 197 3359 198
rect 3379 202 3383 203
rect 3379 197 3383 198
rect 3491 202 3495 203
rect 3491 197 3495 198
rect 3515 202 3519 203
rect 3515 197 3519 198
rect 3627 202 3631 203
rect 3627 197 3631 198
rect 3651 202 3655 203
rect 3651 197 3655 198
rect 3799 202 3803 203
rect 3839 201 3843 202
rect 4291 206 4295 207
rect 4291 201 4295 202
rect 4427 206 4431 207
rect 4427 201 4431 202
rect 4563 206 4567 207
rect 4563 201 4567 202
rect 4699 206 4703 207
rect 4699 201 4703 202
rect 4723 206 4727 207
rect 4723 201 4727 202
rect 4835 206 4839 207
rect 4835 201 4839 202
rect 4883 206 4887 207
rect 4883 201 4887 202
rect 4971 206 4975 207
rect 4971 201 4975 202
rect 5043 206 5047 207
rect 5043 201 5047 202
rect 5107 206 5111 207
rect 5107 201 5111 202
rect 5203 206 5207 207
rect 5203 201 5207 202
rect 5243 206 5247 207
rect 5243 201 5247 202
rect 5371 206 5375 207
rect 5371 201 5375 202
rect 5379 206 5383 207
rect 5379 201 5383 202
rect 5515 206 5519 207
rect 5515 201 5519 202
rect 5663 206 5667 207
rect 5663 201 5667 202
rect 3799 197 3803 198
rect 1934 156 1940 157
rect 110 152 111 156
rect 115 152 116 156
rect 110 151 116 152
rect 146 155 152 156
rect 146 151 147 155
rect 151 151 152 155
rect 146 150 152 151
rect 282 155 288 156
rect 282 151 283 155
rect 287 151 288 155
rect 282 150 288 151
rect 418 155 424 156
rect 418 151 419 155
rect 423 151 424 155
rect 418 150 424 151
rect 554 155 560 156
rect 554 151 555 155
rect 559 151 560 155
rect 554 150 560 151
rect 690 155 696 156
rect 690 151 691 155
rect 695 151 696 155
rect 690 150 696 151
rect 826 155 832 156
rect 826 151 827 155
rect 831 151 832 155
rect 826 150 832 151
rect 962 155 968 156
rect 962 151 963 155
rect 967 151 968 155
rect 962 150 968 151
rect 1098 155 1104 156
rect 1098 151 1099 155
rect 1103 151 1104 155
rect 1934 152 1935 156
rect 1939 152 1940 156
rect 1934 151 1940 152
rect 1098 150 1104 151
rect 174 140 180 141
rect 110 139 116 140
rect 110 135 111 139
rect 115 135 116 139
rect 174 136 175 140
rect 179 136 180 140
rect 174 135 180 136
rect 310 140 316 141
rect 310 136 311 140
rect 315 136 316 140
rect 310 135 316 136
rect 446 140 452 141
rect 446 136 447 140
rect 451 136 452 140
rect 446 135 452 136
rect 582 140 588 141
rect 582 136 583 140
rect 587 136 588 140
rect 582 135 588 136
rect 718 140 724 141
rect 718 136 719 140
rect 723 136 724 140
rect 718 135 724 136
rect 854 140 860 141
rect 854 136 855 140
rect 859 136 860 140
rect 854 135 860 136
rect 990 140 996 141
rect 990 136 991 140
rect 995 136 996 140
rect 990 135 996 136
rect 1126 140 1132 141
rect 1126 136 1127 140
rect 1131 136 1132 140
rect 1126 135 1132 136
rect 1934 139 1940 140
rect 1934 135 1935 139
rect 1939 135 1940 139
rect 1976 137 1978 197
rect 110 134 116 135
rect 112 111 114 134
rect 176 111 178 135
rect 312 111 314 135
rect 448 111 450 135
rect 584 111 586 135
rect 720 111 722 135
rect 856 111 858 135
rect 992 111 994 135
rect 1128 111 1130 135
rect 1934 134 1940 135
rect 1974 136 1980 137
rect 1996 136 1998 197
rect 2132 136 2134 197
rect 2268 136 2270 197
rect 2404 136 2406 197
rect 2540 136 2542 197
rect 2676 136 2678 197
rect 2812 136 2814 197
rect 2948 136 2950 197
rect 3084 136 3086 197
rect 3220 136 3222 197
rect 3356 136 3358 197
rect 3492 136 3494 197
rect 3628 136 3630 197
rect 3800 137 3802 197
rect 3840 141 3842 201
rect 3838 140 3844 141
rect 4292 140 4294 201
rect 4428 140 4430 201
rect 4564 140 4566 201
rect 4700 140 4702 201
rect 4836 140 4838 201
rect 4972 140 4974 201
rect 5108 140 5110 201
rect 5244 140 5246 201
rect 5380 140 5382 201
rect 5516 140 5518 201
rect 5664 141 5666 201
rect 5662 140 5668 141
rect 3798 136 3804 137
rect 1936 111 1938 134
rect 1974 132 1975 136
rect 1979 132 1980 136
rect 1974 131 1980 132
rect 1994 135 2000 136
rect 1994 131 1995 135
rect 1999 131 2000 135
rect 1994 130 2000 131
rect 2130 135 2136 136
rect 2130 131 2131 135
rect 2135 131 2136 135
rect 2130 130 2136 131
rect 2266 135 2272 136
rect 2266 131 2267 135
rect 2271 131 2272 135
rect 2266 130 2272 131
rect 2402 135 2408 136
rect 2402 131 2403 135
rect 2407 131 2408 135
rect 2402 130 2408 131
rect 2538 135 2544 136
rect 2538 131 2539 135
rect 2543 131 2544 135
rect 2538 130 2544 131
rect 2674 135 2680 136
rect 2674 131 2675 135
rect 2679 131 2680 135
rect 2674 130 2680 131
rect 2810 135 2816 136
rect 2810 131 2811 135
rect 2815 131 2816 135
rect 2810 130 2816 131
rect 2946 135 2952 136
rect 2946 131 2947 135
rect 2951 131 2952 135
rect 2946 130 2952 131
rect 3082 135 3088 136
rect 3082 131 3083 135
rect 3087 131 3088 135
rect 3082 130 3088 131
rect 3218 135 3224 136
rect 3218 131 3219 135
rect 3223 131 3224 135
rect 3218 130 3224 131
rect 3354 135 3360 136
rect 3354 131 3355 135
rect 3359 131 3360 135
rect 3354 130 3360 131
rect 3490 135 3496 136
rect 3490 131 3491 135
rect 3495 131 3496 135
rect 3490 130 3496 131
rect 3626 135 3632 136
rect 3626 131 3627 135
rect 3631 131 3632 135
rect 3798 132 3799 136
rect 3803 132 3804 136
rect 3838 136 3839 140
rect 3843 136 3844 140
rect 3838 135 3844 136
rect 4290 139 4296 140
rect 4290 135 4291 139
rect 4295 135 4296 139
rect 4290 134 4296 135
rect 4426 139 4432 140
rect 4426 135 4427 139
rect 4431 135 4432 139
rect 4426 134 4432 135
rect 4562 139 4568 140
rect 4562 135 4563 139
rect 4567 135 4568 139
rect 4562 134 4568 135
rect 4698 139 4704 140
rect 4698 135 4699 139
rect 4703 135 4704 139
rect 4698 134 4704 135
rect 4834 139 4840 140
rect 4834 135 4835 139
rect 4839 135 4840 139
rect 4834 134 4840 135
rect 4970 139 4976 140
rect 4970 135 4971 139
rect 4975 135 4976 139
rect 4970 134 4976 135
rect 5106 139 5112 140
rect 5106 135 5107 139
rect 5111 135 5112 139
rect 5106 134 5112 135
rect 5242 139 5248 140
rect 5242 135 5243 139
rect 5247 135 5248 139
rect 5242 134 5248 135
rect 5378 139 5384 140
rect 5378 135 5379 139
rect 5383 135 5384 139
rect 5378 134 5384 135
rect 5514 139 5520 140
rect 5514 135 5515 139
rect 5519 135 5520 139
rect 5662 136 5663 140
rect 5667 136 5668 140
rect 5662 135 5668 136
rect 5514 134 5520 135
rect 3798 131 3804 132
rect 3626 130 3632 131
rect 4318 124 4324 125
rect 3838 123 3844 124
rect 2022 120 2028 121
rect 1974 119 1980 120
rect 1974 115 1975 119
rect 1979 115 1980 119
rect 2022 116 2023 120
rect 2027 116 2028 120
rect 2022 115 2028 116
rect 2158 120 2164 121
rect 2158 116 2159 120
rect 2163 116 2164 120
rect 2158 115 2164 116
rect 2294 120 2300 121
rect 2294 116 2295 120
rect 2299 116 2300 120
rect 2294 115 2300 116
rect 2430 120 2436 121
rect 2430 116 2431 120
rect 2435 116 2436 120
rect 2430 115 2436 116
rect 2566 120 2572 121
rect 2566 116 2567 120
rect 2571 116 2572 120
rect 2566 115 2572 116
rect 2702 120 2708 121
rect 2702 116 2703 120
rect 2707 116 2708 120
rect 2702 115 2708 116
rect 2838 120 2844 121
rect 2838 116 2839 120
rect 2843 116 2844 120
rect 2838 115 2844 116
rect 2974 120 2980 121
rect 2974 116 2975 120
rect 2979 116 2980 120
rect 2974 115 2980 116
rect 3110 120 3116 121
rect 3110 116 3111 120
rect 3115 116 3116 120
rect 3110 115 3116 116
rect 3246 120 3252 121
rect 3246 116 3247 120
rect 3251 116 3252 120
rect 3246 115 3252 116
rect 3382 120 3388 121
rect 3382 116 3383 120
rect 3387 116 3388 120
rect 3382 115 3388 116
rect 3518 120 3524 121
rect 3518 116 3519 120
rect 3523 116 3524 120
rect 3518 115 3524 116
rect 3654 120 3660 121
rect 3654 116 3655 120
rect 3659 116 3660 120
rect 3654 115 3660 116
rect 3798 119 3804 120
rect 3798 115 3799 119
rect 3803 115 3804 119
rect 3838 119 3839 123
rect 3843 119 3844 123
rect 4318 120 4319 124
rect 4323 120 4324 124
rect 4318 119 4324 120
rect 4454 124 4460 125
rect 4454 120 4455 124
rect 4459 120 4460 124
rect 4454 119 4460 120
rect 4590 124 4596 125
rect 4590 120 4591 124
rect 4595 120 4596 124
rect 4590 119 4596 120
rect 4726 124 4732 125
rect 4726 120 4727 124
rect 4731 120 4732 124
rect 4726 119 4732 120
rect 4862 124 4868 125
rect 4862 120 4863 124
rect 4867 120 4868 124
rect 4862 119 4868 120
rect 4998 124 5004 125
rect 4998 120 4999 124
rect 5003 120 5004 124
rect 4998 119 5004 120
rect 5134 124 5140 125
rect 5134 120 5135 124
rect 5139 120 5140 124
rect 5134 119 5140 120
rect 5270 124 5276 125
rect 5270 120 5271 124
rect 5275 120 5276 124
rect 5270 119 5276 120
rect 5406 124 5412 125
rect 5406 120 5407 124
rect 5411 120 5412 124
rect 5406 119 5412 120
rect 5542 124 5548 125
rect 5542 120 5543 124
rect 5547 120 5548 124
rect 5542 119 5548 120
rect 5662 123 5668 124
rect 5662 119 5663 123
rect 5667 119 5668 123
rect 3838 118 3844 119
rect 1974 114 1980 115
rect 111 110 115 111
rect 111 105 115 106
rect 175 110 179 111
rect 175 105 179 106
rect 311 110 315 111
rect 311 105 315 106
rect 447 110 451 111
rect 447 105 451 106
rect 583 110 587 111
rect 583 105 587 106
rect 719 110 723 111
rect 719 105 723 106
rect 855 110 859 111
rect 855 105 859 106
rect 991 110 995 111
rect 991 105 995 106
rect 1127 110 1131 111
rect 1127 105 1131 106
rect 1935 110 1939 111
rect 1935 105 1939 106
rect 1976 91 1978 114
rect 2024 91 2026 115
rect 2160 91 2162 115
rect 2296 91 2298 115
rect 2432 91 2434 115
rect 2568 91 2570 115
rect 2704 91 2706 115
rect 2840 91 2842 115
rect 2976 91 2978 115
rect 3112 91 3114 115
rect 3248 91 3250 115
rect 3384 91 3386 115
rect 3520 91 3522 115
rect 3656 91 3658 115
rect 3798 114 3804 115
rect 3800 91 3802 114
rect 3840 95 3842 118
rect 4320 95 4322 119
rect 4456 95 4458 119
rect 4592 95 4594 119
rect 4728 95 4730 119
rect 4864 95 4866 119
rect 5000 95 5002 119
rect 5136 95 5138 119
rect 5272 95 5274 119
rect 5408 95 5410 119
rect 5544 95 5546 119
rect 5662 118 5668 119
rect 5664 95 5666 118
rect 3839 94 3843 95
rect 1975 90 1979 91
rect 1975 85 1979 86
rect 2023 90 2027 91
rect 2023 85 2027 86
rect 2159 90 2163 91
rect 2159 85 2163 86
rect 2295 90 2299 91
rect 2295 85 2299 86
rect 2431 90 2435 91
rect 2431 85 2435 86
rect 2567 90 2571 91
rect 2567 85 2571 86
rect 2703 90 2707 91
rect 2703 85 2707 86
rect 2839 90 2843 91
rect 2839 85 2843 86
rect 2975 90 2979 91
rect 2975 85 2979 86
rect 3111 90 3115 91
rect 3111 85 3115 86
rect 3247 90 3251 91
rect 3247 85 3251 86
rect 3383 90 3387 91
rect 3383 85 3387 86
rect 3519 90 3523 91
rect 3519 85 3523 86
rect 3655 90 3659 91
rect 3655 85 3659 86
rect 3799 90 3803 91
rect 3839 89 3843 90
rect 4319 94 4323 95
rect 4319 89 4323 90
rect 4455 94 4459 95
rect 4455 89 4459 90
rect 4591 94 4595 95
rect 4591 89 4595 90
rect 4727 94 4731 95
rect 4727 89 4731 90
rect 4863 94 4867 95
rect 4863 89 4867 90
rect 4999 94 5003 95
rect 4999 89 5003 90
rect 5135 94 5139 95
rect 5135 89 5139 90
rect 5271 94 5275 95
rect 5271 89 5275 90
rect 5407 94 5411 95
rect 5407 89 5411 90
rect 5543 94 5547 95
rect 5543 89 5547 90
rect 5663 94 5667 95
rect 5663 89 5667 90
rect 3799 85 3803 86
<< m4c >>
rect 111 5754 115 5758
rect 131 5754 135 5758
rect 267 5754 271 5758
rect 403 5754 407 5758
rect 1935 5754 1939 5758
rect 1975 5686 1979 5690
rect 1995 5686 1999 5690
rect 2171 5686 2175 5690
rect 2371 5686 2375 5690
rect 2563 5686 2567 5690
rect 2747 5686 2751 5690
rect 2931 5686 2935 5690
rect 3107 5686 3111 5690
rect 3275 5686 3279 5690
rect 3443 5686 3447 5690
rect 3619 5686 3623 5690
rect 3799 5686 3803 5690
rect 3839 5690 3843 5694
rect 4467 5690 4471 5694
rect 4603 5690 4607 5694
rect 4739 5690 4743 5694
rect 4875 5690 4879 5694
rect 5663 5690 5667 5694
rect 111 5642 115 5646
rect 159 5642 163 5646
rect 295 5642 299 5646
rect 343 5642 347 5646
rect 431 5642 435 5646
rect 535 5642 539 5646
rect 735 5642 739 5646
rect 943 5642 947 5646
rect 1159 5642 1163 5646
rect 1383 5642 1387 5646
rect 1607 5642 1611 5646
rect 1815 5642 1819 5646
rect 1935 5642 1939 5646
rect 1975 5574 1979 5578
rect 2023 5574 2027 5578
rect 2199 5574 2203 5578
rect 2375 5574 2379 5578
rect 2399 5574 2403 5578
rect 2591 5574 2595 5578
rect 2607 5574 2611 5578
rect 2775 5574 2779 5578
rect 2831 5574 2835 5578
rect 2959 5574 2963 5578
rect 3047 5574 3051 5578
rect 3135 5574 3139 5578
rect 3263 5574 3267 5578
rect 3303 5574 3307 5578
rect 3471 5574 3475 5578
rect 3479 5574 3483 5578
rect 3647 5574 3651 5578
rect 3679 5574 3683 5578
rect 3799 5574 3803 5578
rect 3839 5578 3843 5582
rect 4431 5578 4435 5582
rect 4495 5578 4499 5582
rect 4567 5578 4571 5582
rect 4631 5578 4635 5582
rect 4703 5578 4707 5582
rect 4767 5578 4771 5582
rect 4839 5578 4843 5582
rect 4903 5578 4907 5582
rect 4975 5578 4979 5582
rect 5111 5578 5115 5582
rect 5663 5578 5667 5582
rect 111 5530 115 5534
rect 315 5530 319 5534
rect 507 5530 511 5534
rect 707 5530 711 5534
rect 875 5530 879 5534
rect 915 5530 919 5534
rect 1011 5530 1015 5534
rect 1131 5530 1135 5534
rect 1147 5530 1151 5534
rect 1291 5530 1295 5534
rect 1355 5530 1359 5534
rect 1435 5530 1439 5534
rect 1579 5530 1583 5534
rect 1723 5530 1727 5534
rect 1787 5530 1791 5534
rect 1935 5530 1939 5534
rect 3839 5466 3843 5470
rect 4403 5466 4407 5470
rect 4427 5466 4431 5470
rect 4539 5466 4543 5470
rect 4587 5466 4591 5470
rect 4675 5466 4679 5470
rect 4747 5466 4751 5470
rect 4811 5466 4815 5470
rect 4907 5466 4911 5470
rect 4947 5466 4951 5470
rect 5075 5466 5079 5470
rect 5083 5466 5087 5470
rect 5663 5466 5667 5470
rect 1975 5458 1979 5462
rect 2347 5458 2351 5462
rect 2451 5458 2455 5462
rect 2579 5458 2583 5462
rect 2699 5458 2703 5462
rect 2803 5458 2807 5462
rect 2947 5458 2951 5462
rect 3019 5458 3023 5462
rect 3187 5458 3191 5462
rect 3235 5458 3239 5462
rect 3427 5458 3431 5462
rect 3451 5458 3455 5462
rect 3651 5458 3655 5462
rect 3799 5458 3803 5462
rect 111 5418 115 5422
rect 719 5418 723 5422
rect 855 5418 859 5422
rect 903 5418 907 5422
rect 991 5418 995 5422
rect 1039 5418 1043 5422
rect 1127 5418 1131 5422
rect 1175 5418 1179 5422
rect 1263 5418 1267 5422
rect 1319 5418 1323 5422
rect 1399 5418 1403 5422
rect 1463 5418 1467 5422
rect 1535 5418 1539 5422
rect 1607 5418 1611 5422
rect 1671 5418 1675 5422
rect 1751 5418 1755 5422
rect 1807 5418 1811 5422
rect 1935 5418 1939 5422
rect 1975 5346 1979 5350
rect 2319 5346 2323 5350
rect 2479 5346 2483 5350
rect 2519 5346 2523 5350
rect 2719 5346 2723 5350
rect 2727 5346 2731 5350
rect 2919 5346 2923 5350
rect 2975 5346 2979 5350
rect 3119 5346 3123 5350
rect 3215 5346 3219 5350
rect 3327 5346 3331 5350
rect 3455 5346 3459 5350
rect 3535 5346 3539 5350
rect 3679 5346 3683 5350
rect 3799 5346 3803 5350
rect 3839 5346 3843 5350
rect 4431 5346 4435 5350
rect 4455 5346 4459 5350
rect 4615 5346 4619 5350
rect 4775 5346 4779 5350
rect 4799 5346 4803 5350
rect 4935 5346 4939 5350
rect 4983 5346 4987 5350
rect 5103 5346 5107 5350
rect 5175 5346 5179 5350
rect 5663 5346 5667 5350
rect 111 5306 115 5310
rect 691 5306 695 5310
rect 723 5306 727 5310
rect 827 5306 831 5310
rect 875 5306 879 5310
rect 963 5306 967 5310
rect 1027 5306 1031 5310
rect 1099 5306 1103 5310
rect 1187 5306 1191 5310
rect 1235 5306 1239 5310
rect 1355 5306 1359 5310
rect 1371 5306 1375 5310
rect 1507 5306 1511 5310
rect 1523 5306 1527 5310
rect 1643 5306 1647 5310
rect 1779 5306 1783 5310
rect 1935 5306 1939 5310
rect 1975 5230 1979 5234
rect 2275 5230 2279 5234
rect 2291 5230 2295 5234
rect 2475 5230 2479 5234
rect 2491 5230 2495 5234
rect 2683 5230 2687 5234
rect 2691 5230 2695 5234
rect 2891 5230 2895 5234
rect 3091 5230 3095 5234
rect 3099 5230 3103 5234
rect 3299 5230 3303 5234
rect 3307 5230 3311 5234
rect 3507 5230 3511 5234
rect 3799 5230 3803 5234
rect 111 5194 115 5198
rect 447 5194 451 5198
rect 623 5194 627 5198
rect 751 5194 755 5198
rect 807 5194 811 5198
rect 903 5194 907 5198
rect 999 5194 1003 5198
rect 1055 5194 1059 5198
rect 1199 5194 1203 5198
rect 1215 5194 1219 5198
rect 1383 5194 1387 5198
rect 1399 5194 1403 5198
rect 1551 5194 1555 5198
rect 1607 5194 1611 5198
rect 1815 5194 1819 5198
rect 1935 5194 1939 5198
rect 3839 5218 3843 5222
rect 4403 5218 4407 5222
rect 4435 5218 4439 5222
rect 4587 5218 4591 5222
rect 4595 5218 4599 5222
rect 4755 5218 4759 5222
rect 4771 5218 4775 5222
rect 4915 5218 4919 5222
rect 4955 5218 4959 5222
rect 5067 5218 5071 5222
rect 5147 5218 5151 5222
rect 5219 5218 5223 5222
rect 5379 5218 5383 5222
rect 5515 5218 5519 5222
rect 5663 5218 5667 5222
rect 1975 5102 1979 5106
rect 2119 5102 2123 5106
rect 2303 5102 2307 5106
rect 2327 5102 2331 5106
rect 2503 5102 2507 5106
rect 2535 5102 2539 5106
rect 2711 5102 2715 5106
rect 2751 5102 2755 5106
rect 2919 5102 2923 5106
rect 2975 5102 2979 5106
rect 3127 5102 3131 5106
rect 3207 5102 3211 5106
rect 3335 5102 3339 5106
rect 3799 5102 3803 5106
rect 111 5074 115 5078
rect 155 5074 159 5078
rect 379 5074 383 5078
rect 419 5074 423 5078
rect 595 5074 599 5078
rect 627 5074 631 5078
rect 779 5074 783 5078
rect 899 5074 903 5078
rect 971 5074 975 5078
rect 1171 5074 1175 5078
rect 1195 5074 1199 5078
rect 1371 5074 1375 5078
rect 1499 5074 1503 5078
rect 1579 5074 1583 5078
rect 1787 5074 1791 5078
rect 1935 5074 1939 5078
rect 3839 5098 3843 5102
rect 3887 5098 3891 5102
rect 4087 5098 4091 5102
rect 4327 5098 4331 5102
rect 4463 5098 4467 5102
rect 4567 5098 4571 5102
rect 4623 5098 4627 5102
rect 4783 5098 4787 5102
rect 4815 5098 4819 5102
rect 4943 5098 4947 5102
rect 5063 5098 5067 5102
rect 5095 5098 5099 5102
rect 5247 5098 5251 5102
rect 5311 5098 5315 5102
rect 5407 5098 5411 5102
rect 5543 5098 5547 5102
rect 5663 5098 5667 5102
rect 1975 4982 1979 4986
rect 1995 4982 1999 4986
rect 2091 4982 2095 4986
rect 2131 4982 2135 4986
rect 2267 4982 2271 4986
rect 2299 4982 2303 4986
rect 2419 4982 2423 4986
rect 2507 4982 2511 4986
rect 2619 4982 2623 4986
rect 2723 4982 2727 4986
rect 2859 4982 2863 4986
rect 2947 4982 2951 4986
rect 3123 4982 3127 4986
rect 3179 4982 3183 4986
rect 3395 4982 3399 4986
rect 3651 4982 3655 4986
rect 3799 4982 3803 4986
rect 3839 4986 3843 4990
rect 3859 4986 3863 4990
rect 3995 4986 3999 4990
rect 4059 4986 4063 4990
rect 4131 4986 4135 4990
rect 4267 4986 4271 4990
rect 4299 4986 4303 4990
rect 4403 4986 4407 4990
rect 4539 4986 4543 4990
rect 4675 4986 4679 4990
rect 4787 4986 4791 4990
rect 4811 4986 4815 4990
rect 4947 4986 4951 4990
rect 5035 4986 5039 4990
rect 5083 4986 5087 4990
rect 5227 4986 5231 4990
rect 5283 4986 5287 4990
rect 5379 4986 5383 4990
rect 5515 4986 5519 4990
rect 5663 4986 5667 4990
rect 111 4934 115 4938
rect 159 4934 163 4938
rect 183 4934 187 4938
rect 295 4934 299 4938
rect 407 4934 411 4938
rect 431 4934 435 4938
rect 567 4934 571 4938
rect 655 4934 659 4938
rect 703 4934 707 4938
rect 927 4934 931 4938
rect 1223 4934 1227 4938
rect 1527 4934 1531 4938
rect 1815 4934 1819 4938
rect 1935 4934 1939 4938
rect 1975 4862 1979 4866
rect 2023 4862 2027 4866
rect 2159 4862 2163 4866
rect 2295 4862 2299 4866
rect 2327 4862 2331 4866
rect 2447 4862 2451 4866
rect 2559 4862 2563 4866
rect 2647 4862 2651 4866
rect 2823 4862 2827 4866
rect 2887 4862 2891 4866
rect 3103 4862 3107 4866
rect 3151 4862 3155 4866
rect 3399 4862 3403 4866
rect 3423 4862 3427 4866
rect 3679 4862 3683 4866
rect 3799 4862 3803 4866
rect 111 4810 115 4814
rect 131 4810 135 4814
rect 267 4810 271 4814
rect 403 4810 407 4814
rect 539 4810 543 4814
rect 675 4810 679 4814
rect 1935 4810 1939 4814
rect 3839 4798 3843 4802
rect 3887 4798 3891 4802
rect 4023 4798 4027 4802
rect 4071 4798 4075 4802
rect 4159 4798 4163 4802
rect 4295 4798 4299 4802
rect 4431 4798 4435 4802
rect 4535 4798 4539 4802
rect 4567 4798 4571 4802
rect 4703 4798 4707 4802
rect 4783 4798 4787 4802
rect 4839 4798 4843 4802
rect 4975 4798 4979 4802
rect 5039 4798 5043 4802
rect 5111 4798 5115 4802
rect 5255 4798 5259 4802
rect 5303 4798 5307 4802
rect 5407 4798 5411 4802
rect 5543 4798 5547 4802
rect 5663 4798 5667 4802
rect 1975 4738 1979 4742
rect 2019 4738 2023 4742
rect 2195 4738 2199 4742
rect 2299 4738 2303 4742
rect 2371 4738 2375 4742
rect 2531 4738 2535 4742
rect 2547 4738 2551 4742
rect 2723 4738 2727 4742
rect 2795 4738 2799 4742
rect 3075 4738 3079 4742
rect 3371 4738 3375 4742
rect 3651 4738 3655 4742
rect 3799 4738 3803 4742
rect 111 4694 115 4698
rect 159 4694 163 4698
rect 295 4694 299 4698
rect 431 4694 435 4698
rect 567 4694 571 4698
rect 703 4694 707 4698
rect 1935 4694 1939 4698
rect 3839 4686 3843 4690
rect 3859 4686 3863 4690
rect 3995 4686 3999 4690
rect 4043 4686 4047 4690
rect 4131 4686 4135 4690
rect 4267 4686 4271 4690
rect 4403 4686 4407 4690
rect 4507 4686 4511 4690
rect 4539 4686 4543 4690
rect 4675 4686 4679 4690
rect 4755 4686 4759 4690
rect 4819 4686 4823 4690
rect 4963 4686 4967 4690
rect 5011 4686 5015 4690
rect 5107 4686 5111 4690
rect 5243 4686 5247 4690
rect 5275 4686 5279 4690
rect 5379 4686 5383 4690
rect 5515 4686 5519 4690
rect 5663 4686 5667 4690
rect 1975 4622 1979 4626
rect 2023 4622 2027 4626
rect 2047 4622 2051 4626
rect 2223 4622 2227 4626
rect 2263 4622 2267 4626
rect 2399 4622 2403 4626
rect 2527 4622 2531 4626
rect 2575 4622 2579 4626
rect 2751 4622 2755 4626
rect 2775 4622 2779 4626
rect 3015 4622 3019 4626
rect 3247 4622 3251 4626
rect 3471 4622 3475 4626
rect 3679 4622 3683 4626
rect 3799 4622 3803 4626
rect 111 4570 115 4574
rect 131 4570 135 4574
rect 251 4570 255 4574
rect 267 4570 271 4574
rect 403 4570 407 4574
rect 443 4570 447 4574
rect 539 4570 543 4574
rect 651 4570 655 4574
rect 675 4570 679 4574
rect 875 4570 879 4574
rect 1099 4570 1103 4574
rect 1331 4570 1335 4574
rect 1571 4570 1575 4574
rect 1787 4570 1791 4574
rect 1935 4570 1939 4574
rect 3839 4574 3843 4578
rect 3887 4574 3891 4578
rect 4023 4574 4027 4578
rect 4159 4574 4163 4578
rect 4295 4574 4299 4578
rect 4431 4574 4435 4578
rect 4567 4574 4571 4578
rect 4671 4574 4675 4578
rect 4703 4574 4707 4578
rect 4807 4574 4811 4578
rect 4847 4574 4851 4578
rect 4943 4574 4947 4578
rect 4991 4574 4995 4578
rect 5079 4574 5083 4578
rect 5135 4574 5139 4578
rect 5271 4574 5275 4578
rect 5407 4574 5411 4578
rect 5543 4574 5547 4578
rect 5663 4574 5667 4578
rect 1975 4498 1979 4502
rect 1995 4498 1999 4502
rect 2235 4498 2239 4502
rect 2267 4498 2271 4502
rect 2499 4498 2503 4502
rect 2515 4498 2519 4502
rect 2747 4498 2751 4502
rect 2971 4498 2975 4502
rect 2987 4498 2991 4502
rect 3187 4498 3191 4502
rect 3219 4498 3223 4502
rect 3395 4498 3399 4502
rect 3443 4498 3447 4502
rect 3611 4498 3615 4502
rect 3651 4498 3655 4502
rect 3799 4498 3803 4502
rect 111 4458 115 4462
rect 279 4458 283 4462
rect 471 4458 475 4462
rect 511 4458 515 4462
rect 679 4458 683 4462
rect 687 4458 691 4462
rect 871 4458 875 4462
rect 903 4458 907 4462
rect 1071 4458 1075 4462
rect 1127 4458 1131 4462
rect 1279 4458 1283 4462
rect 1359 4458 1363 4462
rect 1495 4458 1499 4462
rect 1599 4458 1603 4462
rect 1719 4458 1723 4462
rect 1815 4458 1819 4462
rect 1935 4458 1939 4462
rect 3839 4458 3843 4462
rect 4347 4458 4351 4462
rect 4483 4458 4487 4462
rect 4619 4458 4623 4462
rect 4643 4458 4647 4462
rect 4755 4458 4759 4462
rect 4779 4458 4783 4462
rect 4891 4458 4895 4462
rect 4915 4458 4919 4462
rect 5051 4458 5055 4462
rect 5663 4458 5667 4462
rect 1975 4374 1979 4378
rect 2023 4374 2027 4378
rect 2199 4374 2203 4378
rect 2295 4374 2299 4378
rect 2399 4374 2403 4378
rect 2543 4374 2547 4378
rect 2591 4374 2595 4378
rect 2775 4374 2779 4378
rect 2951 4374 2955 4378
rect 2999 4374 3003 4378
rect 3135 4374 3139 4378
rect 3215 4374 3219 4378
rect 3319 4374 3323 4378
rect 3423 4374 3427 4378
rect 3639 4374 3643 4378
rect 3799 4374 3803 4378
rect 111 4342 115 4346
rect 483 4342 487 4346
rect 659 4342 663 4346
rect 715 4342 719 4346
rect 843 4342 847 4346
rect 851 4342 855 4346
rect 987 4342 991 4346
rect 1043 4342 1047 4346
rect 1123 4342 1127 4346
rect 1251 4342 1255 4346
rect 1259 4342 1263 4346
rect 1395 4342 1399 4346
rect 1467 4342 1471 4346
rect 1531 4342 1535 4346
rect 1667 4342 1671 4346
rect 1691 4342 1695 4346
rect 1935 4342 1939 4346
rect 3839 4330 3843 4334
rect 4135 4330 4139 4334
rect 4271 4330 4275 4334
rect 4375 4330 4379 4334
rect 4407 4330 4411 4334
rect 4511 4330 4515 4334
rect 4543 4330 4547 4334
rect 4647 4330 4651 4334
rect 4679 4330 4683 4334
rect 4783 4330 4787 4334
rect 4919 4330 4923 4334
rect 5663 4330 5667 4334
rect 1975 4258 1979 4262
rect 1995 4258 1999 4262
rect 2171 4258 2175 4262
rect 2243 4258 2247 4262
rect 2371 4258 2375 4262
rect 2507 4258 2511 4262
rect 2563 4258 2567 4262
rect 2747 4258 2751 4262
rect 2763 4258 2767 4262
rect 2923 4258 2927 4262
rect 3019 4258 3023 4262
rect 3107 4258 3111 4262
rect 3283 4258 3287 4262
rect 3291 4258 3295 4262
rect 3799 4258 3803 4262
rect 111 4222 115 4226
rect 727 4222 731 4226
rect 743 4222 747 4226
rect 863 4222 867 4226
rect 879 4222 883 4226
rect 999 4222 1003 4226
rect 1015 4222 1019 4226
rect 1135 4222 1139 4226
rect 1151 4222 1155 4226
rect 1271 4222 1275 4226
rect 1287 4222 1291 4226
rect 1407 4222 1411 4226
rect 1423 4222 1427 4226
rect 1543 4222 1547 4226
rect 1559 4222 1563 4226
rect 1679 4222 1683 4226
rect 1695 4222 1699 4226
rect 1815 4222 1819 4226
rect 1935 4222 1939 4226
rect 3839 4206 3843 4210
rect 3971 4206 3975 4210
rect 4107 4206 4111 4210
rect 4243 4206 4247 4210
rect 4379 4206 4383 4210
rect 4515 4206 4519 4210
rect 4651 4206 4655 4210
rect 5663 4206 5667 4210
rect 1975 4134 1979 4138
rect 2023 4134 2027 4138
rect 2271 4134 2275 4138
rect 2535 4134 2539 4138
rect 2791 4134 2795 4138
rect 3047 4134 3051 4138
rect 3135 4134 3139 4138
rect 3271 4134 3275 4138
rect 3311 4134 3315 4138
rect 3407 4134 3411 4138
rect 3543 4134 3547 4138
rect 3679 4134 3683 4138
rect 3799 4134 3803 4138
rect 111 4110 115 4114
rect 563 4110 567 4114
rect 699 4110 703 4114
rect 835 4110 839 4114
rect 971 4110 975 4114
rect 1107 4110 1111 4114
rect 1243 4110 1247 4114
rect 1379 4110 1383 4114
rect 1515 4110 1519 4114
rect 1651 4110 1655 4114
rect 1787 4110 1791 4114
rect 1935 4110 1939 4114
rect 111 3998 115 4002
rect 159 3998 163 4002
rect 327 3998 331 4002
rect 535 3998 539 4002
rect 591 3998 595 4002
rect 727 3998 731 4002
rect 751 3998 755 4002
rect 863 3998 867 4002
rect 967 3998 971 4002
rect 999 3998 1003 4002
rect 1135 3998 1139 4002
rect 1183 3998 1187 4002
rect 1271 3998 1275 4002
rect 1399 3998 1403 4002
rect 1407 3998 1411 4002
rect 1543 3998 1547 4002
rect 1615 3998 1619 4002
rect 1679 3998 1683 4002
rect 1815 3998 1819 4002
rect 1935 3998 1939 4002
rect 3839 4070 3843 4074
rect 3887 4070 3891 4074
rect 3999 4070 4003 4074
rect 4023 4070 4027 4074
rect 4135 4070 4139 4074
rect 4159 4070 4163 4074
rect 4271 4070 4275 4074
rect 4295 4070 4299 4074
rect 4407 4070 4411 4074
rect 4431 4070 4435 4074
rect 4543 4070 4547 4074
rect 4567 4070 4571 4074
rect 4703 4070 4707 4074
rect 4839 4070 4843 4074
rect 5663 4070 5667 4074
rect 3839 3958 3843 3962
rect 3859 3958 3863 3962
rect 3995 3958 3999 3962
rect 4131 3958 4135 3962
rect 4147 3958 4151 3962
rect 4267 3958 4271 3962
rect 4299 3958 4303 3962
rect 4403 3958 4407 3962
rect 4459 3958 4463 3962
rect 4539 3958 4543 3962
rect 4619 3958 4623 3962
rect 4675 3958 4679 3962
rect 4779 3958 4783 3962
rect 4811 3958 4815 3962
rect 5663 3958 5667 3962
rect 1975 3930 1979 3934
rect 1995 3930 1999 3934
rect 2403 3930 2407 3934
rect 2827 3930 2831 3934
rect 3107 3930 3111 3934
rect 3243 3930 3247 3934
rect 3251 3930 3255 3934
rect 3379 3930 3383 3934
rect 3515 3930 3519 3934
rect 3651 3930 3655 3934
rect 3799 3930 3803 3934
rect 111 3886 115 3890
rect 131 3886 135 3890
rect 299 3886 303 3890
rect 355 3886 359 3890
rect 507 3886 511 3890
rect 619 3886 623 3890
rect 723 3886 727 3890
rect 899 3886 903 3890
rect 939 3886 943 3890
rect 1155 3886 1159 3890
rect 1195 3886 1199 3890
rect 1371 3886 1375 3890
rect 1499 3886 1503 3890
rect 1587 3886 1591 3890
rect 1787 3886 1791 3890
rect 1935 3886 1939 3890
rect 1975 3818 1979 3822
rect 2023 3818 2027 3822
rect 2175 3818 2179 3822
rect 2351 3818 2355 3822
rect 2431 3818 2435 3822
rect 2535 3818 2539 3822
rect 2719 3818 2723 3822
rect 2855 3818 2859 3822
rect 2895 3818 2899 3822
rect 3071 3818 3075 3822
rect 3247 3818 3251 3822
rect 3279 3818 3283 3822
rect 3423 3818 3427 3822
rect 3607 3818 3611 3822
rect 3679 3818 3683 3822
rect 3799 3818 3803 3822
rect 3839 3818 3843 3822
rect 3887 3818 3891 3822
rect 4023 3818 4027 3822
rect 4175 3818 4179 3822
rect 4327 3818 4331 3822
rect 4487 3818 4491 3822
rect 4503 3818 4507 3822
rect 4639 3818 4643 3822
rect 4647 3818 4651 3822
rect 4775 3818 4779 3822
rect 4807 3818 4811 3822
rect 4911 3818 4915 3822
rect 5047 3818 5051 3822
rect 5663 3818 5667 3822
rect 111 3762 115 3766
rect 159 3762 163 3766
rect 247 3762 251 3766
rect 383 3762 387 3766
rect 519 3762 523 3766
rect 647 3762 651 3766
rect 791 3762 795 3766
rect 927 3762 931 3766
rect 1063 3762 1067 3766
rect 1223 3762 1227 3766
rect 1343 3762 1347 3766
rect 1527 3762 1531 3766
rect 1815 3762 1819 3766
rect 1935 3762 1939 3766
rect 1975 3698 1979 3702
rect 1995 3698 1999 3702
rect 2011 3698 2015 3702
rect 2147 3698 2151 3702
rect 2291 3698 2295 3702
rect 2323 3698 2327 3702
rect 2435 3698 2439 3702
rect 2507 3698 2511 3702
rect 2579 3698 2583 3702
rect 2691 3698 2695 3702
rect 2723 3698 2727 3702
rect 2867 3698 2871 3702
rect 3011 3698 3015 3702
rect 3043 3698 3047 3702
rect 3155 3698 3159 3702
rect 3219 3698 3223 3702
rect 3299 3698 3303 3702
rect 3395 3698 3399 3702
rect 3579 3698 3583 3702
rect 3799 3698 3803 3702
rect 111 3634 115 3638
rect 219 3634 223 3638
rect 491 3634 495 3638
rect 635 3634 639 3638
rect 763 3634 767 3638
rect 779 3634 783 3638
rect 923 3634 927 3638
rect 1035 3634 1039 3638
rect 1067 3634 1071 3638
rect 1211 3634 1215 3638
rect 1315 3634 1319 3638
rect 1935 3634 1939 3638
rect 3839 3686 3843 3690
rect 4019 3686 4023 3690
rect 4155 3686 4159 3690
rect 4291 3686 4295 3690
rect 4427 3686 4431 3690
rect 4475 3686 4479 3690
rect 4563 3686 4567 3690
rect 4611 3686 4615 3690
rect 4699 3686 4703 3690
rect 4747 3686 4751 3690
rect 4835 3686 4839 3690
rect 4883 3686 4887 3690
rect 4971 3686 4975 3690
rect 5019 3686 5023 3690
rect 5107 3686 5111 3690
rect 5243 3686 5247 3690
rect 5379 3686 5383 3690
rect 5515 3686 5519 3690
rect 5663 3686 5667 3690
rect 1975 3578 1979 3582
rect 2039 3578 2043 3582
rect 2175 3578 2179 3582
rect 2239 3578 2243 3582
rect 2319 3578 2323 3582
rect 2375 3578 2379 3582
rect 2463 3578 2467 3582
rect 2511 3578 2515 3582
rect 2607 3578 2611 3582
rect 2647 3578 2651 3582
rect 2751 3578 2755 3582
rect 2783 3578 2787 3582
rect 2895 3578 2899 3582
rect 2919 3578 2923 3582
rect 3039 3578 3043 3582
rect 3055 3578 3059 3582
rect 3183 3578 3187 3582
rect 3191 3578 3195 3582
rect 3327 3578 3331 3582
rect 3463 3578 3467 3582
rect 3799 3578 3803 3582
rect 111 3502 115 3506
rect 431 3502 435 3506
rect 519 3502 523 3506
rect 567 3502 571 3506
rect 663 3502 667 3506
rect 703 3502 707 3506
rect 807 3502 811 3506
rect 839 3502 843 3506
rect 951 3502 955 3506
rect 975 3502 979 3506
rect 1095 3502 1099 3506
rect 1239 3502 1243 3506
rect 1935 3502 1939 3506
rect 3839 3526 3843 3530
rect 4047 3526 4051 3530
rect 4183 3526 4187 3530
rect 4319 3526 4323 3530
rect 4455 3526 4459 3530
rect 4591 3526 4595 3530
rect 4727 3526 4731 3530
rect 4863 3526 4867 3530
rect 4999 3526 5003 3530
rect 5135 3526 5139 3530
rect 5271 3526 5275 3530
rect 5407 3526 5411 3530
rect 5543 3526 5547 3530
rect 5663 3526 5667 3530
rect 1975 3462 1979 3466
rect 2171 3462 2175 3466
rect 2211 3462 2215 3466
rect 2347 3462 2351 3466
rect 2483 3462 2487 3466
rect 2531 3462 2535 3466
rect 2619 3462 2623 3466
rect 2715 3462 2719 3466
rect 2755 3462 2759 3466
rect 2891 3462 2895 3466
rect 2907 3462 2911 3466
rect 3027 3462 3031 3466
rect 3099 3462 3103 3466
rect 3163 3462 3167 3466
rect 3291 3462 3295 3466
rect 3299 3462 3303 3466
rect 3435 3462 3439 3466
rect 3483 3462 3487 3466
rect 3651 3462 3655 3466
rect 3799 3462 3803 3466
rect 3839 3406 3843 3410
rect 3859 3406 3863 3410
rect 4099 3406 4103 3410
rect 4347 3406 4351 3410
rect 4587 3406 4591 3410
rect 4811 3406 4815 3410
rect 5027 3406 5031 3410
rect 5235 3406 5239 3410
rect 5379 3406 5383 3410
rect 5451 3406 5455 3410
rect 5515 3406 5519 3410
rect 5663 3406 5667 3410
rect 111 3382 115 3386
rect 323 3382 327 3386
rect 403 3382 407 3386
rect 459 3382 463 3386
rect 539 3382 543 3386
rect 595 3382 599 3386
rect 675 3382 679 3386
rect 731 3382 735 3386
rect 811 3382 815 3386
rect 867 3382 871 3386
rect 947 3382 951 3386
rect 1935 3382 1939 3386
rect 1975 3326 1979 3330
rect 2151 3326 2155 3330
rect 2199 3326 2203 3330
rect 2375 3326 2379 3330
rect 2399 3326 2403 3330
rect 2559 3326 2563 3330
rect 2687 3326 2691 3330
rect 2743 3326 2747 3330
rect 2935 3326 2939 3330
rect 3015 3326 3019 3330
rect 3127 3326 3131 3330
rect 3319 3326 3323 3330
rect 3359 3326 3363 3330
rect 3511 3326 3515 3330
rect 3679 3326 3683 3330
rect 3799 3326 3803 3330
rect 3839 3294 3843 3298
rect 3887 3294 3891 3298
rect 4127 3294 4131 3298
rect 4375 3294 4379 3298
rect 4607 3294 4611 3298
rect 4615 3294 4619 3298
rect 4815 3294 4819 3298
rect 4839 3294 4843 3298
rect 5015 3294 5019 3298
rect 5055 3294 5059 3298
rect 5199 3294 5203 3298
rect 5263 3294 5267 3298
rect 5383 3294 5387 3298
rect 5479 3294 5483 3298
rect 5543 3294 5547 3298
rect 5663 3294 5667 3298
rect 111 3262 115 3266
rect 159 3262 163 3266
rect 335 3262 339 3266
rect 351 3262 355 3266
rect 487 3262 491 3266
rect 543 3262 547 3266
rect 623 3262 627 3266
rect 751 3262 755 3266
rect 759 3262 763 3266
rect 895 3262 899 3266
rect 959 3262 963 3266
rect 1935 3262 1939 3266
rect 1975 3214 1979 3218
rect 1995 3214 1999 3218
rect 2123 3214 2127 3218
rect 2147 3214 2151 3218
rect 2347 3214 2351 3218
rect 2371 3214 2375 3218
rect 2555 3214 2559 3218
rect 2659 3214 2663 3218
rect 2771 3214 2775 3218
rect 2987 3214 2991 3218
rect 3211 3214 3215 3218
rect 3331 3214 3335 3218
rect 3443 3214 3447 3218
rect 3651 3214 3655 3218
rect 3799 3214 3803 3218
rect 3839 3166 3843 3170
rect 3859 3166 3863 3170
rect 4099 3166 4103 3170
rect 4347 3166 4351 3170
rect 4467 3166 4471 3170
rect 4579 3166 4583 3170
rect 4651 3166 4655 3170
rect 4787 3166 4791 3170
rect 4859 3166 4863 3170
rect 4987 3166 4991 3170
rect 5075 3166 5079 3170
rect 5171 3166 5175 3170
rect 5307 3166 5311 3170
rect 5355 3166 5359 3170
rect 5515 3166 5519 3170
rect 5663 3166 5667 3170
rect 111 3134 115 3138
rect 131 3134 135 3138
rect 307 3134 311 3138
rect 371 3134 375 3138
rect 515 3134 519 3138
rect 627 3134 631 3138
rect 723 3134 727 3138
rect 875 3134 879 3138
rect 931 3134 935 3138
rect 1115 3134 1119 3138
rect 1347 3134 1351 3138
rect 1579 3134 1583 3138
rect 1787 3134 1791 3138
rect 1935 3134 1939 3138
rect 1975 3102 1979 3106
rect 2023 3102 2027 3106
rect 2175 3102 2179 3106
rect 2375 3102 2379 3106
rect 2583 3102 2587 3106
rect 2647 3102 2651 3106
rect 2783 3102 2787 3106
rect 2799 3102 2803 3106
rect 2927 3102 2931 3106
rect 3015 3102 3019 3106
rect 3079 3102 3083 3106
rect 3239 3102 3243 3106
rect 3399 3102 3403 3106
rect 3471 3102 3475 3106
rect 3567 3102 3571 3106
rect 3679 3102 3683 3106
rect 3799 3102 3803 3106
rect 111 3022 115 3026
rect 159 3022 163 3026
rect 175 3022 179 3026
rect 399 3022 403 3026
rect 407 3022 411 3026
rect 623 3022 627 3026
rect 655 3022 659 3026
rect 823 3022 827 3026
rect 903 3022 907 3026
rect 1007 3022 1011 3026
rect 1143 3022 1147 3026
rect 1183 3022 1187 3026
rect 1351 3022 1355 3026
rect 1375 3022 1379 3026
rect 1511 3022 1515 3026
rect 1607 3022 1611 3026
rect 1671 3022 1675 3026
rect 1815 3022 1819 3026
rect 1935 3022 1939 3026
rect 3839 3054 3843 3058
rect 4255 3054 4259 3058
rect 4455 3054 4459 3058
rect 4495 3054 4499 3058
rect 4671 3054 4675 3058
rect 4679 3054 4683 3058
rect 4887 3054 4891 3058
rect 4911 3054 4915 3058
rect 5103 3054 5107 3058
rect 5167 3054 5171 3058
rect 5335 3054 5339 3058
rect 5423 3054 5427 3058
rect 5543 3054 5547 3058
rect 5663 3054 5667 3058
rect 1975 2990 1979 2994
rect 2619 2990 2623 2994
rect 2755 2990 2759 2994
rect 2803 2990 2807 2994
rect 2899 2990 2903 2994
rect 2939 2990 2943 2994
rect 3051 2990 3055 2994
rect 3075 2990 3079 2994
rect 3211 2990 3215 2994
rect 3347 2990 3351 2994
rect 3371 2990 3375 2994
rect 3483 2990 3487 2994
rect 3539 2990 3543 2994
rect 3799 2990 3803 2994
rect 3839 2918 3843 2922
rect 3995 2918 3999 2922
rect 4211 2918 4215 2922
rect 4227 2918 4231 2922
rect 4427 2918 4431 2922
rect 4443 2918 4447 2922
rect 4643 2918 4647 2922
rect 4699 2918 4703 2922
rect 4883 2918 4887 2922
rect 4971 2918 4975 2922
rect 5139 2918 5143 2922
rect 5251 2918 5255 2922
rect 5395 2918 5399 2922
rect 5515 2918 5519 2922
rect 5663 2918 5667 2922
rect 111 2906 115 2910
rect 147 2906 151 2910
rect 379 2906 383 2910
rect 395 2906 399 2910
rect 595 2906 599 2910
rect 787 2906 791 2910
rect 795 2906 799 2910
rect 971 2906 975 2910
rect 979 2906 983 2910
rect 1147 2906 1151 2910
rect 1155 2906 1159 2910
rect 1315 2906 1319 2910
rect 1323 2906 1327 2910
rect 1483 2906 1487 2910
rect 1643 2906 1647 2910
rect 1787 2906 1791 2910
rect 1935 2906 1939 2910
rect 1975 2826 1979 2830
rect 2023 2826 2027 2830
rect 2167 2826 2171 2830
rect 2335 2826 2339 2830
rect 2495 2826 2499 2830
rect 2663 2826 2667 2830
rect 2831 2826 2835 2830
rect 2967 2826 2971 2830
rect 2999 2826 3003 2830
rect 3103 2826 3107 2830
rect 3167 2826 3171 2830
rect 3239 2826 3243 2830
rect 3375 2826 3379 2830
rect 3511 2826 3515 2830
rect 3799 2826 3803 2830
rect 3839 2802 3843 2806
rect 3919 2802 3923 2806
rect 4023 2802 4027 2806
rect 4055 2802 4059 2806
rect 4191 2802 4195 2806
rect 4239 2802 4243 2806
rect 4327 2802 4331 2806
rect 4463 2802 4467 2806
rect 4471 2802 4475 2806
rect 4727 2802 4731 2806
rect 4999 2802 5003 2806
rect 5279 2802 5283 2806
rect 5543 2802 5547 2806
rect 5663 2802 5667 2806
rect 111 2782 115 2786
rect 423 2782 427 2786
rect 623 2782 627 2786
rect 655 2782 659 2786
rect 815 2782 819 2786
rect 975 2782 979 2786
rect 999 2782 1003 2786
rect 1143 2782 1147 2786
rect 1175 2782 1179 2786
rect 1311 2782 1315 2786
rect 1343 2782 1347 2786
rect 1479 2782 1483 2786
rect 1511 2782 1515 2786
rect 1671 2782 1675 2786
rect 1815 2782 1819 2786
rect 1935 2782 1939 2786
rect 1975 2714 1979 2718
rect 1995 2714 1999 2718
rect 2139 2714 2143 2718
rect 2307 2714 2311 2718
rect 2379 2714 2383 2718
rect 2467 2714 2471 2718
rect 2515 2714 2519 2718
rect 2635 2714 2639 2718
rect 2659 2714 2663 2718
rect 2803 2714 2807 2718
rect 2947 2714 2951 2718
rect 2971 2714 2975 2718
rect 3091 2714 3095 2718
rect 3139 2714 3143 2718
rect 3235 2714 3239 2718
rect 3799 2714 3803 2718
rect 111 2670 115 2674
rect 627 2670 631 2674
rect 771 2670 775 2674
rect 787 2670 791 2674
rect 907 2670 911 2674
rect 947 2670 951 2674
rect 1043 2670 1047 2674
rect 1115 2670 1119 2674
rect 1179 2670 1183 2674
rect 1283 2670 1287 2674
rect 1315 2670 1319 2674
rect 1451 2670 1455 2674
rect 1587 2670 1591 2674
rect 1723 2670 1727 2674
rect 1935 2670 1939 2674
rect 3839 2678 3843 2682
rect 3891 2678 3895 2682
rect 4027 2678 4031 2682
rect 4099 2678 4103 2682
rect 4163 2678 4167 2682
rect 4299 2678 4303 2682
rect 4435 2678 4439 2682
rect 4515 2678 4519 2682
rect 4755 2678 4759 2682
rect 5011 2678 5015 2682
rect 5275 2678 5279 2682
rect 5515 2678 5519 2682
rect 5663 2678 5667 2682
rect 1975 2598 1979 2602
rect 2407 2598 2411 2602
rect 2511 2598 2515 2602
rect 2543 2598 2547 2602
rect 2647 2598 2651 2602
rect 2687 2598 2691 2602
rect 2783 2598 2787 2602
rect 2831 2598 2835 2602
rect 2919 2598 2923 2602
rect 2975 2598 2979 2602
rect 3055 2598 3059 2602
rect 3119 2598 3123 2602
rect 3191 2598 3195 2602
rect 3263 2598 3267 2602
rect 3327 2598 3331 2602
rect 3463 2598 3467 2602
rect 3799 2598 3803 2602
rect 3839 2562 3843 2566
rect 4127 2562 4131 2566
rect 4327 2562 4331 2566
rect 4495 2562 4499 2566
rect 4543 2562 4547 2566
rect 4631 2562 4635 2566
rect 4767 2562 4771 2566
rect 4783 2562 4787 2566
rect 4903 2562 4907 2566
rect 5039 2562 5043 2566
rect 5303 2562 5307 2566
rect 5543 2562 5547 2566
rect 5663 2562 5667 2566
rect 111 2542 115 2546
rect 551 2542 555 2546
rect 687 2542 691 2546
rect 799 2542 803 2546
rect 831 2542 835 2546
rect 935 2542 939 2546
rect 983 2542 987 2546
rect 1071 2542 1075 2546
rect 1135 2542 1139 2546
rect 1207 2542 1211 2546
rect 1295 2542 1299 2546
rect 1343 2542 1347 2546
rect 1455 2542 1459 2546
rect 1479 2542 1483 2546
rect 1615 2542 1619 2546
rect 1751 2542 1755 2546
rect 1783 2542 1787 2546
rect 1935 2542 1939 2546
rect 1975 2470 1979 2474
rect 2307 2470 2311 2474
rect 2483 2470 2487 2474
rect 2515 2470 2519 2474
rect 2619 2470 2623 2474
rect 2715 2470 2719 2474
rect 2755 2470 2759 2474
rect 2891 2470 2895 2474
rect 2907 2470 2911 2474
rect 3027 2470 3031 2474
rect 3099 2470 3103 2474
rect 3163 2470 3167 2474
rect 3283 2470 3287 2474
rect 3299 2470 3303 2474
rect 3435 2470 3439 2474
rect 3467 2470 3471 2474
rect 3651 2470 3655 2474
rect 3799 2470 3803 2474
rect 111 2418 115 2422
rect 131 2418 135 2422
rect 339 2418 343 2422
rect 523 2418 527 2422
rect 563 2418 567 2422
rect 659 2418 663 2422
rect 803 2418 807 2422
rect 955 2418 959 2422
rect 1043 2418 1047 2422
rect 1107 2418 1111 2422
rect 1267 2418 1271 2422
rect 1291 2418 1295 2422
rect 1427 2418 1431 2422
rect 1547 2418 1551 2422
rect 1587 2418 1591 2422
rect 1755 2418 1759 2422
rect 1787 2418 1791 2422
rect 1935 2418 1939 2422
rect 3839 2434 3843 2438
rect 4467 2434 4471 2438
rect 4603 2434 4607 2438
rect 4699 2434 4703 2438
rect 4739 2434 4743 2438
rect 4835 2434 4839 2438
rect 4875 2434 4879 2438
rect 4971 2434 4975 2438
rect 5011 2434 5015 2438
rect 5107 2434 5111 2438
rect 5243 2434 5247 2438
rect 5379 2434 5383 2438
rect 5515 2434 5519 2438
rect 5663 2434 5667 2438
rect 1975 2350 1979 2354
rect 2223 2350 2227 2354
rect 2335 2350 2339 2354
rect 2503 2350 2507 2354
rect 2543 2350 2547 2354
rect 2743 2350 2747 2354
rect 2767 2350 2771 2354
rect 2935 2350 2939 2354
rect 3007 2350 3011 2354
rect 3127 2350 3131 2354
rect 3239 2350 3243 2354
rect 3311 2350 3315 2354
rect 3471 2350 3475 2354
rect 3495 2350 3499 2354
rect 3679 2350 3683 2354
rect 3799 2350 3803 2354
rect 3839 2310 3843 2314
rect 111 2302 115 2306
rect 159 2302 163 2306
rect 319 2302 323 2306
rect 367 2302 371 2306
rect 551 2302 555 2306
rect 591 2302 595 2306
rect 831 2302 835 2306
rect 1071 2302 1075 2306
rect 1151 2302 1155 2306
rect 1319 2302 1323 2306
rect 1495 2302 1499 2306
rect 1575 2302 1579 2306
rect 1815 2302 1819 2306
rect 1935 2302 1939 2306
rect 3887 2310 3891 2314
rect 4183 2310 4187 2314
rect 4495 2310 4499 2314
rect 4727 2310 4731 2314
rect 4791 2310 4795 2314
rect 4863 2310 4867 2314
rect 4999 2310 5003 2314
rect 5087 2310 5091 2314
rect 5135 2310 5139 2314
rect 5271 2310 5275 2314
rect 5383 2310 5387 2314
rect 5407 2310 5411 2314
rect 5543 2310 5547 2314
rect 5663 2310 5667 2314
rect 1975 2238 1979 2242
rect 1995 2238 1999 2242
rect 2155 2238 2159 2242
rect 2195 2238 2199 2242
rect 2387 2238 2391 2242
rect 2475 2238 2479 2242
rect 2667 2238 2671 2242
rect 2739 2238 2743 2242
rect 2979 2238 2983 2242
rect 2987 2238 2991 2242
rect 3211 2238 3215 2242
rect 3331 2238 3335 2242
rect 3443 2238 3447 2242
rect 3651 2238 3655 2242
rect 3799 2238 3803 2242
rect 3839 2194 3843 2198
rect 3859 2194 3863 2198
rect 3995 2194 3999 2198
rect 4131 2194 4135 2198
rect 4155 2194 4159 2198
rect 4267 2194 4271 2198
rect 4403 2194 4407 2198
rect 4467 2194 4471 2198
rect 4539 2194 4543 2198
rect 4699 2194 4703 2198
rect 4763 2194 4767 2198
rect 4891 2194 4895 2198
rect 5059 2194 5063 2198
rect 5099 2194 5103 2198
rect 5315 2194 5319 2198
rect 5355 2194 5359 2198
rect 5515 2194 5519 2198
rect 5663 2194 5667 2198
rect 111 2166 115 2170
rect 131 2166 135 2170
rect 291 2166 295 2170
rect 483 2166 487 2170
rect 523 2166 527 2170
rect 691 2166 695 2170
rect 803 2166 807 2170
rect 915 2166 919 2170
rect 1123 2166 1127 2170
rect 1147 2166 1151 2170
rect 1387 2166 1391 2170
rect 1467 2166 1471 2170
rect 1635 2166 1639 2170
rect 1787 2166 1791 2170
rect 1935 2166 1939 2170
rect 111 2050 115 2054
rect 263 2050 267 2054
rect 319 2050 323 2054
rect 399 2050 403 2054
rect 511 2050 515 2054
rect 535 2050 539 2054
rect 679 2050 683 2054
rect 719 2050 723 2054
rect 823 2050 827 2054
rect 943 2050 947 2054
rect 967 2050 971 2054
rect 1111 2050 1115 2054
rect 1175 2050 1179 2054
rect 1255 2050 1259 2054
rect 1399 2050 1403 2054
rect 1415 2050 1419 2054
rect 1543 2050 1547 2054
rect 1663 2050 1667 2054
rect 1679 2050 1683 2054
rect 1815 2050 1819 2054
rect 1935 2050 1939 2054
rect 3839 2062 3843 2066
rect 3887 2062 3891 2066
rect 4023 2062 4027 2066
rect 4159 2062 4163 2066
rect 4295 2062 4299 2066
rect 4431 2062 4435 2066
rect 4567 2062 4571 2066
rect 4719 2062 4723 2066
rect 4727 2062 4731 2066
rect 4895 2062 4899 2066
rect 4919 2062 4923 2066
rect 5087 2062 5091 2066
rect 5127 2062 5131 2066
rect 5279 2062 5283 2066
rect 5343 2062 5347 2066
rect 5479 2062 5483 2066
rect 5543 2062 5547 2066
rect 5663 2062 5667 2066
rect 3839 1950 3843 1954
rect 3859 1950 3863 1954
rect 3995 1950 3999 1954
rect 4043 1950 4047 1954
rect 4131 1950 4135 1954
rect 4267 1950 4271 1954
rect 4283 1950 4287 1954
rect 4403 1950 4407 1954
rect 4539 1950 4543 1954
rect 4563 1950 4567 1954
rect 4691 1950 4695 1954
rect 4867 1950 4871 1954
rect 4875 1950 4879 1954
rect 5059 1950 5063 1954
rect 5203 1950 5207 1954
rect 5251 1950 5255 1954
rect 5451 1950 5455 1954
rect 5515 1950 5519 1954
rect 5663 1950 5667 1954
rect 111 1926 115 1930
rect 235 1926 239 1930
rect 371 1926 375 1930
rect 435 1926 439 1930
rect 507 1926 511 1930
rect 627 1926 631 1930
rect 651 1926 655 1930
rect 795 1926 799 1930
rect 811 1926 815 1930
rect 939 1926 943 1930
rect 987 1926 991 1930
rect 1083 1926 1087 1930
rect 1155 1926 1159 1930
rect 1227 1926 1231 1930
rect 1323 1926 1327 1930
rect 1371 1926 1375 1930
rect 1483 1926 1487 1930
rect 1515 1926 1519 1930
rect 1643 1926 1647 1930
rect 1651 1926 1655 1930
rect 1787 1926 1791 1930
rect 1935 1926 1939 1930
rect 1975 1926 1979 1930
rect 2023 1926 2027 1930
rect 2183 1926 2187 1930
rect 2415 1926 2419 1930
rect 2695 1926 2699 1930
rect 3015 1926 3019 1930
rect 3135 1926 3139 1930
rect 3271 1926 3275 1930
rect 3359 1926 3363 1930
rect 3407 1926 3411 1930
rect 3543 1926 3547 1930
rect 3679 1926 3683 1930
rect 3799 1926 3803 1930
rect 3839 1838 3843 1842
rect 3887 1838 3891 1842
rect 4071 1838 4075 1842
rect 4311 1838 4315 1842
rect 4407 1838 4411 1842
rect 4543 1838 4547 1842
rect 4591 1838 4595 1842
rect 4679 1838 4683 1842
rect 4815 1838 4819 1842
rect 4903 1838 4907 1842
rect 4951 1838 4955 1842
rect 5231 1838 5235 1842
rect 5543 1838 5547 1842
rect 5663 1838 5667 1842
rect 111 1802 115 1806
rect 223 1802 227 1806
rect 263 1802 267 1806
rect 463 1802 467 1806
rect 655 1802 659 1806
rect 695 1802 699 1806
rect 839 1802 843 1806
rect 927 1802 931 1806
rect 1015 1802 1019 1806
rect 1159 1802 1163 1806
rect 1183 1802 1187 1806
rect 1351 1802 1355 1806
rect 1391 1802 1395 1806
rect 1511 1802 1515 1806
rect 1671 1802 1675 1806
rect 1815 1802 1819 1806
rect 1935 1802 1939 1806
rect 1975 1802 1979 1806
rect 1995 1802 1999 1806
rect 2131 1802 2135 1806
rect 2267 1802 2271 1806
rect 2419 1802 2423 1806
rect 2579 1802 2583 1806
rect 2739 1802 2743 1806
rect 2899 1802 2903 1806
rect 3051 1802 3055 1806
rect 3107 1802 3111 1806
rect 3203 1802 3207 1806
rect 3243 1802 3247 1806
rect 3355 1802 3359 1806
rect 3379 1802 3383 1806
rect 3515 1802 3519 1806
rect 3651 1802 3655 1806
rect 3799 1802 3803 1806
rect 3839 1710 3843 1714
rect 4379 1710 4383 1714
rect 4515 1710 4519 1714
rect 4563 1710 4567 1714
rect 4651 1710 4655 1714
rect 4699 1710 4703 1714
rect 4787 1710 4791 1714
rect 4835 1710 4839 1714
rect 4923 1710 4927 1714
rect 4971 1710 4975 1714
rect 5107 1710 5111 1714
rect 5243 1710 5247 1714
rect 5379 1710 5383 1714
rect 5515 1710 5519 1714
rect 5663 1710 5667 1714
rect 111 1678 115 1682
rect 131 1678 135 1682
rect 195 1678 199 1682
rect 363 1678 367 1682
rect 435 1678 439 1682
rect 619 1678 623 1682
rect 667 1678 671 1682
rect 875 1678 879 1682
rect 899 1678 903 1682
rect 1131 1678 1135 1682
rect 1139 1678 1143 1682
rect 1363 1678 1367 1682
rect 1935 1678 1939 1682
rect 1975 1678 1979 1682
rect 2023 1678 2027 1682
rect 2159 1678 2163 1682
rect 2167 1678 2171 1682
rect 2295 1678 2299 1682
rect 2319 1678 2323 1682
rect 2447 1678 2451 1682
rect 2479 1678 2483 1682
rect 2607 1678 2611 1682
rect 2639 1678 2643 1682
rect 2767 1678 2771 1682
rect 2791 1678 2795 1682
rect 2927 1678 2931 1682
rect 2943 1678 2947 1682
rect 3079 1678 3083 1682
rect 3103 1678 3107 1682
rect 3231 1678 3235 1682
rect 3263 1678 3267 1682
rect 3383 1678 3387 1682
rect 3423 1678 3427 1682
rect 3543 1678 3547 1682
rect 3679 1678 3683 1682
rect 3799 1678 3803 1682
rect 3839 1582 3843 1586
rect 4591 1582 4595 1586
rect 4727 1582 4731 1586
rect 4863 1582 4867 1586
rect 4999 1582 5003 1586
rect 5135 1582 5139 1586
rect 5271 1582 5275 1586
rect 5407 1582 5411 1586
rect 5543 1582 5547 1586
rect 5663 1582 5667 1586
rect 111 1554 115 1558
rect 159 1554 163 1558
rect 327 1554 331 1558
rect 391 1554 395 1558
rect 511 1554 515 1558
rect 647 1554 651 1558
rect 695 1554 699 1558
rect 887 1554 891 1558
rect 903 1554 907 1558
rect 1079 1554 1083 1558
rect 1167 1554 1171 1558
rect 1935 1554 1939 1558
rect 1975 1554 1979 1558
rect 1995 1554 1999 1558
rect 2131 1554 2135 1558
rect 2139 1554 2143 1558
rect 2267 1554 2271 1558
rect 2291 1554 2295 1558
rect 2403 1554 2407 1558
rect 2451 1554 2455 1558
rect 2539 1554 2543 1558
rect 2611 1554 2615 1558
rect 2675 1554 2679 1558
rect 2763 1554 2767 1558
rect 2811 1554 2815 1558
rect 2915 1554 2919 1558
rect 2947 1554 2951 1558
rect 3075 1554 3079 1558
rect 3083 1554 3087 1558
rect 3219 1554 3223 1558
rect 3235 1554 3239 1558
rect 3355 1554 3359 1558
rect 3395 1554 3399 1558
rect 3491 1554 3495 1558
rect 3799 1554 3803 1558
rect 111 1430 115 1434
rect 131 1430 135 1434
rect 299 1430 303 1434
rect 395 1430 399 1434
rect 483 1430 487 1434
rect 667 1430 671 1434
rect 683 1430 687 1434
rect 859 1430 863 1434
rect 971 1430 975 1434
rect 1051 1430 1055 1434
rect 1259 1430 1263 1434
rect 1935 1430 1939 1434
rect 1975 1430 1979 1434
rect 2023 1430 2027 1434
rect 2159 1430 2163 1434
rect 2167 1430 2171 1434
rect 2295 1430 2299 1434
rect 2303 1430 2307 1434
rect 2431 1430 2435 1434
rect 2439 1430 2443 1434
rect 2567 1430 2571 1434
rect 2575 1430 2579 1434
rect 2703 1430 2707 1434
rect 2711 1430 2715 1434
rect 2839 1430 2843 1434
rect 2847 1430 2851 1434
rect 2975 1430 2979 1434
rect 2983 1430 2987 1434
rect 3111 1430 3115 1434
rect 3119 1430 3123 1434
rect 3247 1430 3251 1434
rect 3255 1430 3259 1434
rect 3383 1430 3387 1434
rect 3519 1430 3523 1434
rect 3799 1430 3803 1434
rect 3839 1398 3843 1402
rect 4563 1398 4567 1402
rect 4699 1398 4703 1402
rect 4811 1398 4815 1402
rect 4835 1398 4839 1402
rect 4947 1398 4951 1402
rect 4971 1398 4975 1402
rect 5083 1398 5087 1402
rect 5107 1398 5111 1402
rect 5219 1398 5223 1402
rect 5243 1398 5247 1402
rect 5355 1398 5359 1402
rect 5379 1398 5383 1402
rect 5491 1398 5495 1402
rect 5515 1398 5519 1402
rect 5663 1398 5667 1402
rect 111 1318 115 1322
rect 159 1318 163 1322
rect 423 1318 427 1322
rect 455 1318 459 1322
rect 711 1318 715 1322
rect 775 1318 779 1322
rect 999 1318 1003 1322
rect 1095 1318 1099 1322
rect 1287 1318 1291 1322
rect 1423 1318 1427 1322
rect 1935 1318 1939 1322
rect 1975 1318 1979 1322
rect 2131 1318 2135 1322
rect 2139 1318 2143 1322
rect 2267 1318 2271 1322
rect 2275 1318 2279 1322
rect 2403 1318 2407 1322
rect 2411 1318 2415 1322
rect 2547 1318 2551 1322
rect 2555 1318 2559 1322
rect 2683 1318 2687 1322
rect 2715 1318 2719 1322
rect 2819 1318 2823 1322
rect 2891 1318 2895 1322
rect 2955 1318 2959 1322
rect 3075 1318 3079 1322
rect 3091 1318 3095 1322
rect 3227 1318 3231 1322
rect 3267 1318 3271 1322
rect 3467 1318 3471 1322
rect 3651 1318 3655 1322
rect 3799 1318 3803 1322
rect 3839 1282 3843 1286
rect 4735 1282 4739 1286
rect 4839 1282 4843 1286
rect 4879 1282 4883 1286
rect 4975 1282 4979 1286
rect 5031 1282 5035 1286
rect 5111 1282 5115 1286
rect 5191 1282 5195 1286
rect 5247 1282 5251 1286
rect 5359 1282 5363 1286
rect 5383 1282 5387 1286
rect 5519 1282 5523 1286
rect 5527 1282 5531 1286
rect 5663 1282 5667 1286
rect 1975 1206 1979 1210
rect 2023 1206 2027 1210
rect 2159 1206 2163 1210
rect 2239 1206 2243 1210
rect 2295 1206 2299 1210
rect 2431 1206 2435 1210
rect 2479 1206 2483 1210
rect 2583 1206 2587 1210
rect 2719 1206 2723 1210
rect 2743 1206 2747 1210
rect 2919 1206 2923 1210
rect 2959 1206 2963 1210
rect 3103 1206 3107 1210
rect 3207 1206 3211 1210
rect 3295 1206 3299 1210
rect 3455 1206 3459 1210
rect 3495 1206 3499 1210
rect 3679 1206 3683 1210
rect 3799 1206 3803 1210
rect 111 1182 115 1186
rect 131 1182 135 1186
rect 331 1182 335 1186
rect 427 1182 431 1186
rect 563 1182 567 1186
rect 747 1182 751 1186
rect 803 1182 807 1186
rect 1043 1182 1047 1186
rect 1067 1182 1071 1186
rect 1283 1182 1287 1186
rect 1395 1182 1399 1186
rect 1523 1182 1527 1186
rect 1771 1182 1775 1186
rect 1935 1182 1939 1186
rect 3839 1162 3843 1166
rect 3859 1162 3863 1166
rect 4067 1162 4071 1166
rect 4299 1162 4303 1166
rect 4539 1162 4543 1166
rect 4707 1162 4711 1166
rect 4779 1162 4783 1166
rect 4851 1162 4855 1166
rect 5003 1162 5007 1166
rect 5027 1162 5031 1166
rect 5163 1162 5167 1166
rect 5283 1162 5287 1166
rect 5331 1162 5335 1166
rect 5499 1162 5503 1166
rect 5515 1162 5519 1166
rect 5663 1162 5667 1166
rect 111 1070 115 1074
rect 159 1070 163 1074
rect 263 1070 267 1074
rect 359 1070 363 1074
rect 439 1070 443 1074
rect 591 1070 595 1074
rect 615 1070 619 1074
rect 783 1070 787 1074
rect 831 1070 835 1074
rect 951 1070 955 1074
rect 1071 1070 1075 1074
rect 1111 1070 1115 1074
rect 1271 1070 1275 1074
rect 1311 1070 1315 1074
rect 1431 1070 1435 1074
rect 1551 1070 1555 1074
rect 1591 1070 1595 1074
rect 1751 1070 1755 1074
rect 1799 1070 1803 1074
rect 1935 1070 1939 1074
rect 1975 1070 1979 1074
rect 1995 1070 1999 1074
rect 2211 1070 2215 1074
rect 2451 1070 2455 1074
rect 2691 1070 2695 1074
rect 2931 1070 2935 1074
rect 3091 1070 3095 1074
rect 3179 1070 3183 1074
rect 3243 1070 3247 1074
rect 3395 1070 3399 1074
rect 3427 1070 3431 1074
rect 3651 1070 3655 1074
rect 3799 1070 3803 1074
rect 3839 1050 3843 1054
rect 3887 1050 3891 1054
rect 4071 1050 4075 1054
rect 4095 1050 4099 1054
rect 4279 1050 4283 1054
rect 4327 1050 4331 1054
rect 4511 1050 4515 1054
rect 4567 1050 4571 1054
rect 4759 1050 4763 1054
rect 4807 1050 4811 1054
rect 5023 1050 5027 1054
rect 5055 1050 5059 1054
rect 5295 1050 5299 1054
rect 5311 1050 5315 1054
rect 5543 1050 5547 1054
rect 5663 1050 5667 1054
rect 111 954 115 958
rect 227 954 231 958
rect 235 954 239 958
rect 379 954 383 958
rect 411 954 415 958
rect 539 954 543 958
rect 587 954 591 958
rect 715 954 719 958
rect 755 954 759 958
rect 891 954 895 958
rect 923 954 927 958
rect 1075 954 1079 958
rect 1083 954 1087 958
rect 1243 954 1247 958
rect 1259 954 1263 958
rect 1403 954 1407 958
rect 1443 954 1447 958
rect 1563 954 1567 958
rect 1627 954 1631 958
rect 1723 954 1727 958
rect 1787 954 1791 958
rect 1935 954 1939 958
rect 3839 938 3843 942
rect 3859 938 3863 942
rect 3971 938 3975 942
rect 4043 938 4047 942
rect 4179 938 4183 942
rect 4251 938 4255 942
rect 4403 938 4407 942
rect 4483 938 4487 942
rect 4643 938 4647 942
rect 4731 938 4735 942
rect 4899 938 4903 942
rect 4995 938 4999 942
rect 5171 938 5175 942
rect 5267 938 5271 942
rect 5443 938 5447 942
rect 5515 938 5519 942
rect 5663 938 5667 942
rect 1975 930 1979 934
rect 2047 930 2051 934
rect 2351 930 2355 934
rect 2647 930 2651 934
rect 2927 930 2931 934
rect 3119 930 3123 934
rect 3207 930 3211 934
rect 3271 930 3275 934
rect 3423 930 3427 934
rect 3495 930 3499 934
rect 3799 930 3803 934
rect 111 826 115 830
rect 255 826 259 830
rect 375 826 379 830
rect 407 826 411 830
rect 567 826 571 830
rect 655 826 659 830
rect 743 826 747 830
rect 919 826 923 830
rect 943 826 947 830
rect 1103 826 1107 830
rect 1239 826 1243 830
rect 1287 826 1291 830
rect 1471 826 1475 830
rect 1535 826 1539 830
rect 1655 826 1659 830
rect 1815 826 1819 830
rect 1935 826 1939 830
rect 3839 826 3843 830
rect 3887 826 3891 830
rect 3999 826 4003 830
rect 4047 826 4051 830
rect 4207 826 4211 830
rect 4279 826 4283 830
rect 4431 826 4435 830
rect 4559 826 4563 830
rect 4671 826 4675 830
rect 4879 826 4883 830
rect 4927 826 4931 830
rect 5199 826 5203 830
rect 5223 826 5227 830
rect 5471 826 5475 830
rect 5543 826 5547 830
rect 5663 826 5667 830
rect 1975 818 1979 822
rect 1995 818 1999 822
rect 2019 818 2023 822
rect 2251 818 2255 822
rect 2323 818 2327 822
rect 2523 818 2527 822
rect 2619 818 2623 822
rect 2771 818 2775 822
rect 2899 818 2903 822
rect 3003 818 3007 822
rect 3179 818 3183 822
rect 3227 818 3231 822
rect 3451 818 3455 822
rect 3467 818 3471 822
rect 3651 818 3655 822
rect 3799 818 3803 822
rect 111 714 115 718
rect 131 714 135 718
rect 307 714 311 718
rect 347 714 351 718
rect 499 714 503 718
rect 627 714 631 718
rect 683 714 687 718
rect 859 714 863 718
rect 915 714 919 718
rect 1027 714 1031 718
rect 1187 714 1191 718
rect 1211 714 1215 718
rect 1339 714 1343 718
rect 1491 714 1495 718
rect 1507 714 1511 718
rect 1651 714 1655 718
rect 1787 714 1791 718
rect 1935 714 1939 718
rect 111 602 115 606
rect 159 602 163 606
rect 335 602 339 606
rect 375 602 379 606
rect 527 602 531 606
rect 599 602 603 606
rect 711 602 715 606
rect 807 602 811 606
rect 887 602 891 606
rect 999 602 1003 606
rect 1055 602 1059 606
rect 1175 602 1179 606
rect 1215 602 1219 606
rect 1343 602 1347 606
rect 1367 602 1371 606
rect 1511 602 1515 606
rect 1519 602 1523 606
rect 1671 602 1675 606
rect 1679 602 1683 606
rect 1815 602 1819 606
rect 1935 602 1939 606
rect 3839 706 3843 710
rect 3859 706 3863 710
rect 3995 706 3999 710
rect 4019 706 4023 710
rect 4131 706 4135 710
rect 4251 706 4255 710
rect 4267 706 4271 710
rect 4403 706 4407 710
rect 4531 706 4535 710
rect 4571 706 4575 710
rect 4771 706 4775 710
rect 4851 706 4855 710
rect 4995 706 4999 710
rect 5195 706 5199 710
rect 5227 706 5231 710
rect 5459 706 5463 710
rect 5515 706 5519 710
rect 5663 706 5667 710
rect 3839 594 3843 598
rect 3887 594 3891 598
rect 4023 594 4027 598
rect 4159 594 4163 598
rect 4295 594 4299 598
rect 4431 594 4435 598
rect 4479 594 4483 598
rect 4599 594 4603 598
rect 4695 594 4699 598
rect 4799 594 4803 598
rect 4935 594 4939 598
rect 5023 594 5027 598
rect 5191 594 5195 598
rect 5255 594 5259 598
rect 5447 594 5451 598
rect 5487 594 5491 598
rect 5663 594 5667 598
rect 1975 574 1979 578
rect 2023 574 2027 578
rect 2279 574 2283 578
rect 2551 574 2555 578
rect 2799 574 2803 578
rect 3031 574 3035 578
rect 3255 574 3259 578
rect 3311 574 3315 578
rect 3447 574 3451 578
rect 3479 574 3483 578
rect 3583 574 3587 578
rect 3679 574 3683 578
rect 3799 574 3803 578
rect 111 490 115 494
rect 131 490 135 494
rect 347 490 351 494
rect 427 490 431 494
rect 571 490 575 494
rect 763 490 767 494
rect 779 490 783 494
rect 971 490 975 494
rect 1107 490 1111 494
rect 1147 490 1151 494
rect 1315 490 1319 494
rect 1459 490 1463 494
rect 1483 490 1487 494
rect 1643 490 1647 494
rect 1787 490 1791 494
rect 1935 490 1939 494
rect 3839 470 3843 474
rect 3859 470 3863 474
rect 3995 470 3999 474
rect 4131 470 4135 474
rect 4267 470 4271 474
rect 4451 470 4455 474
rect 4651 470 4655 474
rect 4667 470 4671 474
rect 4859 470 4863 474
rect 4907 470 4911 474
rect 5067 470 5071 474
rect 5163 470 5167 474
rect 5283 470 5287 474
rect 5419 470 5423 474
rect 5507 470 5511 474
rect 5663 470 5667 474
rect 1975 462 1979 466
rect 1995 462 1999 466
rect 2155 462 2159 466
rect 2347 462 2351 466
rect 2539 462 2543 466
rect 2731 462 2735 466
rect 2923 462 2927 466
rect 3115 462 3119 466
rect 3283 462 3287 466
rect 3299 462 3303 466
rect 3419 462 3423 466
rect 3483 462 3487 466
rect 3555 462 3559 466
rect 3651 462 3655 466
rect 3799 462 3803 466
rect 111 362 115 366
rect 159 362 163 366
rect 239 362 243 366
rect 391 362 395 366
rect 455 362 459 366
rect 551 362 555 366
rect 711 362 715 366
rect 791 362 795 366
rect 871 362 875 366
rect 1031 362 1035 366
rect 1135 362 1139 366
rect 1487 362 1491 366
rect 1815 362 1819 366
rect 1935 362 1939 366
rect 3839 354 3843 358
rect 4479 354 4483 358
rect 4679 354 4683 358
rect 4751 354 4755 358
rect 4887 354 4891 358
rect 4911 354 4915 358
rect 5071 354 5075 358
rect 5095 354 5099 358
rect 5231 354 5235 358
rect 5311 354 5315 358
rect 5399 354 5403 358
rect 5535 354 5539 358
rect 5543 354 5547 358
rect 5663 354 5667 358
rect 1975 326 1979 330
rect 2023 326 2027 330
rect 2047 326 2051 330
rect 2183 326 2187 330
rect 2319 326 2323 330
rect 2375 326 2379 330
rect 2455 326 2459 330
rect 2567 326 2571 330
rect 2591 326 2595 330
rect 2727 326 2731 330
rect 2759 326 2763 330
rect 2863 326 2867 330
rect 2951 326 2955 330
rect 2999 326 3003 330
rect 3135 326 3139 330
rect 3143 326 3147 330
rect 3271 326 3275 330
rect 3327 326 3331 330
rect 3407 326 3411 330
rect 3511 326 3515 330
rect 3543 326 3547 330
rect 3679 326 3683 330
rect 3799 326 3803 330
rect 111 218 115 222
rect 147 218 151 222
rect 211 218 215 222
rect 283 218 287 222
rect 363 218 367 222
rect 419 218 423 222
rect 523 218 527 222
rect 555 218 559 222
rect 683 218 687 222
rect 691 218 695 222
rect 827 218 831 222
rect 843 218 847 222
rect 963 218 967 222
rect 1003 218 1007 222
rect 1099 218 1103 222
rect 1935 218 1939 222
rect 1975 198 1979 202
rect 1995 198 1999 202
rect 2019 198 2023 202
rect 2131 198 2135 202
rect 2155 198 2159 202
rect 2267 198 2271 202
rect 2291 198 2295 202
rect 2403 198 2407 202
rect 2427 198 2431 202
rect 2539 198 2543 202
rect 2563 198 2567 202
rect 2675 198 2679 202
rect 2699 198 2703 202
rect 2811 198 2815 202
rect 2835 198 2839 202
rect 2947 198 2951 202
rect 2971 198 2975 202
rect 3083 198 3087 202
rect 3107 198 3111 202
rect 3219 198 3223 202
rect 3243 198 3247 202
rect 3355 198 3359 202
rect 3379 198 3383 202
rect 3491 198 3495 202
rect 3515 198 3519 202
rect 3627 198 3631 202
rect 3651 198 3655 202
rect 3799 198 3803 202
rect 3839 202 3843 206
rect 4291 202 4295 206
rect 4427 202 4431 206
rect 4563 202 4567 206
rect 4699 202 4703 206
rect 4723 202 4727 206
rect 4835 202 4839 206
rect 4883 202 4887 206
rect 4971 202 4975 206
rect 5043 202 5047 206
rect 5107 202 5111 206
rect 5203 202 5207 206
rect 5243 202 5247 206
rect 5371 202 5375 206
rect 5379 202 5383 206
rect 5515 202 5519 206
rect 5663 202 5667 206
rect 111 106 115 110
rect 175 106 179 110
rect 311 106 315 110
rect 447 106 451 110
rect 583 106 587 110
rect 719 106 723 110
rect 855 106 859 110
rect 991 106 995 110
rect 1127 106 1131 110
rect 1935 106 1939 110
rect 1975 86 1979 90
rect 2023 86 2027 90
rect 2159 86 2163 90
rect 2295 86 2299 90
rect 2431 86 2435 90
rect 2567 86 2571 90
rect 2703 86 2707 90
rect 2839 86 2843 90
rect 2975 86 2979 90
rect 3111 86 3115 90
rect 3247 86 3251 90
rect 3383 86 3387 90
rect 3519 86 3523 90
rect 3655 86 3659 90
rect 3799 86 3803 90
rect 3839 90 3843 94
rect 4319 90 4323 94
rect 4455 90 4459 94
rect 4591 90 4595 94
rect 4727 90 4731 94
rect 4863 90 4867 94
rect 4999 90 5003 94
rect 5135 90 5139 94
rect 5271 90 5275 94
rect 5407 90 5411 94
rect 5543 90 5547 94
rect 5663 90 5667 94
<< m4 >>
rect 96 5753 97 5759
rect 103 5758 1959 5759
rect 103 5754 111 5758
rect 115 5754 131 5758
rect 135 5754 267 5758
rect 271 5754 403 5758
rect 407 5754 1935 5758
rect 1939 5754 1959 5758
rect 103 5753 1959 5754
rect 1965 5753 1966 5759
rect 3822 5694 5714 5695
rect 3822 5691 3839 5694
rect 1958 5685 1959 5691
rect 1965 5690 3823 5691
rect 1965 5686 1975 5690
rect 1979 5686 1995 5690
rect 1999 5686 2171 5690
rect 2175 5686 2371 5690
rect 2375 5686 2563 5690
rect 2567 5686 2747 5690
rect 2751 5686 2931 5690
rect 2935 5686 3107 5690
rect 3111 5686 3275 5690
rect 3279 5686 3443 5690
rect 3447 5686 3619 5690
rect 3623 5686 3799 5690
rect 3803 5686 3823 5690
rect 1965 5685 3823 5686
rect 3829 5690 3839 5691
rect 3843 5690 4467 5694
rect 4471 5690 4603 5694
rect 4607 5690 4739 5694
rect 4743 5690 4875 5694
rect 4879 5690 5663 5694
rect 5667 5690 5714 5694
rect 3829 5689 5714 5690
rect 3829 5685 3830 5689
rect 84 5641 85 5647
rect 91 5646 1947 5647
rect 91 5642 111 5646
rect 115 5642 159 5646
rect 163 5642 295 5646
rect 299 5642 343 5646
rect 347 5642 431 5646
rect 435 5642 535 5646
rect 539 5642 735 5646
rect 739 5642 943 5646
rect 947 5642 1159 5646
rect 1163 5642 1383 5646
rect 1387 5642 1607 5646
rect 1611 5642 1815 5646
rect 1819 5642 1935 5646
rect 1939 5642 1947 5646
rect 91 5641 1947 5642
rect 1953 5641 1954 5647
rect 3810 5582 5702 5583
rect 3810 5579 3839 5582
rect 1946 5573 1947 5579
rect 1953 5578 3811 5579
rect 1953 5574 1975 5578
rect 1979 5574 2023 5578
rect 2027 5574 2199 5578
rect 2203 5574 2375 5578
rect 2379 5574 2399 5578
rect 2403 5574 2591 5578
rect 2595 5574 2607 5578
rect 2611 5574 2775 5578
rect 2779 5574 2831 5578
rect 2835 5574 2959 5578
rect 2963 5574 3047 5578
rect 3051 5574 3135 5578
rect 3139 5574 3263 5578
rect 3267 5574 3303 5578
rect 3307 5574 3471 5578
rect 3475 5574 3479 5578
rect 3483 5574 3647 5578
rect 3651 5574 3679 5578
rect 3683 5574 3799 5578
rect 3803 5574 3811 5578
rect 1953 5573 3811 5574
rect 3817 5578 3839 5579
rect 3843 5578 4431 5582
rect 4435 5578 4495 5582
rect 4499 5578 4567 5582
rect 4571 5578 4631 5582
rect 4635 5578 4703 5582
rect 4707 5578 4767 5582
rect 4771 5578 4839 5582
rect 4843 5578 4903 5582
rect 4907 5578 4975 5582
rect 4979 5578 5111 5582
rect 5115 5578 5663 5582
rect 5667 5578 5702 5582
rect 3817 5577 5702 5578
rect 3817 5573 3818 5577
rect 96 5529 97 5535
rect 103 5534 1959 5535
rect 103 5530 111 5534
rect 115 5530 315 5534
rect 319 5530 507 5534
rect 511 5530 707 5534
rect 711 5530 875 5534
rect 879 5530 915 5534
rect 919 5530 1011 5534
rect 1015 5530 1131 5534
rect 1135 5530 1147 5534
rect 1151 5530 1291 5534
rect 1295 5530 1355 5534
rect 1359 5530 1435 5534
rect 1439 5530 1579 5534
rect 1583 5530 1723 5534
rect 1727 5530 1787 5534
rect 1791 5530 1935 5534
rect 1939 5530 1959 5534
rect 103 5529 1959 5530
rect 1965 5529 1966 5535
rect 3822 5465 3823 5471
rect 3829 5470 5707 5471
rect 3829 5466 3839 5470
rect 3843 5466 4403 5470
rect 4407 5466 4427 5470
rect 4431 5466 4539 5470
rect 4543 5466 4587 5470
rect 4591 5466 4675 5470
rect 4679 5466 4747 5470
rect 4751 5466 4811 5470
rect 4815 5466 4907 5470
rect 4911 5466 4947 5470
rect 4951 5466 5075 5470
rect 5079 5466 5083 5470
rect 5087 5466 5663 5470
rect 5667 5466 5707 5470
rect 3829 5465 5707 5466
rect 5713 5465 5714 5471
rect 3822 5463 3830 5465
rect 1958 5457 1959 5463
rect 1965 5462 3823 5463
rect 1965 5458 1975 5462
rect 1979 5458 2347 5462
rect 2351 5458 2451 5462
rect 2455 5458 2579 5462
rect 2583 5458 2699 5462
rect 2703 5458 2803 5462
rect 2807 5458 2947 5462
rect 2951 5458 3019 5462
rect 3023 5458 3187 5462
rect 3191 5458 3235 5462
rect 3239 5458 3427 5462
rect 3431 5458 3451 5462
rect 3455 5458 3651 5462
rect 3655 5458 3799 5462
rect 3803 5458 3823 5462
rect 1965 5457 3823 5458
rect 3829 5457 3830 5463
rect 84 5417 85 5423
rect 91 5422 1947 5423
rect 91 5418 111 5422
rect 115 5418 719 5422
rect 723 5418 855 5422
rect 859 5418 903 5422
rect 907 5418 991 5422
rect 995 5418 1039 5422
rect 1043 5418 1127 5422
rect 1131 5418 1175 5422
rect 1179 5418 1263 5422
rect 1267 5418 1319 5422
rect 1323 5418 1399 5422
rect 1403 5418 1463 5422
rect 1467 5418 1535 5422
rect 1539 5418 1607 5422
rect 1611 5418 1671 5422
rect 1675 5418 1751 5422
rect 1755 5418 1807 5422
rect 1811 5418 1935 5422
rect 1939 5418 1947 5422
rect 91 5417 1947 5418
rect 1953 5417 1954 5423
rect 1946 5345 1947 5351
rect 1953 5350 3811 5351
rect 1953 5346 1975 5350
rect 1979 5346 2319 5350
rect 2323 5346 2479 5350
rect 2483 5346 2519 5350
rect 2523 5346 2719 5350
rect 2723 5346 2727 5350
rect 2731 5346 2919 5350
rect 2923 5346 2975 5350
rect 2979 5346 3119 5350
rect 3123 5346 3215 5350
rect 3219 5346 3327 5350
rect 3331 5346 3455 5350
rect 3459 5346 3535 5350
rect 3539 5346 3679 5350
rect 3683 5346 3799 5350
rect 3803 5346 3811 5350
rect 1953 5345 3811 5346
rect 3817 5350 5702 5351
rect 3817 5346 3839 5350
rect 3843 5346 4431 5350
rect 4435 5346 4455 5350
rect 4459 5346 4615 5350
rect 4619 5346 4775 5350
rect 4779 5346 4799 5350
rect 4803 5346 4935 5350
rect 4939 5346 4983 5350
rect 4987 5346 5103 5350
rect 5107 5346 5175 5350
rect 5179 5346 5663 5350
rect 5667 5346 5702 5350
rect 3817 5345 5702 5346
rect 96 5305 97 5311
rect 103 5310 1959 5311
rect 103 5306 111 5310
rect 115 5306 691 5310
rect 695 5306 723 5310
rect 727 5306 827 5310
rect 831 5306 875 5310
rect 879 5306 963 5310
rect 967 5306 1027 5310
rect 1031 5306 1099 5310
rect 1103 5306 1187 5310
rect 1191 5306 1235 5310
rect 1239 5306 1355 5310
rect 1359 5306 1371 5310
rect 1375 5306 1507 5310
rect 1511 5306 1523 5310
rect 1527 5306 1643 5310
rect 1647 5306 1779 5310
rect 1783 5306 1935 5310
rect 1939 5306 1959 5310
rect 103 5305 1959 5306
rect 1965 5305 1966 5311
rect 1958 5229 1959 5235
rect 1965 5234 3823 5235
rect 1965 5230 1975 5234
rect 1979 5230 2275 5234
rect 2279 5230 2291 5234
rect 2295 5230 2475 5234
rect 2479 5230 2491 5234
rect 2495 5230 2683 5234
rect 2687 5230 2691 5234
rect 2695 5230 2891 5234
rect 2895 5230 3091 5234
rect 3095 5230 3099 5234
rect 3103 5230 3299 5234
rect 3303 5230 3307 5234
rect 3311 5230 3507 5234
rect 3511 5230 3799 5234
rect 3803 5230 3823 5234
rect 1965 5229 3823 5230
rect 3829 5229 3830 5235
rect 3822 5217 3823 5223
rect 3829 5222 5707 5223
rect 3829 5218 3839 5222
rect 3843 5218 4403 5222
rect 4407 5218 4435 5222
rect 4439 5218 4587 5222
rect 4591 5218 4595 5222
rect 4599 5218 4755 5222
rect 4759 5218 4771 5222
rect 4775 5218 4915 5222
rect 4919 5218 4955 5222
rect 4959 5218 5067 5222
rect 5071 5218 5147 5222
rect 5151 5218 5219 5222
rect 5223 5218 5379 5222
rect 5383 5218 5515 5222
rect 5519 5218 5663 5222
rect 5667 5218 5707 5222
rect 3829 5217 5707 5218
rect 5713 5217 5714 5223
rect 84 5193 85 5199
rect 91 5198 1947 5199
rect 91 5194 111 5198
rect 115 5194 447 5198
rect 451 5194 623 5198
rect 627 5194 751 5198
rect 755 5194 807 5198
rect 811 5194 903 5198
rect 907 5194 999 5198
rect 1003 5194 1055 5198
rect 1059 5194 1199 5198
rect 1203 5194 1215 5198
rect 1219 5194 1383 5198
rect 1387 5194 1399 5198
rect 1403 5194 1551 5198
rect 1555 5194 1607 5198
rect 1611 5194 1815 5198
rect 1819 5194 1935 5198
rect 1939 5194 1947 5198
rect 91 5193 1947 5194
rect 1953 5193 1954 5199
rect 1946 5101 1947 5107
rect 1953 5106 3811 5107
rect 1953 5102 1975 5106
rect 1979 5102 2119 5106
rect 2123 5102 2303 5106
rect 2307 5102 2327 5106
rect 2331 5102 2503 5106
rect 2507 5102 2535 5106
rect 2539 5102 2711 5106
rect 2715 5102 2751 5106
rect 2755 5102 2919 5106
rect 2923 5102 2975 5106
rect 2979 5102 3127 5106
rect 3131 5102 3207 5106
rect 3211 5102 3335 5106
rect 3339 5102 3799 5106
rect 3803 5102 3811 5106
rect 1953 5101 3811 5102
rect 3817 5103 3818 5107
rect 3817 5102 5702 5103
rect 3817 5101 3839 5102
rect 3810 5098 3839 5101
rect 3843 5098 3887 5102
rect 3891 5098 4087 5102
rect 4091 5098 4327 5102
rect 4331 5098 4463 5102
rect 4467 5098 4567 5102
rect 4571 5098 4623 5102
rect 4627 5098 4783 5102
rect 4787 5098 4815 5102
rect 4819 5098 4943 5102
rect 4947 5098 5063 5102
rect 5067 5098 5095 5102
rect 5099 5098 5247 5102
rect 5251 5098 5311 5102
rect 5315 5098 5407 5102
rect 5411 5098 5543 5102
rect 5547 5098 5663 5102
rect 5667 5098 5702 5102
rect 3810 5097 5702 5098
rect 96 5073 97 5079
rect 103 5078 1959 5079
rect 103 5074 111 5078
rect 115 5074 155 5078
rect 159 5074 379 5078
rect 383 5074 419 5078
rect 423 5074 595 5078
rect 599 5074 627 5078
rect 631 5074 779 5078
rect 783 5074 899 5078
rect 903 5074 971 5078
rect 975 5074 1171 5078
rect 1175 5074 1195 5078
rect 1199 5074 1371 5078
rect 1375 5074 1499 5078
rect 1503 5074 1579 5078
rect 1583 5074 1787 5078
rect 1791 5074 1935 5078
rect 1939 5074 1959 5078
rect 103 5073 1959 5074
rect 1965 5073 1966 5079
rect 3822 4990 5714 4991
rect 3822 4987 3839 4990
rect 1958 4981 1959 4987
rect 1965 4986 3823 4987
rect 1965 4982 1975 4986
rect 1979 4982 1995 4986
rect 1999 4982 2091 4986
rect 2095 4982 2131 4986
rect 2135 4982 2267 4986
rect 2271 4982 2299 4986
rect 2303 4982 2419 4986
rect 2423 4982 2507 4986
rect 2511 4982 2619 4986
rect 2623 4982 2723 4986
rect 2727 4982 2859 4986
rect 2863 4982 2947 4986
rect 2951 4982 3123 4986
rect 3127 4982 3179 4986
rect 3183 4982 3395 4986
rect 3399 4982 3651 4986
rect 3655 4982 3799 4986
rect 3803 4982 3823 4986
rect 1965 4981 3823 4982
rect 3829 4986 3839 4987
rect 3843 4986 3859 4990
rect 3863 4986 3995 4990
rect 3999 4986 4059 4990
rect 4063 4986 4131 4990
rect 4135 4986 4267 4990
rect 4271 4986 4299 4990
rect 4303 4986 4403 4990
rect 4407 4986 4539 4990
rect 4543 4986 4675 4990
rect 4679 4986 4787 4990
rect 4791 4986 4811 4990
rect 4815 4986 4947 4990
rect 4951 4986 5035 4990
rect 5039 4986 5083 4990
rect 5087 4986 5227 4990
rect 5231 4986 5283 4990
rect 5287 4986 5379 4990
rect 5383 4986 5515 4990
rect 5519 4986 5663 4990
rect 5667 4986 5714 4990
rect 3829 4985 5714 4986
rect 3829 4981 3830 4985
rect 84 4933 85 4939
rect 91 4938 1947 4939
rect 91 4934 111 4938
rect 115 4934 159 4938
rect 163 4934 183 4938
rect 187 4934 295 4938
rect 299 4934 407 4938
rect 411 4934 431 4938
rect 435 4934 567 4938
rect 571 4934 655 4938
rect 659 4934 703 4938
rect 707 4934 927 4938
rect 931 4934 1223 4938
rect 1227 4934 1527 4938
rect 1531 4934 1815 4938
rect 1819 4934 1935 4938
rect 1939 4934 1947 4938
rect 91 4933 1947 4934
rect 1953 4933 1954 4939
rect 1946 4861 1947 4867
rect 1953 4866 3811 4867
rect 1953 4862 1975 4866
rect 1979 4862 2023 4866
rect 2027 4862 2159 4866
rect 2163 4862 2295 4866
rect 2299 4862 2327 4866
rect 2331 4862 2447 4866
rect 2451 4862 2559 4866
rect 2563 4862 2647 4866
rect 2651 4862 2823 4866
rect 2827 4862 2887 4866
rect 2891 4862 3103 4866
rect 3107 4862 3151 4866
rect 3155 4862 3399 4866
rect 3403 4862 3423 4866
rect 3427 4862 3679 4866
rect 3683 4862 3799 4866
rect 3803 4862 3811 4866
rect 1953 4861 3811 4862
rect 3817 4861 3818 4867
rect 96 4809 97 4815
rect 103 4814 1959 4815
rect 103 4810 111 4814
rect 115 4810 131 4814
rect 135 4810 267 4814
rect 271 4810 403 4814
rect 407 4810 539 4814
rect 543 4810 675 4814
rect 679 4810 1935 4814
rect 1939 4810 1959 4814
rect 103 4809 1959 4810
rect 1965 4809 1966 4815
rect 3810 4797 3811 4803
rect 3817 4802 5695 4803
rect 3817 4798 3839 4802
rect 3843 4798 3887 4802
rect 3891 4798 4023 4802
rect 4027 4798 4071 4802
rect 4075 4798 4159 4802
rect 4163 4798 4295 4802
rect 4299 4798 4431 4802
rect 4435 4798 4535 4802
rect 4539 4798 4567 4802
rect 4571 4798 4703 4802
rect 4707 4798 4783 4802
rect 4787 4798 4839 4802
rect 4843 4798 4975 4802
rect 4979 4798 5039 4802
rect 5043 4798 5111 4802
rect 5115 4798 5255 4802
rect 5259 4798 5303 4802
rect 5307 4798 5407 4802
rect 5411 4798 5543 4802
rect 5547 4798 5663 4802
rect 5667 4798 5695 4802
rect 3817 4797 5695 4798
rect 5701 4797 5702 4803
rect 1958 4737 1959 4743
rect 1965 4742 3823 4743
rect 1965 4738 1975 4742
rect 1979 4738 2019 4742
rect 2023 4738 2195 4742
rect 2199 4738 2299 4742
rect 2303 4738 2371 4742
rect 2375 4738 2531 4742
rect 2535 4738 2547 4742
rect 2551 4738 2723 4742
rect 2727 4738 2795 4742
rect 2799 4738 3075 4742
rect 3079 4738 3371 4742
rect 3375 4738 3651 4742
rect 3655 4738 3799 4742
rect 3803 4738 3823 4742
rect 1965 4737 3823 4738
rect 3829 4737 3830 4743
rect 84 4693 85 4699
rect 91 4698 1947 4699
rect 91 4694 111 4698
rect 115 4694 159 4698
rect 163 4694 295 4698
rect 299 4694 431 4698
rect 435 4694 567 4698
rect 571 4694 703 4698
rect 707 4694 1935 4698
rect 1939 4694 1947 4698
rect 91 4693 1947 4694
rect 1953 4693 1954 4699
rect 3822 4685 3823 4691
rect 3829 4690 5707 4691
rect 3829 4686 3839 4690
rect 3843 4686 3859 4690
rect 3863 4686 3995 4690
rect 3999 4686 4043 4690
rect 4047 4686 4131 4690
rect 4135 4686 4267 4690
rect 4271 4686 4403 4690
rect 4407 4686 4507 4690
rect 4511 4686 4539 4690
rect 4543 4686 4675 4690
rect 4679 4686 4755 4690
rect 4759 4686 4819 4690
rect 4823 4686 4963 4690
rect 4967 4686 5011 4690
rect 5015 4686 5107 4690
rect 5111 4686 5243 4690
rect 5247 4686 5275 4690
rect 5279 4686 5379 4690
rect 5383 4686 5515 4690
rect 5519 4686 5663 4690
rect 5667 4686 5707 4690
rect 3829 4685 5707 4686
rect 5713 4685 5714 4691
rect 1946 4621 1947 4627
rect 1953 4626 3811 4627
rect 1953 4622 1975 4626
rect 1979 4622 2023 4626
rect 2027 4622 2047 4626
rect 2051 4622 2223 4626
rect 2227 4622 2263 4626
rect 2267 4622 2399 4626
rect 2403 4622 2527 4626
rect 2531 4622 2575 4626
rect 2579 4622 2751 4626
rect 2755 4622 2775 4626
rect 2779 4622 3015 4626
rect 3019 4622 3247 4626
rect 3251 4622 3471 4626
rect 3475 4622 3679 4626
rect 3683 4622 3799 4626
rect 3803 4622 3811 4626
rect 1953 4621 3811 4622
rect 3817 4621 3818 4627
rect 96 4569 97 4575
rect 103 4574 1959 4575
rect 103 4570 111 4574
rect 115 4570 131 4574
rect 135 4570 251 4574
rect 255 4570 267 4574
rect 271 4570 403 4574
rect 407 4570 443 4574
rect 447 4570 539 4574
rect 543 4570 651 4574
rect 655 4570 675 4574
rect 679 4570 875 4574
rect 879 4570 1099 4574
rect 1103 4570 1331 4574
rect 1335 4570 1571 4574
rect 1575 4570 1787 4574
rect 1791 4570 1935 4574
rect 1939 4570 1959 4574
rect 103 4569 1959 4570
rect 1965 4569 1966 4575
rect 3810 4573 3811 4579
rect 3817 4578 5695 4579
rect 3817 4574 3839 4578
rect 3843 4574 3887 4578
rect 3891 4574 4023 4578
rect 4027 4574 4159 4578
rect 4163 4574 4295 4578
rect 4299 4574 4431 4578
rect 4435 4574 4567 4578
rect 4571 4574 4671 4578
rect 4675 4574 4703 4578
rect 4707 4574 4807 4578
rect 4811 4574 4847 4578
rect 4851 4574 4943 4578
rect 4947 4574 4991 4578
rect 4995 4574 5079 4578
rect 5083 4574 5135 4578
rect 5139 4574 5271 4578
rect 5275 4574 5407 4578
rect 5411 4574 5543 4578
rect 5547 4574 5663 4578
rect 5667 4574 5695 4578
rect 3817 4573 5695 4574
rect 5701 4573 5702 4579
rect 1958 4497 1959 4503
rect 1965 4502 3823 4503
rect 1965 4498 1975 4502
rect 1979 4498 1995 4502
rect 1999 4498 2235 4502
rect 2239 4498 2267 4502
rect 2271 4498 2499 4502
rect 2503 4498 2515 4502
rect 2519 4498 2747 4502
rect 2751 4498 2971 4502
rect 2975 4498 2987 4502
rect 2991 4498 3187 4502
rect 3191 4498 3219 4502
rect 3223 4498 3395 4502
rect 3399 4498 3443 4502
rect 3447 4498 3611 4502
rect 3615 4498 3651 4502
rect 3655 4498 3799 4502
rect 3803 4498 3823 4502
rect 1965 4497 3823 4498
rect 3829 4497 3830 4503
rect 84 4457 85 4463
rect 91 4462 1947 4463
rect 91 4458 111 4462
rect 115 4458 279 4462
rect 283 4458 471 4462
rect 475 4458 511 4462
rect 515 4458 679 4462
rect 683 4458 687 4462
rect 691 4458 871 4462
rect 875 4458 903 4462
rect 907 4458 1071 4462
rect 1075 4458 1127 4462
rect 1131 4458 1279 4462
rect 1283 4458 1359 4462
rect 1363 4458 1495 4462
rect 1499 4458 1599 4462
rect 1603 4458 1719 4462
rect 1723 4458 1815 4462
rect 1819 4458 1935 4462
rect 1939 4458 1947 4462
rect 91 4457 1947 4458
rect 1953 4457 1954 4463
rect 3822 4457 3823 4463
rect 3829 4462 5707 4463
rect 3829 4458 3839 4462
rect 3843 4458 4347 4462
rect 4351 4458 4483 4462
rect 4487 4458 4619 4462
rect 4623 4458 4643 4462
rect 4647 4458 4755 4462
rect 4759 4458 4779 4462
rect 4783 4458 4891 4462
rect 4895 4458 4915 4462
rect 4919 4458 5051 4462
rect 5055 4458 5663 4462
rect 5667 4458 5707 4462
rect 3829 4457 5707 4458
rect 5713 4457 5714 4463
rect 1946 4373 1947 4379
rect 1953 4378 3811 4379
rect 1953 4374 1975 4378
rect 1979 4374 2023 4378
rect 2027 4374 2199 4378
rect 2203 4374 2295 4378
rect 2299 4374 2399 4378
rect 2403 4374 2543 4378
rect 2547 4374 2591 4378
rect 2595 4374 2775 4378
rect 2779 4374 2951 4378
rect 2955 4374 2999 4378
rect 3003 4374 3135 4378
rect 3139 4374 3215 4378
rect 3219 4374 3319 4378
rect 3323 4374 3423 4378
rect 3427 4374 3639 4378
rect 3643 4374 3799 4378
rect 3803 4374 3811 4378
rect 1953 4373 3811 4374
rect 3817 4373 3818 4379
rect 96 4341 97 4347
rect 103 4346 1959 4347
rect 103 4342 111 4346
rect 115 4342 483 4346
rect 487 4342 659 4346
rect 663 4342 715 4346
rect 719 4342 843 4346
rect 847 4342 851 4346
rect 855 4342 987 4346
rect 991 4342 1043 4346
rect 1047 4342 1123 4346
rect 1127 4342 1251 4346
rect 1255 4342 1259 4346
rect 1263 4342 1395 4346
rect 1399 4342 1467 4346
rect 1471 4342 1531 4346
rect 1535 4342 1667 4346
rect 1671 4342 1691 4346
rect 1695 4342 1935 4346
rect 1939 4342 1959 4346
rect 103 4341 1959 4342
rect 1965 4341 1966 4347
rect 3810 4329 3811 4335
rect 3817 4334 5695 4335
rect 3817 4330 3839 4334
rect 3843 4330 4135 4334
rect 4139 4330 4271 4334
rect 4275 4330 4375 4334
rect 4379 4330 4407 4334
rect 4411 4330 4511 4334
rect 4515 4330 4543 4334
rect 4547 4330 4647 4334
rect 4651 4330 4679 4334
rect 4683 4330 4783 4334
rect 4787 4330 4919 4334
rect 4923 4330 5663 4334
rect 5667 4330 5695 4334
rect 3817 4329 5695 4330
rect 5701 4329 5702 4335
rect 1958 4257 1959 4263
rect 1965 4262 3823 4263
rect 1965 4258 1975 4262
rect 1979 4258 1995 4262
rect 1999 4258 2171 4262
rect 2175 4258 2243 4262
rect 2247 4258 2371 4262
rect 2375 4258 2507 4262
rect 2511 4258 2563 4262
rect 2567 4258 2747 4262
rect 2751 4258 2763 4262
rect 2767 4258 2923 4262
rect 2927 4258 3019 4262
rect 3023 4258 3107 4262
rect 3111 4258 3283 4262
rect 3287 4258 3291 4262
rect 3295 4258 3799 4262
rect 3803 4258 3823 4262
rect 1965 4257 3823 4258
rect 3829 4257 3830 4263
rect 84 4221 85 4227
rect 91 4226 1947 4227
rect 91 4222 111 4226
rect 115 4222 727 4226
rect 731 4222 743 4226
rect 747 4222 863 4226
rect 867 4222 879 4226
rect 883 4222 999 4226
rect 1003 4222 1015 4226
rect 1019 4222 1135 4226
rect 1139 4222 1151 4226
rect 1155 4222 1271 4226
rect 1275 4222 1287 4226
rect 1291 4222 1407 4226
rect 1411 4222 1423 4226
rect 1427 4222 1543 4226
rect 1547 4222 1559 4226
rect 1563 4222 1679 4226
rect 1683 4222 1695 4226
rect 1699 4222 1815 4226
rect 1819 4222 1935 4226
rect 1939 4222 1947 4226
rect 91 4221 1947 4222
rect 1953 4221 1954 4227
rect 3822 4205 3823 4211
rect 3829 4210 5707 4211
rect 3829 4206 3839 4210
rect 3843 4206 3971 4210
rect 3975 4206 4107 4210
rect 4111 4206 4243 4210
rect 4247 4206 4379 4210
rect 4383 4206 4515 4210
rect 4519 4206 4651 4210
rect 4655 4206 5663 4210
rect 5667 4206 5707 4210
rect 3829 4205 5707 4206
rect 5713 4205 5714 4211
rect 1946 4133 1947 4139
rect 1953 4138 3811 4139
rect 1953 4134 1975 4138
rect 1979 4134 2023 4138
rect 2027 4134 2271 4138
rect 2275 4134 2535 4138
rect 2539 4134 2791 4138
rect 2795 4134 3047 4138
rect 3051 4134 3135 4138
rect 3139 4134 3271 4138
rect 3275 4134 3311 4138
rect 3315 4134 3407 4138
rect 3411 4134 3543 4138
rect 3547 4134 3679 4138
rect 3683 4134 3799 4138
rect 3803 4134 3811 4138
rect 1953 4133 3811 4134
rect 3817 4133 3818 4139
rect 96 4109 97 4115
rect 103 4114 1959 4115
rect 103 4110 111 4114
rect 115 4110 563 4114
rect 567 4110 699 4114
rect 703 4110 835 4114
rect 839 4110 971 4114
rect 975 4110 1107 4114
rect 1111 4110 1243 4114
rect 1247 4110 1379 4114
rect 1383 4110 1515 4114
rect 1519 4110 1651 4114
rect 1655 4110 1787 4114
rect 1791 4110 1935 4114
rect 1939 4110 1959 4114
rect 103 4109 1959 4110
rect 1965 4109 1966 4115
rect 3810 4069 3811 4075
rect 3817 4074 5695 4075
rect 3817 4070 3839 4074
rect 3843 4070 3887 4074
rect 3891 4070 3999 4074
rect 4003 4070 4023 4074
rect 4027 4070 4135 4074
rect 4139 4070 4159 4074
rect 4163 4070 4271 4074
rect 4275 4070 4295 4074
rect 4299 4070 4407 4074
rect 4411 4070 4431 4074
rect 4435 4070 4543 4074
rect 4547 4070 4567 4074
rect 4571 4070 4703 4074
rect 4707 4070 4839 4074
rect 4843 4070 5663 4074
rect 5667 4070 5695 4074
rect 3817 4069 5695 4070
rect 5701 4069 5702 4075
rect 84 3997 85 4003
rect 91 4002 1947 4003
rect 91 3998 111 4002
rect 115 3998 159 4002
rect 163 3998 327 4002
rect 331 3998 535 4002
rect 539 3998 591 4002
rect 595 3998 727 4002
rect 731 3998 751 4002
rect 755 3998 863 4002
rect 867 3998 967 4002
rect 971 3998 999 4002
rect 1003 3998 1135 4002
rect 1139 3998 1183 4002
rect 1187 3998 1271 4002
rect 1275 3998 1399 4002
rect 1403 3998 1407 4002
rect 1411 3998 1543 4002
rect 1547 3998 1615 4002
rect 1619 3998 1679 4002
rect 1683 3998 1815 4002
rect 1819 3998 1935 4002
rect 1939 3998 1947 4002
rect 91 3997 1947 3998
rect 1953 3997 1954 4003
rect 3822 3957 3823 3963
rect 3829 3962 5707 3963
rect 3829 3958 3839 3962
rect 3843 3958 3859 3962
rect 3863 3958 3995 3962
rect 3999 3958 4131 3962
rect 4135 3958 4147 3962
rect 4151 3958 4267 3962
rect 4271 3958 4299 3962
rect 4303 3958 4403 3962
rect 4407 3958 4459 3962
rect 4463 3958 4539 3962
rect 4543 3958 4619 3962
rect 4623 3958 4675 3962
rect 4679 3958 4779 3962
rect 4783 3958 4811 3962
rect 4815 3958 5663 3962
rect 5667 3958 5707 3962
rect 3829 3957 5707 3958
rect 5713 3957 5714 3963
rect 1958 3929 1959 3935
rect 1965 3934 3823 3935
rect 1965 3930 1975 3934
rect 1979 3930 1995 3934
rect 1999 3930 2403 3934
rect 2407 3930 2827 3934
rect 2831 3930 3107 3934
rect 3111 3930 3243 3934
rect 3247 3930 3251 3934
rect 3255 3930 3379 3934
rect 3383 3930 3515 3934
rect 3519 3930 3651 3934
rect 3655 3930 3799 3934
rect 3803 3930 3823 3934
rect 1965 3929 3823 3930
rect 3829 3929 3830 3935
rect 96 3885 97 3891
rect 103 3890 1959 3891
rect 103 3886 111 3890
rect 115 3886 131 3890
rect 135 3886 299 3890
rect 303 3886 355 3890
rect 359 3886 507 3890
rect 511 3886 619 3890
rect 623 3886 723 3890
rect 727 3886 899 3890
rect 903 3886 939 3890
rect 943 3886 1155 3890
rect 1159 3886 1195 3890
rect 1199 3886 1371 3890
rect 1375 3886 1499 3890
rect 1503 3886 1587 3890
rect 1591 3886 1787 3890
rect 1791 3886 1935 3890
rect 1939 3886 1959 3890
rect 103 3885 1959 3886
rect 1965 3885 1966 3891
rect 1946 3817 1947 3823
rect 1953 3822 3811 3823
rect 1953 3818 1975 3822
rect 1979 3818 2023 3822
rect 2027 3818 2175 3822
rect 2179 3818 2351 3822
rect 2355 3818 2431 3822
rect 2435 3818 2535 3822
rect 2539 3818 2719 3822
rect 2723 3818 2855 3822
rect 2859 3818 2895 3822
rect 2899 3818 3071 3822
rect 3075 3818 3247 3822
rect 3251 3818 3279 3822
rect 3283 3818 3423 3822
rect 3427 3818 3607 3822
rect 3611 3818 3679 3822
rect 3683 3818 3799 3822
rect 3803 3818 3811 3822
rect 1953 3817 3811 3818
rect 3817 3822 5702 3823
rect 3817 3818 3839 3822
rect 3843 3818 3887 3822
rect 3891 3818 4023 3822
rect 4027 3818 4175 3822
rect 4179 3818 4327 3822
rect 4331 3818 4487 3822
rect 4491 3818 4503 3822
rect 4507 3818 4639 3822
rect 4643 3818 4647 3822
rect 4651 3818 4775 3822
rect 4779 3818 4807 3822
rect 4811 3818 4911 3822
rect 4915 3818 5047 3822
rect 5051 3818 5663 3822
rect 5667 3818 5702 3822
rect 3817 3817 5702 3818
rect 84 3761 85 3767
rect 91 3766 1947 3767
rect 91 3762 111 3766
rect 115 3762 159 3766
rect 163 3762 247 3766
rect 251 3762 383 3766
rect 387 3762 519 3766
rect 523 3762 647 3766
rect 651 3762 791 3766
rect 795 3762 927 3766
rect 931 3762 1063 3766
rect 1067 3762 1223 3766
rect 1227 3762 1343 3766
rect 1347 3762 1527 3766
rect 1531 3762 1815 3766
rect 1819 3762 1935 3766
rect 1939 3762 1947 3766
rect 91 3761 1947 3762
rect 1953 3761 1954 3767
rect 1958 3697 1959 3703
rect 1965 3702 3823 3703
rect 1965 3698 1975 3702
rect 1979 3698 1995 3702
rect 1999 3698 2011 3702
rect 2015 3698 2147 3702
rect 2151 3698 2291 3702
rect 2295 3698 2323 3702
rect 2327 3698 2435 3702
rect 2439 3698 2507 3702
rect 2511 3698 2579 3702
rect 2583 3698 2691 3702
rect 2695 3698 2723 3702
rect 2727 3698 2867 3702
rect 2871 3698 3011 3702
rect 3015 3698 3043 3702
rect 3047 3698 3155 3702
rect 3159 3698 3219 3702
rect 3223 3698 3299 3702
rect 3303 3698 3395 3702
rect 3399 3698 3579 3702
rect 3583 3698 3799 3702
rect 3803 3698 3823 3702
rect 1965 3697 3823 3698
rect 3829 3697 3830 3703
rect 3822 3685 3823 3691
rect 3829 3690 5707 3691
rect 3829 3686 3839 3690
rect 3843 3686 4019 3690
rect 4023 3686 4155 3690
rect 4159 3686 4291 3690
rect 4295 3686 4427 3690
rect 4431 3686 4475 3690
rect 4479 3686 4563 3690
rect 4567 3686 4611 3690
rect 4615 3686 4699 3690
rect 4703 3686 4747 3690
rect 4751 3686 4835 3690
rect 4839 3686 4883 3690
rect 4887 3686 4971 3690
rect 4975 3686 5019 3690
rect 5023 3686 5107 3690
rect 5111 3686 5243 3690
rect 5247 3686 5379 3690
rect 5383 3686 5515 3690
rect 5519 3686 5663 3690
rect 5667 3686 5707 3690
rect 3829 3685 5707 3686
rect 5713 3685 5714 3691
rect 96 3633 97 3639
rect 103 3638 1959 3639
rect 103 3634 111 3638
rect 115 3634 219 3638
rect 223 3634 491 3638
rect 495 3634 635 3638
rect 639 3634 763 3638
rect 767 3634 779 3638
rect 783 3634 923 3638
rect 927 3634 1035 3638
rect 1039 3634 1067 3638
rect 1071 3634 1211 3638
rect 1215 3634 1315 3638
rect 1319 3634 1935 3638
rect 1939 3634 1959 3638
rect 103 3633 1959 3634
rect 1965 3633 1966 3639
rect 1946 3577 1947 3583
rect 1953 3582 3811 3583
rect 1953 3578 1975 3582
rect 1979 3578 2039 3582
rect 2043 3578 2175 3582
rect 2179 3578 2239 3582
rect 2243 3578 2319 3582
rect 2323 3578 2375 3582
rect 2379 3578 2463 3582
rect 2467 3578 2511 3582
rect 2515 3578 2607 3582
rect 2611 3578 2647 3582
rect 2651 3578 2751 3582
rect 2755 3578 2783 3582
rect 2787 3578 2895 3582
rect 2899 3578 2919 3582
rect 2923 3578 3039 3582
rect 3043 3578 3055 3582
rect 3059 3578 3183 3582
rect 3187 3578 3191 3582
rect 3195 3578 3327 3582
rect 3331 3578 3463 3582
rect 3467 3578 3799 3582
rect 3803 3578 3811 3582
rect 1953 3577 3811 3578
rect 3817 3577 3818 3583
rect 3810 3525 3811 3531
rect 3817 3530 5695 3531
rect 3817 3526 3839 3530
rect 3843 3526 4047 3530
rect 4051 3526 4183 3530
rect 4187 3526 4319 3530
rect 4323 3526 4455 3530
rect 4459 3526 4591 3530
rect 4595 3526 4727 3530
rect 4731 3526 4863 3530
rect 4867 3526 4999 3530
rect 5003 3526 5135 3530
rect 5139 3526 5271 3530
rect 5275 3526 5407 3530
rect 5411 3526 5543 3530
rect 5547 3526 5663 3530
rect 5667 3526 5695 3530
rect 3817 3525 5695 3526
rect 5701 3525 5702 3531
rect 84 3501 85 3507
rect 91 3506 1947 3507
rect 91 3502 111 3506
rect 115 3502 431 3506
rect 435 3502 519 3506
rect 523 3502 567 3506
rect 571 3502 663 3506
rect 667 3502 703 3506
rect 707 3502 807 3506
rect 811 3502 839 3506
rect 843 3502 951 3506
rect 955 3502 975 3506
rect 979 3502 1095 3506
rect 1099 3502 1239 3506
rect 1243 3502 1935 3506
rect 1939 3502 1947 3506
rect 91 3501 1947 3502
rect 1953 3501 1954 3507
rect 1958 3461 1959 3467
rect 1965 3466 3823 3467
rect 1965 3462 1975 3466
rect 1979 3462 2171 3466
rect 2175 3462 2211 3466
rect 2215 3462 2347 3466
rect 2351 3462 2483 3466
rect 2487 3462 2531 3466
rect 2535 3462 2619 3466
rect 2623 3462 2715 3466
rect 2719 3462 2755 3466
rect 2759 3462 2891 3466
rect 2895 3462 2907 3466
rect 2911 3462 3027 3466
rect 3031 3462 3099 3466
rect 3103 3462 3163 3466
rect 3167 3462 3291 3466
rect 3295 3462 3299 3466
rect 3303 3462 3435 3466
rect 3439 3462 3483 3466
rect 3487 3462 3651 3466
rect 3655 3462 3799 3466
rect 3803 3462 3823 3466
rect 1965 3461 3823 3462
rect 3829 3461 3830 3467
rect 3822 3405 3823 3411
rect 3829 3410 5707 3411
rect 3829 3406 3839 3410
rect 3843 3406 3859 3410
rect 3863 3406 4099 3410
rect 4103 3406 4347 3410
rect 4351 3406 4587 3410
rect 4591 3406 4811 3410
rect 4815 3406 5027 3410
rect 5031 3406 5235 3410
rect 5239 3406 5379 3410
rect 5383 3406 5451 3410
rect 5455 3406 5515 3410
rect 5519 3406 5663 3410
rect 5667 3406 5707 3410
rect 3829 3405 5707 3406
rect 5713 3405 5714 3411
rect 96 3381 97 3387
rect 103 3386 1959 3387
rect 103 3382 111 3386
rect 115 3382 323 3386
rect 327 3382 403 3386
rect 407 3382 459 3386
rect 463 3382 539 3386
rect 543 3382 595 3386
rect 599 3382 675 3386
rect 679 3382 731 3386
rect 735 3382 811 3386
rect 815 3382 867 3386
rect 871 3382 947 3386
rect 951 3382 1935 3386
rect 1939 3382 1959 3386
rect 103 3381 1959 3382
rect 1965 3381 1966 3387
rect 1946 3325 1947 3331
rect 1953 3330 3811 3331
rect 1953 3326 1975 3330
rect 1979 3326 2151 3330
rect 2155 3326 2199 3330
rect 2203 3326 2375 3330
rect 2379 3326 2399 3330
rect 2403 3326 2559 3330
rect 2563 3326 2687 3330
rect 2691 3326 2743 3330
rect 2747 3326 2935 3330
rect 2939 3326 3015 3330
rect 3019 3326 3127 3330
rect 3131 3326 3319 3330
rect 3323 3326 3359 3330
rect 3363 3326 3511 3330
rect 3515 3326 3679 3330
rect 3683 3326 3799 3330
rect 3803 3326 3811 3330
rect 1953 3325 3811 3326
rect 3817 3325 3818 3331
rect 3810 3293 3811 3299
rect 3817 3298 5695 3299
rect 3817 3294 3839 3298
rect 3843 3294 3887 3298
rect 3891 3294 4127 3298
rect 4131 3294 4375 3298
rect 4379 3294 4607 3298
rect 4611 3294 4615 3298
rect 4619 3294 4815 3298
rect 4819 3294 4839 3298
rect 4843 3294 5015 3298
rect 5019 3294 5055 3298
rect 5059 3294 5199 3298
rect 5203 3294 5263 3298
rect 5267 3294 5383 3298
rect 5387 3294 5479 3298
rect 5483 3294 5543 3298
rect 5547 3294 5663 3298
rect 5667 3294 5695 3298
rect 3817 3293 5695 3294
rect 5701 3293 5702 3299
rect 84 3261 85 3267
rect 91 3266 1947 3267
rect 91 3262 111 3266
rect 115 3262 159 3266
rect 163 3262 335 3266
rect 339 3262 351 3266
rect 355 3262 487 3266
rect 491 3262 543 3266
rect 547 3262 623 3266
rect 627 3262 751 3266
rect 755 3262 759 3266
rect 763 3262 895 3266
rect 899 3262 959 3266
rect 963 3262 1935 3266
rect 1939 3262 1947 3266
rect 91 3261 1947 3262
rect 1953 3261 1954 3267
rect 1958 3213 1959 3219
rect 1965 3218 3823 3219
rect 1965 3214 1975 3218
rect 1979 3214 1995 3218
rect 1999 3214 2123 3218
rect 2127 3214 2147 3218
rect 2151 3214 2347 3218
rect 2351 3214 2371 3218
rect 2375 3214 2555 3218
rect 2559 3214 2659 3218
rect 2663 3214 2771 3218
rect 2775 3214 2987 3218
rect 2991 3214 3211 3218
rect 3215 3214 3331 3218
rect 3335 3214 3443 3218
rect 3447 3214 3651 3218
rect 3655 3214 3799 3218
rect 3803 3214 3823 3218
rect 1965 3213 3823 3214
rect 3829 3213 3830 3219
rect 3822 3165 3823 3171
rect 3829 3170 5707 3171
rect 3829 3166 3839 3170
rect 3843 3166 3859 3170
rect 3863 3166 4099 3170
rect 4103 3166 4347 3170
rect 4351 3166 4467 3170
rect 4471 3166 4579 3170
rect 4583 3166 4651 3170
rect 4655 3166 4787 3170
rect 4791 3166 4859 3170
rect 4863 3166 4987 3170
rect 4991 3166 5075 3170
rect 5079 3166 5171 3170
rect 5175 3166 5307 3170
rect 5311 3166 5355 3170
rect 5359 3166 5515 3170
rect 5519 3166 5663 3170
rect 5667 3166 5707 3170
rect 3829 3165 5707 3166
rect 5713 3165 5714 3171
rect 96 3133 97 3139
rect 103 3138 1959 3139
rect 103 3134 111 3138
rect 115 3134 131 3138
rect 135 3134 307 3138
rect 311 3134 371 3138
rect 375 3134 515 3138
rect 519 3134 627 3138
rect 631 3134 723 3138
rect 727 3134 875 3138
rect 879 3134 931 3138
rect 935 3134 1115 3138
rect 1119 3134 1347 3138
rect 1351 3134 1579 3138
rect 1583 3134 1787 3138
rect 1791 3134 1935 3138
rect 1939 3134 1959 3138
rect 103 3133 1959 3134
rect 1965 3133 1966 3139
rect 1946 3101 1947 3107
rect 1953 3106 3811 3107
rect 1953 3102 1975 3106
rect 1979 3102 2023 3106
rect 2027 3102 2175 3106
rect 2179 3102 2375 3106
rect 2379 3102 2583 3106
rect 2587 3102 2647 3106
rect 2651 3102 2783 3106
rect 2787 3102 2799 3106
rect 2803 3102 2927 3106
rect 2931 3102 3015 3106
rect 3019 3102 3079 3106
rect 3083 3102 3239 3106
rect 3243 3102 3399 3106
rect 3403 3102 3471 3106
rect 3475 3102 3567 3106
rect 3571 3102 3679 3106
rect 3683 3102 3799 3106
rect 3803 3102 3811 3106
rect 1953 3101 3811 3102
rect 3817 3101 3818 3107
rect 3810 3053 3811 3059
rect 3817 3058 5695 3059
rect 3817 3054 3839 3058
rect 3843 3054 4255 3058
rect 4259 3054 4455 3058
rect 4459 3054 4495 3058
rect 4499 3054 4671 3058
rect 4675 3054 4679 3058
rect 4683 3054 4887 3058
rect 4891 3054 4911 3058
rect 4915 3054 5103 3058
rect 5107 3054 5167 3058
rect 5171 3054 5335 3058
rect 5339 3054 5423 3058
rect 5427 3054 5543 3058
rect 5547 3054 5663 3058
rect 5667 3054 5695 3058
rect 3817 3053 5695 3054
rect 5701 3053 5702 3059
rect 84 3021 85 3027
rect 91 3026 1947 3027
rect 91 3022 111 3026
rect 115 3022 159 3026
rect 163 3022 175 3026
rect 179 3022 399 3026
rect 403 3022 407 3026
rect 411 3022 623 3026
rect 627 3022 655 3026
rect 659 3022 823 3026
rect 827 3022 903 3026
rect 907 3022 1007 3026
rect 1011 3022 1143 3026
rect 1147 3022 1183 3026
rect 1187 3022 1351 3026
rect 1355 3022 1375 3026
rect 1379 3022 1511 3026
rect 1515 3022 1607 3026
rect 1611 3022 1671 3026
rect 1675 3022 1815 3026
rect 1819 3022 1935 3026
rect 1939 3022 1947 3026
rect 91 3021 1947 3022
rect 1953 3021 1954 3027
rect 1958 2989 1959 2995
rect 1965 2994 3823 2995
rect 1965 2990 1975 2994
rect 1979 2990 2619 2994
rect 2623 2990 2755 2994
rect 2759 2990 2803 2994
rect 2807 2990 2899 2994
rect 2903 2990 2939 2994
rect 2943 2990 3051 2994
rect 3055 2990 3075 2994
rect 3079 2990 3211 2994
rect 3215 2990 3347 2994
rect 3351 2990 3371 2994
rect 3375 2990 3483 2994
rect 3487 2990 3539 2994
rect 3543 2990 3799 2994
rect 3803 2990 3823 2994
rect 1965 2989 3823 2990
rect 3829 2989 3830 2995
rect 3822 2917 3823 2923
rect 3829 2922 5707 2923
rect 3829 2918 3839 2922
rect 3843 2918 3995 2922
rect 3999 2918 4211 2922
rect 4215 2918 4227 2922
rect 4231 2918 4427 2922
rect 4431 2918 4443 2922
rect 4447 2918 4643 2922
rect 4647 2918 4699 2922
rect 4703 2918 4883 2922
rect 4887 2918 4971 2922
rect 4975 2918 5139 2922
rect 5143 2918 5251 2922
rect 5255 2918 5395 2922
rect 5399 2918 5515 2922
rect 5519 2918 5663 2922
rect 5667 2918 5707 2922
rect 3829 2917 5707 2918
rect 5713 2917 5714 2923
rect 96 2905 97 2911
rect 103 2910 1959 2911
rect 103 2906 111 2910
rect 115 2906 147 2910
rect 151 2906 379 2910
rect 383 2906 395 2910
rect 399 2906 595 2910
rect 599 2906 787 2910
rect 791 2906 795 2910
rect 799 2906 971 2910
rect 975 2906 979 2910
rect 983 2906 1147 2910
rect 1151 2906 1155 2910
rect 1159 2906 1315 2910
rect 1319 2906 1323 2910
rect 1327 2906 1483 2910
rect 1487 2906 1643 2910
rect 1647 2906 1787 2910
rect 1791 2906 1935 2910
rect 1939 2906 1959 2910
rect 103 2905 1959 2906
rect 1965 2905 1966 2911
rect 1946 2825 1947 2831
rect 1953 2830 3811 2831
rect 1953 2826 1975 2830
rect 1979 2826 2023 2830
rect 2027 2826 2167 2830
rect 2171 2826 2335 2830
rect 2339 2826 2495 2830
rect 2499 2826 2663 2830
rect 2667 2826 2831 2830
rect 2835 2826 2967 2830
rect 2971 2826 2999 2830
rect 3003 2826 3103 2830
rect 3107 2826 3167 2830
rect 3171 2826 3239 2830
rect 3243 2826 3375 2830
rect 3379 2826 3511 2830
rect 3515 2826 3799 2830
rect 3803 2826 3811 2830
rect 1953 2825 3811 2826
rect 3817 2825 3818 2831
rect 3810 2801 3811 2807
rect 3817 2806 5695 2807
rect 3817 2802 3839 2806
rect 3843 2802 3919 2806
rect 3923 2802 4023 2806
rect 4027 2802 4055 2806
rect 4059 2802 4191 2806
rect 4195 2802 4239 2806
rect 4243 2802 4327 2806
rect 4331 2802 4463 2806
rect 4467 2802 4471 2806
rect 4475 2802 4727 2806
rect 4731 2802 4999 2806
rect 5003 2802 5279 2806
rect 5283 2802 5543 2806
rect 5547 2802 5663 2806
rect 5667 2802 5695 2806
rect 3817 2801 5695 2802
rect 5701 2801 5702 2807
rect 84 2781 85 2787
rect 91 2786 1947 2787
rect 91 2782 111 2786
rect 115 2782 423 2786
rect 427 2782 623 2786
rect 627 2782 655 2786
rect 659 2782 815 2786
rect 819 2782 975 2786
rect 979 2782 999 2786
rect 1003 2782 1143 2786
rect 1147 2782 1175 2786
rect 1179 2782 1311 2786
rect 1315 2782 1343 2786
rect 1347 2782 1479 2786
rect 1483 2782 1511 2786
rect 1515 2782 1671 2786
rect 1675 2782 1815 2786
rect 1819 2782 1935 2786
rect 1939 2782 1947 2786
rect 91 2781 1947 2782
rect 1953 2781 1954 2787
rect 1958 2713 1959 2719
rect 1965 2718 3823 2719
rect 1965 2714 1975 2718
rect 1979 2714 1995 2718
rect 1999 2714 2139 2718
rect 2143 2714 2307 2718
rect 2311 2714 2379 2718
rect 2383 2714 2467 2718
rect 2471 2714 2515 2718
rect 2519 2714 2635 2718
rect 2639 2714 2659 2718
rect 2663 2714 2803 2718
rect 2807 2714 2947 2718
rect 2951 2714 2971 2718
rect 2975 2714 3091 2718
rect 3095 2714 3139 2718
rect 3143 2714 3235 2718
rect 3239 2714 3799 2718
rect 3803 2714 3823 2718
rect 1965 2713 3823 2714
rect 3829 2713 3830 2719
rect 3822 2677 3823 2683
rect 3829 2682 5707 2683
rect 3829 2678 3839 2682
rect 3843 2678 3891 2682
rect 3895 2678 4027 2682
rect 4031 2678 4099 2682
rect 4103 2678 4163 2682
rect 4167 2678 4299 2682
rect 4303 2678 4435 2682
rect 4439 2678 4515 2682
rect 4519 2678 4755 2682
rect 4759 2678 5011 2682
rect 5015 2678 5275 2682
rect 5279 2678 5515 2682
rect 5519 2678 5663 2682
rect 5667 2678 5707 2682
rect 3829 2677 5707 2678
rect 5713 2677 5714 2683
rect 96 2669 97 2675
rect 103 2674 1959 2675
rect 103 2670 111 2674
rect 115 2670 627 2674
rect 631 2670 771 2674
rect 775 2670 787 2674
rect 791 2670 907 2674
rect 911 2670 947 2674
rect 951 2670 1043 2674
rect 1047 2670 1115 2674
rect 1119 2670 1179 2674
rect 1183 2670 1283 2674
rect 1287 2670 1315 2674
rect 1319 2670 1451 2674
rect 1455 2670 1587 2674
rect 1591 2670 1723 2674
rect 1727 2670 1935 2674
rect 1939 2670 1959 2674
rect 103 2669 1959 2670
rect 1965 2669 1966 2675
rect 1946 2597 1947 2603
rect 1953 2602 3811 2603
rect 1953 2598 1975 2602
rect 1979 2598 2407 2602
rect 2411 2598 2511 2602
rect 2515 2598 2543 2602
rect 2547 2598 2647 2602
rect 2651 2598 2687 2602
rect 2691 2598 2783 2602
rect 2787 2598 2831 2602
rect 2835 2598 2919 2602
rect 2923 2598 2975 2602
rect 2979 2598 3055 2602
rect 3059 2598 3119 2602
rect 3123 2598 3191 2602
rect 3195 2598 3263 2602
rect 3267 2598 3327 2602
rect 3331 2598 3463 2602
rect 3467 2598 3799 2602
rect 3803 2598 3811 2602
rect 1953 2597 3811 2598
rect 3817 2597 3818 2603
rect 3810 2561 3811 2567
rect 3817 2566 5695 2567
rect 3817 2562 3839 2566
rect 3843 2562 4127 2566
rect 4131 2562 4327 2566
rect 4331 2562 4495 2566
rect 4499 2562 4543 2566
rect 4547 2562 4631 2566
rect 4635 2562 4767 2566
rect 4771 2562 4783 2566
rect 4787 2562 4903 2566
rect 4907 2562 5039 2566
rect 5043 2562 5303 2566
rect 5307 2562 5543 2566
rect 5547 2562 5663 2566
rect 5667 2562 5695 2566
rect 3817 2561 5695 2562
rect 5701 2561 5702 2567
rect 84 2541 85 2547
rect 91 2546 1947 2547
rect 91 2542 111 2546
rect 115 2542 551 2546
rect 555 2542 687 2546
rect 691 2542 799 2546
rect 803 2542 831 2546
rect 835 2542 935 2546
rect 939 2542 983 2546
rect 987 2542 1071 2546
rect 1075 2542 1135 2546
rect 1139 2542 1207 2546
rect 1211 2542 1295 2546
rect 1299 2542 1343 2546
rect 1347 2542 1455 2546
rect 1459 2542 1479 2546
rect 1483 2542 1615 2546
rect 1619 2542 1751 2546
rect 1755 2542 1783 2546
rect 1787 2542 1935 2546
rect 1939 2542 1947 2546
rect 91 2541 1947 2542
rect 1953 2541 1954 2547
rect 1958 2469 1959 2475
rect 1965 2474 3823 2475
rect 1965 2470 1975 2474
rect 1979 2470 2307 2474
rect 2311 2470 2483 2474
rect 2487 2470 2515 2474
rect 2519 2470 2619 2474
rect 2623 2470 2715 2474
rect 2719 2470 2755 2474
rect 2759 2470 2891 2474
rect 2895 2470 2907 2474
rect 2911 2470 3027 2474
rect 3031 2470 3099 2474
rect 3103 2470 3163 2474
rect 3167 2470 3283 2474
rect 3287 2470 3299 2474
rect 3303 2470 3435 2474
rect 3439 2470 3467 2474
rect 3471 2470 3651 2474
rect 3655 2470 3799 2474
rect 3803 2470 3823 2474
rect 1965 2469 3823 2470
rect 3829 2469 3830 2475
rect 3822 2433 3823 2439
rect 3829 2438 5707 2439
rect 3829 2434 3839 2438
rect 3843 2434 4467 2438
rect 4471 2434 4603 2438
rect 4607 2434 4699 2438
rect 4703 2434 4739 2438
rect 4743 2434 4835 2438
rect 4839 2434 4875 2438
rect 4879 2434 4971 2438
rect 4975 2434 5011 2438
rect 5015 2434 5107 2438
rect 5111 2434 5243 2438
rect 5247 2434 5379 2438
rect 5383 2434 5515 2438
rect 5519 2434 5663 2438
rect 5667 2434 5707 2438
rect 3829 2433 5707 2434
rect 5713 2433 5714 2439
rect 96 2417 97 2423
rect 103 2422 1959 2423
rect 103 2418 111 2422
rect 115 2418 131 2422
rect 135 2418 339 2422
rect 343 2418 523 2422
rect 527 2418 563 2422
rect 567 2418 659 2422
rect 663 2418 803 2422
rect 807 2418 955 2422
rect 959 2418 1043 2422
rect 1047 2418 1107 2422
rect 1111 2418 1267 2422
rect 1271 2418 1291 2422
rect 1295 2418 1427 2422
rect 1431 2418 1547 2422
rect 1551 2418 1587 2422
rect 1591 2418 1755 2422
rect 1759 2418 1787 2422
rect 1791 2418 1935 2422
rect 1939 2418 1959 2422
rect 103 2417 1959 2418
rect 1965 2417 1966 2423
rect 1946 2349 1947 2355
rect 1953 2354 3811 2355
rect 1953 2350 1975 2354
rect 1979 2350 2223 2354
rect 2227 2350 2335 2354
rect 2339 2350 2503 2354
rect 2507 2350 2543 2354
rect 2547 2350 2743 2354
rect 2747 2350 2767 2354
rect 2771 2350 2935 2354
rect 2939 2350 3007 2354
rect 3011 2350 3127 2354
rect 3131 2350 3239 2354
rect 3243 2350 3311 2354
rect 3315 2350 3471 2354
rect 3475 2350 3495 2354
rect 3499 2350 3679 2354
rect 3683 2350 3799 2354
rect 3803 2350 3811 2354
rect 1953 2349 3811 2350
rect 3817 2349 3818 2355
rect 3810 2309 3811 2315
rect 3817 2314 5695 2315
rect 3817 2310 3839 2314
rect 3843 2310 3887 2314
rect 3891 2310 4183 2314
rect 4187 2310 4495 2314
rect 4499 2310 4727 2314
rect 4731 2310 4791 2314
rect 4795 2310 4863 2314
rect 4867 2310 4999 2314
rect 5003 2310 5087 2314
rect 5091 2310 5135 2314
rect 5139 2310 5271 2314
rect 5275 2310 5383 2314
rect 5387 2310 5407 2314
rect 5411 2310 5543 2314
rect 5547 2310 5663 2314
rect 5667 2310 5695 2314
rect 3817 2309 5695 2310
rect 5701 2309 5702 2315
rect 84 2301 85 2307
rect 91 2306 1947 2307
rect 91 2302 111 2306
rect 115 2302 159 2306
rect 163 2302 319 2306
rect 323 2302 367 2306
rect 371 2302 551 2306
rect 555 2302 591 2306
rect 595 2302 831 2306
rect 835 2302 1071 2306
rect 1075 2302 1151 2306
rect 1155 2302 1319 2306
rect 1323 2302 1495 2306
rect 1499 2302 1575 2306
rect 1579 2302 1815 2306
rect 1819 2302 1935 2306
rect 1939 2302 1947 2306
rect 91 2301 1947 2302
rect 1953 2301 1954 2307
rect 1958 2237 1959 2243
rect 1965 2242 3823 2243
rect 1965 2238 1975 2242
rect 1979 2238 1995 2242
rect 1999 2238 2155 2242
rect 2159 2238 2195 2242
rect 2199 2238 2387 2242
rect 2391 2238 2475 2242
rect 2479 2238 2667 2242
rect 2671 2238 2739 2242
rect 2743 2238 2979 2242
rect 2983 2238 2987 2242
rect 2991 2238 3211 2242
rect 3215 2238 3331 2242
rect 3335 2238 3443 2242
rect 3447 2238 3651 2242
rect 3655 2238 3799 2242
rect 3803 2238 3823 2242
rect 1965 2237 3823 2238
rect 3829 2237 3830 2243
rect 3822 2193 3823 2199
rect 3829 2198 5707 2199
rect 3829 2194 3839 2198
rect 3843 2194 3859 2198
rect 3863 2194 3995 2198
rect 3999 2194 4131 2198
rect 4135 2194 4155 2198
rect 4159 2194 4267 2198
rect 4271 2194 4403 2198
rect 4407 2194 4467 2198
rect 4471 2194 4539 2198
rect 4543 2194 4699 2198
rect 4703 2194 4763 2198
rect 4767 2194 4891 2198
rect 4895 2194 5059 2198
rect 5063 2194 5099 2198
rect 5103 2194 5315 2198
rect 5319 2194 5355 2198
rect 5359 2194 5515 2198
rect 5519 2194 5663 2198
rect 5667 2194 5707 2198
rect 3829 2193 5707 2194
rect 5713 2193 5714 2199
rect 96 2165 97 2171
rect 103 2170 1959 2171
rect 103 2166 111 2170
rect 115 2166 131 2170
rect 135 2166 291 2170
rect 295 2166 483 2170
rect 487 2166 523 2170
rect 527 2166 691 2170
rect 695 2166 803 2170
rect 807 2166 915 2170
rect 919 2166 1123 2170
rect 1127 2166 1147 2170
rect 1151 2166 1387 2170
rect 1391 2166 1467 2170
rect 1471 2166 1635 2170
rect 1639 2166 1787 2170
rect 1791 2166 1935 2170
rect 1939 2166 1959 2170
rect 103 2165 1959 2166
rect 1965 2165 1966 2171
rect 3810 2061 3811 2067
rect 3817 2066 5695 2067
rect 3817 2062 3839 2066
rect 3843 2062 3887 2066
rect 3891 2062 4023 2066
rect 4027 2062 4159 2066
rect 4163 2062 4295 2066
rect 4299 2062 4431 2066
rect 4435 2062 4567 2066
rect 4571 2062 4719 2066
rect 4723 2062 4727 2066
rect 4731 2062 4895 2066
rect 4899 2062 4919 2066
rect 4923 2062 5087 2066
rect 5091 2062 5127 2066
rect 5131 2062 5279 2066
rect 5283 2062 5343 2066
rect 5347 2062 5479 2066
rect 5483 2062 5543 2066
rect 5547 2062 5663 2066
rect 5667 2062 5695 2066
rect 3817 2061 5695 2062
rect 5701 2061 5702 2067
rect 84 2049 85 2055
rect 91 2054 1947 2055
rect 91 2050 111 2054
rect 115 2050 263 2054
rect 267 2050 319 2054
rect 323 2050 399 2054
rect 403 2050 511 2054
rect 515 2050 535 2054
rect 539 2050 679 2054
rect 683 2050 719 2054
rect 723 2050 823 2054
rect 827 2050 943 2054
rect 947 2050 967 2054
rect 971 2050 1111 2054
rect 1115 2050 1175 2054
rect 1179 2050 1255 2054
rect 1259 2050 1399 2054
rect 1403 2050 1415 2054
rect 1419 2050 1543 2054
rect 1547 2050 1663 2054
rect 1667 2050 1679 2054
rect 1683 2050 1815 2054
rect 1819 2050 1935 2054
rect 1939 2050 1947 2054
rect 91 2049 1947 2050
rect 1953 2049 1954 2055
rect 3822 1949 3823 1955
rect 3829 1954 5707 1955
rect 3829 1950 3839 1954
rect 3843 1950 3859 1954
rect 3863 1950 3995 1954
rect 3999 1950 4043 1954
rect 4047 1950 4131 1954
rect 4135 1950 4267 1954
rect 4271 1950 4283 1954
rect 4287 1950 4403 1954
rect 4407 1950 4539 1954
rect 4543 1950 4563 1954
rect 4567 1950 4691 1954
rect 4695 1950 4867 1954
rect 4871 1950 4875 1954
rect 4879 1950 5059 1954
rect 5063 1950 5203 1954
rect 5207 1950 5251 1954
rect 5255 1950 5451 1954
rect 5455 1950 5515 1954
rect 5519 1950 5663 1954
rect 5667 1950 5707 1954
rect 3829 1949 5707 1950
rect 5713 1949 5714 1955
rect 1946 1935 1947 1941
rect 1953 1935 1978 1941
rect 1972 1931 1978 1935
rect 96 1925 97 1931
rect 103 1930 1959 1931
rect 103 1926 111 1930
rect 115 1926 235 1930
rect 239 1926 371 1930
rect 375 1926 435 1930
rect 439 1926 507 1930
rect 511 1926 627 1930
rect 631 1926 651 1930
rect 655 1926 795 1930
rect 799 1926 811 1930
rect 815 1926 939 1930
rect 943 1926 987 1930
rect 991 1926 1083 1930
rect 1087 1926 1155 1930
rect 1159 1926 1227 1930
rect 1231 1926 1323 1930
rect 1327 1926 1371 1930
rect 1375 1926 1483 1930
rect 1487 1926 1515 1930
rect 1519 1926 1643 1930
rect 1647 1926 1651 1930
rect 1655 1926 1787 1930
rect 1791 1926 1935 1930
rect 1939 1926 1959 1930
rect 103 1925 1959 1926
rect 1965 1925 1966 1931
rect 1972 1930 3811 1931
rect 1972 1926 1975 1930
rect 1979 1926 2023 1930
rect 2027 1926 2183 1930
rect 2187 1926 2415 1930
rect 2419 1926 2695 1930
rect 2699 1926 3015 1930
rect 3019 1926 3135 1930
rect 3139 1926 3271 1930
rect 3275 1926 3359 1930
rect 3363 1926 3407 1930
rect 3411 1926 3543 1930
rect 3547 1926 3679 1930
rect 3683 1926 3799 1930
rect 3803 1926 3811 1930
rect 1972 1925 3811 1926
rect 3817 1925 3818 1931
rect 3810 1837 3811 1843
rect 3817 1842 5695 1843
rect 3817 1838 3839 1842
rect 3843 1838 3887 1842
rect 3891 1838 4071 1842
rect 4075 1838 4311 1842
rect 4315 1838 4407 1842
rect 4411 1838 4543 1842
rect 4547 1838 4591 1842
rect 4595 1838 4679 1842
rect 4683 1838 4815 1842
rect 4819 1838 4903 1842
rect 4907 1838 4951 1842
rect 4955 1838 5231 1842
rect 5235 1838 5543 1842
rect 5547 1838 5663 1842
rect 5667 1838 5695 1842
rect 3817 1837 5695 1838
rect 5701 1837 5702 1843
rect 84 1801 85 1807
rect 91 1806 1947 1807
rect 91 1802 111 1806
rect 115 1802 223 1806
rect 227 1802 263 1806
rect 267 1802 463 1806
rect 467 1802 655 1806
rect 659 1802 695 1806
rect 699 1802 839 1806
rect 843 1802 927 1806
rect 931 1802 1015 1806
rect 1019 1802 1159 1806
rect 1163 1802 1183 1806
rect 1187 1802 1351 1806
rect 1355 1802 1391 1806
rect 1395 1802 1511 1806
rect 1515 1802 1671 1806
rect 1675 1802 1815 1806
rect 1819 1802 1935 1806
rect 1939 1802 1947 1806
rect 91 1801 1947 1802
rect 1953 1801 1954 1807
rect 1958 1801 1959 1807
rect 1965 1806 3823 1807
rect 1965 1802 1975 1806
rect 1979 1802 1995 1806
rect 1999 1802 2131 1806
rect 2135 1802 2267 1806
rect 2271 1802 2419 1806
rect 2423 1802 2579 1806
rect 2583 1802 2739 1806
rect 2743 1802 2899 1806
rect 2903 1802 3051 1806
rect 3055 1802 3107 1806
rect 3111 1802 3203 1806
rect 3207 1802 3243 1806
rect 3247 1802 3355 1806
rect 3359 1802 3379 1806
rect 3383 1802 3515 1806
rect 3519 1802 3651 1806
rect 3655 1802 3799 1806
rect 3803 1802 3823 1806
rect 1965 1801 3823 1802
rect 3829 1801 3830 1807
rect 3822 1709 3823 1715
rect 3829 1714 5707 1715
rect 3829 1710 3839 1714
rect 3843 1710 4379 1714
rect 4383 1710 4515 1714
rect 4519 1710 4563 1714
rect 4567 1710 4651 1714
rect 4655 1710 4699 1714
rect 4703 1710 4787 1714
rect 4791 1710 4835 1714
rect 4839 1710 4923 1714
rect 4927 1710 4971 1714
rect 4975 1710 5107 1714
rect 5111 1710 5243 1714
rect 5247 1710 5379 1714
rect 5383 1710 5515 1714
rect 5519 1710 5663 1714
rect 5667 1710 5707 1714
rect 3829 1709 5707 1710
rect 5713 1709 5714 1715
rect 1946 1687 1947 1693
rect 1953 1687 1978 1693
rect 1972 1683 1978 1687
rect 96 1677 97 1683
rect 103 1682 1959 1683
rect 103 1678 111 1682
rect 115 1678 131 1682
rect 135 1678 195 1682
rect 199 1678 363 1682
rect 367 1678 435 1682
rect 439 1678 619 1682
rect 623 1678 667 1682
rect 671 1678 875 1682
rect 879 1678 899 1682
rect 903 1678 1131 1682
rect 1135 1678 1139 1682
rect 1143 1678 1363 1682
rect 1367 1678 1935 1682
rect 1939 1678 1959 1682
rect 103 1677 1959 1678
rect 1965 1677 1966 1683
rect 1972 1682 3811 1683
rect 1972 1678 1975 1682
rect 1979 1678 2023 1682
rect 2027 1678 2159 1682
rect 2163 1678 2167 1682
rect 2171 1678 2295 1682
rect 2299 1678 2319 1682
rect 2323 1678 2447 1682
rect 2451 1678 2479 1682
rect 2483 1678 2607 1682
rect 2611 1678 2639 1682
rect 2643 1678 2767 1682
rect 2771 1678 2791 1682
rect 2795 1678 2927 1682
rect 2931 1678 2943 1682
rect 2947 1678 3079 1682
rect 3083 1678 3103 1682
rect 3107 1678 3231 1682
rect 3235 1678 3263 1682
rect 3267 1678 3383 1682
rect 3387 1678 3423 1682
rect 3427 1678 3543 1682
rect 3547 1678 3679 1682
rect 3683 1678 3799 1682
rect 3803 1678 3811 1682
rect 1972 1677 3811 1678
rect 3817 1677 3818 1683
rect 3810 1581 3811 1587
rect 3817 1586 5695 1587
rect 3817 1582 3839 1586
rect 3843 1582 4591 1586
rect 4595 1582 4727 1586
rect 4731 1582 4863 1586
rect 4867 1582 4999 1586
rect 5003 1582 5135 1586
rect 5139 1582 5271 1586
rect 5275 1582 5407 1586
rect 5411 1582 5543 1586
rect 5547 1582 5663 1586
rect 5667 1582 5695 1586
rect 3817 1581 5695 1582
rect 5701 1581 5702 1587
rect 84 1553 85 1559
rect 91 1558 1947 1559
rect 91 1554 111 1558
rect 115 1554 159 1558
rect 163 1554 327 1558
rect 331 1554 391 1558
rect 395 1554 511 1558
rect 515 1554 647 1558
rect 651 1554 695 1558
rect 699 1554 887 1558
rect 891 1554 903 1558
rect 907 1554 1079 1558
rect 1083 1554 1167 1558
rect 1171 1554 1935 1558
rect 1939 1554 1947 1558
rect 91 1553 1947 1554
rect 1953 1553 1954 1559
rect 1958 1553 1959 1559
rect 1965 1558 3823 1559
rect 1965 1554 1975 1558
rect 1979 1554 1995 1558
rect 1999 1554 2131 1558
rect 2135 1554 2139 1558
rect 2143 1554 2267 1558
rect 2271 1554 2291 1558
rect 2295 1554 2403 1558
rect 2407 1554 2451 1558
rect 2455 1554 2539 1558
rect 2543 1554 2611 1558
rect 2615 1554 2675 1558
rect 2679 1554 2763 1558
rect 2767 1554 2811 1558
rect 2815 1554 2915 1558
rect 2919 1554 2947 1558
rect 2951 1554 3075 1558
rect 3079 1554 3083 1558
rect 3087 1554 3219 1558
rect 3223 1554 3235 1558
rect 3239 1554 3355 1558
rect 3359 1554 3395 1558
rect 3399 1554 3491 1558
rect 3495 1554 3799 1558
rect 3803 1554 3823 1558
rect 1965 1553 3823 1554
rect 3829 1553 3830 1559
rect 1946 1439 1947 1445
rect 1953 1439 1978 1445
rect 1972 1435 1978 1439
rect 96 1429 97 1435
rect 103 1434 1959 1435
rect 103 1430 111 1434
rect 115 1430 131 1434
rect 135 1430 299 1434
rect 303 1430 395 1434
rect 399 1430 483 1434
rect 487 1430 667 1434
rect 671 1430 683 1434
rect 687 1430 859 1434
rect 863 1430 971 1434
rect 975 1430 1051 1434
rect 1055 1430 1259 1434
rect 1263 1430 1935 1434
rect 1939 1430 1959 1434
rect 103 1429 1959 1430
rect 1965 1429 1966 1435
rect 1972 1434 3811 1435
rect 1972 1430 1975 1434
rect 1979 1430 2023 1434
rect 2027 1430 2159 1434
rect 2163 1430 2167 1434
rect 2171 1430 2295 1434
rect 2299 1430 2303 1434
rect 2307 1430 2431 1434
rect 2435 1430 2439 1434
rect 2443 1430 2567 1434
rect 2571 1430 2575 1434
rect 2579 1430 2703 1434
rect 2707 1430 2711 1434
rect 2715 1430 2839 1434
rect 2843 1430 2847 1434
rect 2851 1430 2975 1434
rect 2979 1430 2983 1434
rect 2987 1430 3111 1434
rect 3115 1430 3119 1434
rect 3123 1430 3247 1434
rect 3251 1430 3255 1434
rect 3259 1430 3383 1434
rect 3387 1430 3519 1434
rect 3523 1430 3799 1434
rect 3803 1430 3811 1434
rect 1972 1429 3811 1430
rect 3817 1429 3818 1435
rect 3822 1397 3823 1403
rect 3829 1402 5707 1403
rect 3829 1398 3839 1402
rect 3843 1398 4563 1402
rect 4567 1398 4699 1402
rect 4703 1398 4811 1402
rect 4815 1398 4835 1402
rect 4839 1398 4947 1402
rect 4951 1398 4971 1402
rect 4975 1398 5083 1402
rect 5087 1398 5107 1402
rect 5111 1398 5219 1402
rect 5223 1398 5243 1402
rect 5247 1398 5355 1402
rect 5359 1398 5379 1402
rect 5383 1398 5491 1402
rect 5495 1398 5515 1402
rect 5519 1398 5663 1402
rect 5667 1398 5707 1402
rect 3829 1397 5707 1398
rect 5713 1397 5714 1403
rect 84 1317 85 1323
rect 91 1322 1947 1323
rect 91 1318 111 1322
rect 115 1318 159 1322
rect 163 1318 423 1322
rect 427 1318 455 1322
rect 459 1318 711 1322
rect 715 1318 775 1322
rect 779 1318 999 1322
rect 1003 1318 1095 1322
rect 1099 1318 1287 1322
rect 1291 1318 1423 1322
rect 1427 1318 1935 1322
rect 1939 1318 1947 1322
rect 91 1317 1947 1318
rect 1953 1317 1954 1323
rect 1958 1317 1959 1323
rect 1965 1322 3823 1323
rect 1965 1318 1975 1322
rect 1979 1318 2131 1322
rect 2135 1318 2139 1322
rect 2143 1318 2267 1322
rect 2271 1318 2275 1322
rect 2279 1318 2403 1322
rect 2407 1318 2411 1322
rect 2415 1318 2547 1322
rect 2551 1318 2555 1322
rect 2559 1318 2683 1322
rect 2687 1318 2715 1322
rect 2719 1318 2819 1322
rect 2823 1318 2891 1322
rect 2895 1318 2955 1322
rect 2959 1318 3075 1322
rect 3079 1318 3091 1322
rect 3095 1318 3227 1322
rect 3231 1318 3267 1322
rect 3271 1318 3467 1322
rect 3471 1318 3651 1322
rect 3655 1318 3799 1322
rect 3803 1318 3823 1322
rect 1965 1317 3823 1318
rect 3829 1317 3830 1323
rect 3810 1281 3811 1287
rect 3817 1286 5695 1287
rect 3817 1282 3839 1286
rect 3843 1282 4735 1286
rect 4739 1282 4839 1286
rect 4843 1282 4879 1286
rect 4883 1282 4975 1286
rect 4979 1282 5031 1286
rect 5035 1282 5111 1286
rect 5115 1282 5191 1286
rect 5195 1282 5247 1286
rect 5251 1282 5359 1286
rect 5363 1282 5383 1286
rect 5387 1282 5519 1286
rect 5523 1282 5527 1286
rect 5531 1282 5663 1286
rect 5667 1282 5695 1286
rect 3817 1281 5695 1282
rect 5701 1281 5702 1287
rect 1946 1205 1947 1211
rect 1953 1210 3811 1211
rect 1953 1206 1975 1210
rect 1979 1206 2023 1210
rect 2027 1206 2159 1210
rect 2163 1206 2239 1210
rect 2243 1206 2295 1210
rect 2299 1206 2431 1210
rect 2435 1206 2479 1210
rect 2483 1206 2583 1210
rect 2587 1206 2719 1210
rect 2723 1206 2743 1210
rect 2747 1206 2919 1210
rect 2923 1206 2959 1210
rect 2963 1206 3103 1210
rect 3107 1206 3207 1210
rect 3211 1206 3295 1210
rect 3299 1206 3455 1210
rect 3459 1206 3495 1210
rect 3499 1206 3679 1210
rect 3683 1206 3799 1210
rect 3803 1206 3811 1210
rect 1953 1205 3811 1206
rect 3817 1205 3818 1211
rect 96 1181 97 1187
rect 103 1186 1959 1187
rect 103 1182 111 1186
rect 115 1182 131 1186
rect 135 1182 331 1186
rect 335 1182 427 1186
rect 431 1182 563 1186
rect 567 1182 747 1186
rect 751 1182 803 1186
rect 807 1182 1043 1186
rect 1047 1182 1067 1186
rect 1071 1182 1283 1186
rect 1287 1182 1395 1186
rect 1399 1182 1523 1186
rect 1527 1182 1771 1186
rect 1775 1182 1935 1186
rect 1939 1182 1959 1186
rect 103 1181 1959 1182
rect 1965 1181 1966 1187
rect 3822 1161 3823 1167
rect 3829 1166 5707 1167
rect 3829 1162 3839 1166
rect 3843 1162 3859 1166
rect 3863 1162 4067 1166
rect 4071 1162 4299 1166
rect 4303 1162 4539 1166
rect 4543 1162 4707 1166
rect 4711 1162 4779 1166
rect 4783 1162 4851 1166
rect 4855 1162 5003 1166
rect 5007 1162 5027 1166
rect 5031 1162 5163 1166
rect 5167 1162 5283 1166
rect 5287 1162 5331 1166
rect 5335 1162 5499 1166
rect 5503 1162 5515 1166
rect 5519 1162 5663 1166
rect 5667 1162 5707 1166
rect 3829 1161 5707 1162
rect 5713 1161 5714 1167
rect 84 1069 85 1075
rect 91 1074 1947 1075
rect 91 1070 111 1074
rect 115 1070 159 1074
rect 163 1070 263 1074
rect 267 1070 359 1074
rect 363 1070 439 1074
rect 443 1070 591 1074
rect 595 1070 615 1074
rect 619 1070 783 1074
rect 787 1070 831 1074
rect 835 1070 951 1074
rect 955 1070 1071 1074
rect 1075 1070 1111 1074
rect 1115 1070 1271 1074
rect 1275 1070 1311 1074
rect 1315 1070 1431 1074
rect 1435 1070 1551 1074
rect 1555 1070 1591 1074
rect 1595 1070 1751 1074
rect 1755 1070 1799 1074
rect 1803 1070 1935 1074
rect 1939 1070 1947 1074
rect 91 1069 1947 1070
rect 1953 1069 1954 1075
rect 1958 1069 1959 1075
rect 1965 1074 3823 1075
rect 1965 1070 1975 1074
rect 1979 1070 1995 1074
rect 1999 1070 2211 1074
rect 2215 1070 2451 1074
rect 2455 1070 2691 1074
rect 2695 1070 2931 1074
rect 2935 1070 3091 1074
rect 3095 1070 3179 1074
rect 3183 1070 3243 1074
rect 3247 1070 3395 1074
rect 3399 1070 3427 1074
rect 3431 1070 3651 1074
rect 3655 1070 3799 1074
rect 3803 1070 3823 1074
rect 1965 1069 3823 1070
rect 3829 1069 3830 1075
rect 3810 1049 3811 1055
rect 3817 1054 5695 1055
rect 3817 1050 3839 1054
rect 3843 1050 3887 1054
rect 3891 1050 4071 1054
rect 4075 1050 4095 1054
rect 4099 1050 4279 1054
rect 4283 1050 4327 1054
rect 4331 1050 4511 1054
rect 4515 1050 4567 1054
rect 4571 1050 4759 1054
rect 4763 1050 4807 1054
rect 4811 1050 5023 1054
rect 5027 1050 5055 1054
rect 5059 1050 5295 1054
rect 5299 1050 5311 1054
rect 5315 1050 5543 1054
rect 5547 1050 5663 1054
rect 5667 1050 5695 1054
rect 3817 1049 5695 1050
rect 5701 1049 5702 1055
rect 96 953 97 959
rect 103 958 1959 959
rect 103 954 111 958
rect 115 954 227 958
rect 231 954 235 958
rect 239 954 379 958
rect 383 954 411 958
rect 415 954 539 958
rect 543 954 587 958
rect 591 954 715 958
rect 719 954 755 958
rect 759 954 891 958
rect 895 954 923 958
rect 927 954 1075 958
rect 1079 954 1083 958
rect 1087 954 1243 958
rect 1247 954 1259 958
rect 1263 954 1403 958
rect 1407 954 1443 958
rect 1447 954 1563 958
rect 1567 954 1627 958
rect 1631 954 1723 958
rect 1727 954 1787 958
rect 1791 954 1935 958
rect 1939 954 1959 958
rect 103 953 1959 954
rect 1965 953 1966 959
rect 3822 937 3823 943
rect 3829 942 5707 943
rect 3829 938 3839 942
rect 3843 938 3859 942
rect 3863 938 3971 942
rect 3975 938 4043 942
rect 4047 938 4179 942
rect 4183 938 4251 942
rect 4255 938 4403 942
rect 4407 938 4483 942
rect 4487 938 4643 942
rect 4647 938 4731 942
rect 4735 938 4899 942
rect 4903 938 4995 942
rect 4999 938 5171 942
rect 5175 938 5267 942
rect 5271 938 5443 942
rect 5447 938 5515 942
rect 5519 938 5663 942
rect 5667 938 5707 942
rect 3829 937 5707 938
rect 5713 937 5714 943
rect 1946 929 1947 935
rect 1953 934 3811 935
rect 1953 930 1975 934
rect 1979 930 2047 934
rect 2051 930 2351 934
rect 2355 930 2647 934
rect 2651 930 2927 934
rect 2931 930 3119 934
rect 3123 930 3207 934
rect 3211 930 3271 934
rect 3275 930 3423 934
rect 3427 930 3495 934
rect 3499 930 3799 934
rect 3803 930 3811 934
rect 1953 929 3811 930
rect 3817 929 3818 935
rect 84 825 85 831
rect 91 830 1947 831
rect 91 826 111 830
rect 115 826 255 830
rect 259 826 375 830
rect 379 826 407 830
rect 411 826 567 830
rect 571 826 655 830
rect 659 826 743 830
rect 747 826 919 830
rect 923 826 943 830
rect 947 826 1103 830
rect 1107 826 1239 830
rect 1243 826 1287 830
rect 1291 826 1471 830
rect 1475 826 1535 830
rect 1539 826 1655 830
rect 1659 826 1815 830
rect 1819 826 1935 830
rect 1939 826 1947 830
rect 91 825 1947 826
rect 1953 825 1954 831
rect 3810 827 3811 833
rect 3817 831 3842 833
rect 3817 830 5695 831
rect 3817 827 3839 830
rect 3836 826 3839 827
rect 3843 826 3887 830
rect 3891 826 3999 830
rect 4003 826 4047 830
rect 4051 826 4207 830
rect 4211 826 4279 830
rect 4283 826 4431 830
rect 4435 826 4559 830
rect 4563 826 4671 830
rect 4675 826 4879 830
rect 4883 826 4927 830
rect 4931 826 5199 830
rect 5203 826 5223 830
rect 5227 826 5471 830
rect 5475 826 5543 830
rect 5547 826 5663 830
rect 5667 826 5695 830
rect 3836 825 5695 826
rect 5701 825 5702 831
rect 1958 817 1959 823
rect 1965 822 3823 823
rect 1965 818 1975 822
rect 1979 818 1995 822
rect 1999 818 2019 822
rect 2023 818 2251 822
rect 2255 818 2323 822
rect 2327 818 2523 822
rect 2527 818 2619 822
rect 2623 818 2771 822
rect 2775 818 2899 822
rect 2903 818 3003 822
rect 3007 818 3179 822
rect 3183 818 3227 822
rect 3231 818 3451 822
rect 3455 818 3467 822
rect 3471 818 3651 822
rect 3655 818 3799 822
rect 3803 818 3823 822
rect 1965 817 3823 818
rect 3829 817 3830 823
rect 96 713 97 719
rect 103 718 1959 719
rect 103 714 111 718
rect 115 714 131 718
rect 135 714 307 718
rect 311 714 347 718
rect 351 714 499 718
rect 503 714 627 718
rect 631 714 683 718
rect 687 714 859 718
rect 863 714 915 718
rect 919 714 1027 718
rect 1031 714 1187 718
rect 1191 714 1211 718
rect 1215 714 1339 718
rect 1343 714 1491 718
rect 1495 714 1507 718
rect 1511 714 1651 718
rect 1655 714 1787 718
rect 1791 714 1935 718
rect 1939 714 1959 718
rect 103 713 1959 714
rect 1965 713 1966 719
rect 3822 705 3823 711
rect 3829 710 5707 711
rect 3829 706 3839 710
rect 3843 706 3859 710
rect 3863 706 3995 710
rect 3999 706 4019 710
rect 4023 706 4131 710
rect 4135 706 4251 710
rect 4255 706 4267 710
rect 4271 706 4403 710
rect 4407 706 4531 710
rect 4535 706 4571 710
rect 4575 706 4771 710
rect 4775 706 4851 710
rect 4855 706 4995 710
rect 4999 706 5195 710
rect 5199 706 5227 710
rect 5231 706 5459 710
rect 5463 706 5515 710
rect 5519 706 5663 710
rect 5667 706 5707 710
rect 3829 705 5707 706
rect 5713 705 5714 711
rect 84 601 85 607
rect 91 606 1947 607
rect 91 602 111 606
rect 115 602 159 606
rect 163 602 335 606
rect 339 602 375 606
rect 379 602 527 606
rect 531 602 599 606
rect 603 602 711 606
rect 715 602 807 606
rect 811 602 887 606
rect 891 602 999 606
rect 1003 602 1055 606
rect 1059 602 1175 606
rect 1179 602 1215 606
rect 1219 602 1343 606
rect 1347 602 1367 606
rect 1371 602 1511 606
rect 1515 602 1519 606
rect 1523 602 1671 606
rect 1675 602 1679 606
rect 1683 602 1815 606
rect 1819 602 1935 606
rect 1939 602 1947 606
rect 91 601 1947 602
rect 1953 601 1954 607
rect 3810 593 3811 599
rect 3817 598 5695 599
rect 3817 594 3839 598
rect 3843 594 3887 598
rect 3891 594 4023 598
rect 4027 594 4159 598
rect 4163 594 4295 598
rect 4299 594 4431 598
rect 4435 594 4479 598
rect 4483 594 4599 598
rect 4603 594 4695 598
rect 4699 594 4799 598
rect 4803 594 4935 598
rect 4939 594 5023 598
rect 5027 594 5191 598
rect 5195 594 5255 598
rect 5259 594 5447 598
rect 5451 594 5487 598
rect 5491 594 5663 598
rect 5667 594 5695 598
rect 3817 593 5695 594
rect 5701 593 5702 599
rect 1946 573 1947 579
rect 1953 578 3811 579
rect 1953 574 1975 578
rect 1979 574 2023 578
rect 2027 574 2279 578
rect 2283 574 2551 578
rect 2555 574 2799 578
rect 2803 574 3031 578
rect 3035 574 3255 578
rect 3259 574 3311 578
rect 3315 574 3447 578
rect 3451 574 3479 578
rect 3483 574 3583 578
rect 3587 574 3679 578
rect 3683 574 3799 578
rect 3803 574 3811 578
rect 1953 573 3811 574
rect 3817 573 3818 579
rect 96 489 97 495
rect 103 494 1959 495
rect 103 490 111 494
rect 115 490 131 494
rect 135 490 347 494
rect 351 490 427 494
rect 431 490 571 494
rect 575 490 763 494
rect 767 490 779 494
rect 783 490 971 494
rect 975 490 1107 494
rect 1111 490 1147 494
rect 1151 490 1315 494
rect 1319 490 1459 494
rect 1463 490 1483 494
rect 1487 490 1643 494
rect 1647 490 1787 494
rect 1791 490 1935 494
rect 1939 490 1959 494
rect 103 489 1959 490
rect 1965 489 1966 495
rect 3822 469 3823 475
rect 3829 474 5707 475
rect 3829 470 3839 474
rect 3843 470 3859 474
rect 3863 470 3995 474
rect 3999 470 4131 474
rect 4135 470 4267 474
rect 4271 470 4451 474
rect 4455 470 4651 474
rect 4655 470 4667 474
rect 4671 470 4859 474
rect 4863 470 4907 474
rect 4911 470 5067 474
rect 5071 470 5163 474
rect 5167 470 5283 474
rect 5287 470 5419 474
rect 5423 470 5507 474
rect 5511 470 5663 474
rect 5667 470 5707 474
rect 3829 469 5707 470
rect 5713 469 5714 475
rect 3822 467 3830 469
rect 1958 461 1959 467
rect 1965 466 3823 467
rect 1965 462 1975 466
rect 1979 462 1995 466
rect 1999 462 2155 466
rect 2159 462 2347 466
rect 2351 462 2539 466
rect 2543 462 2731 466
rect 2735 462 2923 466
rect 2927 462 3115 466
rect 3119 462 3283 466
rect 3287 462 3299 466
rect 3303 462 3419 466
rect 3423 462 3483 466
rect 3487 462 3555 466
rect 3559 462 3651 466
rect 3655 462 3799 466
rect 3803 462 3823 466
rect 1965 461 3823 462
rect 3829 461 3830 467
rect 84 361 85 367
rect 91 366 1947 367
rect 91 362 111 366
rect 115 362 159 366
rect 163 362 239 366
rect 243 362 391 366
rect 395 362 455 366
rect 459 362 551 366
rect 555 362 711 366
rect 715 362 791 366
rect 795 362 871 366
rect 875 362 1031 366
rect 1035 362 1135 366
rect 1139 362 1487 366
rect 1491 362 1815 366
rect 1819 362 1935 366
rect 1939 362 1947 366
rect 91 361 1947 362
rect 1953 361 1954 367
rect 3810 353 3811 359
rect 3817 358 5695 359
rect 3817 354 3839 358
rect 3843 354 4479 358
rect 4483 354 4679 358
rect 4683 354 4751 358
rect 4755 354 4887 358
rect 4891 354 4911 358
rect 4915 354 5071 358
rect 5075 354 5095 358
rect 5099 354 5231 358
rect 5235 354 5311 358
rect 5315 354 5399 358
rect 5403 354 5535 358
rect 5539 354 5543 358
rect 5547 354 5663 358
rect 5667 354 5695 358
rect 3817 353 5695 354
rect 5701 353 5702 359
rect 1946 325 1947 331
rect 1953 330 3811 331
rect 1953 326 1975 330
rect 1979 326 2023 330
rect 2027 326 2047 330
rect 2051 326 2183 330
rect 2187 326 2319 330
rect 2323 326 2375 330
rect 2379 326 2455 330
rect 2459 326 2567 330
rect 2571 326 2591 330
rect 2595 326 2727 330
rect 2731 326 2759 330
rect 2763 326 2863 330
rect 2867 326 2951 330
rect 2955 326 2999 330
rect 3003 326 3135 330
rect 3139 326 3143 330
rect 3147 326 3271 330
rect 3275 326 3327 330
rect 3331 326 3407 330
rect 3411 326 3511 330
rect 3515 326 3543 330
rect 3547 326 3679 330
rect 3683 326 3799 330
rect 3803 326 3811 330
rect 1953 325 3811 326
rect 3817 325 3818 331
rect 96 217 97 223
rect 103 222 1959 223
rect 103 218 111 222
rect 115 218 147 222
rect 151 218 211 222
rect 215 218 283 222
rect 287 218 363 222
rect 367 218 419 222
rect 423 218 523 222
rect 527 218 555 222
rect 559 218 683 222
rect 687 218 691 222
rect 695 218 827 222
rect 831 218 843 222
rect 847 218 963 222
rect 967 218 1003 222
rect 1007 218 1099 222
rect 1103 218 1935 222
rect 1939 218 1959 222
rect 103 217 1959 218
rect 1965 217 1966 223
rect 3822 206 5714 207
rect 3822 203 3839 206
rect 1958 197 1959 203
rect 1965 202 3823 203
rect 1965 198 1975 202
rect 1979 198 1995 202
rect 1999 198 2019 202
rect 2023 198 2131 202
rect 2135 198 2155 202
rect 2159 198 2267 202
rect 2271 198 2291 202
rect 2295 198 2403 202
rect 2407 198 2427 202
rect 2431 198 2539 202
rect 2543 198 2563 202
rect 2567 198 2675 202
rect 2679 198 2699 202
rect 2703 198 2811 202
rect 2815 198 2835 202
rect 2839 198 2947 202
rect 2951 198 2971 202
rect 2975 198 3083 202
rect 3087 198 3107 202
rect 3111 198 3219 202
rect 3223 198 3243 202
rect 3247 198 3355 202
rect 3359 198 3379 202
rect 3383 198 3491 202
rect 3495 198 3515 202
rect 3519 198 3627 202
rect 3631 198 3651 202
rect 3655 198 3799 202
rect 3803 198 3823 202
rect 1965 197 3823 198
rect 3829 202 3839 203
rect 3843 202 4291 206
rect 4295 202 4427 206
rect 4431 202 4563 206
rect 4567 202 4699 206
rect 4703 202 4723 206
rect 4727 202 4835 206
rect 4839 202 4883 206
rect 4887 202 4971 206
rect 4975 202 5043 206
rect 5047 202 5107 206
rect 5111 202 5203 206
rect 5207 202 5243 206
rect 5247 202 5371 206
rect 5375 202 5379 206
rect 5383 202 5515 206
rect 5519 202 5663 206
rect 5667 202 5714 206
rect 3829 201 5714 202
rect 3829 197 3830 201
rect 84 105 85 111
rect 91 110 1947 111
rect 91 106 111 110
rect 115 106 175 110
rect 179 106 311 110
rect 315 106 447 110
rect 451 106 583 110
rect 587 106 719 110
rect 723 106 855 110
rect 859 106 991 110
rect 995 106 1127 110
rect 1131 106 1935 110
rect 1939 106 1947 110
rect 91 105 1947 106
rect 1953 105 1954 111
rect 3810 94 5702 95
rect 3810 91 3839 94
rect 1946 85 1947 91
rect 1953 90 3811 91
rect 1953 86 1975 90
rect 1979 86 2023 90
rect 2027 86 2159 90
rect 2163 86 2295 90
rect 2299 86 2431 90
rect 2435 86 2567 90
rect 2571 86 2703 90
rect 2707 86 2839 90
rect 2843 86 2975 90
rect 2979 86 3111 90
rect 3115 86 3247 90
rect 3251 86 3383 90
rect 3387 86 3519 90
rect 3523 86 3655 90
rect 3659 86 3799 90
rect 3803 86 3811 90
rect 1953 85 3811 86
rect 3817 90 3839 91
rect 3843 90 4319 94
rect 4323 90 4455 94
rect 4459 90 4591 94
rect 4595 90 4727 94
rect 4731 90 4863 94
rect 4867 90 4999 94
rect 5003 90 5135 94
rect 5139 90 5271 94
rect 5275 90 5407 94
rect 5411 90 5543 94
rect 5547 90 5663 94
rect 5667 90 5702 94
rect 3817 89 5702 90
rect 3817 85 3818 89
<< m5c >>
rect 97 5753 103 5759
rect 1959 5753 1965 5759
rect 1959 5685 1965 5691
rect 3823 5685 3829 5691
rect 85 5641 91 5647
rect 1947 5641 1953 5647
rect 1947 5573 1953 5579
rect 3811 5573 3817 5579
rect 97 5529 103 5535
rect 1959 5529 1965 5535
rect 3823 5465 3829 5471
rect 5707 5465 5713 5471
rect 1959 5457 1965 5463
rect 3823 5457 3829 5463
rect 85 5417 91 5423
rect 1947 5417 1953 5423
rect 1947 5345 1953 5351
rect 3811 5345 3817 5351
rect 97 5305 103 5311
rect 1959 5305 1965 5311
rect 1959 5229 1965 5235
rect 3823 5229 3829 5235
rect 3823 5217 3829 5223
rect 5707 5217 5713 5223
rect 85 5193 91 5199
rect 1947 5193 1953 5199
rect 1947 5101 1953 5107
rect 3811 5101 3817 5107
rect 97 5073 103 5079
rect 1959 5073 1965 5079
rect 1959 4981 1965 4987
rect 3823 4981 3829 4987
rect 85 4933 91 4939
rect 1947 4933 1953 4939
rect 1947 4861 1953 4867
rect 3811 4861 3817 4867
rect 97 4809 103 4815
rect 1959 4809 1965 4815
rect 3811 4797 3817 4803
rect 5695 4797 5701 4803
rect 1959 4737 1965 4743
rect 3823 4737 3829 4743
rect 85 4693 91 4699
rect 1947 4693 1953 4699
rect 3823 4685 3829 4691
rect 5707 4685 5713 4691
rect 1947 4621 1953 4627
rect 3811 4621 3817 4627
rect 97 4569 103 4575
rect 1959 4569 1965 4575
rect 3811 4573 3817 4579
rect 5695 4573 5701 4579
rect 1959 4497 1965 4503
rect 3823 4497 3829 4503
rect 85 4457 91 4463
rect 1947 4457 1953 4463
rect 3823 4457 3829 4463
rect 5707 4457 5713 4463
rect 1947 4373 1953 4379
rect 3811 4373 3817 4379
rect 97 4341 103 4347
rect 1959 4341 1965 4347
rect 3811 4329 3817 4335
rect 5695 4329 5701 4335
rect 1959 4257 1965 4263
rect 3823 4257 3829 4263
rect 85 4221 91 4227
rect 1947 4221 1953 4227
rect 3823 4205 3829 4211
rect 5707 4205 5713 4211
rect 1947 4133 1953 4139
rect 3811 4133 3817 4139
rect 97 4109 103 4115
rect 1959 4109 1965 4115
rect 3811 4069 3817 4075
rect 5695 4069 5701 4075
rect 85 3997 91 4003
rect 1947 3997 1953 4003
rect 3823 3957 3829 3963
rect 5707 3957 5713 3963
rect 1959 3929 1965 3935
rect 3823 3929 3829 3935
rect 97 3885 103 3891
rect 1959 3885 1965 3891
rect 1947 3817 1953 3823
rect 3811 3817 3817 3823
rect 85 3761 91 3767
rect 1947 3761 1953 3767
rect 1959 3697 1965 3703
rect 3823 3697 3829 3703
rect 3823 3685 3829 3691
rect 5707 3685 5713 3691
rect 97 3633 103 3639
rect 1959 3633 1965 3639
rect 1947 3577 1953 3583
rect 3811 3577 3817 3583
rect 3811 3525 3817 3531
rect 5695 3525 5701 3531
rect 85 3501 91 3507
rect 1947 3501 1953 3507
rect 1959 3461 1965 3467
rect 3823 3461 3829 3467
rect 3823 3405 3829 3411
rect 5707 3405 5713 3411
rect 97 3381 103 3387
rect 1959 3381 1965 3387
rect 1947 3325 1953 3331
rect 3811 3325 3817 3331
rect 3811 3293 3817 3299
rect 5695 3293 5701 3299
rect 85 3261 91 3267
rect 1947 3261 1953 3267
rect 1959 3213 1965 3219
rect 3823 3213 3829 3219
rect 3823 3165 3829 3171
rect 5707 3165 5713 3171
rect 97 3133 103 3139
rect 1959 3133 1965 3139
rect 1947 3101 1953 3107
rect 3811 3101 3817 3107
rect 3811 3053 3817 3059
rect 5695 3053 5701 3059
rect 85 3021 91 3027
rect 1947 3021 1953 3027
rect 1959 2989 1965 2995
rect 3823 2989 3829 2995
rect 3823 2917 3829 2923
rect 5707 2917 5713 2923
rect 97 2905 103 2911
rect 1959 2905 1965 2911
rect 1947 2825 1953 2831
rect 3811 2825 3817 2831
rect 3811 2801 3817 2807
rect 5695 2801 5701 2807
rect 85 2781 91 2787
rect 1947 2781 1953 2787
rect 1959 2713 1965 2719
rect 3823 2713 3829 2719
rect 3823 2677 3829 2683
rect 5707 2677 5713 2683
rect 97 2669 103 2675
rect 1959 2669 1965 2675
rect 1947 2597 1953 2603
rect 3811 2597 3817 2603
rect 3811 2561 3817 2567
rect 5695 2561 5701 2567
rect 85 2541 91 2547
rect 1947 2541 1953 2547
rect 1959 2469 1965 2475
rect 3823 2469 3829 2475
rect 3823 2433 3829 2439
rect 5707 2433 5713 2439
rect 97 2417 103 2423
rect 1959 2417 1965 2423
rect 1947 2349 1953 2355
rect 3811 2349 3817 2355
rect 3811 2309 3817 2315
rect 5695 2309 5701 2315
rect 85 2301 91 2307
rect 1947 2301 1953 2307
rect 1959 2237 1965 2243
rect 3823 2237 3829 2243
rect 3823 2193 3829 2199
rect 5707 2193 5713 2199
rect 97 2165 103 2171
rect 1959 2165 1965 2171
rect 3811 2061 3817 2067
rect 5695 2061 5701 2067
rect 85 2049 91 2055
rect 1947 2049 1953 2055
rect 3823 1949 3829 1955
rect 5707 1949 5713 1955
rect 1947 1935 1953 1941
rect 97 1925 103 1931
rect 1959 1925 1965 1931
rect 3811 1925 3817 1931
rect 3811 1837 3817 1843
rect 5695 1837 5701 1843
rect 85 1801 91 1807
rect 1947 1801 1953 1807
rect 1959 1801 1965 1807
rect 3823 1801 3829 1807
rect 3823 1709 3829 1715
rect 5707 1709 5713 1715
rect 1947 1687 1953 1693
rect 97 1677 103 1683
rect 1959 1677 1965 1683
rect 3811 1677 3817 1683
rect 3811 1581 3817 1587
rect 5695 1581 5701 1587
rect 85 1553 91 1559
rect 1947 1553 1953 1559
rect 1959 1553 1965 1559
rect 3823 1553 3829 1559
rect 1947 1439 1953 1445
rect 97 1429 103 1435
rect 1959 1429 1965 1435
rect 3811 1429 3817 1435
rect 3823 1397 3829 1403
rect 5707 1397 5713 1403
rect 85 1317 91 1323
rect 1947 1317 1953 1323
rect 1959 1317 1965 1323
rect 3823 1317 3829 1323
rect 3811 1281 3817 1287
rect 5695 1281 5701 1287
rect 1947 1205 1953 1211
rect 3811 1205 3817 1211
rect 97 1181 103 1187
rect 1959 1181 1965 1187
rect 3823 1161 3829 1167
rect 5707 1161 5713 1167
rect 85 1069 91 1075
rect 1947 1069 1953 1075
rect 1959 1069 1965 1075
rect 3823 1069 3829 1075
rect 3811 1049 3817 1055
rect 5695 1049 5701 1055
rect 97 953 103 959
rect 1959 953 1965 959
rect 3823 937 3829 943
rect 5707 937 5713 943
rect 1947 929 1953 935
rect 3811 929 3817 935
rect 85 825 91 831
rect 1947 825 1953 831
rect 3811 827 3817 833
rect 5695 825 5701 831
rect 1959 817 1965 823
rect 3823 817 3829 823
rect 97 713 103 719
rect 1959 713 1965 719
rect 3823 705 3829 711
rect 5707 705 5713 711
rect 85 601 91 607
rect 1947 601 1953 607
rect 3811 593 3817 599
rect 5695 593 5701 599
rect 1947 573 1953 579
rect 3811 573 3817 579
rect 97 489 103 495
rect 1959 489 1965 495
rect 3823 469 3829 475
rect 5707 469 5713 475
rect 1959 461 1965 467
rect 3823 461 3829 467
rect 85 361 91 367
rect 1947 361 1953 367
rect 3811 353 3817 359
rect 5695 353 5701 359
rect 1947 325 1953 331
rect 3811 325 3817 331
rect 97 217 103 223
rect 1959 217 1965 223
rect 1959 197 1965 203
rect 3823 197 3829 203
rect 85 105 91 111
rect 1947 105 1953 111
rect 1947 85 1953 91
rect 3811 85 3817 91
<< m5 >>
rect 84 5647 92 5760
rect 84 5641 85 5647
rect 91 5641 92 5647
rect 84 5423 92 5641
rect 84 5417 85 5423
rect 91 5417 92 5423
rect 84 5199 92 5417
rect 84 5193 85 5199
rect 91 5193 92 5199
rect 84 4939 92 5193
rect 84 4933 85 4939
rect 91 4933 92 4939
rect 84 4699 92 4933
rect 84 4693 85 4699
rect 91 4693 92 4699
rect 84 4463 92 4693
rect 84 4457 85 4463
rect 91 4457 92 4463
rect 84 4227 92 4457
rect 84 4221 85 4227
rect 91 4221 92 4227
rect 84 4003 92 4221
rect 84 3997 85 4003
rect 91 3997 92 4003
rect 84 3767 92 3997
rect 84 3761 85 3767
rect 91 3761 92 3767
rect 84 3507 92 3761
rect 84 3501 85 3507
rect 91 3501 92 3507
rect 84 3267 92 3501
rect 84 3261 85 3267
rect 91 3261 92 3267
rect 84 3027 92 3261
rect 84 3021 85 3027
rect 91 3021 92 3027
rect 84 2787 92 3021
rect 84 2781 85 2787
rect 91 2781 92 2787
rect 84 2547 92 2781
rect 84 2541 85 2547
rect 91 2541 92 2547
rect 84 2307 92 2541
rect 84 2301 85 2307
rect 91 2301 92 2307
rect 84 2055 92 2301
rect 84 2049 85 2055
rect 91 2049 92 2055
rect 84 1807 92 2049
rect 84 1801 85 1807
rect 91 1801 92 1807
rect 84 1559 92 1801
rect 84 1553 85 1559
rect 91 1553 92 1559
rect 84 1323 92 1553
rect 84 1317 85 1323
rect 91 1317 92 1323
rect 84 1075 92 1317
rect 84 1069 85 1075
rect 91 1069 92 1075
rect 84 831 92 1069
rect 84 825 85 831
rect 91 825 92 831
rect 84 607 92 825
rect 84 601 85 607
rect 91 601 92 607
rect 84 367 92 601
rect 84 361 85 367
rect 91 361 92 367
rect 84 111 92 361
rect 84 105 85 111
rect 91 105 92 111
rect 84 72 92 105
rect 96 5759 104 5760
rect 96 5753 97 5759
rect 103 5753 104 5759
rect 96 5535 104 5753
rect 96 5529 97 5535
rect 103 5529 104 5535
rect 96 5311 104 5529
rect 96 5305 97 5311
rect 103 5305 104 5311
rect 96 5079 104 5305
rect 96 5073 97 5079
rect 103 5073 104 5079
rect 96 4815 104 5073
rect 96 4809 97 4815
rect 103 4809 104 4815
rect 96 4575 104 4809
rect 96 4569 97 4575
rect 103 4569 104 4575
rect 96 4347 104 4569
rect 96 4341 97 4347
rect 103 4341 104 4347
rect 96 4115 104 4341
rect 96 4109 97 4115
rect 103 4109 104 4115
rect 96 3891 104 4109
rect 96 3885 97 3891
rect 103 3885 104 3891
rect 96 3639 104 3885
rect 96 3633 97 3639
rect 103 3633 104 3639
rect 96 3387 104 3633
rect 96 3381 97 3387
rect 103 3381 104 3387
rect 96 3139 104 3381
rect 96 3133 97 3139
rect 103 3133 104 3139
rect 96 2911 104 3133
rect 96 2905 97 2911
rect 103 2905 104 2911
rect 96 2675 104 2905
rect 96 2669 97 2675
rect 103 2669 104 2675
rect 96 2423 104 2669
rect 96 2417 97 2423
rect 103 2417 104 2423
rect 96 2171 104 2417
rect 96 2165 97 2171
rect 103 2165 104 2171
rect 96 1931 104 2165
rect 96 1925 97 1931
rect 103 1925 104 1931
rect 96 1683 104 1925
rect 96 1677 97 1683
rect 103 1677 104 1683
rect 96 1435 104 1677
rect 96 1429 97 1435
rect 103 1429 104 1435
rect 96 1187 104 1429
rect 96 1181 97 1187
rect 103 1181 104 1187
rect 96 959 104 1181
rect 96 953 97 959
rect 103 953 104 959
rect 96 719 104 953
rect 96 713 97 719
rect 103 713 104 719
rect 96 495 104 713
rect 96 489 97 495
rect 103 489 104 495
rect 96 223 104 489
rect 96 217 97 223
rect 103 217 104 223
rect 96 72 104 217
rect 1946 5647 1954 5760
rect 1946 5641 1947 5647
rect 1953 5641 1954 5647
rect 1946 5579 1954 5641
rect 1946 5573 1947 5579
rect 1953 5573 1954 5579
rect 1946 5423 1954 5573
rect 1946 5417 1947 5423
rect 1953 5417 1954 5423
rect 1946 5351 1954 5417
rect 1946 5345 1947 5351
rect 1953 5345 1954 5351
rect 1946 5199 1954 5345
rect 1946 5193 1947 5199
rect 1953 5193 1954 5199
rect 1946 5107 1954 5193
rect 1946 5101 1947 5107
rect 1953 5101 1954 5107
rect 1946 4939 1954 5101
rect 1946 4933 1947 4939
rect 1953 4933 1954 4939
rect 1946 4867 1954 4933
rect 1946 4861 1947 4867
rect 1953 4861 1954 4867
rect 1946 4699 1954 4861
rect 1946 4693 1947 4699
rect 1953 4693 1954 4699
rect 1946 4627 1954 4693
rect 1946 4621 1947 4627
rect 1953 4621 1954 4627
rect 1946 4463 1954 4621
rect 1946 4457 1947 4463
rect 1953 4457 1954 4463
rect 1946 4379 1954 4457
rect 1946 4373 1947 4379
rect 1953 4373 1954 4379
rect 1946 4227 1954 4373
rect 1946 4221 1947 4227
rect 1953 4221 1954 4227
rect 1946 4139 1954 4221
rect 1946 4133 1947 4139
rect 1953 4133 1954 4139
rect 1946 4003 1954 4133
rect 1946 3997 1947 4003
rect 1953 3997 1954 4003
rect 1946 3823 1954 3997
rect 1946 3817 1947 3823
rect 1953 3817 1954 3823
rect 1946 3767 1954 3817
rect 1946 3761 1947 3767
rect 1953 3761 1954 3767
rect 1946 3583 1954 3761
rect 1946 3577 1947 3583
rect 1953 3577 1954 3583
rect 1946 3507 1954 3577
rect 1946 3501 1947 3507
rect 1953 3501 1954 3507
rect 1946 3331 1954 3501
rect 1946 3325 1947 3331
rect 1953 3325 1954 3331
rect 1946 3267 1954 3325
rect 1946 3261 1947 3267
rect 1953 3261 1954 3267
rect 1946 3107 1954 3261
rect 1946 3101 1947 3107
rect 1953 3101 1954 3107
rect 1946 3027 1954 3101
rect 1946 3021 1947 3027
rect 1953 3021 1954 3027
rect 1946 2831 1954 3021
rect 1946 2825 1947 2831
rect 1953 2825 1954 2831
rect 1946 2787 1954 2825
rect 1946 2781 1947 2787
rect 1953 2781 1954 2787
rect 1946 2603 1954 2781
rect 1946 2597 1947 2603
rect 1953 2597 1954 2603
rect 1946 2547 1954 2597
rect 1946 2541 1947 2547
rect 1953 2541 1954 2547
rect 1946 2355 1954 2541
rect 1946 2349 1947 2355
rect 1953 2349 1954 2355
rect 1946 2307 1954 2349
rect 1946 2301 1947 2307
rect 1953 2301 1954 2307
rect 1946 2055 1954 2301
rect 1946 2049 1947 2055
rect 1953 2049 1954 2055
rect 1946 1941 1954 2049
rect 1946 1935 1947 1941
rect 1953 1935 1954 1941
rect 1946 1807 1954 1935
rect 1946 1801 1947 1807
rect 1953 1801 1954 1807
rect 1946 1693 1954 1801
rect 1946 1687 1947 1693
rect 1953 1687 1954 1693
rect 1946 1559 1954 1687
rect 1946 1553 1947 1559
rect 1953 1553 1954 1559
rect 1946 1445 1954 1553
rect 1946 1439 1947 1445
rect 1953 1439 1954 1445
rect 1946 1323 1954 1439
rect 1946 1317 1947 1323
rect 1953 1317 1954 1323
rect 1946 1211 1954 1317
rect 1946 1205 1947 1211
rect 1953 1205 1954 1211
rect 1946 1075 1954 1205
rect 1946 1069 1947 1075
rect 1953 1069 1954 1075
rect 1946 935 1954 1069
rect 1946 929 1947 935
rect 1953 929 1954 935
rect 1946 831 1954 929
rect 1946 825 1947 831
rect 1953 825 1954 831
rect 1946 607 1954 825
rect 1946 601 1947 607
rect 1953 601 1954 607
rect 1946 579 1954 601
rect 1946 573 1947 579
rect 1953 573 1954 579
rect 1946 367 1954 573
rect 1946 361 1947 367
rect 1953 361 1954 367
rect 1946 331 1954 361
rect 1946 325 1947 331
rect 1953 325 1954 331
rect 1946 111 1954 325
rect 1946 105 1947 111
rect 1953 105 1954 111
rect 1946 91 1954 105
rect 1946 85 1947 91
rect 1953 85 1954 91
rect 1946 72 1954 85
rect 1958 5759 1966 5760
rect 1958 5753 1959 5759
rect 1965 5753 1966 5759
rect 1958 5691 1966 5753
rect 1958 5685 1959 5691
rect 1965 5685 1966 5691
rect 1958 5535 1966 5685
rect 1958 5529 1959 5535
rect 1965 5529 1966 5535
rect 1958 5463 1966 5529
rect 1958 5457 1959 5463
rect 1965 5457 1966 5463
rect 1958 5311 1966 5457
rect 1958 5305 1959 5311
rect 1965 5305 1966 5311
rect 1958 5235 1966 5305
rect 1958 5229 1959 5235
rect 1965 5229 1966 5235
rect 1958 5079 1966 5229
rect 1958 5073 1959 5079
rect 1965 5073 1966 5079
rect 1958 4987 1966 5073
rect 1958 4981 1959 4987
rect 1965 4981 1966 4987
rect 1958 4815 1966 4981
rect 1958 4809 1959 4815
rect 1965 4809 1966 4815
rect 1958 4743 1966 4809
rect 1958 4737 1959 4743
rect 1965 4737 1966 4743
rect 1958 4575 1966 4737
rect 1958 4569 1959 4575
rect 1965 4569 1966 4575
rect 1958 4503 1966 4569
rect 1958 4497 1959 4503
rect 1965 4497 1966 4503
rect 1958 4347 1966 4497
rect 1958 4341 1959 4347
rect 1965 4341 1966 4347
rect 1958 4263 1966 4341
rect 1958 4257 1959 4263
rect 1965 4257 1966 4263
rect 1958 4115 1966 4257
rect 1958 4109 1959 4115
rect 1965 4109 1966 4115
rect 1958 3935 1966 4109
rect 1958 3929 1959 3935
rect 1965 3929 1966 3935
rect 1958 3891 1966 3929
rect 1958 3885 1959 3891
rect 1965 3885 1966 3891
rect 1958 3703 1966 3885
rect 1958 3697 1959 3703
rect 1965 3697 1966 3703
rect 1958 3639 1966 3697
rect 1958 3633 1959 3639
rect 1965 3633 1966 3639
rect 1958 3467 1966 3633
rect 1958 3461 1959 3467
rect 1965 3461 1966 3467
rect 1958 3387 1966 3461
rect 1958 3381 1959 3387
rect 1965 3381 1966 3387
rect 1958 3219 1966 3381
rect 1958 3213 1959 3219
rect 1965 3213 1966 3219
rect 1958 3139 1966 3213
rect 1958 3133 1959 3139
rect 1965 3133 1966 3139
rect 1958 2995 1966 3133
rect 1958 2989 1959 2995
rect 1965 2989 1966 2995
rect 1958 2911 1966 2989
rect 1958 2905 1959 2911
rect 1965 2905 1966 2911
rect 1958 2719 1966 2905
rect 1958 2713 1959 2719
rect 1965 2713 1966 2719
rect 1958 2675 1966 2713
rect 1958 2669 1959 2675
rect 1965 2669 1966 2675
rect 1958 2475 1966 2669
rect 1958 2469 1959 2475
rect 1965 2469 1966 2475
rect 1958 2423 1966 2469
rect 1958 2417 1959 2423
rect 1965 2417 1966 2423
rect 1958 2243 1966 2417
rect 1958 2237 1959 2243
rect 1965 2237 1966 2243
rect 1958 2171 1966 2237
rect 1958 2165 1959 2171
rect 1965 2165 1966 2171
rect 1958 1931 1966 2165
rect 1958 1925 1959 1931
rect 1965 1925 1966 1931
rect 1958 1807 1966 1925
rect 1958 1801 1959 1807
rect 1965 1801 1966 1807
rect 1958 1683 1966 1801
rect 1958 1677 1959 1683
rect 1965 1677 1966 1683
rect 1958 1559 1966 1677
rect 1958 1553 1959 1559
rect 1965 1553 1966 1559
rect 1958 1435 1966 1553
rect 1958 1429 1959 1435
rect 1965 1429 1966 1435
rect 1958 1323 1966 1429
rect 1958 1317 1959 1323
rect 1965 1317 1966 1323
rect 1958 1187 1966 1317
rect 1958 1181 1959 1187
rect 1965 1181 1966 1187
rect 1958 1075 1966 1181
rect 1958 1069 1959 1075
rect 1965 1069 1966 1075
rect 1958 959 1966 1069
rect 1958 953 1959 959
rect 1965 953 1966 959
rect 1958 823 1966 953
rect 1958 817 1959 823
rect 1965 817 1966 823
rect 1958 719 1966 817
rect 1958 713 1959 719
rect 1965 713 1966 719
rect 1958 495 1966 713
rect 1958 489 1959 495
rect 1965 489 1966 495
rect 1958 467 1966 489
rect 1958 461 1959 467
rect 1965 461 1966 467
rect 1958 223 1966 461
rect 1958 217 1959 223
rect 1965 217 1966 223
rect 1958 203 1966 217
rect 1958 197 1959 203
rect 1965 197 1966 203
rect 1958 72 1966 197
rect 3810 5579 3818 5760
rect 3810 5573 3811 5579
rect 3817 5573 3818 5579
rect 3810 5351 3818 5573
rect 3810 5345 3811 5351
rect 3817 5345 3818 5351
rect 3810 5107 3818 5345
rect 3810 5101 3811 5107
rect 3817 5101 3818 5107
rect 3810 4867 3818 5101
rect 3810 4861 3811 4867
rect 3817 4861 3818 4867
rect 3810 4803 3818 4861
rect 3810 4797 3811 4803
rect 3817 4797 3818 4803
rect 3810 4627 3818 4797
rect 3810 4621 3811 4627
rect 3817 4621 3818 4627
rect 3810 4579 3818 4621
rect 3810 4573 3811 4579
rect 3817 4573 3818 4579
rect 3810 4379 3818 4573
rect 3810 4373 3811 4379
rect 3817 4373 3818 4379
rect 3810 4335 3818 4373
rect 3810 4329 3811 4335
rect 3817 4329 3818 4335
rect 3810 4139 3818 4329
rect 3810 4133 3811 4139
rect 3817 4133 3818 4139
rect 3810 4075 3818 4133
rect 3810 4069 3811 4075
rect 3817 4069 3818 4075
rect 3810 3823 3818 4069
rect 3810 3817 3811 3823
rect 3817 3817 3818 3823
rect 3810 3583 3818 3817
rect 3810 3577 3811 3583
rect 3817 3577 3818 3583
rect 3810 3531 3818 3577
rect 3810 3525 3811 3531
rect 3817 3525 3818 3531
rect 3810 3331 3818 3525
rect 3810 3325 3811 3331
rect 3817 3325 3818 3331
rect 3810 3299 3818 3325
rect 3810 3293 3811 3299
rect 3817 3293 3818 3299
rect 3810 3107 3818 3293
rect 3810 3101 3811 3107
rect 3817 3101 3818 3107
rect 3810 3059 3818 3101
rect 3810 3053 3811 3059
rect 3817 3053 3818 3059
rect 3810 2831 3818 3053
rect 3810 2825 3811 2831
rect 3817 2825 3818 2831
rect 3810 2807 3818 2825
rect 3810 2801 3811 2807
rect 3817 2801 3818 2807
rect 3810 2603 3818 2801
rect 3810 2597 3811 2603
rect 3817 2597 3818 2603
rect 3810 2567 3818 2597
rect 3810 2561 3811 2567
rect 3817 2561 3818 2567
rect 3810 2355 3818 2561
rect 3810 2349 3811 2355
rect 3817 2349 3818 2355
rect 3810 2315 3818 2349
rect 3810 2309 3811 2315
rect 3817 2309 3818 2315
rect 3810 2067 3818 2309
rect 3810 2061 3811 2067
rect 3817 2061 3818 2067
rect 3810 1931 3818 2061
rect 3810 1925 3811 1931
rect 3817 1925 3818 1931
rect 3810 1843 3818 1925
rect 3810 1837 3811 1843
rect 3817 1837 3818 1843
rect 3810 1683 3818 1837
rect 3810 1677 3811 1683
rect 3817 1677 3818 1683
rect 3810 1587 3818 1677
rect 3810 1581 3811 1587
rect 3817 1581 3818 1587
rect 3810 1435 3818 1581
rect 3810 1429 3811 1435
rect 3817 1429 3818 1435
rect 3810 1287 3818 1429
rect 3810 1281 3811 1287
rect 3817 1281 3818 1287
rect 3810 1211 3818 1281
rect 3810 1205 3811 1211
rect 3817 1205 3818 1211
rect 3810 1055 3818 1205
rect 3810 1049 3811 1055
rect 3817 1049 3818 1055
rect 3810 935 3818 1049
rect 3810 929 3811 935
rect 3817 929 3818 935
rect 3810 833 3818 929
rect 3810 827 3811 833
rect 3817 827 3818 833
rect 3810 599 3818 827
rect 3810 593 3811 599
rect 3817 593 3818 599
rect 3810 579 3818 593
rect 3810 573 3811 579
rect 3817 573 3818 579
rect 3810 359 3818 573
rect 3810 353 3811 359
rect 3817 353 3818 359
rect 3810 331 3818 353
rect 3810 325 3811 331
rect 3817 325 3818 331
rect 3810 91 3818 325
rect 3810 85 3811 91
rect 3817 85 3818 91
rect 3810 72 3818 85
rect 3822 5691 3830 5760
rect 3822 5685 3823 5691
rect 3829 5685 3830 5691
rect 3822 5471 3830 5685
rect 3822 5465 3823 5471
rect 3829 5465 3830 5471
rect 3822 5463 3830 5465
rect 3822 5457 3823 5463
rect 3829 5457 3830 5463
rect 3822 5235 3830 5457
rect 3822 5229 3823 5235
rect 3829 5229 3830 5235
rect 3822 5223 3830 5229
rect 3822 5217 3823 5223
rect 3829 5217 3830 5223
rect 3822 4987 3830 5217
rect 3822 4981 3823 4987
rect 3829 4981 3830 4987
rect 3822 4743 3830 4981
rect 3822 4737 3823 4743
rect 3829 4737 3830 4743
rect 3822 4691 3830 4737
rect 3822 4685 3823 4691
rect 3829 4685 3830 4691
rect 3822 4503 3830 4685
rect 3822 4497 3823 4503
rect 3829 4497 3830 4503
rect 3822 4463 3830 4497
rect 3822 4457 3823 4463
rect 3829 4457 3830 4463
rect 3822 4263 3830 4457
rect 3822 4257 3823 4263
rect 3829 4257 3830 4263
rect 3822 4211 3830 4257
rect 3822 4205 3823 4211
rect 3829 4205 3830 4211
rect 3822 3963 3830 4205
rect 3822 3957 3823 3963
rect 3829 3957 3830 3963
rect 3822 3935 3830 3957
rect 3822 3929 3823 3935
rect 3829 3929 3830 3935
rect 3822 3703 3830 3929
rect 3822 3697 3823 3703
rect 3829 3697 3830 3703
rect 3822 3691 3830 3697
rect 3822 3685 3823 3691
rect 3829 3685 3830 3691
rect 3822 3467 3830 3685
rect 3822 3461 3823 3467
rect 3829 3461 3830 3467
rect 3822 3411 3830 3461
rect 3822 3405 3823 3411
rect 3829 3405 3830 3411
rect 3822 3219 3830 3405
rect 3822 3213 3823 3219
rect 3829 3213 3830 3219
rect 3822 3171 3830 3213
rect 3822 3165 3823 3171
rect 3829 3165 3830 3171
rect 3822 2995 3830 3165
rect 3822 2989 3823 2995
rect 3829 2989 3830 2995
rect 3822 2923 3830 2989
rect 3822 2917 3823 2923
rect 3829 2917 3830 2923
rect 3822 2719 3830 2917
rect 3822 2713 3823 2719
rect 3829 2713 3830 2719
rect 3822 2683 3830 2713
rect 3822 2677 3823 2683
rect 3829 2677 3830 2683
rect 3822 2475 3830 2677
rect 3822 2469 3823 2475
rect 3829 2469 3830 2475
rect 3822 2439 3830 2469
rect 3822 2433 3823 2439
rect 3829 2433 3830 2439
rect 3822 2243 3830 2433
rect 3822 2237 3823 2243
rect 3829 2237 3830 2243
rect 3822 2199 3830 2237
rect 3822 2193 3823 2199
rect 3829 2193 3830 2199
rect 3822 1955 3830 2193
rect 3822 1949 3823 1955
rect 3829 1949 3830 1955
rect 3822 1807 3830 1949
rect 3822 1801 3823 1807
rect 3829 1801 3830 1807
rect 3822 1715 3830 1801
rect 3822 1709 3823 1715
rect 3829 1709 3830 1715
rect 3822 1559 3830 1709
rect 3822 1553 3823 1559
rect 3829 1553 3830 1559
rect 3822 1403 3830 1553
rect 3822 1397 3823 1403
rect 3829 1397 3830 1403
rect 3822 1323 3830 1397
rect 3822 1317 3823 1323
rect 3829 1317 3830 1323
rect 3822 1167 3830 1317
rect 3822 1161 3823 1167
rect 3829 1161 3830 1167
rect 3822 1075 3830 1161
rect 3822 1069 3823 1075
rect 3829 1069 3830 1075
rect 3822 943 3830 1069
rect 3822 937 3823 943
rect 3829 937 3830 943
rect 3822 823 3830 937
rect 3822 817 3823 823
rect 3829 817 3830 823
rect 3822 711 3830 817
rect 3822 705 3823 711
rect 3829 705 3830 711
rect 3822 475 3830 705
rect 3822 469 3823 475
rect 3829 469 3830 475
rect 3822 467 3830 469
rect 3822 461 3823 467
rect 3829 461 3830 467
rect 3822 203 3830 461
rect 3822 197 3823 203
rect 3829 197 3830 203
rect 3822 72 3830 197
rect 5694 4803 5702 5760
rect 5694 4797 5695 4803
rect 5701 4797 5702 4803
rect 5694 4579 5702 4797
rect 5694 4573 5695 4579
rect 5701 4573 5702 4579
rect 5694 4335 5702 4573
rect 5694 4329 5695 4335
rect 5701 4329 5702 4335
rect 5694 4075 5702 4329
rect 5694 4069 5695 4075
rect 5701 4069 5702 4075
rect 5694 3531 5702 4069
rect 5694 3525 5695 3531
rect 5701 3525 5702 3531
rect 5694 3299 5702 3525
rect 5694 3293 5695 3299
rect 5701 3293 5702 3299
rect 5694 3059 5702 3293
rect 5694 3053 5695 3059
rect 5701 3053 5702 3059
rect 5694 2807 5702 3053
rect 5694 2801 5695 2807
rect 5701 2801 5702 2807
rect 5694 2567 5702 2801
rect 5694 2561 5695 2567
rect 5701 2561 5702 2567
rect 5694 2315 5702 2561
rect 5694 2309 5695 2315
rect 5701 2309 5702 2315
rect 5694 2067 5702 2309
rect 5694 2061 5695 2067
rect 5701 2061 5702 2067
rect 5694 1843 5702 2061
rect 5694 1837 5695 1843
rect 5701 1837 5702 1843
rect 5694 1587 5702 1837
rect 5694 1581 5695 1587
rect 5701 1581 5702 1587
rect 5694 1287 5702 1581
rect 5694 1281 5695 1287
rect 5701 1281 5702 1287
rect 5694 1055 5702 1281
rect 5694 1049 5695 1055
rect 5701 1049 5702 1055
rect 5694 831 5702 1049
rect 5694 825 5695 831
rect 5701 825 5702 831
rect 5694 599 5702 825
rect 5694 593 5695 599
rect 5701 593 5702 599
rect 5694 359 5702 593
rect 5694 353 5695 359
rect 5701 353 5702 359
rect 5694 72 5702 353
rect 5706 5471 5714 5760
rect 5706 5465 5707 5471
rect 5713 5465 5714 5471
rect 5706 5223 5714 5465
rect 5706 5217 5707 5223
rect 5713 5217 5714 5223
rect 5706 4691 5714 5217
rect 5706 4685 5707 4691
rect 5713 4685 5714 4691
rect 5706 4463 5714 4685
rect 5706 4457 5707 4463
rect 5713 4457 5714 4463
rect 5706 4211 5714 4457
rect 5706 4205 5707 4211
rect 5713 4205 5714 4211
rect 5706 3963 5714 4205
rect 5706 3957 5707 3963
rect 5713 3957 5714 3963
rect 5706 3691 5714 3957
rect 5706 3685 5707 3691
rect 5713 3685 5714 3691
rect 5706 3411 5714 3685
rect 5706 3405 5707 3411
rect 5713 3405 5714 3411
rect 5706 3171 5714 3405
rect 5706 3165 5707 3171
rect 5713 3165 5714 3171
rect 5706 2923 5714 3165
rect 5706 2917 5707 2923
rect 5713 2917 5714 2923
rect 5706 2683 5714 2917
rect 5706 2677 5707 2683
rect 5713 2677 5714 2683
rect 5706 2439 5714 2677
rect 5706 2433 5707 2439
rect 5713 2433 5714 2439
rect 5706 2199 5714 2433
rect 5706 2193 5707 2199
rect 5713 2193 5714 2199
rect 5706 1955 5714 2193
rect 5706 1949 5707 1955
rect 5713 1949 5714 1955
rect 5706 1715 5714 1949
rect 5706 1709 5707 1715
rect 5713 1709 5714 1715
rect 5706 1403 5714 1709
rect 5706 1397 5707 1403
rect 5713 1397 5714 1403
rect 5706 1167 5714 1397
rect 5706 1161 5707 1167
rect 5713 1161 5714 1167
rect 5706 943 5714 1161
rect 5706 937 5707 943
rect 5713 937 5714 943
rect 5706 711 5714 937
rect 5706 705 5707 711
rect 5713 705 5714 711
rect 5706 475 5714 705
rect 5706 469 5707 475
rect 5713 469 5714 475
rect 5706 72 5714 469
use circuitwell  npwells
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use circuitppnp  ppnps
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use welltap_svt  __well_tap__269
timestamp 1731220421
transform 1 0 5656 0 1 5604
box 7 3 12 24
use welltap_svt  __well_tap__268
timestamp 1731220421
transform 1 0 3832 0 1 5604
box 7 3 12 24
use welltap_svt  __well_tap__267
timestamp 1731220421
transform 1 0 5656 0 -1 5556
box 7 3 12 24
use welltap_svt  __well_tap__266
timestamp 1731220421
transform 1 0 3832 0 -1 5556
box 7 3 12 24
use welltap_svt  __well_tap__265
timestamp 1731220421
transform 1 0 5656 0 1 5380
box 7 3 12 24
use welltap_svt  __well_tap__264
timestamp 1731220421
transform 1 0 3832 0 1 5380
box 7 3 12 24
use welltap_svt  __well_tap__263
timestamp 1731220421
transform 1 0 5656 0 -1 5324
box 7 3 12 24
use welltap_svt  __well_tap__262
timestamp 1731220421
transform 1 0 3832 0 -1 5324
box 7 3 12 24
use welltap_svt  __well_tap__261
timestamp 1731220421
transform 1 0 5656 0 1 5132
box 7 3 12 24
use welltap_svt  __well_tap__260
timestamp 1731220421
transform 1 0 3832 0 1 5132
box 7 3 12 24
use welltap_svt  __well_tap__259
timestamp 1731220421
transform 1 0 5656 0 -1 5076
box 7 3 12 24
use welltap_svt  __well_tap__258
timestamp 1731220421
transform 1 0 3832 0 -1 5076
box 7 3 12 24
use welltap_svt  __well_tap__257
timestamp 1731220421
transform 1 0 5656 0 1 4900
box 7 3 12 24
use welltap_svt  __well_tap__256
timestamp 1731220421
transform 1 0 3832 0 1 4900
box 7 3 12 24
use welltap_svt  __well_tap__255
timestamp 1731220421
transform 1 0 5656 0 -1 4776
box 7 3 12 24
use welltap_svt  __well_tap__254
timestamp 1731220421
transform 1 0 3832 0 -1 4776
box 7 3 12 24
use welltap_svt  __well_tap__253
timestamp 1731220421
transform 1 0 5656 0 1 4600
box 7 3 12 24
use welltap_svt  __well_tap__252
timestamp 1731220421
transform 1 0 3832 0 1 4600
box 7 3 12 24
use welltap_svt  __well_tap__251
timestamp 1731220421
transform 1 0 5656 0 -1 4552
box 7 3 12 24
use welltap_svt  __well_tap__250
timestamp 1731220421
transform 1 0 3832 0 -1 4552
box 7 3 12 24
use welltap_svt  __well_tap__249
timestamp 1731220421
transform 1 0 5656 0 1 4372
box 7 3 12 24
use welltap_svt  __well_tap__248
timestamp 1731220421
transform 1 0 3832 0 1 4372
box 7 3 12 24
use welltap_svt  __well_tap__247
timestamp 1731220421
transform 1 0 5656 0 -1 4308
box 7 3 12 24
use welltap_svt  __well_tap__246
timestamp 1731220421
transform 1 0 3832 0 -1 4308
box 7 3 12 24
use welltap_svt  __well_tap__245
timestamp 1731220421
transform 1 0 5656 0 1 4120
box 7 3 12 24
use welltap_svt  __well_tap__244
timestamp 1731220421
transform 1 0 3832 0 1 4120
box 7 3 12 24
use welltap_svt  __well_tap__243
timestamp 1731220421
transform 1 0 5656 0 -1 4048
box 7 3 12 24
use welltap_svt  __well_tap__242
timestamp 1731220421
transform 1 0 3832 0 -1 4048
box 7 3 12 24
use welltap_svt  __well_tap__241
timestamp 1731220421
transform 1 0 5656 0 1 3872
box 7 3 12 24
use welltap_svt  __well_tap__240
timestamp 1731220421
transform 1 0 3832 0 1 3872
box 7 3 12 24
use welltap_svt  __well_tap__239
timestamp 1731220421
transform 1 0 5656 0 -1 3796
box 7 3 12 24
use welltap_svt  __well_tap__238
timestamp 1731220421
transform 1 0 3832 0 -1 3796
box 7 3 12 24
use welltap_svt  __well_tap__237
timestamp 1731220421
transform 1 0 5656 0 1 3600
box 7 3 12 24
use welltap_svt  __well_tap__236
timestamp 1731220421
transform 1 0 3832 0 1 3600
box 7 3 12 24
use welltap_svt  __well_tap__235
timestamp 1731220421
transform 1 0 5656 0 -1 3504
box 7 3 12 24
use welltap_svt  __well_tap__234
timestamp 1731220421
transform 1 0 3832 0 -1 3504
box 7 3 12 24
use welltap_svt  __well_tap__233
timestamp 1731220421
transform 1 0 5656 0 1 3320
box 7 3 12 24
use welltap_svt  __well_tap__232
timestamp 1731220421
transform 1 0 3832 0 1 3320
box 7 3 12 24
use welltap_svt  __well_tap__231
timestamp 1731220421
transform 1 0 5656 0 -1 3272
box 7 3 12 24
use welltap_svt  __well_tap__230
timestamp 1731220421
transform 1 0 3832 0 -1 3272
box 7 3 12 24
use welltap_svt  __well_tap__229
timestamp 1731220421
transform 1 0 5656 0 1 3080
box 7 3 12 24
use welltap_svt  __well_tap__228
timestamp 1731220421
transform 1 0 3832 0 1 3080
box 7 3 12 24
use welltap_svt  __well_tap__227
timestamp 1731220421
transform 1 0 5656 0 -1 3032
box 7 3 12 24
use welltap_svt  __well_tap__226
timestamp 1731220421
transform 1 0 3832 0 -1 3032
box 7 3 12 24
use welltap_svt  __well_tap__225
timestamp 1731220421
transform 1 0 5656 0 1 2832
box 7 3 12 24
use welltap_svt  __well_tap__224
timestamp 1731220421
transform 1 0 3832 0 1 2832
box 7 3 12 24
use welltap_svt  __well_tap__223
timestamp 1731220421
transform 1 0 5656 0 -1 2780
box 7 3 12 24
use welltap_svt  __well_tap__222
timestamp 1731220421
transform 1 0 3832 0 -1 2780
box 7 3 12 24
use welltap_svt  __well_tap__221
timestamp 1731220421
transform 1 0 5656 0 1 2592
box 7 3 12 24
use welltap_svt  __well_tap__220
timestamp 1731220421
transform 1 0 3832 0 1 2592
box 7 3 12 24
use welltap_svt  __well_tap__219
timestamp 1731220421
transform 1 0 5656 0 -1 2540
box 7 3 12 24
use welltap_svt  __well_tap__218
timestamp 1731220421
transform 1 0 3832 0 -1 2540
box 7 3 12 24
use welltap_svt  __well_tap__217
timestamp 1731220421
transform 1 0 5656 0 1 2348
box 7 3 12 24
use welltap_svt  __well_tap__216
timestamp 1731220421
transform 1 0 3832 0 1 2348
box 7 3 12 24
use welltap_svt  __well_tap__215
timestamp 1731220421
transform 1 0 5656 0 -1 2288
box 7 3 12 24
use welltap_svt  __well_tap__214
timestamp 1731220421
transform 1 0 3832 0 -1 2288
box 7 3 12 24
use welltap_svt  __well_tap__213
timestamp 1731220421
transform 1 0 5656 0 1 2108
box 7 3 12 24
use welltap_svt  __well_tap__212
timestamp 1731220421
transform 1 0 3832 0 1 2108
box 7 3 12 24
use welltap_svt  __well_tap__211
timestamp 1731220421
transform 1 0 5656 0 -1 2040
box 7 3 12 24
use welltap_svt  __well_tap__210
timestamp 1731220421
transform 1 0 3832 0 -1 2040
box 7 3 12 24
use welltap_svt  __well_tap__209
timestamp 1731220421
transform 1 0 5656 0 1 1864
box 7 3 12 24
use welltap_svt  __well_tap__208
timestamp 1731220421
transform 1 0 3832 0 1 1864
box 7 3 12 24
use welltap_svt  __well_tap__207
timestamp 1731220421
transform 1 0 5656 0 -1 1816
box 7 3 12 24
use welltap_svt  __well_tap__206
timestamp 1731220421
transform 1 0 3832 0 -1 1816
box 7 3 12 24
use welltap_svt  __well_tap__205
timestamp 1731220421
transform 1 0 5656 0 1 1624
box 7 3 12 24
use welltap_svt  __well_tap__204
timestamp 1731220421
transform 1 0 3832 0 1 1624
box 7 3 12 24
use welltap_svt  __well_tap__203
timestamp 1731220421
transform 1 0 5656 0 -1 1560
box 7 3 12 24
use welltap_svt  __well_tap__202
timestamp 1731220421
transform 1 0 3832 0 -1 1560
box 7 3 12 24
use welltap_svt  __well_tap__201
timestamp 1731220421
transform 1 0 5656 0 1 1312
box 7 3 12 24
use welltap_svt  __well_tap__200
timestamp 1731220421
transform 1 0 3832 0 1 1312
box 7 3 12 24
use welltap_svt  __well_tap__199
timestamp 1731220421
transform 1 0 5656 0 -1 1260
box 7 3 12 24
use welltap_svt  __well_tap__198
timestamp 1731220421
transform 1 0 3832 0 -1 1260
box 7 3 12 24
use welltap_svt  __well_tap__197
timestamp 1731220421
transform 1 0 5656 0 1 1076
box 7 3 12 24
use welltap_svt  __well_tap__196
timestamp 1731220421
transform 1 0 3832 0 1 1076
box 7 3 12 24
use welltap_svt  __well_tap__195
timestamp 1731220421
transform 1 0 5656 0 -1 1028
box 7 3 12 24
use welltap_svt  __well_tap__194
timestamp 1731220421
transform 1 0 3832 0 -1 1028
box 7 3 12 24
use welltap_svt  __well_tap__193
timestamp 1731220421
transform 1 0 5656 0 1 852
box 7 3 12 24
use welltap_svt  __well_tap__192
timestamp 1731220421
transform 1 0 3832 0 1 852
box 7 3 12 24
use welltap_svt  __well_tap__191
timestamp 1731220421
transform 1 0 5656 0 -1 804
box 7 3 12 24
use welltap_svt  __well_tap__190
timestamp 1731220421
transform 1 0 3832 0 -1 804
box 7 3 12 24
use welltap_svt  __well_tap__189
timestamp 1731220421
transform 1 0 5656 0 1 620
box 7 3 12 24
use welltap_svt  __well_tap__188
timestamp 1731220421
transform 1 0 3832 0 1 620
box 7 3 12 24
use welltap_svt  __well_tap__187
timestamp 1731220421
transform 1 0 5656 0 -1 572
box 7 3 12 24
use welltap_svt  __well_tap__186
timestamp 1731220421
transform 1 0 3832 0 -1 572
box 7 3 12 24
use welltap_svt  __well_tap__185
timestamp 1731220421
transform 1 0 5656 0 1 384
box 7 3 12 24
use welltap_svt  __well_tap__184
timestamp 1731220421
transform 1 0 3832 0 1 384
box 7 3 12 24
use welltap_svt  __well_tap__183
timestamp 1731220421
transform 1 0 5656 0 -1 332
box 7 3 12 24
use welltap_svt  __well_tap__182
timestamp 1731220421
transform 1 0 3832 0 -1 332
box 7 3 12 24
use welltap_svt  __well_tap__181
timestamp 1731220421
transform 1 0 5656 0 1 116
box 7 3 12 24
use welltap_svt  __well_tap__180
timestamp 1731220421
transform 1 0 3832 0 1 116
box 7 3 12 24
use welltap_svt  __well_tap__179
timestamp 1731220421
transform 1 0 3792 0 1 5600
box 7 3 12 24
use welltap_svt  __well_tap__178
timestamp 1731220421
transform 1 0 1968 0 1 5600
box 7 3 12 24
use welltap_svt  __well_tap__177
timestamp 1731220421
transform 1 0 3792 0 -1 5552
box 7 3 12 24
use welltap_svt  __well_tap__176
timestamp 1731220421
transform 1 0 1968 0 -1 5552
box 7 3 12 24
use welltap_svt  __well_tap__175
timestamp 1731220421
transform 1 0 3792 0 1 5372
box 7 3 12 24
use welltap_svt  __well_tap__174
timestamp 1731220421
transform 1 0 1968 0 1 5372
box 7 3 12 24
use welltap_svt  __well_tap__173
timestamp 1731220421
transform 1 0 3792 0 -1 5324
box 7 3 12 24
use welltap_svt  __well_tap__172
timestamp 1731220421
transform 1 0 1968 0 -1 5324
box 7 3 12 24
use welltap_svt  __well_tap__171
timestamp 1731220421
transform 1 0 3792 0 1 5144
box 7 3 12 24
use welltap_svt  __well_tap__170
timestamp 1731220421
transform 1 0 1968 0 1 5144
box 7 3 12 24
use welltap_svt  __well_tap__169
timestamp 1731220421
transform 1 0 3792 0 -1 5080
box 7 3 12 24
use welltap_svt  __well_tap__168
timestamp 1731220421
transform 1 0 1968 0 -1 5080
box 7 3 12 24
use welltap_svt  __well_tap__167
timestamp 1731220421
transform 1 0 3792 0 1 4896
box 7 3 12 24
use welltap_svt  __well_tap__166
timestamp 1731220421
transform 1 0 1968 0 1 4896
box 7 3 12 24
use welltap_svt  __well_tap__165
timestamp 1731220421
transform 1 0 3792 0 -1 4840
box 7 3 12 24
use welltap_svt  __well_tap__164
timestamp 1731220421
transform 1 0 1968 0 -1 4840
box 7 3 12 24
use welltap_svt  __well_tap__163
timestamp 1731220421
transform 1 0 3792 0 1 4652
box 7 3 12 24
use welltap_svt  __well_tap__162
timestamp 1731220421
transform 1 0 1968 0 1 4652
box 7 3 12 24
use welltap_svt  __well_tap__161
timestamp 1731220421
transform 1 0 3792 0 -1 4600
box 7 3 12 24
use welltap_svt  __well_tap__160
timestamp 1731220421
transform 1 0 1968 0 -1 4600
box 7 3 12 24
use welltap_svt  __well_tap__159
timestamp 1731220421
transform 1 0 3792 0 1 4412
box 7 3 12 24
use welltap_svt  __well_tap__158
timestamp 1731220421
transform 1 0 1968 0 1 4412
box 7 3 12 24
use welltap_svt  __well_tap__157
timestamp 1731220421
transform 1 0 3792 0 -1 4352
box 7 3 12 24
use welltap_svt  __well_tap__156
timestamp 1731220421
transform 1 0 1968 0 -1 4352
box 7 3 12 24
use welltap_svt  __well_tap__155
timestamp 1731220421
transform 1 0 3792 0 1 4172
box 7 3 12 24
use welltap_svt  __well_tap__154
timestamp 1731220421
transform 1 0 1968 0 1 4172
box 7 3 12 24
use welltap_svt  __well_tap__153
timestamp 1731220421
transform 1 0 3792 0 -1 4112
box 7 3 12 24
use welltap_svt  __well_tap__152
timestamp 1731220421
transform 1 0 1968 0 -1 4112
box 7 3 12 24
use welltap_svt  __well_tap__151
timestamp 1731220421
transform 1 0 3792 0 1 3844
box 7 3 12 24
use welltap_svt  __well_tap__150
timestamp 1731220421
transform 1 0 1968 0 1 3844
box 7 3 12 24
use welltap_svt  __well_tap__149
timestamp 1731220421
transform 1 0 3792 0 -1 3796
box 7 3 12 24
use welltap_svt  __well_tap__148
timestamp 1731220421
transform 1 0 1968 0 -1 3796
box 7 3 12 24
use welltap_svt  __well_tap__147
timestamp 1731220421
transform 1 0 3792 0 1 3612
box 7 3 12 24
use welltap_svt  __well_tap__146
timestamp 1731220421
transform 1 0 1968 0 1 3612
box 7 3 12 24
use welltap_svt  __well_tap__145
timestamp 1731220421
transform 1 0 3792 0 -1 3556
box 7 3 12 24
use welltap_svt  __well_tap__144
timestamp 1731220421
transform 1 0 1968 0 -1 3556
box 7 3 12 24
use welltap_svt  __well_tap__143
timestamp 1731220421
transform 1 0 3792 0 1 3376
box 7 3 12 24
use welltap_svt  __well_tap__142
timestamp 1731220421
transform 1 0 1968 0 1 3376
box 7 3 12 24
use welltap_svt  __well_tap__141
timestamp 1731220421
transform 1 0 3792 0 -1 3304
box 7 3 12 24
use welltap_svt  __well_tap__140
timestamp 1731220421
transform 1 0 1968 0 -1 3304
box 7 3 12 24
use welltap_svt  __well_tap__139
timestamp 1731220421
transform 1 0 3792 0 1 3128
box 7 3 12 24
use welltap_svt  __well_tap__138
timestamp 1731220421
transform 1 0 1968 0 1 3128
box 7 3 12 24
use welltap_svt  __well_tap__137
timestamp 1731220421
transform 1 0 3792 0 -1 3080
box 7 3 12 24
use welltap_svt  __well_tap__136
timestamp 1731220421
transform 1 0 1968 0 -1 3080
box 7 3 12 24
use welltap_svt  __well_tap__135
timestamp 1731220421
transform 1 0 3792 0 1 2904
box 7 3 12 24
use welltap_svt  __well_tap__134
timestamp 1731220421
transform 1 0 1968 0 1 2904
box 7 3 12 24
use welltap_svt  __well_tap__133
timestamp 1731220421
transform 1 0 3792 0 -1 2804
box 7 3 12 24
use welltap_svt  __well_tap__132
timestamp 1731220421
transform 1 0 1968 0 -1 2804
box 7 3 12 24
use welltap_svt  __well_tap__131
timestamp 1731220421
transform 1 0 3792 0 1 2628
box 7 3 12 24
use welltap_svt  __well_tap__130
timestamp 1731220421
transform 1 0 1968 0 1 2628
box 7 3 12 24
use welltap_svt  __well_tap__129
timestamp 1731220421
transform 1 0 3792 0 -1 2576
box 7 3 12 24
use welltap_svt  __well_tap__128
timestamp 1731220421
transform 1 0 1968 0 -1 2576
box 7 3 12 24
use welltap_svt  __well_tap__127
timestamp 1731220421
transform 1 0 3792 0 1 2384
box 7 3 12 24
use welltap_svt  __well_tap__126
timestamp 1731220421
transform 1 0 1968 0 1 2384
box 7 3 12 24
use welltap_svt  __well_tap__125
timestamp 1731220421
transform 1 0 3792 0 -1 2328
box 7 3 12 24
use welltap_svt  __well_tap__124
timestamp 1731220421
transform 1 0 1968 0 -1 2328
box 7 3 12 24
use welltap_svt  __well_tap__123
timestamp 1731220421
transform 1 0 3792 0 1 2152
box 7 3 12 24
use welltap_svt  __well_tap__122
timestamp 1731220421
transform 1 0 1968 0 1 2152
box 7 3 12 24
use welltap_svt  __well_tap__121
timestamp 1731220421
transform 1 0 3792 0 -1 1904
box 7 3 12 24
use welltap_svt  __well_tap__120
timestamp 1731220421
transform 1 0 1968 0 -1 1904
box 7 3 12 24
use welltap_svt  __well_tap__119
timestamp 1731220421
transform 1 0 3792 0 1 1716
box 7 3 12 24
use welltap_svt  __well_tap__118
timestamp 1731220421
transform 1 0 1968 0 1 1716
box 7 3 12 24
use welltap_svt  __well_tap__117
timestamp 1731220421
transform 1 0 3792 0 -1 1656
box 7 3 12 24
use welltap_svt  __well_tap__116
timestamp 1731220421
transform 1 0 1968 0 -1 1656
box 7 3 12 24
use welltap_svt  __well_tap__115
timestamp 1731220421
transform 1 0 3792 0 1 1468
box 7 3 12 24
use welltap_svt  __well_tap__114
timestamp 1731220421
transform 1 0 1968 0 1 1468
box 7 3 12 24
use welltap_svt  __well_tap__113
timestamp 1731220421
transform 1 0 3792 0 -1 1408
box 7 3 12 24
use welltap_svt  __well_tap__112
timestamp 1731220421
transform 1 0 1968 0 -1 1408
box 7 3 12 24
use welltap_svt  __well_tap__111
timestamp 1731220421
transform 1 0 3792 0 1 1232
box 7 3 12 24
use welltap_svt  __well_tap__110
timestamp 1731220421
transform 1 0 1968 0 1 1232
box 7 3 12 24
use welltap_svt  __well_tap__109
timestamp 1731220421
transform 1 0 3792 0 -1 1184
box 7 3 12 24
use welltap_svt  __well_tap__108
timestamp 1731220421
transform 1 0 1968 0 -1 1184
box 7 3 12 24
use welltap_svt  __well_tap__107
timestamp 1731220421
transform 1 0 3792 0 1 984
box 7 3 12 24
use welltap_svt  __well_tap__106
timestamp 1731220421
transform 1 0 1968 0 1 984
box 7 3 12 24
use welltap_svt  __well_tap__105
timestamp 1731220421
transform 1 0 3792 0 -1 908
box 7 3 12 24
use welltap_svt  __well_tap__104
timestamp 1731220421
transform 1 0 1968 0 -1 908
box 7 3 12 24
use welltap_svt  __well_tap__103
timestamp 1731220421
transform 1 0 3792 0 1 732
box 7 3 12 24
use welltap_svt  __well_tap__102
timestamp 1731220421
transform 1 0 1968 0 1 732
box 7 3 12 24
use welltap_svt  __well_tap__101
timestamp 1731220421
transform 1 0 3792 0 -1 552
box 7 3 12 24
use welltap_svt  __well_tap__100
timestamp 1731220421
transform 1 0 1968 0 -1 552
box 7 3 12 24
use welltap_svt  __well_tap__99
timestamp 1731220421
transform 1 0 3792 0 1 376
box 7 3 12 24
use welltap_svt  __well_tap__98
timestamp 1731220421
transform 1 0 1968 0 1 376
box 7 3 12 24
use welltap_svt  __well_tap__97
timestamp 1731220421
transform 1 0 3792 0 -1 304
box 7 3 12 24
use welltap_svt  __well_tap__96
timestamp 1731220421
transform 1 0 1968 0 -1 304
box 7 3 12 24
use welltap_svt  __well_tap__95
timestamp 1731220421
transform 1 0 3792 0 1 112
box 7 3 12 24
use welltap_svt  __well_tap__94
timestamp 1731220421
transform 1 0 1968 0 1 112
box 7 3 12 24
use welltap_svt  __well_tap__93
timestamp 1731220421
transform 1 0 1928 0 1 5668
box 7 3 12 24
use welltap_svt  __well_tap__92
timestamp 1731220421
transform 1 0 104 0 1 5668
box 7 3 12 24
use welltap_svt  __well_tap__91
timestamp 1731220421
transform 1 0 1928 0 -1 5620
box 7 3 12 24
use welltap_svt  __well_tap__90
timestamp 1731220421
transform 1 0 104 0 -1 5620
box 7 3 12 24
use welltap_svt  __well_tap__89
timestamp 1731220421
transform 1 0 1928 0 1 5444
box 7 3 12 24
use welltap_svt  __well_tap__88
timestamp 1731220421
transform 1 0 104 0 1 5444
box 7 3 12 24
use welltap_svt  __well_tap__87
timestamp 1731220421
transform 1 0 1928 0 -1 5396
box 7 3 12 24
use welltap_svt  __well_tap__86
timestamp 1731220421
transform 1 0 104 0 -1 5396
box 7 3 12 24
use welltap_svt  __well_tap__85
timestamp 1731220421
transform 1 0 1928 0 1 5220
box 7 3 12 24
use welltap_svt  __well_tap__84
timestamp 1731220421
transform 1 0 104 0 1 5220
box 7 3 12 24
use welltap_svt  __well_tap__83
timestamp 1731220421
transform 1 0 1928 0 -1 5172
box 7 3 12 24
use welltap_svt  __well_tap__82
timestamp 1731220421
transform 1 0 104 0 -1 5172
box 7 3 12 24
use welltap_svt  __well_tap__81
timestamp 1731220421
transform 1 0 1928 0 1 4988
box 7 3 12 24
use welltap_svt  __well_tap__80
timestamp 1731220421
transform 1 0 104 0 1 4988
box 7 3 12 24
use welltap_svt  __well_tap__79
timestamp 1731220421
transform 1 0 1928 0 -1 4912
box 7 3 12 24
use welltap_svt  __well_tap__78
timestamp 1731220421
transform 1 0 104 0 -1 4912
box 7 3 12 24
use welltap_svt  __well_tap__77
timestamp 1731220421
transform 1 0 1928 0 1 4724
box 7 3 12 24
use welltap_svt  __well_tap__76
timestamp 1731220421
transform 1 0 104 0 1 4724
box 7 3 12 24
use welltap_svt  __well_tap__75
timestamp 1731220421
transform 1 0 1928 0 -1 4672
box 7 3 12 24
use welltap_svt  __well_tap__74
timestamp 1731220421
transform 1 0 104 0 -1 4672
box 7 3 12 24
use welltap_svt  __well_tap__73
timestamp 1731220421
transform 1 0 1928 0 1 4484
box 7 3 12 24
use welltap_svt  __well_tap__72
timestamp 1731220421
transform 1 0 104 0 1 4484
box 7 3 12 24
use welltap_svt  __well_tap__71
timestamp 1731220421
transform 1 0 1928 0 -1 4436
box 7 3 12 24
use welltap_svt  __well_tap__70
timestamp 1731220421
transform 1 0 104 0 -1 4436
box 7 3 12 24
use welltap_svt  __well_tap__69
timestamp 1731220421
transform 1 0 1928 0 1 4256
box 7 3 12 24
use welltap_svt  __well_tap__68
timestamp 1731220421
transform 1 0 104 0 1 4256
box 7 3 12 24
use welltap_svt  __well_tap__67
timestamp 1731220421
transform 1 0 1928 0 -1 4200
box 7 3 12 24
use welltap_svt  __well_tap__66
timestamp 1731220421
transform 1 0 104 0 -1 4200
box 7 3 12 24
use welltap_svt  __well_tap__65
timestamp 1731220421
transform 1 0 1928 0 1 4024
box 7 3 12 24
use welltap_svt  __well_tap__64
timestamp 1731220421
transform 1 0 104 0 1 4024
box 7 3 12 24
use welltap_svt  __well_tap__63
timestamp 1731220421
transform 1 0 1928 0 -1 3976
box 7 3 12 24
use welltap_svt  __well_tap__62
timestamp 1731220421
transform 1 0 104 0 -1 3976
box 7 3 12 24
use welltap_svt  __well_tap__61
timestamp 1731220421
transform 1 0 1928 0 1 3800
box 7 3 12 24
use welltap_svt  __well_tap__60
timestamp 1731220421
transform 1 0 104 0 1 3800
box 7 3 12 24
use welltap_svt  __well_tap__59
timestamp 1731220421
transform 1 0 1928 0 -1 3740
box 7 3 12 24
use welltap_svt  __well_tap__58
timestamp 1731220421
transform 1 0 104 0 -1 3740
box 7 3 12 24
use welltap_svt  __well_tap__57
timestamp 1731220421
transform 1 0 1928 0 1 3548
box 7 3 12 24
use welltap_svt  __well_tap__56
timestamp 1731220421
transform 1 0 104 0 1 3548
box 7 3 12 24
use welltap_svt  __well_tap__55
timestamp 1731220421
transform 1 0 1928 0 -1 3480
box 7 3 12 24
use welltap_svt  __well_tap__54
timestamp 1731220421
transform 1 0 104 0 -1 3480
box 7 3 12 24
use welltap_svt  __well_tap__53
timestamp 1731220421
transform 1 0 1928 0 1 3296
box 7 3 12 24
use welltap_svt  __well_tap__52
timestamp 1731220421
transform 1 0 104 0 1 3296
box 7 3 12 24
use welltap_svt  __well_tap__51
timestamp 1731220421
transform 1 0 1928 0 -1 3240
box 7 3 12 24
use welltap_svt  __well_tap__50
timestamp 1731220421
transform 1 0 104 0 -1 3240
box 7 3 12 24
use welltap_svt  __well_tap__49
timestamp 1731220421
transform 1 0 1928 0 1 3048
box 7 3 12 24
use welltap_svt  __well_tap__48
timestamp 1731220421
transform 1 0 104 0 1 3048
box 7 3 12 24
use welltap_svt  __well_tap__47
timestamp 1731220421
transform 1 0 1928 0 -1 3000
box 7 3 12 24
use welltap_svt  __well_tap__46
timestamp 1731220421
transform 1 0 104 0 -1 3000
box 7 3 12 24
use welltap_svt  __well_tap__45
timestamp 1731220421
transform 1 0 1928 0 1 2820
box 7 3 12 24
use welltap_svt  __well_tap__44
timestamp 1731220421
transform 1 0 104 0 1 2820
box 7 3 12 24
use welltap_svt  __well_tap__43
timestamp 1731220421
transform 1 0 1928 0 -1 2760
box 7 3 12 24
use welltap_svt  __well_tap__42
timestamp 1731220421
transform 1 0 104 0 -1 2760
box 7 3 12 24
use welltap_svt  __well_tap__41
timestamp 1731220421
transform 1 0 1928 0 1 2584
box 7 3 12 24
use welltap_svt  __well_tap__40
timestamp 1731220421
transform 1 0 104 0 1 2584
box 7 3 12 24
use welltap_svt  __well_tap__39
timestamp 1731220421
transform 1 0 1928 0 -1 2520
box 7 3 12 24
use welltap_svt  __well_tap__38
timestamp 1731220421
transform 1 0 104 0 -1 2520
box 7 3 12 24
use welltap_svt  __well_tap__37
timestamp 1731220421
transform 1 0 1928 0 1 2332
box 7 3 12 24
use welltap_svt  __well_tap__36
timestamp 1731220421
transform 1 0 104 0 1 2332
box 7 3 12 24
use welltap_svt  __well_tap__35
timestamp 1731220421
transform 1 0 1928 0 -1 2280
box 7 3 12 24
use welltap_svt  __well_tap__34
timestamp 1731220421
transform 1 0 104 0 -1 2280
box 7 3 12 24
use welltap_svt  __well_tap__33
timestamp 1731220421
transform 1 0 1928 0 1 2080
box 7 3 12 24
use welltap_svt  __well_tap__32
timestamp 1731220421
transform 1 0 104 0 1 2080
box 7 3 12 24
use welltap_svt  __well_tap__31
timestamp 1731220421
transform 1 0 1928 0 -1 2028
box 7 3 12 24
use welltap_svt  __well_tap__30
timestamp 1731220421
transform 1 0 104 0 -1 2028
box 7 3 12 24
use welltap_svt  __well_tap__29
timestamp 1731220421
transform 1 0 1928 0 1 1840
box 7 3 12 24
use welltap_svt  __well_tap__28
timestamp 1731220421
transform 1 0 104 0 1 1840
box 7 3 12 24
use welltap_svt  __well_tap__27
timestamp 1731220421
transform 1 0 1928 0 -1 1780
box 7 3 12 24
use welltap_svt  __well_tap__26
timestamp 1731220421
transform 1 0 104 0 -1 1780
box 7 3 12 24
use welltap_svt  __well_tap__25
timestamp 1731220421
transform 1 0 1928 0 1 1592
box 7 3 12 24
use welltap_svt  __well_tap__24
timestamp 1731220421
transform 1 0 104 0 1 1592
box 7 3 12 24
use welltap_svt  __well_tap__23
timestamp 1731220421
transform 1 0 1928 0 -1 1532
box 7 3 12 24
use welltap_svt  __well_tap__22
timestamp 1731220421
transform 1 0 104 0 -1 1532
box 7 3 12 24
use welltap_svt  __well_tap__21
timestamp 1731220421
transform 1 0 1928 0 1 1344
box 7 3 12 24
use welltap_svt  __well_tap__20
timestamp 1731220421
transform 1 0 104 0 1 1344
box 7 3 12 24
use welltap_svt  __well_tap__19
timestamp 1731220421
transform 1 0 1928 0 -1 1296
box 7 3 12 24
use welltap_svt  __well_tap__18
timestamp 1731220421
transform 1 0 104 0 -1 1296
box 7 3 12 24
use welltap_svt  __well_tap__17
timestamp 1731220421
transform 1 0 1928 0 1 1096
box 7 3 12 24
use welltap_svt  __well_tap__16
timestamp 1731220421
transform 1 0 104 0 1 1096
box 7 3 12 24
use welltap_svt  __well_tap__15
timestamp 1731220421
transform 1 0 1928 0 -1 1048
box 7 3 12 24
use welltap_svt  __well_tap__14
timestamp 1731220421
transform 1 0 104 0 -1 1048
box 7 3 12 24
use welltap_svt  __well_tap__13
timestamp 1731220421
transform 1 0 1928 0 1 868
box 7 3 12 24
use welltap_svt  __well_tap__12
timestamp 1731220421
transform 1 0 104 0 1 868
box 7 3 12 24
use welltap_svt  __well_tap__11
timestamp 1731220421
transform 1 0 1928 0 -1 804
box 7 3 12 24
use welltap_svt  __well_tap__10
timestamp 1731220421
transform 1 0 104 0 -1 804
box 7 3 12 24
use welltap_svt  __well_tap__9
timestamp 1731220421
transform 1 0 1928 0 1 628
box 7 3 12 24
use welltap_svt  __well_tap__8
timestamp 1731220421
transform 1 0 104 0 1 628
box 7 3 12 24
use welltap_svt  __well_tap__7
timestamp 1731220421
transform 1 0 1928 0 -1 580
box 7 3 12 24
use welltap_svt  __well_tap__6
timestamp 1731220421
transform 1 0 104 0 -1 580
box 7 3 12 24
use welltap_svt  __well_tap__5
timestamp 1731220421
transform 1 0 1928 0 1 404
box 7 3 12 24
use welltap_svt  __well_tap__4
timestamp 1731220421
transform 1 0 104 0 1 404
box 7 3 12 24
use welltap_svt  __well_tap__3
timestamp 1731220421
transform 1 0 1928 0 -1 340
box 7 3 12 24
use welltap_svt  __well_tap__2
timestamp 1731220421
transform 1 0 104 0 -1 340
box 7 3 12 24
use welltap_svt  __well_tap__1
timestamp 1731220421
transform 1 0 1928 0 1 132
box 7 3 12 24
use welltap_svt  __well_tap__0
timestamp 1731220421
transform 1 0 104 0 1 132
box 7 3 12 24
use _0_0std_0_0cells_0_0FAX1  tst_5999_6
timestamp 1731220421
transform 1 0 5376 0 1 92
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5998_6
timestamp 1731220421
transform 1 0 5512 0 1 92
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5997_6
timestamp 1731220421
transform 1 0 5512 0 -1 356
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5996_6
timestamp 1731220421
transform 1 0 5504 0 1 360
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5995_6
timestamp 1731220421
transform 1 0 5456 0 1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5994_6
timestamp 1731220421
transform 1 0 5416 0 -1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5993_6
timestamp 1731220421
transform 1 0 5280 0 1 360
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5992_6
timestamp 1731220421
transform 1 0 5200 0 -1 356
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5991_6
timestamp 1731220421
transform 1 0 5040 0 -1 356
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5990_6
timestamp 1731220421
transform 1 0 5368 0 -1 356
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5989_6
timestamp 1731220421
transform 1 0 5240 0 1 92
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5988_6
timestamp 1731220421
transform 1 0 5104 0 1 92
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5987_6
timestamp 1731220421
transform 1 0 4968 0 1 92
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5986_6
timestamp 1731220421
transform 1 0 4832 0 1 92
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5985_6
timestamp 1731220421
transform 1 0 4696 0 1 92
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5984_6
timestamp 1731220421
transform 1 0 4560 0 1 92
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5983_6
timestamp 1731220421
transform 1 0 4424 0 1 92
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5982_6
timestamp 1731220421
transform 1 0 4288 0 1 92
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5981_6
timestamp 1731220421
transform 1 0 4720 0 -1 356
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5980_6
timestamp 1731220421
transform 1 0 4880 0 -1 356
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5979_6
timestamp 1731220421
transform 1 0 5064 0 1 360
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5978_6
timestamp 1731220421
transform 1 0 4856 0 1 360
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5977_6
timestamp 1731220421
transform 1 0 4648 0 1 360
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5976_6
timestamp 1731220421
transform 1 0 4448 0 1 360
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5975_6
timestamp 1731220421
transform 1 0 5160 0 -1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5974_6
timestamp 1731220421
transform 1 0 4904 0 -1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5973_6
timestamp 1731220421
transform 1 0 4664 0 -1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5972_6
timestamp 1731220421
transform 1 0 4448 0 -1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5971_6
timestamp 1731220421
transform 1 0 4264 0 -1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5970_6
timestamp 1731220421
transform 1 0 5224 0 1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5969_6
timestamp 1731220421
transform 1 0 4992 0 1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5968_6
timestamp 1731220421
transform 1 0 4768 0 1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5967_6
timestamp 1731220421
transform 1 0 4568 0 1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5966_6
timestamp 1731220421
transform 1 0 4248 0 -1 828
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5965_6
timestamp 1731220421
transform 1 0 3968 0 1 828
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5964_6
timestamp 1731220421
transform 1 0 3856 0 -1 1052
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5963_6
timestamp 1731220421
transform 1 0 4040 0 -1 1052
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5962_6
timestamp 1731220421
transform 1 0 4064 0 1 1052
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5961_6
timestamp 1731220421
transform 1 0 3856 0 1 1052
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5960_6
timestamp 1731220421
transform 1 0 3648 0 -1 1208
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5959_6
timestamp 1731220421
transform 1 0 3648 0 1 1208
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5958_6
timestamp 1731220421
transform 1 0 3464 0 1 1208
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5957_6
timestamp 1731220421
transform 1 0 3424 0 -1 1208
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5956_6
timestamp 1731220421
transform 1 0 3176 0 -1 1208
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5955_6
timestamp 1731220421
transform 1 0 3392 0 1 960
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5954_6
timestamp 1731220421
transform 1 0 3240 0 1 960
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5953_6
timestamp 1731220421
transform 1 0 3176 0 -1 932
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5952_6
timestamp 1731220421
transform 1 0 3464 0 -1 932
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5951_6
timestamp 1731220421
transform 1 0 3448 0 1 708
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5950_6
timestamp 1731220421
transform 1 0 3224 0 1 708
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5949_6
timestamp 1731220421
transform 1 0 3648 0 1 708
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5948_6
timestamp 1731220421
transform 1 0 3856 0 1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5947_6
timestamp 1731220421
transform 1 0 3856 0 -1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5946_6
timestamp 1731220421
transform 1 0 3992 0 -1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5945_6
timestamp 1731220421
transform 1 0 4128 0 -1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5944_6
timestamp 1731220421
transform 1 0 4400 0 1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5943_6
timestamp 1731220421
transform 1 0 4264 0 1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5942_6
timestamp 1731220421
transform 1 0 4128 0 1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5941_6
timestamp 1731220421
transform 1 0 3992 0 1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5940_6
timestamp 1731220421
transform 1 0 3856 0 -1 828
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5939_6
timestamp 1731220421
transform 1 0 4016 0 -1 828
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5938_6
timestamp 1731220421
transform 1 0 5192 0 -1 828
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5937_6
timestamp 1731220421
transform 1 0 4848 0 -1 828
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5936_6
timestamp 1731220421
transform 1 0 4528 0 -1 828
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5935_6
timestamp 1731220421
transform 1 0 4400 0 1 828
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5934_6
timestamp 1731220421
transform 1 0 4176 0 1 828
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5933_6
timestamp 1731220421
transform 1 0 4896 0 1 828
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5932_6
timestamp 1731220421
transform 1 0 4640 0 1 828
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5931_6
timestamp 1731220421
transform 1 0 4480 0 -1 1052
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5930_6
timestamp 1731220421
transform 1 0 4248 0 -1 1052
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5929_6
timestamp 1731220421
transform 1 0 4992 0 -1 1052
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5928_6
timestamp 1731220421
transform 1 0 4728 0 -1 1052
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5927_6
timestamp 1731220421
transform 1 0 4536 0 1 1052
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5926_6
timestamp 1731220421
transform 1 0 4296 0 1 1052
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5925_6
timestamp 1731220421
transform 1 0 5024 0 1 1052
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5924_6
timestamp 1731220421
transform 1 0 4776 0 1 1052
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5923_6
timestamp 1731220421
transform 1 0 4704 0 -1 1284
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5922_6
timestamp 1731220421
transform 1 0 5000 0 -1 1284
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5921_6
timestamp 1731220421
transform 1 0 4848 0 -1 1284
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5920_6
timestamp 1731220421
transform 1 0 4808 0 1 1288
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5919_6
timestamp 1731220421
transform 1 0 4944 0 1 1288
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5918_6
timestamp 1731220421
transform 1 0 5080 0 1 1288
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5917_6
timestamp 1731220421
transform 1 0 5216 0 1 1288
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5916_6
timestamp 1731220421
transform 1 0 5160 0 -1 1284
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5915_6
timestamp 1731220421
transform 1 0 5328 0 -1 1284
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5914_6
timestamp 1731220421
transform 1 0 5280 0 1 1052
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5913_6
timestamp 1731220421
transform 1 0 5264 0 -1 1052
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5912_6
timestamp 1731220421
transform 1 0 5168 0 1 828
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5911_6
timestamp 1731220421
transform 1 0 5440 0 1 828
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5910_6
timestamp 1731220421
transform 1 0 5512 0 -1 828
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5909_6
timestamp 1731220421
transform 1 0 5512 0 -1 1052
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5908_6
timestamp 1731220421
transform 1 0 5512 0 1 1052
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5907_6
timestamp 1731220421
transform 1 0 5496 0 -1 1284
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5906_6
timestamp 1731220421
transform 1 0 5488 0 1 1288
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5905_6
timestamp 1731220421
transform 1 0 5352 0 1 1288
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5904_6
timestamp 1731220421
transform 1 0 5512 0 -1 1584
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5903_6
timestamp 1731220421
transform 1 0 5376 0 -1 1584
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5902_6
timestamp 1731220421
transform 1 0 5104 0 1 1600
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5901_6
timestamp 1731220421
transform 1 0 4968 0 1 1600
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5900_6
timestamp 1731220421
transform 1 0 5240 0 -1 1584
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5899_6
timestamp 1731220421
transform 1 0 5104 0 -1 1584
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5898_6
timestamp 1731220421
transform 1 0 4968 0 -1 1584
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5897_6
timestamp 1731220421
transform 1 0 4832 0 -1 1584
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5896_6
timestamp 1731220421
transform 1 0 4696 0 -1 1584
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5895_6
timestamp 1731220421
transform 1 0 4560 0 -1 1584
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5894_6
timestamp 1731220421
transform 1 0 4560 0 1 1600
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5893_6
timestamp 1731220421
transform 1 0 4696 0 1 1600
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5892_6
timestamp 1731220421
transform 1 0 4832 0 1 1600
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5891_6
timestamp 1731220421
transform 1 0 4920 0 -1 1840
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5890_6
timestamp 1731220421
transform 1 0 4784 0 -1 1840
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5889_6
timestamp 1731220421
transform 1 0 4648 0 -1 1840
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5888_6
timestamp 1731220421
transform 1 0 4512 0 -1 1840
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5887_6
timestamp 1731220421
transform 1 0 4376 0 -1 1840
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5886_6
timestamp 1731220421
transform 1 0 5200 0 1 1840
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5885_6
timestamp 1731220421
transform 1 0 4872 0 1 1840
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5884_6
timestamp 1731220421
transform 1 0 4560 0 1 1840
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5883_6
timestamp 1731220421
transform 1 0 4280 0 1 1840
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5882_6
timestamp 1731220421
transform 1 0 4040 0 1 1840
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5881_6
timestamp 1731220421
transform 1 0 4536 0 -1 2064
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5880_6
timestamp 1731220421
transform 1 0 4688 0 -1 2064
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5879_6
timestamp 1731220421
transform 1 0 4864 0 -1 2064
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5878_6
timestamp 1731220421
transform 1 0 5056 0 -1 2064
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5877_6
timestamp 1731220421
transform 1 0 5248 0 -1 2064
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5876_6
timestamp 1731220421
transform 1 0 5312 0 1 2084
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5875_6
timestamp 1731220421
transform 1 0 5096 0 1 2084
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5874_6
timestamp 1731220421
transform 1 0 4888 0 1 2084
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5873_6
timestamp 1731220421
transform 1 0 4696 0 1 2084
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5872_6
timestamp 1731220421
transform 1 0 4536 0 1 2084
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5871_6
timestamp 1731220421
transform 1 0 4464 0 -1 2312
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5870_6
timestamp 1731220421
transform 1 0 4152 0 -1 2312
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5869_6
timestamp 1731220421
transform 1 0 4760 0 -1 2312
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5868_6
timestamp 1731220421
transform 1 0 5056 0 -1 2312
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5867_6
timestamp 1731220421
transform 1 0 5352 0 -1 2312
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5866_6
timestamp 1731220421
transform 1 0 5240 0 1 2324
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5865_6
timestamp 1731220421
transform 1 0 5104 0 1 2324
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5864_6
timestamp 1731220421
transform 1 0 4968 0 1 2324
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5863_6
timestamp 1731220421
transform 1 0 4832 0 1 2324
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5862_6
timestamp 1731220421
transform 1 0 4696 0 1 2324
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5861_6
timestamp 1731220421
transform 1 0 5008 0 -1 2564
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5860_6
timestamp 1731220421
transform 1 0 4872 0 -1 2564
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5859_6
timestamp 1731220421
transform 1 0 4736 0 -1 2564
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5858_6
timestamp 1731220421
transform 1 0 4600 0 -1 2564
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5857_6
timestamp 1731220421
transform 1 0 4464 0 -1 2564
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5856_6
timestamp 1731220421
transform 1 0 5008 0 1 2568
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5855_6
timestamp 1731220421
transform 1 0 4752 0 1 2568
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5854_6
timestamp 1731220421
transform 1 0 4512 0 1 2568
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5853_6
timestamp 1731220421
transform 1 0 4296 0 1 2568
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5852_6
timestamp 1731220421
transform 1 0 4096 0 1 2568
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5851_6
timestamp 1731220421
transform 1 0 4432 0 -1 2804
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5850_6
timestamp 1731220421
transform 1 0 4296 0 -1 2804
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5849_6
timestamp 1731220421
transform 1 0 4160 0 -1 2804
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5848_6
timestamp 1731220421
transform 1 0 4024 0 -1 2804
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5847_6
timestamp 1731220421
transform 1 0 3888 0 -1 2804
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5846_6
timestamp 1731220421
transform 1 0 3992 0 1 2808
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5845_6
timestamp 1731220421
transform 1 0 4208 0 1 2808
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5844_6
timestamp 1731220421
transform 1 0 4968 0 1 2808
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5843_6
timestamp 1731220421
transform 1 0 4696 0 1 2808
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5842_6
timestamp 1731220421
transform 1 0 4440 0 1 2808
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5841_6
timestamp 1731220421
transform 1 0 4424 0 -1 3056
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5840_6
timestamp 1731220421
transform 1 0 4224 0 -1 3056
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5839_6
timestamp 1731220421
transform 1 0 5136 0 -1 3056
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5838_6
timestamp 1731220421
transform 1 0 4880 0 -1 3056
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5837_6
timestamp 1731220421
transform 1 0 4640 0 -1 3056
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5836_6
timestamp 1731220421
transform 1 0 4464 0 1 3056
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5835_6
timestamp 1731220421
transform 1 0 4648 0 1 3056
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5834_6
timestamp 1731220421
transform 1 0 5304 0 1 3056
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5833_6
timestamp 1731220421
transform 1 0 5072 0 1 3056
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5832_6
timestamp 1731220421
transform 1 0 4856 0 1 3056
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5831_6
timestamp 1731220421
transform 1 0 4576 0 -1 3296
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5830_6
timestamp 1731220421
transform 1 0 4344 0 -1 3296
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5829_6
timestamp 1731220421
transform 1 0 4984 0 -1 3296
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5828_6
timestamp 1731220421
transform 1 0 4784 0 -1 3296
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5827_6
timestamp 1731220421
transform 1 0 4584 0 1 3296
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5826_6
timestamp 1731220421
transform 1 0 4808 0 1 3296
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5825_6
timestamp 1731220421
transform 1 0 5024 0 1 3296
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5824_6
timestamp 1731220421
transform 1 0 5232 0 1 3296
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5823_6
timestamp 1731220421
transform 1 0 5448 0 1 3296
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5822_6
timestamp 1731220421
transform 1 0 5352 0 -1 3296
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5821_6
timestamp 1731220421
transform 1 0 5168 0 -1 3296
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5820_6
timestamp 1731220421
transform 1 0 5392 0 -1 3056
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5819_6
timestamp 1731220421
transform 1 0 5248 0 1 2808
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5818_6
timestamp 1731220421
transform 1 0 5272 0 1 2568
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5817_6
timestamp 1731220421
transform 1 0 5376 0 1 2324
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5816_6
timestamp 1731220421
transform 1 0 5448 0 -1 2064
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5815_6
timestamp 1731220421
transform 1 0 5376 0 1 1600
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5814_6
timestamp 1731220421
transform 1 0 5240 0 1 1600
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5813_6
timestamp 1731220421
transform 1 0 5512 0 1 1600
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5812_6
timestamp 1731220421
transform 1 0 5512 0 1 1840
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5811_6
timestamp 1731220421
transform 1 0 5512 0 1 2084
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5810_6
timestamp 1731220421
transform 1 0 5512 0 1 2324
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5809_6
timestamp 1731220421
transform 1 0 5512 0 1 2568
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5808_6
timestamp 1731220421
transform 1 0 5512 0 1 2808
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5807_6
timestamp 1731220421
transform 1 0 5512 0 1 3056
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5806_6
timestamp 1731220421
transform 1 0 5512 0 -1 3296
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5805_6
timestamp 1731220421
transform 1 0 5512 0 -1 3528
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5804_6
timestamp 1731220421
transform 1 0 5376 0 -1 3528
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5803_6
timestamp 1731220421
transform 1 0 5512 0 1 3576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5802_6
timestamp 1731220421
transform 1 0 5376 0 1 3576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5801_6
timestamp 1731220421
transform 1 0 5240 0 1 3576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5800_6
timestamp 1731220421
transform 1 0 5104 0 1 3576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5799_6
timestamp 1731220421
transform 1 0 4968 0 1 3576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5798_6
timestamp 1731220421
transform 1 0 4832 0 1 3576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5797_6
timestamp 1731220421
transform 1 0 4696 0 1 3576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5796_6
timestamp 1731220421
transform 1 0 4560 0 1 3576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5795_6
timestamp 1731220421
transform 1 0 4424 0 1 3576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5794_6
timestamp 1731220421
transform 1 0 4288 0 1 3576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5793_6
timestamp 1731220421
transform 1 0 4152 0 1 3576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5792_6
timestamp 1731220421
transform 1 0 4016 0 1 3576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5791_6
timestamp 1731220421
transform 1 0 5016 0 -1 3820
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5790_6
timestamp 1731220421
transform 1 0 4880 0 -1 3820
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5789_6
timestamp 1731220421
transform 1 0 4744 0 -1 3820
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5788_6
timestamp 1731220421
transform 1 0 4608 0 -1 3820
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5787_6
timestamp 1731220421
transform 1 0 4472 0 -1 3820
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5786_6
timestamp 1731220421
transform 1 0 4776 0 1 3848
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5785_6
timestamp 1731220421
transform 1 0 4616 0 1 3848
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5784_6
timestamp 1731220421
transform 1 0 4456 0 1 3848
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5783_6
timestamp 1731220421
transform 1 0 4296 0 1 3848
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5782_6
timestamp 1731220421
transform 1 0 4144 0 1 3848
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5781_6
timestamp 1731220421
transform 1 0 4808 0 -1 4072
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5780_6
timestamp 1731220421
transform 1 0 4672 0 -1 4072
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5779_6
timestamp 1731220421
transform 1 0 4536 0 -1 4072
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5778_6
timestamp 1731220421
transform 1 0 4400 0 -1 4072
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5777_6
timestamp 1731220421
transform 1 0 4264 0 -1 4072
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5776_6
timestamp 1731220421
transform 1 0 4104 0 1 4096
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5775_6
timestamp 1731220421
transform 1 0 3968 0 1 4096
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5774_6
timestamp 1731220421
transform 1 0 4512 0 1 4096
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5773_6
timestamp 1731220421
transform 1 0 4376 0 1 4096
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5772_6
timestamp 1731220421
transform 1 0 4240 0 1 4096
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5771_6
timestamp 1731220421
transform 1 0 4104 0 -1 4332
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5770_6
timestamp 1731220421
transform 1 0 4240 0 -1 4332
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5769_6
timestamp 1731220421
transform 1 0 4648 0 -1 4332
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5768_6
timestamp 1731220421
transform 1 0 4512 0 -1 4332
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5767_6
timestamp 1731220421
transform 1 0 4376 0 -1 4332
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5766_6
timestamp 1731220421
transform 1 0 4344 0 1 4348
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5765_6
timestamp 1731220421
transform 1 0 4480 0 1 4348
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5764_6
timestamp 1731220421
transform 1 0 4616 0 1 4348
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5763_6
timestamp 1731220421
transform 1 0 4752 0 1 4348
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5762_6
timestamp 1731220421
transform 1 0 4888 0 1 4348
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5761_6
timestamp 1731220421
transform 1 0 5048 0 -1 4576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5760_6
timestamp 1731220421
transform 1 0 4912 0 -1 4576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5759_6
timestamp 1731220421
transform 1 0 4776 0 -1 4576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5758_6
timestamp 1731220421
transform 1 0 4640 0 -1 4576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5757_6
timestamp 1731220421
transform 1 0 4400 0 1 4576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5756_6
timestamp 1731220421
transform 1 0 4264 0 1 4576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5755_6
timestamp 1731220421
transform 1 0 4128 0 1 4576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5754_6
timestamp 1731220421
transform 1 0 4536 0 1 4576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5753_6
timestamp 1731220421
transform 1 0 4672 0 1 4576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5752_6
timestamp 1731220421
transform 1 0 4816 0 1 4576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5751_6
timestamp 1731220421
transform 1 0 4960 0 1 4576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5750_6
timestamp 1731220421
transform 1 0 5104 0 1 4576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5749_6
timestamp 1731220421
transform 1 0 5240 0 1 4576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5748_6
timestamp 1731220421
transform 1 0 5512 0 1 4576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5747_6
timestamp 1731220421
transform 1 0 5376 0 1 4576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5746_6
timestamp 1731220421
transform 1 0 5272 0 -1 4800
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5745_6
timestamp 1731220421
transform 1 0 5008 0 -1 4800
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5744_6
timestamp 1731220421
transform 1 0 5512 0 -1 4800
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5743_6
timestamp 1731220421
transform 1 0 5512 0 1 4876
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5742_6
timestamp 1731220421
transform 1 0 5376 0 1 4876
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5741_6
timestamp 1731220421
transform 1 0 5280 0 -1 5100
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5740_6
timestamp 1731220421
transform 1 0 5032 0 -1 5100
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5739_6
timestamp 1731220421
transform 1 0 5512 0 -1 5100
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5738_6
timestamp 1731220421
transform 1 0 5512 0 1 5108
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5737_6
timestamp 1731220421
transform 1 0 5376 0 1 5108
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5736_6
timestamp 1731220421
transform 1 0 5216 0 1 5108
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5735_6
timestamp 1731220421
transform 1 0 5064 0 1 5108
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5734_6
timestamp 1731220421
transform 1 0 4912 0 1 5108
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5733_6
timestamp 1731220421
transform 1 0 4752 0 1 5108
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5732_6
timestamp 1731220421
transform 1 0 4592 0 1 5108
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5731_6
timestamp 1731220421
transform 1 0 4768 0 -1 5348
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5730_6
timestamp 1731220421
transform 1 0 4952 0 -1 5348
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5729_6
timestamp 1731220421
transform 1 0 5144 0 -1 5348
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5728_6
timestamp 1731220421
transform 1 0 5072 0 1 5356
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5727_6
timestamp 1731220421
transform 1 0 4904 0 1 5356
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5726_6
timestamp 1731220421
transform 1 0 4744 0 1 5356
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5725_6
timestamp 1731220421
transform 1 0 5080 0 -1 5580
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5724_6
timestamp 1731220421
transform 1 0 4944 0 -1 5580
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5723_6
timestamp 1731220421
transform 1 0 4808 0 -1 5580
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5722_6
timestamp 1731220421
transform 1 0 4672 0 -1 5580
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5721_6
timestamp 1731220421
transform 1 0 4872 0 1 5580
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5720_6
timestamp 1731220421
transform 1 0 4736 0 1 5580
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5719_6
timestamp 1731220421
transform 1 0 4600 0 1 5580
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5718_6
timestamp 1731220421
transform 1 0 4464 0 1 5580
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5717_6
timestamp 1731220421
transform 1 0 4400 0 -1 5580
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5716_6
timestamp 1731220421
transform 1 0 4536 0 -1 5580
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5715_6
timestamp 1731220421
transform 1 0 4584 0 1 5356
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5714_6
timestamp 1731220421
transform 1 0 4424 0 1 5356
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5713_6
timestamp 1731220421
transform 1 0 4400 0 -1 5348
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5712_6
timestamp 1731220421
transform 1 0 4584 0 -1 5348
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5711_6
timestamp 1731220421
transform 1 0 4432 0 1 5108
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5710_6
timestamp 1731220421
transform 1 0 4296 0 -1 5100
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5709_6
timestamp 1731220421
transform 1 0 4536 0 -1 5100
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5708_6
timestamp 1731220421
transform 1 0 4784 0 -1 5100
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5707_6
timestamp 1731220421
transform 1 0 5224 0 1 4876
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5706_6
timestamp 1731220421
transform 1 0 5080 0 1 4876
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5705_6
timestamp 1731220421
transform 1 0 4944 0 1 4876
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5704_6
timestamp 1731220421
transform 1 0 4808 0 1 4876
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5703_6
timestamp 1731220421
transform 1 0 4672 0 1 4876
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5702_6
timestamp 1731220421
transform 1 0 4536 0 1 4876
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5701_6
timestamp 1731220421
transform 1 0 4400 0 1 4876
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5700_6
timestamp 1731220421
transform 1 0 4264 0 1 4876
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5699_6
timestamp 1731220421
transform 1 0 4128 0 1 4876
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5698_6
timestamp 1731220421
transform 1 0 4056 0 -1 5100
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5697_6
timestamp 1731220421
transform 1 0 3856 0 -1 5100
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5696_6
timestamp 1731220421
transform 1 0 3992 0 1 4876
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5695_6
timestamp 1731220421
transform 1 0 3856 0 1 4876
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5694_6
timestamp 1731220421
transform 1 0 3648 0 1 4872
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5693_6
timestamp 1731220421
transform 1 0 3648 0 -1 4864
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5692_6
timestamp 1731220421
transform 1 0 3856 0 -1 4800
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5691_6
timestamp 1731220421
transform 1 0 4040 0 -1 4800
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5690_6
timestamp 1731220421
transform 1 0 4752 0 -1 4800
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5689_6
timestamp 1731220421
transform 1 0 4504 0 -1 4800
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5688_6
timestamp 1731220421
transform 1 0 4264 0 -1 4800
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5687_6
timestamp 1731220421
transform 1 0 3992 0 1 4576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5686_6
timestamp 1731220421
transform 1 0 3856 0 1 4576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5685_6
timestamp 1731220421
transform 1 0 3648 0 -1 4624
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5684_6
timestamp 1731220421
transform 1 0 3440 0 -1 4624
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5683_6
timestamp 1731220421
transform 1 0 3216 0 -1 4624
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5682_6
timestamp 1731220421
transform 1 0 2984 0 -1 4624
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5681_6
timestamp 1731220421
transform 1 0 3608 0 1 4388
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5680_6
timestamp 1731220421
transform 1 0 3392 0 1 4388
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5679_6
timestamp 1731220421
transform 1 0 3184 0 1 4388
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5678_6
timestamp 1731220421
transform 1 0 2968 0 1 4388
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5677_6
timestamp 1731220421
transform 1 0 2744 0 1 4388
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5676_6
timestamp 1731220421
transform 1 0 3288 0 -1 4376
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5675_6
timestamp 1731220421
transform 1 0 3104 0 -1 4376
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5674_6
timestamp 1731220421
transform 1 0 2920 0 -1 4376
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5673_6
timestamp 1731220421
transform 1 0 2744 0 -1 4376
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5672_6
timestamp 1731220421
transform 1 0 2560 0 -1 4376
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5671_6
timestamp 1731220421
transform 1 0 2504 0 1 4148
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5670_6
timestamp 1731220421
transform 1 0 2240 0 1 4148
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5669_6
timestamp 1731220421
transform 1 0 2760 0 1 4148
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5668_6
timestamp 1731220421
transform 1 0 3016 0 1 4148
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5667_6
timestamp 1731220421
transform 1 0 3280 0 1 4148
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5666_6
timestamp 1731220421
transform 1 0 3240 0 -1 4136
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5665_6
timestamp 1731220421
transform 1 0 3104 0 -1 4136
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5664_6
timestamp 1731220421
transform 1 0 3376 0 -1 4136
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5663_6
timestamp 1731220421
transform 1 0 3512 0 -1 4136
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5662_6
timestamp 1731220421
transform 1 0 3648 0 -1 4136
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5661_6
timestamp 1731220421
transform 1 0 3856 0 -1 4072
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5660_6
timestamp 1731220421
transform 1 0 3992 0 -1 4072
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5659_6
timestamp 1731220421
transform 1 0 4128 0 -1 4072
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5658_6
timestamp 1731220421
transform 1 0 3992 0 1 3848
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5657_6
timestamp 1731220421
transform 1 0 3856 0 1 3848
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5656_6
timestamp 1731220421
transform 1 0 3648 0 1 3820
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5655_6
timestamp 1731220421
transform 1 0 3248 0 1 3820
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5654_6
timestamp 1731220421
transform 1 0 2824 0 1 3820
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5653_6
timestamp 1731220421
transform 1 0 2400 0 1 3820
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5652_6
timestamp 1731220421
transform 1 0 3576 0 -1 3820
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5651_6
timestamp 1731220421
transform 1 0 3392 0 -1 3820
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5650_6
timestamp 1731220421
transform 1 0 3216 0 -1 3820
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5649_6
timestamp 1731220421
transform 1 0 3040 0 -1 3820
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5648_6
timestamp 1731220421
transform 1 0 2864 0 -1 3820
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5647_6
timestamp 1731220421
transform 1 0 3296 0 1 3588
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5646_6
timestamp 1731220421
transform 1 0 3152 0 1 3588
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5645_6
timestamp 1731220421
transform 1 0 3008 0 1 3588
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5644_6
timestamp 1731220421
transform 1 0 2864 0 1 3588
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5643_6
timestamp 1731220421
transform 1 0 2720 0 1 3588
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5642_6
timestamp 1731220421
transform 1 0 2888 0 -1 3580
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5641_6
timestamp 1731220421
transform 1 0 3024 0 -1 3580
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5640_6
timestamp 1731220421
transform 1 0 3160 0 -1 3580
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5639_6
timestamp 1731220421
transform 1 0 3432 0 -1 3580
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5638_6
timestamp 1731220421
transform 1 0 3296 0 -1 3580
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5637_6
timestamp 1731220421
transform 1 0 3288 0 1 3352
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5636_6
timestamp 1731220421
transform 1 0 3096 0 1 3352
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5635_6
timestamp 1731220421
transform 1 0 3480 0 1 3352
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5634_6
timestamp 1731220421
transform 1 0 3648 0 1 3352
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5633_6
timestamp 1731220421
transform 1 0 3856 0 1 3296
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5632_6
timestamp 1731220421
transform 1 0 4096 0 1 3296
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5631_6
timestamp 1731220421
transform 1 0 4344 0 1 3296
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5630_6
timestamp 1731220421
transform 1 0 4096 0 -1 3296
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5629_6
timestamp 1731220421
transform 1 0 3856 0 -1 3296
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5628_6
timestamp 1731220421
transform 1 0 3648 0 -1 3328
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5627_6
timestamp 1731220421
transform 1 0 3648 0 1 3104
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5626_6
timestamp 1731220421
transform 1 0 3440 0 1 3104
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5625_6
timestamp 1731220421
transform 1 0 3208 0 1 3104
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5624_6
timestamp 1731220421
transform 1 0 3368 0 -1 3104
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5623_6
timestamp 1731220421
transform 1 0 3536 0 -1 3104
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5622_6
timestamp 1731220421
transform 1 0 3480 0 1 2880
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5621_6
timestamp 1731220421
transform 1 0 3344 0 1 2880
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5620_6
timestamp 1731220421
transform 1 0 3208 0 1 2880
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5619_6
timestamp 1731220421
transform 1 0 3072 0 1 2880
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5618_6
timestamp 1731220421
transform 1 0 3208 0 -1 3104
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5617_6
timestamp 1731220421
transform 1 0 3048 0 -1 3104
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5616_6
timestamp 1731220421
transform 1 0 2896 0 -1 3104
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5615_6
timestamp 1731220421
transform 1 0 2768 0 1 3104
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5614_6
timestamp 1731220421
transform 1 0 2552 0 1 3104
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5613_6
timestamp 1731220421
transform 1 0 2656 0 -1 3328
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5612_6
timestamp 1731220421
transform 1 0 2368 0 -1 3328
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5611_6
timestamp 1731220421
transform 1 0 2120 0 -1 3328
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5610_6
timestamp 1731220421
transform 1 0 2344 0 1 3104
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5609_6
timestamp 1731220421
transform 1 0 2144 0 1 3104
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5608_6
timestamp 1731220421
transform 1 0 1992 0 1 3104
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5607_6
timestamp 1731220421
transform 1 0 1784 0 1 3024
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5606_6
timestamp 1731220421
transform 1 0 1576 0 1 3024
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5605_6
timestamp 1731220421
transform 1 0 1344 0 1 3024
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5604_6
timestamp 1731220421
transform 1 0 1784 0 -1 3024
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5603_6
timestamp 1731220421
transform 1 0 1640 0 -1 3024
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5602_6
timestamp 1731220421
transform 1 0 1480 0 -1 3024
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5601_6
timestamp 1731220421
transform 1 0 1320 0 -1 3024
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5600_6
timestamp 1731220421
transform 1 0 1152 0 -1 3024
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5599_6
timestamp 1731220421
transform 1 0 1312 0 1 2796
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5598_6
timestamp 1731220421
transform 1 0 1480 0 1 2796
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5597_6
timestamp 1731220421
transform 1 0 1640 0 1 2796
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5596_6
timestamp 1731220421
transform 1 0 1784 0 1 2796
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5595_6
timestamp 1731220421
transform 1 0 1992 0 -1 2828
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5594_6
timestamp 1731220421
transform 1 0 2136 0 -1 2828
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5593_6
timestamp 1731220421
transform 1 0 2304 0 -1 2828
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5592_6
timestamp 1731220421
transform 1 0 2464 0 -1 2828
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5591_6
timestamp 1731220421
transform 1 0 2376 0 1 2604
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5590_6
timestamp 1731220421
transform 1 0 2512 0 1 2604
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5589_6
timestamp 1731220421
transform 1 0 2480 0 -1 2600
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5588_6
timestamp 1731220421
transform 1 0 2616 0 -1 2600
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5587_6
timestamp 1731220421
transform 1 0 2752 0 -1 2600
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5586_6
timestamp 1731220421
transform 1 0 2712 0 1 2360
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5585_6
timestamp 1731220421
transform 1 0 2512 0 1 2360
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5584_6
timestamp 1731220421
transform 1 0 2304 0 1 2360
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5583_6
timestamp 1731220421
transform 1 0 2192 0 -1 2352
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5582_6
timestamp 1731220421
transform 1 0 2472 0 -1 2352
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5581_6
timestamp 1731220421
transform 1 0 3328 0 1 2128
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5580_6
timestamp 1731220421
transform 1 0 2984 0 1 2128
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5579_6
timestamp 1731220421
transform 1 0 2664 0 1 2128
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5578_6
timestamp 1731220421
transform 1 0 2384 0 1 2128
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5577_6
timestamp 1731220421
transform 1 0 2152 0 1 2128
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5576_6
timestamp 1731220421
transform 1 0 1992 0 1 2128
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5575_6
timestamp 1731220421
transform 1 0 1784 0 -1 2304
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5574_6
timestamp 1731220421
transform 1 0 1784 0 1 2308
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5573_6
timestamp 1731220421
transform 1 0 1544 0 1 2308
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5572_6
timestamp 1731220421
transform 1 0 1288 0 1 2308
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5571_6
timestamp 1731220421
transform 1 0 1424 0 -1 2544
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5570_6
timestamp 1731220421
transform 1 0 1584 0 -1 2544
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5569_6
timestamp 1731220421
transform 1 0 1752 0 -1 2544
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5568_6
timestamp 1731220421
transform 1 0 1720 0 1 2560
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5567_6
timestamp 1731220421
transform 1 0 1584 0 1 2560
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5566_6
timestamp 1731220421
transform 1 0 1448 0 1 2560
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5565_6
timestamp 1731220421
transform 1 0 1448 0 -1 2784
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5564_6
timestamp 1731220421
transform 1 0 1280 0 -1 2784
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5563_6
timestamp 1731220421
transform 1 0 1112 0 -1 2784
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5562_6
timestamp 1731220421
transform 1 0 1144 0 1 2796
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5561_6
timestamp 1731220421
transform 1 0 968 0 1 2796
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5560_6
timestamp 1731220421
transform 1 0 784 0 1 2796
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5559_6
timestamp 1731220421
transform 1 0 976 0 -1 3024
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5558_6
timestamp 1731220421
transform 1 0 792 0 -1 3024
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5557_6
timestamp 1731220421
transform 1 0 592 0 -1 3024
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5556_6
timestamp 1731220421
transform 1 0 624 0 1 3024
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5555_6
timestamp 1731220421
transform 1 0 872 0 1 3024
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5554_6
timestamp 1731220421
transform 1 0 1112 0 1 3024
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5553_6
timestamp 1731220421
transform 1 0 928 0 -1 3264
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5552_6
timestamp 1731220421
transform 1 0 720 0 -1 3264
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5551_6
timestamp 1731220421
transform 1 0 592 0 1 3272
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5550_6
timestamp 1731220421
transform 1 0 864 0 1 3272
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5549_6
timestamp 1731220421
transform 1 0 728 0 1 3272
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5548_6
timestamp 1731220421
transform 1 0 672 0 -1 3504
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5547_6
timestamp 1731220421
transform 1 0 536 0 -1 3504
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5546_6
timestamp 1731220421
transform 1 0 400 0 -1 3504
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5545_6
timestamp 1731220421
transform 1 0 320 0 1 3272
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5544_6
timestamp 1731220421
transform 1 0 456 0 1 3272
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5543_6
timestamp 1731220421
transform 1 0 512 0 -1 3264
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5542_6
timestamp 1731220421
transform 1 0 304 0 -1 3264
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5541_6
timestamp 1731220421
transform 1 0 128 0 -1 3264
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5540_6
timestamp 1731220421
transform 1 0 128 0 1 3024
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5539_6
timestamp 1731220421
transform 1 0 368 0 1 3024
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5538_6
timestamp 1731220421
transform 1 0 144 0 -1 3024
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5537_6
timestamp 1731220421
transform 1 0 376 0 -1 3024
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5536_6
timestamp 1731220421
transform 1 0 392 0 1 2796
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5535_6
timestamp 1731220421
transform 1 0 592 0 1 2796
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5534_6
timestamp 1731220421
transform 1 0 624 0 -1 2784
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5533_6
timestamp 1731220421
transform 1 0 784 0 -1 2784
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5532_6
timestamp 1731220421
transform 1 0 944 0 -1 2784
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5531_6
timestamp 1731220421
transform 1 0 904 0 1 2560
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5530_6
timestamp 1731220421
transform 1 0 768 0 1 2560
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5529_6
timestamp 1731220421
transform 1 0 1040 0 1 2560
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5528_6
timestamp 1731220421
transform 1 0 1176 0 1 2560
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5527_6
timestamp 1731220421
transform 1 0 1312 0 1 2560
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5526_6
timestamp 1731220421
transform 1 0 1264 0 -1 2544
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5525_6
timestamp 1731220421
transform 1 0 1104 0 -1 2544
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5524_6
timestamp 1731220421
transform 1 0 952 0 -1 2544
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5523_6
timestamp 1731220421
transform 1 0 800 0 -1 2544
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5522_6
timestamp 1731220421
transform 1 0 656 0 -1 2544
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5521_6
timestamp 1731220421
transform 1 0 520 0 -1 2544
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5520_6
timestamp 1731220421
transform 1 0 1040 0 1 2308
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5519_6
timestamp 1731220421
transform 1 0 800 0 1 2308
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5518_6
timestamp 1731220421
transform 1 0 560 0 1 2308
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5517_6
timestamp 1731220421
transform 1 0 336 0 1 2308
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5516_6
timestamp 1731220421
transform 1 0 128 0 1 2308
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5515_6
timestamp 1731220421
transform 1 0 800 0 -1 2304
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5514_6
timestamp 1731220421
transform 1 0 520 0 -1 2304
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5513_6
timestamp 1731220421
transform 1 0 288 0 -1 2304
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5512_6
timestamp 1731220421
transform 1 0 128 0 -1 2304
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5511_6
timestamp 1731220421
transform 1 0 1120 0 -1 2304
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5510_6
timestamp 1731220421
transform 1 0 1464 0 -1 2304
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5509_6
timestamp 1731220421
transform 1 0 1144 0 1 2056
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5508_6
timestamp 1731220421
transform 1 0 480 0 1 2056
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5507_6
timestamp 1731220421
transform 1 0 288 0 1 2056
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5506_6
timestamp 1731220421
transform 1 0 688 0 1 2056
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5505_6
timestamp 1731220421
transform 1 0 912 0 1 2056
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5504_6
timestamp 1731220421
transform 1 0 936 0 -1 2052
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5503_6
timestamp 1731220421
transform 1 0 792 0 -1 2052
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5502_6
timestamp 1731220421
transform 1 0 648 0 -1 2052
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5501_6
timestamp 1731220421
transform 1 0 504 0 -1 2052
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5500_6
timestamp 1731220421
transform 1 0 368 0 -1 2052
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5499_6
timestamp 1731220421
transform 1 0 232 0 -1 2052
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5498_6
timestamp 1731220421
transform 1 0 624 0 1 1816
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5497_6
timestamp 1731220421
transform 1 0 432 0 1 1816
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5496_6
timestamp 1731220421
transform 1 0 232 0 1 1816
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5495_6
timestamp 1731220421
transform 1 0 192 0 -1 1804
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5494_6
timestamp 1731220421
transform 1 0 432 0 -1 1804
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5493_6
timestamp 1731220421
transform 1 0 360 0 1 1568
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5492_6
timestamp 1731220421
transform 1 0 128 0 1 1568
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5491_6
timestamp 1731220421
transform 1 0 128 0 -1 1556
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5490_6
timestamp 1731220421
transform 1 0 296 0 -1 1556
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5489_6
timestamp 1731220421
transform 1 0 392 0 1 1320
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5488_6
timestamp 1731220421
transform 1 0 128 0 1 1320
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5487_6
timestamp 1731220421
transform 1 0 128 0 -1 1320
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5486_6
timestamp 1731220421
transform 1 0 424 0 -1 1320
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5485_6
timestamp 1731220421
transform 1 0 560 0 1 1072
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5484_6
timestamp 1731220421
transform 1 0 328 0 1 1072
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5483_6
timestamp 1731220421
transform 1 0 128 0 1 1072
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5482_6
timestamp 1731220421
transform 1 0 232 0 -1 1072
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5481_6
timestamp 1731220421
transform 1 0 408 0 -1 1072
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5480_6
timestamp 1731220421
transform 1 0 376 0 1 844
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5479_6
timestamp 1731220421
transform 1 0 224 0 1 844
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5478_6
timestamp 1731220421
transform 1 0 624 0 -1 828
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5477_6
timestamp 1731220421
transform 1 0 344 0 -1 828
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5476_6
timestamp 1731220421
transform 1 0 304 0 1 604
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5475_6
timestamp 1731220421
transform 1 0 128 0 1 604
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5474_6
timestamp 1731220421
transform 1 0 496 0 1 604
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5473_6
timestamp 1731220421
transform 1 0 344 0 -1 604
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5472_6
timestamp 1731220421
transform 1 0 128 0 -1 604
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5471_6
timestamp 1731220421
transform 1 0 128 0 1 380
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5470_6
timestamp 1731220421
transform 1 0 424 0 1 380
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5469_6
timestamp 1731220421
transform 1 0 520 0 -1 364
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5468_6
timestamp 1731220421
transform 1 0 360 0 -1 364
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5467_6
timestamp 1731220421
transform 1 0 208 0 -1 364
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5466_6
timestamp 1731220421
transform 1 0 144 0 1 108
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5465_6
timestamp 1731220421
transform 1 0 280 0 1 108
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5464_6
timestamp 1731220421
transform 1 0 416 0 1 108
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5463_6
timestamp 1731220421
transform 1 0 552 0 1 108
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5462_6
timestamp 1731220421
transform 1 0 688 0 1 108
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5461_6
timestamp 1731220421
transform 1 0 1096 0 1 108
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5460_6
timestamp 1731220421
transform 1 0 960 0 1 108
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5459_6
timestamp 1731220421
transform 1 0 824 0 1 108
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5458_6
timestamp 1731220421
transform 1 0 680 0 -1 364
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5457_6
timestamp 1731220421
transform 1 0 840 0 -1 364
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5456_6
timestamp 1731220421
transform 1 0 1000 0 -1 364
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5455_6
timestamp 1731220421
transform 1 0 1456 0 1 380
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5454_6
timestamp 1731220421
transform 1 0 1104 0 1 380
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5453_6
timestamp 1731220421
transform 1 0 760 0 1 380
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5452_6
timestamp 1731220421
transform 1 0 568 0 -1 604
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5451_6
timestamp 1731220421
transform 1 0 776 0 -1 604
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5450_6
timestamp 1731220421
transform 1 0 968 0 -1 604
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5449_6
timestamp 1731220421
transform 1 0 856 0 1 604
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5448_6
timestamp 1731220421
transform 1 0 680 0 1 604
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5447_6
timestamp 1731220421
transform 1 0 1024 0 1 604
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5446_6
timestamp 1731220421
transform 1 0 912 0 -1 828
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5445_6
timestamp 1731220421
transform 1 0 1208 0 -1 828
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5444_6
timestamp 1731220421
transform 1 0 1072 0 1 844
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5443_6
timestamp 1731220421
transform 1 0 888 0 1 844
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5442_6
timestamp 1731220421
transform 1 0 712 0 1 844
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5441_6
timestamp 1731220421
transform 1 0 536 0 1 844
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5440_6
timestamp 1731220421
transform 1 0 584 0 -1 1072
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5439_6
timestamp 1731220421
transform 1 0 752 0 -1 1072
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5438_6
timestamp 1731220421
transform 1 0 920 0 -1 1072
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5437_6
timestamp 1731220421
transform 1 0 800 0 1 1072
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5436_6
timestamp 1731220421
transform 1 0 1040 0 1 1072
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5435_6
timestamp 1731220421
transform 1 0 1280 0 1 1072
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5434_6
timestamp 1731220421
transform 1 0 1064 0 -1 1320
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5433_6
timestamp 1731220421
transform 1 0 744 0 -1 1320
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5432_6
timestamp 1731220421
transform 1 0 1392 0 -1 1320
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5431_6
timestamp 1731220421
transform 1 0 1256 0 1 1320
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5430_6
timestamp 1731220421
transform 1 0 968 0 1 1320
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5429_6
timestamp 1731220421
transform 1 0 680 0 1 1320
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5428_6
timestamp 1731220421
transform 1 0 1048 0 -1 1556
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5427_6
timestamp 1731220421
transform 1 0 856 0 -1 1556
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5426_6
timestamp 1731220421
transform 1 0 664 0 -1 1556
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5425_6
timestamp 1731220421
transform 1 0 480 0 -1 1556
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5424_6
timestamp 1731220421
transform 1 0 616 0 1 1568
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5423_6
timestamp 1731220421
transform 1 0 872 0 1 1568
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5422_6
timestamp 1731220421
transform 1 0 1136 0 1 1568
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5421_6
timestamp 1731220421
transform 1 0 1128 0 -1 1804
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5420_6
timestamp 1731220421
transform 1 0 896 0 -1 1804
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5419_6
timestamp 1731220421
transform 1 0 664 0 -1 1804
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5418_6
timestamp 1731220421
transform 1 0 1360 0 -1 1804
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5417_6
timestamp 1731220421
transform 1 0 1152 0 1 1816
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5416_6
timestamp 1731220421
transform 1 0 984 0 1 1816
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5415_6
timestamp 1731220421
transform 1 0 808 0 1 1816
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5414_6
timestamp 1731220421
transform 1 0 1080 0 -1 2052
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5413_6
timestamp 1731220421
transform 1 0 1224 0 -1 2052
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5412_6
timestamp 1731220421
transform 1 0 1368 0 -1 2052
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5411_6
timestamp 1731220421
transform 1 0 1384 0 1 2056
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5410_6
timestamp 1731220421
transform 1 0 1632 0 1 2056
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5409_6
timestamp 1731220421
transform 1 0 1512 0 -1 2052
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5408_6
timestamp 1731220421
transform 1 0 1784 0 -1 2052
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5407_6
timestamp 1731220421
transform 1 0 1648 0 -1 2052
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5406_6
timestamp 1731220421
transform 1 0 1640 0 1 1816
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5405_6
timestamp 1731220421
transform 1 0 1480 0 1 1816
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5404_6
timestamp 1731220421
transform 1 0 1320 0 1 1816
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5403_6
timestamp 1731220421
transform 1 0 1784 0 1 1816
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5402_6
timestamp 1731220421
transform 1 0 1992 0 1 1692
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5401_6
timestamp 1731220421
transform 1 0 2128 0 1 1692
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5400_6
timestamp 1731220421
transform 1 0 2264 0 1 1692
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5399_6
timestamp 1731220421
transform 1 0 2416 0 1 1692
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5398_6
timestamp 1731220421
transform 1 0 2576 0 1 1692
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5397_6
timestamp 1731220421
transform 1 0 2736 0 1 1692
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5396_6
timestamp 1731220421
transform 1 0 2608 0 -1 1680
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5395_6
timestamp 1731220421
transform 1 0 2448 0 -1 1680
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5394_6
timestamp 1731220421
transform 1 0 2288 0 -1 1680
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5393_6
timestamp 1731220421
transform 1 0 2136 0 -1 1680
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5392_6
timestamp 1731220421
transform 1 0 1992 0 -1 1680
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5391_6
timestamp 1731220421
transform 1 0 1992 0 1 1444
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5390_6
timestamp 1731220421
transform 1 0 2128 0 1 1444
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5389_6
timestamp 1731220421
transform 1 0 2264 0 1 1444
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5388_6
timestamp 1731220421
transform 1 0 2136 0 -1 1432
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5387_6
timestamp 1731220421
transform 1 0 2272 0 -1 1432
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5386_6
timestamp 1731220421
transform 1 0 2408 0 -1 1432
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5385_6
timestamp 1731220421
transform 1 0 2712 0 1 1208
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5384_6
timestamp 1731220421
transform 1 0 2552 0 1 1208
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5383_6
timestamp 1731220421
transform 1 0 2400 0 1 1208
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5382_6
timestamp 1731220421
transform 1 0 2264 0 1 1208
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5381_6
timestamp 1731220421
transform 1 0 2128 0 1 1208
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5380_6
timestamp 1731220421
transform 1 0 2688 0 -1 1208
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5379_6
timestamp 1731220421
transform 1 0 2448 0 -1 1208
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5378_6
timestamp 1731220421
transform 1 0 2208 0 -1 1208
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5377_6
timestamp 1731220421
transform 1 0 1992 0 -1 1208
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5376_6
timestamp 1731220421
transform 1 0 1768 0 1 1072
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5375_6
timestamp 1731220421
transform 1 0 1520 0 1 1072
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5374_6
timestamp 1731220421
transform 1 0 1720 0 -1 1072
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5373_6
timestamp 1731220421
transform 1 0 1560 0 -1 1072
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5372_6
timestamp 1731220421
transform 1 0 1400 0 -1 1072
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5371_6
timestamp 1731220421
transform 1 0 1240 0 -1 1072
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5370_6
timestamp 1731220421
transform 1 0 1080 0 -1 1072
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5369_6
timestamp 1731220421
transform 1 0 1256 0 1 844
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5368_6
timestamp 1731220421
transform 1 0 1440 0 1 844
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5367_6
timestamp 1731220421
transform 1 0 1624 0 1 844
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5366_6
timestamp 1731220421
transform 1 0 1784 0 1 844
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5365_6
timestamp 1731220421
transform 1 0 2016 0 -1 932
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5364_6
timestamp 1731220421
transform 1 0 2320 0 -1 932
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5363_6
timestamp 1731220421
transform 1 0 2520 0 1 708
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5362_6
timestamp 1731220421
transform 1 0 2248 0 1 708
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5361_6
timestamp 1731220421
transform 1 0 1992 0 1 708
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5360_6
timestamp 1731220421
transform 1 0 1784 0 -1 828
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5359_6
timestamp 1731220421
transform 1 0 1504 0 -1 828
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5358_6
timestamp 1731220421
transform 1 0 1784 0 1 604
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5357_6
timestamp 1731220421
transform 1 0 1648 0 1 604
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5356_6
timestamp 1731220421
transform 1 0 1488 0 1 604
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5355_6
timestamp 1731220421
transform 1 0 1336 0 1 604
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5354_6
timestamp 1731220421
transform 1 0 1184 0 1 604
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5353_6
timestamp 1731220421
transform 1 0 1144 0 -1 604
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5352_6
timestamp 1731220421
transform 1 0 1312 0 -1 604
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5351_6
timestamp 1731220421
transform 1 0 1480 0 -1 604
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5350_6
timestamp 1731220421
transform 1 0 1640 0 -1 604
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5349_6
timestamp 1731220421
transform 1 0 1784 0 -1 604
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5348_6
timestamp 1731220421
transform 1 0 1784 0 1 380
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5347_6
timestamp 1731220421
transform 1 0 1992 0 1 352
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5346_6
timestamp 1731220421
transform 1 0 2152 0 1 352
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5345_6
timestamp 1731220421
transform 1 0 2728 0 1 352
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5344_6
timestamp 1731220421
transform 1 0 2536 0 1 352
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5343_6
timestamp 1731220421
transform 1 0 2344 0 1 352
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5342_6
timestamp 1731220421
transform 1 0 2016 0 -1 328
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5341_6
timestamp 1731220421
transform 1 0 1992 0 1 88
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5340_6
timestamp 1731220421
transform 1 0 2128 0 1 88
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5339_6
timestamp 1731220421
transform 1 0 2264 0 1 88
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5338_6
timestamp 1731220421
transform 1 0 2400 0 1 88
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5337_6
timestamp 1731220421
transform 1 0 2808 0 1 88
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5336_6
timestamp 1731220421
transform 1 0 2672 0 1 88
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5335_6
timestamp 1731220421
transform 1 0 2536 0 1 88
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5334_6
timestamp 1731220421
transform 1 0 2424 0 -1 328
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5333_6
timestamp 1731220421
transform 1 0 2288 0 -1 328
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5332_6
timestamp 1731220421
transform 1 0 2152 0 -1 328
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5331_6
timestamp 1731220421
transform 1 0 2560 0 -1 328
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5330_6
timestamp 1731220421
transform 1 0 2696 0 -1 328
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5329_6
timestamp 1731220421
transform 1 0 2944 0 1 88
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5328_6
timestamp 1731220421
transform 1 0 3080 0 1 88
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5327_6
timestamp 1731220421
transform 1 0 3216 0 1 88
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5326_6
timestamp 1731220421
transform 1 0 3624 0 1 88
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5325_6
timestamp 1731220421
transform 1 0 3488 0 1 88
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5324_6
timestamp 1731220421
transform 1 0 3352 0 1 88
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5323_6
timestamp 1731220421
transform 1 0 3104 0 -1 328
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5322_6
timestamp 1731220421
transform 1 0 2968 0 -1 328
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5321_6
timestamp 1731220421
transform 1 0 2832 0 -1 328
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5320_6
timestamp 1731220421
transform 1 0 3240 0 -1 328
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5319_6
timestamp 1731220421
transform 1 0 3648 0 -1 328
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5318_6
timestamp 1731220421
transform 1 0 3512 0 -1 328
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5317_6
timestamp 1731220421
transform 1 0 3376 0 -1 328
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5316_6
timestamp 1731220421
transform 1 0 3296 0 1 352
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5315_6
timestamp 1731220421
transform 1 0 3112 0 1 352
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5314_6
timestamp 1731220421
transform 1 0 2920 0 1 352
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5313_6
timestamp 1731220421
transform 1 0 3480 0 1 352
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5312_6
timestamp 1731220421
transform 1 0 3648 0 1 352
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5311_6
timestamp 1731220421
transform 1 0 3552 0 -1 576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5310_6
timestamp 1731220421
transform 1 0 3416 0 -1 576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5309_6
timestamp 1731220421
transform 1 0 3280 0 -1 576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5308_6
timestamp 1731220421
transform 1 0 3000 0 1 708
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5307_6
timestamp 1731220421
transform 1 0 2768 0 1 708
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5306_6
timestamp 1731220421
transform 1 0 2616 0 -1 932
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5305_6
timestamp 1731220421
transform 1 0 2896 0 -1 932
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5304_6
timestamp 1731220421
transform 1 0 3088 0 1 960
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5303_6
timestamp 1731220421
transform 1 0 2928 0 -1 1208
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5302_6
timestamp 1731220421
transform 1 0 2888 0 1 1208
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5301_6
timestamp 1731220421
transform 1 0 3072 0 1 1208
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5300_6
timestamp 1731220421
transform 1 0 3264 0 1 1208
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5299_6
timestamp 1731220421
transform 1 0 3224 0 -1 1432
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5298_6
timestamp 1731220421
transform 1 0 3088 0 -1 1432
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5297_6
timestamp 1731220421
transform 1 0 2952 0 -1 1432
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5296_6
timestamp 1731220421
transform 1 0 2816 0 -1 1432
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5295_6
timestamp 1731220421
transform 1 0 2680 0 -1 1432
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5294_6
timestamp 1731220421
transform 1 0 2544 0 -1 1432
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5293_6
timestamp 1731220421
transform 1 0 2536 0 1 1444
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5292_6
timestamp 1731220421
transform 1 0 2400 0 1 1444
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5291_6
timestamp 1731220421
transform 1 0 2672 0 1 1444
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5290_6
timestamp 1731220421
transform 1 0 2808 0 1 1444
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5289_6
timestamp 1731220421
transform 1 0 2944 0 1 1444
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5288_6
timestamp 1731220421
transform 1 0 3080 0 1 1444
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5287_6
timestamp 1731220421
transform 1 0 3488 0 1 1444
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5286_6
timestamp 1731220421
transform 1 0 3352 0 1 1444
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5285_6
timestamp 1731220421
transform 1 0 3216 0 1 1444
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5284_6
timestamp 1731220421
transform 1 0 3072 0 -1 1680
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5283_6
timestamp 1731220421
transform 1 0 2912 0 -1 1680
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5282_6
timestamp 1731220421
transform 1 0 2760 0 -1 1680
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5281_6
timestamp 1731220421
transform 1 0 3392 0 -1 1680
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5280_6
timestamp 1731220421
transform 1 0 3232 0 -1 1680
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5279_6
timestamp 1731220421
transform 1 0 3200 0 1 1692
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5278_6
timestamp 1731220421
transform 1 0 3048 0 1 1692
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5277_6
timestamp 1731220421
transform 1 0 2896 0 1 1692
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5276_6
timestamp 1731220421
transform 1 0 3648 0 1 1692
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5275_6
timestamp 1731220421
transform 1 0 3512 0 1 1692
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5274_6
timestamp 1731220421
transform 1 0 3352 0 1 1692
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5273_6
timestamp 1731220421
transform 1 0 3240 0 -1 1928
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5272_6
timestamp 1731220421
transform 1 0 3104 0 -1 1928
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5271_6
timestamp 1731220421
transform 1 0 3376 0 -1 1928
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5270_6
timestamp 1731220421
transform 1 0 3512 0 -1 1928
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5269_6
timestamp 1731220421
transform 1 0 3648 0 -1 1928
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5268_6
timestamp 1731220421
transform 1 0 3856 0 1 1840
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5267_6
timestamp 1731220421
transform 1 0 3856 0 -1 2064
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5266_6
timestamp 1731220421
transform 1 0 3992 0 -1 2064
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5265_6
timestamp 1731220421
transform 1 0 4128 0 -1 2064
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5264_6
timestamp 1731220421
transform 1 0 4264 0 -1 2064
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5263_6
timestamp 1731220421
transform 1 0 4400 0 -1 2064
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5262_6
timestamp 1731220421
transform 1 0 4400 0 1 2084
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5261_6
timestamp 1731220421
transform 1 0 4264 0 1 2084
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5260_6
timestamp 1731220421
transform 1 0 4128 0 1 2084
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5259_6
timestamp 1731220421
transform 1 0 3992 0 1 2084
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5258_6
timestamp 1731220421
transform 1 0 3856 0 1 2084
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5257_6
timestamp 1731220421
transform 1 0 3856 0 -1 2312
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5256_6
timestamp 1731220421
transform 1 0 3648 0 1 2128
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5255_6
timestamp 1731220421
transform 1 0 3648 0 -1 2352
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5254_6
timestamp 1731220421
transform 1 0 3440 0 -1 2352
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5253_6
timestamp 1731220421
transform 1 0 3208 0 -1 2352
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5252_6
timestamp 1731220421
transform 1 0 2976 0 -1 2352
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5251_6
timestamp 1731220421
transform 1 0 2736 0 -1 2352
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5250_6
timestamp 1731220421
transform 1 0 3648 0 1 2360
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5249_6
timestamp 1731220421
transform 1 0 3464 0 1 2360
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5248_6
timestamp 1731220421
transform 1 0 3280 0 1 2360
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5247_6
timestamp 1731220421
transform 1 0 3096 0 1 2360
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5246_6
timestamp 1731220421
transform 1 0 2904 0 1 2360
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5245_6
timestamp 1731220421
transform 1 0 3432 0 -1 2600
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5244_6
timestamp 1731220421
transform 1 0 3296 0 -1 2600
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5243_6
timestamp 1731220421
transform 1 0 3160 0 -1 2600
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5242_6
timestamp 1731220421
transform 1 0 3024 0 -1 2600
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5241_6
timestamp 1731220421
transform 1 0 2888 0 -1 2600
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5240_6
timestamp 1731220421
transform 1 0 3232 0 1 2604
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5239_6
timestamp 1731220421
transform 1 0 3088 0 1 2604
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5238_6
timestamp 1731220421
transform 1 0 2944 0 1 2604
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5237_6
timestamp 1731220421
transform 1 0 2800 0 1 2604
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5236_6
timestamp 1731220421
transform 1 0 2656 0 1 2604
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5235_6
timestamp 1731220421
transform 1 0 2632 0 -1 2828
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5234_6
timestamp 1731220421
transform 1 0 2800 0 -1 2828
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5233_6
timestamp 1731220421
transform 1 0 3136 0 -1 2828
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5232_6
timestamp 1731220421
transform 1 0 2968 0 -1 2828
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5231_6
timestamp 1731220421
transform 1 0 2936 0 1 2880
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5230_6
timestamp 1731220421
transform 1 0 2800 0 1 2880
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5229_6
timestamp 1731220421
transform 1 0 2752 0 -1 3104
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5228_6
timestamp 1731220421
transform 1 0 2616 0 -1 3104
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5227_6
timestamp 1731220421
transform 1 0 2984 0 1 3104
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5226_6
timestamp 1731220421
transform 1 0 3328 0 -1 3328
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5225_6
timestamp 1731220421
transform 1 0 2984 0 -1 3328
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5224_6
timestamp 1731220421
transform 1 0 2904 0 1 3352
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5223_6
timestamp 1731220421
transform 1 0 2528 0 1 3352
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5222_6
timestamp 1731220421
transform 1 0 2344 0 1 3352
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5221_6
timestamp 1731220421
transform 1 0 2168 0 1 3352
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5220_6
timestamp 1731220421
transform 1 0 2712 0 1 3352
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5219_6
timestamp 1731220421
transform 1 0 2752 0 -1 3580
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5218_6
timestamp 1731220421
transform 1 0 2616 0 -1 3580
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5217_6
timestamp 1731220421
transform 1 0 2480 0 -1 3580
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5216_6
timestamp 1731220421
transform 1 0 2344 0 -1 3580
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5215_6
timestamp 1731220421
transform 1 0 2208 0 -1 3580
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5214_6
timestamp 1731220421
transform 1 0 2576 0 1 3588
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5213_6
timestamp 1731220421
transform 1 0 2432 0 1 3588
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5212_6
timestamp 1731220421
transform 1 0 2288 0 1 3588
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5211_6
timestamp 1731220421
transform 1 0 2144 0 1 3588
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5210_6
timestamp 1731220421
transform 1 0 2008 0 1 3588
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5209_6
timestamp 1731220421
transform 1 0 2688 0 -1 3820
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5208_6
timestamp 1731220421
transform 1 0 2504 0 -1 3820
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5207_6
timestamp 1731220421
transform 1 0 2320 0 -1 3820
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5206_6
timestamp 1731220421
transform 1 0 2144 0 -1 3820
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5205_6
timestamp 1731220421
transform 1 0 1992 0 -1 3820
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5204_6
timestamp 1731220421
transform 1 0 1992 0 1 3820
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5203_6
timestamp 1731220421
transform 1 0 1784 0 1 3776
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5202_6
timestamp 1731220421
transform 1 0 1784 0 -1 4000
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5201_6
timestamp 1731220421
transform 1 0 1584 0 -1 4000
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5200_6
timestamp 1731220421
transform 1 0 1512 0 1 4000
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5199_6
timestamp 1731220421
transform 1 0 1648 0 1 4000
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5198_6
timestamp 1731220421
transform 1 0 1784 0 1 4000
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5197_6
timestamp 1731220421
transform 1 0 1648 0 -1 4224
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5196_6
timestamp 1731220421
transform 1 0 1784 0 -1 4224
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5195_6
timestamp 1731220421
transform 1 0 1992 0 1 4148
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5194_6
timestamp 1731220421
transform 1 0 1992 0 -1 4376
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5193_6
timestamp 1731220421
transform 1 0 2168 0 -1 4376
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5192_6
timestamp 1731220421
transform 1 0 2368 0 -1 4376
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5191_6
timestamp 1731220421
transform 1 0 2264 0 1 4388
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5190_6
timestamp 1731220421
transform 1 0 2512 0 1 4388
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5189_6
timestamp 1731220421
transform 1 0 2496 0 -1 4624
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5188_6
timestamp 1731220421
transform 1 0 2232 0 -1 4624
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5187_6
timestamp 1731220421
transform 1 0 2744 0 -1 4624
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5186_6
timestamp 1731220421
transform 1 0 2720 0 1 4628
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5185_6
timestamp 1731220421
transform 1 0 2544 0 1 4628
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5184_6
timestamp 1731220421
transform 1 0 3072 0 -1 4864
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5183_6
timestamp 1731220421
transform 1 0 3368 0 -1 4864
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5182_6
timestamp 1731220421
transform 1 0 3392 0 1 4872
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5181_6
timestamp 1731220421
transform 1 0 3176 0 -1 5104
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5180_6
timestamp 1731220421
transform 1 0 2944 0 -1 5104
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5179_6
timestamp 1731220421
transform 1 0 3096 0 1 5120
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5178_6
timestamp 1731220421
transform 1 0 3304 0 1 5120
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5177_6
timestamp 1731220421
transform 1 0 3296 0 -1 5348
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5176_6
timestamp 1731220421
transform 1 0 3088 0 -1 5348
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5175_6
timestamp 1731220421
transform 1 0 3504 0 -1 5348
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5174_6
timestamp 1731220421
transform 1 0 3424 0 1 5348
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5173_6
timestamp 1731220421
transform 1 0 3184 0 1 5348
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5172_6
timestamp 1731220421
transform 1 0 3648 0 1 5348
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5171_6
timestamp 1731220421
transform 1 0 3448 0 -1 5576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5170_6
timestamp 1731220421
transform 1 0 3232 0 -1 5576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5169_6
timestamp 1731220421
transform 1 0 3648 0 -1 5576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5168_6
timestamp 1731220421
transform 1 0 3616 0 1 5576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5167_6
timestamp 1731220421
transform 1 0 3440 0 1 5576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5166_6
timestamp 1731220421
transform 1 0 3272 0 1 5576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5165_6
timestamp 1731220421
transform 1 0 3104 0 1 5576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5164_6
timestamp 1731220421
transform 1 0 2928 0 1 5576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5163_6
timestamp 1731220421
transform 1 0 2744 0 1 5576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5162_6
timestamp 1731220421
transform 1 0 3016 0 -1 5576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5161_6
timestamp 1731220421
transform 1 0 2800 0 -1 5576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5160_6
timestamp 1731220421
transform 1 0 2696 0 1 5348
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5159_6
timestamp 1731220421
transform 1 0 2944 0 1 5348
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5158_6
timestamp 1731220421
transform 1 0 2888 0 -1 5348
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5157_6
timestamp 1731220421
transform 1 0 2888 0 1 5120
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5156_6
timestamp 1731220421
transform 1 0 2680 0 1 5120
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5155_6
timestamp 1731220421
transform 1 0 2720 0 -1 5104
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5154_6
timestamp 1731220421
transform 1 0 3120 0 1 4872
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5153_6
timestamp 1731220421
transform 1 0 2792 0 -1 4864
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5152_6
timestamp 1731220421
transform 1 0 2528 0 -1 4864
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5151_6
timestamp 1731220421
transform 1 0 2296 0 -1 4864
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5150_6
timestamp 1731220421
transform 1 0 2368 0 1 4628
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5149_6
timestamp 1731220421
transform 1 0 2192 0 1 4628
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5148_6
timestamp 1731220421
transform 1 0 2016 0 1 4628
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5147_6
timestamp 1731220421
transform 1 0 1992 0 -1 4624
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5146_6
timestamp 1731220421
transform 1 0 1784 0 1 4460
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5145_6
timestamp 1731220421
transform 1 0 1568 0 1 4460
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5144_6
timestamp 1731220421
transform 1 0 1328 0 1 4460
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5143_6
timestamp 1731220421
transform 1 0 1464 0 -1 4460
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5142_6
timestamp 1731220421
transform 1 0 1688 0 -1 4460
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5141_6
timestamp 1731220421
transform 1 0 1664 0 1 4232
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5140_6
timestamp 1731220421
transform 1 0 1528 0 1 4232
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5139_6
timestamp 1731220421
transform 1 0 1392 0 1 4232
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5138_6
timestamp 1731220421
transform 1 0 1512 0 -1 4224
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5137_6
timestamp 1731220421
transform 1 0 1376 0 -1 4224
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5136_6
timestamp 1731220421
transform 1 0 1376 0 1 4000
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5135_6
timestamp 1731220421
transform 1 0 1240 0 1 4000
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5134_6
timestamp 1731220421
transform 1 0 1368 0 -1 4000
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5133_6
timestamp 1731220421
transform 1 0 1152 0 -1 4000
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5132_6
timestamp 1731220421
transform 1 0 1192 0 1 3776
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5131_6
timestamp 1731220421
transform 1 0 1496 0 1 3776
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5130_6
timestamp 1731220421
transform 1 0 1312 0 -1 3764
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5129_6
timestamp 1731220421
transform 1 0 1032 0 -1 3764
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5128_6
timestamp 1731220421
transform 1 0 1208 0 1 3524
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5127_6
timestamp 1731220421
transform 1 0 1064 0 1 3524
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5126_6
timestamp 1731220421
transform 1 0 920 0 1 3524
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5125_6
timestamp 1731220421
transform 1 0 944 0 -1 3504
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5124_6
timestamp 1731220421
transform 1 0 808 0 -1 3504
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5123_6
timestamp 1731220421
transform 1 0 776 0 1 3524
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5122_6
timestamp 1731220421
transform 1 0 632 0 1 3524
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5121_6
timestamp 1731220421
transform 1 0 488 0 1 3524
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5120_6
timestamp 1731220421
transform 1 0 488 0 -1 3764
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5119_6
timestamp 1731220421
transform 1 0 216 0 -1 3764
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5118_6
timestamp 1731220421
transform 1 0 760 0 -1 3764
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5117_6
timestamp 1731220421
transform 1 0 896 0 1 3776
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5116_6
timestamp 1731220421
transform 1 0 616 0 1 3776
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5115_6
timestamp 1731220421
transform 1 0 352 0 1 3776
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5114_6
timestamp 1731220421
transform 1 0 128 0 1 3776
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5113_6
timestamp 1731220421
transform 1 0 128 0 -1 4000
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5112_6
timestamp 1731220421
transform 1 0 296 0 -1 4000
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5111_6
timestamp 1731220421
transform 1 0 504 0 -1 4000
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5110_6
timestamp 1731220421
transform 1 0 720 0 -1 4000
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5109_6
timestamp 1731220421
transform 1 0 936 0 -1 4000
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5108_6
timestamp 1731220421
transform 1 0 832 0 1 4000
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5107_6
timestamp 1731220421
transform 1 0 696 0 1 4000
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5106_6
timestamp 1731220421
transform 1 0 560 0 1 4000
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5105_6
timestamp 1731220421
transform 1 0 1104 0 1 4000
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5104_6
timestamp 1731220421
transform 1 0 968 0 1 4000
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5103_6
timestamp 1731220421
transform 1 0 832 0 -1 4224
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5102_6
timestamp 1731220421
transform 1 0 696 0 -1 4224
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5101_6
timestamp 1731220421
transform 1 0 968 0 -1 4224
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5100_6
timestamp 1731220421
transform 1 0 1104 0 -1 4224
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_599_6
timestamp 1731220421
transform 1 0 1240 0 -1 4224
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_598_6
timestamp 1731220421
transform 1 0 1256 0 1 4232
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_597_6
timestamp 1731220421
transform 1 0 1120 0 1 4232
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_596_6
timestamp 1731220421
transform 1 0 984 0 1 4232
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_595_6
timestamp 1731220421
transform 1 0 848 0 1 4232
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_594_6
timestamp 1731220421
transform 1 0 712 0 1 4232
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_593_6
timestamp 1731220421
transform 1 0 1248 0 -1 4460
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_592_6
timestamp 1731220421
transform 1 0 1040 0 -1 4460
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_591_6
timestamp 1731220421
transform 1 0 840 0 -1 4460
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_590_6
timestamp 1731220421
transform 1 0 656 0 -1 4460
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_589_6
timestamp 1731220421
transform 1 0 480 0 -1 4460
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_588_6
timestamp 1731220421
transform 1 0 1096 0 1 4460
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_587_6
timestamp 1731220421
transform 1 0 872 0 1 4460
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_586_6
timestamp 1731220421
transform 1 0 648 0 1 4460
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_585_6
timestamp 1731220421
transform 1 0 440 0 1 4460
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_584_6
timestamp 1731220421
transform 1 0 248 0 1 4460
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_583_6
timestamp 1731220421
transform 1 0 672 0 -1 4696
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_582_6
timestamp 1731220421
transform 1 0 536 0 -1 4696
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_581_6
timestamp 1731220421
transform 1 0 400 0 -1 4696
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_580_6
timestamp 1731220421
transform 1 0 264 0 -1 4696
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_579_6
timestamp 1731220421
transform 1 0 128 0 -1 4696
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_578_6
timestamp 1731220421
transform 1 0 672 0 1 4700
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_577_6
timestamp 1731220421
transform 1 0 536 0 1 4700
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_576_6
timestamp 1731220421
transform 1 0 400 0 1 4700
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_575_6
timestamp 1731220421
transform 1 0 264 0 1 4700
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_574_6
timestamp 1731220421
transform 1 0 128 0 1 4700
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_573_6
timestamp 1731220421
transform 1 0 128 0 -1 4936
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_572_6
timestamp 1731220421
transform 1 0 264 0 -1 4936
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_571_6
timestamp 1731220421
transform 1 0 672 0 -1 4936
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_570_6
timestamp 1731220421
transform 1 0 536 0 -1 4936
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_569_6
timestamp 1731220421
transform 1 0 400 0 -1 4936
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_568_6
timestamp 1731220421
transform 1 0 376 0 1 4964
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_567_6
timestamp 1731220421
transform 1 0 152 0 1 4964
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_566_6
timestamp 1731220421
transform 1 0 1192 0 1 4964
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_565_6
timestamp 1731220421
transform 1 0 896 0 1 4964
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_564_6
timestamp 1731220421
transform 1 0 624 0 1 4964
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_563_6
timestamp 1731220421
transform 1 0 592 0 -1 5196
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_562_6
timestamp 1731220421
transform 1 0 416 0 -1 5196
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_561_6
timestamp 1731220421
transform 1 0 776 0 -1 5196
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_560_6
timestamp 1731220421
transform 1 0 968 0 -1 5196
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_559_6
timestamp 1731220421
transform 1 0 1168 0 -1 5196
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_558_6
timestamp 1731220421
transform 1 0 1184 0 1 5196
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_557_6
timestamp 1731220421
transform 1 0 1024 0 1 5196
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_556_6
timestamp 1731220421
transform 1 0 872 0 1 5196
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_555_6
timestamp 1731220421
transform 1 0 720 0 1 5196
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_554_6
timestamp 1731220421
transform 1 0 688 0 -1 5420
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_553_6
timestamp 1731220421
transform 1 0 824 0 -1 5420
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_552_6
timestamp 1731220421
transform 1 0 960 0 -1 5420
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_551_6
timestamp 1731220421
transform 1 0 1096 0 -1 5420
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_550_6
timestamp 1731220421
transform 1 0 1776 0 -1 5420
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_549_6
timestamp 1731220421
transform 1 0 1640 0 -1 5420
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_548_6
timestamp 1731220421
transform 1 0 1504 0 -1 5420
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_547_6
timestamp 1731220421
transform 1 0 1432 0 1 5420
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_546_6
timestamp 1731220421
transform 1 0 1288 0 1 5420
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_545_6
timestamp 1731220421
transform 1 0 1720 0 1 5420
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_544_6
timestamp 1731220421
transform 1 0 1576 0 1 5420
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_543_6
timestamp 1731220421
transform 1 0 1352 0 -1 5644
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_542_6
timestamp 1731220421
transform 1 0 1576 0 -1 5644
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_541_6
timestamp 1731220421
transform 1 0 1784 0 -1 5644
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_540_6
timestamp 1731220421
transform 1 0 1992 0 1 5576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_539_6
timestamp 1731220421
transform 1 0 2168 0 1 5576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_538_6
timestamp 1731220421
transform 1 0 2368 0 1 5576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_537_6
timestamp 1731220421
transform 1 0 2560 0 1 5576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_536_6
timestamp 1731220421
transform 1 0 2576 0 -1 5576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_535_6
timestamp 1731220421
transform 1 0 2344 0 -1 5576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_534_6
timestamp 1731220421
transform 1 0 2448 0 1 5348
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_533_6
timestamp 1731220421
transform 1 0 2288 0 -1 5348
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_532_6
timestamp 1731220421
transform 1 0 2688 0 -1 5348
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_531_6
timestamp 1731220421
transform 1 0 2488 0 -1 5348
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_530_6
timestamp 1731220421
transform 1 0 2472 0 1 5120
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_529_6
timestamp 1731220421
transform 1 0 2272 0 1 5120
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_528_6
timestamp 1731220421
transform 1 0 2088 0 -1 5104
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_527_6
timestamp 1731220421
transform 1 0 2296 0 -1 5104
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_526_6
timestamp 1731220421
transform 1 0 2504 0 -1 5104
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_525_6
timestamp 1731220421
transform 1 0 2856 0 1 4872
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_524_6
timestamp 1731220421
transform 1 0 2616 0 1 4872
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_523_6
timestamp 1731220421
transform 1 0 2416 0 1 4872
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_522_6
timestamp 1731220421
transform 1 0 2264 0 1 4872
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_521_6
timestamp 1731220421
transform 1 0 2128 0 1 4872
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_520_6
timestamp 1731220421
transform 1 0 1992 0 1 4872
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_519_6
timestamp 1731220421
transform 1 0 1784 0 1 4964
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_518_6
timestamp 1731220421
transform 1 0 1496 0 1 4964
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_517_6
timestamp 1731220421
transform 1 0 1368 0 -1 5196
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_516_6
timestamp 1731220421
transform 1 0 1784 0 -1 5196
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_515_6
timestamp 1731220421
transform 1 0 1576 0 -1 5196
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_514_6
timestamp 1731220421
transform 1 0 1520 0 1 5196
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_513_6
timestamp 1731220421
transform 1 0 1352 0 1 5196
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_512_6
timestamp 1731220421
transform 1 0 1368 0 -1 5420
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_511_6
timestamp 1731220421
transform 1 0 1232 0 -1 5420
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_510_6
timestamp 1731220421
transform 1 0 1144 0 1 5420
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_59_6
timestamp 1731220421
transform 1 0 1008 0 1 5420
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_58_6
timestamp 1731220421
transform 1 0 872 0 1 5420
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_57_6
timestamp 1731220421
transform 1 0 1128 0 -1 5644
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_56_6
timestamp 1731220421
transform 1 0 912 0 -1 5644
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_55_6
timestamp 1731220421
transform 1 0 704 0 -1 5644
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_54_6
timestamp 1731220421
transform 1 0 504 0 -1 5644
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_53_6
timestamp 1731220421
transform 1 0 312 0 -1 5644
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_52_6
timestamp 1731220421
transform 1 0 400 0 1 5644
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_51_6
timestamp 1731220421
transform 1 0 264 0 1 5644
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_50_6
timestamp 1731220421
transform 1 0 128 0 1 5644
box 3 5 132 108
<< end >>
