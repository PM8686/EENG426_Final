magic
tech sky130l
timestamp 1731220359
<< m1 >>
rect 1608 3963 1612 3991
rect 1600 3915 1604 3955
rect 2256 3875 2260 3975
rect 440 3811 444 3839
rect 568 3811 572 3839
rect 1472 3811 1476 3839
rect 2768 3819 2772 3847
rect 2960 3819 2964 3863
rect 2328 3715 2332 3739
rect 2296 3663 2300 3691
rect 728 3591 732 3619
rect 2440 3551 2444 3575
rect 1312 3475 1316 3503
rect 2192 3503 2196 3531
rect 2432 3503 2436 3543
rect 2760 3503 2764 3531
rect 2976 3395 2980 3423
rect 2352 3331 2356 3387
rect 608 3267 612 3295
rect 2368 3219 2372 3243
rect 1232 3163 1236 3191
rect 864 3111 868 3155
rect 1216 3111 1220 3139
rect 1192 2999 1196 3027
rect 2272 3007 2276 3035
rect 1288 2843 1292 2943
rect 3800 2931 3804 3035
rect 2280 2899 2284 2927
rect 3792 2691 3796 2719
rect 1120 2623 1124 2651
rect 2880 2579 2884 2607
rect 3752 2419 3756 2447
rect 440 2179 444 2207
rect 584 2179 588 2207
rect 760 2179 764 2207
rect 1400 2179 1404 2207
rect 1552 2179 1556 2207
rect 784 2131 788 2171
rect 1976 2163 1980 2187
rect 792 2131 796 2151
rect 1072 2059 1076 2159
rect 1216 2131 1220 2159
rect 1480 2131 1484 2159
rect 2744 2067 2748 2095
rect 1504 2027 1508 2051
rect 648 1855 652 1899
rect 840 1871 844 1899
rect 1032 1871 1036 1899
rect 696 1823 700 1851
rect 2272 1843 2276 1871
rect 2376 1843 2380 1871
rect 3624 1843 3628 1895
rect 2216 1735 2220 1763
rect 2400 1735 2404 1763
rect 2968 1735 2972 1763
rect 656 1407 660 1435
rect 1096 1383 1100 1435
rect 3504 1299 3508 1351
rect 928 1199 932 1227
rect 1528 1199 1532 1227
rect 2792 1187 2796 1215
rect 3640 1187 3644 1215
rect 1704 1091 1708 1115
rect 1456 1035 1460 1083
rect 2424 1023 2428 1067
rect 2800 1023 2804 1051
rect 408 931 412 959
rect 2784 859 2788 887
rect 432 779 436 807
rect 792 779 796 807
rect 1592 731 1596 759
rect 3024 755 3028 783
rect 3336 703 3340 731
rect 3488 703 3492 731
rect 960 627 964 655
rect 1160 627 1164 655
rect 872 579 876 607
rect 968 579 972 619
rect 2104 571 2108 619
rect 2360 591 2364 619
rect 2640 539 2644 567
rect 1240 427 1244 483
rect 1528 463 1532 483
rect 3456 435 3460 463
rect 784 395 788 423
rect 888 395 892 423
rect 1096 395 1100 423
rect 824 231 828 259
rect 832 231 836 275
rect 2800 231 2804 259
<< m2c >>
rect 2124 4005 2128 4009
rect 2220 4007 2224 4011
rect 2316 4007 2320 4011
rect 1608 3991 1612 3995
rect 2256 3975 2260 3979
rect 1608 3959 1612 3963
rect 1668 3959 1672 3963
rect 1764 3959 1768 3963
rect 1860 3959 1864 3963
rect 1956 3959 1960 3963
rect 1572 3955 1576 3959
rect 1600 3955 1604 3959
rect 252 3943 256 3947
rect 348 3943 352 3947
rect 444 3943 448 3947
rect 548 3943 552 3947
rect 668 3943 672 3947
rect 796 3943 800 3947
rect 924 3943 928 3947
rect 1052 3943 1056 3947
rect 1180 3943 1184 3947
rect 1308 3943 1312 3947
rect 1436 3943 1440 3947
rect 1564 3943 1568 3947
rect 1700 3943 1704 3947
rect 1600 3911 1604 3915
rect 2212 3871 2216 3875
rect 2256 3871 2260 3875
rect 2340 3871 2344 3875
rect 2468 3871 2472 3875
rect 2604 3871 2608 3875
rect 2740 3871 2744 3875
rect 3004 3871 3008 3875
rect 3124 3871 3128 3875
rect 3244 3871 3248 3875
rect 3356 3871 3360 3875
rect 3460 3871 3464 3875
rect 3572 3871 3576 3875
rect 3684 3871 3688 3875
rect 3796 3871 3800 3875
rect 2876 3867 2880 3871
rect 2960 3863 2964 3867
rect 2260 3847 2264 3851
rect 2396 3847 2400 3851
rect 2540 3847 2544 3851
rect 2700 3847 2704 3851
rect 2768 3847 2772 3851
rect 2876 3847 2880 3851
rect 440 3839 444 3843
rect 568 3839 572 3843
rect 1472 3839 1476 3843
rect 2768 3815 2772 3819
rect 3068 3847 3072 3851
rect 3276 3847 3280 3851
rect 3492 3847 3496 3851
rect 3708 3847 3712 3851
rect 2960 3815 2964 3819
rect 388 3807 392 3811
rect 440 3807 444 3811
rect 508 3807 512 3811
rect 568 3807 572 3811
rect 772 3807 776 3811
rect 900 3807 904 3811
rect 1028 3807 1032 3811
rect 1156 3807 1160 3811
rect 1284 3807 1288 3811
rect 1412 3807 1416 3811
rect 1472 3807 1476 3811
rect 636 3803 640 3807
rect 1540 3803 1544 3807
rect 556 3787 560 3791
rect 668 3787 672 3791
rect 788 3787 792 3791
rect 916 3787 920 3791
rect 1052 3787 1056 3791
rect 1196 3787 1200 3791
rect 1340 3785 1344 3789
rect 1484 3787 1488 3791
rect 1636 3787 1640 3791
rect 2328 3739 2332 3743
rect 2244 3711 2248 3715
rect 2328 3711 2332 3715
rect 2428 3711 2432 3715
rect 2612 3711 2616 3715
rect 2796 3711 2800 3715
rect 2988 3711 2992 3715
rect 3180 3711 3184 3715
rect 3372 3711 3376 3715
rect 3764 3711 3768 3715
rect 3564 3707 3568 3711
rect 2180 3691 2184 3695
rect 2296 3691 2300 3695
rect 2404 3691 2408 3695
rect 2636 3691 2640 3695
rect 2868 3691 2872 3695
rect 3100 3689 3104 3693
rect 3332 3691 3336 3695
rect 3564 3691 3568 3695
rect 3804 3691 3808 3695
rect 2296 3659 2300 3663
rect 644 3643 648 3647
rect 740 3643 744 3647
rect 844 3643 848 3647
rect 964 3643 968 3647
rect 1092 3643 1096 3647
rect 1236 3643 1240 3647
rect 1388 3643 1392 3647
rect 1548 3643 1552 3647
rect 548 3639 552 3643
rect 1708 3639 1712 3643
rect 388 3617 392 3621
rect 516 3619 520 3623
rect 660 3619 664 3623
rect 728 3619 732 3623
rect 812 3619 816 3623
rect 980 3619 984 3623
rect 1148 3619 1152 3623
rect 1316 3619 1320 3623
rect 1492 3617 1496 3621
rect 1668 3619 1672 3623
rect 1844 3619 1848 3623
rect 728 3587 732 3591
rect 2440 3575 2444 3579
rect 2244 3547 2248 3551
rect 2440 3547 2444 3551
rect 2508 3547 2512 3551
rect 2636 3547 2640 3551
rect 2772 3547 2776 3551
rect 2908 3547 2912 3551
rect 3052 3547 3056 3551
rect 3196 3547 3200 3551
rect 3348 3547 3352 3551
rect 3508 3547 3512 3551
rect 2380 3543 2384 3547
rect 2432 3543 2436 3547
rect 3676 3543 3680 3547
rect 2156 3531 2160 3535
rect 2192 3531 2196 3535
rect 2324 3531 2328 3535
rect 1312 3503 1316 3507
rect 2192 3499 2196 3503
rect 2500 3531 2504 3535
rect 2684 3531 2688 3535
rect 2760 3531 2764 3535
rect 2868 3531 2872 3535
rect 3052 3533 3056 3537
rect 3228 3531 3232 3535
rect 3404 3531 3408 3535
rect 3572 3531 3576 3535
rect 3740 3531 3744 3535
rect 3892 3531 3896 3535
rect 2432 3499 2436 3503
rect 2760 3499 2764 3503
rect 356 3471 360 3475
rect 516 3471 520 3475
rect 692 3471 696 3475
rect 868 3471 872 3475
rect 1052 3471 1056 3475
rect 1228 3471 1232 3475
rect 1312 3471 1316 3475
rect 1404 3471 1408 3475
rect 1756 3471 1760 3475
rect 1932 3471 1936 3475
rect 212 3467 216 3471
rect 1580 3467 1584 3471
rect 188 3447 192 3451
rect 372 3447 376 3451
rect 588 3447 592 3451
rect 804 3447 808 3451
rect 1012 3447 1016 3451
rect 1212 3447 1216 3451
rect 1404 3447 1408 3451
rect 1588 3447 1592 3451
rect 1772 3447 1776 3451
rect 1956 3447 1960 3451
rect 2976 3423 2980 3427
rect 2180 3391 2184 3395
rect 2548 3391 2552 3395
rect 2732 3391 2736 3395
rect 2916 3391 2920 3395
rect 2976 3391 2980 3395
rect 3100 3391 3104 3395
rect 3276 3391 3280 3395
rect 3460 3391 3464 3395
rect 3828 3391 3832 3395
rect 2352 3387 2356 3391
rect 2364 3387 2368 3391
rect 3644 3387 3648 3391
rect 2124 3359 2128 3363
rect 2268 3359 2272 3363
rect 2412 3359 2416 3363
rect 2564 3359 2568 3363
rect 2708 3359 2712 3363
rect 2852 3359 2856 3363
rect 2988 3359 2992 3363
rect 3132 3359 3136 3363
rect 3276 3359 3280 3363
rect 3428 3359 3432 3363
rect 3588 3359 3592 3363
rect 3748 3359 3752 3363
rect 3892 3359 3896 3363
rect 2352 3327 2356 3331
rect 284 3311 288 3315
rect 428 3311 432 3315
rect 588 3311 592 3315
rect 756 3311 760 3315
rect 924 3311 928 3315
rect 1100 3311 1104 3315
rect 1268 3311 1272 3315
rect 1436 3311 1440 3315
rect 1756 3311 1760 3315
rect 1924 3311 1928 3315
rect 188 3307 192 3311
rect 1596 3307 1600 3311
rect 188 3295 192 3299
rect 332 3293 336 3297
rect 516 3295 520 3299
rect 608 3295 612 3299
rect 716 3295 720 3299
rect 924 3295 928 3299
rect 1132 3295 1136 3299
rect 1348 3295 1352 3299
rect 1572 3295 1576 3299
rect 1796 3295 1800 3299
rect 608 3263 612 3267
rect 2368 3243 2372 3247
rect 2164 3215 2168 3219
rect 2368 3215 2372 3219
rect 2452 3215 2456 3219
rect 2628 3215 2632 3219
rect 2836 3215 2840 3219
rect 3068 3215 3072 3219
rect 3580 3215 3584 3219
rect 3844 3215 3848 3219
rect 2300 3211 2304 3215
rect 3316 3211 3320 3215
rect 2124 3199 2128 3203
rect 2220 3197 2224 3201
rect 2316 3199 2320 3203
rect 2412 3199 2416 3203
rect 2508 3199 2512 3203
rect 2604 3199 2608 3203
rect 2700 3199 2704 3203
rect 2796 3199 2800 3203
rect 2892 3199 2896 3203
rect 2988 3199 2992 3203
rect 3084 3199 3088 3203
rect 3180 3199 3184 3203
rect 3276 3199 3280 3203
rect 3372 3199 3376 3203
rect 3492 3197 3496 3201
rect 3628 3199 3632 3203
rect 3772 3199 3776 3203
rect 3892 3199 3896 3203
rect 1232 3191 1236 3195
rect 188 3159 192 3163
rect 500 3159 504 3163
rect 668 3159 672 3163
rect 1020 3159 1024 3163
rect 1196 3159 1200 3163
rect 1232 3159 1236 3163
rect 1380 3159 1384 3163
rect 1748 3159 1752 3163
rect 340 3155 344 3159
rect 844 3155 848 3159
rect 864 3155 868 3159
rect 1564 3155 1568 3159
rect 364 3139 368 3143
rect 492 3139 496 3143
rect 636 3139 640 3143
rect 796 3139 800 3143
rect 956 3139 960 3143
rect 1116 3139 1120 3143
rect 1216 3139 1220 3143
rect 1276 3139 1280 3143
rect 1444 3139 1448 3143
rect 1612 3139 1616 3143
rect 1780 3139 1784 3143
rect 864 3107 868 3111
rect 1216 3107 1220 3111
rect 2124 3051 2128 3055
rect 2388 3051 2392 3055
rect 2964 3051 2968 3055
rect 3260 3051 3264 3055
rect 3556 3051 3560 3055
rect 3852 3051 3856 3055
rect 2676 3047 2680 3051
rect 2124 3035 2128 3039
rect 2272 3035 2276 3039
rect 2436 3035 2440 3039
rect 2756 3035 2760 3039
rect 3052 3035 3056 3039
rect 3340 3035 3344 3039
rect 3628 3035 3632 3039
rect 3800 3035 3804 3039
rect 3892 3035 3896 3039
rect 1192 3027 1196 3031
rect 2272 3003 2276 3007
rect 556 2995 560 2999
rect 652 2995 656 2999
rect 756 2995 760 2999
rect 868 2995 872 2999
rect 1124 2995 1128 2999
rect 1192 2995 1196 2999
rect 1276 2995 1280 2999
rect 1436 2995 1440 2999
rect 1772 2995 1776 2999
rect 988 2991 992 2995
rect 1604 2991 1608 2995
rect 604 2973 608 2977
rect 700 2975 704 2979
rect 812 2975 816 2979
rect 940 2975 944 2979
rect 1076 2975 1080 2979
rect 1228 2975 1232 2979
rect 1380 2975 1384 2979
rect 1540 2975 1544 2979
rect 1708 2975 1712 2979
rect 1876 2975 1880 2979
rect 1288 2943 1292 2947
rect 2280 2927 2284 2931
rect 3800 2927 3804 2931
rect 2124 2895 2128 2899
rect 2280 2895 2284 2899
rect 2444 2895 2448 2899
rect 2756 2895 2760 2899
rect 3268 2895 3272 2899
rect 3492 2895 3496 2899
rect 3700 2895 3704 2899
rect 3892 2895 3896 2899
rect 3028 2891 3032 2895
rect 2124 2879 2128 2883
rect 2348 2879 2352 2883
rect 2588 2879 2592 2883
rect 2820 2879 2824 2883
rect 3044 2877 3048 2881
rect 3268 2879 3272 2883
rect 3484 2879 3488 2883
rect 3700 2879 3704 2883
rect 3892 2879 3896 2883
rect 1288 2839 1292 2843
rect 628 2831 632 2835
rect 748 2831 752 2835
rect 892 2831 896 2835
rect 1044 2831 1048 2835
rect 1204 2831 1208 2835
rect 1372 2831 1376 2835
rect 1724 2831 1728 2835
rect 1900 2831 1904 2835
rect 524 2827 528 2831
rect 1548 2827 1552 2831
rect 532 2811 536 2815
rect 628 2811 632 2815
rect 732 2811 736 2815
rect 852 2811 856 2815
rect 988 2811 992 2815
rect 1132 2811 1136 2815
rect 1292 2811 1296 2815
rect 1468 2811 1472 2815
rect 1652 2811 1656 2815
rect 1836 2811 1840 2815
rect 2124 2739 2128 2743
rect 2252 2739 2256 2743
rect 2420 2739 2424 2743
rect 2604 2739 2608 2743
rect 2788 2739 2792 2743
rect 3164 2739 3168 2743
rect 3348 2739 3352 2743
rect 3532 2739 3536 2743
rect 3724 2739 3728 2743
rect 2980 2735 2984 2739
rect 3892 2735 3896 2739
rect 2124 2721 2128 2725
rect 2244 2719 2248 2723
rect 2372 2719 2376 2723
rect 2500 2719 2504 2723
rect 2636 2719 2640 2723
rect 2780 2719 2784 2723
rect 2940 2719 2944 2723
rect 3116 2719 3120 2723
rect 3308 2719 3312 2723
rect 3508 2719 3512 2723
rect 3708 2719 3712 2723
rect 3792 2719 3796 2723
rect 3892 2719 3896 2723
rect 3792 2687 3796 2691
rect 676 2671 680 2675
rect 796 2671 800 2675
rect 932 2671 936 2675
rect 1068 2671 1072 2675
rect 1212 2671 1216 2675
rect 1364 2671 1368 2675
rect 1676 2671 1680 2675
rect 1836 2671 1840 2675
rect 564 2667 568 2671
rect 1516 2667 1520 2671
rect 420 2649 424 2653
rect 540 2651 544 2655
rect 668 2651 672 2655
rect 804 2651 808 2655
rect 948 2651 952 2655
rect 1084 2651 1088 2655
rect 1120 2651 1124 2655
rect 1220 2651 1224 2655
rect 1356 2651 1360 2655
rect 1484 2651 1488 2655
rect 1620 2651 1624 2655
rect 1756 2651 1760 2655
rect 1120 2619 1124 2623
rect 2880 2607 2884 2611
rect 2284 2575 2288 2579
rect 2388 2575 2392 2579
rect 2500 2575 2504 2579
rect 2612 2575 2616 2579
rect 2724 2575 2728 2579
rect 2844 2575 2848 2579
rect 2880 2575 2884 2579
rect 2964 2575 2968 2579
rect 3204 2575 3208 2579
rect 3084 2571 3088 2575
rect 2436 2557 2440 2561
rect 2548 2555 2552 2559
rect 2668 2555 2672 2559
rect 2796 2555 2800 2559
rect 2924 2555 2928 2559
rect 3044 2555 3048 2559
rect 3164 2555 3168 2559
rect 3284 2555 3288 2559
rect 3412 2555 3416 2559
rect 3540 2553 3544 2557
rect 340 2515 344 2519
rect 500 2515 504 2519
rect 660 2515 664 2519
rect 820 2515 824 2519
rect 972 2515 976 2519
rect 1116 2515 1120 2519
rect 1252 2515 1256 2519
rect 1388 2515 1392 2519
rect 1516 2515 1520 2519
rect 1644 2515 1648 2519
rect 1780 2515 1784 2519
rect 188 2511 192 2515
rect 188 2483 192 2487
rect 284 2483 288 2487
rect 380 2483 384 2487
rect 476 2483 480 2487
rect 572 2483 576 2487
rect 3752 2447 3756 2451
rect 2588 2415 2592 2419
rect 2764 2415 2768 2419
rect 2932 2415 2936 2419
rect 3100 2415 3104 2419
rect 3260 2415 3264 2419
rect 3412 2415 3416 2419
rect 3556 2415 3560 2419
rect 3708 2415 3712 2419
rect 3752 2415 3756 2419
rect 3860 2411 3864 2415
rect 2660 2385 2664 2389
rect 2868 2387 2872 2391
rect 3060 2387 3064 2391
rect 3244 2385 3248 2389
rect 3412 2387 3416 2391
rect 3572 2387 3576 2391
rect 3732 2387 3736 2391
rect 3892 2387 3896 2391
rect 188 2331 192 2335
rect 308 2331 312 2335
rect 468 2331 472 2335
rect 628 2331 632 2335
rect 940 2331 944 2335
rect 1092 2331 1096 2335
rect 1236 2331 1240 2335
rect 1380 2331 1384 2335
rect 788 2327 792 2331
rect 1532 2327 1536 2331
rect 188 2315 192 2319
rect 316 2315 320 2319
rect 476 2315 480 2319
rect 636 2315 640 2319
rect 796 2315 800 2319
rect 948 2315 952 2319
rect 1100 2315 1104 2319
rect 1252 2315 1256 2319
rect 1404 2315 1408 2319
rect 1556 2315 1560 2319
rect 2124 2235 2128 2239
rect 2220 2235 2224 2239
rect 2324 2235 2328 2239
rect 2468 2235 2472 2239
rect 2628 2235 2632 2239
rect 2964 2235 2968 2239
rect 3124 2235 3128 2239
rect 3284 2235 3288 2239
rect 3436 2235 3440 2239
rect 3588 2235 3592 2239
rect 3748 2235 3752 2239
rect 2796 2231 2800 2235
rect 2124 2219 2128 2223
rect 2228 2219 2232 2223
rect 2372 2219 2376 2223
rect 2524 2219 2528 2223
rect 2676 2219 2680 2223
rect 2836 2219 2840 2223
rect 2988 2219 2992 2223
rect 3132 2219 3136 2223
rect 3276 2219 3280 2223
rect 3420 2219 3424 2223
rect 3572 2219 3576 2223
rect 440 2207 444 2211
rect 584 2207 588 2211
rect 760 2207 764 2211
rect 1400 2207 1404 2211
rect 1552 2207 1556 2211
rect 276 2175 280 2179
rect 404 2175 408 2179
rect 440 2175 444 2179
rect 548 2175 552 2179
rect 584 2175 588 2179
rect 700 2175 704 2179
rect 760 2175 764 2179
rect 1012 2175 1016 2179
rect 1172 2175 1176 2179
rect 1332 2175 1336 2179
rect 1400 2175 1404 2179
rect 1492 2175 1496 2179
rect 1552 2175 1556 2179
rect 1976 2187 1980 2191
rect 784 2171 788 2175
rect 852 2171 856 2175
rect 1652 2171 1656 2175
rect 524 2157 528 2161
rect 620 2159 624 2163
rect 732 2159 736 2163
rect 860 2159 864 2163
rect 996 2159 1000 2163
rect 1072 2159 1076 2163
rect 1132 2159 1136 2163
rect 1216 2159 1220 2163
rect 1276 2159 1280 2163
rect 784 2127 788 2131
rect 792 2151 796 2155
rect 792 2127 796 2131
rect 1420 2157 1424 2161
rect 1480 2159 1484 2163
rect 1556 2159 1560 2163
rect 1692 2159 1696 2163
rect 1836 2159 1840 2163
rect 1956 2159 1960 2163
rect 1976 2159 1980 2163
rect 1216 2127 1220 2131
rect 1480 2127 1484 2131
rect 2744 2095 2748 2099
rect 2332 2063 2336 2067
rect 2444 2063 2448 2067
rect 2684 2063 2688 2067
rect 2744 2063 2748 2067
rect 2812 2063 2816 2067
rect 3092 2063 3096 2067
rect 3244 2063 3248 2067
rect 3404 2063 3408 2067
rect 3572 2063 3576 2067
rect 3892 2063 3896 2067
rect 2564 2059 2568 2063
rect 2948 2059 2952 2063
rect 3740 2059 3744 2063
rect 1072 2055 1076 2059
rect 1504 2051 1508 2055
rect 2380 2037 2384 2041
rect 2484 2039 2488 2043
rect 2588 2039 2592 2043
rect 2700 2039 2704 2043
rect 2828 2039 2832 2043
rect 2972 2039 2976 2043
rect 3132 2039 3136 2043
rect 3316 2039 3320 2043
rect 3508 2039 3512 2043
rect 3708 2039 3712 2043
rect 3892 2039 3896 2043
rect 788 2023 792 2027
rect 908 2023 912 2027
rect 1036 2023 1040 2027
rect 1172 2023 1176 2027
rect 1308 2023 1312 2027
rect 1504 2023 1508 2027
rect 1580 2023 1584 2027
rect 1708 2023 1712 2027
rect 1844 2023 1848 2027
rect 1956 2023 1960 2027
rect 676 2019 680 2023
rect 1444 2019 1448 2023
rect 500 2003 504 2007
rect 628 2003 632 2007
rect 780 2003 784 2007
rect 940 2003 944 2007
rect 1108 2003 1112 2007
rect 1284 2003 1288 2007
rect 1452 2003 1456 2007
rect 1628 2003 1632 2007
rect 1804 2003 1808 2007
rect 1956 2003 1960 2007
rect 648 1899 652 1903
rect 840 1899 844 1903
rect 1032 1899 1036 1903
rect 2404 1899 2408 1903
rect 2500 1899 2504 1903
rect 2596 1899 2600 1903
rect 2700 1899 2704 1903
rect 2820 1899 2824 1903
rect 2972 1899 2976 1903
rect 3156 1899 3160 1903
rect 3372 1899 3376 1903
rect 3828 1899 3832 1903
rect 2308 1895 2312 1899
rect 3596 1895 3600 1899
rect 3624 1895 3628 1899
rect 2236 1871 2240 1875
rect 2272 1871 2276 1875
rect 2332 1871 2336 1875
rect 2376 1871 2380 1875
rect 2436 1871 2440 1875
rect 2540 1871 2544 1875
rect 2644 1871 2648 1875
rect 2756 1871 2760 1875
rect 2884 1871 2888 1875
rect 3044 1871 3048 1875
rect 3236 1871 3240 1875
rect 3452 1871 3456 1875
rect 708 1867 712 1871
rect 804 1867 808 1871
rect 840 1867 844 1871
rect 900 1867 904 1871
rect 996 1867 1000 1871
rect 1032 1867 1036 1871
rect 1092 1867 1096 1871
rect 1188 1867 1192 1871
rect 1380 1867 1384 1871
rect 1476 1867 1480 1871
rect 1284 1863 1288 1867
rect 372 1851 376 1855
rect 500 1851 504 1855
rect 636 1851 640 1855
rect 648 1851 652 1855
rect 696 1851 700 1855
rect 772 1851 776 1855
rect 908 1851 912 1855
rect 1044 1849 1048 1853
rect 1180 1851 1184 1855
rect 1316 1851 1320 1855
rect 1452 1851 1456 1855
rect 1588 1851 1592 1855
rect 2272 1839 2276 1843
rect 2376 1839 2380 1843
rect 3684 1871 3688 1875
rect 3892 1871 3896 1875
rect 3624 1839 3628 1843
rect 696 1819 700 1823
rect 2216 1763 2220 1767
rect 2400 1763 2404 1767
rect 2968 1763 2972 1767
rect 2180 1731 2184 1735
rect 2216 1731 2220 1735
rect 2364 1731 2368 1735
rect 2400 1731 2404 1735
rect 2740 1731 2744 1735
rect 2932 1731 2936 1735
rect 2968 1731 2972 1735
rect 3124 1731 3128 1735
rect 3316 1731 3320 1735
rect 3716 1731 3720 1735
rect 2548 1727 2552 1731
rect 3516 1727 3520 1731
rect 3892 1727 3896 1731
rect 308 1711 312 1715
rect 588 1711 592 1715
rect 748 1711 752 1715
rect 916 1711 920 1715
rect 1260 1711 1264 1715
rect 1436 1711 1440 1715
rect 1612 1711 1616 1715
rect 1796 1711 1800 1715
rect 444 1707 448 1711
rect 1084 1707 1088 1711
rect 2124 1709 2128 1713
rect 2244 1711 2248 1715
rect 2396 1711 2400 1715
rect 2564 1711 2568 1715
rect 2740 1711 2744 1715
rect 2924 1711 2928 1715
rect 3116 1711 3120 1715
rect 3308 1711 3312 1715
rect 3500 1711 3504 1715
rect 3700 1711 3704 1715
rect 3892 1711 3896 1715
rect 188 1695 192 1699
rect 316 1695 320 1699
rect 484 1695 488 1699
rect 660 1695 664 1699
rect 852 1695 856 1699
rect 1052 1693 1056 1697
rect 1252 1695 1256 1699
rect 1460 1695 1464 1699
rect 1676 1695 1680 1699
rect 1892 1695 1896 1699
rect 2124 1575 2128 1579
rect 2388 1575 2392 1579
rect 2652 1575 2656 1579
rect 2892 1575 2896 1579
rect 3100 1575 3104 1579
rect 3284 1575 3288 1579
rect 3604 1575 3608 1579
rect 3748 1575 3752 1579
rect 3452 1571 3456 1575
rect 3892 1571 3896 1575
rect 188 1559 192 1563
rect 524 1559 528 1563
rect 708 1559 712 1563
rect 892 1559 896 1563
rect 1068 1559 1072 1563
rect 1236 1559 1240 1563
rect 1548 1559 1552 1563
rect 1692 1559 1696 1563
rect 1836 1559 1840 1563
rect 1956 1559 1960 1563
rect 340 1555 344 1559
rect 1396 1555 1400 1559
rect 2636 1555 2640 1559
rect 2796 1555 2800 1559
rect 2956 1555 2960 1559
rect 3116 1555 3120 1559
rect 3276 1553 3280 1557
rect 3436 1555 3440 1559
rect 3596 1555 3600 1559
rect 3756 1555 3760 1559
rect 188 1539 192 1543
rect 348 1539 352 1543
rect 540 1539 544 1543
rect 740 1539 744 1543
rect 940 1539 944 1543
rect 1132 1537 1136 1541
rect 1316 1539 1320 1543
rect 1500 1539 1504 1543
rect 1676 1539 1680 1543
rect 1860 1539 1864 1543
rect 656 1435 660 1439
rect 1096 1435 1100 1439
rect 228 1403 232 1407
rect 620 1403 624 1407
rect 656 1403 660 1407
rect 836 1403 840 1407
rect 412 1399 416 1403
rect 1060 1399 1064 1403
rect 380 1387 384 1391
rect 516 1387 520 1391
rect 652 1387 656 1391
rect 780 1387 784 1391
rect 908 1387 912 1391
rect 1036 1385 1040 1389
rect 2564 1419 2568 1423
rect 2660 1419 2664 1423
rect 2756 1419 2760 1423
rect 2852 1419 2856 1423
rect 2972 1419 2976 1423
rect 3116 1419 3120 1423
rect 3284 1419 3288 1423
rect 3468 1419 3472 1423
rect 3668 1419 3672 1423
rect 2468 1415 2472 1419
rect 3868 1415 3872 1419
rect 1284 1403 1288 1407
rect 1748 1403 1752 1407
rect 1956 1403 1960 1407
rect 1516 1399 1520 1403
rect 1172 1387 1176 1391
rect 1316 1387 1320 1391
rect 1476 1387 1480 1391
rect 1636 1385 1640 1389
rect 1804 1387 1808 1391
rect 1956 1387 1960 1391
rect 2124 1383 2128 1387
rect 2356 1383 2360 1387
rect 2612 1383 2616 1387
rect 2860 1383 2864 1387
rect 3108 1383 3112 1387
rect 3356 1383 3360 1387
rect 3612 1383 3616 1387
rect 3868 1383 3872 1387
rect 1096 1379 1100 1383
rect 3504 1351 3508 1355
rect 3504 1295 3508 1299
rect 708 1243 712 1247
rect 820 1243 824 1247
rect 932 1243 936 1247
rect 1044 1243 1048 1247
rect 1156 1243 1160 1247
rect 1380 1243 1384 1247
rect 1492 1243 1496 1247
rect 1612 1243 1616 1247
rect 604 1239 608 1243
rect 1268 1239 1272 1243
rect 2124 1239 2128 1243
rect 2276 1239 2280 1243
rect 2468 1239 2472 1243
rect 2868 1239 2872 1243
rect 3052 1239 3056 1243
rect 3228 1239 3232 1243
rect 3396 1239 3400 1243
rect 3556 1239 3560 1243
rect 3716 1239 3720 1243
rect 2668 1235 2672 1239
rect 3884 1235 3888 1239
rect 444 1225 448 1229
rect 572 1227 576 1231
rect 716 1227 720 1231
rect 860 1227 864 1231
rect 928 1227 932 1231
rect 1012 1227 1016 1231
rect 1164 1227 1168 1231
rect 1308 1227 1312 1231
rect 1460 1227 1464 1231
rect 1528 1227 1532 1231
rect 1612 1227 1616 1231
rect 1764 1227 1768 1231
rect 928 1195 932 1199
rect 2188 1213 2192 1217
rect 2364 1215 2368 1219
rect 2556 1215 2560 1219
rect 2748 1215 2752 1219
rect 2792 1215 2796 1219
rect 2940 1215 2944 1219
rect 1528 1195 1532 1199
rect 3124 1213 3128 1217
rect 3292 1215 3296 1219
rect 3452 1215 3456 1219
rect 3604 1215 3608 1219
rect 3640 1215 3644 1219
rect 3756 1215 3760 1219
rect 3892 1215 3896 1219
rect 2792 1183 2796 1187
rect 3640 1183 3644 1187
rect 1704 1115 1708 1119
rect 380 1087 384 1091
rect 548 1087 552 1091
rect 724 1087 728 1091
rect 900 1087 904 1091
rect 1084 1087 1088 1091
rect 1260 1087 1264 1091
rect 1620 1087 1624 1091
rect 1704 1087 1708 1091
rect 1804 1087 1808 1091
rect 228 1083 232 1087
rect 1436 1083 1440 1087
rect 1456 1083 1460 1087
rect 188 1063 192 1067
rect 284 1063 288 1067
rect 428 1063 432 1067
rect 596 1063 600 1067
rect 780 1063 784 1067
rect 964 1063 968 1067
rect 1148 1063 1152 1067
rect 1332 1063 1336 1067
rect 2476 1071 2480 1075
rect 2612 1071 2616 1075
rect 2748 1071 2752 1075
rect 2892 1071 2896 1075
rect 3044 1071 3048 1075
rect 3204 1071 3208 1075
rect 3372 1071 3376 1075
rect 3548 1071 3552 1075
rect 3732 1071 3736 1075
rect 2348 1067 2352 1071
rect 2424 1067 2428 1071
rect 3892 1067 3896 1071
rect 1516 1063 1520 1067
rect 1700 1063 1704 1067
rect 1884 1063 1888 1067
rect 1456 1031 1460 1035
rect 2548 1051 2552 1055
rect 2652 1051 2656 1055
rect 2764 1051 2768 1055
rect 2800 1051 2804 1055
rect 2900 1051 2904 1055
rect 3060 1051 3064 1055
rect 3252 1051 3256 1055
rect 3460 1051 3464 1055
rect 3684 1051 3688 1055
rect 3892 1051 3896 1055
rect 2424 1019 2428 1023
rect 2800 1019 2804 1023
rect 408 959 412 963
rect 188 927 192 931
rect 324 927 328 931
rect 408 927 412 931
rect 500 927 504 931
rect 684 927 688 931
rect 1060 927 1064 931
rect 1388 927 1392 931
rect 1540 927 1544 931
rect 1684 927 1688 931
rect 1828 927 1832 931
rect 1956 927 1960 931
rect 876 923 880 927
rect 1228 923 1232 927
rect 188 911 192 915
rect 324 911 328 915
rect 508 911 512 915
rect 708 911 712 915
rect 908 911 912 915
rect 1108 911 1112 915
rect 1292 911 1296 915
rect 1468 911 1472 915
rect 1636 911 1640 915
rect 1804 913 1808 917
rect 2796 915 2800 919
rect 2900 915 2904 919
rect 3020 915 3024 919
rect 3164 915 3168 919
rect 3332 915 3336 919
rect 3516 915 3520 919
rect 3716 915 3720 919
rect 1956 911 1960 915
rect 2700 911 2704 915
rect 3892 911 3896 915
rect 2124 885 2128 889
rect 2308 887 2312 891
rect 2516 887 2520 891
rect 2732 887 2736 891
rect 2784 887 2788 891
rect 3180 889 3184 893
rect 2948 885 2952 889
rect 3420 887 3424 891
rect 3668 887 3672 891
rect 3892 887 3896 891
rect 2784 855 2788 859
rect 432 807 436 811
rect 792 807 796 811
rect 3024 783 3028 787
rect 268 775 272 779
rect 396 775 400 779
rect 432 775 436 779
rect 548 775 552 779
rect 708 775 712 779
rect 792 775 796 779
rect 1060 775 1064 779
rect 1236 775 1240 779
rect 1412 775 1416 779
rect 1588 775 1592 779
rect 884 771 888 775
rect 1772 771 1776 775
rect 428 757 432 761
rect 548 759 552 763
rect 676 759 680 763
rect 804 759 808 763
rect 940 757 944 761
rect 1076 759 1080 763
rect 1220 759 1224 763
rect 1364 759 1368 763
rect 1508 759 1512 763
rect 1592 759 1596 763
rect 1652 759 1656 763
rect 2268 751 2272 755
rect 2380 751 2384 755
rect 2500 751 2504 755
rect 2636 751 2640 755
rect 2788 751 2792 755
rect 2948 751 2952 755
rect 3024 751 3028 755
rect 3300 751 3304 755
rect 3500 751 3504 755
rect 3708 751 3712 755
rect 3116 747 3120 751
rect 3892 747 3896 751
rect 1592 727 1596 731
rect 2428 729 2432 733
rect 2548 731 2552 735
rect 2676 729 2680 733
rect 2820 731 2824 735
rect 2964 731 2968 735
rect 3116 731 3120 735
rect 3268 731 3272 735
rect 3336 731 3340 735
rect 3420 731 3424 735
rect 3488 731 3492 735
rect 3572 731 3576 735
rect 3732 731 3736 735
rect 3892 731 3896 735
rect 3336 699 3340 703
rect 3488 699 3492 703
rect 960 655 964 659
rect 1160 655 1164 659
rect 580 623 584 627
rect 684 623 688 627
rect 796 623 800 627
rect 908 623 912 627
rect 960 623 964 627
rect 1124 623 1128 627
rect 1160 623 1164 627
rect 1236 623 1240 627
rect 1348 623 1352 627
rect 1460 623 1464 627
rect 968 619 972 623
rect 1020 619 1024 623
rect 1572 619 1576 623
rect 2104 619 2108 623
rect 740 605 744 609
rect 836 607 840 611
rect 872 607 876 611
rect 932 607 936 611
rect 872 575 876 579
rect 1028 607 1032 611
rect 1124 605 1128 609
rect 1220 607 1224 611
rect 1316 607 1320 611
rect 1412 607 1416 611
rect 1508 607 1512 611
rect 968 575 972 579
rect 2360 619 2364 623
rect 2164 587 2168 591
rect 2300 587 2304 591
rect 2360 587 2364 591
rect 2452 587 2456 591
rect 2628 587 2632 591
rect 2812 587 2816 591
rect 3180 587 3184 591
rect 3356 587 3360 591
rect 3532 587 3536 591
rect 3708 587 3712 591
rect 2996 583 3000 587
rect 3884 583 3888 587
rect 2104 567 2108 571
rect 2124 567 2128 571
rect 2236 567 2240 571
rect 2388 567 2392 571
rect 2556 567 2560 571
rect 2640 567 2644 571
rect 2740 567 2744 571
rect 2932 567 2936 571
rect 3124 567 3128 571
rect 3316 567 3320 571
rect 3508 567 3512 571
rect 3700 567 3704 571
rect 3892 567 3896 571
rect 2640 535 2644 539
rect 1240 483 1244 487
rect 532 451 536 455
rect 628 451 632 455
rect 724 451 728 455
rect 820 451 824 455
rect 916 451 920 455
rect 1012 451 1016 455
rect 1108 451 1112 455
rect 1204 451 1208 455
rect 436 447 440 451
rect 1528 483 1532 487
rect 1528 459 1532 463
rect 3456 463 3460 467
rect 1300 451 1304 455
rect 1396 451 1400 455
rect 1588 451 1592 455
rect 1492 447 1496 451
rect 2236 431 2240 435
rect 2372 431 2376 435
rect 2516 431 2520 435
rect 2668 431 2672 435
rect 2828 431 2832 435
rect 3012 431 3016 435
rect 3212 431 3216 435
rect 3420 431 3424 435
rect 3456 431 3460 435
rect 3636 427 3640 431
rect 3860 427 3864 431
rect 540 421 544 425
rect 636 423 640 427
rect 740 423 744 427
rect 784 423 788 427
rect 844 423 848 427
rect 888 423 892 427
rect 948 423 952 427
rect 1052 423 1056 427
rect 1096 423 1100 427
rect 1156 423 1160 427
rect 1240 423 1244 427
rect 1260 423 1264 427
rect 1372 423 1376 427
rect 784 391 788 395
rect 888 391 892 395
rect 1484 421 1488 425
rect 2396 417 2400 421
rect 2540 415 2544 419
rect 2692 415 2696 419
rect 2852 415 2856 419
rect 3012 415 3016 419
rect 3164 413 3168 417
rect 3316 415 3320 419
rect 3468 415 3472 419
rect 3612 415 3616 419
rect 3764 415 3768 419
rect 3892 415 3896 419
rect 1096 391 1100 395
rect 516 283 520 287
rect 668 283 672 287
rect 820 283 824 287
rect 972 283 976 287
rect 1116 283 1120 287
rect 1260 283 1264 287
rect 1404 283 1408 287
rect 1548 283 1552 287
rect 380 279 384 283
rect 1692 279 1696 283
rect 832 275 836 279
rect 2548 275 2552 279
rect 2692 275 2696 279
rect 2852 275 2856 279
rect 3012 275 3016 279
rect 3172 275 3176 279
rect 3476 275 3480 279
rect 3620 275 3624 279
rect 3764 275 3768 279
rect 220 257 224 261
rect 380 259 384 263
rect 556 259 560 263
rect 740 259 744 263
rect 824 259 828 263
rect 824 227 828 231
rect 3324 271 3328 275
rect 3892 271 3896 275
rect 924 259 928 263
rect 1100 257 1104 261
rect 1268 259 1272 263
rect 1420 259 1424 263
rect 1564 259 1568 263
rect 1700 259 1704 263
rect 1836 259 1840 263
rect 1956 259 1960 263
rect 2124 259 2128 263
rect 2324 259 2328 263
rect 2548 259 2552 263
rect 2756 259 2760 263
rect 2800 259 2804 263
rect 2956 259 2960 263
rect 832 227 836 231
rect 3148 257 3152 261
rect 3340 259 3344 263
rect 3532 259 3536 263
rect 3724 259 3728 263
rect 3892 259 3896 263
rect 2800 227 2804 231
rect 2124 99 2128 103
rect 2220 99 2224 103
rect 2316 99 2320 103
rect 2412 99 2416 103
rect 2508 99 2512 103
rect 2604 99 2608 103
rect 2708 99 2712 103
rect 2812 99 2816 103
rect 2916 99 2920 103
rect 3028 99 3032 103
rect 3156 99 3160 103
rect 3292 99 3296 103
rect 3436 99 3440 103
rect 3588 99 3592 103
rect 3748 99 3752 103
rect 3892 99 3896 103
rect 284 95 288 99
rect 380 95 384 99
rect 476 95 480 99
rect 580 95 584 99
rect 700 95 704 99
rect 828 95 832 99
rect 956 95 960 99
rect 1084 95 1088 99
rect 1204 95 1208 99
rect 1324 95 1328 99
rect 1436 95 1440 99
rect 1540 95 1544 99
rect 1644 95 1648 99
rect 1756 95 1760 99
rect 1860 95 1864 99
rect 1956 95 1960 99
<< m2 >>
rect 2146 4011 2152 4012
rect 2123 4009 2129 4010
rect 2123 4005 2124 4009
rect 2128 4005 2129 4009
rect 2146 4007 2147 4011
rect 2151 4010 2152 4011
rect 2219 4011 2225 4012
rect 2219 4010 2220 4011
rect 2151 4008 2220 4010
rect 2151 4007 2152 4008
rect 2146 4006 2152 4007
rect 2219 4007 2220 4008
rect 2224 4007 2225 4011
rect 2219 4006 2225 4007
rect 2242 4011 2248 4012
rect 2242 4007 2243 4011
rect 2247 4010 2248 4011
rect 2315 4011 2321 4012
rect 2315 4010 2316 4011
rect 2247 4008 2316 4010
rect 2247 4007 2248 4008
rect 2242 4006 2248 4007
rect 2315 4007 2316 4008
rect 2320 4007 2321 4011
rect 2315 4006 2321 4007
rect 110 4004 116 4005
rect 2006 4004 2012 4005
rect 2123 4004 2129 4005
rect 110 4000 111 4004
rect 115 4000 116 4004
rect 110 3999 116 4000
rect 1518 4003 1524 4004
rect 1518 3999 1519 4003
rect 1523 3999 1524 4003
rect 1518 3998 1524 3999
rect 1614 4003 1620 4004
rect 1614 3999 1615 4003
rect 1619 3999 1620 4003
rect 1614 3998 1620 3999
rect 1710 4003 1716 4004
rect 1710 3999 1711 4003
rect 1715 3999 1716 4003
rect 1710 3998 1716 3999
rect 1806 4003 1812 4004
rect 1806 3999 1807 4003
rect 1811 3999 1812 4003
rect 1806 3998 1812 3999
rect 1902 4003 1908 4004
rect 1902 3999 1903 4003
rect 1907 3999 1908 4003
rect 2006 4000 2007 4004
rect 2011 4000 2012 4004
rect 2006 3999 2012 4000
rect 1902 3998 1908 3999
rect 1607 3995 1613 3996
rect 1607 3994 1608 3995
rect 1597 3992 1608 3994
rect 1607 3991 1608 3992
rect 1612 3991 1613 3995
rect 2124 3994 2126 4004
rect 1981 3992 2126 3994
rect 1607 3990 1613 3991
rect 1690 3991 1696 3992
rect 110 3987 116 3988
rect 110 3983 111 3987
rect 115 3983 116 3987
rect 1690 3987 1691 3991
rect 1695 3987 1696 3991
rect 1690 3986 1696 3987
rect 1786 3991 1792 3992
rect 1786 3987 1787 3991
rect 1791 3987 1792 3991
rect 1786 3986 1792 3987
rect 1882 3991 1888 3992
rect 1882 3987 1883 3991
rect 1887 3987 1888 3991
rect 2070 3988 2076 3989
rect 1882 3986 1888 3987
rect 2006 3987 2012 3988
rect 110 3982 116 3983
rect 1518 3984 1524 3985
rect 1518 3980 1519 3984
rect 1523 3980 1524 3984
rect 1518 3979 1524 3980
rect 1614 3984 1620 3985
rect 1614 3980 1615 3984
rect 1619 3980 1620 3984
rect 1614 3979 1620 3980
rect 1710 3984 1716 3985
rect 1710 3980 1711 3984
rect 1715 3980 1716 3984
rect 1710 3979 1716 3980
rect 1806 3984 1812 3985
rect 1806 3980 1807 3984
rect 1811 3980 1812 3984
rect 1806 3979 1812 3980
rect 1902 3984 1908 3985
rect 1902 3980 1903 3984
rect 1907 3980 1908 3984
rect 2006 3983 2007 3987
rect 2011 3983 2012 3987
rect 2006 3982 2012 3983
rect 2046 3985 2052 3986
rect 2046 3981 2047 3985
rect 2051 3981 2052 3985
rect 2070 3984 2071 3988
rect 2075 3984 2076 3988
rect 2070 3983 2076 3984
rect 2166 3988 2172 3989
rect 2166 3984 2167 3988
rect 2171 3984 2172 3988
rect 2166 3983 2172 3984
rect 2262 3988 2268 3989
rect 2262 3984 2263 3988
rect 2267 3984 2268 3988
rect 2262 3983 2268 3984
rect 3942 3985 3948 3986
rect 2046 3980 2052 3981
rect 3942 3981 3943 3985
rect 3947 3981 3948 3985
rect 3942 3980 3948 3981
rect 1902 3979 1908 3980
rect 2146 3979 2152 3980
rect 2146 3975 2147 3979
rect 2151 3975 2152 3979
rect 2146 3974 2152 3975
rect 2242 3979 2248 3980
rect 2242 3975 2243 3979
rect 2247 3975 2248 3979
rect 2242 3974 2248 3975
rect 2255 3979 2261 3980
rect 2255 3975 2256 3979
rect 2260 3978 2261 3979
rect 2260 3976 2305 3978
rect 2260 3975 2261 3976
rect 2255 3974 2261 3975
rect 2070 3969 2076 3970
rect 2046 3968 2052 3969
rect 2046 3964 2047 3968
rect 2051 3964 2052 3968
rect 2070 3965 2071 3969
rect 2075 3965 2076 3969
rect 2070 3964 2076 3965
rect 2166 3969 2172 3970
rect 2166 3965 2167 3969
rect 2171 3965 2172 3969
rect 2166 3964 2172 3965
rect 2262 3969 2268 3970
rect 2262 3965 2263 3969
rect 2267 3965 2268 3969
rect 2262 3964 2268 3965
rect 3942 3968 3948 3969
rect 3942 3964 3943 3968
rect 3947 3964 3948 3968
rect 1607 3963 1613 3964
rect 1571 3959 1577 3960
rect 1571 3955 1572 3959
rect 1576 3958 1577 3959
rect 1599 3959 1605 3960
rect 1599 3958 1600 3959
rect 1576 3956 1600 3958
rect 1576 3955 1577 3956
rect 1571 3954 1577 3955
rect 1599 3955 1600 3956
rect 1604 3955 1605 3959
rect 1607 3959 1608 3963
rect 1612 3962 1613 3963
rect 1667 3963 1673 3964
rect 1667 3962 1668 3963
rect 1612 3960 1668 3962
rect 1612 3959 1613 3960
rect 1607 3958 1613 3959
rect 1667 3959 1668 3960
rect 1672 3959 1673 3963
rect 1667 3958 1673 3959
rect 1690 3963 1696 3964
rect 1690 3959 1691 3963
rect 1695 3962 1696 3963
rect 1763 3963 1769 3964
rect 1763 3962 1764 3963
rect 1695 3960 1764 3962
rect 1695 3959 1696 3960
rect 1690 3958 1696 3959
rect 1763 3959 1764 3960
rect 1768 3959 1769 3963
rect 1763 3958 1769 3959
rect 1786 3963 1792 3964
rect 1786 3959 1787 3963
rect 1791 3962 1792 3963
rect 1859 3963 1865 3964
rect 1859 3962 1860 3963
rect 1791 3960 1860 3962
rect 1791 3959 1792 3960
rect 1786 3958 1792 3959
rect 1859 3959 1860 3960
rect 1864 3959 1865 3963
rect 1859 3958 1865 3959
rect 1882 3963 1888 3964
rect 1882 3959 1883 3963
rect 1887 3962 1888 3963
rect 1955 3963 1961 3964
rect 2046 3963 2052 3964
rect 3942 3963 3948 3964
rect 1955 3962 1956 3963
rect 1887 3960 1956 3962
rect 1887 3959 1888 3960
rect 1882 3958 1888 3959
rect 1955 3959 1956 3960
rect 1960 3959 1961 3963
rect 1955 3958 1961 3959
rect 1599 3954 1605 3955
rect 251 3947 257 3948
rect 251 3943 252 3947
rect 256 3946 257 3947
rect 266 3947 272 3948
rect 266 3946 267 3947
rect 256 3944 267 3946
rect 256 3943 257 3944
rect 251 3942 257 3943
rect 266 3943 267 3944
rect 271 3943 272 3947
rect 266 3942 272 3943
rect 274 3947 280 3948
rect 274 3943 275 3947
rect 279 3946 280 3947
rect 347 3947 353 3948
rect 347 3946 348 3947
rect 279 3944 348 3946
rect 279 3943 280 3944
rect 274 3942 280 3943
rect 347 3943 348 3944
rect 352 3943 353 3947
rect 347 3942 353 3943
rect 370 3947 376 3948
rect 370 3943 371 3947
rect 375 3946 376 3947
rect 443 3947 449 3948
rect 443 3946 444 3947
rect 375 3944 444 3946
rect 375 3943 376 3944
rect 370 3942 376 3943
rect 443 3943 444 3944
rect 448 3943 449 3947
rect 443 3942 449 3943
rect 466 3947 472 3948
rect 466 3943 467 3947
rect 471 3946 472 3947
rect 547 3947 553 3948
rect 547 3946 548 3947
rect 471 3944 548 3946
rect 471 3943 472 3944
rect 466 3942 472 3943
rect 547 3943 548 3944
rect 552 3943 553 3947
rect 547 3942 553 3943
rect 570 3947 576 3948
rect 570 3943 571 3947
rect 575 3946 576 3947
rect 667 3947 673 3948
rect 667 3946 668 3947
rect 575 3944 668 3946
rect 575 3943 576 3944
rect 570 3942 576 3943
rect 667 3943 668 3944
rect 672 3943 673 3947
rect 667 3942 673 3943
rect 690 3947 696 3948
rect 690 3943 691 3947
rect 695 3946 696 3947
rect 795 3947 801 3948
rect 795 3946 796 3947
rect 695 3944 796 3946
rect 695 3943 696 3944
rect 690 3942 696 3943
rect 795 3943 796 3944
rect 800 3943 801 3947
rect 795 3942 801 3943
rect 818 3947 824 3948
rect 818 3943 819 3947
rect 823 3946 824 3947
rect 923 3947 929 3948
rect 923 3946 924 3947
rect 823 3944 924 3946
rect 823 3943 824 3944
rect 818 3942 824 3943
rect 923 3943 924 3944
rect 928 3943 929 3947
rect 923 3942 929 3943
rect 946 3947 952 3948
rect 946 3943 947 3947
rect 951 3946 952 3947
rect 1051 3947 1057 3948
rect 1051 3946 1052 3947
rect 951 3944 1052 3946
rect 951 3943 952 3944
rect 946 3942 952 3943
rect 1051 3943 1052 3944
rect 1056 3943 1057 3947
rect 1051 3942 1057 3943
rect 1178 3947 1185 3948
rect 1178 3943 1179 3947
rect 1184 3943 1185 3947
rect 1178 3942 1185 3943
rect 1202 3947 1208 3948
rect 1202 3943 1203 3947
rect 1207 3946 1208 3947
rect 1307 3947 1313 3948
rect 1307 3946 1308 3947
rect 1207 3944 1308 3946
rect 1207 3943 1208 3944
rect 1202 3942 1208 3943
rect 1307 3943 1308 3944
rect 1312 3943 1313 3947
rect 1307 3942 1313 3943
rect 1330 3947 1336 3948
rect 1330 3943 1331 3947
rect 1335 3946 1336 3947
rect 1435 3947 1441 3948
rect 1435 3946 1436 3947
rect 1335 3944 1436 3946
rect 1335 3943 1336 3944
rect 1330 3942 1336 3943
rect 1435 3943 1436 3944
rect 1440 3943 1441 3947
rect 1435 3942 1441 3943
rect 1458 3947 1464 3948
rect 1458 3943 1459 3947
rect 1463 3946 1464 3947
rect 1563 3947 1569 3948
rect 1563 3946 1564 3947
rect 1463 3944 1564 3946
rect 1463 3943 1464 3944
rect 1458 3942 1464 3943
rect 1563 3943 1564 3944
rect 1568 3943 1569 3947
rect 1563 3942 1569 3943
rect 1586 3947 1592 3948
rect 1586 3943 1587 3947
rect 1591 3946 1592 3947
rect 1699 3947 1705 3948
rect 1699 3946 1700 3947
rect 1591 3944 1700 3946
rect 1591 3943 1592 3944
rect 1586 3942 1592 3943
rect 1699 3943 1700 3944
rect 1704 3943 1705 3947
rect 1699 3942 1705 3943
rect 198 3924 204 3925
rect 110 3921 116 3922
rect 110 3917 111 3921
rect 115 3917 116 3921
rect 198 3920 199 3924
rect 203 3920 204 3924
rect 198 3919 204 3920
rect 294 3924 300 3925
rect 294 3920 295 3924
rect 299 3920 300 3924
rect 294 3919 300 3920
rect 390 3924 396 3925
rect 390 3920 391 3924
rect 395 3920 396 3924
rect 390 3919 396 3920
rect 494 3924 500 3925
rect 494 3920 495 3924
rect 499 3920 500 3924
rect 494 3919 500 3920
rect 614 3924 620 3925
rect 614 3920 615 3924
rect 619 3920 620 3924
rect 614 3919 620 3920
rect 742 3924 748 3925
rect 742 3920 743 3924
rect 747 3920 748 3924
rect 742 3919 748 3920
rect 870 3924 876 3925
rect 870 3920 871 3924
rect 875 3920 876 3924
rect 870 3919 876 3920
rect 998 3924 1004 3925
rect 998 3920 999 3924
rect 1003 3920 1004 3924
rect 998 3919 1004 3920
rect 1126 3924 1132 3925
rect 1126 3920 1127 3924
rect 1131 3920 1132 3924
rect 1126 3919 1132 3920
rect 1254 3924 1260 3925
rect 1254 3920 1255 3924
rect 1259 3920 1260 3924
rect 1254 3919 1260 3920
rect 1382 3924 1388 3925
rect 1382 3920 1383 3924
rect 1387 3920 1388 3924
rect 1382 3919 1388 3920
rect 1510 3924 1516 3925
rect 1510 3920 1511 3924
rect 1515 3920 1516 3924
rect 1510 3919 1516 3920
rect 1646 3924 1652 3925
rect 1646 3920 1647 3924
rect 1651 3920 1652 3924
rect 1646 3919 1652 3920
rect 2006 3921 2012 3922
rect 110 3916 116 3917
rect 2006 3917 2007 3921
rect 2011 3917 2012 3921
rect 2006 3916 2012 3917
rect 2046 3916 2052 3917
rect 3942 3916 3948 3917
rect 274 3915 280 3916
rect 274 3911 275 3915
rect 279 3911 280 3915
rect 274 3910 280 3911
rect 370 3915 376 3916
rect 370 3911 371 3915
rect 375 3911 376 3915
rect 370 3910 376 3911
rect 466 3915 472 3916
rect 466 3911 467 3915
rect 471 3911 472 3915
rect 466 3910 472 3911
rect 570 3915 576 3916
rect 570 3911 571 3915
rect 575 3911 576 3915
rect 570 3910 576 3911
rect 690 3915 696 3916
rect 690 3911 691 3915
rect 695 3911 696 3915
rect 690 3910 696 3911
rect 818 3915 824 3916
rect 818 3911 819 3915
rect 823 3911 824 3915
rect 818 3910 824 3911
rect 946 3915 952 3916
rect 946 3911 947 3915
rect 951 3911 952 3915
rect 946 3910 952 3911
rect 954 3915 960 3916
rect 954 3911 955 3915
rect 959 3914 960 3915
rect 1202 3915 1208 3916
rect 959 3912 1041 3914
rect 959 3911 960 3912
rect 954 3910 960 3911
rect 1202 3911 1203 3915
rect 1207 3911 1208 3915
rect 1202 3910 1208 3911
rect 1330 3915 1336 3916
rect 1330 3911 1331 3915
rect 1335 3911 1336 3915
rect 1330 3910 1336 3911
rect 1458 3915 1464 3916
rect 1458 3911 1459 3915
rect 1463 3911 1464 3915
rect 1458 3910 1464 3911
rect 1586 3915 1592 3916
rect 1586 3911 1587 3915
rect 1591 3911 1592 3915
rect 1586 3910 1592 3911
rect 1599 3915 1605 3916
rect 1599 3911 1600 3915
rect 1604 3914 1605 3915
rect 1604 3912 1689 3914
rect 2046 3912 2047 3916
rect 2051 3912 2052 3916
rect 1604 3911 1605 3912
rect 2046 3911 2052 3912
rect 2158 3915 2164 3916
rect 2158 3911 2159 3915
rect 2163 3911 2164 3915
rect 1599 3910 1605 3911
rect 2158 3910 2164 3911
rect 2286 3915 2292 3916
rect 2286 3911 2287 3915
rect 2291 3911 2292 3915
rect 2286 3910 2292 3911
rect 2414 3915 2420 3916
rect 2414 3911 2415 3915
rect 2419 3911 2420 3915
rect 2414 3910 2420 3911
rect 2550 3915 2556 3916
rect 2550 3911 2551 3915
rect 2555 3911 2556 3915
rect 2550 3910 2556 3911
rect 2686 3915 2692 3916
rect 2686 3911 2687 3915
rect 2691 3911 2692 3915
rect 2686 3910 2692 3911
rect 2822 3915 2828 3916
rect 2822 3911 2823 3915
rect 2827 3911 2828 3915
rect 2822 3910 2828 3911
rect 2950 3915 2956 3916
rect 2950 3911 2951 3915
rect 2955 3911 2956 3915
rect 2950 3910 2956 3911
rect 3070 3915 3076 3916
rect 3070 3911 3071 3915
rect 3075 3911 3076 3915
rect 3070 3910 3076 3911
rect 3190 3915 3196 3916
rect 3190 3911 3191 3915
rect 3195 3911 3196 3915
rect 3190 3910 3196 3911
rect 3302 3915 3308 3916
rect 3302 3911 3303 3915
rect 3307 3911 3308 3915
rect 3302 3910 3308 3911
rect 3406 3915 3412 3916
rect 3406 3911 3407 3915
rect 3411 3911 3412 3915
rect 3406 3910 3412 3911
rect 3518 3915 3524 3916
rect 3518 3911 3519 3915
rect 3523 3911 3524 3915
rect 3518 3910 3524 3911
rect 3630 3915 3636 3916
rect 3630 3911 3631 3915
rect 3635 3911 3636 3915
rect 3630 3910 3636 3911
rect 3742 3915 3748 3916
rect 3742 3911 3743 3915
rect 3747 3911 3748 3915
rect 3942 3912 3943 3916
rect 3947 3912 3948 3916
rect 3942 3911 3948 3912
rect 3742 3910 3748 3911
rect 3714 3907 3720 3908
rect 198 3905 204 3906
rect 110 3904 116 3905
rect 110 3900 111 3904
rect 115 3900 116 3904
rect 198 3901 199 3905
rect 203 3901 204 3905
rect 198 3900 204 3901
rect 294 3905 300 3906
rect 294 3901 295 3905
rect 299 3901 300 3905
rect 294 3900 300 3901
rect 390 3905 396 3906
rect 390 3901 391 3905
rect 395 3901 396 3905
rect 390 3900 396 3901
rect 494 3905 500 3906
rect 494 3901 495 3905
rect 499 3901 500 3905
rect 494 3900 500 3901
rect 614 3905 620 3906
rect 614 3901 615 3905
rect 619 3901 620 3905
rect 614 3900 620 3901
rect 742 3905 748 3906
rect 742 3901 743 3905
rect 747 3901 748 3905
rect 742 3900 748 3901
rect 870 3905 876 3906
rect 870 3901 871 3905
rect 875 3901 876 3905
rect 870 3900 876 3901
rect 998 3905 1004 3906
rect 998 3901 999 3905
rect 1003 3901 1004 3905
rect 998 3900 1004 3901
rect 1126 3905 1132 3906
rect 1126 3901 1127 3905
rect 1131 3901 1132 3905
rect 1126 3900 1132 3901
rect 1254 3905 1260 3906
rect 1254 3901 1255 3905
rect 1259 3901 1260 3905
rect 1254 3900 1260 3901
rect 1382 3905 1388 3906
rect 1382 3901 1383 3905
rect 1387 3901 1388 3905
rect 1382 3900 1388 3901
rect 1510 3905 1516 3906
rect 1510 3901 1511 3905
rect 1515 3901 1516 3905
rect 1510 3900 1516 3901
rect 1646 3905 1652 3906
rect 1646 3901 1647 3905
rect 1651 3901 1652 3905
rect 1646 3900 1652 3901
rect 2006 3904 2012 3905
rect 2006 3900 2007 3904
rect 2011 3900 2012 3904
rect 2270 3903 2276 3904
rect 2270 3902 2271 3903
rect 2237 3900 2271 3902
rect 110 3899 116 3900
rect 2006 3899 2012 3900
rect 2046 3899 2052 3900
rect 2046 3895 2047 3899
rect 2051 3895 2052 3899
rect 2270 3899 2271 3900
rect 2275 3899 2276 3903
rect 2270 3898 2276 3899
rect 2362 3903 2368 3904
rect 2362 3899 2363 3903
rect 2367 3899 2368 3903
rect 2362 3898 2368 3899
rect 2490 3903 2496 3904
rect 2490 3899 2491 3903
rect 2495 3899 2496 3903
rect 2490 3898 2496 3899
rect 2626 3903 2632 3904
rect 2626 3899 2627 3903
rect 2631 3899 2632 3903
rect 2782 3903 2788 3904
rect 2782 3902 2783 3903
rect 2765 3900 2783 3902
rect 2626 3898 2632 3899
rect 2782 3899 2783 3900
rect 2787 3899 2788 3903
rect 2782 3898 2788 3899
rect 2898 3903 2904 3904
rect 2898 3899 2899 3903
rect 2903 3899 2904 3903
rect 2898 3898 2904 3899
rect 3026 3903 3032 3904
rect 3026 3899 3027 3903
rect 3031 3899 3032 3903
rect 3026 3898 3032 3899
rect 3146 3903 3152 3904
rect 3146 3899 3147 3903
rect 3151 3899 3152 3903
rect 3146 3898 3152 3899
rect 3266 3903 3272 3904
rect 3266 3899 3267 3903
rect 3271 3899 3272 3903
rect 3266 3898 3272 3899
rect 3378 3903 3384 3904
rect 3378 3899 3379 3903
rect 3383 3899 3384 3903
rect 3378 3898 3384 3899
rect 3482 3903 3488 3904
rect 3482 3899 3483 3903
rect 3487 3899 3488 3903
rect 3482 3898 3488 3899
rect 3594 3903 3600 3904
rect 3594 3899 3595 3903
rect 3599 3899 3600 3903
rect 3594 3898 3600 3899
rect 3706 3903 3712 3904
rect 3706 3899 3707 3903
rect 3711 3899 3712 3903
rect 3714 3903 3715 3907
rect 3719 3906 3720 3907
rect 3719 3904 3785 3906
rect 3719 3903 3720 3904
rect 3714 3902 3720 3903
rect 3706 3898 3712 3899
rect 3942 3899 3948 3900
rect 2046 3894 2052 3895
rect 2158 3896 2164 3897
rect 2158 3892 2159 3896
rect 2163 3892 2164 3896
rect 2158 3891 2164 3892
rect 2286 3896 2292 3897
rect 2286 3892 2287 3896
rect 2291 3892 2292 3896
rect 2286 3891 2292 3892
rect 2414 3896 2420 3897
rect 2414 3892 2415 3896
rect 2419 3892 2420 3896
rect 2414 3891 2420 3892
rect 2550 3896 2556 3897
rect 2550 3892 2551 3896
rect 2555 3892 2556 3896
rect 2550 3891 2556 3892
rect 2686 3896 2692 3897
rect 2686 3892 2687 3896
rect 2691 3892 2692 3896
rect 2686 3891 2692 3892
rect 2822 3896 2828 3897
rect 2822 3892 2823 3896
rect 2827 3892 2828 3896
rect 2822 3891 2828 3892
rect 2950 3896 2956 3897
rect 2950 3892 2951 3896
rect 2955 3892 2956 3896
rect 2950 3891 2956 3892
rect 3070 3896 3076 3897
rect 3070 3892 3071 3896
rect 3075 3892 3076 3896
rect 3070 3891 3076 3892
rect 3190 3896 3196 3897
rect 3190 3892 3191 3896
rect 3195 3892 3196 3896
rect 3190 3891 3196 3892
rect 3302 3896 3308 3897
rect 3302 3892 3303 3896
rect 3307 3892 3308 3896
rect 3302 3891 3308 3892
rect 3406 3896 3412 3897
rect 3406 3892 3407 3896
rect 3411 3892 3412 3896
rect 3406 3891 3412 3892
rect 3518 3896 3524 3897
rect 3518 3892 3519 3896
rect 3523 3892 3524 3896
rect 3518 3891 3524 3892
rect 3630 3896 3636 3897
rect 3630 3892 3631 3896
rect 3635 3892 3636 3896
rect 3630 3891 3636 3892
rect 3742 3896 3748 3897
rect 3742 3892 3743 3896
rect 3747 3892 3748 3896
rect 3942 3895 3943 3899
rect 3947 3895 3948 3899
rect 3942 3894 3948 3895
rect 3742 3891 3748 3892
rect 2211 3875 2217 3876
rect 2211 3871 2212 3875
rect 2216 3874 2217 3875
rect 2255 3875 2261 3876
rect 2255 3874 2256 3875
rect 2216 3872 2256 3874
rect 2216 3871 2217 3872
rect 2211 3870 2217 3871
rect 2255 3871 2256 3872
rect 2260 3871 2261 3875
rect 2255 3870 2261 3871
rect 2270 3875 2276 3876
rect 2270 3871 2271 3875
rect 2275 3874 2276 3875
rect 2339 3875 2345 3876
rect 2339 3874 2340 3875
rect 2275 3872 2340 3874
rect 2275 3871 2276 3872
rect 2270 3870 2276 3871
rect 2339 3871 2340 3872
rect 2344 3871 2345 3875
rect 2339 3870 2345 3871
rect 2362 3875 2368 3876
rect 2362 3871 2363 3875
rect 2367 3874 2368 3875
rect 2467 3875 2473 3876
rect 2467 3874 2468 3875
rect 2367 3872 2468 3874
rect 2367 3871 2368 3872
rect 2362 3870 2368 3871
rect 2467 3871 2468 3872
rect 2472 3871 2473 3875
rect 2467 3870 2473 3871
rect 2490 3875 2496 3876
rect 2490 3871 2491 3875
rect 2495 3874 2496 3875
rect 2603 3875 2609 3876
rect 2603 3874 2604 3875
rect 2495 3872 2604 3874
rect 2495 3871 2496 3872
rect 2490 3870 2496 3871
rect 2603 3871 2604 3872
rect 2608 3871 2609 3875
rect 2603 3870 2609 3871
rect 2626 3875 2632 3876
rect 2626 3871 2627 3875
rect 2631 3874 2632 3875
rect 2739 3875 2745 3876
rect 2739 3874 2740 3875
rect 2631 3872 2740 3874
rect 2631 3871 2632 3872
rect 2626 3870 2632 3871
rect 2739 3871 2740 3872
rect 2744 3871 2745 3875
rect 2898 3875 2904 3876
rect 2739 3870 2745 3871
rect 2875 3871 2881 3872
rect 2875 3867 2876 3871
rect 2880 3870 2881 3871
rect 2898 3871 2899 3875
rect 2903 3874 2904 3875
rect 3003 3875 3009 3876
rect 3003 3874 3004 3875
rect 2903 3872 3004 3874
rect 2903 3871 2904 3872
rect 2898 3870 2904 3871
rect 3003 3871 3004 3872
rect 3008 3871 3009 3875
rect 3003 3870 3009 3871
rect 3026 3875 3032 3876
rect 3026 3871 3027 3875
rect 3031 3874 3032 3875
rect 3123 3875 3129 3876
rect 3123 3874 3124 3875
rect 3031 3872 3124 3874
rect 3031 3871 3032 3872
rect 3026 3870 3032 3871
rect 3123 3871 3124 3872
rect 3128 3871 3129 3875
rect 3123 3870 3129 3871
rect 3146 3875 3152 3876
rect 3146 3871 3147 3875
rect 3151 3874 3152 3875
rect 3243 3875 3249 3876
rect 3243 3874 3244 3875
rect 3151 3872 3244 3874
rect 3151 3871 3152 3872
rect 3146 3870 3152 3871
rect 3243 3871 3244 3872
rect 3248 3871 3249 3875
rect 3243 3870 3249 3871
rect 3266 3875 3272 3876
rect 3266 3871 3267 3875
rect 3271 3874 3272 3875
rect 3355 3875 3361 3876
rect 3355 3874 3356 3875
rect 3271 3872 3356 3874
rect 3271 3871 3272 3872
rect 3266 3870 3272 3871
rect 3355 3871 3356 3872
rect 3360 3871 3361 3875
rect 3355 3870 3361 3871
rect 3378 3875 3384 3876
rect 3378 3871 3379 3875
rect 3383 3874 3384 3875
rect 3459 3875 3465 3876
rect 3459 3874 3460 3875
rect 3383 3872 3460 3874
rect 3383 3871 3384 3872
rect 3378 3870 3384 3871
rect 3459 3871 3460 3872
rect 3464 3871 3465 3875
rect 3459 3870 3465 3871
rect 3482 3875 3488 3876
rect 3482 3871 3483 3875
rect 3487 3874 3488 3875
rect 3571 3875 3577 3876
rect 3571 3874 3572 3875
rect 3487 3872 3572 3874
rect 3487 3871 3488 3872
rect 3482 3870 3488 3871
rect 3571 3871 3572 3872
rect 3576 3871 3577 3875
rect 3571 3870 3577 3871
rect 3594 3875 3600 3876
rect 3594 3871 3595 3875
rect 3599 3874 3600 3875
rect 3683 3875 3689 3876
rect 3683 3874 3684 3875
rect 3599 3872 3684 3874
rect 3599 3871 3600 3872
rect 3594 3870 3600 3871
rect 3683 3871 3684 3872
rect 3688 3871 3689 3875
rect 3683 3870 3689 3871
rect 3706 3875 3712 3876
rect 3706 3871 3707 3875
rect 3711 3874 3712 3875
rect 3795 3875 3801 3876
rect 3795 3874 3796 3875
rect 3711 3872 3796 3874
rect 3711 3871 3712 3872
rect 3706 3870 3712 3871
rect 3795 3871 3796 3872
rect 3800 3871 3801 3875
rect 3795 3870 3801 3871
rect 2880 3868 2894 3870
rect 2880 3867 2881 3868
rect 2875 3866 2881 3867
rect 2892 3866 2894 3868
rect 2959 3867 2965 3868
rect 2959 3866 2960 3867
rect 2892 3864 2960 3866
rect 2959 3863 2960 3864
rect 2964 3863 2965 3867
rect 2959 3862 2965 3863
rect 110 3852 116 3853
rect 2006 3852 2012 3853
rect 110 3848 111 3852
rect 115 3848 116 3852
rect 110 3847 116 3848
rect 334 3851 340 3852
rect 334 3847 335 3851
rect 339 3847 340 3851
rect 334 3846 340 3847
rect 454 3851 460 3852
rect 454 3847 455 3851
rect 459 3847 460 3851
rect 454 3846 460 3847
rect 582 3851 588 3852
rect 582 3847 583 3851
rect 587 3847 588 3851
rect 582 3846 588 3847
rect 718 3851 724 3852
rect 718 3847 719 3851
rect 723 3847 724 3851
rect 718 3846 724 3847
rect 846 3851 852 3852
rect 846 3847 847 3851
rect 851 3847 852 3851
rect 846 3846 852 3847
rect 974 3851 980 3852
rect 974 3847 975 3851
rect 979 3847 980 3851
rect 974 3846 980 3847
rect 1102 3851 1108 3852
rect 1102 3847 1103 3851
rect 1107 3847 1108 3851
rect 1102 3846 1108 3847
rect 1230 3851 1236 3852
rect 1230 3847 1231 3851
rect 1235 3847 1236 3851
rect 1230 3846 1236 3847
rect 1358 3851 1364 3852
rect 1358 3847 1359 3851
rect 1363 3847 1364 3851
rect 1358 3846 1364 3847
rect 1486 3851 1492 3852
rect 1486 3847 1487 3851
rect 1491 3847 1492 3851
rect 2006 3848 2007 3852
rect 2011 3848 2012 3852
rect 2006 3847 2012 3848
rect 2259 3851 2265 3852
rect 2259 3847 2260 3851
rect 2264 3850 2265 3851
rect 2294 3851 2300 3852
rect 2294 3850 2295 3851
rect 2264 3848 2295 3850
rect 2264 3847 2265 3848
rect 1486 3846 1492 3847
rect 2259 3846 2265 3847
rect 2294 3847 2295 3848
rect 2299 3847 2300 3851
rect 2294 3846 2300 3847
rect 2395 3851 2401 3852
rect 2395 3847 2396 3851
rect 2400 3850 2401 3851
rect 2426 3851 2432 3852
rect 2426 3850 2427 3851
rect 2400 3848 2427 3850
rect 2400 3847 2401 3848
rect 2395 3846 2401 3847
rect 2426 3847 2427 3848
rect 2431 3847 2432 3851
rect 2426 3846 2432 3847
rect 2539 3851 2545 3852
rect 2539 3847 2540 3851
rect 2544 3850 2545 3851
rect 2570 3851 2576 3852
rect 2570 3850 2571 3851
rect 2544 3848 2571 3850
rect 2544 3847 2545 3848
rect 2539 3846 2545 3847
rect 2570 3847 2571 3848
rect 2575 3847 2576 3851
rect 2570 3846 2576 3847
rect 2699 3851 2705 3852
rect 2699 3847 2700 3851
rect 2704 3850 2705 3851
rect 2767 3851 2773 3852
rect 2767 3850 2768 3851
rect 2704 3848 2768 3850
rect 2704 3847 2705 3848
rect 2699 3846 2705 3847
rect 2767 3847 2768 3848
rect 2772 3847 2773 3851
rect 2767 3846 2773 3847
rect 2782 3851 2788 3852
rect 2782 3847 2783 3851
rect 2787 3850 2788 3851
rect 2875 3851 2881 3852
rect 2875 3850 2876 3851
rect 2787 3848 2876 3850
rect 2787 3847 2788 3848
rect 2782 3846 2788 3847
rect 2875 3847 2876 3848
rect 2880 3847 2881 3851
rect 2875 3846 2881 3847
rect 3067 3851 3073 3852
rect 3067 3847 3068 3851
rect 3072 3850 3073 3851
rect 3098 3851 3104 3852
rect 3098 3850 3099 3851
rect 3072 3848 3099 3850
rect 3072 3847 3073 3848
rect 3067 3846 3073 3847
rect 3098 3847 3099 3848
rect 3103 3847 3104 3851
rect 3098 3846 3104 3847
rect 3275 3851 3281 3852
rect 3275 3847 3276 3851
rect 3280 3850 3281 3851
rect 3310 3851 3316 3852
rect 3310 3850 3311 3851
rect 3280 3848 3311 3850
rect 3280 3847 3281 3848
rect 3275 3846 3281 3847
rect 3310 3847 3311 3848
rect 3315 3847 3316 3851
rect 3310 3846 3316 3847
rect 3394 3851 3400 3852
rect 3394 3847 3395 3851
rect 3399 3850 3400 3851
rect 3491 3851 3497 3852
rect 3491 3850 3492 3851
rect 3399 3848 3492 3850
rect 3399 3847 3400 3848
rect 3394 3846 3400 3847
rect 3491 3847 3492 3848
rect 3496 3847 3497 3851
rect 3491 3846 3497 3847
rect 3707 3851 3716 3852
rect 3707 3847 3708 3851
rect 3715 3847 3716 3851
rect 3707 3846 3716 3847
rect 266 3843 272 3844
rect 266 3839 267 3843
rect 271 3842 272 3843
rect 439 3843 445 3844
rect 271 3840 377 3842
rect 271 3839 272 3840
rect 266 3838 272 3839
rect 439 3839 440 3843
rect 444 3842 445 3843
rect 567 3843 573 3844
rect 444 3840 497 3842
rect 444 3839 445 3840
rect 439 3838 445 3839
rect 567 3839 568 3843
rect 572 3842 573 3843
rect 1178 3843 1184 3844
rect 572 3840 625 3842
rect 572 3839 573 3840
rect 567 3838 573 3839
rect 794 3839 800 3840
rect 110 3835 116 3836
rect 110 3831 111 3835
rect 115 3831 116 3835
rect 794 3835 795 3839
rect 799 3835 800 3839
rect 794 3834 800 3835
rect 922 3839 928 3840
rect 922 3835 923 3839
rect 927 3835 928 3839
rect 922 3834 928 3835
rect 1050 3839 1056 3840
rect 1050 3835 1051 3839
rect 1055 3835 1056 3839
rect 1178 3839 1179 3843
rect 1183 3839 1184 3843
rect 1178 3838 1184 3839
rect 1214 3843 1220 3844
rect 1214 3839 1215 3843
rect 1219 3842 1220 3843
rect 1342 3843 1348 3844
rect 1219 3840 1273 3842
rect 1219 3839 1220 3840
rect 1214 3838 1220 3839
rect 1342 3839 1343 3843
rect 1347 3842 1348 3843
rect 1471 3843 1477 3844
rect 1347 3840 1401 3842
rect 1347 3839 1348 3840
rect 1342 3838 1348 3839
rect 1471 3839 1472 3843
rect 1476 3842 1477 3843
rect 1476 3840 1529 3842
rect 1476 3839 1477 3840
rect 1471 3838 1477 3839
rect 1050 3834 1056 3835
rect 2006 3835 2012 3836
rect 110 3830 116 3831
rect 334 3832 340 3833
rect 334 3828 335 3832
rect 339 3828 340 3832
rect 334 3827 340 3828
rect 454 3832 460 3833
rect 454 3828 455 3832
rect 459 3828 460 3832
rect 454 3827 460 3828
rect 582 3832 588 3833
rect 582 3828 583 3832
rect 587 3828 588 3832
rect 582 3827 588 3828
rect 718 3832 724 3833
rect 718 3828 719 3832
rect 723 3828 724 3832
rect 718 3827 724 3828
rect 846 3832 852 3833
rect 846 3828 847 3832
rect 851 3828 852 3832
rect 846 3827 852 3828
rect 974 3832 980 3833
rect 974 3828 975 3832
rect 979 3828 980 3832
rect 974 3827 980 3828
rect 1102 3832 1108 3833
rect 1102 3828 1103 3832
rect 1107 3828 1108 3832
rect 1102 3827 1108 3828
rect 1230 3832 1236 3833
rect 1230 3828 1231 3832
rect 1235 3828 1236 3832
rect 1230 3827 1236 3828
rect 1358 3832 1364 3833
rect 1358 3828 1359 3832
rect 1363 3828 1364 3832
rect 1358 3827 1364 3828
rect 1486 3832 1492 3833
rect 1486 3828 1487 3832
rect 1491 3828 1492 3832
rect 2006 3831 2007 3835
rect 2011 3831 2012 3835
rect 2006 3830 2012 3831
rect 1486 3827 1492 3828
rect 2206 3828 2212 3829
rect 2046 3825 2052 3826
rect 2046 3821 2047 3825
rect 2051 3821 2052 3825
rect 2206 3824 2207 3828
rect 2211 3824 2212 3828
rect 2206 3823 2212 3824
rect 2342 3828 2348 3829
rect 2342 3824 2343 3828
rect 2347 3824 2348 3828
rect 2342 3823 2348 3824
rect 2486 3828 2492 3829
rect 2486 3824 2487 3828
rect 2491 3824 2492 3828
rect 2486 3823 2492 3824
rect 2646 3828 2652 3829
rect 2646 3824 2647 3828
rect 2651 3824 2652 3828
rect 2646 3823 2652 3824
rect 2822 3828 2828 3829
rect 2822 3824 2823 3828
rect 2827 3824 2828 3828
rect 2822 3823 2828 3824
rect 3014 3828 3020 3829
rect 3014 3824 3015 3828
rect 3019 3824 3020 3828
rect 3014 3823 3020 3824
rect 3222 3828 3228 3829
rect 3222 3824 3223 3828
rect 3227 3824 3228 3828
rect 3222 3823 3228 3824
rect 3438 3828 3444 3829
rect 3438 3824 3439 3828
rect 3443 3824 3444 3828
rect 3438 3823 3444 3824
rect 3654 3828 3660 3829
rect 3654 3824 3655 3828
rect 3659 3824 3660 3828
rect 3654 3823 3660 3824
rect 3942 3825 3948 3826
rect 2046 3820 2052 3821
rect 3942 3821 3943 3825
rect 3947 3821 3948 3825
rect 3942 3820 3948 3821
rect 954 3819 960 3820
rect 954 3818 955 3819
rect 788 3816 955 3818
rect 387 3811 393 3812
rect 387 3807 388 3811
rect 392 3810 393 3811
rect 439 3811 445 3812
rect 439 3810 440 3811
rect 392 3808 440 3810
rect 392 3807 393 3808
rect 387 3806 393 3807
rect 439 3807 440 3808
rect 444 3807 445 3811
rect 439 3806 445 3807
rect 507 3811 513 3812
rect 507 3807 508 3811
rect 512 3810 513 3811
rect 567 3811 573 3812
rect 567 3810 568 3811
rect 512 3808 568 3810
rect 512 3807 513 3808
rect 507 3806 513 3807
rect 567 3807 568 3808
rect 572 3807 573 3811
rect 771 3811 777 3812
rect 567 3806 573 3807
rect 635 3807 641 3808
rect 635 3806 636 3807
rect 584 3804 636 3806
rect 574 3803 580 3804
rect 574 3799 575 3803
rect 579 3802 580 3803
rect 584 3802 586 3804
rect 635 3803 636 3804
rect 640 3803 641 3807
rect 771 3807 772 3811
rect 776 3810 777 3811
rect 788 3810 790 3816
rect 954 3815 955 3816
rect 959 3815 960 3819
rect 954 3814 960 3815
rect 2274 3819 2280 3820
rect 2274 3815 2275 3819
rect 2279 3815 2280 3819
rect 2274 3814 2280 3815
rect 2294 3819 2300 3820
rect 2294 3815 2295 3819
rect 2299 3818 2300 3819
rect 2426 3819 2432 3820
rect 2299 3816 2385 3818
rect 2299 3815 2300 3816
rect 2294 3814 2300 3815
rect 2426 3815 2427 3819
rect 2431 3818 2432 3819
rect 2570 3819 2576 3820
rect 2431 3816 2529 3818
rect 2431 3815 2432 3816
rect 2426 3814 2432 3815
rect 2570 3815 2571 3819
rect 2575 3818 2576 3819
rect 2767 3819 2773 3820
rect 2575 3816 2689 3818
rect 2575 3815 2576 3816
rect 2570 3814 2576 3815
rect 2767 3815 2768 3819
rect 2772 3818 2773 3819
rect 2959 3819 2965 3820
rect 2772 3816 2865 3818
rect 2772 3815 2773 3816
rect 2767 3814 2773 3815
rect 2959 3815 2960 3819
rect 2964 3818 2965 3819
rect 3098 3819 3104 3820
rect 2964 3816 3057 3818
rect 2964 3815 2965 3816
rect 2959 3814 2965 3815
rect 3098 3815 3099 3819
rect 3103 3818 3104 3819
rect 3310 3819 3316 3820
rect 3103 3816 3265 3818
rect 3103 3815 3104 3816
rect 3098 3814 3104 3815
rect 3310 3815 3311 3819
rect 3315 3818 3316 3819
rect 3730 3819 3736 3820
rect 3315 3816 3481 3818
rect 3315 3815 3316 3816
rect 3310 3814 3316 3815
rect 3730 3815 3731 3819
rect 3735 3815 3736 3819
rect 3730 3814 3736 3815
rect 776 3808 790 3810
rect 794 3811 800 3812
rect 776 3807 777 3808
rect 771 3806 777 3807
rect 794 3807 795 3811
rect 799 3810 800 3811
rect 899 3811 905 3812
rect 899 3810 900 3811
rect 799 3808 900 3810
rect 799 3807 800 3808
rect 794 3806 800 3807
rect 899 3807 900 3808
rect 904 3807 905 3811
rect 899 3806 905 3807
rect 922 3811 928 3812
rect 922 3807 923 3811
rect 927 3810 928 3811
rect 1027 3811 1033 3812
rect 1027 3810 1028 3811
rect 927 3808 1028 3810
rect 927 3807 928 3808
rect 922 3806 928 3807
rect 1027 3807 1028 3808
rect 1032 3807 1033 3811
rect 1027 3806 1033 3807
rect 1155 3811 1161 3812
rect 1155 3807 1156 3811
rect 1160 3810 1161 3811
rect 1214 3811 1220 3812
rect 1214 3810 1215 3811
rect 1160 3808 1215 3810
rect 1160 3807 1161 3808
rect 1155 3806 1161 3807
rect 1214 3807 1215 3808
rect 1219 3807 1220 3811
rect 1214 3806 1220 3807
rect 1283 3811 1289 3812
rect 1283 3807 1284 3811
rect 1288 3810 1289 3811
rect 1342 3811 1348 3812
rect 1342 3810 1343 3811
rect 1288 3808 1343 3810
rect 1288 3807 1289 3808
rect 1283 3806 1289 3807
rect 1342 3807 1343 3808
rect 1347 3807 1348 3811
rect 1342 3806 1348 3807
rect 1411 3811 1417 3812
rect 1411 3807 1412 3811
rect 1416 3810 1417 3811
rect 1471 3811 1477 3812
rect 1471 3810 1472 3811
rect 1416 3808 1472 3810
rect 1416 3807 1417 3808
rect 1411 3806 1417 3807
rect 1471 3807 1472 3808
rect 1476 3807 1477 3811
rect 2206 3809 2212 3810
rect 2046 3808 2052 3809
rect 1471 3806 1477 3807
rect 1506 3807 1512 3808
rect 635 3802 641 3803
rect 1506 3803 1507 3807
rect 1511 3806 1512 3807
rect 1539 3807 1545 3808
rect 1539 3806 1540 3807
rect 1511 3804 1540 3806
rect 1511 3803 1512 3804
rect 1506 3802 1512 3803
rect 1539 3803 1540 3804
rect 1544 3803 1545 3807
rect 2046 3804 2047 3808
rect 2051 3804 2052 3808
rect 2206 3805 2207 3809
rect 2211 3805 2212 3809
rect 2206 3804 2212 3805
rect 2342 3809 2348 3810
rect 2342 3805 2343 3809
rect 2347 3805 2348 3809
rect 2342 3804 2348 3805
rect 2486 3809 2492 3810
rect 2486 3805 2487 3809
rect 2491 3805 2492 3809
rect 2486 3804 2492 3805
rect 2646 3809 2652 3810
rect 2646 3805 2647 3809
rect 2651 3805 2652 3809
rect 2646 3804 2652 3805
rect 2822 3809 2828 3810
rect 2822 3805 2823 3809
rect 2827 3805 2828 3809
rect 2822 3804 2828 3805
rect 3014 3809 3020 3810
rect 3014 3805 3015 3809
rect 3019 3805 3020 3809
rect 3014 3804 3020 3805
rect 3222 3809 3228 3810
rect 3222 3805 3223 3809
rect 3227 3805 3228 3809
rect 3222 3804 3228 3805
rect 3438 3809 3444 3810
rect 3438 3805 3439 3809
rect 3443 3805 3444 3809
rect 3438 3804 3444 3805
rect 3654 3809 3660 3810
rect 3654 3805 3655 3809
rect 3659 3805 3660 3809
rect 3654 3804 3660 3805
rect 3942 3808 3948 3809
rect 3942 3804 3943 3808
rect 3947 3804 3948 3808
rect 2046 3803 2052 3804
rect 3942 3803 3948 3804
rect 1539 3802 1545 3803
rect 579 3800 586 3802
rect 579 3799 580 3800
rect 574 3798 580 3799
rect 555 3791 561 3792
rect 555 3787 556 3791
rect 560 3790 561 3791
rect 590 3791 596 3792
rect 590 3790 591 3791
rect 560 3788 591 3790
rect 560 3787 561 3788
rect 555 3786 561 3787
rect 590 3787 591 3788
rect 595 3787 596 3791
rect 590 3786 596 3787
rect 667 3791 673 3792
rect 667 3787 668 3791
rect 672 3790 673 3791
rect 698 3791 704 3792
rect 698 3790 699 3791
rect 672 3788 699 3790
rect 672 3787 673 3788
rect 667 3786 673 3787
rect 698 3787 699 3788
rect 703 3787 704 3791
rect 698 3786 704 3787
rect 787 3791 793 3792
rect 787 3787 788 3791
rect 792 3790 793 3791
rect 818 3791 824 3792
rect 818 3790 819 3791
rect 792 3788 819 3790
rect 792 3787 793 3788
rect 787 3786 793 3787
rect 818 3787 819 3788
rect 823 3787 824 3791
rect 818 3786 824 3787
rect 902 3791 908 3792
rect 902 3787 903 3791
rect 907 3790 908 3791
rect 915 3791 921 3792
rect 915 3790 916 3791
rect 907 3788 916 3790
rect 907 3787 908 3788
rect 902 3786 908 3787
rect 915 3787 916 3788
rect 920 3787 921 3791
rect 915 3786 921 3787
rect 1050 3791 1057 3792
rect 1050 3787 1051 3791
rect 1056 3787 1057 3791
rect 1050 3786 1057 3787
rect 1074 3791 1080 3792
rect 1074 3787 1075 3791
rect 1079 3790 1080 3791
rect 1195 3791 1201 3792
rect 1195 3790 1196 3791
rect 1079 3788 1196 3790
rect 1079 3787 1080 3788
rect 1074 3786 1080 3787
rect 1195 3787 1196 3788
rect 1200 3787 1201 3791
rect 1406 3791 1412 3792
rect 1195 3786 1201 3787
rect 1339 3789 1345 3790
rect 1339 3785 1340 3789
rect 1344 3785 1345 3789
rect 1406 3787 1407 3791
rect 1411 3790 1412 3791
rect 1483 3791 1489 3792
rect 1483 3790 1484 3791
rect 1411 3788 1484 3790
rect 1411 3787 1412 3788
rect 1406 3786 1412 3787
rect 1483 3787 1484 3788
rect 1488 3787 1489 3791
rect 1483 3786 1489 3787
rect 1570 3791 1576 3792
rect 1570 3787 1571 3791
rect 1575 3790 1576 3791
rect 1635 3791 1641 3792
rect 1635 3790 1636 3791
rect 1575 3788 1636 3790
rect 1575 3787 1576 3788
rect 1570 3786 1576 3787
rect 1635 3787 1636 3788
rect 1640 3787 1641 3791
rect 1635 3786 1641 3787
rect 1339 3784 1345 3785
rect 1340 3782 1342 3784
rect 1514 3783 1520 3784
rect 1514 3782 1515 3783
rect 1340 3780 1515 3782
rect 1514 3779 1515 3780
rect 1519 3779 1520 3783
rect 1514 3778 1520 3779
rect 502 3768 508 3769
rect 110 3765 116 3766
rect 110 3761 111 3765
rect 115 3761 116 3765
rect 502 3764 503 3768
rect 507 3764 508 3768
rect 502 3763 508 3764
rect 614 3768 620 3769
rect 614 3764 615 3768
rect 619 3764 620 3768
rect 614 3763 620 3764
rect 734 3768 740 3769
rect 734 3764 735 3768
rect 739 3764 740 3768
rect 734 3763 740 3764
rect 862 3768 868 3769
rect 862 3764 863 3768
rect 867 3764 868 3768
rect 862 3763 868 3764
rect 998 3768 1004 3769
rect 998 3764 999 3768
rect 1003 3764 1004 3768
rect 998 3763 1004 3764
rect 1142 3768 1148 3769
rect 1142 3764 1143 3768
rect 1147 3764 1148 3768
rect 1142 3763 1148 3764
rect 1286 3768 1292 3769
rect 1286 3764 1287 3768
rect 1291 3764 1292 3768
rect 1286 3763 1292 3764
rect 1430 3768 1436 3769
rect 1430 3764 1431 3768
rect 1435 3764 1436 3768
rect 1430 3763 1436 3764
rect 1582 3768 1588 3769
rect 1582 3764 1583 3768
rect 1587 3764 1588 3768
rect 1582 3763 1588 3764
rect 2006 3765 2012 3766
rect 110 3760 116 3761
rect 2006 3761 2007 3765
rect 2011 3761 2012 3765
rect 2006 3760 2012 3761
rect 574 3759 580 3760
rect 574 3755 575 3759
rect 579 3755 580 3759
rect 574 3754 580 3755
rect 590 3759 596 3760
rect 590 3755 591 3759
rect 595 3758 596 3759
rect 698 3759 704 3760
rect 595 3756 657 3758
rect 595 3755 596 3756
rect 590 3754 596 3755
rect 698 3755 699 3759
rect 703 3758 704 3759
rect 818 3759 824 3760
rect 703 3756 777 3758
rect 703 3755 704 3756
rect 698 3754 704 3755
rect 818 3755 819 3759
rect 823 3758 824 3759
rect 1074 3759 1080 3760
rect 823 3756 905 3758
rect 823 3755 824 3756
rect 818 3754 824 3755
rect 1074 3755 1075 3759
rect 1079 3755 1080 3759
rect 1074 3754 1080 3755
rect 1218 3759 1224 3760
rect 1218 3755 1219 3759
rect 1223 3755 1224 3759
rect 1406 3759 1412 3760
rect 1406 3758 1407 3759
rect 1365 3756 1407 3758
rect 1218 3754 1224 3755
rect 1406 3755 1407 3756
rect 1411 3755 1412 3759
rect 1406 3754 1412 3755
rect 1506 3759 1512 3760
rect 1506 3755 1507 3759
rect 1511 3755 1512 3759
rect 1506 3754 1512 3755
rect 1514 3759 1520 3760
rect 1514 3755 1515 3759
rect 1519 3758 1520 3759
rect 1519 3756 1625 3758
rect 2046 3756 2052 3757
rect 3942 3756 3948 3757
rect 1519 3755 1520 3756
rect 1514 3754 1520 3755
rect 2046 3752 2047 3756
rect 2051 3752 2052 3756
rect 2046 3751 2052 3752
rect 2190 3755 2196 3756
rect 2190 3751 2191 3755
rect 2195 3751 2196 3755
rect 2190 3750 2196 3751
rect 2374 3755 2380 3756
rect 2374 3751 2375 3755
rect 2379 3751 2380 3755
rect 2374 3750 2380 3751
rect 2558 3755 2564 3756
rect 2558 3751 2559 3755
rect 2563 3751 2564 3755
rect 2558 3750 2564 3751
rect 2742 3755 2748 3756
rect 2742 3751 2743 3755
rect 2747 3751 2748 3755
rect 2742 3750 2748 3751
rect 2934 3755 2940 3756
rect 2934 3751 2935 3755
rect 2939 3751 2940 3755
rect 2934 3750 2940 3751
rect 3126 3755 3132 3756
rect 3126 3751 3127 3755
rect 3131 3751 3132 3755
rect 3126 3750 3132 3751
rect 3318 3755 3324 3756
rect 3318 3751 3319 3755
rect 3323 3751 3324 3755
rect 3318 3750 3324 3751
rect 3510 3755 3516 3756
rect 3510 3751 3511 3755
rect 3515 3751 3516 3755
rect 3510 3750 3516 3751
rect 3710 3755 3716 3756
rect 3710 3751 3711 3755
rect 3715 3751 3716 3755
rect 3942 3752 3943 3756
rect 3947 3752 3948 3756
rect 3942 3751 3948 3752
rect 3710 3750 3716 3751
rect 502 3749 508 3750
rect 110 3748 116 3749
rect 110 3744 111 3748
rect 115 3744 116 3748
rect 502 3745 503 3749
rect 507 3745 508 3749
rect 502 3744 508 3745
rect 614 3749 620 3750
rect 614 3745 615 3749
rect 619 3745 620 3749
rect 614 3744 620 3745
rect 734 3749 740 3750
rect 734 3745 735 3749
rect 739 3745 740 3749
rect 734 3744 740 3745
rect 862 3749 868 3750
rect 862 3745 863 3749
rect 867 3745 868 3749
rect 862 3744 868 3745
rect 998 3749 1004 3750
rect 998 3745 999 3749
rect 1003 3745 1004 3749
rect 998 3744 1004 3745
rect 1142 3749 1148 3750
rect 1142 3745 1143 3749
rect 1147 3745 1148 3749
rect 1142 3744 1148 3745
rect 1286 3749 1292 3750
rect 1286 3745 1287 3749
rect 1291 3745 1292 3749
rect 1286 3744 1292 3745
rect 1430 3749 1436 3750
rect 1430 3745 1431 3749
rect 1435 3745 1436 3749
rect 1430 3744 1436 3745
rect 1582 3749 1588 3750
rect 1582 3745 1583 3749
rect 1587 3745 1588 3749
rect 1582 3744 1588 3745
rect 2006 3748 2012 3749
rect 2006 3744 2007 3748
rect 2011 3744 2012 3748
rect 3394 3747 3400 3748
rect 110 3743 116 3744
rect 2006 3743 2012 3744
rect 2327 3743 2333 3744
rect 2327 3742 2328 3743
rect 2269 3740 2328 3742
rect 2046 3739 2052 3740
rect 2046 3735 2047 3739
rect 2051 3735 2052 3739
rect 2327 3739 2328 3740
rect 2332 3739 2333 3743
rect 2327 3738 2333 3739
rect 2450 3743 2456 3744
rect 2450 3739 2451 3743
rect 2455 3739 2456 3743
rect 2450 3738 2456 3739
rect 2634 3743 2640 3744
rect 2634 3739 2635 3743
rect 2639 3739 2640 3743
rect 2826 3743 2832 3744
rect 2826 3742 2827 3743
rect 2821 3740 2827 3742
rect 2634 3738 2640 3739
rect 2826 3739 2827 3740
rect 2831 3739 2832 3743
rect 2826 3738 2832 3739
rect 3010 3743 3016 3744
rect 3010 3739 3011 3743
rect 3015 3739 3016 3743
rect 3010 3738 3016 3739
rect 3202 3743 3208 3744
rect 3202 3739 3203 3743
rect 3207 3739 3208 3743
rect 3394 3743 3395 3747
rect 3399 3743 3400 3747
rect 3394 3742 3400 3743
rect 3438 3747 3444 3748
rect 3438 3743 3439 3747
rect 3443 3746 3444 3747
rect 3443 3744 3553 3746
rect 3443 3743 3444 3744
rect 3438 3742 3444 3743
rect 3786 3743 3792 3744
rect 3202 3738 3208 3739
rect 3786 3739 3787 3743
rect 3791 3739 3792 3743
rect 3786 3738 3792 3739
rect 3942 3739 3948 3740
rect 2046 3734 2052 3735
rect 2190 3736 2196 3737
rect 2190 3732 2191 3736
rect 2195 3732 2196 3736
rect 2190 3731 2196 3732
rect 2374 3736 2380 3737
rect 2374 3732 2375 3736
rect 2379 3732 2380 3736
rect 2374 3731 2380 3732
rect 2558 3736 2564 3737
rect 2558 3732 2559 3736
rect 2563 3732 2564 3736
rect 2558 3731 2564 3732
rect 2742 3736 2748 3737
rect 2742 3732 2743 3736
rect 2747 3732 2748 3736
rect 2742 3731 2748 3732
rect 2934 3736 2940 3737
rect 2934 3732 2935 3736
rect 2939 3732 2940 3736
rect 2934 3731 2940 3732
rect 3126 3736 3132 3737
rect 3126 3732 3127 3736
rect 3131 3732 3132 3736
rect 3126 3731 3132 3732
rect 3318 3736 3324 3737
rect 3318 3732 3319 3736
rect 3323 3732 3324 3736
rect 3318 3731 3324 3732
rect 3510 3736 3516 3737
rect 3510 3732 3511 3736
rect 3515 3732 3516 3736
rect 3510 3731 3516 3732
rect 3710 3736 3716 3737
rect 3710 3732 3711 3736
rect 3715 3732 3716 3736
rect 3942 3735 3943 3739
rect 3947 3735 3948 3739
rect 3942 3734 3948 3735
rect 3710 3731 3716 3732
rect 3438 3723 3444 3724
rect 3438 3722 3439 3723
rect 3004 3720 3439 3722
rect 2243 3715 2249 3716
rect 2243 3711 2244 3715
rect 2248 3714 2249 3715
rect 2274 3715 2280 3716
rect 2274 3714 2275 3715
rect 2248 3712 2275 3714
rect 2248 3711 2249 3712
rect 2243 3710 2249 3711
rect 2274 3711 2275 3712
rect 2279 3711 2280 3715
rect 2274 3710 2280 3711
rect 2327 3715 2333 3716
rect 2327 3711 2328 3715
rect 2332 3714 2333 3715
rect 2427 3715 2433 3716
rect 2427 3714 2428 3715
rect 2332 3712 2428 3714
rect 2332 3711 2333 3712
rect 2327 3710 2333 3711
rect 2427 3711 2428 3712
rect 2432 3711 2433 3715
rect 2427 3710 2433 3711
rect 2450 3715 2456 3716
rect 2450 3711 2451 3715
rect 2455 3714 2456 3715
rect 2611 3715 2617 3716
rect 2611 3714 2612 3715
rect 2455 3712 2612 3714
rect 2455 3711 2456 3712
rect 2450 3710 2456 3711
rect 2611 3711 2612 3712
rect 2616 3711 2617 3715
rect 2611 3710 2617 3711
rect 2634 3715 2640 3716
rect 2634 3711 2635 3715
rect 2639 3714 2640 3715
rect 2795 3715 2801 3716
rect 2795 3714 2796 3715
rect 2639 3712 2796 3714
rect 2639 3711 2640 3712
rect 2634 3710 2640 3711
rect 2795 3711 2796 3712
rect 2800 3711 2801 3715
rect 2795 3710 2801 3711
rect 2987 3715 2993 3716
rect 2987 3711 2988 3715
rect 2992 3714 2993 3715
rect 3004 3714 3006 3720
rect 3438 3719 3439 3720
rect 3443 3719 3444 3723
rect 3438 3718 3444 3719
rect 2992 3712 3006 3714
rect 3010 3715 3016 3716
rect 2992 3711 2993 3712
rect 2987 3710 2993 3711
rect 3010 3711 3011 3715
rect 3015 3714 3016 3715
rect 3179 3715 3185 3716
rect 3179 3714 3180 3715
rect 3015 3712 3180 3714
rect 3015 3711 3016 3712
rect 3010 3710 3016 3711
rect 3179 3711 3180 3712
rect 3184 3711 3185 3715
rect 3179 3710 3185 3711
rect 3202 3715 3208 3716
rect 3202 3711 3203 3715
rect 3207 3714 3208 3715
rect 3371 3715 3377 3716
rect 3371 3714 3372 3715
rect 3207 3712 3372 3714
rect 3207 3711 3208 3712
rect 3202 3710 3208 3711
rect 3371 3711 3372 3712
rect 3376 3711 3377 3715
rect 3730 3715 3736 3716
rect 3371 3710 3377 3711
rect 3563 3711 3569 3712
rect 3563 3707 3564 3711
rect 3568 3710 3569 3711
rect 3578 3711 3584 3712
rect 3578 3710 3579 3711
rect 3568 3708 3579 3710
rect 3568 3707 3569 3708
rect 3563 3706 3569 3707
rect 3578 3707 3579 3708
rect 3583 3707 3584 3711
rect 3730 3711 3731 3715
rect 3735 3714 3736 3715
rect 3763 3715 3769 3716
rect 3763 3714 3764 3715
rect 3735 3712 3764 3714
rect 3735 3711 3736 3712
rect 3730 3710 3736 3711
rect 3763 3711 3764 3712
rect 3768 3711 3769 3715
rect 3763 3710 3769 3711
rect 3578 3706 3584 3707
rect 2179 3695 2185 3696
rect 2179 3691 2180 3695
rect 2184 3694 2185 3695
rect 2295 3695 2301 3696
rect 2295 3694 2296 3695
rect 2184 3692 2296 3694
rect 2184 3691 2185 3692
rect 2179 3690 2185 3691
rect 2295 3691 2296 3692
rect 2300 3691 2301 3695
rect 2295 3690 2301 3691
rect 2403 3695 2409 3696
rect 2403 3691 2404 3695
rect 2408 3694 2409 3695
rect 2434 3695 2440 3696
rect 2434 3694 2435 3695
rect 2408 3692 2435 3694
rect 2408 3691 2409 3692
rect 2403 3690 2409 3691
rect 2434 3691 2435 3692
rect 2439 3691 2440 3695
rect 2434 3690 2440 3691
rect 2635 3695 2641 3696
rect 2635 3691 2636 3695
rect 2640 3694 2641 3695
rect 2666 3695 2672 3696
rect 2666 3694 2667 3695
rect 2640 3692 2667 3694
rect 2640 3691 2641 3692
rect 2635 3690 2641 3691
rect 2666 3691 2667 3692
rect 2671 3691 2672 3695
rect 2666 3690 2672 3691
rect 2826 3695 2832 3696
rect 2826 3691 2827 3695
rect 2831 3694 2832 3695
rect 2867 3695 2873 3696
rect 2867 3694 2868 3695
rect 2831 3692 2868 3694
rect 2831 3691 2832 3692
rect 2826 3690 2832 3691
rect 2867 3691 2868 3692
rect 2872 3691 2873 3695
rect 3142 3695 3148 3696
rect 2867 3690 2873 3691
rect 3099 3693 3105 3694
rect 3099 3689 3100 3693
rect 3104 3689 3105 3693
rect 3142 3691 3143 3695
rect 3147 3694 3148 3695
rect 3331 3695 3337 3696
rect 3331 3694 3332 3695
rect 3147 3692 3332 3694
rect 3147 3691 3148 3692
rect 3142 3690 3148 3691
rect 3331 3691 3332 3692
rect 3336 3691 3337 3695
rect 3331 3690 3337 3691
rect 3354 3695 3360 3696
rect 3354 3691 3355 3695
rect 3359 3694 3360 3695
rect 3563 3695 3569 3696
rect 3563 3694 3564 3695
rect 3359 3692 3564 3694
rect 3359 3691 3360 3692
rect 3354 3690 3360 3691
rect 3563 3691 3564 3692
rect 3568 3691 3569 3695
rect 3563 3690 3569 3691
rect 3786 3695 3792 3696
rect 3786 3691 3787 3695
rect 3791 3694 3792 3695
rect 3803 3695 3809 3696
rect 3803 3694 3804 3695
rect 3791 3692 3804 3694
rect 3791 3691 3792 3692
rect 3786 3690 3792 3691
rect 3803 3691 3804 3692
rect 3808 3691 3809 3695
rect 3803 3690 3809 3691
rect 110 3688 116 3689
rect 2006 3688 2012 3689
rect 3099 3688 3105 3689
rect 110 3684 111 3688
rect 115 3684 116 3688
rect 110 3683 116 3684
rect 494 3687 500 3688
rect 494 3683 495 3687
rect 499 3683 500 3687
rect 494 3682 500 3683
rect 590 3687 596 3688
rect 590 3683 591 3687
rect 595 3683 596 3687
rect 590 3682 596 3683
rect 686 3687 692 3688
rect 686 3683 687 3687
rect 691 3683 692 3687
rect 686 3682 692 3683
rect 790 3687 796 3688
rect 790 3683 791 3687
rect 795 3683 796 3687
rect 790 3682 796 3683
rect 910 3687 916 3688
rect 910 3683 911 3687
rect 915 3683 916 3687
rect 910 3682 916 3683
rect 1038 3687 1044 3688
rect 1038 3683 1039 3687
rect 1043 3683 1044 3687
rect 1038 3682 1044 3683
rect 1182 3687 1188 3688
rect 1182 3683 1183 3687
rect 1187 3683 1188 3687
rect 1182 3682 1188 3683
rect 1334 3687 1340 3688
rect 1334 3683 1335 3687
rect 1339 3683 1340 3687
rect 1334 3682 1340 3683
rect 1494 3687 1500 3688
rect 1494 3683 1495 3687
rect 1499 3683 1500 3687
rect 1494 3682 1500 3683
rect 1654 3687 1660 3688
rect 1654 3683 1655 3687
rect 1659 3683 1660 3687
rect 2006 3684 2007 3688
rect 2011 3684 2012 3688
rect 3100 3686 3102 3688
rect 3378 3687 3384 3688
rect 3378 3686 3379 3687
rect 3100 3684 3379 3686
rect 2006 3683 2012 3684
rect 3378 3683 3379 3684
rect 3383 3683 3384 3687
rect 1654 3682 1660 3683
rect 3378 3682 3384 3683
rect 902 3679 908 3680
rect 570 3675 576 3676
rect 110 3671 116 3672
rect 110 3667 111 3671
rect 115 3667 116 3671
rect 570 3671 571 3675
rect 575 3671 576 3675
rect 570 3670 576 3671
rect 666 3675 672 3676
rect 666 3671 667 3675
rect 671 3671 672 3675
rect 666 3670 672 3671
rect 762 3675 768 3676
rect 762 3671 763 3675
rect 767 3671 768 3675
rect 762 3670 768 3671
rect 866 3675 872 3676
rect 866 3671 867 3675
rect 871 3671 872 3675
rect 902 3675 903 3679
rect 907 3678 908 3679
rect 1266 3679 1272 3680
rect 907 3676 953 3678
rect 907 3675 908 3676
rect 902 3674 908 3675
rect 1114 3675 1120 3676
rect 866 3670 872 3671
rect 1114 3671 1115 3675
rect 1119 3671 1120 3675
rect 1114 3670 1120 3671
rect 1258 3675 1264 3676
rect 1258 3671 1259 3675
rect 1263 3671 1264 3675
rect 1266 3675 1267 3679
rect 1271 3678 1272 3679
rect 1570 3679 1576 3680
rect 1271 3676 1377 3678
rect 1271 3675 1272 3676
rect 1266 3674 1272 3675
rect 1570 3675 1571 3679
rect 1575 3675 1576 3679
rect 1570 3674 1576 3675
rect 1614 3679 1620 3680
rect 1614 3675 1615 3679
rect 1619 3678 1620 3679
rect 1619 3676 1697 3678
rect 1619 3675 1620 3676
rect 1614 3674 1620 3675
rect 2126 3672 2132 3673
rect 1258 3670 1264 3671
rect 2006 3671 2012 3672
rect 110 3666 116 3667
rect 494 3668 500 3669
rect 494 3664 495 3668
rect 499 3664 500 3668
rect 494 3663 500 3664
rect 590 3668 596 3669
rect 590 3664 591 3668
rect 595 3664 596 3668
rect 590 3663 596 3664
rect 686 3668 692 3669
rect 686 3664 687 3668
rect 691 3664 692 3668
rect 686 3663 692 3664
rect 790 3668 796 3669
rect 790 3664 791 3668
rect 795 3664 796 3668
rect 790 3663 796 3664
rect 910 3668 916 3669
rect 910 3664 911 3668
rect 915 3664 916 3668
rect 910 3663 916 3664
rect 1038 3668 1044 3669
rect 1038 3664 1039 3668
rect 1043 3664 1044 3668
rect 1038 3663 1044 3664
rect 1182 3668 1188 3669
rect 1182 3664 1183 3668
rect 1187 3664 1188 3668
rect 1182 3663 1188 3664
rect 1334 3668 1340 3669
rect 1334 3664 1335 3668
rect 1339 3664 1340 3668
rect 1334 3663 1340 3664
rect 1494 3668 1500 3669
rect 1494 3664 1495 3668
rect 1499 3664 1500 3668
rect 1494 3663 1500 3664
rect 1654 3668 1660 3669
rect 1654 3664 1655 3668
rect 1659 3664 1660 3668
rect 2006 3667 2007 3671
rect 2011 3667 2012 3671
rect 2006 3666 2012 3667
rect 2046 3669 2052 3670
rect 2046 3665 2047 3669
rect 2051 3665 2052 3669
rect 2126 3668 2127 3672
rect 2131 3668 2132 3672
rect 2126 3667 2132 3668
rect 2350 3672 2356 3673
rect 2350 3668 2351 3672
rect 2355 3668 2356 3672
rect 2350 3667 2356 3668
rect 2582 3672 2588 3673
rect 2582 3668 2583 3672
rect 2587 3668 2588 3672
rect 2582 3667 2588 3668
rect 2814 3672 2820 3673
rect 2814 3668 2815 3672
rect 2819 3668 2820 3672
rect 2814 3667 2820 3668
rect 3046 3672 3052 3673
rect 3046 3668 3047 3672
rect 3051 3668 3052 3672
rect 3046 3667 3052 3668
rect 3278 3672 3284 3673
rect 3278 3668 3279 3672
rect 3283 3668 3284 3672
rect 3278 3667 3284 3668
rect 3510 3672 3516 3673
rect 3510 3668 3511 3672
rect 3515 3668 3516 3672
rect 3510 3667 3516 3668
rect 3750 3672 3756 3673
rect 3750 3668 3751 3672
rect 3755 3668 3756 3672
rect 3750 3667 3756 3668
rect 3942 3669 3948 3670
rect 2046 3664 2052 3665
rect 3942 3665 3943 3669
rect 3947 3665 3948 3669
rect 3942 3664 3948 3665
rect 1654 3663 1660 3664
rect 2202 3663 2208 3664
rect 2202 3659 2203 3663
rect 2207 3659 2208 3663
rect 2202 3658 2208 3659
rect 2295 3663 2301 3664
rect 2295 3659 2296 3663
rect 2300 3662 2301 3663
rect 2434 3663 2440 3664
rect 2300 3660 2393 3662
rect 2300 3659 2301 3660
rect 2295 3658 2301 3659
rect 2434 3659 2435 3663
rect 2439 3662 2440 3663
rect 2666 3663 2672 3664
rect 2439 3660 2625 3662
rect 2439 3659 2440 3660
rect 2434 3658 2440 3659
rect 2666 3659 2667 3663
rect 2671 3662 2672 3663
rect 3142 3663 3148 3664
rect 3142 3662 3143 3663
rect 2671 3660 2857 3662
rect 3125 3660 3143 3662
rect 2671 3659 2672 3660
rect 2666 3658 2672 3659
rect 3142 3659 3143 3660
rect 3147 3659 3148 3663
rect 3142 3658 3148 3659
rect 3354 3663 3360 3664
rect 3354 3659 3355 3663
rect 3359 3659 3360 3663
rect 3354 3658 3360 3659
rect 3578 3663 3584 3664
rect 3578 3659 3579 3663
rect 3583 3659 3584 3663
rect 3578 3658 3584 3659
rect 3826 3663 3832 3664
rect 3826 3659 3827 3663
rect 3831 3659 3832 3663
rect 3826 3658 3832 3659
rect 1266 3655 1272 3656
rect 1266 3654 1267 3655
rect 1159 3652 1267 3654
rect 570 3647 576 3648
rect 547 3643 553 3644
rect 547 3639 548 3643
rect 552 3642 553 3643
rect 570 3643 571 3647
rect 575 3646 576 3647
rect 643 3647 649 3648
rect 643 3646 644 3647
rect 575 3644 644 3646
rect 575 3643 576 3644
rect 570 3642 576 3643
rect 643 3643 644 3644
rect 648 3643 649 3647
rect 643 3642 649 3643
rect 666 3647 672 3648
rect 666 3643 667 3647
rect 671 3646 672 3647
rect 739 3647 745 3648
rect 739 3646 740 3647
rect 671 3644 740 3646
rect 671 3643 672 3644
rect 666 3642 672 3643
rect 739 3643 740 3644
rect 744 3643 745 3647
rect 739 3642 745 3643
rect 762 3647 768 3648
rect 762 3643 763 3647
rect 767 3646 768 3647
rect 843 3647 849 3648
rect 843 3646 844 3647
rect 767 3644 844 3646
rect 767 3643 768 3644
rect 762 3642 768 3643
rect 843 3643 844 3644
rect 848 3643 849 3647
rect 843 3642 849 3643
rect 866 3647 872 3648
rect 866 3643 867 3647
rect 871 3646 872 3647
rect 963 3647 969 3648
rect 963 3646 964 3647
rect 871 3644 964 3646
rect 871 3643 872 3644
rect 866 3642 872 3643
rect 963 3643 964 3644
rect 968 3643 969 3647
rect 963 3642 969 3643
rect 1091 3647 1097 3648
rect 1091 3643 1092 3647
rect 1096 3646 1097 3647
rect 1159 3646 1161 3652
rect 1266 3651 1267 3652
rect 1271 3651 1272 3655
rect 2126 3653 2132 3654
rect 1266 3650 1272 3651
rect 2046 3652 2052 3653
rect 2046 3648 2047 3652
rect 2051 3648 2052 3652
rect 2126 3649 2127 3653
rect 2131 3649 2132 3653
rect 2126 3648 2132 3649
rect 2350 3653 2356 3654
rect 2350 3649 2351 3653
rect 2355 3649 2356 3653
rect 2350 3648 2356 3649
rect 2582 3653 2588 3654
rect 2582 3649 2583 3653
rect 2587 3649 2588 3653
rect 2582 3648 2588 3649
rect 2814 3653 2820 3654
rect 2814 3649 2815 3653
rect 2819 3649 2820 3653
rect 2814 3648 2820 3649
rect 3046 3653 3052 3654
rect 3046 3649 3047 3653
rect 3051 3649 3052 3653
rect 3046 3648 3052 3649
rect 3278 3653 3284 3654
rect 3278 3649 3279 3653
rect 3283 3649 3284 3653
rect 3278 3648 3284 3649
rect 3510 3653 3516 3654
rect 3510 3649 3511 3653
rect 3515 3649 3516 3653
rect 3510 3648 3516 3649
rect 3750 3653 3756 3654
rect 3750 3649 3751 3653
rect 3755 3649 3756 3653
rect 3750 3648 3756 3649
rect 3942 3652 3948 3653
rect 3942 3648 3943 3652
rect 3947 3648 3948 3652
rect 1096 3644 1161 3646
rect 1218 3647 1224 3648
rect 1096 3643 1097 3644
rect 1091 3642 1097 3643
rect 1218 3643 1219 3647
rect 1223 3646 1224 3647
rect 1235 3647 1241 3648
rect 1235 3646 1236 3647
rect 1223 3644 1236 3646
rect 1223 3643 1224 3644
rect 1218 3642 1224 3643
rect 1235 3643 1236 3644
rect 1240 3643 1241 3647
rect 1235 3642 1241 3643
rect 1258 3647 1264 3648
rect 1258 3643 1259 3647
rect 1263 3646 1264 3647
rect 1387 3647 1393 3648
rect 1387 3646 1388 3647
rect 1263 3644 1388 3646
rect 1263 3643 1264 3644
rect 1258 3642 1264 3643
rect 1387 3643 1388 3644
rect 1392 3643 1393 3647
rect 1387 3642 1393 3643
rect 1547 3647 1553 3648
rect 1547 3643 1548 3647
rect 1552 3646 1553 3647
rect 1614 3647 1620 3648
rect 2046 3647 2052 3648
rect 3942 3647 3948 3648
rect 1614 3646 1615 3647
rect 1552 3644 1615 3646
rect 1552 3643 1553 3644
rect 1547 3642 1553 3643
rect 1614 3643 1615 3644
rect 1619 3643 1620 3647
rect 1614 3642 1620 3643
rect 1690 3643 1696 3644
rect 552 3640 566 3642
rect 552 3639 553 3640
rect 547 3638 553 3639
rect 564 3638 566 3640
rect 858 3639 864 3640
rect 858 3638 859 3639
rect 564 3636 859 3638
rect 858 3635 859 3636
rect 863 3635 864 3639
rect 1690 3639 1691 3643
rect 1695 3642 1696 3643
rect 1707 3643 1713 3644
rect 1707 3642 1708 3643
rect 1695 3640 1708 3642
rect 1695 3639 1696 3640
rect 1690 3638 1696 3639
rect 1707 3639 1708 3640
rect 1712 3639 1713 3643
rect 1707 3638 1713 3639
rect 858 3634 864 3635
rect 410 3623 416 3624
rect 387 3621 393 3622
rect 387 3617 388 3621
rect 392 3617 393 3621
rect 410 3619 411 3623
rect 415 3622 416 3623
rect 515 3623 521 3624
rect 515 3622 516 3623
rect 415 3620 516 3622
rect 415 3619 416 3620
rect 410 3618 416 3619
rect 515 3619 516 3620
rect 520 3619 521 3623
rect 515 3618 521 3619
rect 538 3623 544 3624
rect 538 3619 539 3623
rect 543 3622 544 3623
rect 659 3623 665 3624
rect 659 3622 660 3623
rect 543 3620 660 3622
rect 543 3619 544 3620
rect 538 3618 544 3619
rect 659 3619 660 3620
rect 664 3619 665 3623
rect 659 3618 665 3619
rect 727 3623 733 3624
rect 727 3619 728 3623
rect 732 3622 733 3623
rect 811 3623 817 3624
rect 811 3622 812 3623
rect 732 3620 812 3622
rect 732 3619 733 3620
rect 727 3618 733 3619
rect 811 3619 812 3620
rect 816 3619 817 3623
rect 811 3618 817 3619
rect 834 3623 840 3624
rect 834 3619 835 3623
rect 839 3622 840 3623
rect 979 3623 985 3624
rect 979 3622 980 3623
rect 839 3620 980 3622
rect 839 3619 840 3620
rect 834 3618 840 3619
rect 979 3619 980 3620
rect 984 3619 985 3623
rect 979 3618 985 3619
rect 1114 3623 1120 3624
rect 1114 3619 1115 3623
rect 1119 3622 1120 3623
rect 1147 3623 1153 3624
rect 1147 3622 1148 3623
rect 1119 3620 1148 3622
rect 1119 3619 1120 3620
rect 1114 3618 1120 3619
rect 1147 3619 1148 3620
rect 1152 3619 1153 3623
rect 1147 3618 1153 3619
rect 1170 3623 1176 3624
rect 1170 3619 1171 3623
rect 1175 3622 1176 3623
rect 1315 3623 1321 3624
rect 1315 3622 1316 3623
rect 1175 3620 1316 3622
rect 1175 3619 1176 3620
rect 1170 3618 1176 3619
rect 1315 3619 1316 3620
rect 1320 3619 1321 3623
rect 1514 3623 1520 3624
rect 1315 3618 1321 3619
rect 1491 3621 1497 3622
rect 387 3616 393 3617
rect 1491 3617 1492 3621
rect 1496 3617 1497 3621
rect 1514 3619 1515 3623
rect 1519 3622 1520 3623
rect 1667 3623 1673 3624
rect 1667 3622 1668 3623
rect 1519 3620 1668 3622
rect 1519 3619 1520 3620
rect 1514 3618 1520 3619
rect 1667 3619 1668 3620
rect 1672 3619 1673 3623
rect 1667 3618 1673 3619
rect 1843 3623 1852 3624
rect 1843 3619 1844 3623
rect 1851 3619 1852 3623
rect 1843 3618 1852 3619
rect 1491 3616 1497 3617
rect 388 3614 390 3616
rect 738 3615 744 3616
rect 738 3614 739 3615
rect 388 3612 739 3614
rect 738 3611 739 3612
rect 743 3611 744 3615
rect 1492 3614 1494 3616
rect 1758 3615 1764 3616
rect 1758 3614 1759 3615
rect 1492 3612 1759 3614
rect 738 3610 744 3611
rect 1758 3611 1759 3612
rect 1763 3611 1764 3615
rect 1758 3610 1764 3611
rect 334 3600 340 3601
rect 110 3597 116 3598
rect 110 3593 111 3597
rect 115 3593 116 3597
rect 334 3596 335 3600
rect 339 3596 340 3600
rect 334 3595 340 3596
rect 462 3600 468 3601
rect 462 3596 463 3600
rect 467 3596 468 3600
rect 462 3595 468 3596
rect 606 3600 612 3601
rect 606 3596 607 3600
rect 611 3596 612 3600
rect 606 3595 612 3596
rect 758 3600 764 3601
rect 758 3596 759 3600
rect 763 3596 764 3600
rect 758 3595 764 3596
rect 926 3600 932 3601
rect 926 3596 927 3600
rect 931 3596 932 3600
rect 926 3595 932 3596
rect 1094 3600 1100 3601
rect 1094 3596 1095 3600
rect 1099 3596 1100 3600
rect 1094 3595 1100 3596
rect 1262 3600 1268 3601
rect 1262 3596 1263 3600
rect 1267 3596 1268 3600
rect 1262 3595 1268 3596
rect 1438 3600 1444 3601
rect 1438 3596 1439 3600
rect 1443 3596 1444 3600
rect 1438 3595 1444 3596
rect 1614 3600 1620 3601
rect 1614 3596 1615 3600
rect 1619 3596 1620 3600
rect 1614 3595 1620 3596
rect 1790 3600 1796 3601
rect 1790 3596 1791 3600
rect 1795 3596 1796 3600
rect 1790 3595 1796 3596
rect 2006 3597 2012 3598
rect 110 3592 116 3593
rect 2006 3593 2007 3597
rect 2011 3593 2012 3597
rect 2006 3592 2012 3593
rect 2046 3592 2052 3593
rect 3942 3592 3948 3593
rect 410 3591 416 3592
rect 410 3587 411 3591
rect 415 3587 416 3591
rect 410 3586 416 3587
rect 538 3591 544 3592
rect 538 3587 539 3591
rect 543 3587 544 3591
rect 727 3591 733 3592
rect 727 3590 728 3591
rect 685 3588 728 3590
rect 538 3586 544 3587
rect 727 3587 728 3588
rect 732 3587 733 3591
rect 727 3586 733 3587
rect 834 3591 840 3592
rect 834 3587 835 3591
rect 839 3587 840 3591
rect 834 3586 840 3587
rect 858 3591 864 3592
rect 858 3587 859 3591
rect 863 3590 864 3591
rect 1170 3591 1176 3592
rect 863 3588 969 3590
rect 863 3587 864 3588
rect 858 3586 864 3587
rect 1170 3587 1171 3591
rect 1175 3587 1176 3591
rect 1170 3586 1176 3587
rect 1338 3591 1344 3592
rect 1338 3587 1339 3591
rect 1343 3587 1344 3591
rect 1338 3586 1344 3587
rect 1514 3591 1520 3592
rect 1514 3587 1515 3591
rect 1519 3587 1520 3591
rect 1514 3586 1520 3587
rect 1690 3591 1696 3592
rect 1690 3587 1691 3591
rect 1695 3587 1696 3591
rect 1690 3586 1696 3587
rect 1758 3591 1764 3592
rect 1758 3587 1759 3591
rect 1763 3590 1764 3591
rect 1763 3588 1833 3590
rect 2046 3588 2047 3592
rect 2051 3588 2052 3592
rect 1763 3587 1764 3588
rect 2046 3587 2052 3588
rect 2190 3591 2196 3592
rect 2190 3587 2191 3591
rect 2195 3587 2196 3591
rect 1758 3586 1764 3587
rect 2190 3586 2196 3587
rect 2326 3591 2332 3592
rect 2326 3587 2327 3591
rect 2331 3587 2332 3591
rect 2326 3586 2332 3587
rect 2454 3591 2460 3592
rect 2454 3587 2455 3591
rect 2459 3587 2460 3591
rect 2454 3586 2460 3587
rect 2582 3591 2588 3592
rect 2582 3587 2583 3591
rect 2587 3587 2588 3591
rect 2582 3586 2588 3587
rect 2718 3591 2724 3592
rect 2718 3587 2719 3591
rect 2723 3587 2724 3591
rect 2718 3586 2724 3587
rect 2854 3591 2860 3592
rect 2854 3587 2855 3591
rect 2859 3587 2860 3591
rect 2854 3586 2860 3587
rect 2998 3591 3004 3592
rect 2998 3587 2999 3591
rect 3003 3587 3004 3591
rect 2998 3586 3004 3587
rect 3142 3591 3148 3592
rect 3142 3587 3143 3591
rect 3147 3587 3148 3591
rect 3142 3586 3148 3587
rect 3294 3591 3300 3592
rect 3294 3587 3295 3591
rect 3299 3587 3300 3591
rect 3294 3586 3300 3587
rect 3454 3591 3460 3592
rect 3454 3587 3455 3591
rect 3459 3587 3460 3591
rect 3454 3586 3460 3587
rect 3622 3591 3628 3592
rect 3622 3587 3623 3591
rect 3627 3587 3628 3591
rect 3942 3588 3943 3592
rect 3947 3588 3948 3592
rect 3942 3587 3948 3588
rect 3622 3586 3628 3587
rect 3258 3583 3264 3584
rect 334 3581 340 3582
rect 110 3580 116 3581
rect 110 3576 111 3580
rect 115 3576 116 3580
rect 334 3577 335 3581
rect 339 3577 340 3581
rect 334 3576 340 3577
rect 462 3581 468 3582
rect 462 3577 463 3581
rect 467 3577 468 3581
rect 462 3576 468 3577
rect 606 3581 612 3582
rect 606 3577 607 3581
rect 611 3577 612 3581
rect 606 3576 612 3577
rect 758 3581 764 3582
rect 758 3577 759 3581
rect 763 3577 764 3581
rect 758 3576 764 3577
rect 926 3581 932 3582
rect 926 3577 927 3581
rect 931 3577 932 3581
rect 926 3576 932 3577
rect 1094 3581 1100 3582
rect 1094 3577 1095 3581
rect 1099 3577 1100 3581
rect 1094 3576 1100 3577
rect 1262 3581 1268 3582
rect 1262 3577 1263 3581
rect 1267 3577 1268 3581
rect 1262 3576 1268 3577
rect 1438 3581 1444 3582
rect 1438 3577 1439 3581
rect 1443 3577 1444 3581
rect 1438 3576 1444 3577
rect 1614 3581 1620 3582
rect 1614 3577 1615 3581
rect 1619 3577 1620 3581
rect 1614 3576 1620 3577
rect 1790 3581 1796 3582
rect 1790 3577 1791 3581
rect 1795 3577 1796 3581
rect 1790 3576 1796 3577
rect 2006 3580 2012 3581
rect 2006 3576 2007 3580
rect 2011 3576 2012 3580
rect 2278 3579 2284 3580
rect 2278 3578 2279 3579
rect 2269 3576 2279 3578
rect 110 3575 116 3576
rect 2006 3575 2012 3576
rect 2046 3575 2052 3576
rect 2046 3571 2047 3575
rect 2051 3571 2052 3575
rect 2278 3575 2279 3576
rect 2283 3575 2284 3579
rect 2439 3579 2445 3580
rect 2439 3578 2440 3579
rect 2405 3576 2440 3578
rect 2278 3574 2284 3575
rect 2439 3575 2440 3576
rect 2444 3575 2445 3579
rect 2439 3574 2445 3575
rect 2530 3579 2536 3580
rect 2530 3575 2531 3579
rect 2535 3575 2536 3579
rect 2530 3574 2536 3575
rect 2658 3579 2664 3580
rect 2658 3575 2659 3579
rect 2663 3575 2664 3579
rect 2658 3574 2664 3575
rect 2794 3579 2800 3580
rect 2794 3575 2795 3579
rect 2799 3575 2800 3579
rect 2794 3574 2800 3575
rect 2930 3579 2936 3580
rect 2930 3575 2931 3579
rect 2935 3575 2936 3579
rect 2930 3574 2936 3575
rect 3074 3579 3080 3580
rect 3074 3575 3075 3579
rect 3079 3575 3080 3579
rect 3074 3574 3080 3575
rect 3218 3579 3224 3580
rect 3218 3575 3219 3579
rect 3223 3575 3224 3579
rect 3258 3579 3259 3583
rect 3263 3582 3264 3583
rect 3378 3583 3384 3584
rect 3263 3580 3337 3582
rect 3263 3579 3264 3580
rect 3258 3578 3264 3579
rect 3378 3579 3379 3583
rect 3383 3582 3384 3583
rect 3586 3583 3592 3584
rect 3383 3580 3497 3582
rect 3383 3579 3384 3580
rect 3378 3578 3384 3579
rect 3586 3579 3587 3583
rect 3591 3582 3592 3583
rect 3591 3580 3665 3582
rect 3591 3579 3592 3580
rect 3586 3578 3592 3579
rect 3218 3574 3224 3575
rect 3942 3575 3948 3576
rect 2046 3570 2052 3571
rect 2190 3572 2196 3573
rect 2190 3568 2191 3572
rect 2195 3568 2196 3572
rect 2190 3567 2196 3568
rect 2326 3572 2332 3573
rect 2326 3568 2327 3572
rect 2331 3568 2332 3572
rect 2326 3567 2332 3568
rect 2454 3572 2460 3573
rect 2454 3568 2455 3572
rect 2459 3568 2460 3572
rect 2454 3567 2460 3568
rect 2582 3572 2588 3573
rect 2582 3568 2583 3572
rect 2587 3568 2588 3572
rect 2582 3567 2588 3568
rect 2718 3572 2724 3573
rect 2718 3568 2719 3572
rect 2723 3568 2724 3572
rect 2718 3567 2724 3568
rect 2854 3572 2860 3573
rect 2854 3568 2855 3572
rect 2859 3568 2860 3572
rect 2854 3567 2860 3568
rect 2998 3572 3004 3573
rect 2998 3568 2999 3572
rect 3003 3568 3004 3572
rect 2998 3567 3004 3568
rect 3142 3572 3148 3573
rect 3142 3568 3143 3572
rect 3147 3568 3148 3572
rect 3142 3567 3148 3568
rect 3294 3572 3300 3573
rect 3294 3568 3295 3572
rect 3299 3568 3300 3572
rect 3294 3567 3300 3568
rect 3454 3572 3460 3573
rect 3454 3568 3455 3572
rect 3459 3568 3460 3572
rect 3454 3567 3460 3568
rect 3622 3572 3628 3573
rect 3622 3568 3623 3572
rect 3627 3568 3628 3572
rect 3942 3571 3943 3575
rect 3947 3571 3948 3575
rect 3942 3570 3948 3571
rect 3622 3567 3628 3568
rect 2202 3551 2208 3552
rect 2202 3547 2203 3551
rect 2207 3550 2208 3551
rect 2243 3551 2249 3552
rect 2243 3550 2244 3551
rect 2207 3548 2244 3550
rect 2207 3547 2208 3548
rect 2202 3546 2208 3547
rect 2243 3547 2244 3548
rect 2248 3547 2249 3551
rect 2439 3551 2445 3552
rect 2243 3546 2249 3547
rect 2379 3547 2385 3548
rect 2379 3543 2380 3547
rect 2384 3546 2385 3547
rect 2431 3547 2437 3548
rect 2431 3546 2432 3547
rect 2384 3544 2432 3546
rect 2384 3543 2385 3544
rect 2379 3542 2385 3543
rect 2431 3543 2432 3544
rect 2436 3543 2437 3547
rect 2439 3547 2440 3551
rect 2444 3550 2445 3551
rect 2507 3551 2513 3552
rect 2507 3550 2508 3551
rect 2444 3548 2508 3550
rect 2444 3547 2445 3548
rect 2439 3546 2445 3547
rect 2507 3547 2508 3548
rect 2512 3547 2513 3551
rect 2507 3546 2513 3547
rect 2530 3551 2536 3552
rect 2530 3547 2531 3551
rect 2535 3550 2536 3551
rect 2635 3551 2641 3552
rect 2635 3550 2636 3551
rect 2535 3548 2636 3550
rect 2535 3547 2536 3548
rect 2530 3546 2536 3547
rect 2635 3547 2636 3548
rect 2640 3547 2641 3551
rect 2635 3546 2641 3547
rect 2658 3551 2664 3552
rect 2658 3547 2659 3551
rect 2663 3550 2664 3551
rect 2771 3551 2777 3552
rect 2771 3550 2772 3551
rect 2663 3548 2772 3550
rect 2663 3547 2664 3548
rect 2658 3546 2664 3547
rect 2771 3547 2772 3548
rect 2776 3547 2777 3551
rect 2771 3546 2777 3547
rect 2794 3551 2800 3552
rect 2794 3547 2795 3551
rect 2799 3550 2800 3551
rect 2907 3551 2913 3552
rect 2907 3550 2908 3551
rect 2799 3548 2908 3550
rect 2799 3547 2800 3548
rect 2794 3546 2800 3547
rect 2907 3547 2908 3548
rect 2912 3547 2913 3551
rect 2907 3546 2913 3547
rect 2930 3551 2936 3552
rect 2930 3547 2931 3551
rect 2935 3550 2936 3551
rect 3051 3551 3057 3552
rect 3051 3550 3052 3551
rect 2935 3548 3052 3550
rect 2935 3547 2936 3548
rect 2930 3546 2936 3547
rect 3051 3547 3052 3548
rect 3056 3547 3057 3551
rect 3051 3546 3057 3547
rect 3074 3551 3080 3552
rect 3074 3547 3075 3551
rect 3079 3550 3080 3551
rect 3195 3551 3201 3552
rect 3195 3550 3196 3551
rect 3079 3548 3196 3550
rect 3079 3547 3080 3548
rect 3074 3546 3080 3547
rect 3195 3547 3196 3548
rect 3200 3547 3201 3551
rect 3195 3546 3201 3547
rect 3218 3551 3224 3552
rect 3218 3547 3219 3551
rect 3223 3550 3224 3551
rect 3347 3551 3353 3552
rect 3347 3550 3348 3551
rect 3223 3548 3348 3550
rect 3223 3547 3224 3548
rect 3218 3546 3224 3547
rect 3347 3547 3348 3548
rect 3352 3547 3353 3551
rect 3347 3546 3353 3547
rect 3507 3551 3513 3552
rect 3507 3547 3508 3551
rect 3512 3550 3513 3551
rect 3586 3551 3592 3552
rect 3586 3550 3587 3551
rect 3512 3548 3587 3550
rect 3512 3547 3513 3548
rect 3507 3546 3513 3547
rect 3586 3547 3587 3548
rect 3591 3547 3592 3551
rect 3586 3546 3592 3547
rect 3594 3547 3600 3548
rect 2431 3542 2437 3543
rect 3258 3543 3264 3544
rect 3258 3542 3259 3543
rect 3052 3540 3259 3542
rect 3052 3538 3054 3540
rect 3258 3539 3259 3540
rect 3263 3539 3264 3543
rect 3594 3543 3595 3547
rect 3599 3546 3600 3547
rect 3675 3547 3681 3548
rect 3675 3546 3676 3547
rect 3599 3544 3676 3546
rect 3599 3543 3600 3544
rect 3594 3542 3600 3543
rect 3675 3543 3676 3544
rect 3680 3543 3681 3547
rect 3675 3542 3681 3543
rect 3258 3538 3264 3539
rect 3051 3537 3057 3538
rect 2155 3535 2161 3536
rect 2155 3531 2156 3535
rect 2160 3534 2161 3535
rect 2191 3535 2197 3536
rect 2191 3534 2192 3535
rect 2160 3532 2192 3534
rect 2160 3531 2161 3532
rect 2155 3530 2161 3531
rect 2191 3531 2192 3532
rect 2196 3531 2197 3535
rect 2191 3530 2197 3531
rect 2278 3535 2284 3536
rect 2278 3531 2279 3535
rect 2283 3534 2284 3535
rect 2323 3535 2329 3536
rect 2323 3534 2324 3535
rect 2283 3532 2324 3534
rect 2283 3531 2284 3532
rect 2278 3530 2284 3531
rect 2323 3531 2324 3532
rect 2328 3531 2329 3535
rect 2323 3530 2329 3531
rect 2499 3535 2505 3536
rect 2499 3531 2500 3535
rect 2504 3534 2505 3535
rect 2530 3535 2536 3536
rect 2530 3534 2531 3535
rect 2504 3532 2531 3534
rect 2504 3531 2505 3532
rect 2499 3530 2505 3531
rect 2530 3531 2531 3532
rect 2535 3531 2536 3535
rect 2530 3530 2536 3531
rect 2683 3535 2689 3536
rect 2683 3531 2684 3535
rect 2688 3534 2689 3535
rect 2759 3535 2765 3536
rect 2759 3534 2760 3535
rect 2688 3532 2760 3534
rect 2688 3531 2689 3532
rect 2683 3530 2689 3531
rect 2759 3531 2760 3532
rect 2764 3531 2765 3535
rect 2759 3530 2765 3531
rect 2778 3535 2784 3536
rect 2778 3531 2779 3535
rect 2783 3534 2784 3535
rect 2867 3535 2873 3536
rect 2867 3534 2868 3535
rect 2783 3532 2868 3534
rect 2783 3531 2784 3532
rect 2778 3530 2784 3531
rect 2867 3531 2868 3532
rect 2872 3531 2873 3535
rect 3051 3533 3052 3537
rect 3056 3533 3057 3537
rect 3051 3532 3057 3533
rect 3074 3535 3080 3536
rect 2867 3530 2873 3531
rect 3074 3531 3075 3535
rect 3079 3534 3080 3535
rect 3227 3535 3233 3536
rect 3227 3534 3228 3535
rect 3079 3532 3228 3534
rect 3079 3531 3080 3532
rect 3074 3530 3080 3531
rect 3227 3531 3228 3532
rect 3232 3531 3233 3535
rect 3227 3530 3233 3531
rect 3398 3535 3409 3536
rect 3398 3531 3399 3535
rect 3403 3531 3404 3535
rect 3408 3531 3409 3535
rect 3398 3530 3409 3531
rect 3426 3535 3432 3536
rect 3426 3531 3427 3535
rect 3431 3534 3432 3535
rect 3571 3535 3577 3536
rect 3571 3534 3572 3535
rect 3431 3532 3572 3534
rect 3431 3531 3432 3532
rect 3426 3530 3432 3531
rect 3571 3531 3572 3532
rect 3576 3531 3577 3535
rect 3571 3530 3577 3531
rect 3739 3535 3745 3536
rect 3739 3531 3740 3535
rect 3744 3534 3745 3535
rect 3770 3535 3776 3536
rect 3770 3534 3771 3535
rect 3744 3532 3771 3534
rect 3744 3531 3745 3532
rect 3739 3530 3745 3531
rect 3770 3531 3771 3532
rect 3775 3531 3776 3535
rect 3770 3530 3776 3531
rect 3891 3535 3897 3536
rect 3891 3531 3892 3535
rect 3896 3534 3897 3535
rect 3914 3535 3920 3536
rect 3914 3534 3915 3535
rect 3896 3532 3915 3534
rect 3896 3531 3897 3532
rect 3891 3530 3897 3531
rect 3914 3531 3915 3532
rect 3919 3531 3920 3535
rect 3914 3530 3920 3531
rect 110 3516 116 3517
rect 2006 3516 2012 3517
rect 110 3512 111 3516
rect 115 3512 116 3516
rect 110 3511 116 3512
rect 158 3515 164 3516
rect 158 3511 159 3515
rect 163 3511 164 3515
rect 158 3510 164 3511
rect 302 3515 308 3516
rect 302 3511 303 3515
rect 307 3511 308 3515
rect 302 3510 308 3511
rect 462 3515 468 3516
rect 462 3511 463 3515
rect 467 3511 468 3515
rect 462 3510 468 3511
rect 638 3515 644 3516
rect 638 3511 639 3515
rect 643 3511 644 3515
rect 638 3510 644 3511
rect 814 3515 820 3516
rect 814 3511 815 3515
rect 819 3511 820 3515
rect 814 3510 820 3511
rect 998 3515 1004 3516
rect 998 3511 999 3515
rect 1003 3511 1004 3515
rect 998 3510 1004 3511
rect 1174 3515 1180 3516
rect 1174 3511 1175 3515
rect 1179 3511 1180 3515
rect 1174 3510 1180 3511
rect 1350 3515 1356 3516
rect 1350 3511 1351 3515
rect 1355 3511 1356 3515
rect 1350 3510 1356 3511
rect 1526 3515 1532 3516
rect 1526 3511 1527 3515
rect 1531 3511 1532 3515
rect 1526 3510 1532 3511
rect 1702 3515 1708 3516
rect 1702 3511 1703 3515
rect 1707 3511 1708 3515
rect 1702 3510 1708 3511
rect 1878 3515 1884 3516
rect 1878 3511 1879 3515
rect 1883 3511 1884 3515
rect 2006 3512 2007 3516
rect 2011 3512 2012 3516
rect 2006 3511 2012 3512
rect 2102 3512 2108 3513
rect 1878 3510 1884 3511
rect 2046 3509 2052 3510
rect 738 3507 744 3508
rect 234 3503 240 3504
rect 110 3499 116 3500
rect 110 3495 111 3499
rect 115 3495 116 3499
rect 234 3499 235 3503
rect 239 3499 240 3503
rect 234 3498 240 3499
rect 378 3503 384 3504
rect 378 3499 379 3503
rect 383 3499 384 3503
rect 378 3498 384 3499
rect 538 3503 544 3504
rect 538 3499 539 3503
rect 543 3499 544 3503
rect 538 3498 544 3499
rect 714 3503 720 3504
rect 714 3499 715 3503
rect 719 3499 720 3503
rect 738 3503 739 3507
rect 743 3506 744 3507
rect 1082 3507 1088 3508
rect 743 3504 857 3506
rect 743 3503 744 3504
rect 738 3502 744 3503
rect 1074 3503 1080 3504
rect 714 3498 720 3499
rect 1074 3499 1075 3503
rect 1079 3499 1080 3503
rect 1082 3503 1083 3507
rect 1087 3506 1088 3507
rect 1311 3507 1317 3508
rect 1087 3504 1217 3506
rect 1087 3503 1088 3504
rect 1082 3502 1088 3503
rect 1311 3503 1312 3507
rect 1316 3506 1317 3507
rect 1846 3507 1852 3508
rect 1316 3504 1393 3506
rect 1316 3503 1317 3504
rect 1311 3502 1317 3503
rect 1662 3503 1668 3504
rect 1662 3502 1663 3503
rect 1605 3500 1663 3502
rect 1074 3498 1080 3499
rect 1662 3499 1663 3500
rect 1667 3499 1668 3503
rect 1662 3498 1668 3499
rect 1778 3503 1784 3504
rect 1778 3499 1779 3503
rect 1783 3499 1784 3503
rect 1846 3503 1847 3507
rect 1851 3506 1852 3507
rect 1851 3504 1921 3506
rect 2046 3505 2047 3509
rect 2051 3505 2052 3509
rect 2102 3508 2103 3512
rect 2107 3508 2108 3512
rect 2102 3507 2108 3508
rect 2270 3512 2276 3513
rect 2270 3508 2271 3512
rect 2275 3508 2276 3512
rect 2270 3507 2276 3508
rect 2446 3512 2452 3513
rect 2446 3508 2447 3512
rect 2451 3508 2452 3512
rect 2446 3507 2452 3508
rect 2630 3512 2636 3513
rect 2630 3508 2631 3512
rect 2635 3508 2636 3512
rect 2630 3507 2636 3508
rect 2814 3512 2820 3513
rect 2814 3508 2815 3512
rect 2819 3508 2820 3512
rect 2814 3507 2820 3508
rect 2998 3512 3004 3513
rect 2998 3508 2999 3512
rect 3003 3508 3004 3512
rect 2998 3507 3004 3508
rect 3174 3512 3180 3513
rect 3174 3508 3175 3512
rect 3179 3508 3180 3512
rect 3174 3507 3180 3508
rect 3350 3512 3356 3513
rect 3350 3508 3351 3512
rect 3355 3508 3356 3512
rect 3350 3507 3356 3508
rect 3518 3512 3524 3513
rect 3518 3508 3519 3512
rect 3523 3508 3524 3512
rect 3518 3507 3524 3508
rect 3686 3512 3692 3513
rect 3686 3508 3687 3512
rect 3691 3508 3692 3512
rect 3686 3507 3692 3508
rect 3838 3512 3844 3513
rect 3838 3508 3839 3512
rect 3843 3508 3844 3512
rect 3838 3507 3844 3508
rect 3942 3509 3948 3510
rect 2046 3504 2052 3505
rect 3942 3505 3943 3509
rect 3947 3505 3948 3509
rect 3942 3504 3948 3505
rect 1851 3503 1852 3504
rect 1846 3502 1852 3503
rect 2178 3503 2184 3504
rect 1778 3498 1784 3499
rect 2006 3499 2012 3500
rect 110 3494 116 3495
rect 158 3496 164 3497
rect 158 3492 159 3496
rect 163 3492 164 3496
rect 158 3491 164 3492
rect 302 3496 308 3497
rect 302 3492 303 3496
rect 307 3492 308 3496
rect 302 3491 308 3492
rect 462 3496 468 3497
rect 462 3492 463 3496
rect 467 3492 468 3496
rect 462 3491 468 3492
rect 638 3496 644 3497
rect 638 3492 639 3496
rect 643 3492 644 3496
rect 638 3491 644 3492
rect 814 3496 820 3497
rect 814 3492 815 3496
rect 819 3492 820 3496
rect 814 3491 820 3492
rect 998 3496 1004 3497
rect 998 3492 999 3496
rect 1003 3492 1004 3496
rect 998 3491 1004 3492
rect 1174 3496 1180 3497
rect 1174 3492 1175 3496
rect 1179 3492 1180 3496
rect 1174 3491 1180 3492
rect 1350 3496 1356 3497
rect 1350 3492 1351 3496
rect 1355 3492 1356 3496
rect 1350 3491 1356 3492
rect 1526 3496 1532 3497
rect 1526 3492 1527 3496
rect 1531 3492 1532 3496
rect 1526 3491 1532 3492
rect 1702 3496 1708 3497
rect 1702 3492 1703 3496
rect 1707 3492 1708 3496
rect 1702 3491 1708 3492
rect 1878 3496 1884 3497
rect 1878 3492 1879 3496
rect 1883 3492 1884 3496
rect 2006 3495 2007 3499
rect 2011 3495 2012 3499
rect 2178 3499 2179 3503
rect 2183 3499 2184 3503
rect 2178 3498 2184 3499
rect 2191 3503 2197 3504
rect 2191 3499 2192 3503
rect 2196 3502 2197 3503
rect 2431 3503 2437 3504
rect 2196 3500 2313 3502
rect 2196 3499 2197 3500
rect 2191 3498 2197 3499
rect 2431 3499 2432 3503
rect 2436 3502 2437 3503
rect 2530 3503 2536 3504
rect 2436 3500 2489 3502
rect 2436 3499 2437 3500
rect 2431 3498 2437 3499
rect 2530 3499 2531 3503
rect 2535 3502 2536 3503
rect 2759 3503 2765 3504
rect 2535 3500 2673 3502
rect 2535 3499 2536 3500
rect 2530 3498 2536 3499
rect 2759 3499 2760 3503
rect 2764 3502 2765 3503
rect 3074 3503 3080 3504
rect 2764 3500 2857 3502
rect 2764 3499 2765 3500
rect 2759 3498 2765 3499
rect 3074 3499 3075 3503
rect 3079 3499 3080 3503
rect 3074 3498 3080 3499
rect 3250 3503 3256 3504
rect 3250 3499 3251 3503
rect 3255 3499 3256 3503
rect 3250 3498 3256 3499
rect 3426 3503 3432 3504
rect 3426 3499 3427 3503
rect 3431 3499 3432 3503
rect 3426 3498 3432 3499
rect 3594 3503 3600 3504
rect 3594 3499 3595 3503
rect 3599 3499 3600 3503
rect 3594 3498 3600 3499
rect 3770 3503 3776 3504
rect 3770 3499 3771 3503
rect 3775 3502 3776 3503
rect 3775 3500 3881 3502
rect 3775 3499 3776 3500
rect 3770 3498 3776 3499
rect 2006 3494 2012 3495
rect 2102 3493 2108 3494
rect 1878 3491 1884 3492
rect 2046 3492 2052 3493
rect 2046 3488 2047 3492
rect 2051 3488 2052 3492
rect 2102 3489 2103 3493
rect 2107 3489 2108 3493
rect 2102 3488 2108 3489
rect 2270 3493 2276 3494
rect 2270 3489 2271 3493
rect 2275 3489 2276 3493
rect 2270 3488 2276 3489
rect 2446 3493 2452 3494
rect 2446 3489 2447 3493
rect 2451 3489 2452 3493
rect 2446 3488 2452 3489
rect 2630 3493 2636 3494
rect 2630 3489 2631 3493
rect 2635 3489 2636 3493
rect 2630 3488 2636 3489
rect 2814 3493 2820 3494
rect 2814 3489 2815 3493
rect 2819 3489 2820 3493
rect 2814 3488 2820 3489
rect 2998 3493 3004 3494
rect 2998 3489 2999 3493
rect 3003 3489 3004 3493
rect 2998 3488 3004 3489
rect 3174 3493 3180 3494
rect 3174 3489 3175 3493
rect 3179 3489 3180 3493
rect 3174 3488 3180 3489
rect 3350 3493 3356 3494
rect 3350 3489 3351 3493
rect 3355 3489 3356 3493
rect 3350 3488 3356 3489
rect 3518 3493 3524 3494
rect 3518 3489 3519 3493
rect 3523 3489 3524 3493
rect 3518 3488 3524 3489
rect 3686 3493 3692 3494
rect 3686 3489 3687 3493
rect 3691 3489 3692 3493
rect 3686 3488 3692 3489
rect 3838 3493 3844 3494
rect 3838 3489 3839 3493
rect 3843 3489 3844 3493
rect 3838 3488 3844 3489
rect 3942 3492 3948 3493
rect 3942 3488 3943 3492
rect 3947 3488 3948 3492
rect 2046 3487 2052 3488
rect 3942 3487 3948 3488
rect 234 3479 240 3480
rect 234 3475 235 3479
rect 239 3478 240 3479
rect 239 3476 321 3478
rect 239 3475 240 3476
rect 234 3474 240 3475
rect 319 3474 321 3476
rect 355 3475 361 3476
rect 355 3474 356 3475
rect 319 3472 356 3474
rect 211 3471 217 3472
rect 211 3467 212 3471
rect 216 3470 217 3471
rect 355 3471 356 3472
rect 360 3471 361 3475
rect 355 3470 361 3471
rect 378 3475 384 3476
rect 378 3471 379 3475
rect 383 3474 384 3475
rect 515 3475 521 3476
rect 515 3474 516 3475
rect 383 3472 516 3474
rect 383 3471 384 3472
rect 378 3470 384 3471
rect 515 3471 516 3472
rect 520 3471 521 3475
rect 515 3470 521 3471
rect 538 3475 544 3476
rect 538 3471 539 3475
rect 543 3474 544 3475
rect 691 3475 697 3476
rect 691 3474 692 3475
rect 543 3472 692 3474
rect 543 3471 544 3472
rect 538 3470 544 3471
rect 691 3471 692 3472
rect 696 3471 697 3475
rect 691 3470 697 3471
rect 714 3475 720 3476
rect 714 3471 715 3475
rect 719 3474 720 3475
rect 867 3475 873 3476
rect 867 3474 868 3475
rect 719 3472 868 3474
rect 719 3471 720 3472
rect 714 3470 720 3471
rect 867 3471 868 3472
rect 872 3471 873 3475
rect 867 3470 873 3471
rect 1051 3475 1057 3476
rect 1051 3471 1052 3475
rect 1056 3474 1057 3475
rect 1082 3475 1088 3476
rect 1082 3474 1083 3475
rect 1056 3472 1083 3474
rect 1056 3471 1057 3472
rect 1051 3470 1057 3471
rect 1082 3471 1083 3472
rect 1087 3471 1088 3475
rect 1082 3470 1088 3471
rect 1227 3475 1233 3476
rect 1227 3471 1228 3475
rect 1232 3474 1233 3475
rect 1311 3475 1317 3476
rect 1311 3474 1312 3475
rect 1232 3472 1312 3474
rect 1232 3471 1233 3472
rect 1227 3470 1233 3471
rect 1311 3471 1312 3472
rect 1316 3471 1317 3475
rect 1311 3470 1317 3471
rect 1338 3475 1344 3476
rect 1338 3471 1339 3475
rect 1343 3474 1344 3475
rect 1403 3475 1409 3476
rect 1403 3474 1404 3475
rect 1343 3472 1404 3474
rect 1343 3471 1344 3472
rect 1338 3470 1344 3471
rect 1403 3471 1404 3472
rect 1408 3471 1409 3475
rect 1662 3475 1668 3476
rect 1403 3470 1409 3471
rect 1579 3471 1585 3472
rect 216 3468 321 3470
rect 216 3467 217 3468
rect 211 3466 217 3467
rect 319 3466 321 3468
rect 678 3467 684 3468
rect 678 3466 679 3467
rect 319 3464 679 3466
rect 678 3463 679 3464
rect 683 3463 684 3467
rect 1579 3467 1580 3471
rect 1584 3470 1585 3471
rect 1602 3471 1608 3472
rect 1602 3470 1603 3471
rect 1584 3468 1603 3470
rect 1584 3467 1585 3468
rect 1579 3466 1585 3467
rect 1602 3467 1603 3468
rect 1607 3467 1608 3471
rect 1662 3471 1663 3475
rect 1667 3474 1668 3475
rect 1755 3475 1761 3476
rect 1755 3474 1756 3475
rect 1667 3472 1756 3474
rect 1667 3471 1668 3472
rect 1662 3470 1668 3471
rect 1755 3471 1756 3472
rect 1760 3471 1761 3475
rect 1755 3470 1761 3471
rect 1778 3475 1784 3476
rect 1778 3471 1779 3475
rect 1783 3474 1784 3475
rect 1931 3475 1937 3476
rect 1931 3474 1932 3475
rect 1783 3472 1932 3474
rect 1783 3471 1784 3472
rect 1778 3470 1784 3471
rect 1931 3471 1932 3472
rect 1936 3471 1937 3475
rect 1931 3470 1937 3471
rect 1602 3466 1608 3467
rect 678 3462 684 3463
rect 187 3451 193 3452
rect 187 3447 188 3451
rect 192 3450 193 3451
rect 254 3451 260 3452
rect 254 3450 255 3451
rect 192 3448 255 3450
rect 192 3447 193 3448
rect 187 3446 193 3447
rect 254 3447 255 3448
rect 259 3447 260 3451
rect 254 3446 260 3447
rect 262 3451 268 3452
rect 262 3447 263 3451
rect 267 3450 268 3451
rect 371 3451 377 3452
rect 371 3450 372 3451
rect 267 3448 372 3450
rect 267 3447 268 3448
rect 262 3446 268 3447
rect 371 3447 372 3448
rect 376 3447 377 3451
rect 371 3446 377 3447
rect 394 3451 400 3452
rect 394 3447 395 3451
rect 399 3450 400 3451
rect 587 3451 593 3452
rect 587 3450 588 3451
rect 399 3448 588 3450
rect 399 3447 400 3448
rect 394 3446 400 3447
rect 587 3447 588 3448
rect 592 3447 593 3451
rect 587 3446 593 3447
rect 610 3451 616 3452
rect 610 3447 611 3451
rect 615 3450 616 3451
rect 803 3451 809 3452
rect 803 3450 804 3451
rect 615 3448 804 3450
rect 615 3447 616 3448
rect 610 3446 616 3447
rect 803 3447 804 3448
rect 808 3447 809 3451
rect 803 3446 809 3447
rect 1011 3451 1017 3452
rect 1011 3447 1012 3451
rect 1016 3450 1017 3451
rect 1074 3451 1080 3452
rect 1074 3450 1075 3451
rect 1016 3448 1075 3450
rect 1016 3447 1017 3448
rect 1011 3446 1017 3447
rect 1074 3447 1075 3448
rect 1079 3447 1080 3451
rect 1074 3446 1080 3447
rect 1082 3451 1088 3452
rect 1082 3447 1083 3451
rect 1087 3450 1088 3451
rect 1211 3451 1217 3452
rect 1211 3450 1212 3451
rect 1087 3448 1212 3450
rect 1087 3447 1088 3448
rect 1082 3446 1088 3447
rect 1211 3447 1212 3448
rect 1216 3447 1217 3451
rect 1211 3446 1217 3447
rect 1234 3451 1240 3452
rect 1234 3447 1235 3451
rect 1239 3450 1240 3451
rect 1403 3451 1409 3452
rect 1403 3450 1404 3451
rect 1239 3448 1404 3450
rect 1239 3447 1240 3448
rect 1234 3446 1240 3447
rect 1403 3447 1404 3448
rect 1408 3447 1409 3451
rect 1403 3446 1409 3447
rect 1587 3451 1593 3452
rect 1587 3447 1588 3451
rect 1592 3450 1593 3451
rect 1618 3451 1624 3452
rect 1618 3450 1619 3451
rect 1592 3448 1619 3450
rect 1592 3447 1593 3448
rect 1587 3446 1593 3447
rect 1618 3447 1619 3448
rect 1623 3447 1624 3451
rect 1618 3446 1624 3447
rect 1771 3451 1777 3452
rect 1771 3447 1772 3451
rect 1776 3450 1777 3451
rect 1802 3451 1808 3452
rect 1802 3450 1803 3451
rect 1776 3448 1803 3450
rect 1776 3447 1777 3448
rect 1771 3446 1777 3447
rect 1802 3447 1803 3448
rect 1807 3447 1808 3451
rect 1802 3446 1808 3447
rect 1946 3451 1952 3452
rect 1946 3447 1947 3451
rect 1951 3450 1952 3451
rect 1955 3451 1961 3452
rect 1955 3450 1956 3451
rect 1951 3448 1956 3450
rect 1951 3447 1952 3448
rect 1946 3446 1952 3447
rect 1955 3447 1956 3448
rect 1960 3447 1961 3451
rect 1955 3446 1961 3447
rect 2046 3436 2052 3437
rect 3942 3436 3948 3437
rect 2046 3432 2047 3436
rect 2051 3432 2052 3436
rect 2046 3431 2052 3432
rect 2126 3435 2132 3436
rect 2126 3431 2127 3435
rect 2131 3431 2132 3435
rect 2126 3430 2132 3431
rect 2310 3435 2316 3436
rect 2310 3431 2311 3435
rect 2315 3431 2316 3435
rect 2310 3430 2316 3431
rect 2494 3435 2500 3436
rect 2494 3431 2495 3435
rect 2499 3431 2500 3435
rect 2494 3430 2500 3431
rect 2678 3435 2684 3436
rect 2678 3431 2679 3435
rect 2683 3431 2684 3435
rect 2678 3430 2684 3431
rect 2862 3435 2868 3436
rect 2862 3431 2863 3435
rect 2867 3431 2868 3435
rect 2862 3430 2868 3431
rect 3046 3435 3052 3436
rect 3046 3431 3047 3435
rect 3051 3431 3052 3435
rect 3046 3430 3052 3431
rect 3222 3435 3228 3436
rect 3222 3431 3223 3435
rect 3227 3431 3228 3435
rect 3222 3430 3228 3431
rect 3406 3435 3412 3436
rect 3406 3431 3407 3435
rect 3411 3431 3412 3435
rect 3406 3430 3412 3431
rect 3590 3435 3596 3436
rect 3590 3431 3591 3435
rect 3595 3431 3596 3435
rect 3590 3430 3596 3431
rect 3774 3435 3780 3436
rect 3774 3431 3775 3435
rect 3779 3431 3780 3435
rect 3942 3432 3943 3436
rect 3947 3432 3948 3436
rect 3942 3431 3948 3432
rect 3774 3430 3780 3431
rect 134 3428 140 3429
rect 110 3425 116 3426
rect 110 3421 111 3425
rect 115 3421 116 3425
rect 134 3424 135 3428
rect 139 3424 140 3428
rect 134 3423 140 3424
rect 318 3428 324 3429
rect 318 3424 319 3428
rect 323 3424 324 3428
rect 318 3423 324 3424
rect 534 3428 540 3429
rect 534 3424 535 3428
rect 539 3424 540 3428
rect 534 3423 540 3424
rect 750 3428 756 3429
rect 750 3424 751 3428
rect 755 3424 756 3428
rect 750 3423 756 3424
rect 958 3428 964 3429
rect 958 3424 959 3428
rect 963 3424 964 3428
rect 958 3423 964 3424
rect 1158 3428 1164 3429
rect 1158 3424 1159 3428
rect 1163 3424 1164 3428
rect 1158 3423 1164 3424
rect 1350 3428 1356 3429
rect 1350 3424 1351 3428
rect 1355 3424 1356 3428
rect 1350 3423 1356 3424
rect 1534 3428 1540 3429
rect 1534 3424 1535 3428
rect 1539 3424 1540 3428
rect 1534 3423 1540 3424
rect 1718 3428 1724 3429
rect 1718 3424 1719 3428
rect 1723 3424 1724 3428
rect 1718 3423 1724 3424
rect 1902 3428 1908 3429
rect 1902 3424 1903 3428
rect 1907 3424 1908 3428
rect 2778 3427 2784 3428
rect 2778 3426 2779 3427
rect 1902 3423 1908 3424
rect 2006 3425 2012 3426
rect 110 3420 116 3421
rect 2006 3421 2007 3425
rect 2011 3421 2012 3425
rect 2757 3424 2779 3426
rect 2006 3420 2012 3421
rect 2202 3423 2208 3424
rect 262 3419 268 3420
rect 262 3418 263 3419
rect 213 3416 263 3418
rect 262 3415 263 3416
rect 267 3415 268 3419
rect 262 3414 268 3415
rect 394 3419 400 3420
rect 394 3415 395 3419
rect 399 3415 400 3419
rect 394 3414 400 3415
rect 610 3419 616 3420
rect 610 3415 611 3419
rect 615 3415 616 3419
rect 610 3414 616 3415
rect 678 3419 684 3420
rect 678 3415 679 3419
rect 683 3418 684 3419
rect 1082 3419 1088 3420
rect 1082 3418 1083 3419
rect 683 3416 793 3418
rect 1037 3416 1083 3418
rect 683 3415 684 3416
rect 678 3414 684 3415
rect 1082 3415 1083 3416
rect 1087 3415 1088 3419
rect 1082 3414 1088 3415
rect 1234 3419 1240 3420
rect 1234 3415 1235 3419
rect 1239 3415 1240 3419
rect 1234 3414 1240 3415
rect 1426 3419 1432 3420
rect 1426 3415 1427 3419
rect 1431 3415 1432 3419
rect 1426 3414 1432 3415
rect 1602 3419 1608 3420
rect 1602 3415 1603 3419
rect 1607 3415 1608 3419
rect 1602 3414 1608 3415
rect 1618 3419 1624 3420
rect 1618 3415 1619 3419
rect 1623 3418 1624 3419
rect 1802 3419 1808 3420
rect 1623 3416 1761 3418
rect 1623 3415 1624 3416
rect 1618 3414 1624 3415
rect 1802 3415 1803 3419
rect 1807 3418 1808 3419
rect 2046 3419 2052 3420
rect 1807 3416 1945 3418
rect 1807 3415 1808 3416
rect 1802 3414 1808 3415
rect 2046 3415 2047 3419
rect 2051 3415 2052 3419
rect 2202 3419 2203 3423
rect 2207 3419 2208 3423
rect 2202 3418 2208 3419
rect 2386 3423 2392 3424
rect 2386 3419 2387 3423
rect 2391 3419 2392 3423
rect 2386 3418 2392 3419
rect 2570 3423 2576 3424
rect 2570 3419 2571 3423
rect 2575 3419 2576 3423
rect 2778 3423 2779 3424
rect 2783 3423 2784 3427
rect 2975 3427 2981 3428
rect 2778 3422 2784 3423
rect 2946 3423 2952 3424
rect 2946 3422 2947 3423
rect 2941 3420 2947 3422
rect 2570 3418 2576 3419
rect 2946 3419 2947 3420
rect 2951 3419 2952 3423
rect 2975 3423 2976 3427
rect 2980 3426 2981 3427
rect 3174 3427 3180 3428
rect 2980 3424 3089 3426
rect 2980 3423 2981 3424
rect 2975 3422 2981 3423
rect 3174 3423 3175 3427
rect 3179 3426 3180 3427
rect 3398 3427 3404 3428
rect 3179 3424 3265 3426
rect 3179 3423 3180 3424
rect 3174 3422 3180 3423
rect 3398 3423 3399 3427
rect 3403 3426 3404 3427
rect 3546 3427 3552 3428
rect 3403 3424 3449 3426
rect 3403 3423 3404 3424
rect 3398 3422 3404 3423
rect 3546 3423 3547 3427
rect 3551 3426 3552 3427
rect 3551 3424 3633 3426
rect 3551 3423 3552 3424
rect 3546 3422 3552 3423
rect 3850 3423 3856 3424
rect 2946 3418 2952 3419
rect 3850 3419 3851 3423
rect 3855 3419 3856 3423
rect 3850 3418 3856 3419
rect 3942 3419 3948 3420
rect 2046 3414 2052 3415
rect 2126 3416 2132 3417
rect 2126 3412 2127 3416
rect 2131 3412 2132 3416
rect 2126 3411 2132 3412
rect 2310 3416 2316 3417
rect 2310 3412 2311 3416
rect 2315 3412 2316 3416
rect 2310 3411 2316 3412
rect 2494 3416 2500 3417
rect 2494 3412 2495 3416
rect 2499 3412 2500 3416
rect 2494 3411 2500 3412
rect 2678 3416 2684 3417
rect 2678 3412 2679 3416
rect 2683 3412 2684 3416
rect 2678 3411 2684 3412
rect 2862 3416 2868 3417
rect 2862 3412 2863 3416
rect 2867 3412 2868 3416
rect 2862 3411 2868 3412
rect 3046 3416 3052 3417
rect 3046 3412 3047 3416
rect 3051 3412 3052 3416
rect 3046 3411 3052 3412
rect 3222 3416 3228 3417
rect 3222 3412 3223 3416
rect 3227 3412 3228 3416
rect 3222 3411 3228 3412
rect 3406 3416 3412 3417
rect 3406 3412 3407 3416
rect 3411 3412 3412 3416
rect 3406 3411 3412 3412
rect 3590 3416 3596 3417
rect 3590 3412 3591 3416
rect 3595 3412 3596 3416
rect 3590 3411 3596 3412
rect 3774 3416 3780 3417
rect 3774 3412 3775 3416
rect 3779 3412 3780 3416
rect 3942 3415 3943 3419
rect 3947 3415 3948 3419
rect 3942 3414 3948 3415
rect 3774 3411 3780 3412
rect 134 3409 140 3410
rect 110 3408 116 3409
rect 110 3404 111 3408
rect 115 3404 116 3408
rect 134 3405 135 3409
rect 139 3405 140 3409
rect 134 3404 140 3405
rect 318 3409 324 3410
rect 318 3405 319 3409
rect 323 3405 324 3409
rect 318 3404 324 3405
rect 534 3409 540 3410
rect 534 3405 535 3409
rect 539 3405 540 3409
rect 534 3404 540 3405
rect 750 3409 756 3410
rect 750 3405 751 3409
rect 755 3405 756 3409
rect 750 3404 756 3405
rect 958 3409 964 3410
rect 958 3405 959 3409
rect 963 3405 964 3409
rect 958 3404 964 3405
rect 1158 3409 1164 3410
rect 1158 3405 1159 3409
rect 1163 3405 1164 3409
rect 1158 3404 1164 3405
rect 1350 3409 1356 3410
rect 1350 3405 1351 3409
rect 1355 3405 1356 3409
rect 1350 3404 1356 3405
rect 1534 3409 1540 3410
rect 1534 3405 1535 3409
rect 1539 3405 1540 3409
rect 1534 3404 1540 3405
rect 1718 3409 1724 3410
rect 1718 3405 1719 3409
rect 1723 3405 1724 3409
rect 1718 3404 1724 3405
rect 1902 3409 1908 3410
rect 1902 3405 1903 3409
rect 1907 3405 1908 3409
rect 1902 3404 1908 3405
rect 2006 3408 2012 3409
rect 2006 3404 2007 3408
rect 2011 3404 2012 3408
rect 110 3403 116 3404
rect 2006 3403 2012 3404
rect 2178 3395 2185 3396
rect 2178 3391 2179 3395
rect 2184 3391 2185 3395
rect 2386 3395 2392 3396
rect 2178 3390 2185 3391
rect 2351 3391 2357 3392
rect 2351 3387 2352 3391
rect 2356 3390 2357 3391
rect 2363 3391 2369 3392
rect 2363 3390 2364 3391
rect 2356 3388 2364 3390
rect 2356 3387 2357 3388
rect 2351 3386 2357 3387
rect 2363 3387 2364 3388
rect 2368 3387 2369 3391
rect 2386 3391 2387 3395
rect 2391 3394 2392 3395
rect 2547 3395 2553 3396
rect 2547 3394 2548 3395
rect 2391 3392 2548 3394
rect 2391 3391 2392 3392
rect 2386 3390 2392 3391
rect 2547 3391 2548 3392
rect 2552 3391 2553 3395
rect 2547 3390 2553 3391
rect 2570 3395 2576 3396
rect 2570 3391 2571 3395
rect 2575 3394 2576 3395
rect 2731 3395 2737 3396
rect 2731 3394 2732 3395
rect 2575 3392 2732 3394
rect 2575 3391 2576 3392
rect 2570 3390 2576 3391
rect 2731 3391 2732 3392
rect 2736 3391 2737 3395
rect 2731 3390 2737 3391
rect 2915 3395 2921 3396
rect 2915 3391 2916 3395
rect 2920 3394 2921 3395
rect 2975 3395 2981 3396
rect 2975 3394 2976 3395
rect 2920 3392 2976 3394
rect 2920 3391 2921 3392
rect 2915 3390 2921 3391
rect 2975 3391 2976 3392
rect 2980 3391 2981 3395
rect 2975 3390 2981 3391
rect 3099 3395 3105 3396
rect 3099 3391 3100 3395
rect 3104 3394 3105 3395
rect 3174 3395 3180 3396
rect 3174 3394 3175 3395
rect 3104 3392 3175 3394
rect 3104 3391 3105 3392
rect 3099 3390 3105 3391
rect 3174 3391 3175 3392
rect 3179 3391 3180 3395
rect 3174 3390 3180 3391
rect 3250 3395 3256 3396
rect 3250 3391 3251 3395
rect 3255 3394 3256 3395
rect 3275 3395 3281 3396
rect 3275 3394 3276 3395
rect 3255 3392 3276 3394
rect 3255 3391 3256 3392
rect 3250 3390 3256 3391
rect 3275 3391 3276 3392
rect 3280 3391 3281 3395
rect 3275 3390 3281 3391
rect 3459 3395 3465 3396
rect 3459 3391 3460 3395
rect 3464 3394 3465 3395
rect 3546 3395 3552 3396
rect 3546 3394 3547 3395
rect 3464 3392 3547 3394
rect 3464 3391 3465 3392
rect 3459 3390 3465 3391
rect 3546 3391 3547 3392
rect 3551 3391 3552 3395
rect 3826 3395 3833 3396
rect 3546 3390 3552 3391
rect 3643 3391 3649 3392
rect 2363 3386 2369 3387
rect 3643 3387 3644 3391
rect 3648 3390 3649 3391
rect 3658 3391 3664 3392
rect 3658 3390 3659 3391
rect 3648 3388 3659 3390
rect 3648 3387 3649 3388
rect 3643 3386 3649 3387
rect 3658 3387 3659 3388
rect 3663 3387 3664 3391
rect 3826 3391 3827 3395
rect 3832 3391 3833 3395
rect 3826 3390 3833 3391
rect 3658 3386 3664 3387
rect 2123 3363 2129 3364
rect 2123 3359 2124 3363
rect 2128 3362 2129 3363
rect 2154 3363 2160 3364
rect 2154 3362 2155 3363
rect 2128 3360 2155 3362
rect 2128 3359 2129 3360
rect 2123 3358 2129 3359
rect 2154 3359 2155 3360
rect 2159 3359 2160 3363
rect 2154 3358 2160 3359
rect 2202 3363 2208 3364
rect 2202 3359 2203 3363
rect 2207 3362 2208 3363
rect 2267 3363 2273 3364
rect 2267 3362 2268 3363
rect 2207 3360 2268 3362
rect 2207 3359 2208 3360
rect 2202 3358 2208 3359
rect 2267 3359 2268 3360
rect 2272 3359 2273 3363
rect 2267 3358 2273 3359
rect 2411 3363 2417 3364
rect 2411 3359 2412 3363
rect 2416 3362 2417 3363
rect 2442 3363 2448 3364
rect 2442 3362 2443 3363
rect 2416 3360 2443 3362
rect 2416 3359 2417 3360
rect 2411 3358 2417 3359
rect 2442 3359 2443 3360
rect 2447 3359 2448 3363
rect 2442 3358 2448 3359
rect 2563 3363 2569 3364
rect 2563 3359 2564 3363
rect 2568 3362 2569 3363
rect 2594 3363 2600 3364
rect 2594 3362 2595 3363
rect 2568 3360 2595 3362
rect 2568 3359 2569 3360
rect 2563 3358 2569 3359
rect 2594 3359 2595 3360
rect 2599 3359 2600 3363
rect 2594 3358 2600 3359
rect 2707 3363 2713 3364
rect 2707 3359 2708 3363
rect 2712 3362 2713 3363
rect 2774 3363 2780 3364
rect 2774 3362 2775 3363
rect 2712 3360 2775 3362
rect 2712 3359 2713 3360
rect 2707 3358 2713 3359
rect 2774 3359 2775 3360
rect 2779 3359 2780 3363
rect 2774 3358 2780 3359
rect 2851 3363 2857 3364
rect 2851 3359 2852 3363
rect 2856 3362 2857 3363
rect 2870 3363 2876 3364
rect 2870 3362 2871 3363
rect 2856 3360 2871 3362
rect 2856 3359 2857 3360
rect 2851 3358 2857 3359
rect 2870 3359 2871 3360
rect 2875 3359 2876 3363
rect 2870 3358 2876 3359
rect 2946 3363 2952 3364
rect 2946 3359 2947 3363
rect 2951 3362 2952 3363
rect 2987 3363 2993 3364
rect 2987 3362 2988 3363
rect 2951 3360 2988 3362
rect 2951 3359 2952 3360
rect 2946 3358 2952 3359
rect 2987 3359 2988 3360
rect 2992 3359 2993 3363
rect 2987 3358 2993 3359
rect 3010 3363 3016 3364
rect 3010 3359 3011 3363
rect 3015 3362 3016 3363
rect 3131 3363 3137 3364
rect 3131 3362 3132 3363
rect 3015 3360 3132 3362
rect 3015 3359 3016 3360
rect 3010 3358 3016 3359
rect 3131 3359 3132 3360
rect 3136 3359 3137 3363
rect 3131 3358 3137 3359
rect 3154 3363 3160 3364
rect 3154 3359 3155 3363
rect 3159 3362 3160 3363
rect 3275 3363 3281 3364
rect 3275 3362 3276 3363
rect 3159 3360 3276 3362
rect 3159 3359 3160 3360
rect 3154 3358 3160 3359
rect 3275 3359 3276 3360
rect 3280 3359 3281 3363
rect 3275 3358 3281 3359
rect 3427 3363 3433 3364
rect 3427 3359 3428 3363
rect 3432 3362 3433 3363
rect 3498 3363 3504 3364
rect 3498 3362 3499 3363
rect 3432 3360 3499 3362
rect 3432 3359 3433 3360
rect 3427 3358 3433 3359
rect 3498 3359 3499 3360
rect 3503 3359 3504 3363
rect 3498 3358 3504 3359
rect 3506 3363 3512 3364
rect 3506 3359 3507 3363
rect 3511 3362 3512 3363
rect 3587 3363 3593 3364
rect 3587 3362 3588 3363
rect 3511 3360 3588 3362
rect 3511 3359 3512 3360
rect 3506 3358 3512 3359
rect 3587 3359 3588 3360
rect 3592 3359 3593 3363
rect 3587 3358 3593 3359
rect 3610 3363 3616 3364
rect 3610 3359 3611 3363
rect 3615 3362 3616 3363
rect 3747 3363 3753 3364
rect 3747 3362 3748 3363
rect 3615 3360 3748 3362
rect 3615 3359 3616 3360
rect 3610 3358 3616 3359
rect 3747 3359 3748 3360
rect 3752 3359 3753 3363
rect 3747 3358 3753 3359
rect 3891 3363 3897 3364
rect 3891 3359 3892 3363
rect 3896 3362 3897 3363
rect 3906 3363 3912 3364
rect 3906 3362 3907 3363
rect 3896 3360 3907 3362
rect 3896 3359 3897 3360
rect 3891 3358 3897 3359
rect 3906 3359 3907 3360
rect 3911 3359 3912 3363
rect 3906 3358 3912 3359
rect 110 3356 116 3357
rect 2006 3356 2012 3357
rect 110 3352 111 3356
rect 115 3352 116 3356
rect 110 3351 116 3352
rect 134 3355 140 3356
rect 134 3351 135 3355
rect 139 3351 140 3355
rect 134 3350 140 3351
rect 230 3355 236 3356
rect 230 3351 231 3355
rect 235 3351 236 3355
rect 230 3350 236 3351
rect 374 3355 380 3356
rect 374 3351 375 3355
rect 379 3351 380 3355
rect 374 3350 380 3351
rect 534 3355 540 3356
rect 534 3351 535 3355
rect 539 3351 540 3355
rect 534 3350 540 3351
rect 702 3355 708 3356
rect 702 3351 703 3355
rect 707 3351 708 3355
rect 702 3350 708 3351
rect 870 3355 876 3356
rect 870 3351 871 3355
rect 875 3351 876 3355
rect 870 3350 876 3351
rect 1046 3355 1052 3356
rect 1046 3351 1047 3355
rect 1051 3351 1052 3355
rect 1046 3350 1052 3351
rect 1214 3355 1220 3356
rect 1214 3351 1215 3355
rect 1219 3351 1220 3355
rect 1214 3350 1220 3351
rect 1382 3355 1388 3356
rect 1382 3351 1383 3355
rect 1387 3351 1388 3355
rect 1382 3350 1388 3351
rect 1542 3355 1548 3356
rect 1542 3351 1543 3355
rect 1547 3351 1548 3355
rect 1542 3350 1548 3351
rect 1702 3355 1708 3356
rect 1702 3351 1703 3355
rect 1707 3351 1708 3355
rect 1702 3350 1708 3351
rect 1870 3355 1876 3356
rect 1870 3351 1871 3355
rect 1875 3351 1876 3355
rect 2006 3352 2007 3356
rect 2011 3352 2012 3356
rect 2006 3351 2012 3352
rect 1870 3350 1876 3351
rect 798 3347 804 3348
rect 210 3343 216 3344
rect 110 3339 116 3340
rect 110 3335 111 3339
rect 115 3335 116 3339
rect 210 3339 211 3343
rect 215 3339 216 3343
rect 210 3338 216 3339
rect 306 3343 312 3344
rect 306 3339 307 3343
rect 311 3339 312 3343
rect 306 3338 312 3339
rect 450 3343 456 3344
rect 450 3339 451 3343
rect 455 3339 456 3343
rect 450 3338 456 3339
rect 610 3343 616 3344
rect 610 3339 611 3343
rect 615 3339 616 3343
rect 610 3338 616 3339
rect 778 3343 784 3344
rect 778 3339 779 3343
rect 783 3339 784 3343
rect 798 3343 799 3347
rect 803 3346 804 3347
rect 1166 3347 1172 3348
rect 803 3344 913 3346
rect 803 3343 804 3344
rect 798 3342 804 3343
rect 1122 3343 1128 3344
rect 778 3338 784 3339
rect 1122 3339 1123 3343
rect 1127 3339 1128 3343
rect 1166 3343 1167 3347
rect 1171 3346 1172 3347
rect 1342 3347 1348 3348
rect 1171 3344 1257 3346
rect 1171 3343 1172 3344
rect 1166 3342 1172 3343
rect 1342 3343 1343 3347
rect 1347 3346 1348 3347
rect 1946 3347 1952 3348
rect 1347 3344 1425 3346
rect 1347 3343 1348 3344
rect 1342 3342 1348 3343
rect 1618 3343 1624 3344
rect 1122 3338 1128 3339
rect 1618 3339 1619 3343
rect 1623 3339 1624 3343
rect 1618 3338 1624 3339
rect 1778 3343 1784 3344
rect 1778 3339 1779 3343
rect 1783 3339 1784 3343
rect 1946 3343 1947 3347
rect 1951 3343 1952 3347
rect 1946 3342 1952 3343
rect 2070 3340 2076 3341
rect 1778 3338 1784 3339
rect 2006 3339 2012 3340
rect 110 3334 116 3335
rect 134 3336 140 3337
rect 134 3332 135 3336
rect 139 3332 140 3336
rect 134 3331 140 3332
rect 230 3336 236 3337
rect 230 3332 231 3336
rect 235 3332 236 3336
rect 230 3331 236 3332
rect 374 3336 380 3337
rect 374 3332 375 3336
rect 379 3332 380 3336
rect 374 3331 380 3332
rect 534 3336 540 3337
rect 534 3332 535 3336
rect 539 3332 540 3336
rect 534 3331 540 3332
rect 702 3336 708 3337
rect 702 3332 703 3336
rect 707 3332 708 3336
rect 702 3331 708 3332
rect 870 3336 876 3337
rect 870 3332 871 3336
rect 875 3332 876 3336
rect 870 3331 876 3332
rect 1046 3336 1052 3337
rect 1046 3332 1047 3336
rect 1051 3332 1052 3336
rect 1046 3331 1052 3332
rect 1214 3336 1220 3337
rect 1214 3332 1215 3336
rect 1219 3332 1220 3336
rect 1214 3331 1220 3332
rect 1382 3336 1388 3337
rect 1382 3332 1383 3336
rect 1387 3332 1388 3336
rect 1382 3331 1388 3332
rect 1542 3336 1548 3337
rect 1542 3332 1543 3336
rect 1547 3332 1548 3336
rect 1542 3331 1548 3332
rect 1702 3336 1708 3337
rect 1702 3332 1703 3336
rect 1707 3332 1708 3336
rect 1702 3331 1708 3332
rect 1870 3336 1876 3337
rect 1870 3332 1871 3336
rect 1875 3332 1876 3336
rect 2006 3335 2007 3339
rect 2011 3335 2012 3339
rect 2006 3334 2012 3335
rect 2046 3337 2052 3338
rect 2046 3333 2047 3337
rect 2051 3333 2052 3337
rect 2070 3336 2071 3340
rect 2075 3336 2076 3340
rect 2070 3335 2076 3336
rect 2214 3340 2220 3341
rect 2214 3336 2215 3340
rect 2219 3336 2220 3340
rect 2214 3335 2220 3336
rect 2358 3340 2364 3341
rect 2358 3336 2359 3340
rect 2363 3336 2364 3340
rect 2358 3335 2364 3336
rect 2510 3340 2516 3341
rect 2510 3336 2511 3340
rect 2515 3336 2516 3340
rect 2510 3335 2516 3336
rect 2654 3340 2660 3341
rect 2654 3336 2655 3340
rect 2659 3336 2660 3340
rect 2654 3335 2660 3336
rect 2798 3340 2804 3341
rect 2798 3336 2799 3340
rect 2803 3336 2804 3340
rect 2798 3335 2804 3336
rect 2934 3340 2940 3341
rect 2934 3336 2935 3340
rect 2939 3336 2940 3340
rect 2934 3335 2940 3336
rect 3078 3340 3084 3341
rect 3078 3336 3079 3340
rect 3083 3336 3084 3340
rect 3078 3335 3084 3336
rect 3222 3340 3228 3341
rect 3222 3336 3223 3340
rect 3227 3336 3228 3340
rect 3222 3335 3228 3336
rect 3374 3340 3380 3341
rect 3374 3336 3375 3340
rect 3379 3336 3380 3340
rect 3374 3335 3380 3336
rect 3534 3340 3540 3341
rect 3534 3336 3535 3340
rect 3539 3336 3540 3340
rect 3534 3335 3540 3336
rect 3694 3340 3700 3341
rect 3694 3336 3695 3340
rect 3699 3336 3700 3340
rect 3694 3335 3700 3336
rect 3838 3340 3844 3341
rect 3838 3336 3839 3340
rect 3843 3336 3844 3340
rect 3838 3335 3844 3336
rect 3942 3337 3948 3338
rect 2046 3332 2052 3333
rect 3942 3333 3943 3337
rect 3947 3333 3948 3337
rect 3942 3332 3948 3333
rect 1870 3331 1876 3332
rect 2146 3331 2152 3332
rect 2146 3327 2147 3331
rect 2151 3327 2152 3331
rect 2146 3326 2152 3327
rect 2154 3331 2160 3332
rect 2154 3327 2155 3331
rect 2159 3330 2160 3331
rect 2351 3331 2357 3332
rect 2159 3328 2257 3330
rect 2159 3327 2160 3328
rect 2154 3326 2160 3327
rect 2351 3327 2352 3331
rect 2356 3330 2357 3331
rect 2442 3331 2448 3332
rect 2356 3328 2401 3330
rect 2356 3327 2357 3328
rect 2351 3326 2357 3327
rect 2442 3327 2443 3331
rect 2447 3330 2448 3331
rect 2594 3331 2600 3332
rect 2447 3328 2553 3330
rect 2447 3327 2448 3328
rect 2442 3326 2448 3327
rect 2594 3327 2595 3331
rect 2599 3330 2600 3331
rect 2774 3331 2780 3332
rect 2599 3328 2697 3330
rect 2599 3327 2600 3328
rect 2594 3326 2600 3327
rect 2774 3327 2775 3331
rect 2779 3330 2780 3331
rect 3010 3331 3016 3332
rect 2779 3328 2841 3330
rect 2779 3327 2780 3328
rect 2774 3326 2780 3327
rect 3010 3327 3011 3331
rect 3015 3327 3016 3331
rect 3010 3326 3016 3327
rect 3154 3331 3160 3332
rect 3154 3327 3155 3331
rect 3159 3327 3160 3331
rect 3154 3326 3160 3327
rect 3298 3331 3304 3332
rect 3298 3327 3299 3331
rect 3303 3327 3304 3331
rect 3506 3331 3512 3332
rect 3506 3330 3507 3331
rect 3453 3328 3507 3330
rect 3298 3326 3304 3327
rect 3506 3327 3507 3328
rect 3511 3327 3512 3331
rect 3506 3326 3512 3327
rect 3610 3331 3616 3332
rect 3610 3327 3611 3331
rect 3615 3327 3616 3331
rect 3610 3326 3616 3327
rect 3658 3331 3664 3332
rect 3658 3327 3659 3331
rect 3663 3330 3664 3331
rect 3914 3331 3920 3332
rect 3663 3328 3737 3330
rect 3663 3327 3664 3328
rect 3658 3326 3664 3327
rect 3914 3327 3915 3331
rect 3919 3327 3920 3331
rect 3914 3326 3920 3327
rect 2070 3321 2076 3322
rect 2046 3320 2052 3321
rect 2046 3316 2047 3320
rect 2051 3316 2052 3320
rect 2070 3317 2071 3321
rect 2075 3317 2076 3321
rect 2070 3316 2076 3317
rect 2214 3321 2220 3322
rect 2214 3317 2215 3321
rect 2219 3317 2220 3321
rect 2214 3316 2220 3317
rect 2358 3321 2364 3322
rect 2358 3317 2359 3321
rect 2363 3317 2364 3321
rect 2358 3316 2364 3317
rect 2510 3321 2516 3322
rect 2510 3317 2511 3321
rect 2515 3317 2516 3321
rect 2510 3316 2516 3317
rect 2654 3321 2660 3322
rect 2654 3317 2655 3321
rect 2659 3317 2660 3321
rect 2654 3316 2660 3317
rect 2798 3321 2804 3322
rect 2798 3317 2799 3321
rect 2803 3317 2804 3321
rect 2798 3316 2804 3317
rect 2934 3321 2940 3322
rect 2934 3317 2935 3321
rect 2939 3317 2940 3321
rect 2934 3316 2940 3317
rect 3078 3321 3084 3322
rect 3078 3317 3079 3321
rect 3083 3317 3084 3321
rect 3078 3316 3084 3317
rect 3222 3321 3228 3322
rect 3222 3317 3223 3321
rect 3227 3317 3228 3321
rect 3222 3316 3228 3317
rect 3374 3321 3380 3322
rect 3374 3317 3375 3321
rect 3379 3317 3380 3321
rect 3374 3316 3380 3317
rect 3534 3321 3540 3322
rect 3534 3317 3535 3321
rect 3539 3317 3540 3321
rect 3534 3316 3540 3317
rect 3694 3321 3700 3322
rect 3694 3317 3695 3321
rect 3699 3317 3700 3321
rect 3694 3316 3700 3317
rect 3838 3321 3844 3322
rect 3838 3317 3839 3321
rect 3843 3317 3844 3321
rect 3838 3316 3844 3317
rect 3942 3320 3948 3321
rect 3942 3316 3943 3320
rect 3947 3316 3948 3320
rect 210 3315 216 3316
rect 187 3311 193 3312
rect 187 3307 188 3311
rect 192 3310 193 3311
rect 202 3311 208 3312
rect 202 3310 203 3311
rect 192 3308 203 3310
rect 192 3307 193 3308
rect 187 3306 193 3307
rect 202 3307 203 3308
rect 207 3307 208 3311
rect 210 3311 211 3315
rect 215 3314 216 3315
rect 283 3315 289 3316
rect 283 3314 284 3315
rect 215 3312 284 3314
rect 215 3311 216 3312
rect 210 3310 216 3311
rect 283 3311 284 3312
rect 288 3311 289 3315
rect 283 3310 289 3311
rect 306 3315 312 3316
rect 306 3311 307 3315
rect 311 3314 312 3315
rect 427 3315 433 3316
rect 427 3314 428 3315
rect 311 3312 428 3314
rect 311 3311 312 3312
rect 306 3310 312 3311
rect 427 3311 428 3312
rect 432 3311 433 3315
rect 427 3310 433 3311
rect 450 3315 456 3316
rect 450 3311 451 3315
rect 455 3314 456 3315
rect 587 3315 593 3316
rect 587 3314 588 3315
rect 455 3312 588 3314
rect 455 3311 456 3312
rect 450 3310 456 3311
rect 587 3311 588 3312
rect 592 3311 593 3315
rect 587 3310 593 3311
rect 610 3315 616 3316
rect 610 3311 611 3315
rect 615 3314 616 3315
rect 755 3315 761 3316
rect 755 3314 756 3315
rect 615 3312 756 3314
rect 615 3311 616 3312
rect 610 3310 616 3311
rect 755 3311 756 3312
rect 760 3311 761 3315
rect 755 3310 761 3311
rect 778 3315 784 3316
rect 778 3311 779 3315
rect 783 3314 784 3315
rect 923 3315 929 3316
rect 923 3314 924 3315
rect 783 3312 924 3314
rect 783 3311 784 3312
rect 778 3310 784 3311
rect 923 3311 924 3312
rect 928 3311 929 3315
rect 923 3310 929 3311
rect 1099 3315 1105 3316
rect 1099 3311 1100 3315
rect 1104 3314 1105 3315
rect 1166 3315 1172 3316
rect 1166 3314 1167 3315
rect 1104 3312 1167 3314
rect 1104 3311 1105 3312
rect 1099 3310 1105 3311
rect 1166 3311 1167 3312
rect 1171 3311 1172 3315
rect 1166 3310 1172 3311
rect 1267 3315 1273 3316
rect 1267 3311 1268 3315
rect 1272 3314 1273 3315
rect 1342 3315 1348 3316
rect 1342 3314 1343 3315
rect 1272 3312 1343 3314
rect 1272 3311 1273 3312
rect 1267 3310 1273 3311
rect 1342 3311 1343 3312
rect 1347 3311 1348 3315
rect 1342 3310 1348 3311
rect 1426 3315 1432 3316
rect 1426 3311 1427 3315
rect 1431 3314 1432 3315
rect 1435 3315 1441 3316
rect 1435 3314 1436 3315
rect 1431 3312 1436 3314
rect 1431 3311 1432 3312
rect 1426 3310 1432 3311
rect 1435 3311 1436 3312
rect 1440 3311 1441 3315
rect 1618 3315 1624 3316
rect 1435 3310 1441 3311
rect 1594 3311 1601 3312
rect 202 3306 208 3307
rect 1594 3307 1595 3311
rect 1600 3307 1601 3311
rect 1618 3311 1619 3315
rect 1623 3314 1624 3315
rect 1755 3315 1761 3316
rect 1755 3314 1756 3315
rect 1623 3312 1756 3314
rect 1623 3311 1624 3312
rect 1618 3310 1624 3311
rect 1755 3311 1756 3312
rect 1760 3311 1761 3315
rect 1755 3310 1761 3311
rect 1778 3315 1784 3316
rect 1778 3311 1779 3315
rect 1783 3314 1784 3315
rect 1923 3315 1929 3316
rect 2046 3315 2052 3316
rect 3942 3315 3948 3316
rect 1923 3314 1924 3315
rect 1783 3312 1924 3314
rect 1783 3311 1784 3312
rect 1778 3310 1784 3311
rect 1923 3311 1924 3312
rect 1928 3311 1929 3315
rect 1923 3310 1929 3311
rect 1594 3306 1601 3307
rect 187 3299 193 3300
rect 187 3295 188 3299
rect 192 3298 193 3299
rect 254 3299 260 3300
rect 254 3298 255 3299
rect 192 3296 255 3298
rect 192 3295 193 3296
rect 187 3294 193 3295
rect 254 3295 255 3296
rect 259 3295 260 3299
rect 515 3299 524 3300
rect 254 3294 260 3295
rect 331 3297 337 3298
rect 331 3293 332 3297
rect 336 3293 337 3297
rect 515 3295 516 3299
rect 523 3295 524 3299
rect 515 3294 524 3295
rect 607 3299 613 3300
rect 607 3295 608 3299
rect 612 3298 613 3299
rect 715 3299 721 3300
rect 715 3298 716 3299
rect 612 3296 716 3298
rect 612 3295 613 3296
rect 607 3294 613 3295
rect 715 3295 716 3296
rect 720 3295 721 3299
rect 715 3294 721 3295
rect 738 3299 744 3300
rect 738 3295 739 3299
rect 743 3298 744 3299
rect 923 3299 929 3300
rect 923 3298 924 3299
rect 743 3296 924 3298
rect 743 3295 744 3296
rect 738 3294 744 3295
rect 923 3295 924 3296
rect 928 3295 929 3299
rect 923 3294 929 3295
rect 1122 3299 1128 3300
rect 1122 3295 1123 3299
rect 1127 3298 1128 3299
rect 1131 3299 1137 3300
rect 1131 3298 1132 3299
rect 1127 3296 1132 3298
rect 1127 3295 1128 3296
rect 1122 3294 1128 3295
rect 1131 3295 1132 3296
rect 1136 3295 1137 3299
rect 1131 3294 1137 3295
rect 1154 3299 1160 3300
rect 1154 3295 1155 3299
rect 1159 3298 1160 3299
rect 1347 3299 1353 3300
rect 1347 3298 1348 3299
rect 1159 3296 1348 3298
rect 1159 3295 1160 3296
rect 1154 3294 1160 3295
rect 1347 3295 1348 3296
rect 1352 3295 1353 3299
rect 1347 3294 1353 3295
rect 1571 3299 1577 3300
rect 1571 3295 1572 3299
rect 1576 3298 1577 3299
rect 1602 3299 1608 3300
rect 1602 3298 1603 3299
rect 1576 3296 1603 3298
rect 1576 3295 1577 3296
rect 1571 3294 1577 3295
rect 1602 3295 1603 3296
rect 1607 3295 1608 3299
rect 1602 3294 1608 3295
rect 1770 3299 1776 3300
rect 1770 3295 1771 3299
rect 1775 3298 1776 3299
rect 1795 3299 1801 3300
rect 1795 3298 1796 3299
rect 1775 3296 1796 3298
rect 1775 3295 1776 3296
rect 1770 3294 1776 3295
rect 1795 3295 1796 3296
rect 1800 3295 1801 3299
rect 1795 3294 1801 3295
rect 331 3292 337 3293
rect 332 3286 334 3292
rect 798 3287 804 3288
rect 798 3286 799 3287
rect 332 3284 799 3286
rect 798 3283 799 3284
rect 803 3283 804 3287
rect 798 3282 804 3283
rect 134 3276 140 3277
rect 110 3273 116 3274
rect 110 3269 111 3273
rect 115 3269 116 3273
rect 134 3272 135 3276
rect 139 3272 140 3276
rect 134 3271 140 3272
rect 278 3276 284 3277
rect 278 3272 279 3276
rect 283 3272 284 3276
rect 278 3271 284 3272
rect 462 3276 468 3277
rect 462 3272 463 3276
rect 467 3272 468 3276
rect 462 3271 468 3272
rect 662 3276 668 3277
rect 662 3272 663 3276
rect 667 3272 668 3276
rect 662 3271 668 3272
rect 870 3276 876 3277
rect 870 3272 871 3276
rect 875 3272 876 3276
rect 870 3271 876 3272
rect 1078 3276 1084 3277
rect 1078 3272 1079 3276
rect 1083 3272 1084 3276
rect 1078 3271 1084 3272
rect 1294 3276 1300 3277
rect 1294 3272 1295 3276
rect 1299 3272 1300 3276
rect 1294 3271 1300 3272
rect 1518 3276 1524 3277
rect 1518 3272 1519 3276
rect 1523 3272 1524 3276
rect 1518 3271 1524 3272
rect 1742 3276 1748 3277
rect 1742 3272 1743 3276
rect 1747 3272 1748 3276
rect 1742 3271 1748 3272
rect 2006 3273 2012 3274
rect 110 3268 116 3269
rect 2006 3269 2007 3273
rect 2011 3269 2012 3273
rect 2006 3268 2012 3269
rect 202 3267 208 3268
rect 202 3263 203 3267
rect 207 3263 208 3267
rect 202 3262 208 3263
rect 254 3267 260 3268
rect 254 3263 255 3267
rect 259 3266 260 3267
rect 607 3267 613 3268
rect 607 3266 608 3267
rect 259 3264 321 3266
rect 541 3264 608 3266
rect 259 3263 260 3264
rect 254 3262 260 3263
rect 607 3263 608 3264
rect 612 3263 613 3267
rect 607 3262 613 3263
rect 738 3267 744 3268
rect 738 3263 739 3267
rect 743 3263 744 3267
rect 738 3262 744 3263
rect 798 3267 804 3268
rect 798 3263 799 3267
rect 803 3266 804 3267
rect 1154 3267 1160 3268
rect 803 3264 913 3266
rect 803 3263 804 3264
rect 798 3262 804 3263
rect 1154 3263 1155 3267
rect 1159 3263 1160 3267
rect 1154 3262 1160 3263
rect 1370 3267 1376 3268
rect 1370 3263 1371 3267
rect 1375 3263 1376 3267
rect 1370 3262 1376 3263
rect 1594 3267 1600 3268
rect 1594 3263 1595 3267
rect 1599 3263 1600 3267
rect 1594 3262 1600 3263
rect 1602 3267 1608 3268
rect 1602 3263 1603 3267
rect 1607 3266 1608 3267
rect 1607 3264 1785 3266
rect 1607 3263 1608 3264
rect 1602 3262 1608 3263
rect 2046 3260 2052 3261
rect 3942 3260 3948 3261
rect 134 3257 140 3258
rect 110 3256 116 3257
rect 110 3252 111 3256
rect 115 3252 116 3256
rect 134 3253 135 3257
rect 139 3253 140 3257
rect 134 3252 140 3253
rect 278 3257 284 3258
rect 278 3253 279 3257
rect 283 3253 284 3257
rect 278 3252 284 3253
rect 462 3257 468 3258
rect 462 3253 463 3257
rect 467 3253 468 3257
rect 462 3252 468 3253
rect 662 3257 668 3258
rect 662 3253 663 3257
rect 667 3253 668 3257
rect 662 3252 668 3253
rect 870 3257 876 3258
rect 870 3253 871 3257
rect 875 3253 876 3257
rect 870 3252 876 3253
rect 1078 3257 1084 3258
rect 1078 3253 1079 3257
rect 1083 3253 1084 3257
rect 1078 3252 1084 3253
rect 1294 3257 1300 3258
rect 1294 3253 1295 3257
rect 1299 3253 1300 3257
rect 1294 3252 1300 3253
rect 1518 3257 1524 3258
rect 1518 3253 1519 3257
rect 1523 3253 1524 3257
rect 1518 3252 1524 3253
rect 1742 3257 1748 3258
rect 1742 3253 1743 3257
rect 1747 3253 1748 3257
rect 1742 3252 1748 3253
rect 2006 3256 2012 3257
rect 2006 3252 2007 3256
rect 2011 3252 2012 3256
rect 2046 3256 2047 3260
rect 2051 3256 2052 3260
rect 2046 3255 2052 3256
rect 2110 3259 2116 3260
rect 2110 3255 2111 3259
rect 2115 3255 2116 3259
rect 2110 3254 2116 3255
rect 2246 3259 2252 3260
rect 2246 3255 2247 3259
rect 2251 3255 2252 3259
rect 2246 3254 2252 3255
rect 2398 3259 2404 3260
rect 2398 3255 2399 3259
rect 2403 3255 2404 3259
rect 2398 3254 2404 3255
rect 2574 3259 2580 3260
rect 2574 3255 2575 3259
rect 2579 3255 2580 3259
rect 2574 3254 2580 3255
rect 2782 3259 2788 3260
rect 2782 3255 2783 3259
rect 2787 3255 2788 3259
rect 3014 3259 3020 3260
rect 2782 3254 2788 3255
rect 2870 3255 2876 3256
rect 110 3251 116 3252
rect 2006 3251 2012 3252
rect 2870 3251 2871 3255
rect 2875 3254 2876 3255
rect 3014 3255 3015 3259
rect 3019 3255 3020 3259
rect 3014 3254 3020 3255
rect 3262 3259 3268 3260
rect 3262 3255 3263 3259
rect 3267 3255 3268 3259
rect 3262 3254 3268 3255
rect 3526 3259 3532 3260
rect 3526 3255 3527 3259
rect 3531 3255 3532 3259
rect 3526 3254 3532 3255
rect 3790 3259 3796 3260
rect 3790 3255 3791 3259
rect 3795 3255 3796 3259
rect 3942 3256 3943 3260
rect 3947 3256 3948 3260
rect 3942 3255 3948 3256
rect 3790 3254 3796 3255
rect 2875 3252 2962 3254
rect 2875 3251 2876 3252
rect 2870 3250 2876 3251
rect 2960 3250 2962 3252
rect 3498 3251 3504 3252
rect 2960 3248 3057 3250
rect 2186 3247 2192 3248
rect 2046 3243 2052 3244
rect 2046 3239 2047 3243
rect 2051 3239 2052 3243
rect 2186 3243 2187 3247
rect 2191 3243 2192 3247
rect 2367 3247 2373 3248
rect 2367 3246 2368 3247
rect 2325 3244 2368 3246
rect 2186 3242 2192 3243
rect 2367 3243 2368 3244
rect 2372 3243 2373 3247
rect 2367 3242 2373 3243
rect 2474 3247 2480 3248
rect 2474 3243 2475 3247
rect 2479 3243 2480 3247
rect 2474 3242 2480 3243
rect 2650 3247 2656 3248
rect 2650 3243 2651 3247
rect 2655 3243 2656 3247
rect 2650 3242 2656 3243
rect 2858 3247 2864 3248
rect 2858 3243 2859 3247
rect 2863 3243 2864 3247
rect 2858 3242 2864 3243
rect 3338 3247 3344 3248
rect 3338 3243 3339 3247
rect 3343 3243 3344 3247
rect 3498 3247 3499 3251
rect 3503 3250 3504 3251
rect 3503 3248 3569 3250
rect 3503 3247 3504 3248
rect 3498 3246 3504 3247
rect 3866 3247 3872 3248
rect 3338 3242 3344 3243
rect 3866 3243 3867 3247
rect 3871 3243 3872 3247
rect 3866 3242 3872 3243
rect 3942 3243 3948 3244
rect 2046 3238 2052 3239
rect 2110 3240 2116 3241
rect 2110 3236 2111 3240
rect 2115 3236 2116 3240
rect 2110 3235 2116 3236
rect 2246 3240 2252 3241
rect 2246 3236 2247 3240
rect 2251 3236 2252 3240
rect 2246 3235 2252 3236
rect 2398 3240 2404 3241
rect 2398 3236 2399 3240
rect 2403 3236 2404 3240
rect 2398 3235 2404 3236
rect 2574 3240 2580 3241
rect 2574 3236 2575 3240
rect 2579 3236 2580 3240
rect 2574 3235 2580 3236
rect 2782 3240 2788 3241
rect 2782 3236 2783 3240
rect 2787 3236 2788 3240
rect 2782 3235 2788 3236
rect 3014 3240 3020 3241
rect 3014 3236 3015 3240
rect 3019 3236 3020 3240
rect 3014 3235 3020 3236
rect 3262 3240 3268 3241
rect 3262 3236 3263 3240
rect 3267 3236 3268 3240
rect 3262 3235 3268 3236
rect 3526 3240 3532 3241
rect 3526 3236 3527 3240
rect 3531 3236 3532 3240
rect 3526 3235 3532 3236
rect 3790 3240 3796 3241
rect 3790 3236 3791 3240
rect 3795 3236 3796 3240
rect 3942 3239 3943 3243
rect 3947 3239 3948 3243
rect 3942 3238 3948 3239
rect 3790 3235 3796 3236
rect 2146 3219 2152 3220
rect 2146 3215 2147 3219
rect 2151 3218 2152 3219
rect 2163 3219 2169 3220
rect 2163 3218 2164 3219
rect 2151 3216 2164 3218
rect 2151 3215 2152 3216
rect 2146 3214 2152 3215
rect 2163 3215 2164 3216
rect 2168 3215 2169 3219
rect 2367 3219 2373 3220
rect 2163 3214 2169 3215
rect 2299 3215 2305 3216
rect 2299 3211 2300 3215
rect 2304 3214 2305 3215
rect 2330 3215 2336 3216
rect 2330 3214 2331 3215
rect 2304 3212 2331 3214
rect 2304 3211 2305 3212
rect 2299 3210 2305 3211
rect 2330 3211 2331 3212
rect 2335 3211 2336 3215
rect 2367 3215 2368 3219
rect 2372 3218 2373 3219
rect 2451 3219 2457 3220
rect 2451 3218 2452 3219
rect 2372 3216 2452 3218
rect 2372 3215 2373 3216
rect 2367 3214 2373 3215
rect 2451 3215 2452 3216
rect 2456 3215 2457 3219
rect 2451 3214 2457 3215
rect 2474 3219 2480 3220
rect 2474 3215 2475 3219
rect 2479 3218 2480 3219
rect 2627 3219 2633 3220
rect 2627 3218 2628 3219
rect 2479 3216 2628 3218
rect 2479 3215 2480 3216
rect 2474 3214 2480 3215
rect 2627 3215 2628 3216
rect 2632 3215 2633 3219
rect 2627 3214 2633 3215
rect 2650 3219 2656 3220
rect 2650 3215 2651 3219
rect 2655 3218 2656 3219
rect 2835 3219 2841 3220
rect 2835 3218 2836 3219
rect 2655 3216 2836 3218
rect 2655 3215 2656 3216
rect 2650 3214 2656 3215
rect 2835 3215 2836 3216
rect 2840 3215 2841 3219
rect 2835 3214 2841 3215
rect 2858 3219 2864 3220
rect 2858 3215 2859 3219
rect 2863 3218 2864 3219
rect 3067 3219 3073 3220
rect 3067 3218 3068 3219
rect 2863 3216 3068 3218
rect 2863 3215 2864 3216
rect 2858 3214 2864 3215
rect 3067 3215 3068 3216
rect 3072 3215 3073 3219
rect 3506 3219 3512 3220
rect 3067 3214 3073 3215
rect 3310 3215 3321 3216
rect 2330 3210 2336 3211
rect 3310 3211 3311 3215
rect 3315 3211 3316 3215
rect 3320 3211 3321 3215
rect 3506 3215 3507 3219
rect 3511 3218 3512 3219
rect 3579 3219 3585 3220
rect 3579 3218 3580 3219
rect 3511 3216 3580 3218
rect 3511 3215 3512 3216
rect 3506 3214 3512 3215
rect 3579 3215 3580 3216
rect 3584 3215 3585 3219
rect 3579 3214 3585 3215
rect 3843 3219 3852 3220
rect 3843 3215 3844 3219
rect 3851 3215 3852 3219
rect 3843 3214 3852 3215
rect 3310 3210 3321 3211
rect 110 3204 116 3205
rect 2006 3204 2012 3205
rect 110 3200 111 3204
rect 115 3200 116 3204
rect 110 3199 116 3200
rect 134 3203 140 3204
rect 134 3199 135 3203
rect 139 3199 140 3203
rect 134 3198 140 3199
rect 286 3203 292 3204
rect 286 3199 287 3203
rect 291 3199 292 3203
rect 286 3198 292 3199
rect 446 3203 452 3204
rect 446 3199 447 3203
rect 451 3199 452 3203
rect 446 3198 452 3199
rect 614 3203 620 3204
rect 614 3199 615 3203
rect 619 3199 620 3203
rect 614 3198 620 3199
rect 790 3203 796 3204
rect 790 3199 791 3203
rect 795 3199 796 3203
rect 790 3198 796 3199
rect 966 3203 972 3204
rect 966 3199 967 3203
rect 971 3199 972 3203
rect 966 3198 972 3199
rect 1142 3203 1148 3204
rect 1142 3199 1143 3203
rect 1147 3199 1148 3203
rect 1142 3198 1148 3199
rect 1326 3203 1332 3204
rect 1326 3199 1327 3203
rect 1331 3199 1332 3203
rect 1326 3198 1332 3199
rect 1510 3203 1516 3204
rect 1510 3199 1511 3203
rect 1515 3199 1516 3203
rect 1510 3198 1516 3199
rect 1694 3203 1700 3204
rect 1694 3199 1695 3203
rect 1699 3199 1700 3203
rect 2006 3200 2007 3204
rect 2011 3200 2012 3204
rect 2006 3199 2012 3200
rect 2123 3203 2129 3204
rect 2123 3199 2124 3203
rect 2128 3202 2129 3203
rect 2186 3203 2192 3204
rect 2186 3202 2187 3203
rect 2128 3200 2187 3202
rect 2128 3199 2129 3200
rect 1694 3198 1700 3199
rect 2123 3198 2129 3199
rect 2186 3199 2187 3200
rect 2191 3199 2192 3203
rect 2315 3203 2321 3204
rect 2186 3198 2192 3199
rect 2219 3201 2225 3202
rect 2219 3197 2220 3201
rect 2224 3197 2225 3201
rect 2315 3199 2316 3203
rect 2320 3202 2321 3203
rect 2346 3203 2352 3204
rect 2346 3202 2347 3203
rect 2320 3200 2347 3202
rect 2320 3199 2321 3200
rect 2315 3198 2321 3199
rect 2346 3199 2347 3200
rect 2351 3199 2352 3203
rect 2346 3198 2352 3199
rect 2411 3203 2417 3204
rect 2411 3199 2412 3203
rect 2416 3202 2417 3203
rect 2442 3203 2448 3204
rect 2442 3202 2443 3203
rect 2416 3200 2443 3202
rect 2416 3199 2417 3200
rect 2411 3198 2417 3199
rect 2442 3199 2443 3200
rect 2447 3199 2448 3203
rect 2442 3198 2448 3199
rect 2507 3203 2513 3204
rect 2507 3199 2508 3203
rect 2512 3202 2513 3203
rect 2538 3203 2544 3204
rect 2538 3202 2539 3203
rect 2512 3200 2539 3202
rect 2512 3199 2513 3200
rect 2507 3198 2513 3199
rect 2538 3199 2539 3200
rect 2543 3199 2544 3203
rect 2538 3198 2544 3199
rect 2603 3203 2609 3204
rect 2603 3199 2604 3203
rect 2608 3202 2609 3203
rect 2634 3203 2640 3204
rect 2634 3202 2635 3203
rect 2608 3200 2635 3202
rect 2608 3199 2609 3200
rect 2603 3198 2609 3199
rect 2634 3199 2635 3200
rect 2639 3199 2640 3203
rect 2634 3198 2640 3199
rect 2699 3203 2705 3204
rect 2699 3199 2700 3203
rect 2704 3202 2705 3203
rect 2730 3203 2736 3204
rect 2730 3202 2731 3203
rect 2704 3200 2731 3202
rect 2704 3199 2705 3200
rect 2699 3198 2705 3199
rect 2730 3199 2731 3200
rect 2735 3199 2736 3203
rect 2730 3198 2736 3199
rect 2795 3203 2801 3204
rect 2795 3199 2796 3203
rect 2800 3202 2801 3203
rect 2826 3203 2832 3204
rect 2826 3202 2827 3203
rect 2800 3200 2827 3202
rect 2800 3199 2801 3200
rect 2795 3198 2801 3199
rect 2826 3199 2827 3200
rect 2831 3199 2832 3203
rect 2826 3198 2832 3199
rect 2891 3203 2897 3204
rect 2891 3199 2892 3203
rect 2896 3202 2897 3203
rect 2922 3203 2928 3204
rect 2922 3202 2923 3203
rect 2896 3200 2923 3202
rect 2896 3199 2897 3200
rect 2891 3198 2897 3199
rect 2922 3199 2923 3200
rect 2927 3199 2928 3203
rect 2922 3198 2928 3199
rect 2987 3203 2993 3204
rect 2987 3199 2988 3203
rect 2992 3202 2993 3203
rect 3022 3203 3028 3204
rect 3022 3202 3023 3203
rect 2992 3200 3023 3202
rect 2992 3199 2993 3200
rect 2987 3198 2993 3199
rect 3022 3199 3023 3200
rect 3027 3199 3028 3203
rect 3022 3198 3028 3199
rect 3083 3203 3089 3204
rect 3083 3199 3084 3203
rect 3088 3202 3089 3203
rect 3114 3203 3120 3204
rect 3114 3202 3115 3203
rect 3088 3200 3115 3202
rect 3088 3199 3089 3200
rect 3083 3198 3089 3199
rect 3114 3199 3115 3200
rect 3119 3199 3120 3203
rect 3114 3198 3120 3199
rect 3179 3203 3185 3204
rect 3179 3199 3180 3203
rect 3184 3202 3185 3203
rect 3210 3203 3216 3204
rect 3210 3202 3211 3203
rect 3184 3200 3211 3202
rect 3184 3199 3185 3200
rect 3179 3198 3185 3199
rect 3210 3199 3211 3200
rect 3215 3199 3216 3203
rect 3210 3198 3216 3199
rect 3275 3203 3281 3204
rect 3275 3199 3276 3203
rect 3280 3202 3281 3203
rect 3338 3203 3344 3204
rect 3338 3202 3339 3203
rect 3280 3200 3339 3202
rect 3280 3199 3281 3200
rect 3275 3198 3281 3199
rect 3338 3199 3339 3200
rect 3343 3199 3344 3203
rect 3338 3198 3344 3199
rect 3371 3203 3377 3204
rect 3371 3199 3372 3203
rect 3376 3202 3377 3203
rect 3402 3203 3408 3204
rect 3402 3202 3403 3203
rect 3376 3200 3403 3202
rect 3376 3199 3377 3200
rect 3371 3198 3377 3199
rect 3402 3199 3403 3200
rect 3407 3199 3408 3203
rect 3586 3203 3592 3204
rect 3402 3198 3408 3199
rect 3491 3201 3497 3202
rect 2219 3196 2225 3197
rect 3491 3197 3492 3201
rect 3496 3197 3497 3201
rect 3586 3199 3587 3203
rect 3591 3202 3592 3203
rect 3627 3203 3633 3204
rect 3627 3202 3628 3203
rect 3591 3200 3628 3202
rect 3591 3199 3592 3200
rect 3586 3198 3592 3199
rect 3627 3199 3628 3200
rect 3632 3199 3633 3203
rect 3627 3198 3633 3199
rect 3650 3203 3656 3204
rect 3650 3199 3651 3203
rect 3655 3202 3656 3203
rect 3771 3203 3777 3204
rect 3771 3202 3772 3203
rect 3655 3200 3772 3202
rect 3655 3199 3656 3200
rect 3650 3198 3656 3199
rect 3771 3199 3772 3200
rect 3776 3199 3777 3203
rect 3771 3198 3777 3199
rect 3891 3203 3897 3204
rect 3891 3199 3892 3203
rect 3896 3202 3897 3203
rect 3914 3203 3920 3204
rect 3914 3202 3915 3203
rect 3896 3200 3915 3202
rect 3896 3199 3897 3200
rect 3891 3198 3897 3199
rect 3914 3199 3915 3200
rect 3919 3199 3920 3203
rect 3914 3198 3920 3199
rect 3491 3196 3497 3197
rect 522 3195 528 3196
rect 258 3191 264 3192
rect 258 3190 259 3191
rect 213 3188 259 3190
rect 110 3187 116 3188
rect 110 3183 111 3187
rect 115 3183 116 3187
rect 258 3187 259 3188
rect 263 3187 264 3191
rect 258 3186 264 3187
rect 362 3191 368 3192
rect 362 3187 363 3191
rect 367 3187 368 3191
rect 522 3191 523 3195
rect 527 3191 528 3195
rect 522 3190 528 3191
rect 558 3195 564 3196
rect 558 3191 559 3195
rect 563 3194 564 3195
rect 750 3195 756 3196
rect 563 3192 657 3194
rect 563 3191 564 3192
rect 558 3190 564 3191
rect 750 3191 751 3195
rect 755 3194 756 3195
rect 1090 3195 1096 3196
rect 755 3192 833 3194
rect 755 3191 756 3192
rect 750 3190 756 3191
rect 1042 3191 1048 3192
rect 362 3186 368 3187
rect 1042 3187 1043 3191
rect 1047 3187 1048 3191
rect 1090 3191 1091 3195
rect 1095 3194 1096 3195
rect 1231 3195 1237 3196
rect 1095 3192 1185 3194
rect 1095 3191 1096 3192
rect 1090 3190 1096 3191
rect 1231 3191 1232 3195
rect 1236 3194 1237 3195
rect 1770 3195 1776 3196
rect 1236 3192 1369 3194
rect 1236 3191 1237 3192
rect 1231 3190 1237 3191
rect 1586 3191 1592 3192
rect 1042 3186 1048 3187
rect 1586 3187 1587 3191
rect 1591 3187 1592 3191
rect 1770 3191 1771 3195
rect 1775 3191 1776 3195
rect 1770 3190 1776 3191
rect 2146 3195 2152 3196
rect 2146 3191 2147 3195
rect 2151 3194 2152 3195
rect 2220 3194 2222 3196
rect 2151 3192 2222 3194
rect 3492 3194 3494 3196
rect 3658 3195 3664 3196
rect 3658 3194 3659 3195
rect 3492 3192 3659 3194
rect 2151 3191 2152 3192
rect 2146 3190 2152 3191
rect 3658 3191 3659 3192
rect 3663 3191 3664 3195
rect 3658 3190 3664 3191
rect 1586 3186 1592 3187
rect 2006 3187 2012 3188
rect 110 3182 116 3183
rect 134 3184 140 3185
rect 134 3180 135 3184
rect 139 3180 140 3184
rect 134 3179 140 3180
rect 286 3184 292 3185
rect 286 3180 287 3184
rect 291 3180 292 3184
rect 286 3179 292 3180
rect 446 3184 452 3185
rect 446 3180 447 3184
rect 451 3180 452 3184
rect 446 3179 452 3180
rect 614 3184 620 3185
rect 614 3180 615 3184
rect 619 3180 620 3184
rect 614 3179 620 3180
rect 790 3184 796 3185
rect 790 3180 791 3184
rect 795 3180 796 3184
rect 790 3179 796 3180
rect 966 3184 972 3185
rect 966 3180 967 3184
rect 971 3180 972 3184
rect 966 3179 972 3180
rect 1142 3184 1148 3185
rect 1142 3180 1143 3184
rect 1147 3180 1148 3184
rect 1142 3179 1148 3180
rect 1326 3184 1332 3185
rect 1326 3180 1327 3184
rect 1331 3180 1332 3184
rect 1326 3179 1332 3180
rect 1510 3184 1516 3185
rect 1510 3180 1511 3184
rect 1515 3180 1516 3184
rect 1510 3179 1516 3180
rect 1694 3184 1700 3185
rect 1694 3180 1695 3184
rect 1699 3180 1700 3184
rect 2006 3183 2007 3187
rect 2011 3183 2012 3187
rect 2006 3182 2012 3183
rect 1694 3179 1700 3180
rect 2070 3180 2076 3181
rect 2046 3177 2052 3178
rect 2046 3173 2047 3177
rect 2051 3173 2052 3177
rect 2070 3176 2071 3180
rect 2075 3176 2076 3180
rect 2070 3175 2076 3176
rect 2166 3180 2172 3181
rect 2166 3176 2167 3180
rect 2171 3176 2172 3180
rect 2166 3175 2172 3176
rect 2262 3180 2268 3181
rect 2262 3176 2263 3180
rect 2267 3176 2268 3180
rect 2262 3175 2268 3176
rect 2358 3180 2364 3181
rect 2358 3176 2359 3180
rect 2363 3176 2364 3180
rect 2358 3175 2364 3176
rect 2454 3180 2460 3181
rect 2454 3176 2455 3180
rect 2459 3176 2460 3180
rect 2454 3175 2460 3176
rect 2550 3180 2556 3181
rect 2550 3176 2551 3180
rect 2555 3176 2556 3180
rect 2550 3175 2556 3176
rect 2646 3180 2652 3181
rect 2646 3176 2647 3180
rect 2651 3176 2652 3180
rect 2646 3175 2652 3176
rect 2742 3180 2748 3181
rect 2742 3176 2743 3180
rect 2747 3176 2748 3180
rect 2742 3175 2748 3176
rect 2838 3180 2844 3181
rect 2838 3176 2839 3180
rect 2843 3176 2844 3180
rect 2838 3175 2844 3176
rect 2934 3180 2940 3181
rect 2934 3176 2935 3180
rect 2939 3176 2940 3180
rect 2934 3175 2940 3176
rect 3030 3180 3036 3181
rect 3030 3176 3031 3180
rect 3035 3176 3036 3180
rect 3030 3175 3036 3176
rect 3126 3180 3132 3181
rect 3126 3176 3127 3180
rect 3131 3176 3132 3180
rect 3126 3175 3132 3176
rect 3222 3180 3228 3181
rect 3222 3176 3223 3180
rect 3227 3176 3228 3180
rect 3222 3175 3228 3176
rect 3318 3180 3324 3181
rect 3318 3176 3319 3180
rect 3323 3176 3324 3180
rect 3318 3175 3324 3176
rect 3438 3180 3444 3181
rect 3438 3176 3439 3180
rect 3443 3176 3444 3180
rect 3438 3175 3444 3176
rect 3574 3180 3580 3181
rect 3574 3176 3575 3180
rect 3579 3176 3580 3180
rect 3574 3175 3580 3176
rect 3718 3180 3724 3181
rect 3718 3176 3719 3180
rect 3723 3176 3724 3180
rect 3718 3175 3724 3176
rect 3838 3180 3844 3181
rect 3838 3176 3839 3180
rect 3843 3176 3844 3180
rect 3838 3175 3844 3176
rect 3942 3177 3948 3178
rect 2046 3172 2052 3173
rect 3942 3173 3943 3177
rect 3947 3173 3948 3177
rect 3942 3172 3948 3173
rect 558 3171 564 3172
rect 558 3170 559 3171
rect 319 3168 559 3170
rect 319 3166 321 3168
rect 558 3167 559 3168
rect 563 3167 564 3171
rect 558 3166 564 3167
rect 2146 3171 2152 3172
rect 2146 3167 2147 3171
rect 2151 3167 2152 3171
rect 2330 3171 2336 3172
rect 2146 3166 2152 3167
rect 252 3164 321 3166
rect 187 3163 193 3164
rect 187 3159 188 3163
rect 192 3162 193 3163
rect 252 3162 254 3164
rect 192 3160 254 3162
rect 362 3163 368 3164
rect 192 3159 193 3160
rect 187 3158 193 3159
rect 258 3159 264 3160
rect 258 3155 259 3159
rect 263 3158 264 3159
rect 339 3159 345 3160
rect 339 3158 340 3159
rect 263 3156 340 3158
rect 263 3155 264 3156
rect 258 3154 264 3155
rect 339 3155 340 3156
rect 344 3155 345 3159
rect 362 3159 363 3163
rect 367 3162 368 3163
rect 499 3163 505 3164
rect 499 3162 500 3163
rect 367 3160 500 3162
rect 367 3159 368 3160
rect 362 3158 368 3159
rect 499 3159 500 3160
rect 504 3159 505 3163
rect 499 3158 505 3159
rect 667 3163 673 3164
rect 667 3159 668 3163
rect 672 3162 673 3163
rect 750 3163 756 3164
rect 750 3162 751 3163
rect 672 3160 751 3162
rect 672 3159 673 3160
rect 667 3158 673 3159
rect 750 3159 751 3160
rect 755 3159 756 3163
rect 1019 3163 1025 3164
rect 750 3158 756 3159
rect 843 3159 849 3160
rect 339 3154 345 3155
rect 843 3155 844 3159
rect 848 3158 849 3159
rect 863 3159 869 3160
rect 863 3158 864 3159
rect 848 3156 864 3158
rect 848 3155 849 3156
rect 843 3154 849 3155
rect 863 3155 864 3156
rect 868 3155 869 3159
rect 1019 3159 1020 3163
rect 1024 3162 1025 3163
rect 1090 3163 1096 3164
rect 1090 3162 1091 3163
rect 1024 3160 1091 3162
rect 1024 3159 1025 3160
rect 1019 3158 1025 3159
rect 1090 3159 1091 3160
rect 1095 3159 1096 3163
rect 1090 3158 1096 3159
rect 1195 3163 1201 3164
rect 1195 3159 1196 3163
rect 1200 3162 1201 3163
rect 1231 3163 1237 3164
rect 1231 3162 1232 3163
rect 1200 3160 1232 3162
rect 1200 3159 1201 3160
rect 1195 3158 1201 3159
rect 1231 3159 1232 3160
rect 1236 3159 1237 3163
rect 1231 3158 1237 3159
rect 1370 3163 1376 3164
rect 1370 3159 1371 3163
rect 1375 3162 1376 3163
rect 1379 3163 1385 3164
rect 1379 3162 1380 3163
rect 1375 3160 1380 3162
rect 1375 3159 1376 3160
rect 1370 3158 1376 3159
rect 1379 3159 1380 3160
rect 1384 3159 1385 3163
rect 1586 3163 1592 3164
rect 1379 3158 1385 3159
rect 1466 3159 1472 3160
rect 863 3154 869 3155
rect 1466 3155 1467 3159
rect 1471 3158 1472 3159
rect 1563 3159 1569 3160
rect 1563 3158 1564 3159
rect 1471 3156 1564 3158
rect 1471 3155 1472 3156
rect 1466 3154 1472 3155
rect 1563 3155 1564 3156
rect 1568 3155 1569 3159
rect 1586 3159 1587 3163
rect 1591 3162 1592 3163
rect 1747 3163 1753 3164
rect 1747 3162 1748 3163
rect 1591 3160 1748 3162
rect 1591 3159 1592 3160
rect 1586 3158 1592 3159
rect 1747 3159 1748 3160
rect 1752 3159 1753 3163
rect 2070 3161 2076 3162
rect 1747 3158 1753 3159
rect 2046 3160 2052 3161
rect 2046 3156 2047 3160
rect 2051 3156 2052 3160
rect 2070 3157 2071 3161
rect 2075 3157 2076 3161
rect 2070 3156 2076 3157
rect 2166 3161 2172 3162
rect 2166 3157 2167 3161
rect 2171 3157 2172 3161
rect 2166 3156 2172 3157
rect 2046 3155 2052 3156
rect 1563 3154 1569 3155
rect 2244 3154 2246 3169
rect 2330 3167 2331 3171
rect 2335 3167 2336 3171
rect 2330 3166 2336 3167
rect 2346 3171 2352 3172
rect 2346 3167 2347 3171
rect 2351 3170 2352 3171
rect 2442 3171 2448 3172
rect 2351 3168 2401 3170
rect 2351 3167 2352 3168
rect 2346 3166 2352 3167
rect 2442 3167 2443 3171
rect 2447 3170 2448 3171
rect 2538 3171 2544 3172
rect 2447 3168 2497 3170
rect 2447 3167 2448 3168
rect 2442 3166 2448 3167
rect 2538 3167 2539 3171
rect 2543 3170 2544 3171
rect 2634 3171 2640 3172
rect 2543 3168 2593 3170
rect 2543 3167 2544 3168
rect 2538 3166 2544 3167
rect 2634 3167 2635 3171
rect 2639 3170 2640 3171
rect 2730 3171 2736 3172
rect 2639 3168 2689 3170
rect 2639 3167 2640 3168
rect 2634 3166 2640 3167
rect 2730 3167 2731 3171
rect 2735 3170 2736 3171
rect 2826 3171 2832 3172
rect 2735 3168 2785 3170
rect 2735 3167 2736 3168
rect 2730 3166 2736 3167
rect 2826 3167 2827 3171
rect 2831 3170 2832 3171
rect 2922 3171 2928 3172
rect 2831 3168 2881 3170
rect 2831 3167 2832 3168
rect 2826 3166 2832 3167
rect 2922 3167 2923 3171
rect 2927 3170 2928 3171
rect 3022 3171 3028 3172
rect 2927 3168 2977 3170
rect 2927 3167 2928 3168
rect 2922 3166 2928 3167
rect 3022 3167 3023 3171
rect 3027 3170 3028 3171
rect 3114 3171 3120 3172
rect 3027 3168 3073 3170
rect 3027 3167 3028 3168
rect 3022 3166 3028 3167
rect 3114 3167 3115 3171
rect 3119 3170 3120 3171
rect 3210 3171 3216 3172
rect 3119 3168 3169 3170
rect 3119 3167 3120 3168
rect 3114 3166 3120 3167
rect 3210 3167 3211 3171
rect 3215 3170 3216 3171
rect 3310 3171 3316 3172
rect 3215 3168 3265 3170
rect 3215 3167 3216 3168
rect 3210 3166 3216 3167
rect 3310 3167 3311 3171
rect 3315 3170 3316 3171
rect 3402 3171 3408 3172
rect 3315 3168 3361 3170
rect 3315 3167 3316 3168
rect 3310 3166 3316 3167
rect 3402 3167 3403 3171
rect 3407 3170 3408 3171
rect 3650 3171 3656 3172
rect 3407 3168 3481 3170
rect 3407 3167 3408 3168
rect 3402 3166 3408 3167
rect 3650 3167 3651 3171
rect 3655 3167 3656 3171
rect 3650 3166 3656 3167
rect 3658 3171 3664 3172
rect 3658 3167 3659 3171
rect 3663 3170 3664 3171
rect 3906 3171 3912 3172
rect 3663 3168 3761 3170
rect 3663 3167 3664 3168
rect 3658 3166 3664 3167
rect 3906 3167 3907 3171
rect 3911 3167 3912 3171
rect 3906 3166 3912 3167
rect 2262 3161 2268 3162
rect 2262 3157 2263 3161
rect 2267 3157 2268 3161
rect 2262 3156 2268 3157
rect 2358 3161 2364 3162
rect 2358 3157 2359 3161
rect 2363 3157 2364 3161
rect 2358 3156 2364 3157
rect 2454 3161 2460 3162
rect 2454 3157 2455 3161
rect 2459 3157 2460 3161
rect 2454 3156 2460 3157
rect 2550 3161 2556 3162
rect 2550 3157 2551 3161
rect 2555 3157 2556 3161
rect 2550 3156 2556 3157
rect 2646 3161 2652 3162
rect 2646 3157 2647 3161
rect 2651 3157 2652 3161
rect 2646 3156 2652 3157
rect 2742 3161 2748 3162
rect 2742 3157 2743 3161
rect 2747 3157 2748 3161
rect 2742 3156 2748 3157
rect 2838 3161 2844 3162
rect 2838 3157 2839 3161
rect 2843 3157 2844 3161
rect 2838 3156 2844 3157
rect 2934 3161 2940 3162
rect 2934 3157 2935 3161
rect 2939 3157 2940 3161
rect 2934 3156 2940 3157
rect 3030 3161 3036 3162
rect 3030 3157 3031 3161
rect 3035 3157 3036 3161
rect 3030 3156 3036 3157
rect 3126 3161 3132 3162
rect 3126 3157 3127 3161
rect 3131 3157 3132 3161
rect 3126 3156 3132 3157
rect 3222 3161 3228 3162
rect 3222 3157 3223 3161
rect 3227 3157 3228 3161
rect 3222 3156 3228 3157
rect 3318 3161 3324 3162
rect 3318 3157 3319 3161
rect 3323 3157 3324 3161
rect 3318 3156 3324 3157
rect 3438 3161 3444 3162
rect 3438 3157 3439 3161
rect 3443 3157 3444 3161
rect 3438 3156 3444 3157
rect 3574 3161 3580 3162
rect 3574 3157 3575 3161
rect 3579 3157 3580 3161
rect 3574 3156 3580 3157
rect 3718 3161 3724 3162
rect 3718 3157 3719 3161
rect 3723 3157 3724 3161
rect 3718 3156 3724 3157
rect 3838 3161 3844 3162
rect 3838 3157 3839 3161
rect 3843 3157 3844 3161
rect 3838 3156 3844 3157
rect 3942 3160 3948 3161
rect 3942 3156 3943 3160
rect 3947 3156 3948 3160
rect 2298 3155 2304 3156
rect 3942 3155 3948 3156
rect 2298 3154 2299 3155
rect 2244 3152 2299 3154
rect 2298 3151 2299 3152
rect 2303 3151 2304 3155
rect 2298 3150 2304 3151
rect 363 3143 372 3144
rect 363 3139 364 3143
rect 371 3139 372 3143
rect 363 3138 372 3139
rect 386 3143 392 3144
rect 386 3139 387 3143
rect 391 3142 392 3143
rect 491 3143 497 3144
rect 491 3142 492 3143
rect 391 3140 492 3142
rect 391 3139 392 3140
rect 386 3138 392 3139
rect 491 3139 492 3140
rect 496 3139 497 3143
rect 491 3138 497 3139
rect 514 3143 520 3144
rect 514 3139 515 3143
rect 519 3142 520 3143
rect 635 3143 641 3144
rect 635 3142 636 3143
rect 519 3140 636 3142
rect 519 3139 520 3140
rect 514 3138 520 3139
rect 635 3139 636 3140
rect 640 3139 641 3143
rect 635 3138 641 3139
rect 658 3143 664 3144
rect 658 3139 659 3143
rect 663 3142 664 3143
rect 795 3143 801 3144
rect 795 3142 796 3143
rect 663 3140 796 3142
rect 663 3139 664 3140
rect 658 3138 664 3139
rect 795 3139 796 3140
rect 800 3139 801 3143
rect 795 3138 801 3139
rect 818 3143 824 3144
rect 818 3139 819 3143
rect 823 3142 824 3143
rect 955 3143 961 3144
rect 955 3142 956 3143
rect 823 3140 956 3142
rect 823 3139 824 3140
rect 818 3138 824 3139
rect 955 3139 956 3140
rect 960 3139 961 3143
rect 955 3138 961 3139
rect 1042 3143 1048 3144
rect 1042 3139 1043 3143
rect 1047 3142 1048 3143
rect 1115 3143 1121 3144
rect 1115 3142 1116 3143
rect 1047 3140 1116 3142
rect 1047 3139 1048 3140
rect 1042 3138 1048 3139
rect 1115 3139 1116 3140
rect 1120 3139 1121 3143
rect 1115 3138 1121 3139
rect 1215 3143 1221 3144
rect 1215 3139 1216 3143
rect 1220 3142 1221 3143
rect 1275 3143 1281 3144
rect 1275 3142 1276 3143
rect 1220 3140 1276 3142
rect 1220 3139 1221 3140
rect 1215 3138 1221 3139
rect 1275 3139 1276 3140
rect 1280 3139 1281 3143
rect 1275 3138 1281 3139
rect 1443 3143 1449 3144
rect 1443 3139 1444 3143
rect 1448 3142 1449 3143
rect 1474 3143 1480 3144
rect 1474 3142 1475 3143
rect 1448 3140 1475 3142
rect 1448 3139 1449 3140
rect 1443 3138 1449 3139
rect 1474 3139 1475 3140
rect 1479 3139 1480 3143
rect 1474 3138 1480 3139
rect 1611 3143 1617 3144
rect 1611 3139 1612 3143
rect 1616 3142 1617 3143
rect 1642 3143 1648 3144
rect 1642 3142 1643 3143
rect 1616 3140 1643 3142
rect 1616 3139 1617 3140
rect 1611 3138 1617 3139
rect 1642 3139 1643 3140
rect 1647 3139 1648 3143
rect 1642 3138 1648 3139
rect 1779 3143 1785 3144
rect 1779 3139 1780 3143
rect 1784 3142 1785 3143
rect 1794 3143 1800 3144
rect 1794 3142 1795 3143
rect 1784 3140 1795 3142
rect 1784 3139 1785 3140
rect 1779 3138 1785 3139
rect 1794 3139 1795 3140
rect 1799 3139 1800 3143
rect 1794 3138 1800 3139
rect 310 3120 316 3121
rect 110 3117 116 3118
rect 110 3113 111 3117
rect 115 3113 116 3117
rect 310 3116 311 3120
rect 315 3116 316 3120
rect 310 3115 316 3116
rect 438 3120 444 3121
rect 438 3116 439 3120
rect 443 3116 444 3120
rect 438 3115 444 3116
rect 582 3120 588 3121
rect 582 3116 583 3120
rect 587 3116 588 3120
rect 582 3115 588 3116
rect 742 3120 748 3121
rect 742 3116 743 3120
rect 747 3116 748 3120
rect 742 3115 748 3116
rect 902 3120 908 3121
rect 902 3116 903 3120
rect 907 3116 908 3120
rect 902 3115 908 3116
rect 1062 3120 1068 3121
rect 1062 3116 1063 3120
rect 1067 3116 1068 3120
rect 1062 3115 1068 3116
rect 1222 3120 1228 3121
rect 1222 3116 1223 3120
rect 1227 3116 1228 3120
rect 1222 3115 1228 3116
rect 1390 3120 1396 3121
rect 1390 3116 1391 3120
rect 1395 3116 1396 3120
rect 1390 3115 1396 3116
rect 1558 3120 1564 3121
rect 1558 3116 1559 3120
rect 1563 3116 1564 3120
rect 1558 3115 1564 3116
rect 1726 3120 1732 3121
rect 1726 3116 1727 3120
rect 1731 3116 1732 3120
rect 1726 3115 1732 3116
rect 2006 3117 2012 3118
rect 110 3112 116 3113
rect 2006 3113 2007 3117
rect 2011 3113 2012 3117
rect 2006 3112 2012 3113
rect 386 3111 392 3112
rect 386 3107 387 3111
rect 391 3107 392 3111
rect 386 3106 392 3107
rect 514 3111 520 3112
rect 514 3107 515 3111
rect 519 3107 520 3111
rect 514 3106 520 3107
rect 658 3111 664 3112
rect 658 3107 659 3111
rect 663 3107 664 3111
rect 658 3106 664 3107
rect 818 3111 824 3112
rect 818 3107 819 3111
rect 823 3107 824 3111
rect 818 3106 824 3107
rect 863 3111 869 3112
rect 863 3107 864 3111
rect 868 3110 869 3111
rect 1215 3111 1221 3112
rect 1215 3110 1216 3111
rect 868 3108 945 3110
rect 1141 3108 1216 3110
rect 868 3107 869 3108
rect 863 3106 869 3107
rect 1215 3107 1216 3108
rect 1220 3107 1221 3111
rect 1350 3111 1356 3112
rect 1350 3110 1351 3111
rect 1301 3108 1351 3110
rect 1215 3106 1221 3107
rect 1350 3107 1351 3108
rect 1355 3107 1356 3111
rect 1350 3106 1356 3107
rect 1466 3111 1472 3112
rect 1466 3107 1467 3111
rect 1471 3107 1472 3111
rect 1466 3106 1472 3107
rect 1474 3111 1480 3112
rect 1474 3107 1475 3111
rect 1479 3110 1480 3111
rect 1642 3111 1648 3112
rect 1479 3108 1601 3110
rect 1479 3107 1480 3108
rect 1474 3106 1480 3107
rect 1642 3107 1643 3111
rect 1647 3110 1648 3111
rect 1647 3108 1769 3110
rect 1647 3107 1648 3108
rect 1642 3106 1648 3107
rect 310 3101 316 3102
rect 110 3100 116 3101
rect 110 3096 111 3100
rect 115 3096 116 3100
rect 310 3097 311 3101
rect 315 3097 316 3101
rect 310 3096 316 3097
rect 438 3101 444 3102
rect 438 3097 439 3101
rect 443 3097 444 3101
rect 438 3096 444 3097
rect 582 3101 588 3102
rect 582 3097 583 3101
rect 587 3097 588 3101
rect 582 3096 588 3097
rect 742 3101 748 3102
rect 742 3097 743 3101
rect 747 3097 748 3101
rect 742 3096 748 3097
rect 902 3101 908 3102
rect 902 3097 903 3101
rect 907 3097 908 3101
rect 902 3096 908 3097
rect 1062 3101 1068 3102
rect 1062 3097 1063 3101
rect 1067 3097 1068 3101
rect 1062 3096 1068 3097
rect 1222 3101 1228 3102
rect 1222 3097 1223 3101
rect 1227 3097 1228 3101
rect 1222 3096 1228 3097
rect 1390 3101 1396 3102
rect 1390 3097 1391 3101
rect 1395 3097 1396 3101
rect 1390 3096 1396 3097
rect 1558 3101 1564 3102
rect 1558 3097 1559 3101
rect 1563 3097 1564 3101
rect 1558 3096 1564 3097
rect 1726 3101 1732 3102
rect 1726 3097 1727 3101
rect 1731 3097 1732 3101
rect 1726 3096 1732 3097
rect 2006 3100 2012 3101
rect 2006 3096 2007 3100
rect 2011 3096 2012 3100
rect 110 3095 116 3096
rect 2006 3095 2012 3096
rect 2046 3096 2052 3097
rect 3942 3096 3948 3097
rect 2046 3092 2047 3096
rect 2051 3092 2052 3096
rect 2046 3091 2052 3092
rect 2070 3095 2076 3096
rect 2070 3091 2071 3095
rect 2075 3091 2076 3095
rect 2070 3090 2076 3091
rect 2334 3095 2340 3096
rect 2334 3091 2335 3095
rect 2339 3091 2340 3095
rect 2334 3090 2340 3091
rect 2622 3095 2628 3096
rect 2622 3091 2623 3095
rect 2627 3091 2628 3095
rect 2622 3090 2628 3091
rect 2910 3095 2916 3096
rect 2910 3091 2911 3095
rect 2915 3091 2916 3095
rect 2910 3090 2916 3091
rect 3206 3095 3212 3096
rect 3206 3091 3207 3095
rect 3211 3091 3212 3095
rect 3206 3090 3212 3091
rect 3502 3095 3508 3096
rect 3502 3091 3503 3095
rect 3507 3091 3508 3095
rect 3502 3090 3508 3091
rect 3798 3095 3804 3096
rect 3798 3091 3799 3095
rect 3803 3091 3804 3095
rect 3942 3092 3943 3096
rect 3947 3092 3948 3096
rect 3942 3091 3948 3092
rect 3798 3090 3804 3091
rect 2182 3087 2188 3088
rect 2146 3083 2152 3084
rect 2046 3079 2052 3080
rect 2046 3075 2047 3079
rect 2051 3075 2052 3079
rect 2146 3079 2147 3083
rect 2151 3079 2152 3083
rect 2182 3083 2183 3087
rect 2187 3086 2188 3087
rect 3586 3087 3592 3088
rect 3586 3086 3587 3087
rect 2187 3084 2377 3086
rect 3581 3084 3587 3086
rect 2187 3083 2188 3084
rect 2182 3082 2188 3083
rect 2698 3083 2704 3084
rect 2146 3078 2152 3079
rect 2698 3079 2699 3083
rect 2703 3079 2704 3083
rect 2698 3078 2704 3079
rect 2986 3083 2992 3084
rect 2986 3079 2987 3083
rect 2991 3079 2992 3083
rect 2986 3078 2992 3079
rect 3282 3083 3288 3084
rect 3282 3079 3283 3083
rect 3287 3079 3288 3083
rect 3586 3083 3587 3084
rect 3591 3083 3592 3087
rect 3586 3082 3592 3083
rect 3874 3083 3880 3084
rect 3282 3078 3288 3079
rect 3874 3079 3875 3083
rect 3879 3079 3880 3083
rect 3874 3078 3880 3079
rect 3942 3079 3948 3080
rect 2046 3074 2052 3075
rect 2070 3076 2076 3077
rect 2070 3072 2071 3076
rect 2075 3072 2076 3076
rect 2070 3071 2076 3072
rect 2334 3076 2340 3077
rect 2334 3072 2335 3076
rect 2339 3072 2340 3076
rect 2334 3071 2340 3072
rect 2622 3076 2628 3077
rect 2622 3072 2623 3076
rect 2627 3072 2628 3076
rect 2622 3071 2628 3072
rect 2910 3076 2916 3077
rect 2910 3072 2911 3076
rect 2915 3072 2916 3076
rect 2910 3071 2916 3072
rect 3206 3076 3212 3077
rect 3206 3072 3207 3076
rect 3211 3072 3212 3076
rect 3206 3071 3212 3072
rect 3502 3076 3508 3077
rect 3502 3072 3503 3076
rect 3507 3072 3508 3076
rect 3502 3071 3508 3072
rect 3798 3076 3804 3077
rect 3798 3072 3799 3076
rect 3803 3072 3804 3076
rect 3942 3075 3943 3079
rect 3947 3075 3948 3079
rect 3942 3074 3948 3075
rect 3798 3071 3804 3072
rect 2123 3055 2129 3056
rect 2123 3051 2124 3055
rect 2128 3054 2129 3055
rect 2182 3055 2188 3056
rect 2182 3054 2183 3055
rect 2128 3052 2183 3054
rect 2128 3051 2129 3052
rect 2123 3050 2129 3051
rect 2182 3051 2183 3052
rect 2187 3051 2188 3055
rect 2182 3050 2188 3051
rect 2298 3055 2304 3056
rect 2298 3051 2299 3055
rect 2303 3054 2304 3055
rect 2387 3055 2393 3056
rect 2387 3054 2388 3055
rect 2303 3052 2388 3054
rect 2303 3051 2304 3052
rect 2298 3050 2304 3051
rect 2387 3051 2388 3052
rect 2392 3051 2393 3055
rect 2698 3055 2704 3056
rect 2387 3050 2393 3051
rect 2674 3051 2681 3052
rect 2674 3047 2675 3051
rect 2680 3047 2681 3051
rect 2698 3051 2699 3055
rect 2703 3054 2704 3055
rect 2963 3055 2969 3056
rect 2963 3054 2964 3055
rect 2703 3052 2964 3054
rect 2703 3051 2704 3052
rect 2698 3050 2704 3051
rect 2963 3051 2964 3052
rect 2968 3051 2969 3055
rect 2963 3050 2969 3051
rect 2986 3055 2992 3056
rect 2986 3051 2987 3055
rect 2991 3054 2992 3055
rect 3259 3055 3265 3056
rect 3259 3054 3260 3055
rect 2991 3052 3260 3054
rect 2991 3051 2992 3052
rect 2986 3050 2992 3051
rect 3259 3051 3260 3052
rect 3264 3051 3265 3055
rect 3259 3050 3265 3051
rect 3282 3055 3288 3056
rect 3282 3051 3283 3055
rect 3287 3054 3288 3055
rect 3555 3055 3561 3056
rect 3555 3054 3556 3055
rect 3287 3052 3556 3054
rect 3287 3051 3288 3052
rect 3282 3050 3288 3051
rect 3555 3051 3556 3052
rect 3560 3051 3561 3055
rect 3555 3050 3561 3051
rect 3851 3055 3857 3056
rect 3851 3051 3852 3055
rect 3856 3054 3857 3055
rect 3866 3055 3872 3056
rect 3866 3054 3867 3055
rect 3856 3052 3867 3054
rect 3856 3051 3857 3052
rect 3851 3050 3857 3051
rect 3866 3051 3867 3052
rect 3871 3051 3872 3055
rect 3866 3050 3872 3051
rect 2674 3046 2681 3047
rect 110 3040 116 3041
rect 2006 3040 2012 3041
rect 110 3036 111 3040
rect 115 3036 116 3040
rect 110 3035 116 3036
rect 502 3039 508 3040
rect 502 3035 503 3039
rect 507 3035 508 3039
rect 502 3034 508 3035
rect 598 3039 604 3040
rect 598 3035 599 3039
rect 603 3035 604 3039
rect 598 3034 604 3035
rect 702 3039 708 3040
rect 702 3035 703 3039
rect 707 3035 708 3039
rect 702 3034 708 3035
rect 814 3039 820 3040
rect 814 3035 815 3039
rect 819 3035 820 3039
rect 814 3034 820 3035
rect 934 3039 940 3040
rect 934 3035 935 3039
rect 939 3035 940 3039
rect 934 3034 940 3035
rect 1070 3039 1076 3040
rect 1070 3035 1071 3039
rect 1075 3035 1076 3039
rect 1070 3034 1076 3035
rect 1222 3039 1228 3040
rect 1222 3035 1223 3039
rect 1227 3035 1228 3039
rect 1222 3034 1228 3035
rect 1382 3039 1388 3040
rect 1382 3035 1383 3039
rect 1387 3035 1388 3039
rect 1382 3034 1388 3035
rect 1550 3039 1556 3040
rect 1550 3035 1551 3039
rect 1555 3035 1556 3039
rect 1550 3034 1556 3035
rect 1718 3039 1724 3040
rect 1718 3035 1719 3039
rect 1723 3035 1724 3039
rect 2006 3036 2007 3040
rect 2011 3036 2012 3040
rect 2006 3035 2012 3036
rect 2123 3039 2129 3040
rect 2123 3035 2124 3039
rect 2128 3038 2129 3039
rect 2146 3039 2152 3040
rect 2146 3038 2147 3039
rect 2128 3036 2147 3038
rect 2128 3035 2129 3036
rect 1718 3034 1724 3035
rect 2123 3034 2129 3035
rect 2146 3035 2147 3036
rect 2151 3035 2152 3039
rect 2146 3034 2152 3035
rect 2271 3039 2277 3040
rect 2271 3035 2272 3039
rect 2276 3038 2277 3039
rect 2435 3039 2441 3040
rect 2435 3038 2436 3039
rect 2276 3036 2436 3038
rect 2276 3035 2277 3036
rect 2271 3034 2277 3035
rect 2435 3035 2436 3036
rect 2440 3035 2441 3039
rect 2435 3034 2441 3035
rect 2755 3039 2761 3040
rect 2755 3035 2756 3039
rect 2760 3038 2761 3039
rect 2958 3039 2964 3040
rect 2958 3038 2959 3039
rect 2760 3036 2959 3038
rect 2760 3035 2761 3036
rect 2755 3034 2761 3035
rect 2958 3035 2959 3036
rect 2963 3035 2964 3039
rect 2958 3034 2964 3035
rect 3051 3039 3057 3040
rect 3051 3035 3052 3039
rect 3056 3038 3057 3039
rect 3258 3039 3264 3040
rect 3258 3038 3259 3039
rect 3056 3036 3259 3038
rect 3056 3035 3057 3036
rect 3051 3034 3057 3035
rect 3258 3035 3259 3036
rect 3263 3035 3264 3039
rect 3258 3034 3264 3035
rect 3339 3039 3345 3040
rect 3339 3035 3340 3039
rect 3344 3038 3345 3039
rect 3370 3039 3376 3040
rect 3370 3038 3371 3039
rect 3344 3036 3371 3038
rect 3344 3035 3345 3036
rect 3339 3034 3345 3035
rect 3370 3035 3371 3036
rect 3375 3035 3376 3039
rect 3370 3034 3376 3035
rect 3627 3039 3633 3040
rect 3627 3035 3628 3039
rect 3632 3038 3633 3039
rect 3799 3039 3805 3040
rect 3799 3038 3800 3039
rect 3632 3036 3800 3038
rect 3632 3035 3633 3036
rect 3627 3034 3633 3035
rect 3799 3035 3800 3036
rect 3804 3035 3805 3039
rect 3799 3034 3805 3035
rect 3891 3039 3897 3040
rect 3891 3035 3892 3039
rect 3896 3038 3897 3039
rect 3922 3039 3928 3040
rect 3922 3038 3923 3039
rect 3896 3036 3923 3038
rect 3896 3035 3897 3036
rect 3891 3034 3897 3035
rect 3922 3035 3923 3036
rect 3927 3035 3928 3039
rect 3922 3034 3928 3035
rect 366 3031 372 3032
rect 366 3027 367 3031
rect 371 3030 372 3031
rect 586 3031 592 3032
rect 371 3028 545 3030
rect 371 3027 372 3028
rect 366 3026 372 3027
rect 586 3027 587 3031
rect 591 3030 592 3031
rect 682 3031 688 3032
rect 591 3028 641 3030
rect 591 3027 592 3028
rect 586 3026 592 3027
rect 682 3027 683 3031
rect 687 3030 688 3031
rect 806 3031 812 3032
rect 687 3028 745 3030
rect 687 3027 688 3028
rect 682 3026 688 3027
rect 806 3027 807 3031
rect 811 3030 812 3031
rect 902 3031 908 3032
rect 811 3028 857 3030
rect 811 3027 812 3028
rect 806 3026 812 3027
rect 902 3027 903 3031
rect 907 3030 908 3031
rect 1191 3031 1197 3032
rect 907 3028 977 3030
rect 907 3027 908 3028
rect 902 3026 908 3027
rect 1146 3027 1152 3028
rect 110 3023 116 3024
rect 110 3019 111 3023
rect 115 3019 116 3023
rect 1146 3023 1147 3027
rect 1151 3023 1152 3027
rect 1191 3027 1192 3031
rect 1196 3030 1197 3031
rect 1342 3031 1348 3032
rect 1196 3028 1265 3030
rect 1196 3027 1197 3028
rect 1191 3026 1197 3027
rect 1342 3027 1343 3031
rect 1347 3030 1348 3031
rect 1794 3031 1800 3032
rect 1347 3028 1425 3030
rect 1347 3027 1348 3028
rect 1342 3026 1348 3027
rect 1626 3027 1632 3028
rect 1146 3022 1152 3023
rect 1626 3023 1627 3027
rect 1631 3023 1632 3027
rect 1794 3027 1795 3031
rect 1799 3027 1800 3031
rect 1794 3026 1800 3027
rect 1626 3022 1632 3023
rect 2006 3023 2012 3024
rect 110 3018 116 3019
rect 502 3020 508 3021
rect 502 3016 503 3020
rect 507 3016 508 3020
rect 502 3015 508 3016
rect 598 3020 604 3021
rect 598 3016 599 3020
rect 603 3016 604 3020
rect 598 3015 604 3016
rect 702 3020 708 3021
rect 702 3016 703 3020
rect 707 3016 708 3020
rect 702 3015 708 3016
rect 814 3020 820 3021
rect 814 3016 815 3020
rect 819 3016 820 3020
rect 814 3015 820 3016
rect 934 3020 940 3021
rect 934 3016 935 3020
rect 939 3016 940 3020
rect 934 3015 940 3016
rect 1070 3020 1076 3021
rect 1070 3016 1071 3020
rect 1075 3016 1076 3020
rect 1070 3015 1076 3016
rect 1222 3020 1228 3021
rect 1222 3016 1223 3020
rect 1227 3016 1228 3020
rect 1222 3015 1228 3016
rect 1382 3020 1388 3021
rect 1382 3016 1383 3020
rect 1387 3016 1388 3020
rect 1382 3015 1388 3016
rect 1550 3020 1556 3021
rect 1550 3016 1551 3020
rect 1555 3016 1556 3020
rect 1550 3015 1556 3016
rect 1718 3020 1724 3021
rect 1718 3016 1719 3020
rect 1723 3016 1724 3020
rect 2006 3019 2007 3023
rect 2011 3019 2012 3023
rect 2006 3018 2012 3019
rect 1718 3015 1724 3016
rect 2070 3016 2076 3017
rect 2046 3013 2052 3014
rect 2046 3009 2047 3013
rect 2051 3009 2052 3013
rect 2070 3012 2071 3016
rect 2075 3012 2076 3016
rect 2070 3011 2076 3012
rect 2382 3016 2388 3017
rect 2382 3012 2383 3016
rect 2387 3012 2388 3016
rect 2382 3011 2388 3012
rect 2702 3016 2708 3017
rect 2702 3012 2703 3016
rect 2707 3012 2708 3016
rect 2702 3011 2708 3012
rect 2998 3016 3004 3017
rect 2998 3012 2999 3016
rect 3003 3012 3004 3016
rect 2998 3011 3004 3012
rect 3286 3016 3292 3017
rect 3286 3012 3287 3016
rect 3291 3012 3292 3016
rect 3286 3011 3292 3012
rect 3574 3016 3580 3017
rect 3574 3012 3575 3016
rect 3579 3012 3580 3016
rect 3574 3011 3580 3012
rect 3838 3016 3844 3017
rect 3838 3012 3839 3016
rect 3843 3012 3844 3016
rect 3838 3011 3844 3012
rect 3942 3013 3948 3014
rect 2046 3008 2052 3009
rect 3942 3009 3943 3013
rect 3947 3009 3948 3013
rect 3942 3008 3948 3009
rect 2271 3007 2277 3008
rect 2271 3006 2272 3007
rect 2149 3004 2272 3006
rect 2271 3003 2272 3004
rect 2276 3003 2277 3007
rect 2271 3002 2277 3003
rect 2450 3007 2456 3008
rect 2450 3003 2451 3007
rect 2455 3003 2456 3007
rect 2450 3002 2456 3003
rect 2674 3007 2680 3008
rect 2674 3003 2675 3007
rect 2679 3006 2680 3007
rect 2958 3007 2964 3008
rect 2679 3004 2745 3006
rect 2679 3003 2680 3004
rect 2674 3002 2680 3003
rect 2958 3003 2959 3007
rect 2963 3006 2964 3007
rect 3258 3007 3264 3008
rect 2963 3004 3041 3006
rect 2963 3003 2964 3004
rect 2958 3002 2964 3003
rect 3258 3003 3259 3007
rect 3263 3006 3264 3007
rect 3370 3007 3376 3008
rect 3263 3004 3329 3006
rect 3263 3003 3264 3004
rect 3258 3002 3264 3003
rect 3370 3003 3371 3007
rect 3375 3006 3376 3007
rect 3914 3007 3920 3008
rect 3375 3004 3617 3006
rect 3375 3003 3376 3004
rect 3370 3002 3376 3003
rect 3914 3003 3915 3007
rect 3919 3003 3920 3007
rect 3914 3002 3920 3003
rect 555 2999 561 3000
rect 555 2995 556 2999
rect 560 2998 561 2999
rect 586 2999 592 3000
rect 586 2998 587 2999
rect 560 2996 587 2998
rect 560 2995 561 2996
rect 555 2994 561 2995
rect 586 2995 587 2996
rect 591 2995 592 2999
rect 586 2994 592 2995
rect 651 2999 657 3000
rect 651 2995 652 2999
rect 656 2998 657 2999
rect 682 2999 688 3000
rect 682 2998 683 2999
rect 656 2996 683 2998
rect 656 2995 657 2996
rect 651 2994 657 2995
rect 682 2995 683 2996
rect 687 2995 688 2999
rect 682 2994 688 2995
rect 755 2999 761 3000
rect 755 2995 756 2999
rect 760 2998 761 2999
rect 806 2999 812 3000
rect 806 2998 807 2999
rect 760 2996 807 2998
rect 760 2995 761 2996
rect 755 2994 761 2995
rect 806 2995 807 2996
rect 811 2995 812 2999
rect 806 2994 812 2995
rect 867 2999 873 3000
rect 867 2995 868 2999
rect 872 2998 873 2999
rect 902 2999 908 3000
rect 902 2998 903 2999
rect 872 2996 903 2998
rect 872 2995 873 2996
rect 867 2994 873 2995
rect 902 2995 903 2996
rect 907 2995 908 2999
rect 1123 2999 1129 3000
rect 902 2994 908 2995
rect 987 2995 996 2996
rect 987 2991 988 2995
rect 995 2991 996 2995
rect 1123 2995 1124 2999
rect 1128 2998 1129 2999
rect 1191 2999 1197 3000
rect 1191 2998 1192 2999
rect 1128 2996 1192 2998
rect 1128 2995 1129 2996
rect 1123 2994 1129 2995
rect 1191 2995 1192 2996
rect 1196 2995 1197 2999
rect 1191 2994 1197 2995
rect 1275 2999 1281 3000
rect 1275 2995 1276 2999
rect 1280 2998 1281 2999
rect 1342 2999 1348 3000
rect 1342 2998 1343 2999
rect 1280 2996 1343 2998
rect 1280 2995 1281 2996
rect 1275 2994 1281 2995
rect 1342 2995 1343 2996
rect 1347 2995 1348 2999
rect 1342 2994 1348 2995
rect 1350 2999 1356 3000
rect 1350 2995 1351 2999
rect 1355 2998 1356 2999
rect 1435 2999 1441 3000
rect 1435 2998 1436 2999
rect 1355 2996 1436 2998
rect 1355 2995 1356 2996
rect 1350 2994 1356 2995
rect 1435 2995 1436 2996
rect 1440 2995 1441 2999
rect 1626 2999 1632 3000
rect 1435 2994 1441 2995
rect 1562 2995 1568 2996
rect 987 2990 996 2991
rect 1562 2991 1563 2995
rect 1567 2994 1568 2995
rect 1603 2995 1609 2996
rect 1603 2994 1604 2995
rect 1567 2992 1604 2994
rect 1567 2991 1568 2992
rect 1562 2990 1568 2991
rect 1603 2991 1604 2992
rect 1608 2991 1609 2995
rect 1626 2995 1627 2999
rect 1631 2998 1632 2999
rect 1771 2999 1777 3000
rect 1771 2998 1772 2999
rect 1631 2996 1772 2998
rect 1631 2995 1632 2996
rect 1626 2994 1632 2995
rect 1771 2995 1772 2996
rect 1776 2995 1777 2999
rect 2070 2997 2076 2998
rect 1771 2994 1777 2995
rect 2046 2996 2052 2997
rect 2046 2992 2047 2996
rect 2051 2992 2052 2996
rect 2070 2993 2071 2997
rect 2075 2993 2076 2997
rect 2070 2992 2076 2993
rect 2382 2997 2388 2998
rect 2382 2993 2383 2997
rect 2387 2993 2388 2997
rect 2382 2992 2388 2993
rect 2702 2997 2708 2998
rect 2702 2993 2703 2997
rect 2707 2993 2708 2997
rect 2702 2992 2708 2993
rect 2998 2997 3004 2998
rect 2998 2993 2999 2997
rect 3003 2993 3004 2997
rect 2998 2992 3004 2993
rect 3286 2997 3292 2998
rect 3286 2993 3287 2997
rect 3291 2993 3292 2997
rect 3286 2992 3292 2993
rect 3574 2997 3580 2998
rect 3574 2993 3575 2997
rect 3579 2993 3580 2997
rect 3574 2992 3580 2993
rect 3838 2997 3844 2998
rect 3838 2993 3839 2997
rect 3843 2993 3844 2997
rect 3838 2992 3844 2993
rect 3942 2996 3948 2997
rect 3942 2992 3943 2996
rect 3947 2992 3948 2996
rect 2046 2991 2052 2992
rect 3942 2991 3948 2992
rect 1603 2990 1609 2991
rect 626 2979 632 2980
rect 603 2977 609 2978
rect 603 2973 604 2977
rect 608 2973 609 2977
rect 626 2975 627 2979
rect 631 2978 632 2979
rect 699 2979 705 2980
rect 699 2978 700 2979
rect 631 2976 700 2978
rect 631 2975 632 2976
rect 626 2974 632 2975
rect 699 2975 700 2976
rect 704 2975 705 2979
rect 699 2974 705 2975
rect 722 2979 728 2980
rect 722 2975 723 2979
rect 727 2978 728 2979
rect 811 2979 817 2980
rect 811 2978 812 2979
rect 727 2976 812 2978
rect 727 2975 728 2976
rect 722 2974 728 2975
rect 811 2975 812 2976
rect 816 2975 817 2979
rect 811 2974 817 2975
rect 834 2979 840 2980
rect 834 2975 835 2979
rect 839 2978 840 2979
rect 939 2979 945 2980
rect 939 2978 940 2979
rect 839 2976 940 2978
rect 839 2975 840 2976
rect 834 2974 840 2975
rect 939 2975 940 2976
rect 944 2975 945 2979
rect 939 2974 945 2975
rect 962 2979 968 2980
rect 962 2975 963 2979
rect 967 2978 968 2979
rect 1075 2979 1081 2980
rect 1075 2978 1076 2979
rect 967 2976 1076 2978
rect 967 2975 968 2976
rect 962 2974 968 2975
rect 1075 2975 1076 2976
rect 1080 2975 1081 2979
rect 1075 2974 1081 2975
rect 1146 2979 1152 2980
rect 1146 2975 1147 2979
rect 1151 2978 1152 2979
rect 1227 2979 1233 2980
rect 1227 2978 1228 2979
rect 1151 2976 1228 2978
rect 1151 2975 1152 2976
rect 1146 2974 1152 2975
rect 1227 2975 1228 2976
rect 1232 2975 1233 2979
rect 1227 2974 1233 2975
rect 1250 2979 1256 2980
rect 1250 2975 1251 2979
rect 1255 2978 1256 2979
rect 1379 2979 1385 2980
rect 1379 2978 1380 2979
rect 1255 2976 1380 2978
rect 1255 2975 1256 2976
rect 1250 2974 1256 2975
rect 1379 2975 1380 2976
rect 1384 2975 1385 2979
rect 1379 2974 1385 2975
rect 1539 2979 1545 2980
rect 1539 2975 1540 2979
rect 1544 2978 1545 2979
rect 1570 2979 1576 2980
rect 1570 2978 1571 2979
rect 1544 2976 1571 2978
rect 1544 2975 1545 2976
rect 1539 2974 1545 2975
rect 1570 2975 1571 2976
rect 1575 2975 1576 2979
rect 1570 2974 1576 2975
rect 1707 2979 1713 2980
rect 1707 2975 1708 2979
rect 1712 2978 1713 2979
rect 1738 2979 1744 2980
rect 1738 2978 1739 2979
rect 1712 2976 1739 2978
rect 1712 2975 1713 2976
rect 1707 2974 1713 2975
rect 1738 2975 1739 2976
rect 1743 2975 1744 2979
rect 1738 2974 1744 2975
rect 1875 2979 1881 2980
rect 1875 2975 1876 2979
rect 1880 2978 1881 2979
rect 1922 2979 1928 2980
rect 1922 2978 1923 2979
rect 1880 2976 1923 2978
rect 1880 2975 1881 2976
rect 1875 2974 1881 2975
rect 1922 2975 1923 2976
rect 1927 2975 1928 2979
rect 1922 2974 1928 2975
rect 603 2972 609 2973
rect 604 2970 606 2972
rect 922 2971 928 2972
rect 922 2970 923 2971
rect 604 2968 923 2970
rect 922 2967 923 2968
rect 927 2967 928 2971
rect 922 2966 928 2967
rect 550 2956 556 2957
rect 110 2953 116 2954
rect 110 2949 111 2953
rect 115 2949 116 2953
rect 550 2952 551 2956
rect 555 2952 556 2956
rect 550 2951 556 2952
rect 646 2956 652 2957
rect 646 2952 647 2956
rect 651 2952 652 2956
rect 646 2951 652 2952
rect 758 2956 764 2957
rect 758 2952 759 2956
rect 763 2952 764 2956
rect 758 2951 764 2952
rect 886 2956 892 2957
rect 886 2952 887 2956
rect 891 2952 892 2956
rect 886 2951 892 2952
rect 1022 2956 1028 2957
rect 1022 2952 1023 2956
rect 1027 2952 1028 2956
rect 1022 2951 1028 2952
rect 1174 2956 1180 2957
rect 1174 2952 1175 2956
rect 1179 2952 1180 2956
rect 1174 2951 1180 2952
rect 1326 2956 1332 2957
rect 1326 2952 1327 2956
rect 1331 2952 1332 2956
rect 1326 2951 1332 2952
rect 1486 2956 1492 2957
rect 1486 2952 1487 2956
rect 1491 2952 1492 2956
rect 1486 2951 1492 2952
rect 1654 2956 1660 2957
rect 1654 2952 1655 2956
rect 1659 2952 1660 2956
rect 1654 2951 1660 2952
rect 1822 2956 1828 2957
rect 1822 2952 1823 2956
rect 1827 2952 1828 2956
rect 1822 2951 1828 2952
rect 2006 2953 2012 2954
rect 110 2948 116 2949
rect 2006 2949 2007 2953
rect 2011 2949 2012 2953
rect 2006 2948 2012 2949
rect 626 2947 632 2948
rect 626 2943 627 2947
rect 631 2943 632 2947
rect 626 2942 632 2943
rect 722 2947 728 2948
rect 722 2943 723 2947
rect 727 2943 728 2947
rect 722 2942 728 2943
rect 834 2947 840 2948
rect 834 2943 835 2947
rect 839 2943 840 2947
rect 834 2942 840 2943
rect 962 2947 968 2948
rect 962 2943 963 2947
rect 967 2943 968 2947
rect 962 2942 968 2943
rect 990 2947 996 2948
rect 990 2943 991 2947
rect 995 2946 996 2947
rect 1250 2947 1256 2948
rect 995 2944 1065 2946
rect 995 2943 996 2944
rect 990 2942 996 2943
rect 1250 2943 1251 2947
rect 1255 2943 1256 2947
rect 1250 2942 1256 2943
rect 1287 2947 1293 2948
rect 1287 2943 1288 2947
rect 1292 2946 1293 2947
rect 1562 2947 1568 2948
rect 1292 2944 1369 2946
rect 1292 2943 1293 2944
rect 1287 2942 1293 2943
rect 1562 2943 1563 2947
rect 1567 2943 1568 2947
rect 1562 2942 1568 2943
rect 1570 2947 1576 2948
rect 1570 2943 1571 2947
rect 1575 2946 1576 2947
rect 1738 2947 1744 2948
rect 1575 2944 1697 2946
rect 1575 2943 1576 2944
rect 1570 2942 1576 2943
rect 1738 2943 1739 2947
rect 1743 2946 1744 2947
rect 1743 2944 1865 2946
rect 1743 2943 1744 2944
rect 1738 2942 1744 2943
rect 2046 2940 2052 2941
rect 3942 2940 3948 2941
rect 550 2937 556 2938
rect 110 2936 116 2937
rect 110 2932 111 2936
rect 115 2932 116 2936
rect 550 2933 551 2937
rect 555 2933 556 2937
rect 550 2932 556 2933
rect 646 2937 652 2938
rect 646 2933 647 2937
rect 651 2933 652 2937
rect 646 2932 652 2933
rect 758 2937 764 2938
rect 758 2933 759 2937
rect 763 2933 764 2937
rect 758 2932 764 2933
rect 886 2937 892 2938
rect 886 2933 887 2937
rect 891 2933 892 2937
rect 886 2932 892 2933
rect 1022 2937 1028 2938
rect 1022 2933 1023 2937
rect 1027 2933 1028 2937
rect 1022 2932 1028 2933
rect 1174 2937 1180 2938
rect 1174 2933 1175 2937
rect 1179 2933 1180 2937
rect 1174 2932 1180 2933
rect 1326 2937 1332 2938
rect 1326 2933 1327 2937
rect 1331 2933 1332 2937
rect 1326 2932 1332 2933
rect 1486 2937 1492 2938
rect 1486 2933 1487 2937
rect 1491 2933 1492 2937
rect 1486 2932 1492 2933
rect 1654 2937 1660 2938
rect 1654 2933 1655 2937
rect 1659 2933 1660 2937
rect 1654 2932 1660 2933
rect 1822 2937 1828 2938
rect 1822 2933 1823 2937
rect 1827 2933 1828 2937
rect 1822 2932 1828 2933
rect 2006 2936 2012 2937
rect 2006 2932 2007 2936
rect 2011 2932 2012 2936
rect 2046 2936 2047 2940
rect 2051 2936 2052 2940
rect 2046 2935 2052 2936
rect 2070 2939 2076 2940
rect 2070 2935 2071 2939
rect 2075 2935 2076 2939
rect 2070 2934 2076 2935
rect 2390 2939 2396 2940
rect 2390 2935 2391 2939
rect 2395 2935 2396 2939
rect 2390 2934 2396 2935
rect 2702 2939 2708 2940
rect 2702 2935 2703 2939
rect 2707 2935 2708 2939
rect 2702 2934 2708 2935
rect 2974 2939 2980 2940
rect 2974 2935 2975 2939
rect 2979 2935 2980 2939
rect 2974 2934 2980 2935
rect 3214 2939 3220 2940
rect 3214 2935 3215 2939
rect 3219 2935 3220 2939
rect 3214 2934 3220 2935
rect 3438 2939 3444 2940
rect 3438 2935 3439 2939
rect 3443 2935 3444 2939
rect 3438 2934 3444 2935
rect 3646 2939 3652 2940
rect 3646 2935 3647 2939
rect 3651 2935 3652 2939
rect 3646 2934 3652 2935
rect 3838 2939 3844 2940
rect 3838 2935 3839 2939
rect 3843 2935 3844 2939
rect 3942 2936 3943 2940
rect 3947 2936 3948 2940
rect 3942 2935 3948 2936
rect 3838 2934 3844 2935
rect 110 2931 116 2932
rect 2006 2931 2012 2932
rect 2279 2931 2285 2932
rect 2146 2927 2152 2928
rect 2046 2923 2052 2924
rect 2046 2919 2047 2923
rect 2051 2919 2052 2923
rect 2146 2923 2147 2927
rect 2151 2923 2152 2927
rect 2279 2927 2280 2931
rect 2284 2930 2285 2931
rect 3799 2931 3805 2932
rect 2284 2928 2433 2930
rect 2284 2927 2285 2928
rect 2279 2926 2285 2927
rect 2778 2927 2784 2928
rect 2146 2922 2152 2923
rect 2778 2923 2779 2927
rect 2783 2923 2784 2927
rect 2778 2922 2784 2923
rect 3050 2927 3056 2928
rect 3050 2923 3051 2927
rect 3055 2923 3056 2927
rect 3050 2922 3056 2923
rect 3290 2927 3296 2928
rect 3290 2923 3291 2927
rect 3295 2923 3296 2927
rect 3290 2922 3296 2923
rect 3514 2927 3520 2928
rect 3514 2923 3515 2927
rect 3519 2923 3520 2927
rect 3514 2922 3520 2923
rect 3722 2927 3728 2928
rect 3722 2923 3723 2927
rect 3727 2923 3728 2927
rect 3799 2927 3800 2931
rect 3804 2930 3805 2931
rect 3804 2928 3881 2930
rect 3804 2927 3805 2928
rect 3799 2926 3805 2927
rect 3722 2922 3728 2923
rect 3942 2923 3948 2924
rect 2046 2918 2052 2919
rect 2070 2920 2076 2921
rect 2070 2916 2071 2920
rect 2075 2916 2076 2920
rect 2070 2915 2076 2916
rect 2390 2920 2396 2921
rect 2390 2916 2391 2920
rect 2395 2916 2396 2920
rect 2390 2915 2396 2916
rect 2702 2920 2708 2921
rect 2702 2916 2703 2920
rect 2707 2916 2708 2920
rect 2702 2915 2708 2916
rect 2974 2920 2980 2921
rect 2974 2916 2975 2920
rect 2979 2916 2980 2920
rect 2974 2915 2980 2916
rect 3214 2920 3220 2921
rect 3214 2916 3215 2920
rect 3219 2916 3220 2920
rect 3214 2915 3220 2916
rect 3438 2920 3444 2921
rect 3438 2916 3439 2920
rect 3443 2916 3444 2920
rect 3438 2915 3444 2916
rect 3646 2920 3652 2921
rect 3646 2916 3647 2920
rect 3651 2916 3652 2920
rect 3646 2915 3652 2916
rect 3838 2920 3844 2921
rect 3838 2916 3839 2920
rect 3843 2916 3844 2920
rect 3942 2919 3943 2923
rect 3947 2919 3948 2923
rect 3942 2918 3948 2919
rect 3838 2915 3844 2916
rect 3618 2907 3624 2908
rect 3618 2906 3619 2907
rect 2839 2904 3619 2906
rect 2123 2899 2129 2900
rect 2123 2895 2124 2899
rect 2128 2898 2129 2899
rect 2279 2899 2285 2900
rect 2279 2898 2280 2899
rect 2128 2896 2280 2898
rect 2128 2895 2129 2896
rect 2123 2894 2129 2895
rect 2279 2895 2280 2896
rect 2284 2895 2285 2899
rect 2279 2894 2285 2895
rect 2443 2899 2452 2900
rect 2443 2895 2444 2899
rect 2451 2895 2452 2899
rect 2443 2894 2452 2895
rect 2755 2899 2761 2900
rect 2755 2895 2756 2899
rect 2760 2898 2761 2899
rect 2839 2898 2841 2904
rect 3618 2903 3619 2904
rect 3623 2903 3624 2907
rect 3618 2902 3624 2903
rect 2760 2896 2841 2898
rect 3050 2899 3056 2900
rect 2760 2895 2761 2896
rect 2755 2894 2761 2895
rect 3027 2895 3033 2896
rect 3027 2894 3028 2895
rect 2839 2892 3028 2894
rect 2778 2891 2784 2892
rect 2778 2887 2779 2891
rect 2783 2890 2784 2891
rect 2839 2890 2841 2892
rect 3027 2891 3028 2892
rect 3032 2891 3033 2895
rect 3050 2895 3051 2899
rect 3055 2898 3056 2899
rect 3267 2899 3273 2900
rect 3267 2898 3268 2899
rect 3055 2896 3268 2898
rect 3055 2895 3056 2896
rect 3050 2894 3056 2895
rect 3267 2895 3268 2896
rect 3272 2895 3273 2899
rect 3267 2894 3273 2895
rect 3290 2899 3296 2900
rect 3290 2895 3291 2899
rect 3295 2898 3296 2899
rect 3491 2899 3497 2900
rect 3491 2898 3492 2899
rect 3295 2896 3492 2898
rect 3295 2895 3296 2896
rect 3290 2894 3296 2895
rect 3491 2895 3492 2896
rect 3496 2895 3497 2899
rect 3491 2894 3497 2895
rect 3514 2899 3520 2900
rect 3514 2895 3515 2899
rect 3519 2898 3520 2899
rect 3699 2899 3705 2900
rect 3699 2898 3700 2899
rect 3519 2896 3700 2898
rect 3519 2895 3520 2896
rect 3514 2894 3520 2895
rect 3699 2895 3700 2896
rect 3704 2895 3705 2899
rect 3699 2894 3705 2895
rect 3722 2899 3728 2900
rect 3722 2895 3723 2899
rect 3727 2898 3728 2899
rect 3891 2899 3897 2900
rect 3891 2898 3892 2899
rect 3727 2896 3892 2898
rect 3727 2895 3728 2896
rect 3722 2894 3728 2895
rect 3891 2895 3892 2896
rect 3896 2895 3897 2899
rect 3891 2894 3897 2895
rect 3027 2890 3033 2891
rect 2783 2888 2841 2890
rect 2783 2887 2784 2888
rect 2778 2886 2784 2887
rect 2123 2883 2129 2884
rect 2123 2879 2124 2883
rect 2128 2882 2129 2883
rect 2146 2883 2152 2884
rect 2146 2882 2147 2883
rect 2128 2880 2147 2882
rect 2128 2879 2129 2880
rect 2123 2878 2129 2879
rect 2146 2879 2147 2880
rect 2151 2879 2152 2883
rect 2146 2878 2152 2879
rect 2230 2883 2236 2884
rect 2230 2879 2231 2883
rect 2235 2882 2236 2883
rect 2347 2883 2353 2884
rect 2347 2882 2348 2883
rect 2235 2880 2348 2882
rect 2235 2879 2236 2880
rect 2230 2878 2236 2879
rect 2347 2879 2348 2880
rect 2352 2879 2353 2883
rect 2347 2878 2353 2879
rect 2370 2883 2376 2884
rect 2370 2879 2371 2883
rect 2375 2882 2376 2883
rect 2587 2883 2593 2884
rect 2587 2882 2588 2883
rect 2375 2880 2588 2882
rect 2375 2879 2376 2880
rect 2370 2878 2376 2879
rect 2587 2879 2588 2880
rect 2592 2879 2593 2883
rect 2587 2878 2593 2879
rect 2610 2883 2616 2884
rect 2610 2879 2611 2883
rect 2615 2882 2616 2883
rect 2819 2883 2825 2884
rect 2819 2882 2820 2883
rect 2615 2880 2820 2882
rect 2615 2879 2616 2880
rect 2610 2878 2616 2879
rect 2819 2879 2820 2880
rect 2824 2879 2825 2883
rect 3066 2883 3072 2884
rect 2819 2878 2825 2879
rect 3043 2881 3049 2882
rect 3043 2877 3044 2881
rect 3048 2877 3049 2881
rect 3066 2879 3067 2883
rect 3071 2882 3072 2883
rect 3267 2883 3273 2884
rect 3267 2882 3268 2883
rect 3071 2880 3268 2882
rect 3071 2879 3072 2880
rect 3066 2878 3072 2879
rect 3267 2879 3268 2880
rect 3272 2879 3273 2883
rect 3267 2878 3273 2879
rect 3290 2883 3296 2884
rect 3290 2879 3291 2883
rect 3295 2882 3296 2883
rect 3483 2883 3489 2884
rect 3483 2882 3484 2883
rect 3295 2880 3484 2882
rect 3295 2879 3296 2880
rect 3290 2878 3296 2879
rect 3483 2879 3484 2880
rect 3488 2879 3489 2883
rect 3483 2878 3489 2879
rect 3506 2883 3512 2884
rect 3506 2879 3507 2883
rect 3511 2882 3512 2883
rect 3699 2883 3705 2884
rect 3699 2882 3700 2883
rect 3511 2880 3700 2882
rect 3511 2879 3512 2880
rect 3506 2878 3512 2879
rect 3699 2879 3700 2880
rect 3704 2879 3705 2883
rect 3699 2878 3705 2879
rect 3891 2883 3897 2884
rect 3891 2879 3892 2883
rect 3896 2882 3897 2883
rect 3906 2883 3912 2884
rect 3906 2882 3907 2883
rect 3896 2880 3907 2882
rect 3896 2879 3897 2880
rect 3891 2878 3897 2879
rect 3906 2879 3907 2880
rect 3911 2879 3912 2883
rect 3906 2878 3912 2879
rect 110 2876 116 2877
rect 2006 2876 2012 2877
rect 3043 2876 3049 2877
rect 110 2872 111 2876
rect 115 2872 116 2876
rect 110 2871 116 2872
rect 470 2875 476 2876
rect 470 2871 471 2875
rect 475 2871 476 2875
rect 470 2870 476 2871
rect 574 2875 580 2876
rect 574 2871 575 2875
rect 579 2871 580 2875
rect 574 2870 580 2871
rect 694 2875 700 2876
rect 694 2871 695 2875
rect 699 2871 700 2875
rect 694 2870 700 2871
rect 838 2875 844 2876
rect 838 2871 839 2875
rect 843 2871 844 2875
rect 838 2870 844 2871
rect 990 2875 996 2876
rect 990 2871 991 2875
rect 995 2871 996 2875
rect 990 2870 996 2871
rect 1150 2875 1156 2876
rect 1150 2871 1151 2875
rect 1155 2871 1156 2875
rect 1150 2870 1156 2871
rect 1318 2875 1324 2876
rect 1318 2871 1319 2875
rect 1323 2871 1324 2875
rect 1318 2870 1324 2871
rect 1494 2875 1500 2876
rect 1494 2871 1495 2875
rect 1499 2871 1500 2875
rect 1494 2870 1500 2871
rect 1670 2875 1676 2876
rect 1670 2871 1671 2875
rect 1675 2871 1676 2875
rect 1670 2870 1676 2871
rect 1846 2875 1852 2876
rect 1846 2871 1847 2875
rect 1851 2871 1852 2875
rect 2006 2872 2007 2876
rect 2011 2872 2012 2876
rect 3044 2874 3046 2876
rect 3438 2875 3444 2876
rect 3438 2874 3439 2875
rect 3044 2872 3439 2874
rect 2006 2871 2012 2872
rect 3438 2871 3439 2872
rect 3443 2871 3444 2875
rect 1846 2870 1852 2871
rect 3438 2870 3444 2871
rect 922 2867 928 2868
rect 566 2863 572 2864
rect 566 2862 567 2863
rect 549 2860 567 2862
rect 110 2859 116 2860
rect 110 2855 111 2859
rect 115 2855 116 2859
rect 566 2859 567 2860
rect 571 2859 572 2863
rect 566 2858 572 2859
rect 650 2863 656 2864
rect 650 2859 651 2863
rect 655 2859 656 2863
rect 650 2858 656 2859
rect 770 2863 776 2864
rect 770 2859 771 2863
rect 775 2859 776 2863
rect 770 2858 776 2859
rect 914 2863 920 2864
rect 914 2859 915 2863
rect 919 2859 920 2863
rect 922 2863 923 2867
rect 927 2866 928 2867
rect 1922 2867 1928 2868
rect 927 2864 1033 2866
rect 927 2863 928 2864
rect 922 2862 928 2863
rect 1226 2863 1232 2864
rect 914 2858 920 2859
rect 1226 2859 1227 2863
rect 1231 2859 1232 2863
rect 1226 2858 1232 2859
rect 1394 2863 1400 2864
rect 1394 2859 1395 2863
rect 1399 2859 1400 2863
rect 1630 2863 1636 2864
rect 1630 2862 1631 2863
rect 1573 2860 1631 2862
rect 1394 2858 1400 2859
rect 1630 2859 1631 2860
rect 1635 2859 1636 2863
rect 1630 2858 1636 2859
rect 1746 2863 1752 2864
rect 1746 2859 1747 2863
rect 1751 2859 1752 2863
rect 1922 2863 1923 2867
rect 1927 2863 1928 2867
rect 1922 2862 1928 2863
rect 2070 2860 2076 2861
rect 1746 2858 1752 2859
rect 2006 2859 2012 2860
rect 110 2854 116 2855
rect 470 2856 476 2857
rect 470 2852 471 2856
rect 475 2852 476 2856
rect 470 2851 476 2852
rect 574 2856 580 2857
rect 574 2852 575 2856
rect 579 2852 580 2856
rect 574 2851 580 2852
rect 694 2856 700 2857
rect 694 2852 695 2856
rect 699 2852 700 2856
rect 694 2851 700 2852
rect 838 2856 844 2857
rect 838 2852 839 2856
rect 843 2852 844 2856
rect 838 2851 844 2852
rect 990 2856 996 2857
rect 990 2852 991 2856
rect 995 2852 996 2856
rect 990 2851 996 2852
rect 1150 2856 1156 2857
rect 1150 2852 1151 2856
rect 1155 2852 1156 2856
rect 1150 2851 1156 2852
rect 1318 2856 1324 2857
rect 1318 2852 1319 2856
rect 1323 2852 1324 2856
rect 1318 2851 1324 2852
rect 1494 2856 1500 2857
rect 1494 2852 1495 2856
rect 1499 2852 1500 2856
rect 1494 2851 1500 2852
rect 1670 2856 1676 2857
rect 1670 2852 1671 2856
rect 1675 2852 1676 2856
rect 1670 2851 1676 2852
rect 1846 2856 1852 2857
rect 1846 2852 1847 2856
rect 1851 2852 1852 2856
rect 2006 2855 2007 2859
rect 2011 2855 2012 2859
rect 2006 2854 2012 2855
rect 2046 2857 2052 2858
rect 2046 2853 2047 2857
rect 2051 2853 2052 2857
rect 2070 2856 2071 2860
rect 2075 2856 2076 2860
rect 2070 2855 2076 2856
rect 2294 2860 2300 2861
rect 2294 2856 2295 2860
rect 2299 2856 2300 2860
rect 2294 2855 2300 2856
rect 2534 2860 2540 2861
rect 2534 2856 2535 2860
rect 2539 2856 2540 2860
rect 2534 2855 2540 2856
rect 2766 2860 2772 2861
rect 2766 2856 2767 2860
rect 2771 2856 2772 2860
rect 2766 2855 2772 2856
rect 2990 2860 2996 2861
rect 2990 2856 2991 2860
rect 2995 2856 2996 2860
rect 2990 2855 2996 2856
rect 3214 2860 3220 2861
rect 3214 2856 3215 2860
rect 3219 2856 3220 2860
rect 3214 2855 3220 2856
rect 3430 2860 3436 2861
rect 3430 2856 3431 2860
rect 3435 2856 3436 2860
rect 3430 2855 3436 2856
rect 3646 2860 3652 2861
rect 3646 2856 3647 2860
rect 3651 2856 3652 2860
rect 3646 2855 3652 2856
rect 3838 2860 3844 2861
rect 3838 2856 3839 2860
rect 3843 2856 3844 2860
rect 3838 2855 3844 2856
rect 3942 2857 3948 2858
rect 2046 2852 2052 2853
rect 3942 2853 3943 2857
rect 3947 2853 3948 2857
rect 3942 2852 3948 2853
rect 1846 2851 1852 2852
rect 2230 2851 2236 2852
rect 2230 2850 2231 2851
rect 2149 2848 2231 2850
rect 2230 2847 2231 2848
rect 2235 2847 2236 2851
rect 2230 2846 2236 2847
rect 2370 2851 2376 2852
rect 2370 2847 2371 2851
rect 2375 2847 2376 2851
rect 2370 2846 2376 2847
rect 2610 2851 2616 2852
rect 2610 2847 2611 2851
rect 2615 2847 2616 2851
rect 2610 2846 2616 2847
rect 2718 2851 2724 2852
rect 2718 2847 2719 2851
rect 2723 2850 2724 2851
rect 3066 2851 3072 2852
rect 2723 2848 2809 2850
rect 2723 2847 2724 2848
rect 2718 2846 2724 2847
rect 3066 2847 3067 2851
rect 3071 2847 3072 2851
rect 3066 2846 3072 2847
rect 3290 2851 3296 2852
rect 3290 2847 3291 2851
rect 3295 2847 3296 2851
rect 3290 2846 3296 2847
rect 3506 2851 3512 2852
rect 3506 2847 3507 2851
rect 3511 2847 3512 2851
rect 3506 2846 3512 2847
rect 3618 2851 3624 2852
rect 3618 2847 3619 2851
rect 3623 2850 3624 2851
rect 3922 2851 3928 2852
rect 3922 2850 3923 2851
rect 3623 2848 3689 2850
rect 3917 2848 3923 2850
rect 3623 2847 3624 2848
rect 3618 2846 3624 2847
rect 3922 2847 3923 2848
rect 3927 2847 3928 2851
rect 3922 2846 3928 2847
rect 1287 2843 1293 2844
rect 1287 2842 1288 2843
rect 1220 2840 1288 2842
rect 566 2835 572 2836
rect 523 2831 529 2832
rect 523 2827 524 2831
rect 528 2830 529 2831
rect 546 2831 552 2832
rect 546 2830 547 2831
rect 528 2828 547 2830
rect 528 2827 529 2828
rect 523 2826 529 2827
rect 546 2827 547 2828
rect 551 2827 552 2831
rect 566 2831 567 2835
rect 571 2834 572 2835
rect 627 2835 633 2836
rect 627 2834 628 2835
rect 571 2832 628 2834
rect 571 2831 572 2832
rect 566 2830 572 2831
rect 627 2831 628 2832
rect 632 2831 633 2835
rect 627 2830 633 2831
rect 650 2835 656 2836
rect 650 2831 651 2835
rect 655 2834 656 2835
rect 747 2835 753 2836
rect 747 2834 748 2835
rect 655 2832 748 2834
rect 655 2831 656 2832
rect 650 2830 656 2831
rect 747 2831 748 2832
rect 752 2831 753 2835
rect 747 2830 753 2831
rect 770 2835 776 2836
rect 770 2831 771 2835
rect 775 2834 776 2835
rect 891 2835 897 2836
rect 891 2834 892 2835
rect 775 2832 892 2834
rect 775 2831 776 2832
rect 770 2830 776 2831
rect 891 2831 892 2832
rect 896 2831 897 2835
rect 891 2830 897 2831
rect 914 2835 920 2836
rect 914 2831 915 2835
rect 919 2834 920 2835
rect 1043 2835 1049 2836
rect 1043 2834 1044 2835
rect 919 2832 1044 2834
rect 919 2831 920 2832
rect 914 2830 920 2831
rect 1043 2831 1044 2832
rect 1048 2831 1049 2835
rect 1043 2830 1049 2831
rect 1203 2835 1209 2836
rect 1203 2831 1204 2835
rect 1208 2834 1209 2835
rect 1220 2834 1222 2840
rect 1287 2839 1288 2840
rect 1292 2839 1293 2843
rect 2070 2841 2076 2842
rect 1287 2838 1293 2839
rect 2046 2840 2052 2841
rect 2046 2836 2047 2840
rect 2051 2836 2052 2840
rect 2070 2837 2071 2841
rect 2075 2837 2076 2841
rect 2070 2836 2076 2837
rect 2294 2841 2300 2842
rect 2294 2837 2295 2841
rect 2299 2837 2300 2841
rect 2294 2836 2300 2837
rect 2534 2841 2540 2842
rect 2534 2837 2535 2841
rect 2539 2837 2540 2841
rect 2534 2836 2540 2837
rect 2766 2841 2772 2842
rect 2766 2837 2767 2841
rect 2771 2837 2772 2841
rect 2766 2836 2772 2837
rect 2990 2841 2996 2842
rect 2990 2837 2991 2841
rect 2995 2837 2996 2841
rect 2990 2836 2996 2837
rect 3214 2841 3220 2842
rect 3214 2837 3215 2841
rect 3219 2837 3220 2841
rect 3214 2836 3220 2837
rect 3430 2841 3436 2842
rect 3430 2837 3431 2841
rect 3435 2837 3436 2841
rect 3430 2836 3436 2837
rect 3646 2841 3652 2842
rect 3646 2837 3647 2841
rect 3651 2837 3652 2841
rect 3646 2836 3652 2837
rect 3838 2841 3844 2842
rect 3838 2837 3839 2841
rect 3843 2837 3844 2841
rect 3838 2836 3844 2837
rect 3942 2840 3948 2841
rect 3942 2836 3943 2840
rect 3947 2836 3948 2840
rect 1208 2832 1222 2834
rect 1226 2835 1232 2836
rect 1208 2831 1209 2832
rect 1203 2830 1209 2831
rect 1226 2831 1227 2835
rect 1231 2834 1232 2835
rect 1371 2835 1377 2836
rect 1371 2834 1372 2835
rect 1231 2832 1372 2834
rect 1231 2831 1232 2832
rect 1226 2830 1232 2831
rect 1371 2831 1372 2832
rect 1376 2831 1377 2835
rect 1630 2835 1636 2836
rect 1371 2830 1377 2831
rect 1547 2831 1556 2832
rect 546 2826 552 2827
rect 1547 2827 1548 2831
rect 1555 2827 1556 2831
rect 1630 2831 1631 2835
rect 1635 2834 1636 2835
rect 1723 2835 1729 2836
rect 1723 2834 1724 2835
rect 1635 2832 1724 2834
rect 1635 2831 1636 2832
rect 1630 2830 1636 2831
rect 1723 2831 1724 2832
rect 1728 2831 1729 2835
rect 1723 2830 1729 2831
rect 1746 2835 1752 2836
rect 1746 2831 1747 2835
rect 1751 2834 1752 2835
rect 1899 2835 1905 2836
rect 2046 2835 2052 2836
rect 3942 2835 3948 2836
rect 1899 2834 1900 2835
rect 1751 2832 1900 2834
rect 1751 2831 1752 2832
rect 1746 2830 1752 2831
rect 1899 2831 1900 2832
rect 1904 2831 1905 2835
rect 1899 2830 1905 2831
rect 1547 2826 1556 2827
rect 531 2815 537 2816
rect 531 2811 532 2815
rect 536 2814 537 2815
rect 562 2815 568 2816
rect 562 2814 563 2815
rect 536 2812 563 2814
rect 536 2811 537 2812
rect 531 2810 537 2811
rect 562 2811 563 2812
rect 567 2811 568 2815
rect 562 2810 568 2811
rect 627 2815 633 2816
rect 627 2811 628 2815
rect 632 2814 633 2815
rect 658 2815 664 2816
rect 658 2814 659 2815
rect 632 2812 659 2814
rect 632 2811 633 2812
rect 627 2810 633 2811
rect 658 2811 659 2812
rect 663 2811 664 2815
rect 658 2810 664 2811
rect 731 2815 737 2816
rect 731 2811 732 2815
rect 736 2814 737 2815
rect 762 2815 768 2816
rect 762 2814 763 2815
rect 736 2812 763 2814
rect 736 2811 737 2812
rect 731 2810 737 2811
rect 762 2811 763 2812
rect 767 2811 768 2815
rect 762 2810 768 2811
rect 851 2815 857 2816
rect 851 2811 852 2815
rect 856 2814 857 2815
rect 882 2815 888 2816
rect 882 2814 883 2815
rect 856 2812 883 2814
rect 856 2811 857 2812
rect 851 2810 857 2811
rect 882 2811 883 2812
rect 887 2811 888 2815
rect 882 2810 888 2811
rect 987 2815 993 2816
rect 987 2811 988 2815
rect 992 2814 993 2815
rect 998 2815 1004 2816
rect 998 2814 999 2815
rect 992 2812 999 2814
rect 992 2811 993 2812
rect 987 2810 993 2811
rect 998 2811 999 2812
rect 1003 2811 1004 2815
rect 998 2810 1004 2811
rect 1131 2815 1137 2816
rect 1131 2811 1132 2815
rect 1136 2814 1137 2815
rect 1190 2815 1196 2816
rect 1190 2814 1191 2815
rect 1136 2812 1191 2814
rect 1136 2811 1137 2812
rect 1131 2810 1137 2811
rect 1190 2811 1191 2812
rect 1195 2811 1196 2815
rect 1190 2810 1196 2811
rect 1291 2815 1297 2816
rect 1291 2811 1292 2815
rect 1296 2814 1297 2815
rect 1326 2815 1332 2816
rect 1326 2814 1327 2815
rect 1296 2812 1327 2814
rect 1296 2811 1297 2812
rect 1291 2810 1297 2811
rect 1326 2811 1327 2812
rect 1331 2811 1332 2815
rect 1326 2810 1332 2811
rect 1394 2815 1400 2816
rect 1394 2811 1395 2815
rect 1399 2814 1400 2815
rect 1467 2815 1473 2816
rect 1467 2814 1468 2815
rect 1399 2812 1468 2814
rect 1399 2811 1400 2812
rect 1394 2810 1400 2811
rect 1467 2811 1468 2812
rect 1472 2811 1473 2815
rect 1467 2810 1473 2811
rect 1651 2815 1657 2816
rect 1651 2811 1652 2815
rect 1656 2814 1657 2815
rect 1682 2815 1688 2816
rect 1682 2814 1683 2815
rect 1656 2812 1683 2814
rect 1656 2811 1657 2812
rect 1651 2810 1657 2811
rect 1682 2811 1683 2812
rect 1687 2811 1688 2815
rect 1682 2810 1688 2811
rect 1835 2815 1841 2816
rect 1835 2811 1836 2815
rect 1840 2814 1841 2815
rect 1858 2815 1864 2816
rect 1858 2814 1859 2815
rect 1840 2812 1859 2814
rect 1840 2811 1841 2812
rect 1835 2810 1841 2811
rect 1858 2811 1859 2812
rect 1863 2811 1864 2815
rect 1858 2810 1864 2811
rect 478 2792 484 2793
rect 110 2789 116 2790
rect 110 2785 111 2789
rect 115 2785 116 2789
rect 478 2788 479 2792
rect 483 2788 484 2792
rect 478 2787 484 2788
rect 574 2792 580 2793
rect 574 2788 575 2792
rect 579 2788 580 2792
rect 574 2787 580 2788
rect 678 2792 684 2793
rect 678 2788 679 2792
rect 683 2788 684 2792
rect 678 2787 684 2788
rect 798 2792 804 2793
rect 798 2788 799 2792
rect 803 2788 804 2792
rect 798 2787 804 2788
rect 934 2792 940 2793
rect 934 2788 935 2792
rect 939 2788 940 2792
rect 934 2787 940 2788
rect 1078 2792 1084 2793
rect 1078 2788 1079 2792
rect 1083 2788 1084 2792
rect 1078 2787 1084 2788
rect 1238 2792 1244 2793
rect 1238 2788 1239 2792
rect 1243 2788 1244 2792
rect 1238 2787 1244 2788
rect 1414 2792 1420 2793
rect 1414 2788 1415 2792
rect 1419 2788 1420 2792
rect 1414 2787 1420 2788
rect 1598 2792 1604 2793
rect 1598 2788 1599 2792
rect 1603 2788 1604 2792
rect 1598 2787 1604 2788
rect 1782 2792 1788 2793
rect 1782 2788 1783 2792
rect 1787 2788 1788 2792
rect 1782 2787 1788 2788
rect 2006 2789 2012 2790
rect 110 2784 116 2785
rect 2006 2785 2007 2789
rect 2011 2785 2012 2789
rect 2006 2784 2012 2785
rect 2046 2784 2052 2785
rect 3942 2784 3948 2785
rect 546 2783 552 2784
rect 546 2779 547 2783
rect 551 2779 552 2783
rect 546 2778 552 2779
rect 562 2783 568 2784
rect 562 2779 563 2783
rect 567 2782 568 2783
rect 658 2783 664 2784
rect 567 2780 617 2782
rect 567 2779 568 2780
rect 562 2778 568 2779
rect 658 2779 659 2783
rect 663 2782 664 2783
rect 762 2783 768 2784
rect 663 2780 721 2782
rect 663 2779 664 2780
rect 658 2778 664 2779
rect 762 2779 763 2783
rect 767 2782 768 2783
rect 882 2783 888 2784
rect 767 2780 841 2782
rect 767 2779 768 2780
rect 762 2778 768 2779
rect 882 2779 883 2783
rect 887 2782 888 2783
rect 1150 2783 1156 2784
rect 887 2780 977 2782
rect 887 2779 888 2780
rect 882 2778 888 2779
rect 1150 2779 1151 2783
rect 1155 2779 1156 2783
rect 1150 2778 1156 2779
rect 1190 2783 1196 2784
rect 1190 2779 1191 2783
rect 1195 2782 1196 2783
rect 1326 2783 1332 2784
rect 1195 2780 1281 2782
rect 1195 2779 1196 2780
rect 1190 2778 1196 2779
rect 1326 2779 1327 2783
rect 1331 2782 1332 2783
rect 1550 2783 1556 2784
rect 1331 2780 1457 2782
rect 1331 2779 1332 2780
rect 1326 2778 1332 2779
rect 1550 2779 1551 2783
rect 1555 2782 1556 2783
rect 1682 2783 1688 2784
rect 1555 2780 1641 2782
rect 1555 2779 1556 2780
rect 1550 2778 1556 2779
rect 1682 2779 1683 2783
rect 1687 2782 1688 2783
rect 1687 2780 1825 2782
rect 2046 2780 2047 2784
rect 2051 2780 2052 2784
rect 1687 2779 1688 2780
rect 2046 2779 2052 2780
rect 2070 2783 2076 2784
rect 2070 2779 2071 2783
rect 2075 2779 2076 2783
rect 1682 2778 1688 2779
rect 2070 2778 2076 2779
rect 2198 2783 2204 2784
rect 2198 2779 2199 2783
rect 2203 2779 2204 2783
rect 2198 2778 2204 2779
rect 2366 2783 2372 2784
rect 2366 2779 2367 2783
rect 2371 2779 2372 2783
rect 2366 2778 2372 2779
rect 2550 2783 2556 2784
rect 2550 2779 2551 2783
rect 2555 2779 2556 2783
rect 2550 2778 2556 2779
rect 2734 2783 2740 2784
rect 2734 2779 2735 2783
rect 2739 2779 2740 2783
rect 2734 2778 2740 2779
rect 2926 2783 2932 2784
rect 2926 2779 2927 2783
rect 2931 2779 2932 2783
rect 2926 2778 2932 2779
rect 3110 2783 3116 2784
rect 3110 2779 3111 2783
rect 3115 2779 3116 2783
rect 3110 2778 3116 2779
rect 3294 2783 3300 2784
rect 3294 2779 3295 2783
rect 3299 2779 3300 2783
rect 3294 2778 3300 2779
rect 3478 2783 3484 2784
rect 3478 2779 3479 2783
rect 3483 2779 3484 2783
rect 3478 2778 3484 2779
rect 3670 2783 3676 2784
rect 3670 2779 3671 2783
rect 3675 2779 3676 2783
rect 3670 2778 3676 2779
rect 3838 2783 3844 2784
rect 3838 2779 3839 2783
rect 3843 2779 3844 2783
rect 3942 2780 3943 2784
rect 3947 2780 3948 2784
rect 3838 2778 3844 2779
rect 3906 2779 3912 2780
rect 3942 2779 3948 2780
rect 2658 2775 2664 2776
rect 478 2773 484 2774
rect 110 2772 116 2773
rect 110 2768 111 2772
rect 115 2768 116 2772
rect 478 2769 479 2773
rect 483 2769 484 2773
rect 478 2768 484 2769
rect 574 2773 580 2774
rect 574 2769 575 2773
rect 579 2769 580 2773
rect 574 2768 580 2769
rect 678 2773 684 2774
rect 678 2769 679 2773
rect 683 2769 684 2773
rect 678 2768 684 2769
rect 798 2773 804 2774
rect 798 2769 799 2773
rect 803 2769 804 2773
rect 798 2768 804 2769
rect 934 2773 940 2774
rect 934 2769 935 2773
rect 939 2769 940 2773
rect 934 2768 940 2769
rect 1078 2773 1084 2774
rect 1078 2769 1079 2773
rect 1083 2769 1084 2773
rect 1078 2768 1084 2769
rect 1238 2773 1244 2774
rect 1238 2769 1239 2773
rect 1243 2769 1244 2773
rect 1238 2768 1244 2769
rect 1414 2773 1420 2774
rect 1414 2769 1415 2773
rect 1419 2769 1420 2773
rect 1414 2768 1420 2769
rect 1598 2773 1604 2774
rect 1598 2769 1599 2773
rect 1603 2769 1604 2773
rect 1598 2768 1604 2769
rect 1782 2773 1788 2774
rect 1782 2769 1783 2773
rect 1787 2769 1788 2773
rect 1782 2768 1788 2769
rect 2006 2772 2012 2773
rect 2006 2768 2007 2772
rect 2011 2768 2012 2772
rect 2146 2771 2152 2772
rect 110 2767 116 2768
rect 2006 2767 2012 2768
rect 2046 2767 2052 2768
rect 2046 2763 2047 2767
rect 2051 2763 2052 2767
rect 2146 2767 2147 2771
rect 2151 2767 2152 2771
rect 2146 2766 2152 2767
rect 2274 2771 2280 2772
rect 2274 2767 2275 2771
rect 2279 2767 2280 2771
rect 2274 2766 2280 2767
rect 2442 2771 2448 2772
rect 2442 2767 2443 2771
rect 2447 2767 2448 2771
rect 2442 2766 2448 2767
rect 2626 2771 2632 2772
rect 2626 2767 2627 2771
rect 2631 2767 2632 2771
rect 2658 2771 2659 2775
rect 2663 2774 2664 2775
rect 3438 2775 3444 2776
rect 2663 2772 2777 2774
rect 2663 2771 2664 2772
rect 2658 2770 2664 2771
rect 3002 2771 3008 2772
rect 2626 2766 2632 2767
rect 3002 2767 3003 2771
rect 3007 2767 3008 2771
rect 3002 2766 3008 2767
rect 3186 2771 3192 2772
rect 3186 2767 3187 2771
rect 3191 2767 3192 2771
rect 3186 2766 3192 2767
rect 3370 2771 3376 2772
rect 3370 2767 3371 2771
rect 3375 2767 3376 2771
rect 3438 2771 3439 2775
rect 3443 2774 3444 2775
rect 3906 2775 3907 2779
rect 3911 2775 3912 2779
rect 3906 2774 3912 2775
rect 3443 2772 3521 2774
rect 3908 2772 3917 2774
rect 3443 2771 3444 2772
rect 3438 2770 3444 2771
rect 3746 2771 3752 2772
rect 3370 2766 3376 2767
rect 3746 2767 3747 2771
rect 3751 2767 3752 2771
rect 3746 2766 3752 2767
rect 3942 2767 3948 2768
rect 2046 2762 2052 2763
rect 2070 2764 2076 2765
rect 2070 2760 2071 2764
rect 2075 2760 2076 2764
rect 2070 2759 2076 2760
rect 2198 2764 2204 2765
rect 2198 2760 2199 2764
rect 2203 2760 2204 2764
rect 2198 2759 2204 2760
rect 2366 2764 2372 2765
rect 2366 2760 2367 2764
rect 2371 2760 2372 2764
rect 2366 2759 2372 2760
rect 2550 2764 2556 2765
rect 2550 2760 2551 2764
rect 2555 2760 2556 2764
rect 2550 2759 2556 2760
rect 2734 2764 2740 2765
rect 2734 2760 2735 2764
rect 2739 2760 2740 2764
rect 2734 2759 2740 2760
rect 2926 2764 2932 2765
rect 2926 2760 2927 2764
rect 2931 2760 2932 2764
rect 2926 2759 2932 2760
rect 3110 2764 3116 2765
rect 3110 2760 3111 2764
rect 3115 2760 3116 2764
rect 3110 2759 3116 2760
rect 3294 2764 3300 2765
rect 3294 2760 3295 2764
rect 3299 2760 3300 2764
rect 3294 2759 3300 2760
rect 3478 2764 3484 2765
rect 3478 2760 3479 2764
rect 3483 2760 3484 2764
rect 3478 2759 3484 2760
rect 3670 2764 3676 2765
rect 3670 2760 3671 2764
rect 3675 2760 3676 2764
rect 3670 2759 3676 2760
rect 3838 2764 3844 2765
rect 3838 2760 3839 2764
rect 3843 2760 3844 2764
rect 3942 2763 3943 2767
rect 3947 2763 3948 2767
rect 3942 2762 3948 2763
rect 3838 2759 3844 2760
rect 2718 2751 2724 2752
rect 2718 2750 2719 2751
rect 2140 2748 2719 2750
rect 2123 2743 2129 2744
rect 2123 2739 2124 2743
rect 2128 2742 2129 2743
rect 2140 2742 2142 2748
rect 2718 2747 2719 2748
rect 2723 2747 2724 2751
rect 2718 2746 2724 2747
rect 2128 2740 2142 2742
rect 2146 2743 2152 2744
rect 2128 2739 2129 2740
rect 2123 2738 2129 2739
rect 2146 2739 2147 2743
rect 2151 2742 2152 2743
rect 2251 2743 2257 2744
rect 2251 2742 2252 2743
rect 2151 2740 2252 2742
rect 2151 2739 2152 2740
rect 2146 2738 2152 2739
rect 2251 2739 2252 2740
rect 2256 2739 2257 2743
rect 2251 2738 2257 2739
rect 2274 2743 2280 2744
rect 2274 2739 2275 2743
rect 2279 2742 2280 2743
rect 2419 2743 2425 2744
rect 2419 2742 2420 2743
rect 2279 2740 2420 2742
rect 2279 2739 2280 2740
rect 2274 2738 2280 2739
rect 2419 2739 2420 2740
rect 2424 2739 2425 2743
rect 2419 2738 2425 2739
rect 2442 2743 2448 2744
rect 2442 2739 2443 2743
rect 2447 2742 2448 2743
rect 2603 2743 2609 2744
rect 2603 2742 2604 2743
rect 2447 2740 2604 2742
rect 2447 2739 2448 2740
rect 2442 2738 2448 2739
rect 2603 2739 2604 2740
rect 2608 2739 2609 2743
rect 2603 2738 2609 2739
rect 2626 2743 2632 2744
rect 2626 2739 2627 2743
rect 2631 2742 2632 2743
rect 2787 2743 2793 2744
rect 2787 2742 2788 2743
rect 2631 2740 2788 2742
rect 2631 2739 2632 2740
rect 2626 2738 2632 2739
rect 2787 2739 2788 2740
rect 2792 2739 2793 2743
rect 3002 2743 3008 2744
rect 2787 2738 2793 2739
rect 2979 2739 2985 2740
rect 2979 2735 2980 2739
rect 2984 2738 2985 2739
rect 3002 2739 3003 2743
rect 3007 2742 3008 2743
rect 3163 2743 3169 2744
rect 3163 2742 3164 2743
rect 3007 2740 3164 2742
rect 3007 2739 3008 2740
rect 3002 2738 3008 2739
rect 3163 2739 3164 2740
rect 3168 2739 3169 2743
rect 3163 2738 3169 2739
rect 3186 2743 3192 2744
rect 3186 2739 3187 2743
rect 3191 2742 3192 2743
rect 3347 2743 3353 2744
rect 3347 2742 3348 2743
rect 3191 2740 3348 2742
rect 3191 2739 3192 2740
rect 3186 2738 3192 2739
rect 3347 2739 3348 2740
rect 3352 2739 3353 2743
rect 3347 2738 3353 2739
rect 3370 2743 3376 2744
rect 3370 2739 3371 2743
rect 3375 2742 3376 2743
rect 3531 2743 3537 2744
rect 3531 2742 3532 2743
rect 3375 2740 3532 2742
rect 3375 2739 3376 2740
rect 3370 2738 3376 2739
rect 3531 2739 3532 2740
rect 3536 2739 3537 2743
rect 3531 2738 3537 2739
rect 3723 2743 3729 2744
rect 3723 2739 3724 2743
rect 3728 2742 3729 2743
rect 3874 2743 3880 2744
rect 3874 2742 3875 2743
rect 3728 2740 3875 2742
rect 3728 2739 3729 2740
rect 3723 2738 3729 2739
rect 3874 2739 3875 2740
rect 3879 2739 3880 2743
rect 3874 2738 3880 2739
rect 3891 2739 3897 2740
rect 2984 2736 2998 2738
rect 2984 2735 2985 2736
rect 2979 2734 2985 2735
rect 2996 2734 2998 2736
rect 3378 2735 3384 2736
rect 3378 2734 3379 2735
rect 2996 2732 3379 2734
rect 2658 2731 2664 2732
rect 2658 2730 2659 2731
rect 2124 2728 2659 2730
rect 2124 2726 2126 2728
rect 2658 2727 2659 2728
rect 2663 2727 2664 2731
rect 3378 2731 3379 2732
rect 3383 2731 3384 2735
rect 3891 2735 3892 2739
rect 3896 2738 3897 2739
rect 3906 2739 3912 2740
rect 3906 2738 3907 2739
rect 3896 2736 3907 2738
rect 3896 2735 3897 2736
rect 3891 2734 3897 2735
rect 3906 2735 3907 2736
rect 3911 2735 3912 2739
rect 3906 2734 3912 2735
rect 3378 2730 3384 2731
rect 2658 2726 2664 2727
rect 2123 2725 2129 2726
rect 2123 2721 2124 2725
rect 2128 2721 2129 2725
rect 2123 2720 2129 2721
rect 2146 2723 2152 2724
rect 2146 2719 2147 2723
rect 2151 2722 2152 2723
rect 2243 2723 2249 2724
rect 2243 2722 2244 2723
rect 2151 2720 2244 2722
rect 2151 2719 2152 2720
rect 2146 2718 2152 2719
rect 2243 2719 2244 2720
rect 2248 2719 2249 2723
rect 2243 2718 2249 2719
rect 2266 2723 2272 2724
rect 2266 2719 2267 2723
rect 2271 2722 2272 2723
rect 2371 2723 2377 2724
rect 2371 2722 2372 2723
rect 2271 2720 2372 2722
rect 2271 2719 2272 2720
rect 2266 2718 2272 2719
rect 2371 2719 2372 2720
rect 2376 2719 2377 2723
rect 2371 2718 2377 2719
rect 2394 2723 2400 2724
rect 2394 2719 2395 2723
rect 2399 2722 2400 2723
rect 2499 2723 2505 2724
rect 2499 2722 2500 2723
rect 2399 2720 2500 2722
rect 2399 2719 2400 2720
rect 2394 2718 2400 2719
rect 2499 2719 2500 2720
rect 2504 2719 2505 2723
rect 2499 2718 2505 2719
rect 2522 2723 2528 2724
rect 2522 2719 2523 2723
rect 2527 2722 2528 2723
rect 2635 2723 2641 2724
rect 2635 2722 2636 2723
rect 2527 2720 2636 2722
rect 2527 2719 2528 2720
rect 2522 2718 2528 2719
rect 2635 2719 2636 2720
rect 2640 2719 2641 2723
rect 2635 2718 2641 2719
rect 2779 2723 2788 2724
rect 2779 2719 2780 2723
rect 2787 2719 2788 2723
rect 2779 2718 2788 2719
rect 2802 2723 2808 2724
rect 2802 2719 2803 2723
rect 2807 2722 2808 2723
rect 2939 2723 2945 2724
rect 2939 2722 2940 2723
rect 2807 2720 2940 2722
rect 2807 2719 2808 2720
rect 2802 2718 2808 2719
rect 2939 2719 2940 2720
rect 2944 2719 2945 2723
rect 2939 2718 2945 2719
rect 2962 2723 2968 2724
rect 2962 2719 2963 2723
rect 2967 2722 2968 2723
rect 3115 2723 3121 2724
rect 3115 2722 3116 2723
rect 2967 2720 3116 2722
rect 2967 2719 2968 2720
rect 2962 2718 2968 2719
rect 3115 2719 3116 2720
rect 3120 2719 3121 2723
rect 3115 2718 3121 2719
rect 3138 2723 3144 2724
rect 3138 2719 3139 2723
rect 3143 2722 3144 2723
rect 3307 2723 3313 2724
rect 3307 2722 3308 2723
rect 3143 2720 3308 2722
rect 3143 2719 3144 2720
rect 3138 2718 3144 2719
rect 3307 2719 3308 2720
rect 3312 2719 3313 2723
rect 3307 2718 3313 2719
rect 3330 2723 3336 2724
rect 3330 2719 3331 2723
rect 3335 2722 3336 2723
rect 3507 2723 3513 2724
rect 3507 2722 3508 2723
rect 3335 2720 3508 2722
rect 3335 2719 3336 2720
rect 3330 2718 3336 2719
rect 3507 2719 3508 2720
rect 3512 2719 3513 2723
rect 3507 2718 3513 2719
rect 3707 2723 3713 2724
rect 3707 2719 3708 2723
rect 3712 2722 3713 2723
rect 3746 2723 3752 2724
rect 3746 2722 3747 2723
rect 3712 2720 3747 2722
rect 3712 2719 3713 2720
rect 3707 2718 3713 2719
rect 3746 2719 3747 2720
rect 3751 2719 3752 2723
rect 3746 2718 3752 2719
rect 3791 2723 3797 2724
rect 3791 2719 3792 2723
rect 3796 2722 3797 2723
rect 3891 2723 3897 2724
rect 3891 2722 3892 2723
rect 3796 2720 3892 2722
rect 3796 2719 3797 2720
rect 3791 2718 3797 2719
rect 3891 2719 3892 2720
rect 3896 2719 3897 2723
rect 3891 2718 3897 2719
rect 110 2716 116 2717
rect 2006 2716 2012 2717
rect 110 2712 111 2716
rect 115 2712 116 2716
rect 110 2711 116 2712
rect 510 2715 516 2716
rect 510 2711 511 2715
rect 515 2711 516 2715
rect 510 2710 516 2711
rect 622 2715 628 2716
rect 622 2711 623 2715
rect 627 2711 628 2715
rect 622 2710 628 2711
rect 742 2715 748 2716
rect 742 2711 743 2715
rect 747 2711 748 2715
rect 742 2710 748 2711
rect 878 2715 884 2716
rect 878 2711 879 2715
rect 883 2711 884 2715
rect 878 2710 884 2711
rect 1014 2715 1020 2716
rect 1014 2711 1015 2715
rect 1019 2711 1020 2715
rect 1014 2710 1020 2711
rect 1158 2715 1164 2716
rect 1158 2711 1159 2715
rect 1163 2711 1164 2715
rect 1158 2710 1164 2711
rect 1310 2715 1316 2716
rect 1310 2711 1311 2715
rect 1315 2711 1316 2715
rect 1310 2710 1316 2711
rect 1462 2715 1468 2716
rect 1462 2711 1463 2715
rect 1467 2711 1468 2715
rect 1462 2710 1468 2711
rect 1622 2715 1628 2716
rect 1622 2711 1623 2715
rect 1627 2711 1628 2715
rect 1622 2710 1628 2711
rect 1782 2715 1788 2716
rect 1782 2711 1783 2715
rect 1787 2711 1788 2715
rect 2006 2712 2007 2716
rect 2011 2712 2012 2716
rect 2006 2711 2012 2712
rect 1782 2710 1788 2711
rect 998 2707 1004 2708
rect 586 2703 592 2704
rect 110 2699 116 2700
rect 110 2695 111 2699
rect 115 2695 116 2699
rect 586 2699 587 2703
rect 591 2699 592 2703
rect 586 2698 592 2699
rect 698 2703 704 2704
rect 698 2699 699 2703
rect 703 2699 704 2703
rect 698 2698 704 2699
rect 818 2703 824 2704
rect 818 2699 819 2703
rect 823 2699 824 2703
rect 818 2698 824 2699
rect 954 2703 960 2704
rect 954 2699 955 2703
rect 959 2699 960 2703
rect 998 2703 999 2707
rect 1003 2706 1004 2707
rect 1858 2707 1864 2708
rect 1003 2704 1057 2706
rect 1003 2703 1004 2704
rect 998 2702 1004 2703
rect 1234 2703 1240 2704
rect 954 2698 960 2699
rect 1234 2699 1235 2703
rect 1239 2699 1240 2703
rect 1234 2698 1240 2699
rect 1386 2703 1392 2704
rect 1386 2699 1387 2703
rect 1391 2699 1392 2703
rect 1386 2698 1392 2699
rect 1538 2703 1544 2704
rect 1538 2699 1539 2703
rect 1543 2699 1544 2703
rect 1538 2698 1544 2699
rect 1698 2703 1704 2704
rect 1698 2699 1699 2703
rect 1703 2699 1704 2703
rect 1858 2703 1859 2707
rect 1863 2703 1864 2707
rect 1858 2702 1864 2703
rect 2070 2700 2076 2701
rect 1698 2698 1704 2699
rect 2006 2699 2012 2700
rect 110 2694 116 2695
rect 510 2696 516 2697
rect 510 2692 511 2696
rect 515 2692 516 2696
rect 510 2691 516 2692
rect 622 2696 628 2697
rect 622 2692 623 2696
rect 627 2692 628 2696
rect 622 2691 628 2692
rect 742 2696 748 2697
rect 742 2692 743 2696
rect 747 2692 748 2696
rect 742 2691 748 2692
rect 878 2696 884 2697
rect 878 2692 879 2696
rect 883 2692 884 2696
rect 878 2691 884 2692
rect 1014 2696 1020 2697
rect 1014 2692 1015 2696
rect 1019 2692 1020 2696
rect 1014 2691 1020 2692
rect 1158 2696 1164 2697
rect 1158 2692 1159 2696
rect 1163 2692 1164 2696
rect 1158 2691 1164 2692
rect 1310 2696 1316 2697
rect 1310 2692 1311 2696
rect 1315 2692 1316 2696
rect 1310 2691 1316 2692
rect 1462 2696 1468 2697
rect 1462 2692 1463 2696
rect 1467 2692 1468 2696
rect 1462 2691 1468 2692
rect 1622 2696 1628 2697
rect 1622 2692 1623 2696
rect 1627 2692 1628 2696
rect 1622 2691 1628 2692
rect 1782 2696 1788 2697
rect 1782 2692 1783 2696
rect 1787 2692 1788 2696
rect 2006 2695 2007 2699
rect 2011 2695 2012 2699
rect 2006 2694 2012 2695
rect 2046 2697 2052 2698
rect 2046 2693 2047 2697
rect 2051 2693 2052 2697
rect 2070 2696 2071 2700
rect 2075 2696 2076 2700
rect 2070 2695 2076 2696
rect 2190 2700 2196 2701
rect 2190 2696 2191 2700
rect 2195 2696 2196 2700
rect 2190 2695 2196 2696
rect 2318 2700 2324 2701
rect 2318 2696 2319 2700
rect 2323 2696 2324 2700
rect 2318 2695 2324 2696
rect 2446 2700 2452 2701
rect 2446 2696 2447 2700
rect 2451 2696 2452 2700
rect 2446 2695 2452 2696
rect 2582 2700 2588 2701
rect 2582 2696 2583 2700
rect 2587 2696 2588 2700
rect 2582 2695 2588 2696
rect 2726 2700 2732 2701
rect 2726 2696 2727 2700
rect 2731 2696 2732 2700
rect 2726 2695 2732 2696
rect 2886 2700 2892 2701
rect 2886 2696 2887 2700
rect 2891 2696 2892 2700
rect 2886 2695 2892 2696
rect 3062 2700 3068 2701
rect 3062 2696 3063 2700
rect 3067 2696 3068 2700
rect 3062 2695 3068 2696
rect 3254 2700 3260 2701
rect 3254 2696 3255 2700
rect 3259 2696 3260 2700
rect 3254 2695 3260 2696
rect 3454 2700 3460 2701
rect 3454 2696 3455 2700
rect 3459 2696 3460 2700
rect 3454 2695 3460 2696
rect 3654 2700 3660 2701
rect 3654 2696 3655 2700
rect 3659 2696 3660 2700
rect 3654 2695 3660 2696
rect 3838 2700 3844 2701
rect 3838 2696 3839 2700
rect 3843 2696 3844 2700
rect 3838 2695 3844 2696
rect 3942 2697 3948 2698
rect 2046 2692 2052 2693
rect 3942 2693 3943 2697
rect 3947 2693 3948 2697
rect 3942 2692 3948 2693
rect 1782 2691 1788 2692
rect 2146 2691 2152 2692
rect 2146 2687 2147 2691
rect 2151 2687 2152 2691
rect 2146 2686 2152 2687
rect 2266 2691 2272 2692
rect 2266 2687 2267 2691
rect 2271 2687 2272 2691
rect 2266 2686 2272 2687
rect 2394 2691 2400 2692
rect 2394 2687 2395 2691
rect 2399 2687 2400 2691
rect 2394 2686 2400 2687
rect 2522 2691 2528 2692
rect 2522 2687 2523 2691
rect 2527 2687 2528 2691
rect 2522 2686 2528 2687
rect 2538 2691 2544 2692
rect 2538 2687 2539 2691
rect 2543 2690 2544 2691
rect 2802 2691 2808 2692
rect 2543 2688 2625 2690
rect 2543 2687 2544 2688
rect 2538 2686 2544 2687
rect 2802 2687 2803 2691
rect 2807 2687 2808 2691
rect 2802 2686 2808 2687
rect 2962 2691 2968 2692
rect 2962 2687 2963 2691
rect 2967 2687 2968 2691
rect 2962 2686 2968 2687
rect 3138 2691 3144 2692
rect 3138 2687 3139 2691
rect 3143 2687 3144 2691
rect 3138 2686 3144 2687
rect 3330 2691 3336 2692
rect 3330 2687 3331 2691
rect 3335 2687 3336 2691
rect 3330 2686 3336 2687
rect 3378 2691 3384 2692
rect 3378 2687 3379 2691
rect 3383 2690 3384 2691
rect 3791 2691 3797 2692
rect 3791 2690 3792 2691
rect 3383 2688 3497 2690
rect 3733 2688 3792 2690
rect 3383 2687 3384 2688
rect 3378 2686 3384 2687
rect 3791 2687 3792 2688
rect 3796 2687 3797 2691
rect 3791 2686 3797 2687
rect 3906 2691 3912 2692
rect 3906 2687 3907 2691
rect 3911 2687 3912 2691
rect 3906 2686 3912 2687
rect 2070 2681 2076 2682
rect 2046 2680 2052 2681
rect 2046 2676 2047 2680
rect 2051 2676 2052 2680
rect 2070 2677 2071 2681
rect 2075 2677 2076 2681
rect 2070 2676 2076 2677
rect 2190 2681 2196 2682
rect 2190 2677 2191 2681
rect 2195 2677 2196 2681
rect 2190 2676 2196 2677
rect 2318 2681 2324 2682
rect 2318 2677 2319 2681
rect 2323 2677 2324 2681
rect 2318 2676 2324 2677
rect 2446 2681 2452 2682
rect 2446 2677 2447 2681
rect 2451 2677 2452 2681
rect 2446 2676 2452 2677
rect 2582 2681 2588 2682
rect 2582 2677 2583 2681
rect 2587 2677 2588 2681
rect 2582 2676 2588 2677
rect 2726 2681 2732 2682
rect 2726 2677 2727 2681
rect 2731 2677 2732 2681
rect 2726 2676 2732 2677
rect 2886 2681 2892 2682
rect 2886 2677 2887 2681
rect 2891 2677 2892 2681
rect 2886 2676 2892 2677
rect 3062 2681 3068 2682
rect 3062 2677 3063 2681
rect 3067 2677 3068 2681
rect 3062 2676 3068 2677
rect 3254 2681 3260 2682
rect 3254 2677 3255 2681
rect 3259 2677 3260 2681
rect 3254 2676 3260 2677
rect 3454 2681 3460 2682
rect 3454 2677 3455 2681
rect 3459 2677 3460 2681
rect 3454 2676 3460 2677
rect 3654 2681 3660 2682
rect 3654 2677 3655 2681
rect 3659 2677 3660 2681
rect 3654 2676 3660 2677
rect 3838 2681 3844 2682
rect 3838 2677 3839 2681
rect 3843 2677 3844 2681
rect 3838 2676 3844 2677
rect 3942 2680 3948 2681
rect 3942 2676 3943 2680
rect 3947 2676 3948 2680
rect 586 2675 592 2676
rect 563 2671 569 2672
rect 563 2667 564 2671
rect 568 2670 569 2671
rect 586 2671 587 2675
rect 591 2674 592 2675
rect 675 2675 681 2676
rect 675 2674 676 2675
rect 591 2672 676 2674
rect 591 2671 592 2672
rect 586 2670 592 2671
rect 675 2671 676 2672
rect 680 2671 681 2675
rect 675 2670 681 2671
rect 698 2675 704 2676
rect 698 2671 699 2675
rect 703 2674 704 2675
rect 795 2675 801 2676
rect 795 2674 796 2675
rect 703 2672 796 2674
rect 703 2671 704 2672
rect 698 2670 704 2671
rect 795 2671 796 2672
rect 800 2671 801 2675
rect 795 2670 801 2671
rect 818 2675 824 2676
rect 818 2671 819 2675
rect 823 2674 824 2675
rect 931 2675 937 2676
rect 931 2674 932 2675
rect 823 2672 932 2674
rect 823 2671 824 2672
rect 818 2670 824 2671
rect 931 2671 932 2672
rect 936 2671 937 2675
rect 931 2670 937 2671
rect 954 2675 960 2676
rect 954 2671 955 2675
rect 959 2674 960 2675
rect 1067 2675 1073 2676
rect 1067 2674 1068 2675
rect 959 2672 1068 2674
rect 959 2671 960 2672
rect 954 2670 960 2671
rect 1067 2671 1068 2672
rect 1072 2671 1073 2675
rect 1067 2670 1073 2671
rect 1150 2675 1156 2676
rect 1150 2671 1151 2675
rect 1155 2674 1156 2675
rect 1211 2675 1217 2676
rect 1211 2674 1212 2675
rect 1155 2672 1212 2674
rect 1155 2671 1156 2672
rect 1150 2670 1156 2671
rect 1211 2671 1212 2672
rect 1216 2671 1217 2675
rect 1211 2670 1217 2671
rect 1234 2675 1240 2676
rect 1234 2671 1235 2675
rect 1239 2674 1240 2675
rect 1363 2675 1369 2676
rect 1363 2674 1364 2675
rect 1239 2672 1364 2674
rect 1239 2671 1240 2672
rect 1234 2670 1240 2671
rect 1363 2671 1364 2672
rect 1368 2671 1369 2675
rect 1538 2675 1544 2676
rect 1363 2670 1369 2671
rect 1506 2671 1512 2672
rect 568 2668 582 2670
rect 568 2667 569 2668
rect 563 2666 569 2667
rect 580 2666 582 2668
rect 858 2667 864 2668
rect 858 2666 859 2667
rect 580 2664 859 2666
rect 858 2663 859 2664
rect 863 2663 864 2667
rect 1506 2667 1507 2671
rect 1511 2670 1512 2671
rect 1515 2671 1521 2672
rect 1515 2670 1516 2671
rect 1511 2668 1516 2670
rect 1511 2667 1512 2668
rect 1506 2666 1512 2667
rect 1515 2667 1516 2668
rect 1520 2667 1521 2671
rect 1538 2671 1539 2675
rect 1543 2674 1544 2675
rect 1675 2675 1681 2676
rect 1675 2674 1676 2675
rect 1543 2672 1676 2674
rect 1543 2671 1544 2672
rect 1538 2670 1544 2671
rect 1675 2671 1676 2672
rect 1680 2671 1681 2675
rect 1675 2670 1681 2671
rect 1698 2675 1704 2676
rect 1698 2671 1699 2675
rect 1703 2674 1704 2675
rect 1835 2675 1841 2676
rect 2046 2675 2052 2676
rect 3942 2675 3948 2676
rect 1835 2674 1836 2675
rect 1703 2672 1836 2674
rect 1703 2671 1704 2672
rect 1698 2670 1704 2671
rect 1835 2671 1836 2672
rect 1840 2671 1841 2675
rect 1835 2670 1841 2671
rect 1515 2666 1521 2667
rect 858 2662 864 2663
rect 442 2655 448 2656
rect 419 2653 425 2654
rect 419 2649 420 2653
rect 424 2649 425 2653
rect 442 2651 443 2655
rect 447 2654 448 2655
rect 539 2655 545 2656
rect 539 2654 540 2655
rect 447 2652 540 2654
rect 447 2651 448 2652
rect 442 2650 448 2651
rect 539 2651 540 2652
rect 544 2651 545 2655
rect 539 2650 545 2651
rect 562 2655 568 2656
rect 562 2651 563 2655
rect 567 2654 568 2655
rect 667 2655 673 2656
rect 667 2654 668 2655
rect 567 2652 668 2654
rect 567 2651 568 2652
rect 562 2650 568 2651
rect 667 2651 668 2652
rect 672 2651 673 2655
rect 667 2650 673 2651
rect 690 2655 696 2656
rect 690 2651 691 2655
rect 695 2654 696 2655
rect 803 2655 809 2656
rect 803 2654 804 2655
rect 695 2652 804 2654
rect 695 2651 696 2652
rect 690 2650 696 2651
rect 803 2651 804 2652
rect 808 2651 809 2655
rect 803 2650 809 2651
rect 826 2655 832 2656
rect 826 2651 827 2655
rect 831 2654 832 2655
rect 947 2655 953 2656
rect 947 2654 948 2655
rect 831 2652 948 2654
rect 831 2651 832 2652
rect 826 2650 832 2651
rect 947 2651 948 2652
rect 952 2651 953 2655
rect 947 2650 953 2651
rect 1083 2655 1089 2656
rect 1083 2651 1084 2655
rect 1088 2654 1089 2655
rect 1119 2655 1125 2656
rect 1119 2654 1120 2655
rect 1088 2652 1120 2654
rect 1088 2651 1089 2652
rect 1083 2650 1089 2651
rect 1119 2651 1120 2652
rect 1124 2651 1125 2655
rect 1119 2650 1125 2651
rect 1219 2655 1225 2656
rect 1219 2651 1220 2655
rect 1224 2654 1225 2655
rect 1250 2655 1256 2656
rect 1250 2654 1251 2655
rect 1224 2652 1251 2654
rect 1224 2651 1225 2652
rect 1219 2650 1225 2651
rect 1250 2651 1251 2652
rect 1255 2651 1256 2655
rect 1250 2650 1256 2651
rect 1355 2655 1361 2656
rect 1355 2651 1356 2655
rect 1360 2654 1361 2655
rect 1386 2655 1392 2656
rect 1386 2654 1387 2655
rect 1360 2652 1387 2654
rect 1360 2651 1361 2652
rect 1355 2650 1361 2651
rect 1386 2651 1387 2652
rect 1391 2651 1392 2655
rect 1386 2650 1392 2651
rect 1483 2655 1489 2656
rect 1483 2651 1484 2655
rect 1488 2654 1489 2655
rect 1514 2655 1520 2656
rect 1514 2654 1515 2655
rect 1488 2652 1515 2654
rect 1488 2651 1489 2652
rect 1483 2650 1489 2651
rect 1514 2651 1515 2652
rect 1519 2651 1520 2655
rect 1514 2650 1520 2651
rect 1619 2655 1625 2656
rect 1619 2651 1620 2655
rect 1624 2654 1625 2655
rect 1650 2655 1656 2656
rect 1650 2654 1651 2655
rect 1624 2652 1651 2654
rect 1624 2651 1625 2652
rect 1619 2650 1625 2651
rect 1650 2651 1651 2652
rect 1655 2651 1656 2655
rect 1650 2650 1656 2651
rect 1755 2655 1761 2656
rect 1755 2651 1756 2655
rect 1760 2654 1761 2655
rect 1802 2655 1808 2656
rect 1802 2654 1803 2655
rect 1760 2652 1803 2654
rect 1760 2651 1761 2652
rect 1755 2650 1761 2651
rect 1802 2651 1803 2652
rect 1807 2651 1808 2655
rect 1802 2650 1808 2651
rect 419 2648 425 2649
rect 420 2646 422 2648
rect 738 2647 744 2648
rect 738 2646 739 2647
rect 420 2644 739 2646
rect 738 2643 739 2644
rect 743 2643 744 2647
rect 738 2642 744 2643
rect 366 2632 372 2633
rect 110 2629 116 2630
rect 110 2625 111 2629
rect 115 2625 116 2629
rect 366 2628 367 2632
rect 371 2628 372 2632
rect 366 2627 372 2628
rect 486 2632 492 2633
rect 486 2628 487 2632
rect 491 2628 492 2632
rect 486 2627 492 2628
rect 614 2632 620 2633
rect 614 2628 615 2632
rect 619 2628 620 2632
rect 614 2627 620 2628
rect 750 2632 756 2633
rect 750 2628 751 2632
rect 755 2628 756 2632
rect 750 2627 756 2628
rect 894 2632 900 2633
rect 894 2628 895 2632
rect 899 2628 900 2632
rect 894 2627 900 2628
rect 1030 2632 1036 2633
rect 1030 2628 1031 2632
rect 1035 2628 1036 2632
rect 1030 2627 1036 2628
rect 1166 2632 1172 2633
rect 1166 2628 1167 2632
rect 1171 2628 1172 2632
rect 1166 2627 1172 2628
rect 1302 2632 1308 2633
rect 1302 2628 1303 2632
rect 1307 2628 1308 2632
rect 1302 2627 1308 2628
rect 1430 2632 1436 2633
rect 1430 2628 1431 2632
rect 1435 2628 1436 2632
rect 1430 2627 1436 2628
rect 1566 2632 1572 2633
rect 1566 2628 1567 2632
rect 1571 2628 1572 2632
rect 1566 2627 1572 2628
rect 1702 2632 1708 2633
rect 1702 2628 1703 2632
rect 1707 2628 1708 2632
rect 1702 2627 1708 2628
rect 2006 2629 2012 2630
rect 110 2624 116 2625
rect 2006 2625 2007 2629
rect 2011 2625 2012 2629
rect 2006 2624 2012 2625
rect 442 2623 448 2624
rect 442 2619 443 2623
rect 447 2619 448 2623
rect 442 2618 448 2619
rect 562 2623 568 2624
rect 562 2619 563 2623
rect 567 2619 568 2623
rect 562 2618 568 2619
rect 690 2623 696 2624
rect 690 2619 691 2623
rect 695 2619 696 2623
rect 690 2618 696 2619
rect 826 2623 832 2624
rect 826 2619 827 2623
rect 831 2619 832 2623
rect 826 2618 832 2619
rect 858 2623 864 2624
rect 858 2619 859 2623
rect 863 2622 864 2623
rect 978 2623 984 2624
rect 863 2620 937 2622
rect 863 2619 864 2620
rect 858 2618 864 2619
rect 978 2619 979 2623
rect 983 2622 984 2623
rect 1119 2623 1125 2624
rect 983 2620 1073 2622
rect 983 2619 984 2620
rect 978 2618 984 2619
rect 1119 2619 1120 2623
rect 1124 2622 1125 2623
rect 1250 2623 1256 2624
rect 1124 2620 1209 2622
rect 1124 2619 1125 2620
rect 1119 2618 1125 2619
rect 1250 2619 1251 2623
rect 1255 2622 1256 2623
rect 1506 2623 1512 2624
rect 1255 2620 1345 2622
rect 1255 2619 1256 2620
rect 1250 2618 1256 2619
rect 1506 2619 1507 2623
rect 1511 2619 1512 2623
rect 1506 2618 1512 2619
rect 1514 2623 1520 2624
rect 1514 2619 1515 2623
rect 1519 2622 1520 2623
rect 1650 2623 1656 2624
rect 1519 2620 1609 2622
rect 1519 2619 1520 2620
rect 1514 2618 1520 2619
rect 1650 2619 1651 2623
rect 1655 2622 1656 2623
rect 1655 2620 1745 2622
rect 2046 2620 2052 2621
rect 3942 2620 3948 2621
rect 1655 2619 1656 2620
rect 1650 2618 1656 2619
rect 2046 2616 2047 2620
rect 2051 2616 2052 2620
rect 2046 2615 2052 2616
rect 2230 2619 2236 2620
rect 2230 2615 2231 2619
rect 2235 2615 2236 2619
rect 2230 2614 2236 2615
rect 2334 2619 2340 2620
rect 2334 2615 2335 2619
rect 2339 2615 2340 2619
rect 2334 2614 2340 2615
rect 2446 2619 2452 2620
rect 2446 2615 2447 2619
rect 2451 2615 2452 2619
rect 2446 2614 2452 2615
rect 2558 2619 2564 2620
rect 2558 2615 2559 2619
rect 2563 2615 2564 2619
rect 2558 2614 2564 2615
rect 2670 2619 2676 2620
rect 2670 2615 2671 2619
rect 2675 2615 2676 2619
rect 2670 2614 2676 2615
rect 2790 2619 2796 2620
rect 2790 2615 2791 2619
rect 2795 2615 2796 2619
rect 2790 2614 2796 2615
rect 2910 2619 2916 2620
rect 2910 2615 2911 2619
rect 2915 2615 2916 2619
rect 2910 2614 2916 2615
rect 3030 2619 3036 2620
rect 3030 2615 3031 2619
rect 3035 2615 3036 2619
rect 3030 2614 3036 2615
rect 3150 2619 3156 2620
rect 3150 2615 3151 2619
rect 3155 2615 3156 2619
rect 3942 2616 3943 2620
rect 3947 2616 3948 2620
rect 3942 2615 3948 2616
rect 3150 2614 3156 2615
rect 366 2613 372 2614
rect 110 2612 116 2613
rect 110 2608 111 2612
rect 115 2608 116 2612
rect 366 2609 367 2613
rect 371 2609 372 2613
rect 366 2608 372 2609
rect 486 2613 492 2614
rect 486 2609 487 2613
rect 491 2609 492 2613
rect 486 2608 492 2609
rect 614 2613 620 2614
rect 614 2609 615 2613
rect 619 2609 620 2613
rect 614 2608 620 2609
rect 750 2613 756 2614
rect 750 2609 751 2613
rect 755 2609 756 2613
rect 750 2608 756 2609
rect 894 2613 900 2614
rect 894 2609 895 2613
rect 899 2609 900 2613
rect 894 2608 900 2609
rect 1030 2613 1036 2614
rect 1030 2609 1031 2613
rect 1035 2609 1036 2613
rect 1030 2608 1036 2609
rect 1166 2613 1172 2614
rect 1166 2609 1167 2613
rect 1171 2609 1172 2613
rect 1166 2608 1172 2609
rect 1302 2613 1308 2614
rect 1302 2609 1303 2613
rect 1307 2609 1308 2613
rect 1302 2608 1308 2609
rect 1430 2613 1436 2614
rect 1430 2609 1431 2613
rect 1435 2609 1436 2613
rect 1430 2608 1436 2609
rect 1566 2613 1572 2614
rect 1566 2609 1567 2613
rect 1571 2609 1572 2613
rect 1566 2608 1572 2609
rect 1702 2613 1708 2614
rect 1702 2609 1703 2613
rect 1707 2609 1708 2613
rect 1702 2608 1708 2609
rect 2006 2612 2012 2613
rect 2006 2608 2007 2612
rect 2011 2608 2012 2612
rect 2642 2611 2648 2612
rect 110 2607 116 2608
rect 2006 2607 2012 2608
rect 2306 2607 2312 2608
rect 2046 2603 2052 2604
rect 2046 2599 2047 2603
rect 2051 2599 2052 2603
rect 2306 2603 2307 2607
rect 2311 2603 2312 2607
rect 2306 2602 2312 2603
rect 2410 2607 2416 2608
rect 2410 2603 2411 2607
rect 2415 2603 2416 2607
rect 2410 2602 2416 2603
rect 2522 2607 2528 2608
rect 2522 2603 2523 2607
rect 2527 2603 2528 2607
rect 2522 2602 2528 2603
rect 2634 2607 2640 2608
rect 2634 2603 2635 2607
rect 2639 2603 2640 2607
rect 2642 2607 2643 2611
rect 2647 2610 2648 2611
rect 2782 2611 2788 2612
rect 2647 2608 2713 2610
rect 2647 2607 2648 2608
rect 2642 2606 2648 2607
rect 2782 2607 2783 2611
rect 2787 2610 2788 2611
rect 2879 2611 2885 2612
rect 2787 2608 2833 2610
rect 2787 2607 2788 2608
rect 2782 2606 2788 2607
rect 2879 2607 2880 2611
rect 2884 2610 2885 2611
rect 3114 2611 3120 2612
rect 2884 2608 2953 2610
rect 2884 2607 2885 2608
rect 2879 2606 2885 2607
rect 3106 2607 3112 2608
rect 2634 2602 2640 2603
rect 3106 2603 3107 2607
rect 3111 2603 3112 2607
rect 3114 2607 3115 2611
rect 3119 2610 3120 2611
rect 3119 2608 3193 2610
rect 3119 2607 3120 2608
rect 3114 2606 3120 2607
rect 3106 2602 3112 2603
rect 3942 2603 3948 2604
rect 2046 2598 2052 2599
rect 2230 2600 2236 2601
rect 2230 2596 2231 2600
rect 2235 2596 2236 2600
rect 2230 2595 2236 2596
rect 2334 2600 2340 2601
rect 2334 2596 2335 2600
rect 2339 2596 2340 2600
rect 2334 2595 2340 2596
rect 2446 2600 2452 2601
rect 2446 2596 2447 2600
rect 2451 2596 2452 2600
rect 2446 2595 2452 2596
rect 2558 2600 2564 2601
rect 2558 2596 2559 2600
rect 2563 2596 2564 2600
rect 2558 2595 2564 2596
rect 2670 2600 2676 2601
rect 2670 2596 2671 2600
rect 2675 2596 2676 2600
rect 2670 2595 2676 2596
rect 2790 2600 2796 2601
rect 2790 2596 2791 2600
rect 2795 2596 2796 2600
rect 2790 2595 2796 2596
rect 2910 2600 2916 2601
rect 2910 2596 2911 2600
rect 2915 2596 2916 2600
rect 2910 2595 2916 2596
rect 3030 2600 3036 2601
rect 3030 2596 3031 2600
rect 3035 2596 3036 2600
rect 3030 2595 3036 2596
rect 3150 2600 3156 2601
rect 3150 2596 3151 2600
rect 3155 2596 3156 2600
rect 3942 2599 3943 2603
rect 3947 2599 3948 2603
rect 3942 2598 3948 2599
rect 3150 2595 3156 2596
rect 2538 2587 2544 2588
rect 2538 2586 2539 2587
rect 2300 2584 2539 2586
rect 2283 2579 2289 2580
rect 2283 2575 2284 2579
rect 2288 2578 2289 2579
rect 2300 2578 2302 2584
rect 2538 2583 2539 2584
rect 2543 2583 2544 2587
rect 3114 2587 3120 2588
rect 3114 2586 3115 2587
rect 2538 2582 2544 2583
rect 3060 2584 3115 2586
rect 2288 2576 2302 2578
rect 2306 2579 2312 2580
rect 2288 2575 2289 2576
rect 2283 2574 2289 2575
rect 2306 2575 2307 2579
rect 2311 2578 2312 2579
rect 2387 2579 2393 2580
rect 2387 2578 2388 2579
rect 2311 2576 2388 2578
rect 2311 2575 2312 2576
rect 2306 2574 2312 2575
rect 2387 2575 2388 2576
rect 2392 2575 2393 2579
rect 2387 2574 2393 2575
rect 2410 2579 2416 2580
rect 2410 2575 2411 2579
rect 2415 2578 2416 2579
rect 2499 2579 2505 2580
rect 2499 2578 2500 2579
rect 2415 2576 2500 2578
rect 2415 2575 2416 2576
rect 2410 2574 2416 2575
rect 2499 2575 2500 2576
rect 2504 2575 2505 2579
rect 2499 2574 2505 2575
rect 2522 2579 2528 2580
rect 2522 2575 2523 2579
rect 2527 2578 2528 2579
rect 2611 2579 2617 2580
rect 2611 2578 2612 2579
rect 2527 2576 2612 2578
rect 2527 2575 2528 2576
rect 2522 2574 2528 2575
rect 2611 2575 2612 2576
rect 2616 2575 2617 2579
rect 2611 2574 2617 2575
rect 2634 2579 2640 2580
rect 2634 2575 2635 2579
rect 2639 2578 2640 2579
rect 2723 2579 2729 2580
rect 2723 2578 2724 2579
rect 2639 2576 2724 2578
rect 2639 2575 2640 2576
rect 2634 2574 2640 2575
rect 2723 2575 2724 2576
rect 2728 2575 2729 2579
rect 2723 2574 2729 2575
rect 2843 2579 2849 2580
rect 2843 2575 2844 2579
rect 2848 2578 2849 2579
rect 2879 2579 2885 2580
rect 2879 2578 2880 2579
rect 2848 2576 2880 2578
rect 2848 2575 2849 2576
rect 2843 2574 2849 2575
rect 2879 2575 2880 2576
rect 2884 2575 2885 2579
rect 2879 2574 2885 2575
rect 2963 2579 2969 2580
rect 2963 2575 2964 2579
rect 2968 2578 2969 2579
rect 3060 2578 3062 2584
rect 3114 2583 3115 2584
rect 3119 2583 3120 2587
rect 3114 2582 3120 2583
rect 2968 2576 3062 2578
rect 3106 2579 3112 2580
rect 2968 2575 2969 2576
rect 2963 2574 2969 2575
rect 3066 2575 3072 2576
rect 3066 2571 3067 2575
rect 3071 2574 3072 2575
rect 3083 2575 3089 2576
rect 3083 2574 3084 2575
rect 3071 2572 3084 2574
rect 3071 2571 3072 2572
rect 3066 2570 3072 2571
rect 3083 2571 3084 2572
rect 3088 2571 3089 2575
rect 3106 2575 3107 2579
rect 3111 2578 3112 2579
rect 3203 2579 3209 2580
rect 3203 2578 3204 2579
rect 3111 2576 3204 2578
rect 3111 2575 3112 2576
rect 3106 2574 3112 2575
rect 3203 2575 3204 2576
rect 3208 2575 3209 2579
rect 3203 2574 3209 2575
rect 3083 2570 3089 2571
rect 2642 2567 2648 2568
rect 2642 2566 2643 2567
rect 2436 2564 2643 2566
rect 2436 2562 2438 2564
rect 2642 2563 2643 2564
rect 2647 2563 2648 2567
rect 2642 2562 2648 2563
rect 2435 2561 2441 2562
rect 110 2560 116 2561
rect 2006 2560 2012 2561
rect 110 2556 111 2560
rect 115 2556 116 2560
rect 110 2555 116 2556
rect 134 2559 140 2560
rect 134 2555 135 2559
rect 139 2555 140 2559
rect 134 2554 140 2555
rect 286 2559 292 2560
rect 286 2555 287 2559
rect 291 2555 292 2559
rect 286 2554 292 2555
rect 446 2559 452 2560
rect 446 2555 447 2559
rect 451 2555 452 2559
rect 446 2554 452 2555
rect 606 2559 612 2560
rect 606 2555 607 2559
rect 611 2555 612 2559
rect 606 2554 612 2555
rect 766 2559 772 2560
rect 766 2555 767 2559
rect 771 2555 772 2559
rect 766 2554 772 2555
rect 918 2559 924 2560
rect 918 2555 919 2559
rect 923 2555 924 2559
rect 918 2554 924 2555
rect 1062 2559 1068 2560
rect 1062 2555 1063 2559
rect 1067 2555 1068 2559
rect 1062 2554 1068 2555
rect 1198 2559 1204 2560
rect 1198 2555 1199 2559
rect 1203 2555 1204 2559
rect 1198 2554 1204 2555
rect 1334 2559 1340 2560
rect 1334 2555 1335 2559
rect 1339 2555 1340 2559
rect 1334 2554 1340 2555
rect 1462 2559 1468 2560
rect 1462 2555 1463 2559
rect 1467 2555 1468 2559
rect 1462 2554 1468 2555
rect 1590 2559 1596 2560
rect 1590 2555 1591 2559
rect 1595 2555 1596 2559
rect 1590 2554 1596 2555
rect 1726 2559 1732 2560
rect 1726 2555 1727 2559
rect 1731 2555 1732 2559
rect 2006 2556 2007 2560
rect 2011 2556 2012 2560
rect 2435 2557 2436 2561
rect 2440 2557 2441 2561
rect 2435 2556 2441 2557
rect 2458 2559 2464 2560
rect 2006 2555 2012 2556
rect 2458 2555 2459 2559
rect 2463 2558 2464 2559
rect 2547 2559 2553 2560
rect 2547 2558 2548 2559
rect 2463 2556 2548 2558
rect 2463 2555 2464 2556
rect 1726 2554 1732 2555
rect 2458 2554 2464 2555
rect 2547 2555 2548 2556
rect 2552 2555 2553 2559
rect 2547 2554 2553 2555
rect 2570 2559 2576 2560
rect 2570 2555 2571 2559
rect 2575 2558 2576 2559
rect 2667 2559 2673 2560
rect 2667 2558 2668 2559
rect 2575 2556 2668 2558
rect 2575 2555 2576 2556
rect 2570 2554 2576 2555
rect 2667 2555 2668 2556
rect 2672 2555 2673 2559
rect 2667 2554 2673 2555
rect 2690 2559 2696 2560
rect 2690 2555 2691 2559
rect 2695 2558 2696 2559
rect 2795 2559 2801 2560
rect 2795 2558 2796 2559
rect 2695 2556 2796 2558
rect 2695 2555 2696 2556
rect 2690 2554 2696 2555
rect 2795 2555 2796 2556
rect 2800 2555 2801 2559
rect 2795 2554 2801 2555
rect 2818 2559 2824 2560
rect 2818 2555 2819 2559
rect 2823 2558 2824 2559
rect 2923 2559 2929 2560
rect 2923 2558 2924 2559
rect 2823 2556 2924 2558
rect 2823 2555 2824 2556
rect 2818 2554 2824 2555
rect 2923 2555 2924 2556
rect 2928 2555 2929 2559
rect 2923 2554 2929 2555
rect 3043 2559 3049 2560
rect 3043 2555 3044 2559
rect 3048 2558 3049 2559
rect 3074 2559 3080 2560
rect 3074 2558 3075 2559
rect 3048 2556 3075 2558
rect 3048 2555 3049 2556
rect 3043 2554 3049 2555
rect 3074 2555 3075 2556
rect 3079 2555 3080 2559
rect 3074 2554 3080 2555
rect 3163 2559 3169 2560
rect 3163 2555 3164 2559
rect 3168 2558 3169 2559
rect 3194 2559 3200 2560
rect 3194 2558 3195 2559
rect 3168 2556 3195 2558
rect 3168 2555 3169 2556
rect 3163 2554 3169 2555
rect 3194 2555 3195 2556
rect 3199 2555 3200 2559
rect 3194 2554 3200 2555
rect 3283 2559 3289 2560
rect 3283 2555 3284 2559
rect 3288 2558 3289 2559
rect 3314 2559 3320 2560
rect 3314 2558 3315 2559
rect 3288 2556 3315 2558
rect 3288 2555 3289 2556
rect 3283 2554 3289 2555
rect 3314 2555 3315 2556
rect 3319 2555 3320 2559
rect 3314 2554 3320 2555
rect 3411 2559 3417 2560
rect 3411 2555 3412 2559
rect 3416 2558 3417 2559
rect 3442 2559 3448 2560
rect 3442 2558 3443 2559
rect 3416 2556 3443 2558
rect 3416 2555 3417 2556
rect 3411 2554 3417 2555
rect 3442 2555 3443 2556
rect 3447 2555 3448 2559
rect 3442 2554 3448 2555
rect 3539 2557 3545 2558
rect 3539 2553 3540 2557
rect 3544 2553 3545 2557
rect 3539 2552 3545 2553
rect 738 2551 744 2552
rect 210 2547 216 2548
rect 110 2543 116 2544
rect 110 2539 111 2543
rect 115 2539 116 2543
rect 210 2543 211 2547
rect 215 2543 216 2547
rect 210 2542 216 2543
rect 362 2547 368 2548
rect 362 2543 363 2547
rect 367 2543 368 2547
rect 362 2542 368 2543
rect 522 2547 528 2548
rect 522 2543 523 2547
rect 527 2543 528 2547
rect 522 2542 528 2543
rect 682 2547 688 2548
rect 682 2543 683 2547
rect 687 2543 688 2547
rect 738 2547 739 2551
rect 743 2550 744 2551
rect 1802 2551 1808 2552
rect 743 2548 809 2550
rect 743 2547 744 2548
rect 738 2546 744 2547
rect 994 2547 1000 2548
rect 682 2542 688 2543
rect 994 2543 995 2547
rect 999 2543 1000 2547
rect 994 2542 1000 2543
rect 1138 2547 1144 2548
rect 1138 2543 1139 2547
rect 1143 2543 1144 2547
rect 1138 2542 1144 2543
rect 1274 2547 1280 2548
rect 1274 2543 1275 2547
rect 1279 2543 1280 2547
rect 1274 2542 1280 2543
rect 1410 2547 1416 2548
rect 1410 2543 1411 2547
rect 1415 2543 1416 2547
rect 1410 2542 1416 2543
rect 1538 2547 1544 2548
rect 1538 2543 1539 2547
rect 1543 2543 1544 2547
rect 1538 2542 1544 2543
rect 1666 2547 1672 2548
rect 1666 2543 1667 2547
rect 1671 2543 1672 2547
rect 1802 2547 1803 2551
rect 1807 2547 1808 2551
rect 1802 2546 1808 2547
rect 3434 2551 3440 2552
rect 3434 2547 3435 2551
rect 3439 2550 3440 2551
rect 3540 2550 3542 2552
rect 3439 2548 3542 2550
rect 3439 2547 3440 2548
rect 3434 2546 3440 2547
rect 1666 2542 1672 2543
rect 2006 2543 2012 2544
rect 110 2538 116 2539
rect 134 2540 140 2541
rect 134 2536 135 2540
rect 139 2536 140 2540
rect 134 2535 140 2536
rect 286 2540 292 2541
rect 286 2536 287 2540
rect 291 2536 292 2540
rect 286 2535 292 2536
rect 446 2540 452 2541
rect 446 2536 447 2540
rect 451 2536 452 2540
rect 446 2535 452 2536
rect 606 2540 612 2541
rect 606 2536 607 2540
rect 611 2536 612 2540
rect 606 2535 612 2536
rect 766 2540 772 2541
rect 766 2536 767 2540
rect 771 2536 772 2540
rect 766 2535 772 2536
rect 918 2540 924 2541
rect 918 2536 919 2540
rect 923 2536 924 2540
rect 918 2535 924 2536
rect 1062 2540 1068 2541
rect 1062 2536 1063 2540
rect 1067 2536 1068 2540
rect 1062 2535 1068 2536
rect 1198 2540 1204 2541
rect 1198 2536 1199 2540
rect 1203 2536 1204 2540
rect 1198 2535 1204 2536
rect 1334 2540 1340 2541
rect 1334 2536 1335 2540
rect 1339 2536 1340 2540
rect 1334 2535 1340 2536
rect 1462 2540 1468 2541
rect 1462 2536 1463 2540
rect 1467 2536 1468 2540
rect 1462 2535 1468 2536
rect 1590 2540 1596 2541
rect 1590 2536 1591 2540
rect 1595 2536 1596 2540
rect 1590 2535 1596 2536
rect 1726 2540 1732 2541
rect 1726 2536 1727 2540
rect 1731 2536 1732 2540
rect 2006 2539 2007 2543
rect 2011 2539 2012 2543
rect 2006 2538 2012 2539
rect 1726 2535 1732 2536
rect 2382 2536 2388 2537
rect 2046 2533 2052 2534
rect 2046 2529 2047 2533
rect 2051 2529 2052 2533
rect 2382 2532 2383 2536
rect 2387 2532 2388 2536
rect 2382 2531 2388 2532
rect 2494 2536 2500 2537
rect 2494 2532 2495 2536
rect 2499 2532 2500 2536
rect 2494 2531 2500 2532
rect 2614 2536 2620 2537
rect 2614 2532 2615 2536
rect 2619 2532 2620 2536
rect 2614 2531 2620 2532
rect 2742 2536 2748 2537
rect 2742 2532 2743 2536
rect 2747 2532 2748 2536
rect 2742 2531 2748 2532
rect 2870 2536 2876 2537
rect 2870 2532 2871 2536
rect 2875 2532 2876 2536
rect 2870 2531 2876 2532
rect 2990 2536 2996 2537
rect 2990 2532 2991 2536
rect 2995 2532 2996 2536
rect 2990 2531 2996 2532
rect 3110 2536 3116 2537
rect 3110 2532 3111 2536
rect 3115 2532 3116 2536
rect 3110 2531 3116 2532
rect 3230 2536 3236 2537
rect 3230 2532 3231 2536
rect 3235 2532 3236 2536
rect 3230 2531 3236 2532
rect 3358 2536 3364 2537
rect 3358 2532 3359 2536
rect 3363 2532 3364 2536
rect 3358 2531 3364 2532
rect 3486 2536 3492 2537
rect 3486 2532 3487 2536
rect 3491 2532 3492 2536
rect 3486 2531 3492 2532
rect 3942 2533 3948 2534
rect 2046 2528 2052 2529
rect 3942 2529 3943 2533
rect 3947 2529 3948 2533
rect 3942 2528 3948 2529
rect 2458 2527 2464 2528
rect 210 2523 216 2524
rect 210 2519 211 2523
rect 215 2519 216 2523
rect 2458 2523 2459 2527
rect 2463 2523 2464 2527
rect 2458 2522 2464 2523
rect 2570 2527 2576 2528
rect 2570 2523 2571 2527
rect 2575 2523 2576 2527
rect 2570 2522 2576 2523
rect 2690 2527 2696 2528
rect 2690 2523 2691 2527
rect 2695 2523 2696 2527
rect 2690 2522 2696 2523
rect 2818 2527 2824 2528
rect 2818 2523 2819 2527
rect 2823 2523 2824 2527
rect 2818 2522 2824 2523
rect 2826 2527 2832 2528
rect 2826 2523 2827 2527
rect 2831 2526 2832 2527
rect 3066 2527 3072 2528
rect 2831 2524 2913 2526
rect 2831 2523 2832 2524
rect 2826 2522 2832 2523
rect 3066 2523 3067 2527
rect 3071 2523 3072 2527
rect 3066 2522 3072 2523
rect 3074 2527 3080 2528
rect 3074 2523 3075 2527
rect 3079 2526 3080 2527
rect 3194 2527 3200 2528
rect 3079 2524 3153 2526
rect 3079 2523 3080 2524
rect 3074 2522 3080 2523
rect 3194 2523 3195 2527
rect 3199 2526 3200 2527
rect 3314 2527 3320 2528
rect 3199 2524 3273 2526
rect 3199 2523 3200 2524
rect 3194 2522 3200 2523
rect 3314 2523 3315 2527
rect 3319 2526 3320 2527
rect 3442 2527 3448 2528
rect 3319 2524 3401 2526
rect 3319 2523 3320 2524
rect 3314 2522 3320 2523
rect 3442 2523 3443 2527
rect 3447 2526 3448 2527
rect 3447 2524 3529 2526
rect 3447 2523 3448 2524
rect 3442 2522 3448 2523
rect 210 2518 216 2519
rect 339 2519 345 2520
rect 339 2518 340 2519
rect 212 2516 340 2518
rect 187 2515 193 2516
rect 187 2511 188 2515
rect 192 2514 193 2515
rect 339 2515 340 2516
rect 344 2515 345 2519
rect 339 2514 345 2515
rect 362 2519 368 2520
rect 362 2515 363 2519
rect 367 2518 368 2519
rect 499 2519 505 2520
rect 499 2518 500 2519
rect 367 2516 500 2518
rect 367 2515 368 2516
rect 362 2514 368 2515
rect 499 2515 500 2516
rect 504 2515 505 2519
rect 499 2514 505 2515
rect 522 2519 528 2520
rect 522 2515 523 2519
rect 527 2518 528 2519
rect 659 2519 665 2520
rect 659 2518 660 2519
rect 527 2516 660 2518
rect 527 2515 528 2516
rect 522 2514 528 2515
rect 659 2515 660 2516
rect 664 2515 665 2519
rect 659 2514 665 2515
rect 682 2519 688 2520
rect 682 2515 683 2519
rect 687 2518 688 2519
rect 819 2519 825 2520
rect 819 2518 820 2519
rect 687 2516 820 2518
rect 687 2515 688 2516
rect 682 2514 688 2515
rect 819 2515 820 2516
rect 824 2515 825 2519
rect 819 2514 825 2515
rect 971 2519 980 2520
rect 971 2515 972 2519
rect 979 2515 980 2519
rect 971 2514 980 2515
rect 994 2519 1000 2520
rect 994 2515 995 2519
rect 999 2518 1000 2519
rect 1115 2519 1121 2520
rect 1115 2518 1116 2519
rect 999 2516 1116 2518
rect 999 2515 1000 2516
rect 994 2514 1000 2515
rect 1115 2515 1116 2516
rect 1120 2515 1121 2519
rect 1115 2514 1121 2515
rect 1138 2519 1144 2520
rect 1138 2515 1139 2519
rect 1143 2518 1144 2519
rect 1251 2519 1257 2520
rect 1251 2518 1252 2519
rect 1143 2516 1252 2518
rect 1143 2515 1144 2516
rect 1138 2514 1144 2515
rect 1251 2515 1252 2516
rect 1256 2515 1257 2519
rect 1251 2514 1257 2515
rect 1274 2519 1280 2520
rect 1274 2515 1275 2519
rect 1279 2518 1280 2519
rect 1387 2519 1393 2520
rect 1387 2518 1388 2519
rect 1279 2516 1388 2518
rect 1279 2515 1280 2516
rect 1274 2514 1280 2515
rect 1387 2515 1388 2516
rect 1392 2515 1393 2519
rect 1387 2514 1393 2515
rect 1410 2519 1416 2520
rect 1410 2515 1411 2519
rect 1415 2518 1416 2519
rect 1515 2519 1521 2520
rect 1515 2518 1516 2519
rect 1415 2516 1516 2518
rect 1415 2515 1416 2516
rect 1410 2514 1416 2515
rect 1515 2515 1516 2516
rect 1520 2515 1521 2519
rect 1515 2514 1521 2515
rect 1538 2519 1544 2520
rect 1538 2515 1539 2519
rect 1543 2518 1544 2519
rect 1643 2519 1649 2520
rect 1643 2518 1644 2519
rect 1543 2516 1644 2518
rect 1543 2515 1544 2516
rect 1538 2514 1544 2515
rect 1643 2515 1644 2516
rect 1648 2515 1649 2519
rect 1643 2514 1649 2515
rect 1666 2519 1672 2520
rect 1666 2515 1667 2519
rect 1671 2518 1672 2519
rect 1779 2519 1785 2520
rect 1779 2518 1780 2519
rect 1671 2516 1780 2518
rect 1671 2515 1672 2516
rect 1666 2514 1672 2515
rect 1779 2515 1780 2516
rect 1784 2515 1785 2519
rect 2382 2517 2388 2518
rect 1779 2514 1785 2515
rect 2046 2516 2052 2517
rect 192 2512 321 2514
rect 2046 2512 2047 2516
rect 2051 2512 2052 2516
rect 2382 2513 2383 2517
rect 2387 2513 2388 2517
rect 2382 2512 2388 2513
rect 2494 2517 2500 2518
rect 2494 2513 2495 2517
rect 2499 2513 2500 2517
rect 2494 2512 2500 2513
rect 2614 2517 2620 2518
rect 2614 2513 2615 2517
rect 2619 2513 2620 2517
rect 2614 2512 2620 2513
rect 2742 2517 2748 2518
rect 2742 2513 2743 2517
rect 2747 2513 2748 2517
rect 2742 2512 2748 2513
rect 2870 2517 2876 2518
rect 2870 2513 2871 2517
rect 2875 2513 2876 2517
rect 2870 2512 2876 2513
rect 2990 2517 2996 2518
rect 2990 2513 2991 2517
rect 2995 2513 2996 2517
rect 2990 2512 2996 2513
rect 3110 2517 3116 2518
rect 3110 2513 3111 2517
rect 3115 2513 3116 2517
rect 3110 2512 3116 2513
rect 3230 2517 3236 2518
rect 3230 2513 3231 2517
rect 3235 2513 3236 2517
rect 3230 2512 3236 2513
rect 3358 2517 3364 2518
rect 3358 2513 3359 2517
rect 3363 2513 3364 2517
rect 3358 2512 3364 2513
rect 3486 2517 3492 2518
rect 3486 2513 3487 2517
rect 3491 2513 3492 2517
rect 3486 2512 3492 2513
rect 3942 2516 3948 2517
rect 3942 2512 3943 2516
rect 3947 2512 3948 2516
rect 192 2511 193 2512
rect 187 2510 193 2511
rect 319 2510 321 2512
rect 506 2511 512 2512
rect 2046 2511 2052 2512
rect 3942 2511 3948 2512
rect 506 2510 507 2511
rect 319 2508 507 2510
rect 506 2507 507 2508
rect 511 2507 512 2511
rect 506 2506 512 2507
rect 187 2487 193 2488
rect 187 2483 188 2487
rect 192 2486 193 2487
rect 202 2487 208 2488
rect 202 2486 203 2487
rect 192 2484 203 2486
rect 192 2483 193 2484
rect 187 2482 193 2483
rect 202 2483 203 2484
rect 207 2483 208 2487
rect 202 2482 208 2483
rect 210 2487 216 2488
rect 210 2483 211 2487
rect 215 2486 216 2487
rect 283 2487 289 2488
rect 283 2486 284 2487
rect 215 2484 284 2486
rect 215 2483 216 2484
rect 210 2482 216 2483
rect 283 2483 284 2484
rect 288 2483 289 2487
rect 283 2482 289 2483
rect 306 2487 312 2488
rect 306 2483 307 2487
rect 311 2486 312 2487
rect 379 2487 385 2488
rect 379 2486 380 2487
rect 311 2484 380 2486
rect 311 2483 312 2484
rect 306 2482 312 2483
rect 379 2483 380 2484
rect 384 2483 385 2487
rect 379 2482 385 2483
rect 402 2487 408 2488
rect 402 2483 403 2487
rect 407 2486 408 2487
rect 475 2487 481 2488
rect 475 2486 476 2487
rect 407 2484 476 2486
rect 407 2483 408 2484
rect 402 2482 408 2483
rect 475 2483 476 2484
rect 480 2483 481 2487
rect 475 2482 481 2483
rect 498 2487 504 2488
rect 498 2483 499 2487
rect 503 2486 504 2487
rect 571 2487 577 2488
rect 571 2486 572 2487
rect 503 2484 572 2486
rect 503 2483 504 2484
rect 498 2482 504 2483
rect 571 2483 572 2484
rect 576 2483 577 2487
rect 571 2482 577 2483
rect 134 2464 140 2465
rect 110 2461 116 2462
rect 110 2457 111 2461
rect 115 2457 116 2461
rect 134 2460 135 2464
rect 139 2460 140 2464
rect 134 2459 140 2460
rect 230 2464 236 2465
rect 230 2460 231 2464
rect 235 2460 236 2464
rect 230 2459 236 2460
rect 326 2464 332 2465
rect 326 2460 327 2464
rect 331 2460 332 2464
rect 326 2459 332 2460
rect 422 2464 428 2465
rect 422 2460 423 2464
rect 427 2460 428 2464
rect 422 2459 428 2460
rect 518 2464 524 2465
rect 518 2460 519 2464
rect 523 2460 524 2464
rect 518 2459 524 2460
rect 2006 2461 2012 2462
rect 110 2456 116 2457
rect 2006 2457 2007 2461
rect 2011 2457 2012 2461
rect 2006 2456 2012 2457
rect 2046 2460 2052 2461
rect 3942 2460 3948 2461
rect 2046 2456 2047 2460
rect 2051 2456 2052 2460
rect 210 2455 216 2456
rect 210 2451 211 2455
rect 215 2451 216 2455
rect 210 2450 216 2451
rect 306 2455 312 2456
rect 306 2451 307 2455
rect 311 2451 312 2455
rect 306 2450 312 2451
rect 402 2455 408 2456
rect 402 2451 403 2455
rect 407 2451 408 2455
rect 402 2450 408 2451
rect 498 2455 504 2456
rect 498 2451 499 2455
rect 503 2451 504 2455
rect 498 2450 504 2451
rect 506 2455 512 2456
rect 2046 2455 2052 2456
rect 2534 2459 2540 2460
rect 2534 2455 2535 2459
rect 2539 2455 2540 2459
rect 506 2451 507 2455
rect 511 2454 512 2455
rect 2534 2454 2540 2455
rect 2710 2459 2716 2460
rect 2710 2455 2711 2459
rect 2715 2455 2716 2459
rect 2710 2454 2716 2455
rect 2878 2459 2884 2460
rect 2878 2455 2879 2459
rect 2883 2455 2884 2459
rect 2878 2454 2884 2455
rect 3046 2459 3052 2460
rect 3046 2455 3047 2459
rect 3051 2455 3052 2459
rect 3046 2454 3052 2455
rect 3206 2459 3212 2460
rect 3206 2455 3207 2459
rect 3211 2455 3212 2459
rect 3206 2454 3212 2455
rect 3358 2459 3364 2460
rect 3358 2455 3359 2459
rect 3363 2455 3364 2459
rect 3358 2454 3364 2455
rect 3502 2459 3508 2460
rect 3502 2455 3503 2459
rect 3507 2455 3508 2459
rect 3502 2454 3508 2455
rect 3654 2459 3660 2460
rect 3654 2455 3655 2459
rect 3659 2455 3660 2459
rect 3654 2454 3660 2455
rect 3806 2459 3812 2460
rect 3806 2455 3807 2459
rect 3811 2455 3812 2459
rect 3942 2456 3943 2460
rect 3947 2456 3948 2460
rect 3942 2455 3948 2456
rect 3806 2454 3812 2455
rect 511 2452 561 2454
rect 511 2451 512 2452
rect 506 2450 512 2451
rect 3434 2451 3440 2452
rect 2610 2447 2616 2448
rect 134 2445 140 2446
rect 110 2444 116 2445
rect 110 2440 111 2444
rect 115 2440 116 2444
rect 134 2441 135 2445
rect 139 2441 140 2445
rect 134 2440 140 2441
rect 230 2445 236 2446
rect 230 2441 231 2445
rect 235 2441 236 2445
rect 230 2440 236 2441
rect 326 2445 332 2446
rect 326 2441 327 2445
rect 331 2441 332 2445
rect 326 2440 332 2441
rect 422 2445 428 2446
rect 422 2441 423 2445
rect 427 2441 428 2445
rect 422 2440 428 2441
rect 518 2445 524 2446
rect 518 2441 519 2445
rect 523 2441 524 2445
rect 518 2440 524 2441
rect 2006 2444 2012 2445
rect 2006 2440 2007 2444
rect 2011 2440 2012 2444
rect 110 2439 116 2440
rect 2006 2439 2012 2440
rect 2046 2443 2052 2444
rect 2046 2439 2047 2443
rect 2051 2439 2052 2443
rect 2610 2443 2611 2447
rect 2615 2443 2616 2447
rect 2610 2442 2616 2443
rect 2786 2447 2792 2448
rect 2786 2443 2787 2447
rect 2791 2443 2792 2447
rect 2786 2442 2792 2443
rect 2954 2447 2960 2448
rect 2954 2443 2955 2447
rect 2959 2443 2960 2447
rect 2954 2442 2960 2443
rect 3122 2447 3128 2448
rect 3122 2443 3123 2447
rect 3127 2443 3128 2447
rect 3122 2442 3128 2443
rect 3282 2447 3288 2448
rect 3282 2443 3283 2447
rect 3287 2443 3288 2447
rect 3434 2447 3435 2451
rect 3439 2447 3440 2451
rect 3434 2446 3440 2447
rect 3442 2451 3448 2452
rect 3442 2447 3443 2451
rect 3447 2450 3448 2451
rect 3586 2451 3592 2452
rect 3447 2448 3545 2450
rect 3447 2447 3448 2448
rect 3442 2446 3448 2447
rect 3586 2447 3587 2451
rect 3591 2450 3592 2451
rect 3751 2451 3757 2452
rect 3591 2448 3697 2450
rect 3591 2447 3592 2448
rect 3586 2446 3592 2447
rect 3751 2447 3752 2451
rect 3756 2450 3757 2451
rect 3756 2448 3849 2450
rect 3756 2447 3757 2448
rect 3751 2446 3757 2447
rect 3282 2442 3288 2443
rect 3942 2443 3948 2444
rect 2046 2438 2052 2439
rect 2534 2440 2540 2441
rect 2534 2436 2535 2440
rect 2539 2436 2540 2440
rect 2534 2435 2540 2436
rect 2710 2440 2716 2441
rect 2710 2436 2711 2440
rect 2715 2436 2716 2440
rect 2710 2435 2716 2436
rect 2878 2440 2884 2441
rect 2878 2436 2879 2440
rect 2883 2436 2884 2440
rect 2878 2435 2884 2436
rect 3046 2440 3052 2441
rect 3046 2436 3047 2440
rect 3051 2436 3052 2440
rect 3046 2435 3052 2436
rect 3206 2440 3212 2441
rect 3206 2436 3207 2440
rect 3211 2436 3212 2440
rect 3206 2435 3212 2436
rect 3358 2440 3364 2441
rect 3358 2436 3359 2440
rect 3363 2436 3364 2440
rect 3358 2435 3364 2436
rect 3502 2440 3508 2441
rect 3502 2436 3503 2440
rect 3507 2436 3508 2440
rect 3502 2435 3508 2436
rect 3654 2440 3660 2441
rect 3654 2436 3655 2440
rect 3659 2436 3660 2440
rect 3654 2435 3660 2436
rect 3806 2440 3812 2441
rect 3806 2436 3807 2440
rect 3811 2436 3812 2440
rect 3942 2439 3943 2443
rect 3947 2439 3948 2443
rect 3942 2438 3948 2439
rect 3806 2435 3812 2436
rect 2826 2427 2832 2428
rect 2826 2426 2827 2427
rect 2604 2424 2827 2426
rect 2587 2419 2593 2420
rect 2587 2415 2588 2419
rect 2592 2418 2593 2419
rect 2604 2418 2606 2424
rect 2826 2423 2827 2424
rect 2831 2423 2832 2427
rect 3442 2427 3448 2428
rect 3442 2426 3443 2427
rect 2826 2422 2832 2423
rect 3276 2424 3443 2426
rect 2592 2416 2606 2418
rect 2610 2419 2616 2420
rect 2592 2415 2593 2416
rect 2587 2414 2593 2415
rect 2610 2415 2611 2419
rect 2615 2418 2616 2419
rect 2763 2419 2769 2420
rect 2763 2418 2764 2419
rect 2615 2416 2764 2418
rect 2615 2415 2616 2416
rect 2610 2414 2616 2415
rect 2763 2415 2764 2416
rect 2768 2415 2769 2419
rect 2763 2414 2769 2415
rect 2786 2419 2792 2420
rect 2786 2415 2787 2419
rect 2791 2418 2792 2419
rect 2931 2419 2937 2420
rect 2931 2418 2932 2419
rect 2791 2416 2932 2418
rect 2791 2415 2792 2416
rect 2786 2414 2792 2415
rect 2931 2415 2932 2416
rect 2936 2415 2937 2419
rect 2931 2414 2937 2415
rect 2954 2419 2960 2420
rect 2954 2415 2955 2419
rect 2959 2418 2960 2419
rect 3099 2419 3105 2420
rect 3099 2418 3100 2419
rect 2959 2416 3100 2418
rect 2959 2415 2960 2416
rect 2954 2414 2960 2415
rect 3099 2415 3100 2416
rect 3104 2415 3105 2419
rect 3099 2414 3105 2415
rect 3259 2419 3265 2420
rect 3259 2415 3260 2419
rect 3264 2418 3265 2419
rect 3276 2418 3278 2424
rect 3442 2423 3443 2424
rect 3447 2423 3448 2427
rect 3442 2422 3448 2423
rect 3264 2416 3278 2418
rect 3282 2419 3288 2420
rect 3264 2415 3265 2416
rect 3259 2414 3265 2415
rect 3282 2415 3283 2419
rect 3287 2418 3288 2419
rect 3411 2419 3417 2420
rect 3411 2418 3412 2419
rect 3287 2416 3412 2418
rect 3287 2415 3288 2416
rect 3282 2414 3288 2415
rect 3411 2415 3412 2416
rect 3416 2415 3417 2419
rect 3411 2414 3417 2415
rect 3555 2419 3561 2420
rect 3555 2415 3556 2419
rect 3560 2418 3561 2419
rect 3586 2419 3592 2420
rect 3586 2418 3587 2419
rect 3560 2416 3587 2418
rect 3560 2415 3561 2416
rect 3555 2414 3561 2415
rect 3586 2415 3587 2416
rect 3591 2415 3592 2419
rect 3586 2414 3592 2415
rect 3707 2419 3713 2420
rect 3707 2415 3708 2419
rect 3712 2418 3713 2419
rect 3751 2419 3757 2420
rect 3751 2418 3752 2419
rect 3712 2416 3752 2418
rect 3712 2415 3713 2416
rect 3707 2414 3713 2415
rect 3751 2415 3752 2416
rect 3756 2415 3757 2419
rect 3751 2414 3757 2415
rect 3859 2415 3865 2416
rect 3859 2411 3860 2415
rect 3864 2414 3865 2415
rect 3906 2415 3912 2416
rect 3906 2414 3907 2415
rect 3864 2412 3907 2414
rect 3864 2411 3865 2412
rect 3859 2410 3865 2411
rect 3906 2411 3907 2412
rect 3911 2411 3912 2415
rect 3906 2410 3912 2411
rect 2682 2391 2688 2392
rect 2659 2389 2665 2390
rect 2659 2385 2660 2389
rect 2664 2385 2665 2389
rect 2682 2387 2683 2391
rect 2687 2390 2688 2391
rect 2867 2391 2873 2392
rect 2867 2390 2868 2391
rect 2687 2388 2868 2390
rect 2687 2387 2688 2388
rect 2682 2386 2688 2387
rect 2867 2387 2868 2388
rect 2872 2387 2873 2391
rect 2867 2386 2873 2387
rect 3059 2391 3065 2392
rect 3059 2387 3060 2391
rect 3064 2390 3065 2391
rect 3122 2391 3128 2392
rect 3122 2390 3123 2391
rect 3064 2388 3123 2390
rect 3064 2387 3065 2388
rect 3059 2386 3065 2387
rect 3122 2387 3123 2388
rect 3127 2387 3128 2391
rect 3266 2391 3272 2392
rect 3122 2386 3128 2387
rect 3243 2389 3249 2390
rect 2659 2384 2665 2385
rect 3243 2385 3244 2389
rect 3248 2385 3249 2389
rect 3266 2387 3267 2391
rect 3271 2390 3272 2391
rect 3411 2391 3417 2392
rect 3411 2390 3412 2391
rect 3271 2388 3412 2390
rect 3271 2387 3272 2388
rect 3266 2386 3272 2387
rect 3411 2387 3412 2388
rect 3416 2387 3417 2391
rect 3411 2386 3417 2387
rect 3434 2391 3440 2392
rect 3434 2387 3435 2391
rect 3439 2390 3440 2391
rect 3571 2391 3577 2392
rect 3571 2390 3572 2391
rect 3439 2388 3572 2390
rect 3439 2387 3440 2388
rect 3434 2386 3440 2387
rect 3571 2387 3572 2388
rect 3576 2387 3577 2391
rect 3571 2386 3577 2387
rect 3594 2391 3600 2392
rect 3594 2387 3595 2391
rect 3599 2390 3600 2391
rect 3731 2391 3737 2392
rect 3731 2390 3732 2391
rect 3599 2388 3732 2390
rect 3599 2387 3600 2388
rect 3594 2386 3600 2387
rect 3731 2387 3732 2388
rect 3736 2387 3737 2391
rect 3731 2386 3737 2387
rect 3754 2391 3760 2392
rect 3754 2387 3755 2391
rect 3759 2390 3760 2391
rect 3891 2391 3897 2392
rect 3891 2390 3892 2391
rect 3759 2388 3892 2390
rect 3759 2387 3760 2388
rect 3754 2386 3760 2387
rect 3891 2387 3892 2388
rect 3896 2387 3897 2391
rect 3891 2386 3897 2387
rect 3243 2384 3249 2385
rect 2660 2382 2662 2384
rect 2942 2383 2948 2384
rect 2942 2382 2943 2383
rect 2660 2380 2943 2382
rect 2942 2379 2943 2380
rect 2947 2379 2948 2383
rect 3244 2382 3246 2384
rect 3618 2383 3624 2384
rect 3618 2382 3619 2383
rect 3244 2380 3619 2382
rect 2942 2378 2948 2379
rect 3618 2379 3619 2380
rect 3623 2379 3624 2383
rect 3618 2378 3624 2379
rect 110 2376 116 2377
rect 2006 2376 2012 2377
rect 110 2372 111 2376
rect 115 2372 116 2376
rect 110 2371 116 2372
rect 134 2375 140 2376
rect 134 2371 135 2375
rect 139 2371 140 2375
rect 254 2375 260 2376
rect 134 2370 140 2371
rect 202 2371 208 2372
rect 202 2367 203 2371
rect 207 2370 208 2371
rect 254 2371 255 2375
rect 259 2371 260 2375
rect 254 2370 260 2371
rect 414 2375 420 2376
rect 414 2371 415 2375
rect 419 2371 420 2375
rect 414 2370 420 2371
rect 574 2375 580 2376
rect 574 2371 575 2375
rect 579 2371 580 2375
rect 574 2370 580 2371
rect 734 2375 740 2376
rect 734 2371 735 2375
rect 739 2371 740 2375
rect 734 2370 740 2371
rect 886 2375 892 2376
rect 886 2371 887 2375
rect 891 2371 892 2375
rect 886 2370 892 2371
rect 1038 2375 1044 2376
rect 1038 2371 1039 2375
rect 1043 2371 1044 2375
rect 1038 2370 1044 2371
rect 1182 2375 1188 2376
rect 1182 2371 1183 2375
rect 1187 2371 1188 2375
rect 1182 2370 1188 2371
rect 1326 2375 1332 2376
rect 1326 2371 1327 2375
rect 1331 2371 1332 2375
rect 1326 2370 1332 2371
rect 1478 2375 1484 2376
rect 1478 2371 1479 2375
rect 1483 2371 1484 2375
rect 2006 2372 2007 2376
rect 2011 2372 2012 2376
rect 2006 2371 2012 2372
rect 1478 2370 1484 2371
rect 207 2368 214 2370
rect 2606 2368 2612 2369
rect 207 2367 208 2368
rect 202 2366 208 2367
rect 212 2365 214 2368
rect 218 2367 224 2368
rect 218 2363 219 2367
rect 223 2366 224 2367
rect 358 2367 364 2368
rect 223 2364 297 2366
rect 223 2363 224 2364
rect 218 2362 224 2363
rect 358 2363 359 2367
rect 363 2366 364 2367
rect 510 2367 516 2368
rect 363 2364 457 2366
rect 363 2363 364 2364
rect 358 2362 364 2363
rect 510 2363 511 2367
rect 515 2366 516 2367
rect 702 2367 708 2368
rect 515 2364 617 2366
rect 515 2363 516 2364
rect 510 2362 516 2363
rect 702 2363 703 2367
rect 707 2366 708 2367
rect 970 2367 976 2368
rect 707 2364 777 2366
rect 707 2363 708 2364
rect 702 2362 708 2363
rect 962 2363 968 2364
rect 110 2359 116 2360
rect 110 2355 111 2359
rect 115 2355 116 2359
rect 962 2359 963 2363
rect 967 2359 968 2363
rect 970 2363 971 2367
rect 975 2366 976 2367
rect 1122 2367 1128 2368
rect 975 2364 1081 2366
rect 975 2363 976 2364
rect 970 2362 976 2363
rect 1122 2363 1123 2367
rect 1127 2366 1128 2367
rect 1266 2367 1272 2368
rect 1127 2364 1225 2366
rect 1127 2363 1128 2364
rect 1122 2362 1128 2363
rect 1266 2363 1267 2367
rect 1271 2366 1272 2367
rect 1414 2367 1420 2368
rect 1271 2364 1369 2366
rect 1271 2363 1272 2364
rect 1266 2362 1272 2363
rect 1414 2363 1415 2367
rect 1419 2366 1420 2367
rect 1419 2364 1521 2366
rect 2046 2365 2052 2366
rect 1419 2363 1420 2364
rect 1414 2362 1420 2363
rect 2046 2361 2047 2365
rect 2051 2361 2052 2365
rect 2606 2364 2607 2368
rect 2611 2364 2612 2368
rect 2606 2363 2612 2364
rect 2814 2368 2820 2369
rect 2814 2364 2815 2368
rect 2819 2364 2820 2368
rect 2814 2363 2820 2364
rect 3006 2368 3012 2369
rect 3006 2364 3007 2368
rect 3011 2364 3012 2368
rect 3006 2363 3012 2364
rect 3190 2368 3196 2369
rect 3190 2364 3191 2368
rect 3195 2364 3196 2368
rect 3190 2363 3196 2364
rect 3358 2368 3364 2369
rect 3358 2364 3359 2368
rect 3363 2364 3364 2368
rect 3358 2363 3364 2364
rect 3518 2368 3524 2369
rect 3518 2364 3519 2368
rect 3523 2364 3524 2368
rect 3518 2363 3524 2364
rect 3678 2368 3684 2369
rect 3678 2364 3679 2368
rect 3683 2364 3684 2368
rect 3678 2363 3684 2364
rect 3838 2368 3844 2369
rect 3838 2364 3839 2368
rect 3843 2364 3844 2368
rect 3838 2363 3844 2364
rect 3942 2365 3948 2366
rect 2046 2360 2052 2361
rect 3942 2361 3943 2365
rect 3947 2361 3948 2365
rect 3942 2360 3948 2361
rect 962 2358 968 2359
rect 2006 2359 2012 2360
rect 110 2354 116 2355
rect 134 2356 140 2357
rect 134 2352 135 2356
rect 139 2352 140 2356
rect 134 2351 140 2352
rect 254 2356 260 2357
rect 254 2352 255 2356
rect 259 2352 260 2356
rect 254 2351 260 2352
rect 414 2356 420 2357
rect 414 2352 415 2356
rect 419 2352 420 2356
rect 414 2351 420 2352
rect 574 2356 580 2357
rect 574 2352 575 2356
rect 579 2352 580 2356
rect 574 2351 580 2352
rect 734 2356 740 2357
rect 734 2352 735 2356
rect 739 2352 740 2356
rect 734 2351 740 2352
rect 886 2356 892 2357
rect 886 2352 887 2356
rect 891 2352 892 2356
rect 886 2351 892 2352
rect 1038 2356 1044 2357
rect 1038 2352 1039 2356
rect 1043 2352 1044 2356
rect 1038 2351 1044 2352
rect 1182 2356 1188 2357
rect 1182 2352 1183 2356
rect 1187 2352 1188 2356
rect 1182 2351 1188 2352
rect 1326 2356 1332 2357
rect 1326 2352 1327 2356
rect 1331 2352 1332 2356
rect 1326 2351 1332 2352
rect 1478 2356 1484 2357
rect 1478 2352 1479 2356
rect 1483 2352 1484 2356
rect 2006 2355 2007 2359
rect 2011 2355 2012 2359
rect 2006 2354 2012 2355
rect 2682 2359 2688 2360
rect 2682 2355 2683 2359
rect 2687 2355 2688 2359
rect 2682 2354 2688 2355
rect 2890 2359 2896 2360
rect 2890 2355 2891 2359
rect 2895 2355 2896 2359
rect 2890 2354 2896 2355
rect 2942 2359 2948 2360
rect 2942 2355 2943 2359
rect 2947 2358 2948 2359
rect 3266 2359 3272 2360
rect 2947 2356 3049 2358
rect 2947 2355 2948 2356
rect 2942 2354 2948 2355
rect 3266 2355 3267 2359
rect 3271 2355 3272 2359
rect 3266 2354 3272 2355
rect 3434 2359 3440 2360
rect 3434 2355 3435 2359
rect 3439 2355 3440 2359
rect 3434 2354 3440 2355
rect 3594 2359 3600 2360
rect 3594 2355 3595 2359
rect 3599 2355 3600 2359
rect 3594 2354 3600 2355
rect 3754 2359 3760 2360
rect 3754 2355 3755 2359
rect 3759 2355 3760 2359
rect 3754 2354 3760 2355
rect 3906 2359 3912 2360
rect 3906 2355 3907 2359
rect 3911 2355 3912 2359
rect 3906 2354 3912 2355
rect 1478 2351 1484 2352
rect 2606 2349 2612 2350
rect 2046 2348 2052 2349
rect 2046 2344 2047 2348
rect 2051 2344 2052 2348
rect 2606 2345 2607 2349
rect 2611 2345 2612 2349
rect 2606 2344 2612 2345
rect 2814 2349 2820 2350
rect 2814 2345 2815 2349
rect 2819 2345 2820 2349
rect 2814 2344 2820 2345
rect 3006 2349 3012 2350
rect 3006 2345 3007 2349
rect 3011 2345 3012 2349
rect 3006 2344 3012 2345
rect 3190 2349 3196 2350
rect 3190 2345 3191 2349
rect 3195 2345 3196 2349
rect 3190 2344 3196 2345
rect 3358 2349 3364 2350
rect 3358 2345 3359 2349
rect 3363 2345 3364 2349
rect 3358 2344 3364 2345
rect 3518 2349 3524 2350
rect 3518 2345 3519 2349
rect 3523 2345 3524 2349
rect 3518 2344 3524 2345
rect 3678 2349 3684 2350
rect 3678 2345 3679 2349
rect 3683 2345 3684 2349
rect 3678 2344 3684 2345
rect 3838 2349 3844 2350
rect 3838 2345 3839 2349
rect 3843 2345 3844 2349
rect 3838 2344 3844 2345
rect 3942 2348 3948 2349
rect 3942 2344 3943 2348
rect 3947 2344 3948 2348
rect 2046 2343 2052 2344
rect 3942 2343 3948 2344
rect 187 2335 193 2336
rect 187 2331 188 2335
rect 192 2334 193 2335
rect 218 2335 224 2336
rect 218 2334 219 2335
rect 192 2332 219 2334
rect 192 2331 193 2332
rect 187 2330 193 2331
rect 218 2331 219 2332
rect 223 2331 224 2335
rect 218 2330 224 2331
rect 307 2335 313 2336
rect 307 2331 308 2335
rect 312 2334 313 2335
rect 358 2335 364 2336
rect 358 2334 359 2335
rect 312 2332 359 2334
rect 312 2331 313 2332
rect 307 2330 313 2331
rect 358 2331 359 2332
rect 363 2331 364 2335
rect 358 2330 364 2331
rect 467 2335 473 2336
rect 467 2331 468 2335
rect 472 2334 473 2335
rect 510 2335 516 2336
rect 510 2334 511 2335
rect 472 2332 511 2334
rect 472 2331 473 2332
rect 467 2330 473 2331
rect 510 2331 511 2332
rect 515 2331 516 2335
rect 510 2330 516 2331
rect 627 2335 633 2336
rect 627 2331 628 2335
rect 632 2334 633 2335
rect 702 2335 708 2336
rect 702 2334 703 2335
rect 632 2332 703 2334
rect 632 2331 633 2332
rect 627 2330 633 2331
rect 702 2331 703 2332
rect 707 2331 708 2335
rect 939 2335 945 2336
rect 702 2330 708 2331
rect 787 2331 793 2332
rect 787 2327 788 2331
rect 792 2330 793 2331
rect 810 2331 816 2332
rect 810 2330 811 2331
rect 792 2328 811 2330
rect 792 2327 793 2328
rect 787 2326 793 2327
rect 810 2327 811 2328
rect 815 2327 816 2331
rect 939 2331 940 2335
rect 944 2334 945 2335
rect 970 2335 976 2336
rect 970 2334 971 2335
rect 944 2332 971 2334
rect 944 2331 945 2332
rect 939 2330 945 2331
rect 970 2331 971 2332
rect 975 2331 976 2335
rect 970 2330 976 2331
rect 1091 2335 1097 2336
rect 1091 2331 1092 2335
rect 1096 2334 1097 2335
rect 1122 2335 1128 2336
rect 1122 2334 1123 2335
rect 1096 2332 1123 2334
rect 1096 2331 1097 2332
rect 1091 2330 1097 2331
rect 1122 2331 1123 2332
rect 1127 2331 1128 2335
rect 1122 2330 1128 2331
rect 1235 2335 1241 2336
rect 1235 2331 1236 2335
rect 1240 2334 1241 2335
rect 1266 2335 1272 2336
rect 1266 2334 1267 2335
rect 1240 2332 1267 2334
rect 1240 2331 1241 2332
rect 1235 2330 1241 2331
rect 1266 2331 1267 2332
rect 1271 2331 1272 2335
rect 1266 2330 1272 2331
rect 1379 2335 1385 2336
rect 1379 2331 1380 2335
rect 1384 2334 1385 2335
rect 1414 2335 1420 2336
rect 1414 2334 1415 2335
rect 1384 2332 1415 2334
rect 1384 2331 1385 2332
rect 1379 2330 1385 2331
rect 1414 2331 1415 2332
rect 1419 2331 1420 2335
rect 1414 2330 1420 2331
rect 1531 2331 1537 2332
rect 810 2326 816 2327
rect 1531 2327 1532 2331
rect 1536 2330 1537 2331
rect 1570 2331 1576 2332
rect 1570 2330 1571 2331
rect 1536 2328 1571 2330
rect 1536 2327 1537 2328
rect 1531 2326 1537 2327
rect 1570 2327 1571 2328
rect 1575 2327 1576 2331
rect 1570 2326 1576 2327
rect 187 2319 196 2320
rect 187 2315 188 2319
rect 195 2315 196 2319
rect 187 2314 196 2315
rect 210 2319 216 2320
rect 210 2315 211 2319
rect 215 2318 216 2319
rect 315 2319 321 2320
rect 315 2318 316 2319
rect 215 2316 316 2318
rect 215 2315 216 2316
rect 210 2314 216 2315
rect 315 2315 316 2316
rect 320 2315 321 2319
rect 315 2314 321 2315
rect 338 2319 344 2320
rect 338 2315 339 2319
rect 343 2318 344 2319
rect 475 2319 481 2320
rect 475 2318 476 2319
rect 343 2316 476 2318
rect 343 2315 344 2316
rect 338 2314 344 2315
rect 475 2315 476 2316
rect 480 2315 481 2319
rect 475 2314 481 2315
rect 498 2319 504 2320
rect 498 2315 499 2319
rect 503 2318 504 2319
rect 635 2319 641 2320
rect 635 2318 636 2319
rect 503 2316 636 2318
rect 503 2315 504 2316
rect 498 2314 504 2315
rect 635 2315 636 2316
rect 640 2315 641 2319
rect 635 2314 641 2315
rect 658 2319 664 2320
rect 658 2315 659 2319
rect 663 2318 664 2319
rect 795 2319 801 2320
rect 795 2318 796 2319
rect 663 2316 796 2318
rect 663 2315 664 2316
rect 658 2314 664 2315
rect 795 2315 796 2316
rect 800 2315 801 2319
rect 795 2314 801 2315
rect 947 2319 953 2320
rect 947 2315 948 2319
rect 952 2318 953 2319
rect 962 2319 968 2320
rect 962 2318 963 2319
rect 952 2316 963 2318
rect 952 2315 953 2316
rect 947 2314 953 2315
rect 962 2315 963 2316
rect 967 2315 968 2319
rect 962 2314 968 2315
rect 970 2319 976 2320
rect 970 2315 971 2319
rect 975 2318 976 2319
rect 1099 2319 1105 2320
rect 1099 2318 1100 2319
rect 975 2316 1100 2318
rect 975 2315 976 2316
rect 970 2314 976 2315
rect 1099 2315 1100 2316
rect 1104 2315 1105 2319
rect 1099 2314 1105 2315
rect 1251 2319 1260 2320
rect 1251 2315 1252 2319
rect 1259 2315 1260 2319
rect 1251 2314 1260 2315
rect 1274 2319 1280 2320
rect 1274 2315 1275 2319
rect 1279 2318 1280 2319
rect 1403 2319 1409 2320
rect 1403 2318 1404 2319
rect 1279 2316 1404 2318
rect 1279 2315 1280 2316
rect 1274 2314 1280 2315
rect 1403 2315 1404 2316
rect 1408 2315 1409 2319
rect 1403 2314 1409 2315
rect 1426 2319 1432 2320
rect 1426 2315 1427 2319
rect 1431 2318 1432 2319
rect 1555 2319 1561 2320
rect 1555 2318 1556 2319
rect 1431 2316 1556 2318
rect 1431 2315 1432 2316
rect 1426 2314 1432 2315
rect 1555 2315 1556 2316
rect 1560 2315 1561 2319
rect 1555 2314 1561 2315
rect 134 2296 140 2297
rect 110 2293 116 2294
rect 110 2289 111 2293
rect 115 2289 116 2293
rect 134 2292 135 2296
rect 139 2292 140 2296
rect 134 2291 140 2292
rect 262 2296 268 2297
rect 262 2292 263 2296
rect 267 2292 268 2296
rect 262 2291 268 2292
rect 422 2296 428 2297
rect 422 2292 423 2296
rect 427 2292 428 2296
rect 422 2291 428 2292
rect 582 2296 588 2297
rect 582 2292 583 2296
rect 587 2292 588 2296
rect 582 2291 588 2292
rect 742 2296 748 2297
rect 742 2292 743 2296
rect 747 2292 748 2296
rect 742 2291 748 2292
rect 894 2296 900 2297
rect 894 2292 895 2296
rect 899 2292 900 2296
rect 894 2291 900 2292
rect 1046 2296 1052 2297
rect 1046 2292 1047 2296
rect 1051 2292 1052 2296
rect 1046 2291 1052 2292
rect 1198 2296 1204 2297
rect 1198 2292 1199 2296
rect 1203 2292 1204 2296
rect 1198 2291 1204 2292
rect 1350 2296 1356 2297
rect 1350 2292 1351 2296
rect 1355 2292 1356 2296
rect 1350 2291 1356 2292
rect 1502 2296 1508 2297
rect 1502 2292 1503 2296
rect 1507 2292 1508 2296
rect 1502 2291 1508 2292
rect 2006 2293 2012 2294
rect 110 2288 116 2289
rect 2006 2289 2007 2293
rect 2011 2289 2012 2293
rect 2006 2288 2012 2289
rect 210 2287 216 2288
rect 210 2283 211 2287
rect 215 2283 216 2287
rect 210 2282 216 2283
rect 338 2287 344 2288
rect 338 2283 339 2287
rect 343 2283 344 2287
rect 338 2282 344 2283
rect 498 2287 504 2288
rect 498 2283 499 2287
rect 503 2283 504 2287
rect 498 2282 504 2283
rect 658 2287 664 2288
rect 658 2283 659 2287
rect 663 2283 664 2287
rect 658 2282 664 2283
rect 810 2287 816 2288
rect 810 2283 811 2287
rect 815 2283 816 2287
rect 810 2282 816 2283
rect 970 2287 976 2288
rect 970 2283 971 2287
rect 975 2283 976 2287
rect 970 2282 976 2283
rect 1014 2287 1020 2288
rect 1014 2283 1015 2287
rect 1019 2286 1020 2287
rect 1274 2287 1280 2288
rect 1019 2284 1089 2286
rect 1019 2283 1020 2284
rect 1014 2282 1020 2283
rect 1274 2283 1275 2287
rect 1279 2283 1280 2287
rect 1274 2282 1280 2283
rect 1426 2287 1432 2288
rect 1426 2283 1427 2287
rect 1431 2283 1432 2287
rect 1426 2282 1432 2283
rect 1570 2287 1576 2288
rect 1570 2283 1571 2287
rect 1575 2283 1576 2287
rect 1570 2282 1576 2283
rect 2046 2280 2052 2281
rect 3942 2280 3948 2281
rect 134 2277 140 2278
rect 110 2276 116 2277
rect 110 2272 111 2276
rect 115 2272 116 2276
rect 134 2273 135 2277
rect 139 2273 140 2277
rect 134 2272 140 2273
rect 262 2277 268 2278
rect 262 2273 263 2277
rect 267 2273 268 2277
rect 262 2272 268 2273
rect 422 2277 428 2278
rect 422 2273 423 2277
rect 427 2273 428 2277
rect 422 2272 428 2273
rect 582 2277 588 2278
rect 582 2273 583 2277
rect 587 2273 588 2277
rect 582 2272 588 2273
rect 742 2277 748 2278
rect 742 2273 743 2277
rect 747 2273 748 2277
rect 742 2272 748 2273
rect 894 2277 900 2278
rect 894 2273 895 2277
rect 899 2273 900 2277
rect 894 2272 900 2273
rect 1046 2277 1052 2278
rect 1046 2273 1047 2277
rect 1051 2273 1052 2277
rect 1046 2272 1052 2273
rect 1198 2277 1204 2278
rect 1198 2273 1199 2277
rect 1203 2273 1204 2277
rect 1198 2272 1204 2273
rect 1350 2277 1356 2278
rect 1350 2273 1351 2277
rect 1355 2273 1356 2277
rect 1350 2272 1356 2273
rect 1502 2277 1508 2278
rect 1502 2273 1503 2277
rect 1507 2273 1508 2277
rect 1502 2272 1508 2273
rect 2006 2276 2012 2277
rect 2006 2272 2007 2276
rect 2011 2272 2012 2276
rect 2046 2276 2047 2280
rect 2051 2276 2052 2280
rect 2046 2275 2052 2276
rect 2070 2279 2076 2280
rect 2070 2275 2071 2279
rect 2075 2275 2076 2279
rect 2070 2274 2076 2275
rect 2166 2279 2172 2280
rect 2166 2275 2167 2279
rect 2171 2275 2172 2279
rect 2166 2274 2172 2275
rect 2270 2279 2276 2280
rect 2270 2275 2271 2279
rect 2275 2275 2276 2279
rect 2270 2274 2276 2275
rect 2414 2279 2420 2280
rect 2414 2275 2415 2279
rect 2419 2275 2420 2279
rect 2414 2274 2420 2275
rect 2574 2279 2580 2280
rect 2574 2275 2575 2279
rect 2579 2275 2580 2279
rect 2574 2274 2580 2275
rect 2742 2279 2748 2280
rect 2742 2275 2743 2279
rect 2747 2275 2748 2279
rect 2742 2274 2748 2275
rect 2910 2279 2916 2280
rect 2910 2275 2911 2279
rect 2915 2275 2916 2279
rect 2910 2274 2916 2275
rect 3070 2279 3076 2280
rect 3070 2275 3071 2279
rect 3075 2275 3076 2279
rect 3070 2274 3076 2275
rect 3230 2279 3236 2280
rect 3230 2275 3231 2279
rect 3235 2275 3236 2279
rect 3230 2274 3236 2275
rect 3382 2279 3388 2280
rect 3382 2275 3383 2279
rect 3387 2275 3388 2279
rect 3382 2274 3388 2275
rect 3534 2279 3540 2280
rect 3534 2275 3535 2279
rect 3539 2275 3540 2279
rect 3534 2274 3540 2275
rect 3694 2279 3700 2280
rect 3694 2275 3695 2279
rect 3699 2275 3700 2279
rect 3942 2276 3943 2280
rect 3947 2276 3948 2280
rect 3942 2275 3948 2276
rect 3694 2274 3700 2275
rect 110 2271 116 2272
rect 2006 2271 2012 2272
rect 2250 2271 2256 2272
rect 2146 2267 2152 2268
rect 2046 2263 2052 2264
rect 2046 2259 2047 2263
rect 2051 2259 2052 2263
rect 2146 2263 2147 2267
rect 2151 2263 2152 2267
rect 2146 2262 2152 2263
rect 2242 2267 2248 2268
rect 2242 2263 2243 2267
rect 2247 2263 2248 2267
rect 2250 2267 2251 2271
rect 2255 2270 2256 2271
rect 2358 2271 2364 2272
rect 2255 2268 2313 2270
rect 2255 2267 2256 2268
rect 2250 2266 2256 2267
rect 2358 2267 2359 2271
rect 2363 2270 2364 2271
rect 2534 2271 2540 2272
rect 2363 2268 2457 2270
rect 2363 2267 2364 2268
rect 2358 2266 2364 2267
rect 2534 2267 2535 2271
rect 2539 2270 2540 2271
rect 2658 2271 2664 2272
rect 2539 2268 2617 2270
rect 2539 2267 2540 2268
rect 2534 2266 2540 2267
rect 2658 2267 2659 2271
rect 2663 2270 2664 2271
rect 2870 2271 2876 2272
rect 2663 2268 2785 2270
rect 2663 2267 2664 2268
rect 2658 2266 2664 2267
rect 2870 2267 2871 2271
rect 2875 2270 2876 2271
rect 3618 2271 3624 2272
rect 2875 2268 2953 2270
rect 2875 2267 2876 2268
rect 2870 2266 2876 2267
rect 3146 2267 3152 2268
rect 2242 2262 2248 2263
rect 3146 2263 3147 2267
rect 3151 2263 3152 2267
rect 3146 2262 3152 2263
rect 3306 2267 3312 2268
rect 3306 2263 3307 2267
rect 3311 2263 3312 2267
rect 3306 2262 3312 2263
rect 3458 2267 3464 2268
rect 3458 2263 3459 2267
rect 3463 2263 3464 2267
rect 3458 2262 3464 2263
rect 3610 2267 3616 2268
rect 3610 2263 3611 2267
rect 3615 2263 3616 2267
rect 3618 2267 3619 2271
rect 3623 2270 3624 2271
rect 3623 2268 3737 2270
rect 3623 2267 3624 2268
rect 3618 2266 3624 2267
rect 3610 2262 3616 2263
rect 3942 2263 3948 2264
rect 2046 2258 2052 2259
rect 2070 2260 2076 2261
rect 2070 2256 2071 2260
rect 2075 2256 2076 2260
rect 2070 2255 2076 2256
rect 2166 2260 2172 2261
rect 2166 2256 2167 2260
rect 2171 2256 2172 2260
rect 2166 2255 2172 2256
rect 2270 2260 2276 2261
rect 2270 2256 2271 2260
rect 2275 2256 2276 2260
rect 2270 2255 2276 2256
rect 2414 2260 2420 2261
rect 2414 2256 2415 2260
rect 2419 2256 2420 2260
rect 2414 2255 2420 2256
rect 2574 2260 2580 2261
rect 2574 2256 2575 2260
rect 2579 2256 2580 2260
rect 2574 2255 2580 2256
rect 2742 2260 2748 2261
rect 2742 2256 2743 2260
rect 2747 2256 2748 2260
rect 2742 2255 2748 2256
rect 2910 2260 2916 2261
rect 2910 2256 2911 2260
rect 2915 2256 2916 2260
rect 2910 2255 2916 2256
rect 3070 2260 3076 2261
rect 3070 2256 3071 2260
rect 3075 2256 3076 2260
rect 3070 2255 3076 2256
rect 3230 2260 3236 2261
rect 3230 2256 3231 2260
rect 3235 2256 3236 2260
rect 3230 2255 3236 2256
rect 3382 2260 3388 2261
rect 3382 2256 3383 2260
rect 3387 2256 3388 2260
rect 3382 2255 3388 2256
rect 3534 2260 3540 2261
rect 3534 2256 3535 2260
rect 3539 2256 3540 2260
rect 3534 2255 3540 2256
rect 3694 2260 3700 2261
rect 3694 2256 3695 2260
rect 3699 2256 3700 2260
rect 3942 2259 3943 2263
rect 3947 2259 3948 2263
rect 3942 2258 3948 2259
rect 3694 2255 3700 2256
rect 2250 2247 2256 2248
rect 2250 2246 2251 2247
rect 2140 2244 2251 2246
rect 2123 2239 2129 2240
rect 2123 2235 2124 2239
rect 2128 2238 2129 2239
rect 2140 2238 2142 2244
rect 2250 2243 2251 2244
rect 2255 2243 2256 2247
rect 3450 2247 3456 2248
rect 3450 2246 3451 2247
rect 2250 2242 2256 2243
rect 3140 2244 3451 2246
rect 2128 2236 2142 2238
rect 2146 2239 2152 2240
rect 2128 2235 2129 2236
rect 2123 2234 2129 2235
rect 2146 2235 2147 2239
rect 2151 2238 2152 2239
rect 2219 2239 2225 2240
rect 2219 2238 2220 2239
rect 2151 2236 2220 2238
rect 2151 2235 2152 2236
rect 2146 2234 2152 2235
rect 2219 2235 2220 2236
rect 2224 2235 2225 2239
rect 2219 2234 2225 2235
rect 2323 2239 2329 2240
rect 2323 2235 2324 2239
rect 2328 2238 2329 2239
rect 2358 2239 2364 2240
rect 2358 2238 2359 2239
rect 2328 2236 2359 2238
rect 2328 2235 2329 2236
rect 2323 2234 2329 2235
rect 2358 2235 2359 2236
rect 2363 2235 2364 2239
rect 2358 2234 2364 2235
rect 2467 2239 2473 2240
rect 2467 2235 2468 2239
rect 2472 2238 2473 2239
rect 2534 2239 2540 2240
rect 2534 2238 2535 2239
rect 2472 2236 2535 2238
rect 2472 2235 2473 2236
rect 2467 2234 2473 2235
rect 2534 2235 2535 2236
rect 2539 2235 2540 2239
rect 2534 2234 2540 2235
rect 2627 2239 2633 2240
rect 2627 2235 2628 2239
rect 2632 2238 2633 2239
rect 2658 2239 2664 2240
rect 2658 2238 2659 2239
rect 2632 2236 2659 2238
rect 2632 2235 2633 2236
rect 2627 2234 2633 2235
rect 2658 2235 2659 2236
rect 2663 2235 2664 2239
rect 2890 2239 2896 2240
rect 2658 2234 2664 2235
rect 2698 2235 2704 2236
rect 2698 2231 2699 2235
rect 2703 2234 2704 2235
rect 2795 2235 2801 2236
rect 2795 2234 2796 2235
rect 2703 2232 2796 2234
rect 2703 2231 2704 2232
rect 2698 2230 2704 2231
rect 2795 2231 2796 2232
rect 2800 2231 2801 2235
rect 2890 2235 2891 2239
rect 2895 2238 2896 2239
rect 2963 2239 2969 2240
rect 2963 2238 2964 2239
rect 2895 2236 2964 2238
rect 2895 2235 2896 2236
rect 2890 2234 2896 2235
rect 2963 2235 2964 2236
rect 2968 2235 2969 2239
rect 2963 2234 2969 2235
rect 3123 2239 3129 2240
rect 3123 2235 3124 2239
rect 3128 2238 3129 2239
rect 3140 2238 3142 2244
rect 3450 2243 3451 2244
rect 3455 2243 3456 2247
rect 3450 2242 3456 2243
rect 3128 2236 3142 2238
rect 3146 2239 3152 2240
rect 3128 2235 3129 2236
rect 3123 2234 3129 2235
rect 3146 2235 3147 2239
rect 3151 2238 3152 2239
rect 3283 2239 3289 2240
rect 3283 2238 3284 2239
rect 3151 2236 3284 2238
rect 3151 2235 3152 2236
rect 3146 2234 3152 2235
rect 3283 2235 3284 2236
rect 3288 2235 3289 2239
rect 3283 2234 3289 2235
rect 3306 2239 3312 2240
rect 3306 2235 3307 2239
rect 3311 2238 3312 2239
rect 3435 2239 3441 2240
rect 3435 2238 3436 2239
rect 3311 2236 3436 2238
rect 3311 2235 3312 2236
rect 3306 2234 3312 2235
rect 3435 2235 3436 2236
rect 3440 2235 3441 2239
rect 3435 2234 3441 2235
rect 3458 2239 3464 2240
rect 3458 2235 3459 2239
rect 3463 2238 3464 2239
rect 3587 2239 3593 2240
rect 3587 2238 3588 2239
rect 3463 2236 3588 2238
rect 3463 2235 3464 2236
rect 3458 2234 3464 2235
rect 3587 2235 3588 2236
rect 3592 2235 3593 2239
rect 3587 2234 3593 2235
rect 3610 2239 3616 2240
rect 3610 2235 3611 2239
rect 3615 2238 3616 2239
rect 3747 2239 3753 2240
rect 3747 2238 3748 2239
rect 3615 2236 3748 2238
rect 3615 2235 3616 2236
rect 3610 2234 3616 2235
rect 3747 2235 3748 2236
rect 3752 2235 3753 2239
rect 3747 2234 3753 2235
rect 2795 2230 2801 2231
rect 2123 2223 2129 2224
rect 110 2220 116 2221
rect 2006 2220 2012 2221
rect 110 2216 111 2220
rect 115 2216 116 2220
rect 110 2215 116 2216
rect 222 2219 228 2220
rect 222 2215 223 2219
rect 227 2215 228 2219
rect 222 2214 228 2215
rect 350 2219 356 2220
rect 350 2215 351 2219
rect 355 2215 356 2219
rect 350 2214 356 2215
rect 494 2219 500 2220
rect 494 2215 495 2219
rect 499 2215 500 2219
rect 494 2214 500 2215
rect 646 2219 652 2220
rect 646 2215 647 2219
rect 651 2215 652 2219
rect 646 2214 652 2215
rect 798 2219 804 2220
rect 798 2215 799 2219
rect 803 2215 804 2219
rect 798 2214 804 2215
rect 958 2219 964 2220
rect 958 2215 959 2219
rect 963 2215 964 2219
rect 958 2214 964 2215
rect 1118 2219 1124 2220
rect 1118 2215 1119 2219
rect 1123 2215 1124 2219
rect 1118 2214 1124 2215
rect 1278 2219 1284 2220
rect 1278 2215 1279 2219
rect 1283 2215 1284 2219
rect 1278 2214 1284 2215
rect 1438 2219 1444 2220
rect 1438 2215 1439 2219
rect 1443 2215 1444 2219
rect 1438 2214 1444 2215
rect 1598 2219 1604 2220
rect 1598 2215 1599 2219
rect 1603 2215 1604 2219
rect 2006 2216 2007 2220
rect 2011 2216 2012 2220
rect 2123 2219 2124 2223
rect 2128 2222 2129 2223
rect 2154 2223 2160 2224
rect 2154 2222 2155 2223
rect 2128 2220 2155 2222
rect 2128 2219 2129 2220
rect 2123 2218 2129 2219
rect 2154 2219 2155 2220
rect 2159 2219 2160 2223
rect 2154 2218 2160 2219
rect 2227 2223 2233 2224
rect 2227 2219 2228 2223
rect 2232 2222 2233 2223
rect 2242 2223 2248 2224
rect 2242 2222 2243 2223
rect 2232 2220 2243 2222
rect 2232 2219 2233 2220
rect 2227 2218 2233 2219
rect 2242 2219 2243 2220
rect 2247 2219 2248 2223
rect 2242 2218 2248 2219
rect 2354 2223 2360 2224
rect 2354 2219 2355 2223
rect 2359 2222 2360 2223
rect 2371 2223 2377 2224
rect 2371 2222 2372 2223
rect 2359 2220 2372 2222
rect 2359 2219 2360 2220
rect 2354 2218 2360 2219
rect 2371 2219 2372 2220
rect 2376 2219 2377 2223
rect 2371 2218 2377 2219
rect 2394 2223 2400 2224
rect 2394 2219 2395 2223
rect 2399 2222 2400 2223
rect 2523 2223 2529 2224
rect 2523 2222 2524 2223
rect 2399 2220 2524 2222
rect 2399 2219 2400 2220
rect 2394 2218 2400 2219
rect 2523 2219 2524 2220
rect 2528 2219 2529 2223
rect 2523 2218 2529 2219
rect 2546 2223 2552 2224
rect 2546 2219 2547 2223
rect 2551 2222 2552 2223
rect 2675 2223 2681 2224
rect 2675 2222 2676 2223
rect 2551 2220 2676 2222
rect 2551 2219 2552 2220
rect 2546 2218 2552 2219
rect 2675 2219 2676 2220
rect 2680 2219 2681 2223
rect 2675 2218 2681 2219
rect 2835 2223 2841 2224
rect 2835 2219 2836 2223
rect 2840 2222 2841 2223
rect 2870 2223 2876 2224
rect 2870 2222 2871 2223
rect 2840 2220 2871 2222
rect 2840 2219 2841 2220
rect 2835 2218 2841 2219
rect 2870 2219 2871 2220
rect 2875 2219 2876 2223
rect 2870 2218 2876 2219
rect 2987 2223 2996 2224
rect 2987 2219 2988 2223
rect 2995 2219 2996 2223
rect 2987 2218 2996 2219
rect 3010 2223 3016 2224
rect 3010 2219 3011 2223
rect 3015 2222 3016 2223
rect 3131 2223 3137 2224
rect 3131 2222 3132 2223
rect 3015 2220 3132 2222
rect 3015 2219 3016 2220
rect 3010 2218 3016 2219
rect 3131 2219 3132 2220
rect 3136 2219 3137 2223
rect 3131 2218 3137 2219
rect 3154 2223 3160 2224
rect 3154 2219 3155 2223
rect 3159 2222 3160 2223
rect 3275 2223 3281 2224
rect 3275 2222 3276 2223
rect 3159 2220 3276 2222
rect 3159 2219 3160 2220
rect 3154 2218 3160 2219
rect 3275 2219 3276 2220
rect 3280 2219 3281 2223
rect 3275 2218 3281 2219
rect 3298 2223 3304 2224
rect 3298 2219 3299 2223
rect 3303 2222 3304 2223
rect 3419 2223 3425 2224
rect 3419 2222 3420 2223
rect 3303 2220 3420 2222
rect 3303 2219 3304 2220
rect 3298 2218 3304 2219
rect 3419 2219 3420 2220
rect 3424 2219 3425 2223
rect 3419 2218 3425 2219
rect 3442 2223 3448 2224
rect 3442 2219 3443 2223
rect 3447 2222 3448 2223
rect 3571 2223 3577 2224
rect 3571 2222 3572 2223
rect 3447 2220 3572 2222
rect 3447 2219 3448 2220
rect 3442 2218 3448 2219
rect 3571 2219 3572 2220
rect 3576 2219 3577 2223
rect 3571 2218 3577 2219
rect 2006 2215 2012 2216
rect 1598 2214 1604 2215
rect 190 2211 196 2212
rect 190 2207 191 2211
rect 195 2210 196 2211
rect 306 2211 312 2212
rect 195 2208 265 2210
rect 195 2207 196 2208
rect 190 2206 196 2207
rect 306 2207 307 2211
rect 311 2210 312 2211
rect 439 2211 445 2212
rect 311 2208 393 2210
rect 311 2207 312 2208
rect 306 2206 312 2207
rect 439 2207 440 2211
rect 444 2210 445 2211
rect 583 2211 589 2212
rect 444 2208 537 2210
rect 444 2207 445 2208
rect 439 2206 445 2207
rect 583 2207 584 2211
rect 588 2210 589 2211
rect 759 2211 765 2212
rect 588 2208 689 2210
rect 588 2207 589 2208
rect 583 2206 589 2207
rect 759 2207 760 2211
rect 764 2210 765 2211
rect 1254 2211 1260 2212
rect 764 2208 841 2210
rect 764 2207 765 2208
rect 759 2206 765 2207
rect 1034 2207 1040 2208
rect 110 2203 116 2204
rect 110 2199 111 2203
rect 115 2199 116 2203
rect 1034 2203 1035 2207
rect 1039 2203 1040 2207
rect 1034 2202 1040 2203
rect 1194 2207 1200 2208
rect 1194 2203 1195 2207
rect 1199 2203 1200 2207
rect 1254 2207 1255 2211
rect 1259 2210 1260 2211
rect 1399 2211 1405 2212
rect 1259 2208 1321 2210
rect 1259 2207 1260 2208
rect 1254 2206 1260 2207
rect 1399 2207 1400 2211
rect 1404 2210 1405 2211
rect 1551 2211 1557 2212
rect 1404 2208 1481 2210
rect 1404 2207 1405 2208
rect 1399 2206 1405 2207
rect 1551 2207 1552 2211
rect 1556 2210 1557 2211
rect 1556 2208 1641 2210
rect 1556 2207 1557 2208
rect 1551 2206 1557 2207
rect 1194 2202 1200 2203
rect 2006 2203 2012 2204
rect 110 2198 116 2199
rect 222 2200 228 2201
rect 222 2196 223 2200
rect 227 2196 228 2200
rect 222 2195 228 2196
rect 350 2200 356 2201
rect 350 2196 351 2200
rect 355 2196 356 2200
rect 350 2195 356 2196
rect 494 2200 500 2201
rect 494 2196 495 2200
rect 499 2196 500 2200
rect 494 2195 500 2196
rect 646 2200 652 2201
rect 646 2196 647 2200
rect 651 2196 652 2200
rect 646 2195 652 2196
rect 798 2200 804 2201
rect 798 2196 799 2200
rect 803 2196 804 2200
rect 798 2195 804 2196
rect 958 2200 964 2201
rect 958 2196 959 2200
rect 963 2196 964 2200
rect 958 2195 964 2196
rect 1118 2200 1124 2201
rect 1118 2196 1119 2200
rect 1123 2196 1124 2200
rect 1118 2195 1124 2196
rect 1278 2200 1284 2201
rect 1278 2196 1279 2200
rect 1283 2196 1284 2200
rect 1278 2195 1284 2196
rect 1438 2200 1444 2201
rect 1438 2196 1439 2200
rect 1443 2196 1444 2200
rect 1438 2195 1444 2196
rect 1598 2200 1604 2201
rect 1598 2196 1599 2200
rect 1603 2196 1604 2200
rect 2006 2199 2007 2203
rect 2011 2199 2012 2203
rect 2006 2198 2012 2199
rect 2070 2200 2076 2201
rect 1598 2195 1604 2196
rect 2046 2197 2052 2198
rect 2046 2193 2047 2197
rect 2051 2193 2052 2197
rect 2070 2196 2071 2200
rect 2075 2196 2076 2200
rect 2070 2195 2076 2196
rect 2174 2200 2180 2201
rect 2174 2196 2175 2200
rect 2179 2196 2180 2200
rect 2174 2195 2180 2196
rect 2318 2200 2324 2201
rect 2318 2196 2319 2200
rect 2323 2196 2324 2200
rect 2318 2195 2324 2196
rect 2470 2200 2476 2201
rect 2470 2196 2471 2200
rect 2475 2196 2476 2200
rect 2470 2195 2476 2196
rect 2622 2200 2628 2201
rect 2622 2196 2623 2200
rect 2627 2196 2628 2200
rect 2622 2195 2628 2196
rect 2782 2200 2788 2201
rect 2782 2196 2783 2200
rect 2787 2196 2788 2200
rect 2782 2195 2788 2196
rect 2934 2200 2940 2201
rect 2934 2196 2935 2200
rect 2939 2196 2940 2200
rect 2934 2195 2940 2196
rect 3078 2200 3084 2201
rect 3078 2196 3079 2200
rect 3083 2196 3084 2200
rect 3078 2195 3084 2196
rect 3222 2200 3228 2201
rect 3222 2196 3223 2200
rect 3227 2196 3228 2200
rect 3222 2195 3228 2196
rect 3366 2200 3372 2201
rect 3366 2196 3367 2200
rect 3371 2196 3372 2200
rect 3366 2195 3372 2196
rect 3518 2200 3524 2201
rect 3518 2196 3519 2200
rect 3523 2196 3524 2200
rect 3518 2195 3524 2196
rect 3942 2197 3948 2198
rect 2046 2192 2052 2193
rect 3942 2193 3943 2197
rect 3947 2193 3948 2197
rect 3942 2192 3948 2193
rect 1975 2191 1981 2192
rect 1975 2187 1976 2191
rect 1980 2190 1981 2191
rect 2154 2191 2160 2192
rect 1980 2188 2113 2190
rect 1980 2187 1981 2188
rect 1975 2186 1981 2187
rect 2154 2187 2155 2191
rect 2159 2190 2160 2191
rect 2394 2191 2400 2192
rect 2159 2188 2217 2190
rect 2159 2187 2160 2188
rect 2154 2186 2160 2187
rect 2394 2187 2395 2191
rect 2399 2187 2400 2191
rect 2394 2186 2400 2187
rect 2546 2191 2552 2192
rect 2546 2187 2547 2191
rect 2551 2187 2552 2191
rect 2546 2186 2552 2187
rect 2698 2191 2704 2192
rect 2698 2187 2699 2191
rect 2703 2187 2704 2191
rect 2698 2186 2704 2187
rect 2850 2191 2856 2192
rect 2850 2187 2851 2191
rect 2855 2187 2856 2191
rect 2850 2186 2856 2187
rect 3010 2191 3016 2192
rect 3010 2187 3011 2191
rect 3015 2187 3016 2191
rect 3010 2186 3016 2187
rect 3154 2191 3160 2192
rect 3154 2187 3155 2191
rect 3159 2187 3160 2191
rect 3154 2186 3160 2187
rect 3298 2191 3304 2192
rect 3298 2187 3299 2191
rect 3303 2187 3304 2191
rect 3298 2186 3304 2187
rect 3442 2191 3448 2192
rect 3442 2187 3443 2191
rect 3447 2187 3448 2191
rect 3442 2186 3448 2187
rect 3450 2191 3456 2192
rect 3450 2187 3451 2191
rect 3455 2190 3456 2191
rect 3455 2188 3561 2190
rect 3455 2187 3456 2188
rect 3450 2186 3456 2187
rect 2070 2181 2076 2182
rect 2046 2180 2052 2181
rect 275 2179 281 2180
rect 275 2175 276 2179
rect 280 2178 281 2179
rect 306 2179 312 2180
rect 306 2178 307 2179
rect 280 2176 307 2178
rect 280 2175 281 2176
rect 275 2174 281 2175
rect 306 2175 307 2176
rect 311 2175 312 2179
rect 306 2174 312 2175
rect 403 2179 409 2180
rect 403 2175 404 2179
rect 408 2178 409 2179
rect 439 2179 445 2180
rect 439 2178 440 2179
rect 408 2176 440 2178
rect 408 2175 409 2176
rect 403 2174 409 2175
rect 439 2175 440 2176
rect 444 2175 445 2179
rect 439 2174 445 2175
rect 547 2179 553 2180
rect 547 2175 548 2179
rect 552 2178 553 2179
rect 583 2179 589 2180
rect 583 2178 584 2179
rect 552 2176 584 2178
rect 552 2175 553 2176
rect 547 2174 553 2175
rect 583 2175 584 2176
rect 588 2175 589 2179
rect 583 2174 589 2175
rect 699 2179 705 2180
rect 699 2175 700 2179
rect 704 2178 705 2179
rect 759 2179 765 2180
rect 759 2178 760 2179
rect 704 2176 760 2178
rect 704 2175 705 2176
rect 699 2174 705 2175
rect 759 2175 760 2176
rect 764 2175 765 2179
rect 1011 2179 1020 2180
rect 759 2174 765 2175
rect 783 2175 789 2176
rect 783 2171 784 2175
rect 788 2174 789 2175
rect 851 2175 857 2176
rect 851 2174 852 2175
rect 788 2172 852 2174
rect 788 2171 789 2172
rect 783 2170 789 2171
rect 851 2171 852 2172
rect 856 2171 857 2175
rect 1011 2175 1012 2179
rect 1019 2175 1020 2179
rect 1011 2174 1020 2175
rect 1034 2179 1040 2180
rect 1034 2175 1035 2179
rect 1039 2178 1040 2179
rect 1171 2179 1177 2180
rect 1171 2178 1172 2179
rect 1039 2176 1172 2178
rect 1039 2175 1040 2176
rect 1034 2174 1040 2175
rect 1171 2175 1172 2176
rect 1176 2175 1177 2179
rect 1171 2174 1177 2175
rect 1331 2179 1337 2180
rect 1331 2175 1332 2179
rect 1336 2178 1337 2179
rect 1399 2179 1405 2180
rect 1399 2178 1400 2179
rect 1336 2176 1400 2178
rect 1336 2175 1337 2176
rect 1331 2174 1337 2175
rect 1399 2175 1400 2176
rect 1404 2175 1405 2179
rect 1399 2174 1405 2175
rect 1491 2179 1497 2180
rect 1491 2175 1492 2179
rect 1496 2178 1497 2179
rect 1551 2179 1557 2180
rect 1551 2178 1552 2179
rect 1496 2176 1552 2178
rect 1496 2175 1497 2176
rect 1491 2174 1497 2175
rect 1551 2175 1552 2176
rect 1556 2175 1557 2179
rect 2046 2176 2047 2180
rect 2051 2176 2052 2180
rect 2070 2177 2071 2181
rect 2075 2177 2076 2181
rect 2070 2176 2076 2177
rect 2174 2181 2180 2182
rect 2174 2177 2175 2181
rect 2179 2177 2180 2181
rect 2174 2176 2180 2177
rect 2318 2181 2324 2182
rect 2318 2177 2319 2181
rect 2323 2177 2324 2181
rect 2318 2176 2324 2177
rect 2470 2181 2476 2182
rect 2470 2177 2471 2181
rect 2475 2177 2476 2181
rect 2470 2176 2476 2177
rect 2622 2181 2628 2182
rect 2622 2177 2623 2181
rect 2627 2177 2628 2181
rect 2622 2176 2628 2177
rect 2782 2181 2788 2182
rect 2782 2177 2783 2181
rect 2787 2177 2788 2181
rect 2782 2176 2788 2177
rect 2934 2181 2940 2182
rect 2934 2177 2935 2181
rect 2939 2177 2940 2181
rect 2934 2176 2940 2177
rect 3078 2181 3084 2182
rect 3078 2177 3079 2181
rect 3083 2177 3084 2181
rect 3078 2176 3084 2177
rect 3222 2181 3228 2182
rect 3222 2177 3223 2181
rect 3227 2177 3228 2181
rect 3222 2176 3228 2177
rect 3366 2181 3372 2182
rect 3366 2177 3367 2181
rect 3371 2177 3372 2181
rect 3366 2176 3372 2177
rect 3518 2181 3524 2182
rect 3518 2177 3519 2181
rect 3523 2177 3524 2181
rect 3518 2176 3524 2177
rect 3942 2180 3948 2181
rect 3942 2176 3943 2180
rect 3947 2176 3948 2180
rect 1551 2174 1557 2175
rect 1578 2175 1584 2176
rect 851 2170 857 2171
rect 1578 2171 1579 2175
rect 1583 2174 1584 2175
rect 1651 2175 1657 2176
rect 2046 2175 2052 2176
rect 3942 2175 3948 2176
rect 1651 2174 1652 2175
rect 1583 2172 1652 2174
rect 1583 2171 1584 2172
rect 1578 2170 1584 2171
rect 1651 2171 1652 2172
rect 1656 2171 1657 2175
rect 1651 2170 1657 2171
rect 546 2163 552 2164
rect 523 2161 529 2162
rect 523 2157 524 2161
rect 528 2157 529 2161
rect 546 2159 547 2163
rect 551 2162 552 2163
rect 619 2163 625 2164
rect 619 2162 620 2163
rect 551 2160 620 2162
rect 551 2159 552 2160
rect 546 2158 552 2159
rect 619 2159 620 2160
rect 624 2159 625 2163
rect 619 2158 625 2159
rect 670 2163 676 2164
rect 670 2159 671 2163
rect 675 2162 676 2163
rect 731 2163 737 2164
rect 731 2162 732 2163
rect 675 2160 732 2162
rect 675 2159 676 2160
rect 670 2158 676 2159
rect 731 2159 732 2160
rect 736 2159 737 2163
rect 731 2158 737 2159
rect 859 2163 865 2164
rect 859 2159 860 2163
rect 864 2162 865 2163
rect 890 2163 896 2164
rect 890 2162 891 2163
rect 864 2160 891 2162
rect 864 2159 865 2160
rect 859 2158 865 2159
rect 890 2159 891 2160
rect 895 2159 896 2163
rect 890 2158 896 2159
rect 995 2163 1001 2164
rect 995 2159 996 2163
rect 1000 2162 1001 2163
rect 1071 2163 1077 2164
rect 1071 2162 1072 2163
rect 1000 2160 1072 2162
rect 1000 2159 1001 2160
rect 995 2158 1001 2159
rect 1071 2159 1072 2160
rect 1076 2159 1077 2163
rect 1071 2158 1077 2159
rect 1131 2163 1137 2164
rect 1131 2159 1132 2163
rect 1136 2162 1137 2163
rect 1194 2163 1200 2164
rect 1194 2162 1195 2163
rect 1136 2160 1195 2162
rect 1136 2159 1137 2160
rect 1131 2158 1137 2159
rect 1194 2159 1195 2160
rect 1199 2159 1200 2163
rect 1194 2158 1200 2159
rect 1215 2163 1221 2164
rect 1215 2159 1216 2163
rect 1220 2162 1221 2163
rect 1275 2163 1281 2164
rect 1275 2162 1276 2163
rect 1220 2160 1276 2162
rect 1220 2159 1221 2160
rect 1215 2158 1221 2159
rect 1275 2159 1276 2160
rect 1280 2159 1281 2163
rect 1479 2163 1485 2164
rect 1275 2158 1281 2159
rect 1419 2161 1425 2162
rect 523 2156 529 2157
rect 1419 2157 1420 2161
rect 1424 2157 1425 2161
rect 1479 2159 1480 2163
rect 1484 2162 1485 2163
rect 1555 2163 1561 2164
rect 1555 2162 1556 2163
rect 1484 2160 1556 2162
rect 1484 2159 1485 2160
rect 1479 2158 1485 2159
rect 1555 2159 1556 2160
rect 1560 2159 1561 2163
rect 1555 2158 1561 2159
rect 1691 2163 1697 2164
rect 1691 2159 1692 2163
rect 1696 2162 1697 2163
rect 1730 2163 1736 2164
rect 1730 2162 1731 2163
rect 1696 2160 1731 2162
rect 1696 2159 1697 2160
rect 1691 2158 1697 2159
rect 1730 2159 1731 2160
rect 1735 2159 1736 2163
rect 1730 2158 1736 2159
rect 1835 2163 1841 2164
rect 1835 2159 1836 2163
rect 1840 2162 1841 2163
rect 1866 2163 1872 2164
rect 1866 2162 1867 2163
rect 1840 2160 1867 2162
rect 1840 2159 1841 2160
rect 1835 2158 1841 2159
rect 1866 2159 1867 2160
rect 1871 2159 1872 2163
rect 1866 2158 1872 2159
rect 1955 2163 1961 2164
rect 1955 2159 1956 2163
rect 1960 2162 1961 2163
rect 1975 2163 1981 2164
rect 1975 2162 1976 2163
rect 1960 2160 1976 2162
rect 1960 2159 1961 2160
rect 1955 2158 1961 2159
rect 1975 2159 1976 2160
rect 1980 2159 1981 2163
rect 1975 2158 1981 2159
rect 1419 2156 1425 2157
rect 524 2154 526 2156
rect 791 2155 797 2156
rect 791 2154 792 2155
rect 524 2152 792 2154
rect 791 2151 792 2152
rect 796 2151 797 2155
rect 1420 2154 1422 2156
rect 1586 2155 1592 2156
rect 1586 2154 1587 2155
rect 1420 2152 1587 2154
rect 791 2150 797 2151
rect 1586 2151 1587 2152
rect 1591 2151 1592 2155
rect 1586 2150 1592 2151
rect 470 2140 476 2141
rect 110 2137 116 2138
rect 110 2133 111 2137
rect 115 2133 116 2137
rect 470 2136 471 2140
rect 475 2136 476 2140
rect 470 2135 476 2136
rect 566 2140 572 2141
rect 566 2136 567 2140
rect 571 2136 572 2140
rect 566 2135 572 2136
rect 678 2140 684 2141
rect 678 2136 679 2140
rect 683 2136 684 2140
rect 678 2135 684 2136
rect 806 2140 812 2141
rect 806 2136 807 2140
rect 811 2136 812 2140
rect 806 2135 812 2136
rect 942 2140 948 2141
rect 942 2136 943 2140
rect 947 2136 948 2140
rect 942 2135 948 2136
rect 1078 2140 1084 2141
rect 1078 2136 1079 2140
rect 1083 2136 1084 2140
rect 1078 2135 1084 2136
rect 1222 2140 1228 2141
rect 1222 2136 1223 2140
rect 1227 2136 1228 2140
rect 1222 2135 1228 2136
rect 1366 2140 1372 2141
rect 1366 2136 1367 2140
rect 1371 2136 1372 2140
rect 1366 2135 1372 2136
rect 1502 2140 1508 2141
rect 1502 2136 1503 2140
rect 1507 2136 1508 2140
rect 1502 2135 1508 2136
rect 1638 2140 1644 2141
rect 1638 2136 1639 2140
rect 1643 2136 1644 2140
rect 1638 2135 1644 2136
rect 1782 2140 1788 2141
rect 1782 2136 1783 2140
rect 1787 2136 1788 2140
rect 1782 2135 1788 2136
rect 1902 2140 1908 2141
rect 1902 2136 1903 2140
rect 1907 2136 1908 2140
rect 1902 2135 1908 2136
rect 2006 2137 2012 2138
rect 110 2132 116 2133
rect 2006 2133 2007 2137
rect 2011 2133 2012 2137
rect 2006 2132 2012 2133
rect 546 2131 552 2132
rect 546 2127 547 2131
rect 551 2127 552 2131
rect 670 2131 676 2132
rect 670 2130 671 2131
rect 645 2128 671 2130
rect 546 2126 552 2127
rect 670 2127 671 2128
rect 675 2127 676 2131
rect 783 2131 789 2132
rect 783 2130 784 2131
rect 757 2128 784 2130
rect 670 2126 676 2127
rect 783 2127 784 2128
rect 788 2127 789 2131
rect 783 2126 789 2127
rect 791 2131 797 2132
rect 791 2127 792 2131
rect 796 2130 797 2131
rect 890 2131 896 2132
rect 796 2128 849 2130
rect 796 2127 797 2128
rect 791 2126 797 2127
rect 890 2127 891 2131
rect 895 2130 896 2131
rect 1215 2131 1221 2132
rect 1215 2130 1216 2131
rect 895 2128 985 2130
rect 1157 2128 1216 2130
rect 895 2127 896 2128
rect 890 2126 896 2127
rect 1215 2127 1216 2128
rect 1220 2127 1221 2131
rect 1215 2126 1221 2127
rect 1298 2131 1304 2132
rect 1298 2127 1299 2131
rect 1303 2127 1304 2131
rect 1479 2131 1485 2132
rect 1479 2130 1480 2131
rect 1445 2128 1480 2130
rect 1298 2126 1304 2127
rect 1479 2127 1480 2128
rect 1484 2127 1485 2131
rect 1479 2126 1485 2127
rect 1578 2131 1584 2132
rect 1578 2127 1579 2131
rect 1583 2127 1584 2131
rect 1578 2126 1584 2127
rect 1586 2131 1592 2132
rect 1586 2127 1587 2131
rect 1591 2130 1592 2131
rect 1850 2131 1856 2132
rect 1591 2128 1681 2130
rect 1591 2127 1592 2128
rect 1586 2126 1592 2127
rect 1850 2127 1851 2131
rect 1855 2127 1856 2131
rect 1850 2126 1856 2127
rect 1866 2131 1872 2132
rect 1866 2127 1867 2131
rect 1871 2130 1872 2131
rect 1871 2128 1945 2130
rect 1871 2127 1872 2128
rect 1866 2126 1872 2127
rect 470 2121 476 2122
rect 110 2120 116 2121
rect 110 2116 111 2120
rect 115 2116 116 2120
rect 470 2117 471 2121
rect 475 2117 476 2121
rect 470 2116 476 2117
rect 566 2121 572 2122
rect 566 2117 567 2121
rect 571 2117 572 2121
rect 566 2116 572 2117
rect 678 2121 684 2122
rect 678 2117 679 2121
rect 683 2117 684 2121
rect 678 2116 684 2117
rect 806 2121 812 2122
rect 806 2117 807 2121
rect 811 2117 812 2121
rect 806 2116 812 2117
rect 942 2121 948 2122
rect 942 2117 943 2121
rect 947 2117 948 2121
rect 942 2116 948 2117
rect 1078 2121 1084 2122
rect 1078 2117 1079 2121
rect 1083 2117 1084 2121
rect 1078 2116 1084 2117
rect 1222 2121 1228 2122
rect 1222 2117 1223 2121
rect 1227 2117 1228 2121
rect 1222 2116 1228 2117
rect 1366 2121 1372 2122
rect 1366 2117 1367 2121
rect 1371 2117 1372 2121
rect 1366 2116 1372 2117
rect 1502 2121 1508 2122
rect 1502 2117 1503 2121
rect 1507 2117 1508 2121
rect 1502 2116 1508 2117
rect 1638 2121 1644 2122
rect 1638 2117 1639 2121
rect 1643 2117 1644 2121
rect 1638 2116 1644 2117
rect 1782 2121 1788 2122
rect 1782 2117 1783 2121
rect 1787 2117 1788 2121
rect 1782 2116 1788 2117
rect 1902 2121 1908 2122
rect 1902 2117 1903 2121
rect 1907 2117 1908 2121
rect 1902 2116 1908 2117
rect 2006 2120 2012 2121
rect 2006 2116 2007 2120
rect 2011 2116 2012 2120
rect 110 2115 116 2116
rect 2006 2115 2012 2116
rect 2990 2115 2996 2116
rect 2990 2111 2991 2115
rect 2995 2114 2996 2115
rect 2995 2112 3438 2114
rect 2995 2111 2996 2112
rect 2990 2110 2996 2111
rect 2046 2108 2052 2109
rect 2046 2104 2047 2108
rect 2051 2104 2052 2108
rect 2046 2103 2052 2104
rect 2278 2107 2284 2108
rect 2278 2103 2279 2107
rect 2283 2103 2284 2107
rect 2278 2102 2284 2103
rect 2390 2107 2396 2108
rect 2390 2103 2391 2107
rect 2395 2103 2396 2107
rect 2390 2102 2396 2103
rect 2510 2107 2516 2108
rect 2510 2103 2511 2107
rect 2515 2103 2516 2107
rect 2510 2102 2516 2103
rect 2630 2107 2636 2108
rect 2630 2103 2631 2107
rect 2635 2103 2636 2107
rect 2630 2102 2636 2103
rect 2758 2107 2764 2108
rect 2758 2103 2759 2107
rect 2763 2103 2764 2107
rect 2758 2102 2764 2103
rect 2894 2107 2900 2108
rect 2894 2103 2895 2107
rect 2899 2103 2900 2107
rect 2894 2102 2900 2103
rect 3038 2107 3044 2108
rect 3038 2103 3039 2107
rect 3043 2103 3044 2107
rect 3038 2102 3044 2103
rect 3190 2107 3196 2108
rect 3190 2103 3191 2107
rect 3195 2103 3196 2107
rect 3190 2102 3196 2103
rect 3350 2107 3356 2108
rect 3350 2103 3351 2107
rect 3355 2103 3356 2107
rect 3350 2102 3356 2103
rect 2354 2099 2360 2100
rect 2354 2095 2355 2099
rect 2359 2095 2360 2099
rect 2354 2094 2360 2095
rect 2382 2099 2388 2100
rect 2382 2095 2383 2099
rect 2387 2098 2388 2099
rect 2498 2099 2504 2100
rect 2387 2096 2433 2098
rect 2387 2095 2388 2096
rect 2382 2094 2388 2095
rect 2498 2095 2499 2099
rect 2503 2098 2504 2099
rect 2743 2099 2749 2100
rect 2503 2096 2553 2098
rect 2503 2095 2504 2096
rect 2498 2094 2504 2095
rect 2706 2095 2712 2096
rect 2046 2091 2052 2092
rect 2046 2087 2047 2091
rect 2051 2087 2052 2091
rect 2706 2091 2707 2095
rect 2711 2091 2712 2095
rect 2743 2095 2744 2099
rect 2748 2098 2749 2099
rect 3436 2098 3438 2112
rect 3942 2108 3948 2109
rect 3518 2107 3524 2108
rect 3518 2103 3519 2107
rect 3523 2103 3524 2107
rect 3518 2102 3524 2103
rect 3686 2107 3692 2108
rect 3686 2103 3687 2107
rect 3691 2103 3692 2107
rect 3686 2102 3692 2103
rect 3838 2107 3844 2108
rect 3838 2103 3839 2107
rect 3843 2103 3844 2107
rect 3942 2104 3943 2108
rect 3947 2104 3948 2108
rect 3942 2103 3948 2104
rect 3838 2102 3844 2103
rect 3830 2099 3836 2100
rect 2748 2096 2801 2098
rect 3436 2096 3561 2098
rect 2748 2095 2749 2096
rect 2743 2094 2749 2095
rect 2970 2095 2976 2096
rect 2706 2090 2712 2091
rect 2970 2091 2971 2095
rect 2975 2091 2976 2095
rect 2970 2090 2976 2091
rect 3114 2095 3120 2096
rect 3114 2091 3115 2095
rect 3119 2091 3120 2095
rect 3114 2090 3120 2091
rect 3266 2095 3272 2096
rect 3266 2091 3267 2095
rect 3271 2091 3272 2095
rect 3266 2090 3272 2091
rect 3426 2095 3432 2096
rect 3426 2091 3427 2095
rect 3431 2091 3432 2095
rect 3426 2090 3432 2091
rect 3762 2095 3768 2096
rect 3762 2091 3763 2095
rect 3767 2091 3768 2095
rect 3830 2095 3831 2099
rect 3835 2098 3836 2099
rect 3835 2096 3881 2098
rect 3835 2095 3836 2096
rect 3830 2094 3836 2095
rect 3762 2090 3768 2091
rect 3942 2091 3948 2092
rect 2046 2086 2052 2087
rect 2278 2088 2284 2089
rect 2278 2084 2279 2088
rect 2283 2084 2284 2088
rect 2278 2083 2284 2084
rect 2390 2088 2396 2089
rect 2390 2084 2391 2088
rect 2395 2084 2396 2088
rect 2390 2083 2396 2084
rect 2510 2088 2516 2089
rect 2510 2084 2511 2088
rect 2515 2084 2516 2088
rect 2510 2083 2516 2084
rect 2630 2088 2636 2089
rect 2630 2084 2631 2088
rect 2635 2084 2636 2088
rect 2630 2083 2636 2084
rect 2758 2088 2764 2089
rect 2758 2084 2759 2088
rect 2763 2084 2764 2088
rect 2758 2083 2764 2084
rect 2894 2088 2900 2089
rect 2894 2084 2895 2088
rect 2899 2084 2900 2088
rect 2894 2083 2900 2084
rect 3038 2088 3044 2089
rect 3038 2084 3039 2088
rect 3043 2084 3044 2088
rect 3038 2083 3044 2084
rect 3190 2088 3196 2089
rect 3190 2084 3191 2088
rect 3195 2084 3196 2088
rect 3190 2083 3196 2084
rect 3350 2088 3356 2089
rect 3350 2084 3351 2088
rect 3355 2084 3356 2088
rect 3350 2083 3356 2084
rect 3518 2088 3524 2089
rect 3518 2084 3519 2088
rect 3523 2084 3524 2088
rect 3518 2083 3524 2084
rect 3686 2088 3692 2089
rect 3686 2084 3687 2088
rect 3691 2084 3692 2088
rect 3686 2083 3692 2084
rect 3838 2088 3844 2089
rect 3838 2084 3839 2088
rect 3843 2084 3844 2088
rect 3942 2087 3943 2091
rect 3947 2087 3948 2091
rect 3942 2086 3948 2087
rect 3838 2083 3844 2084
rect 110 2068 116 2069
rect 2006 2068 2012 2069
rect 110 2064 111 2068
rect 115 2064 116 2068
rect 110 2063 116 2064
rect 622 2067 628 2068
rect 622 2063 623 2067
rect 627 2063 628 2067
rect 622 2062 628 2063
rect 734 2067 740 2068
rect 734 2063 735 2067
rect 739 2063 740 2067
rect 734 2062 740 2063
rect 854 2067 860 2068
rect 854 2063 855 2067
rect 859 2063 860 2067
rect 854 2062 860 2063
rect 982 2067 988 2068
rect 982 2063 983 2067
rect 987 2063 988 2067
rect 982 2062 988 2063
rect 1118 2067 1124 2068
rect 1118 2063 1119 2067
rect 1123 2063 1124 2067
rect 1118 2062 1124 2063
rect 1254 2067 1260 2068
rect 1254 2063 1255 2067
rect 1259 2063 1260 2067
rect 1254 2062 1260 2063
rect 1390 2067 1396 2068
rect 1390 2063 1391 2067
rect 1395 2063 1396 2067
rect 1390 2062 1396 2063
rect 1526 2067 1532 2068
rect 1526 2063 1527 2067
rect 1531 2063 1532 2067
rect 1526 2062 1532 2063
rect 1654 2067 1660 2068
rect 1654 2063 1655 2067
rect 1659 2063 1660 2067
rect 1654 2062 1660 2063
rect 1790 2067 1796 2068
rect 1790 2063 1791 2067
rect 1795 2063 1796 2067
rect 1790 2062 1796 2063
rect 1902 2067 1908 2068
rect 1902 2063 1903 2067
rect 1907 2063 1908 2067
rect 2006 2064 2007 2068
rect 2011 2064 2012 2068
rect 2006 2063 2012 2064
rect 2331 2067 2337 2068
rect 2331 2063 2332 2067
rect 2336 2066 2337 2067
rect 2382 2067 2388 2068
rect 2382 2066 2383 2067
rect 2336 2064 2383 2066
rect 2336 2063 2337 2064
rect 1902 2062 1908 2063
rect 2331 2062 2337 2063
rect 2382 2063 2383 2064
rect 2387 2063 2388 2067
rect 2382 2062 2388 2063
rect 2443 2067 2449 2068
rect 2443 2063 2444 2067
rect 2448 2066 2449 2067
rect 2498 2067 2504 2068
rect 2498 2066 2499 2067
rect 2448 2064 2499 2066
rect 2448 2063 2449 2064
rect 2443 2062 2449 2063
rect 2498 2063 2499 2064
rect 2503 2063 2504 2067
rect 2683 2067 2689 2068
rect 2498 2062 2504 2063
rect 2518 2063 2524 2064
rect 1071 2059 1077 2060
rect 698 2055 704 2056
rect 110 2051 116 2052
rect 110 2047 111 2051
rect 115 2047 116 2051
rect 698 2051 699 2055
rect 703 2051 704 2055
rect 698 2050 704 2051
rect 810 2055 816 2056
rect 810 2051 811 2055
rect 815 2051 816 2055
rect 810 2050 816 2051
rect 930 2055 936 2056
rect 930 2051 931 2055
rect 935 2051 936 2055
rect 930 2050 936 2051
rect 1058 2055 1064 2056
rect 1058 2051 1059 2055
rect 1063 2051 1064 2055
rect 1071 2055 1072 2059
rect 1076 2058 1077 2059
rect 1730 2059 1736 2060
rect 1076 2056 1161 2058
rect 1076 2055 1077 2056
rect 1071 2054 1077 2055
rect 1330 2055 1336 2056
rect 1058 2050 1064 2051
rect 1330 2051 1331 2055
rect 1335 2051 1336 2055
rect 1503 2055 1509 2056
rect 1503 2054 1504 2055
rect 1469 2052 1504 2054
rect 1330 2050 1336 2051
rect 1503 2051 1504 2052
rect 1508 2051 1509 2055
rect 1503 2050 1509 2051
rect 1602 2055 1608 2056
rect 1602 2051 1603 2055
rect 1607 2051 1608 2055
rect 1730 2055 1731 2059
rect 1735 2055 1736 2059
rect 2518 2059 2519 2063
rect 2523 2062 2524 2063
rect 2563 2063 2569 2064
rect 2563 2062 2564 2063
rect 2523 2060 2564 2062
rect 2523 2059 2524 2060
rect 2518 2058 2524 2059
rect 2563 2059 2564 2060
rect 2568 2059 2569 2063
rect 2683 2063 2684 2067
rect 2688 2066 2689 2067
rect 2743 2067 2749 2068
rect 2743 2066 2744 2067
rect 2688 2064 2744 2066
rect 2688 2063 2689 2064
rect 2683 2062 2689 2063
rect 2743 2063 2744 2064
rect 2748 2063 2749 2067
rect 2743 2062 2749 2063
rect 2811 2067 2817 2068
rect 2811 2063 2812 2067
rect 2816 2066 2817 2067
rect 2850 2067 2856 2068
rect 2850 2066 2851 2067
rect 2816 2064 2851 2066
rect 2816 2063 2817 2064
rect 2811 2062 2817 2063
rect 2850 2063 2851 2064
rect 2855 2063 2856 2067
rect 2970 2067 2976 2068
rect 2850 2062 2856 2063
rect 2947 2063 2953 2064
rect 2563 2058 2569 2059
rect 2947 2059 2948 2063
rect 2952 2062 2953 2063
rect 2970 2063 2971 2067
rect 2975 2066 2976 2067
rect 3091 2067 3097 2068
rect 3091 2066 3092 2067
rect 2975 2064 3092 2066
rect 2975 2063 2976 2064
rect 2970 2062 2976 2063
rect 3091 2063 3092 2064
rect 3096 2063 3097 2067
rect 3091 2062 3097 2063
rect 3114 2067 3120 2068
rect 3114 2063 3115 2067
rect 3119 2066 3120 2067
rect 3243 2067 3249 2068
rect 3243 2066 3244 2067
rect 3119 2064 3244 2066
rect 3119 2063 3120 2064
rect 3114 2062 3120 2063
rect 3243 2063 3244 2064
rect 3248 2063 3249 2067
rect 3243 2062 3249 2063
rect 3266 2067 3272 2068
rect 3266 2063 3267 2067
rect 3271 2066 3272 2067
rect 3403 2067 3409 2068
rect 3403 2066 3404 2067
rect 3271 2064 3404 2066
rect 3271 2063 3272 2064
rect 3266 2062 3272 2063
rect 3403 2063 3404 2064
rect 3408 2063 3409 2067
rect 3403 2062 3409 2063
rect 3426 2067 3432 2068
rect 3426 2063 3427 2067
rect 3431 2066 3432 2067
rect 3571 2067 3577 2068
rect 3571 2066 3572 2067
rect 3431 2064 3572 2066
rect 3431 2063 3432 2064
rect 3426 2062 3432 2063
rect 3571 2063 3572 2064
rect 3576 2063 3577 2067
rect 3762 2067 3768 2068
rect 3571 2062 3577 2063
rect 3730 2063 3736 2064
rect 2952 2060 2966 2062
rect 2952 2059 2953 2060
rect 2947 2058 2953 2059
rect 2964 2058 2966 2060
rect 3378 2059 3384 2060
rect 3378 2058 3379 2059
rect 2964 2056 3379 2058
rect 1730 2054 1736 2055
rect 1866 2055 1872 2056
rect 1602 2050 1608 2051
rect 1866 2051 1867 2055
rect 1871 2051 1872 2055
rect 1866 2050 1872 2051
rect 1978 2055 1984 2056
rect 1978 2051 1979 2055
rect 1983 2051 1984 2055
rect 3378 2055 3379 2056
rect 3383 2055 3384 2059
rect 3730 2059 3731 2063
rect 3735 2062 3736 2063
rect 3739 2063 3745 2064
rect 3739 2062 3740 2063
rect 3735 2060 3740 2062
rect 3735 2059 3736 2060
rect 3730 2058 3736 2059
rect 3739 2059 3740 2060
rect 3744 2059 3745 2063
rect 3762 2063 3763 2067
rect 3767 2066 3768 2067
rect 3891 2067 3897 2068
rect 3891 2066 3892 2067
rect 3767 2064 3892 2066
rect 3767 2063 3768 2064
rect 3762 2062 3768 2063
rect 3891 2063 3892 2064
rect 3896 2063 3897 2067
rect 3891 2062 3897 2063
rect 3739 2058 3745 2059
rect 3378 2054 3384 2055
rect 1978 2050 1984 2051
rect 2006 2051 2012 2052
rect 110 2046 116 2047
rect 622 2048 628 2049
rect 622 2044 623 2048
rect 627 2044 628 2048
rect 622 2043 628 2044
rect 734 2048 740 2049
rect 734 2044 735 2048
rect 739 2044 740 2048
rect 734 2043 740 2044
rect 854 2048 860 2049
rect 854 2044 855 2048
rect 859 2044 860 2048
rect 854 2043 860 2044
rect 982 2048 988 2049
rect 982 2044 983 2048
rect 987 2044 988 2048
rect 982 2043 988 2044
rect 1118 2048 1124 2049
rect 1118 2044 1119 2048
rect 1123 2044 1124 2048
rect 1118 2043 1124 2044
rect 1254 2048 1260 2049
rect 1254 2044 1255 2048
rect 1259 2044 1260 2048
rect 1254 2043 1260 2044
rect 1390 2048 1396 2049
rect 1390 2044 1391 2048
rect 1395 2044 1396 2048
rect 1390 2043 1396 2044
rect 1526 2048 1532 2049
rect 1526 2044 1527 2048
rect 1531 2044 1532 2048
rect 1526 2043 1532 2044
rect 1654 2048 1660 2049
rect 1654 2044 1655 2048
rect 1659 2044 1660 2048
rect 1654 2043 1660 2044
rect 1790 2048 1796 2049
rect 1790 2044 1791 2048
rect 1795 2044 1796 2048
rect 1790 2043 1796 2044
rect 1902 2048 1908 2049
rect 1902 2044 1903 2048
rect 1907 2044 1908 2048
rect 2006 2047 2007 2051
rect 2011 2047 2012 2051
rect 2006 2046 2012 2047
rect 1902 2043 1908 2044
rect 2402 2043 2408 2044
rect 2379 2041 2385 2042
rect 2379 2037 2380 2041
rect 2384 2037 2385 2041
rect 2402 2039 2403 2043
rect 2407 2042 2408 2043
rect 2483 2043 2489 2044
rect 2483 2042 2484 2043
rect 2407 2040 2484 2042
rect 2407 2039 2408 2040
rect 2402 2038 2408 2039
rect 2483 2039 2484 2040
rect 2488 2039 2489 2043
rect 2483 2038 2489 2039
rect 2587 2043 2593 2044
rect 2587 2039 2588 2043
rect 2592 2042 2593 2043
rect 2618 2043 2624 2044
rect 2618 2042 2619 2043
rect 2592 2040 2619 2042
rect 2592 2039 2593 2040
rect 2587 2038 2593 2039
rect 2618 2039 2619 2040
rect 2623 2039 2624 2043
rect 2618 2038 2624 2039
rect 2699 2043 2708 2044
rect 2699 2039 2700 2043
rect 2707 2039 2708 2043
rect 2699 2038 2708 2039
rect 2827 2043 2833 2044
rect 2827 2039 2828 2043
rect 2832 2042 2833 2043
rect 2842 2043 2848 2044
rect 2842 2042 2843 2043
rect 2832 2040 2843 2042
rect 2832 2039 2833 2040
rect 2827 2038 2833 2039
rect 2842 2039 2843 2040
rect 2847 2039 2848 2043
rect 2842 2038 2848 2039
rect 2850 2043 2856 2044
rect 2850 2039 2851 2043
rect 2855 2042 2856 2043
rect 2971 2043 2977 2044
rect 2971 2042 2972 2043
rect 2855 2040 2972 2042
rect 2855 2039 2856 2040
rect 2850 2038 2856 2039
rect 2971 2039 2972 2040
rect 2976 2039 2977 2043
rect 2971 2038 2977 2039
rect 2994 2043 3000 2044
rect 2994 2039 2995 2043
rect 2999 2042 3000 2043
rect 3131 2043 3137 2044
rect 3131 2042 3132 2043
rect 2999 2040 3132 2042
rect 2999 2039 3000 2040
rect 2994 2038 3000 2039
rect 3131 2039 3132 2040
rect 3136 2039 3137 2043
rect 3131 2038 3137 2039
rect 3154 2043 3160 2044
rect 3154 2039 3155 2043
rect 3159 2042 3160 2043
rect 3315 2043 3321 2044
rect 3315 2042 3316 2043
rect 3159 2040 3316 2042
rect 3159 2039 3160 2040
rect 3154 2038 3160 2039
rect 3315 2039 3316 2040
rect 3320 2039 3321 2043
rect 3315 2038 3321 2039
rect 3338 2043 3344 2044
rect 3338 2039 3339 2043
rect 3343 2042 3344 2043
rect 3507 2043 3513 2044
rect 3507 2042 3508 2043
rect 3343 2040 3508 2042
rect 3343 2039 3344 2040
rect 3338 2038 3344 2039
rect 3507 2039 3508 2040
rect 3512 2039 3513 2043
rect 3507 2038 3513 2039
rect 3707 2043 3713 2044
rect 3707 2039 3708 2043
rect 3712 2042 3713 2043
rect 3738 2043 3744 2044
rect 3738 2042 3739 2043
rect 3712 2040 3739 2042
rect 3712 2039 3713 2040
rect 3707 2038 3713 2039
rect 3738 2039 3739 2040
rect 3743 2039 3744 2043
rect 3738 2038 3744 2039
rect 3891 2043 3897 2044
rect 3891 2039 3892 2043
rect 3896 2042 3897 2043
rect 3906 2043 3912 2044
rect 3906 2042 3907 2043
rect 3896 2040 3907 2042
rect 3896 2039 3897 2040
rect 3891 2038 3897 2039
rect 3906 2039 3907 2040
rect 3911 2039 3912 2043
rect 3906 2038 3912 2039
rect 2379 2036 2385 2037
rect 2380 2034 2382 2036
rect 2526 2035 2532 2036
rect 2526 2034 2527 2035
rect 2380 2032 2527 2034
rect 2526 2031 2527 2032
rect 2531 2031 2532 2035
rect 2526 2030 2532 2031
rect 698 2027 704 2028
rect 675 2023 681 2024
rect 675 2019 676 2023
rect 680 2022 681 2023
rect 698 2023 699 2027
rect 703 2026 704 2027
rect 787 2027 793 2028
rect 787 2026 788 2027
rect 703 2024 788 2026
rect 703 2023 704 2024
rect 698 2022 704 2023
rect 787 2023 788 2024
rect 792 2023 793 2027
rect 787 2022 793 2023
rect 810 2027 816 2028
rect 810 2023 811 2027
rect 815 2026 816 2027
rect 907 2027 913 2028
rect 907 2026 908 2027
rect 815 2024 908 2026
rect 815 2023 816 2024
rect 810 2022 816 2023
rect 907 2023 908 2024
rect 912 2023 913 2027
rect 907 2022 913 2023
rect 930 2027 936 2028
rect 930 2023 931 2027
rect 935 2026 936 2027
rect 1035 2027 1041 2028
rect 1035 2026 1036 2027
rect 935 2024 1036 2026
rect 935 2023 936 2024
rect 930 2022 936 2023
rect 1035 2023 1036 2024
rect 1040 2023 1041 2027
rect 1035 2022 1041 2023
rect 1058 2027 1064 2028
rect 1058 2023 1059 2027
rect 1063 2026 1064 2027
rect 1171 2027 1177 2028
rect 1171 2026 1172 2027
rect 1063 2024 1172 2026
rect 1063 2023 1064 2024
rect 1058 2022 1064 2023
rect 1171 2023 1172 2024
rect 1176 2023 1177 2027
rect 1171 2022 1177 2023
rect 1298 2027 1304 2028
rect 1298 2023 1299 2027
rect 1303 2026 1304 2027
rect 1307 2027 1313 2028
rect 1307 2026 1308 2027
rect 1303 2024 1308 2026
rect 1303 2023 1304 2024
rect 1298 2022 1304 2023
rect 1307 2023 1308 2024
rect 1312 2023 1313 2027
rect 1503 2027 1509 2028
rect 1307 2022 1313 2023
rect 1443 2023 1449 2024
rect 680 2020 694 2022
rect 680 2019 681 2020
rect 675 2018 681 2019
rect 692 2018 694 2020
rect 810 2019 816 2020
rect 810 2018 811 2019
rect 692 2016 811 2018
rect 810 2015 811 2016
rect 815 2015 816 2019
rect 1443 2019 1444 2023
rect 1448 2022 1449 2023
rect 1466 2023 1472 2024
rect 1466 2022 1467 2023
rect 1448 2020 1467 2022
rect 1448 2019 1449 2020
rect 1443 2018 1449 2019
rect 1466 2019 1467 2020
rect 1471 2019 1472 2023
rect 1503 2023 1504 2027
rect 1508 2026 1509 2027
rect 1579 2027 1585 2028
rect 1579 2026 1580 2027
rect 1508 2024 1580 2026
rect 1508 2023 1509 2024
rect 1503 2022 1509 2023
rect 1579 2023 1580 2024
rect 1584 2023 1585 2027
rect 1579 2022 1585 2023
rect 1602 2027 1608 2028
rect 1602 2023 1603 2027
rect 1607 2026 1608 2027
rect 1707 2027 1713 2028
rect 1707 2026 1708 2027
rect 1607 2024 1708 2026
rect 1607 2023 1608 2024
rect 1602 2022 1608 2023
rect 1707 2023 1708 2024
rect 1712 2023 1713 2027
rect 1707 2022 1713 2023
rect 1843 2027 1852 2028
rect 1843 2023 1844 2027
rect 1851 2023 1852 2027
rect 1843 2022 1852 2023
rect 1866 2027 1872 2028
rect 1866 2023 1867 2027
rect 1871 2026 1872 2027
rect 1955 2027 1961 2028
rect 1955 2026 1956 2027
rect 1871 2024 1956 2026
rect 1871 2023 1872 2024
rect 1866 2022 1872 2023
rect 1955 2023 1956 2024
rect 1960 2023 1961 2027
rect 1955 2022 1961 2023
rect 1466 2018 1472 2019
rect 2326 2020 2332 2021
rect 810 2014 816 2015
rect 2046 2017 2052 2018
rect 2046 2013 2047 2017
rect 2051 2013 2052 2017
rect 2326 2016 2327 2020
rect 2331 2016 2332 2020
rect 2326 2015 2332 2016
rect 2430 2020 2436 2021
rect 2430 2016 2431 2020
rect 2435 2016 2436 2020
rect 2430 2015 2436 2016
rect 2534 2020 2540 2021
rect 2534 2016 2535 2020
rect 2539 2016 2540 2020
rect 2534 2015 2540 2016
rect 2646 2020 2652 2021
rect 2646 2016 2647 2020
rect 2651 2016 2652 2020
rect 2646 2015 2652 2016
rect 2774 2020 2780 2021
rect 2774 2016 2775 2020
rect 2779 2016 2780 2020
rect 2774 2015 2780 2016
rect 2918 2020 2924 2021
rect 2918 2016 2919 2020
rect 2923 2016 2924 2020
rect 2918 2015 2924 2016
rect 3078 2020 3084 2021
rect 3078 2016 3079 2020
rect 3083 2016 3084 2020
rect 3078 2015 3084 2016
rect 3262 2020 3268 2021
rect 3262 2016 3263 2020
rect 3267 2016 3268 2020
rect 3262 2015 3268 2016
rect 3454 2020 3460 2021
rect 3454 2016 3455 2020
rect 3459 2016 3460 2020
rect 3454 2015 3460 2016
rect 3654 2020 3660 2021
rect 3654 2016 3655 2020
rect 3659 2016 3660 2020
rect 3654 2015 3660 2016
rect 3838 2020 3844 2021
rect 3838 2016 3839 2020
rect 3843 2016 3844 2020
rect 3838 2015 3844 2016
rect 3942 2017 3948 2018
rect 2046 2012 2052 2013
rect 3942 2013 3943 2017
rect 3947 2013 3948 2017
rect 3942 2012 3948 2013
rect 2402 2011 2408 2012
rect 499 2007 505 2008
rect 499 2003 500 2007
rect 504 2006 505 2007
rect 514 2007 520 2008
rect 514 2006 515 2007
rect 504 2004 515 2006
rect 504 2003 505 2004
rect 499 2002 505 2003
rect 514 2003 515 2004
rect 519 2003 520 2007
rect 514 2002 520 2003
rect 522 2007 528 2008
rect 522 2003 523 2007
rect 527 2006 528 2007
rect 627 2007 633 2008
rect 627 2006 628 2007
rect 527 2004 628 2006
rect 527 2003 528 2004
rect 522 2002 528 2003
rect 627 2003 628 2004
rect 632 2003 633 2007
rect 627 2002 633 2003
rect 650 2007 656 2008
rect 650 2003 651 2007
rect 655 2006 656 2007
rect 779 2007 785 2008
rect 779 2006 780 2007
rect 655 2004 780 2006
rect 655 2003 656 2004
rect 650 2002 656 2003
rect 779 2003 780 2004
rect 784 2003 785 2007
rect 779 2002 785 2003
rect 802 2007 808 2008
rect 802 2003 803 2007
rect 807 2006 808 2007
rect 939 2007 945 2008
rect 939 2006 940 2007
rect 807 2004 940 2006
rect 807 2003 808 2004
rect 802 2002 808 2003
rect 939 2003 940 2004
rect 944 2003 945 2007
rect 939 2002 945 2003
rect 1106 2007 1113 2008
rect 1106 2003 1107 2007
rect 1112 2003 1113 2007
rect 1106 2002 1113 2003
rect 1283 2007 1289 2008
rect 1283 2003 1284 2007
rect 1288 2006 1289 2007
rect 1330 2007 1336 2008
rect 1330 2006 1331 2007
rect 1288 2004 1331 2006
rect 1288 2003 1289 2004
rect 1283 2002 1289 2003
rect 1330 2003 1331 2004
rect 1335 2003 1336 2007
rect 1330 2002 1336 2003
rect 1451 2007 1457 2008
rect 1451 2003 1452 2007
rect 1456 2006 1457 2007
rect 1486 2007 1492 2008
rect 1486 2006 1487 2007
rect 1456 2004 1487 2006
rect 1456 2003 1457 2004
rect 1451 2002 1457 2003
rect 1486 2003 1487 2004
rect 1491 2003 1492 2007
rect 1486 2002 1492 2003
rect 1627 2007 1633 2008
rect 1627 2003 1628 2007
rect 1632 2006 1633 2007
rect 1662 2007 1668 2008
rect 1662 2006 1663 2007
rect 1632 2004 1663 2006
rect 1632 2003 1633 2004
rect 1627 2002 1633 2003
rect 1662 2003 1663 2004
rect 1667 2003 1668 2007
rect 1662 2002 1668 2003
rect 1803 2007 1809 2008
rect 1803 2003 1804 2007
rect 1808 2006 1809 2007
rect 1834 2007 1840 2008
rect 1834 2006 1835 2007
rect 1808 2004 1835 2006
rect 1808 2003 1809 2004
rect 1803 2002 1809 2003
rect 1834 2003 1835 2004
rect 1839 2003 1840 2007
rect 1834 2002 1840 2003
rect 1955 2007 1961 2008
rect 1955 2003 1956 2007
rect 1960 2006 1961 2007
rect 1978 2007 1984 2008
rect 1978 2006 1979 2007
rect 1960 2004 1979 2006
rect 1960 2003 1961 2004
rect 1955 2002 1961 2003
rect 1978 2003 1979 2004
rect 1983 2003 1984 2007
rect 2402 2007 2403 2011
rect 2407 2007 2408 2011
rect 2518 2011 2524 2012
rect 2518 2010 2519 2011
rect 2509 2008 2519 2010
rect 2402 2006 2408 2007
rect 2518 2007 2519 2008
rect 2523 2007 2524 2011
rect 2518 2006 2524 2007
rect 2526 2011 2532 2012
rect 2526 2007 2527 2011
rect 2531 2010 2532 2011
rect 2714 2011 2720 2012
rect 2531 2008 2577 2010
rect 2531 2007 2532 2008
rect 2526 2006 2532 2007
rect 2714 2007 2715 2011
rect 2719 2007 2720 2011
rect 2714 2006 2720 2007
rect 2850 2011 2856 2012
rect 2850 2007 2851 2011
rect 2855 2007 2856 2011
rect 2850 2006 2856 2007
rect 2994 2011 3000 2012
rect 2994 2007 2995 2011
rect 2999 2007 3000 2011
rect 2994 2006 3000 2007
rect 3154 2011 3160 2012
rect 3154 2007 3155 2011
rect 3159 2007 3160 2011
rect 3154 2006 3160 2007
rect 3338 2011 3344 2012
rect 3338 2007 3339 2011
rect 3343 2007 3344 2011
rect 3338 2006 3344 2007
rect 3378 2011 3384 2012
rect 3378 2007 3379 2011
rect 3383 2010 3384 2011
rect 3730 2011 3736 2012
rect 3383 2008 3497 2010
rect 3383 2007 3384 2008
rect 3378 2006 3384 2007
rect 3730 2007 3731 2011
rect 3735 2007 3736 2011
rect 3730 2006 3736 2007
rect 3738 2011 3744 2012
rect 3738 2007 3739 2011
rect 3743 2010 3744 2011
rect 3743 2008 3881 2010
rect 3743 2007 3744 2008
rect 3738 2006 3744 2007
rect 1978 2002 1984 2003
rect 2326 2001 2332 2002
rect 2046 2000 2052 2001
rect 2046 1996 2047 2000
rect 2051 1996 2052 2000
rect 2326 1997 2327 2001
rect 2331 1997 2332 2001
rect 2326 1996 2332 1997
rect 2430 2001 2436 2002
rect 2430 1997 2431 2001
rect 2435 1997 2436 2001
rect 2430 1996 2436 1997
rect 2534 2001 2540 2002
rect 2534 1997 2535 2001
rect 2539 1997 2540 2001
rect 2534 1996 2540 1997
rect 2646 2001 2652 2002
rect 2646 1997 2647 2001
rect 2651 1997 2652 2001
rect 2646 1996 2652 1997
rect 2774 2001 2780 2002
rect 2774 1997 2775 2001
rect 2779 1997 2780 2001
rect 2774 1996 2780 1997
rect 2918 2001 2924 2002
rect 2918 1997 2919 2001
rect 2923 1997 2924 2001
rect 2918 1996 2924 1997
rect 3078 2001 3084 2002
rect 3078 1997 3079 2001
rect 3083 1997 3084 2001
rect 3078 1996 3084 1997
rect 3262 2001 3268 2002
rect 3262 1997 3263 2001
rect 3267 1997 3268 2001
rect 3262 1996 3268 1997
rect 3454 2001 3460 2002
rect 3454 1997 3455 2001
rect 3459 1997 3460 2001
rect 3454 1996 3460 1997
rect 3654 2001 3660 2002
rect 3654 1997 3655 2001
rect 3659 1997 3660 2001
rect 3654 1996 3660 1997
rect 3838 2001 3844 2002
rect 3838 1997 3839 2001
rect 3843 1997 3844 2001
rect 3838 1996 3844 1997
rect 3942 2000 3948 2001
rect 3942 1996 3943 2000
rect 3947 1996 3948 2000
rect 2046 1995 2052 1996
rect 3942 1995 3948 1996
rect 446 1984 452 1985
rect 110 1981 116 1982
rect 110 1977 111 1981
rect 115 1977 116 1981
rect 446 1980 447 1984
rect 451 1980 452 1984
rect 446 1979 452 1980
rect 574 1984 580 1985
rect 574 1980 575 1984
rect 579 1980 580 1984
rect 574 1979 580 1980
rect 726 1984 732 1985
rect 726 1980 727 1984
rect 731 1980 732 1984
rect 726 1979 732 1980
rect 886 1984 892 1985
rect 886 1980 887 1984
rect 891 1980 892 1984
rect 886 1979 892 1980
rect 1054 1984 1060 1985
rect 1054 1980 1055 1984
rect 1059 1980 1060 1984
rect 1054 1979 1060 1980
rect 1230 1984 1236 1985
rect 1230 1980 1231 1984
rect 1235 1980 1236 1984
rect 1230 1979 1236 1980
rect 1398 1984 1404 1985
rect 1398 1980 1399 1984
rect 1403 1980 1404 1984
rect 1398 1979 1404 1980
rect 1574 1984 1580 1985
rect 1574 1980 1575 1984
rect 1579 1980 1580 1984
rect 1574 1979 1580 1980
rect 1750 1984 1756 1985
rect 1750 1980 1751 1984
rect 1755 1980 1756 1984
rect 1750 1979 1756 1980
rect 1902 1984 1908 1985
rect 1902 1980 1903 1984
rect 1907 1980 1908 1984
rect 1902 1979 1908 1980
rect 2006 1981 2012 1982
rect 110 1976 116 1977
rect 2006 1977 2007 1981
rect 2011 1977 2012 1981
rect 2006 1976 2012 1977
rect 522 1975 528 1976
rect 522 1971 523 1975
rect 527 1971 528 1975
rect 522 1970 528 1971
rect 650 1975 656 1976
rect 650 1971 651 1975
rect 655 1971 656 1975
rect 650 1970 656 1971
rect 802 1975 808 1976
rect 802 1971 803 1975
rect 807 1971 808 1975
rect 802 1970 808 1971
rect 810 1975 816 1976
rect 810 1971 811 1975
rect 815 1974 816 1975
rect 1122 1975 1128 1976
rect 815 1972 929 1974
rect 815 1971 816 1972
rect 810 1970 816 1971
rect 1122 1971 1123 1975
rect 1127 1971 1128 1975
rect 1122 1970 1128 1971
rect 1202 1975 1208 1976
rect 1202 1971 1203 1975
rect 1207 1974 1208 1975
rect 1466 1975 1472 1976
rect 1207 1972 1273 1974
rect 1207 1971 1208 1972
rect 1202 1970 1208 1971
rect 1466 1971 1467 1975
rect 1471 1971 1472 1975
rect 1466 1970 1472 1971
rect 1486 1975 1492 1976
rect 1486 1971 1487 1975
rect 1491 1974 1492 1975
rect 1662 1975 1668 1976
rect 1491 1972 1617 1974
rect 1491 1971 1492 1972
rect 1486 1970 1492 1971
rect 1662 1971 1663 1975
rect 1667 1974 1668 1975
rect 1834 1975 1840 1976
rect 1667 1972 1793 1974
rect 1667 1971 1668 1972
rect 1662 1970 1668 1971
rect 1834 1971 1835 1975
rect 1839 1974 1840 1975
rect 1839 1972 1945 1974
rect 1839 1971 1840 1972
rect 1834 1970 1840 1971
rect 446 1965 452 1966
rect 110 1964 116 1965
rect 110 1960 111 1964
rect 115 1960 116 1964
rect 446 1961 447 1965
rect 451 1961 452 1965
rect 446 1960 452 1961
rect 574 1965 580 1966
rect 574 1961 575 1965
rect 579 1961 580 1965
rect 574 1960 580 1961
rect 726 1965 732 1966
rect 726 1961 727 1965
rect 731 1961 732 1965
rect 726 1960 732 1961
rect 886 1965 892 1966
rect 886 1961 887 1965
rect 891 1961 892 1965
rect 886 1960 892 1961
rect 1054 1965 1060 1966
rect 1054 1961 1055 1965
rect 1059 1961 1060 1965
rect 1054 1960 1060 1961
rect 1230 1965 1236 1966
rect 1230 1961 1231 1965
rect 1235 1961 1236 1965
rect 1230 1960 1236 1961
rect 1398 1965 1404 1966
rect 1398 1961 1399 1965
rect 1403 1961 1404 1965
rect 1398 1960 1404 1961
rect 1574 1965 1580 1966
rect 1574 1961 1575 1965
rect 1579 1961 1580 1965
rect 1574 1960 1580 1961
rect 1750 1965 1756 1966
rect 1750 1961 1751 1965
rect 1755 1961 1756 1965
rect 1750 1960 1756 1961
rect 1902 1965 1908 1966
rect 1902 1961 1903 1965
rect 1907 1961 1908 1965
rect 1902 1960 1908 1961
rect 2006 1964 2012 1965
rect 2006 1960 2007 1964
rect 2011 1960 2012 1964
rect 110 1959 116 1960
rect 2006 1959 2012 1960
rect 2046 1944 2052 1945
rect 3942 1944 3948 1945
rect 2046 1940 2047 1944
rect 2051 1940 2052 1944
rect 2046 1939 2052 1940
rect 2254 1943 2260 1944
rect 2254 1939 2255 1943
rect 2259 1939 2260 1943
rect 2254 1938 2260 1939
rect 2350 1943 2356 1944
rect 2350 1939 2351 1943
rect 2355 1939 2356 1943
rect 2350 1938 2356 1939
rect 2446 1943 2452 1944
rect 2446 1939 2447 1943
rect 2451 1939 2452 1943
rect 2446 1938 2452 1939
rect 2542 1943 2548 1944
rect 2542 1939 2543 1943
rect 2547 1939 2548 1943
rect 2542 1938 2548 1939
rect 2646 1943 2652 1944
rect 2646 1939 2647 1943
rect 2651 1939 2652 1943
rect 2646 1938 2652 1939
rect 2766 1943 2772 1944
rect 2766 1939 2767 1943
rect 2771 1939 2772 1943
rect 2766 1938 2772 1939
rect 2918 1943 2924 1944
rect 2918 1939 2919 1943
rect 2923 1939 2924 1943
rect 2918 1938 2924 1939
rect 3102 1943 3108 1944
rect 3102 1939 3103 1943
rect 3107 1939 3108 1943
rect 3102 1938 3108 1939
rect 3318 1943 3324 1944
rect 3318 1939 3319 1943
rect 3323 1939 3324 1943
rect 3318 1938 3324 1939
rect 3542 1943 3548 1944
rect 3542 1939 3543 1943
rect 3547 1939 3548 1943
rect 3542 1938 3548 1939
rect 3774 1943 3780 1944
rect 3774 1939 3775 1943
rect 3779 1939 3780 1943
rect 3942 1940 3943 1944
rect 3947 1940 3948 1944
rect 3942 1939 3948 1940
rect 3774 1938 3780 1939
rect 2618 1935 2624 1936
rect 2330 1931 2336 1932
rect 2046 1927 2052 1928
rect 2046 1923 2047 1927
rect 2051 1923 2052 1927
rect 2330 1927 2331 1931
rect 2335 1927 2336 1931
rect 2330 1926 2336 1927
rect 2426 1931 2432 1932
rect 2426 1927 2427 1931
rect 2431 1927 2432 1931
rect 2426 1926 2432 1927
rect 2522 1931 2528 1932
rect 2522 1927 2523 1931
rect 2527 1927 2528 1931
rect 2618 1931 2619 1935
rect 2623 1931 2624 1935
rect 2618 1930 2624 1931
rect 2638 1935 2644 1936
rect 2638 1931 2639 1935
rect 2643 1934 2644 1935
rect 2842 1935 2848 1936
rect 2643 1932 2689 1934
rect 2643 1931 2644 1932
rect 2638 1930 2644 1931
rect 2842 1931 2843 1935
rect 2847 1931 2848 1935
rect 2842 1930 2848 1931
rect 2858 1935 2864 1936
rect 2858 1931 2859 1935
rect 2863 1934 2864 1935
rect 3006 1935 3012 1936
rect 2863 1932 2961 1934
rect 2863 1931 2864 1932
rect 2858 1930 2864 1931
rect 3006 1931 3007 1935
rect 3011 1934 3012 1935
rect 3186 1935 3192 1936
rect 3011 1932 3145 1934
rect 3011 1931 3012 1932
rect 3006 1930 3012 1931
rect 3186 1931 3187 1935
rect 3191 1934 3192 1935
rect 3402 1935 3408 1936
rect 3191 1932 3361 1934
rect 3191 1931 3192 1932
rect 3186 1930 3192 1931
rect 3402 1931 3403 1935
rect 3407 1934 3408 1935
rect 3750 1935 3756 1936
rect 3407 1932 3585 1934
rect 3407 1931 3408 1932
rect 3402 1930 3408 1931
rect 3750 1931 3751 1935
rect 3755 1934 3756 1935
rect 3755 1932 3817 1934
rect 3755 1931 3756 1932
rect 3750 1930 3756 1931
rect 2522 1926 2528 1927
rect 3942 1927 3948 1928
rect 2046 1922 2052 1923
rect 2254 1924 2260 1925
rect 2254 1920 2255 1924
rect 2259 1920 2260 1924
rect 2254 1919 2260 1920
rect 2350 1924 2356 1925
rect 2350 1920 2351 1924
rect 2355 1920 2356 1924
rect 2350 1919 2356 1920
rect 2446 1924 2452 1925
rect 2446 1920 2447 1924
rect 2451 1920 2452 1924
rect 2446 1919 2452 1920
rect 2542 1924 2548 1925
rect 2542 1920 2543 1924
rect 2547 1920 2548 1924
rect 2542 1919 2548 1920
rect 2646 1924 2652 1925
rect 2646 1920 2647 1924
rect 2651 1920 2652 1924
rect 2646 1919 2652 1920
rect 2766 1924 2772 1925
rect 2766 1920 2767 1924
rect 2771 1920 2772 1924
rect 2766 1919 2772 1920
rect 2918 1924 2924 1925
rect 2918 1920 2919 1924
rect 2923 1920 2924 1924
rect 2918 1919 2924 1920
rect 3102 1924 3108 1925
rect 3102 1920 3103 1924
rect 3107 1920 3108 1924
rect 3102 1919 3108 1920
rect 3318 1924 3324 1925
rect 3318 1920 3319 1924
rect 3323 1920 3324 1924
rect 3318 1919 3324 1920
rect 3542 1924 3548 1925
rect 3542 1920 3543 1924
rect 3547 1920 3548 1924
rect 3542 1919 3548 1920
rect 3774 1924 3780 1925
rect 3774 1920 3775 1924
rect 3779 1920 3780 1924
rect 3942 1923 3943 1927
rect 3947 1923 3948 1927
rect 3942 1922 3948 1923
rect 3774 1919 3780 1920
rect 110 1912 116 1913
rect 2006 1912 2012 1913
rect 110 1908 111 1912
rect 115 1908 116 1912
rect 110 1907 116 1908
rect 654 1911 660 1912
rect 654 1907 655 1911
rect 659 1907 660 1911
rect 654 1906 660 1907
rect 750 1911 756 1912
rect 750 1907 751 1911
rect 755 1907 756 1911
rect 750 1906 756 1907
rect 846 1911 852 1912
rect 846 1907 847 1911
rect 851 1907 852 1911
rect 846 1906 852 1907
rect 942 1911 948 1912
rect 942 1907 943 1911
rect 947 1907 948 1911
rect 942 1906 948 1907
rect 1038 1911 1044 1912
rect 1038 1907 1039 1911
rect 1043 1907 1044 1911
rect 1134 1911 1140 1912
rect 1038 1906 1044 1907
rect 1106 1907 1112 1908
rect 647 1903 653 1904
rect 647 1899 648 1903
rect 652 1902 653 1903
rect 738 1903 744 1904
rect 652 1900 697 1902
rect 652 1899 653 1900
rect 647 1898 653 1899
rect 738 1899 739 1903
rect 743 1902 744 1903
rect 839 1903 845 1904
rect 743 1900 793 1902
rect 743 1899 744 1900
rect 738 1898 744 1899
rect 839 1899 840 1903
rect 844 1902 845 1903
rect 930 1903 936 1904
rect 844 1900 889 1902
rect 844 1899 845 1900
rect 839 1898 845 1899
rect 930 1899 931 1903
rect 935 1902 936 1903
rect 1031 1903 1037 1904
rect 935 1900 985 1902
rect 935 1899 936 1900
rect 930 1898 936 1899
rect 1031 1899 1032 1903
rect 1036 1902 1037 1903
rect 1106 1903 1107 1907
rect 1111 1906 1112 1907
rect 1134 1907 1135 1911
rect 1139 1907 1140 1911
rect 1134 1906 1140 1907
rect 1230 1911 1236 1912
rect 1230 1907 1231 1911
rect 1235 1907 1236 1911
rect 1230 1906 1236 1907
rect 1326 1911 1332 1912
rect 1326 1907 1327 1911
rect 1331 1907 1332 1911
rect 1326 1906 1332 1907
rect 1422 1911 1428 1912
rect 1422 1907 1423 1911
rect 1427 1907 1428 1911
rect 2006 1908 2007 1912
rect 2011 1908 2012 1912
rect 2006 1907 2012 1908
rect 1422 1906 1428 1907
rect 1111 1904 1126 1906
rect 1111 1903 1112 1904
rect 1106 1902 1112 1903
rect 1124 1902 1126 1904
rect 2330 1903 2336 1904
rect 1036 1900 1081 1902
rect 1124 1900 1177 1902
rect 1036 1899 1037 1900
rect 1031 1898 1037 1899
rect 1306 1899 1312 1900
rect 110 1895 116 1896
rect 110 1891 111 1895
rect 115 1891 116 1895
rect 1306 1895 1307 1899
rect 1311 1895 1312 1899
rect 1306 1894 1312 1895
rect 1402 1899 1408 1900
rect 1402 1895 1403 1899
rect 1407 1895 1408 1899
rect 1402 1894 1408 1895
rect 1498 1899 1504 1900
rect 1498 1895 1499 1899
rect 1503 1895 1504 1899
rect 2307 1899 2313 1900
rect 1498 1894 1504 1895
rect 2006 1895 2012 1896
rect 110 1890 116 1891
rect 654 1892 660 1893
rect 654 1888 655 1892
rect 659 1888 660 1892
rect 654 1887 660 1888
rect 750 1892 756 1893
rect 750 1888 751 1892
rect 755 1888 756 1892
rect 750 1887 756 1888
rect 846 1892 852 1893
rect 846 1888 847 1892
rect 851 1888 852 1892
rect 846 1887 852 1888
rect 942 1892 948 1893
rect 942 1888 943 1892
rect 947 1888 948 1892
rect 942 1887 948 1888
rect 1038 1892 1044 1893
rect 1038 1888 1039 1892
rect 1043 1888 1044 1892
rect 1038 1887 1044 1888
rect 1134 1892 1140 1893
rect 1134 1888 1135 1892
rect 1139 1888 1140 1892
rect 1134 1887 1140 1888
rect 1230 1892 1236 1893
rect 1230 1888 1231 1892
rect 1235 1888 1236 1892
rect 1230 1887 1236 1888
rect 1326 1892 1332 1893
rect 1326 1888 1327 1892
rect 1331 1888 1332 1892
rect 1326 1887 1332 1888
rect 1422 1892 1428 1893
rect 1422 1888 1423 1892
rect 1427 1888 1428 1892
rect 2006 1891 2007 1895
rect 2011 1891 2012 1895
rect 2307 1895 2308 1899
rect 2312 1898 2313 1899
rect 2330 1899 2331 1903
rect 2335 1902 2336 1903
rect 2403 1903 2409 1904
rect 2403 1902 2404 1903
rect 2335 1900 2404 1902
rect 2335 1899 2336 1900
rect 2330 1898 2336 1899
rect 2403 1899 2404 1900
rect 2408 1899 2409 1903
rect 2403 1898 2409 1899
rect 2426 1903 2432 1904
rect 2426 1899 2427 1903
rect 2431 1902 2432 1903
rect 2499 1903 2505 1904
rect 2499 1902 2500 1903
rect 2431 1900 2500 1902
rect 2431 1899 2432 1900
rect 2426 1898 2432 1899
rect 2499 1899 2500 1900
rect 2504 1899 2505 1903
rect 2499 1898 2505 1899
rect 2522 1903 2528 1904
rect 2522 1899 2523 1903
rect 2527 1902 2528 1903
rect 2595 1903 2601 1904
rect 2595 1902 2596 1903
rect 2527 1900 2596 1902
rect 2527 1899 2528 1900
rect 2522 1898 2528 1899
rect 2595 1899 2596 1900
rect 2600 1899 2601 1903
rect 2595 1898 2601 1899
rect 2699 1903 2705 1904
rect 2699 1899 2700 1903
rect 2704 1902 2705 1903
rect 2714 1903 2720 1904
rect 2714 1902 2715 1903
rect 2704 1900 2715 1902
rect 2704 1899 2705 1900
rect 2699 1898 2705 1899
rect 2714 1899 2715 1900
rect 2719 1899 2720 1903
rect 2714 1898 2720 1899
rect 2819 1903 2825 1904
rect 2819 1899 2820 1903
rect 2824 1902 2825 1903
rect 2858 1903 2864 1904
rect 2858 1902 2859 1903
rect 2824 1900 2859 1902
rect 2824 1899 2825 1900
rect 2819 1898 2825 1899
rect 2858 1899 2859 1900
rect 2863 1899 2864 1903
rect 2858 1898 2864 1899
rect 2971 1903 2977 1904
rect 2971 1899 2972 1903
rect 2976 1902 2977 1903
rect 3006 1903 3012 1904
rect 3006 1902 3007 1903
rect 2976 1900 3007 1902
rect 2976 1899 2977 1900
rect 2971 1898 2977 1899
rect 3006 1899 3007 1900
rect 3011 1899 3012 1903
rect 3006 1898 3012 1899
rect 3155 1903 3161 1904
rect 3155 1899 3156 1903
rect 3160 1902 3161 1903
rect 3186 1903 3192 1904
rect 3186 1902 3187 1903
rect 3160 1900 3187 1902
rect 3160 1899 3161 1900
rect 3155 1898 3161 1899
rect 3186 1899 3187 1900
rect 3191 1899 3192 1903
rect 3186 1898 3192 1899
rect 3371 1903 3377 1904
rect 3371 1899 3372 1903
rect 3376 1902 3377 1903
rect 3402 1903 3408 1904
rect 3402 1902 3403 1903
rect 3376 1900 3403 1902
rect 3376 1899 3377 1900
rect 3371 1898 3377 1899
rect 3402 1899 3403 1900
rect 3407 1899 3408 1903
rect 3827 1903 3836 1904
rect 3402 1898 3408 1899
rect 3595 1899 3601 1900
rect 2312 1896 2326 1898
rect 2312 1895 2313 1896
rect 2307 1894 2313 1895
rect 2324 1894 2326 1896
rect 2466 1895 2472 1896
rect 2466 1894 2467 1895
rect 2324 1892 2467 1894
rect 2006 1890 2012 1891
rect 2466 1891 2467 1892
rect 2471 1891 2472 1895
rect 3595 1895 3596 1899
rect 3600 1898 3601 1899
rect 3623 1899 3629 1900
rect 3623 1898 3624 1899
rect 3600 1896 3624 1898
rect 3600 1895 3601 1896
rect 3595 1894 3601 1895
rect 3623 1895 3624 1896
rect 3628 1895 3629 1899
rect 3827 1899 3828 1903
rect 3835 1899 3836 1903
rect 3827 1898 3836 1899
rect 3623 1894 3629 1895
rect 2466 1890 2472 1891
rect 1422 1887 1428 1888
rect 1306 1875 1312 1876
rect 707 1871 713 1872
rect 707 1867 708 1871
rect 712 1870 713 1871
rect 738 1871 744 1872
rect 738 1870 739 1871
rect 712 1868 739 1870
rect 712 1867 713 1868
rect 707 1866 713 1867
rect 738 1867 739 1868
rect 743 1867 744 1871
rect 738 1866 744 1867
rect 803 1871 809 1872
rect 803 1867 804 1871
rect 808 1870 809 1871
rect 839 1871 845 1872
rect 839 1870 840 1871
rect 808 1868 840 1870
rect 808 1867 809 1868
rect 803 1866 809 1867
rect 839 1867 840 1868
rect 844 1867 845 1871
rect 839 1866 845 1867
rect 899 1871 905 1872
rect 899 1867 900 1871
rect 904 1870 905 1871
rect 930 1871 936 1872
rect 930 1870 931 1871
rect 904 1868 931 1870
rect 904 1867 905 1868
rect 899 1866 905 1867
rect 930 1867 931 1868
rect 935 1867 936 1871
rect 930 1866 936 1867
rect 995 1871 1001 1872
rect 995 1867 996 1871
rect 1000 1870 1001 1871
rect 1031 1871 1037 1872
rect 1031 1870 1032 1871
rect 1000 1868 1032 1870
rect 1000 1867 1001 1868
rect 995 1866 1001 1867
rect 1031 1867 1032 1868
rect 1036 1867 1037 1871
rect 1031 1866 1037 1867
rect 1091 1871 1097 1872
rect 1091 1867 1092 1871
rect 1096 1870 1097 1871
rect 1122 1871 1128 1872
rect 1122 1870 1123 1871
rect 1096 1868 1123 1870
rect 1096 1867 1097 1868
rect 1091 1866 1097 1867
rect 1122 1867 1123 1868
rect 1127 1867 1128 1871
rect 1122 1866 1128 1867
rect 1187 1871 1193 1872
rect 1187 1867 1188 1871
rect 1192 1870 1193 1871
rect 1202 1871 1208 1872
rect 1202 1870 1203 1871
rect 1192 1868 1203 1870
rect 1192 1867 1193 1868
rect 1187 1866 1193 1867
rect 1202 1867 1203 1868
rect 1207 1867 1208 1871
rect 1306 1871 1307 1875
rect 1311 1874 1312 1875
rect 2202 1875 2208 1876
rect 1311 1872 1346 1874
rect 1311 1871 1312 1872
rect 1306 1870 1312 1871
rect 1344 1870 1346 1872
rect 1379 1871 1385 1872
rect 1379 1870 1380 1871
rect 1344 1868 1380 1870
rect 1202 1866 1208 1867
rect 1283 1867 1289 1868
rect 1283 1863 1284 1867
rect 1288 1866 1289 1867
rect 1334 1867 1340 1868
rect 1334 1866 1335 1867
rect 1288 1864 1335 1866
rect 1288 1863 1289 1864
rect 1283 1862 1289 1863
rect 1334 1863 1335 1864
rect 1339 1863 1340 1867
rect 1379 1867 1380 1868
rect 1384 1867 1385 1871
rect 1379 1866 1385 1867
rect 1402 1871 1408 1872
rect 1402 1867 1403 1871
rect 1407 1870 1408 1871
rect 1475 1871 1481 1872
rect 1475 1870 1476 1871
rect 1407 1868 1476 1870
rect 1407 1867 1408 1868
rect 1402 1866 1408 1867
rect 1475 1867 1476 1868
rect 1480 1867 1481 1871
rect 2202 1871 2203 1875
rect 2207 1874 2208 1875
rect 2235 1875 2241 1876
rect 2235 1874 2236 1875
rect 2207 1872 2236 1874
rect 2207 1871 2208 1872
rect 2202 1870 2208 1871
rect 2235 1871 2236 1872
rect 2240 1871 2241 1875
rect 2235 1870 2241 1871
rect 2271 1875 2277 1876
rect 2271 1871 2272 1875
rect 2276 1874 2277 1875
rect 2331 1875 2337 1876
rect 2331 1874 2332 1875
rect 2276 1872 2332 1874
rect 2276 1871 2277 1872
rect 2271 1870 2277 1871
rect 2331 1871 2332 1872
rect 2336 1871 2337 1875
rect 2331 1870 2337 1871
rect 2375 1875 2381 1876
rect 2375 1871 2376 1875
rect 2380 1874 2381 1875
rect 2435 1875 2441 1876
rect 2435 1874 2436 1875
rect 2380 1872 2436 1874
rect 2380 1871 2381 1872
rect 2375 1870 2381 1871
rect 2435 1871 2436 1872
rect 2440 1871 2441 1875
rect 2435 1870 2441 1871
rect 2458 1875 2464 1876
rect 2458 1871 2459 1875
rect 2463 1874 2464 1875
rect 2539 1875 2545 1876
rect 2539 1874 2540 1875
rect 2463 1872 2540 1874
rect 2463 1871 2464 1872
rect 2458 1870 2464 1871
rect 2539 1871 2540 1872
rect 2544 1871 2545 1875
rect 2539 1870 2545 1871
rect 2638 1875 2649 1876
rect 2638 1871 2639 1875
rect 2643 1871 2644 1875
rect 2648 1871 2649 1875
rect 2638 1870 2649 1871
rect 2666 1875 2672 1876
rect 2666 1871 2667 1875
rect 2671 1874 2672 1875
rect 2755 1875 2761 1876
rect 2755 1874 2756 1875
rect 2671 1872 2756 1874
rect 2671 1871 2672 1872
rect 2666 1870 2672 1871
rect 2755 1871 2756 1872
rect 2760 1871 2761 1875
rect 2755 1870 2761 1871
rect 2870 1875 2876 1876
rect 2870 1871 2871 1875
rect 2875 1874 2876 1875
rect 2883 1875 2889 1876
rect 2883 1874 2884 1875
rect 2875 1872 2884 1874
rect 2875 1871 2876 1872
rect 2870 1870 2876 1871
rect 2883 1871 2884 1872
rect 2888 1871 2889 1875
rect 2883 1870 2889 1871
rect 2906 1875 2912 1876
rect 2906 1871 2907 1875
rect 2911 1874 2912 1875
rect 3043 1875 3049 1876
rect 3043 1874 3044 1875
rect 2911 1872 3044 1874
rect 2911 1871 2912 1872
rect 2906 1870 2912 1871
rect 3043 1871 3044 1872
rect 3048 1871 3049 1875
rect 3043 1870 3049 1871
rect 3066 1875 3072 1876
rect 3066 1871 3067 1875
rect 3071 1874 3072 1875
rect 3235 1875 3241 1876
rect 3235 1874 3236 1875
rect 3071 1872 3236 1874
rect 3071 1871 3072 1872
rect 3066 1870 3072 1871
rect 3235 1871 3236 1872
rect 3240 1871 3241 1875
rect 3235 1870 3241 1871
rect 3258 1875 3264 1876
rect 3258 1871 3259 1875
rect 3263 1874 3264 1875
rect 3451 1875 3457 1876
rect 3451 1874 3452 1875
rect 3263 1872 3452 1874
rect 3263 1871 3264 1872
rect 3258 1870 3264 1871
rect 3451 1871 3452 1872
rect 3456 1871 3457 1875
rect 3451 1870 3457 1871
rect 3474 1875 3480 1876
rect 3474 1871 3475 1875
rect 3479 1874 3480 1875
rect 3683 1875 3689 1876
rect 3683 1874 3684 1875
rect 3479 1872 3684 1874
rect 3479 1871 3480 1872
rect 3474 1870 3480 1871
rect 3683 1871 3684 1872
rect 3688 1871 3689 1875
rect 3683 1870 3689 1871
rect 3891 1875 3897 1876
rect 3891 1871 3892 1875
rect 3896 1874 3897 1875
rect 3906 1875 3912 1876
rect 3906 1874 3907 1875
rect 3896 1872 3907 1874
rect 3896 1871 3897 1872
rect 3891 1870 3897 1871
rect 3906 1871 3907 1872
rect 3911 1871 3912 1875
rect 3906 1870 3912 1871
rect 1475 1866 1481 1867
rect 1334 1862 1340 1863
rect 330 1855 336 1856
rect 330 1851 331 1855
rect 335 1854 336 1855
rect 371 1855 377 1856
rect 371 1854 372 1855
rect 335 1852 372 1854
rect 335 1851 336 1852
rect 330 1850 336 1851
rect 371 1851 372 1852
rect 376 1851 377 1855
rect 371 1850 377 1851
rect 394 1855 400 1856
rect 394 1851 395 1855
rect 399 1854 400 1855
rect 499 1855 505 1856
rect 499 1854 500 1855
rect 399 1852 500 1854
rect 399 1851 400 1852
rect 394 1850 400 1851
rect 499 1851 500 1852
rect 504 1851 505 1855
rect 499 1850 505 1851
rect 635 1855 641 1856
rect 635 1851 636 1855
rect 640 1854 641 1855
rect 647 1855 653 1856
rect 647 1854 648 1855
rect 640 1852 648 1854
rect 640 1851 641 1852
rect 635 1850 641 1851
rect 647 1851 648 1852
rect 652 1851 653 1855
rect 647 1850 653 1851
rect 695 1855 701 1856
rect 695 1851 696 1855
rect 700 1854 701 1855
rect 771 1855 777 1856
rect 771 1854 772 1855
rect 700 1852 772 1854
rect 700 1851 701 1852
rect 695 1850 701 1851
rect 771 1851 772 1852
rect 776 1851 777 1855
rect 771 1850 777 1851
rect 794 1855 800 1856
rect 794 1851 795 1855
rect 799 1854 800 1855
rect 907 1855 913 1856
rect 907 1854 908 1855
rect 799 1852 908 1854
rect 799 1851 800 1852
rect 794 1850 800 1851
rect 907 1851 908 1852
rect 912 1851 913 1855
rect 1066 1855 1072 1856
rect 907 1850 913 1851
rect 1043 1853 1049 1854
rect 1043 1849 1044 1853
rect 1048 1849 1049 1853
rect 1066 1851 1067 1855
rect 1071 1854 1072 1855
rect 1179 1855 1185 1856
rect 1179 1854 1180 1855
rect 1071 1852 1180 1854
rect 1071 1851 1072 1852
rect 1066 1850 1072 1851
rect 1179 1851 1180 1852
rect 1184 1851 1185 1855
rect 1179 1850 1185 1851
rect 1202 1855 1208 1856
rect 1202 1851 1203 1855
rect 1207 1854 1208 1855
rect 1315 1855 1321 1856
rect 1315 1854 1316 1855
rect 1207 1852 1316 1854
rect 1207 1851 1208 1852
rect 1202 1850 1208 1851
rect 1315 1851 1316 1852
rect 1320 1851 1321 1855
rect 1315 1850 1321 1851
rect 1451 1855 1457 1856
rect 1451 1851 1452 1855
rect 1456 1854 1457 1855
rect 1482 1855 1488 1856
rect 1482 1854 1483 1855
rect 1456 1852 1483 1854
rect 1456 1851 1457 1852
rect 1451 1850 1457 1851
rect 1482 1851 1483 1852
rect 1487 1851 1488 1855
rect 1482 1850 1488 1851
rect 1498 1855 1504 1856
rect 1498 1851 1499 1855
rect 1503 1854 1504 1855
rect 1587 1855 1593 1856
rect 1587 1854 1588 1855
rect 1503 1852 1588 1854
rect 1503 1851 1504 1852
rect 1498 1850 1504 1851
rect 1587 1851 1588 1852
rect 1592 1851 1593 1855
rect 1587 1850 1593 1851
rect 2182 1852 2188 1853
rect 1043 1848 1049 1849
rect 2046 1849 2052 1850
rect 1044 1846 1046 1848
rect 1170 1847 1176 1848
rect 1170 1846 1171 1847
rect 1044 1844 1171 1846
rect 1170 1843 1171 1844
rect 1175 1843 1176 1847
rect 2046 1845 2047 1849
rect 2051 1845 2052 1849
rect 2182 1848 2183 1852
rect 2187 1848 2188 1852
rect 2182 1847 2188 1848
rect 2278 1852 2284 1853
rect 2278 1848 2279 1852
rect 2283 1848 2284 1852
rect 2278 1847 2284 1848
rect 2382 1852 2388 1853
rect 2382 1848 2383 1852
rect 2387 1848 2388 1852
rect 2382 1847 2388 1848
rect 2486 1852 2492 1853
rect 2486 1848 2487 1852
rect 2491 1848 2492 1852
rect 2486 1847 2492 1848
rect 2590 1852 2596 1853
rect 2590 1848 2591 1852
rect 2595 1848 2596 1852
rect 2590 1847 2596 1848
rect 2702 1852 2708 1853
rect 2702 1848 2703 1852
rect 2707 1848 2708 1852
rect 2702 1847 2708 1848
rect 2830 1852 2836 1853
rect 2830 1848 2831 1852
rect 2835 1848 2836 1852
rect 2830 1847 2836 1848
rect 2990 1852 2996 1853
rect 2990 1848 2991 1852
rect 2995 1848 2996 1852
rect 2990 1847 2996 1848
rect 3182 1852 3188 1853
rect 3182 1848 3183 1852
rect 3187 1848 3188 1852
rect 3182 1847 3188 1848
rect 3398 1852 3404 1853
rect 3398 1848 3399 1852
rect 3403 1848 3404 1852
rect 3398 1847 3404 1848
rect 3630 1852 3636 1853
rect 3630 1848 3631 1852
rect 3635 1848 3636 1852
rect 3630 1847 3636 1848
rect 3838 1852 3844 1853
rect 3838 1848 3839 1852
rect 3843 1848 3844 1852
rect 3838 1847 3844 1848
rect 3942 1849 3948 1850
rect 2046 1844 2052 1845
rect 3942 1845 3943 1849
rect 3947 1845 3948 1849
rect 3942 1844 3948 1845
rect 1170 1842 1176 1843
rect 2271 1843 2277 1844
rect 2271 1842 2272 1843
rect 2261 1840 2272 1842
rect 2271 1839 2272 1840
rect 2276 1839 2277 1843
rect 2375 1843 2381 1844
rect 2375 1842 2376 1843
rect 2357 1840 2376 1842
rect 2271 1838 2277 1839
rect 2375 1839 2376 1840
rect 2380 1839 2381 1843
rect 2375 1838 2381 1839
rect 2458 1843 2464 1844
rect 2458 1839 2459 1843
rect 2463 1839 2464 1843
rect 2458 1838 2464 1839
rect 2466 1843 2472 1844
rect 2466 1839 2467 1843
rect 2471 1842 2472 1843
rect 2666 1843 2672 1844
rect 2471 1840 2529 1842
rect 2471 1839 2472 1840
rect 2466 1838 2472 1839
rect 2666 1839 2667 1843
rect 2671 1839 2672 1843
rect 2666 1838 2672 1839
rect 2770 1843 2776 1844
rect 2770 1839 2771 1843
rect 2775 1839 2776 1843
rect 2770 1838 2776 1839
rect 2906 1843 2912 1844
rect 2906 1839 2907 1843
rect 2911 1839 2912 1843
rect 2906 1838 2912 1839
rect 3066 1843 3072 1844
rect 3066 1839 3067 1843
rect 3071 1839 3072 1843
rect 3066 1838 3072 1839
rect 3258 1843 3264 1844
rect 3258 1839 3259 1843
rect 3263 1839 3264 1843
rect 3258 1838 3264 1839
rect 3474 1843 3480 1844
rect 3474 1839 3475 1843
rect 3479 1839 3480 1843
rect 3474 1838 3480 1839
rect 3623 1843 3629 1844
rect 3623 1839 3624 1843
rect 3628 1842 3629 1843
rect 3914 1843 3920 1844
rect 3628 1840 3673 1842
rect 3628 1839 3629 1840
rect 3623 1838 3629 1839
rect 3914 1839 3915 1843
rect 3919 1839 3920 1843
rect 3914 1838 3920 1839
rect 2182 1833 2188 1834
rect 318 1832 324 1833
rect 110 1829 116 1830
rect 110 1825 111 1829
rect 115 1825 116 1829
rect 318 1828 319 1832
rect 323 1828 324 1832
rect 318 1827 324 1828
rect 446 1832 452 1833
rect 446 1828 447 1832
rect 451 1828 452 1832
rect 446 1827 452 1828
rect 582 1832 588 1833
rect 582 1828 583 1832
rect 587 1828 588 1832
rect 582 1827 588 1828
rect 718 1832 724 1833
rect 718 1828 719 1832
rect 723 1828 724 1832
rect 718 1827 724 1828
rect 854 1832 860 1833
rect 854 1828 855 1832
rect 859 1828 860 1832
rect 854 1827 860 1828
rect 990 1832 996 1833
rect 990 1828 991 1832
rect 995 1828 996 1832
rect 990 1827 996 1828
rect 1126 1832 1132 1833
rect 1126 1828 1127 1832
rect 1131 1828 1132 1832
rect 1126 1827 1132 1828
rect 1262 1832 1268 1833
rect 1262 1828 1263 1832
rect 1267 1828 1268 1832
rect 1262 1827 1268 1828
rect 1398 1832 1404 1833
rect 1398 1828 1399 1832
rect 1403 1828 1404 1832
rect 1398 1827 1404 1828
rect 1534 1832 1540 1833
rect 1534 1828 1535 1832
rect 1539 1828 1540 1832
rect 2046 1832 2052 1833
rect 1534 1827 1540 1828
rect 2006 1829 2012 1830
rect 110 1824 116 1825
rect 2006 1825 2007 1829
rect 2011 1825 2012 1829
rect 2046 1828 2047 1832
rect 2051 1828 2052 1832
rect 2182 1829 2183 1833
rect 2187 1829 2188 1833
rect 2182 1828 2188 1829
rect 2278 1833 2284 1834
rect 2278 1829 2279 1833
rect 2283 1829 2284 1833
rect 2278 1828 2284 1829
rect 2382 1833 2388 1834
rect 2382 1829 2383 1833
rect 2387 1829 2388 1833
rect 2382 1828 2388 1829
rect 2486 1833 2492 1834
rect 2486 1829 2487 1833
rect 2491 1829 2492 1833
rect 2486 1828 2492 1829
rect 2590 1833 2596 1834
rect 2590 1829 2591 1833
rect 2595 1829 2596 1833
rect 2590 1828 2596 1829
rect 2702 1833 2708 1834
rect 2702 1829 2703 1833
rect 2707 1829 2708 1833
rect 2702 1828 2708 1829
rect 2830 1833 2836 1834
rect 2830 1829 2831 1833
rect 2835 1829 2836 1833
rect 2830 1828 2836 1829
rect 2990 1833 2996 1834
rect 2990 1829 2991 1833
rect 2995 1829 2996 1833
rect 2990 1828 2996 1829
rect 3182 1833 3188 1834
rect 3182 1829 3183 1833
rect 3187 1829 3188 1833
rect 3182 1828 3188 1829
rect 3398 1833 3404 1834
rect 3398 1829 3399 1833
rect 3403 1829 3404 1833
rect 3398 1828 3404 1829
rect 3630 1833 3636 1834
rect 3630 1829 3631 1833
rect 3635 1829 3636 1833
rect 3630 1828 3636 1829
rect 3838 1833 3844 1834
rect 3838 1829 3839 1833
rect 3843 1829 3844 1833
rect 3838 1828 3844 1829
rect 3942 1832 3948 1833
rect 3942 1828 3943 1832
rect 3947 1828 3948 1832
rect 2046 1827 2052 1828
rect 3942 1827 3948 1828
rect 2006 1824 2012 1825
rect 394 1823 400 1824
rect 394 1819 395 1823
rect 399 1819 400 1823
rect 394 1818 400 1819
rect 514 1823 520 1824
rect 514 1819 515 1823
rect 519 1819 520 1823
rect 695 1823 701 1824
rect 695 1822 696 1823
rect 661 1820 696 1822
rect 514 1818 520 1819
rect 695 1819 696 1820
rect 700 1819 701 1823
rect 695 1818 701 1819
rect 794 1823 800 1824
rect 794 1819 795 1823
rect 799 1819 800 1823
rect 794 1818 800 1819
rect 922 1823 928 1824
rect 922 1819 923 1823
rect 927 1819 928 1823
rect 922 1818 928 1819
rect 1066 1823 1072 1824
rect 1066 1819 1067 1823
rect 1071 1819 1072 1823
rect 1066 1818 1072 1819
rect 1202 1823 1208 1824
rect 1202 1819 1203 1823
rect 1207 1819 1208 1823
rect 1202 1818 1208 1819
rect 1334 1823 1340 1824
rect 1334 1819 1335 1823
rect 1339 1819 1340 1823
rect 1334 1818 1340 1819
rect 1466 1823 1472 1824
rect 1466 1819 1467 1823
rect 1471 1819 1472 1823
rect 1466 1818 1472 1819
rect 1482 1823 1488 1824
rect 1482 1819 1483 1823
rect 1487 1822 1488 1823
rect 1487 1820 1577 1822
rect 1487 1819 1488 1820
rect 1482 1818 1488 1819
rect 318 1813 324 1814
rect 110 1812 116 1813
rect 110 1808 111 1812
rect 115 1808 116 1812
rect 318 1809 319 1813
rect 323 1809 324 1813
rect 318 1808 324 1809
rect 446 1813 452 1814
rect 446 1809 447 1813
rect 451 1809 452 1813
rect 446 1808 452 1809
rect 582 1813 588 1814
rect 582 1809 583 1813
rect 587 1809 588 1813
rect 582 1808 588 1809
rect 718 1813 724 1814
rect 718 1809 719 1813
rect 723 1809 724 1813
rect 718 1808 724 1809
rect 854 1813 860 1814
rect 854 1809 855 1813
rect 859 1809 860 1813
rect 854 1808 860 1809
rect 990 1813 996 1814
rect 990 1809 991 1813
rect 995 1809 996 1813
rect 990 1808 996 1809
rect 1126 1813 1132 1814
rect 1126 1809 1127 1813
rect 1131 1809 1132 1813
rect 1126 1808 1132 1809
rect 1262 1813 1268 1814
rect 1262 1809 1263 1813
rect 1267 1809 1268 1813
rect 1262 1808 1268 1809
rect 1398 1813 1404 1814
rect 1398 1809 1399 1813
rect 1403 1809 1404 1813
rect 1398 1808 1404 1809
rect 1534 1813 1540 1814
rect 1534 1809 1535 1813
rect 1539 1809 1540 1813
rect 1534 1808 1540 1809
rect 2006 1812 2012 1813
rect 2006 1808 2007 1812
rect 2011 1808 2012 1812
rect 110 1807 116 1808
rect 2006 1807 2012 1808
rect 2046 1776 2052 1777
rect 3942 1776 3948 1777
rect 2046 1772 2047 1776
rect 2051 1772 2052 1776
rect 2046 1771 2052 1772
rect 2126 1775 2132 1776
rect 2126 1771 2127 1775
rect 2131 1771 2132 1775
rect 2126 1770 2132 1771
rect 2310 1775 2316 1776
rect 2310 1771 2311 1775
rect 2315 1771 2316 1775
rect 2310 1770 2316 1771
rect 2494 1775 2500 1776
rect 2494 1771 2495 1775
rect 2499 1771 2500 1775
rect 2494 1770 2500 1771
rect 2686 1775 2692 1776
rect 2686 1771 2687 1775
rect 2691 1771 2692 1775
rect 2686 1770 2692 1771
rect 2878 1775 2884 1776
rect 2878 1771 2879 1775
rect 2883 1771 2884 1775
rect 2878 1770 2884 1771
rect 3070 1775 3076 1776
rect 3070 1771 3071 1775
rect 3075 1771 3076 1775
rect 3070 1770 3076 1771
rect 3262 1775 3268 1776
rect 3262 1771 3263 1775
rect 3267 1771 3268 1775
rect 3262 1770 3268 1771
rect 3462 1775 3468 1776
rect 3462 1771 3463 1775
rect 3467 1771 3468 1775
rect 3462 1770 3468 1771
rect 3662 1775 3668 1776
rect 3662 1771 3663 1775
rect 3667 1771 3668 1775
rect 3662 1770 3668 1771
rect 3838 1775 3844 1776
rect 3838 1771 3839 1775
rect 3843 1771 3844 1775
rect 3942 1772 3943 1776
rect 3947 1772 3948 1776
rect 3838 1770 3844 1771
rect 3906 1771 3912 1772
rect 3942 1771 3948 1772
rect 2202 1767 2208 1768
rect 2202 1763 2203 1767
rect 2207 1763 2208 1767
rect 2202 1762 2208 1763
rect 2215 1767 2221 1768
rect 2215 1763 2216 1767
rect 2220 1766 2221 1767
rect 2399 1767 2405 1768
rect 2220 1764 2353 1766
rect 2220 1763 2221 1764
rect 2215 1762 2221 1763
rect 2399 1763 2400 1767
rect 2404 1766 2405 1767
rect 2870 1767 2876 1768
rect 2404 1764 2537 1766
rect 2404 1763 2405 1764
rect 2399 1762 2405 1763
rect 2798 1763 2804 1764
rect 2798 1762 2799 1763
rect 2765 1760 2799 1762
rect 2046 1759 2052 1760
rect 110 1756 116 1757
rect 2006 1756 2012 1757
rect 110 1752 111 1756
rect 115 1752 116 1756
rect 110 1751 116 1752
rect 254 1755 260 1756
rect 254 1751 255 1755
rect 259 1751 260 1755
rect 254 1750 260 1751
rect 390 1755 396 1756
rect 390 1751 391 1755
rect 395 1751 396 1755
rect 390 1750 396 1751
rect 534 1755 540 1756
rect 534 1751 535 1755
rect 539 1751 540 1755
rect 534 1750 540 1751
rect 694 1755 700 1756
rect 694 1751 695 1755
rect 699 1751 700 1755
rect 694 1750 700 1751
rect 862 1755 868 1756
rect 862 1751 863 1755
rect 867 1751 868 1755
rect 862 1750 868 1751
rect 1030 1755 1036 1756
rect 1030 1751 1031 1755
rect 1035 1751 1036 1755
rect 1030 1750 1036 1751
rect 1206 1755 1212 1756
rect 1206 1751 1207 1755
rect 1211 1751 1212 1755
rect 1206 1750 1212 1751
rect 1382 1755 1388 1756
rect 1382 1751 1383 1755
rect 1387 1751 1388 1755
rect 1382 1750 1388 1751
rect 1558 1755 1564 1756
rect 1558 1751 1559 1755
rect 1563 1751 1564 1755
rect 1558 1750 1564 1751
rect 1742 1755 1748 1756
rect 1742 1751 1743 1755
rect 1747 1751 1748 1755
rect 2006 1752 2007 1756
rect 2011 1752 2012 1756
rect 2046 1755 2047 1759
rect 2051 1755 2052 1759
rect 2798 1759 2799 1760
rect 2803 1759 2804 1763
rect 2870 1763 2871 1767
rect 2875 1766 2876 1767
rect 2967 1767 2973 1768
rect 2875 1764 2921 1766
rect 2875 1763 2876 1764
rect 2870 1762 2876 1763
rect 2967 1763 2968 1767
rect 2972 1766 2973 1767
rect 3158 1767 3164 1768
rect 2972 1764 3113 1766
rect 2972 1763 2973 1764
rect 2967 1762 2973 1763
rect 3158 1763 3159 1767
rect 3163 1766 3164 1767
rect 3346 1767 3352 1768
rect 3163 1764 3305 1766
rect 3163 1763 3164 1764
rect 3158 1762 3164 1763
rect 3346 1763 3347 1767
rect 3351 1766 3352 1767
rect 3906 1767 3907 1771
rect 3911 1770 3912 1771
rect 3911 1768 3918 1770
rect 3911 1767 3912 1768
rect 3906 1766 3912 1767
rect 3351 1764 3505 1766
rect 3916 1765 3918 1768
rect 3351 1763 3352 1764
rect 3346 1762 3352 1763
rect 3738 1763 3744 1764
rect 2798 1758 2804 1759
rect 3738 1759 3739 1763
rect 3743 1759 3744 1763
rect 3738 1758 3744 1759
rect 3942 1759 3948 1760
rect 2046 1754 2052 1755
rect 2126 1756 2132 1757
rect 2006 1751 2012 1752
rect 2126 1752 2127 1756
rect 2131 1752 2132 1756
rect 2126 1751 2132 1752
rect 2310 1756 2316 1757
rect 2310 1752 2311 1756
rect 2315 1752 2316 1756
rect 2310 1751 2316 1752
rect 2494 1756 2500 1757
rect 2494 1752 2495 1756
rect 2499 1752 2500 1756
rect 2494 1751 2500 1752
rect 2686 1756 2692 1757
rect 2686 1752 2687 1756
rect 2691 1752 2692 1756
rect 2686 1751 2692 1752
rect 2878 1756 2884 1757
rect 2878 1752 2879 1756
rect 2883 1752 2884 1756
rect 2878 1751 2884 1752
rect 3070 1756 3076 1757
rect 3070 1752 3071 1756
rect 3075 1752 3076 1756
rect 3070 1751 3076 1752
rect 3262 1756 3268 1757
rect 3262 1752 3263 1756
rect 3267 1752 3268 1756
rect 3262 1751 3268 1752
rect 3462 1756 3468 1757
rect 3462 1752 3463 1756
rect 3467 1752 3468 1756
rect 3462 1751 3468 1752
rect 3662 1756 3668 1757
rect 3662 1752 3663 1756
rect 3667 1752 3668 1756
rect 3662 1751 3668 1752
rect 3838 1756 3844 1757
rect 3838 1752 3839 1756
rect 3843 1752 3844 1756
rect 3942 1755 3943 1759
rect 3947 1755 3948 1759
rect 3942 1754 3948 1755
rect 3838 1751 3844 1752
rect 1742 1750 1748 1751
rect 330 1747 336 1748
rect 330 1743 331 1747
rect 335 1743 336 1747
rect 330 1742 336 1743
rect 342 1747 348 1748
rect 342 1743 343 1747
rect 347 1746 348 1747
rect 662 1747 668 1748
rect 347 1744 433 1746
rect 347 1743 348 1744
rect 342 1742 348 1743
rect 618 1743 624 1744
rect 618 1742 619 1743
rect 613 1740 619 1742
rect 110 1739 116 1740
rect 110 1735 111 1739
rect 115 1735 116 1739
rect 618 1739 619 1740
rect 623 1739 624 1743
rect 662 1743 663 1747
rect 667 1746 668 1747
rect 814 1747 820 1748
rect 667 1744 737 1746
rect 667 1743 668 1744
rect 662 1742 668 1743
rect 814 1743 815 1747
rect 819 1746 820 1747
rect 1170 1747 1176 1748
rect 819 1744 905 1746
rect 819 1743 820 1744
rect 814 1742 820 1743
rect 1106 1743 1112 1744
rect 618 1738 624 1739
rect 1106 1739 1107 1743
rect 1111 1739 1112 1743
rect 1170 1743 1171 1747
rect 1175 1746 1176 1747
rect 1175 1744 1249 1746
rect 1175 1743 1176 1744
rect 1170 1742 1176 1743
rect 1518 1743 1524 1744
rect 1518 1742 1519 1743
rect 1461 1740 1519 1742
rect 1106 1738 1112 1739
rect 1518 1739 1519 1740
rect 1523 1739 1524 1743
rect 1518 1738 1524 1739
rect 1634 1743 1640 1744
rect 1634 1739 1635 1743
rect 1639 1739 1640 1743
rect 1634 1738 1640 1739
rect 1818 1743 1824 1744
rect 1818 1739 1819 1743
rect 1823 1739 1824 1743
rect 1818 1738 1824 1739
rect 2006 1739 2012 1740
rect 110 1734 116 1735
rect 254 1736 260 1737
rect 254 1732 255 1736
rect 259 1732 260 1736
rect 254 1731 260 1732
rect 390 1736 396 1737
rect 390 1732 391 1736
rect 395 1732 396 1736
rect 390 1731 396 1732
rect 534 1736 540 1737
rect 534 1732 535 1736
rect 539 1732 540 1736
rect 534 1731 540 1732
rect 694 1736 700 1737
rect 694 1732 695 1736
rect 699 1732 700 1736
rect 694 1731 700 1732
rect 862 1736 868 1737
rect 862 1732 863 1736
rect 867 1732 868 1736
rect 862 1731 868 1732
rect 1030 1736 1036 1737
rect 1030 1732 1031 1736
rect 1035 1732 1036 1736
rect 1030 1731 1036 1732
rect 1206 1736 1212 1737
rect 1206 1732 1207 1736
rect 1211 1732 1212 1736
rect 1206 1731 1212 1732
rect 1382 1736 1388 1737
rect 1382 1732 1383 1736
rect 1387 1732 1388 1736
rect 1382 1731 1388 1732
rect 1558 1736 1564 1737
rect 1558 1732 1559 1736
rect 1563 1732 1564 1736
rect 1558 1731 1564 1732
rect 1742 1736 1748 1737
rect 1742 1732 1743 1736
rect 1747 1732 1748 1736
rect 2006 1735 2007 1739
rect 2011 1735 2012 1739
rect 2006 1734 2012 1735
rect 2179 1735 2185 1736
rect 1742 1731 1748 1732
rect 2179 1731 2180 1735
rect 2184 1734 2185 1735
rect 2215 1735 2221 1736
rect 2215 1734 2216 1735
rect 2184 1732 2216 1734
rect 2184 1731 2185 1732
rect 2179 1730 2185 1731
rect 2215 1731 2216 1732
rect 2220 1731 2221 1735
rect 2215 1730 2221 1731
rect 2363 1735 2369 1736
rect 2363 1731 2364 1735
rect 2368 1734 2369 1735
rect 2399 1735 2405 1736
rect 2399 1734 2400 1735
rect 2368 1732 2400 1734
rect 2368 1731 2369 1732
rect 2363 1730 2369 1731
rect 2399 1731 2400 1732
rect 2404 1731 2405 1735
rect 2739 1735 2745 1736
rect 2399 1730 2405 1731
rect 2547 1731 2553 1732
rect 2547 1727 2548 1731
rect 2552 1730 2553 1731
rect 2578 1731 2584 1732
rect 2578 1730 2579 1731
rect 2552 1728 2579 1730
rect 2552 1727 2553 1728
rect 2547 1726 2553 1727
rect 2578 1727 2579 1728
rect 2583 1727 2584 1731
rect 2739 1731 2740 1735
rect 2744 1734 2745 1735
rect 2770 1735 2776 1736
rect 2770 1734 2771 1735
rect 2744 1732 2771 1734
rect 2744 1731 2745 1732
rect 2739 1730 2745 1731
rect 2770 1731 2771 1732
rect 2775 1731 2776 1735
rect 2770 1730 2776 1731
rect 2931 1735 2937 1736
rect 2931 1731 2932 1735
rect 2936 1734 2937 1735
rect 2967 1735 2973 1736
rect 2967 1734 2968 1735
rect 2936 1732 2968 1734
rect 2936 1731 2937 1732
rect 2931 1730 2937 1731
rect 2967 1731 2968 1732
rect 2972 1731 2973 1735
rect 2967 1730 2973 1731
rect 3123 1735 3129 1736
rect 3123 1731 3124 1735
rect 3128 1734 3129 1735
rect 3158 1735 3164 1736
rect 3158 1734 3159 1735
rect 3128 1732 3159 1734
rect 3128 1731 3129 1732
rect 3123 1730 3129 1731
rect 3158 1731 3159 1732
rect 3163 1731 3164 1735
rect 3158 1730 3164 1731
rect 3315 1735 3321 1736
rect 3315 1731 3316 1735
rect 3320 1734 3321 1735
rect 3346 1735 3352 1736
rect 3346 1734 3347 1735
rect 3320 1732 3347 1734
rect 3320 1731 3321 1732
rect 3315 1730 3321 1731
rect 3346 1731 3347 1732
rect 3351 1731 3352 1735
rect 3715 1735 3721 1736
rect 3346 1730 3352 1731
rect 3514 1731 3521 1732
rect 2578 1726 2584 1727
rect 3514 1727 3515 1731
rect 3520 1727 3521 1731
rect 3715 1731 3716 1735
rect 3720 1734 3721 1735
rect 3750 1735 3756 1736
rect 3750 1734 3751 1735
rect 3720 1732 3751 1734
rect 3720 1731 3721 1732
rect 3715 1730 3721 1731
rect 3750 1731 3751 1732
rect 3755 1731 3756 1735
rect 3750 1730 3756 1731
rect 3891 1731 3897 1732
rect 3514 1726 3521 1727
rect 3891 1727 3892 1731
rect 3896 1730 3897 1731
rect 3906 1731 3912 1732
rect 3906 1730 3907 1731
rect 3896 1728 3907 1730
rect 3896 1727 3897 1728
rect 3891 1726 3897 1727
rect 3906 1727 3907 1728
rect 3911 1727 3912 1731
rect 3906 1726 3912 1727
rect 307 1715 313 1716
rect 307 1711 308 1715
rect 312 1714 313 1715
rect 342 1715 348 1716
rect 342 1714 343 1715
rect 312 1712 343 1714
rect 312 1711 313 1712
rect 307 1710 313 1711
rect 342 1711 343 1712
rect 347 1711 348 1715
rect 587 1715 593 1716
rect 342 1710 348 1711
rect 443 1711 449 1712
rect 443 1707 444 1711
rect 448 1710 449 1711
rect 498 1711 504 1712
rect 498 1710 499 1711
rect 448 1708 499 1710
rect 448 1707 449 1708
rect 443 1706 449 1707
rect 498 1707 499 1708
rect 503 1707 504 1711
rect 587 1711 588 1715
rect 592 1714 593 1715
rect 662 1715 668 1716
rect 662 1714 663 1715
rect 592 1712 663 1714
rect 592 1711 593 1712
rect 587 1710 593 1711
rect 662 1711 663 1712
rect 667 1711 668 1715
rect 662 1710 668 1711
rect 747 1715 753 1716
rect 747 1711 748 1715
rect 752 1714 753 1715
rect 814 1715 820 1716
rect 814 1714 815 1715
rect 752 1712 815 1714
rect 752 1711 753 1712
rect 747 1710 753 1711
rect 814 1711 815 1712
rect 819 1711 820 1715
rect 814 1710 820 1711
rect 915 1715 924 1716
rect 915 1711 916 1715
rect 923 1711 924 1715
rect 1106 1715 1112 1716
rect 915 1710 924 1711
rect 1074 1711 1080 1712
rect 498 1706 504 1707
rect 1074 1707 1075 1711
rect 1079 1710 1080 1711
rect 1083 1711 1089 1712
rect 1083 1710 1084 1711
rect 1079 1708 1084 1710
rect 1079 1707 1080 1708
rect 1074 1706 1080 1707
rect 1083 1707 1084 1708
rect 1088 1707 1089 1711
rect 1106 1711 1107 1715
rect 1111 1714 1112 1715
rect 1259 1715 1265 1716
rect 1259 1714 1260 1715
rect 1111 1712 1260 1714
rect 1111 1711 1112 1712
rect 1106 1710 1112 1711
rect 1259 1711 1260 1712
rect 1264 1711 1265 1715
rect 1259 1710 1265 1711
rect 1435 1715 1441 1716
rect 1435 1711 1436 1715
rect 1440 1714 1441 1715
rect 1466 1715 1472 1716
rect 1466 1714 1467 1715
rect 1440 1712 1467 1714
rect 1440 1711 1441 1712
rect 1435 1710 1441 1711
rect 1466 1711 1467 1712
rect 1471 1711 1472 1715
rect 1466 1710 1472 1711
rect 1518 1715 1524 1716
rect 1518 1711 1519 1715
rect 1523 1714 1524 1715
rect 1611 1715 1617 1716
rect 1611 1714 1612 1715
rect 1523 1712 1612 1714
rect 1523 1711 1524 1712
rect 1518 1710 1524 1711
rect 1611 1711 1612 1712
rect 1616 1711 1617 1715
rect 1611 1710 1617 1711
rect 1634 1715 1640 1716
rect 1634 1711 1635 1715
rect 1639 1714 1640 1715
rect 1795 1715 1801 1716
rect 1795 1714 1796 1715
rect 1639 1712 1796 1714
rect 1639 1711 1640 1712
rect 1634 1710 1640 1711
rect 1795 1711 1796 1712
rect 1800 1711 1801 1715
rect 2146 1715 2152 1716
rect 1795 1710 1801 1711
rect 2123 1713 2129 1714
rect 2123 1709 2124 1713
rect 2128 1709 2129 1713
rect 2146 1711 2147 1715
rect 2151 1714 2152 1715
rect 2243 1715 2249 1716
rect 2243 1714 2244 1715
rect 2151 1712 2244 1714
rect 2151 1711 2152 1712
rect 2146 1710 2152 1711
rect 2243 1711 2244 1712
rect 2248 1711 2249 1715
rect 2243 1710 2249 1711
rect 2266 1715 2272 1716
rect 2266 1711 2267 1715
rect 2271 1714 2272 1715
rect 2395 1715 2401 1716
rect 2395 1714 2396 1715
rect 2271 1712 2396 1714
rect 2271 1711 2272 1712
rect 2266 1710 2272 1711
rect 2395 1711 2396 1712
rect 2400 1711 2401 1715
rect 2395 1710 2401 1711
rect 2418 1715 2424 1716
rect 2418 1711 2419 1715
rect 2423 1714 2424 1715
rect 2563 1715 2569 1716
rect 2563 1714 2564 1715
rect 2423 1712 2564 1714
rect 2423 1711 2424 1712
rect 2418 1710 2424 1711
rect 2563 1711 2564 1712
rect 2568 1711 2569 1715
rect 2563 1710 2569 1711
rect 2739 1715 2745 1716
rect 2739 1711 2740 1715
rect 2744 1714 2745 1715
rect 2790 1715 2796 1716
rect 2790 1714 2791 1715
rect 2744 1712 2791 1714
rect 2744 1711 2745 1712
rect 2739 1710 2745 1711
rect 2790 1711 2791 1712
rect 2795 1711 2796 1715
rect 2790 1710 2796 1711
rect 2798 1715 2804 1716
rect 2798 1711 2799 1715
rect 2803 1714 2804 1715
rect 2923 1715 2929 1716
rect 2923 1714 2924 1715
rect 2803 1712 2924 1714
rect 2803 1711 2804 1712
rect 2798 1710 2804 1711
rect 2923 1711 2924 1712
rect 2928 1711 2929 1715
rect 2923 1710 2929 1711
rect 3115 1715 3124 1716
rect 3115 1711 3116 1715
rect 3123 1711 3124 1715
rect 3115 1710 3124 1711
rect 3138 1715 3144 1716
rect 3138 1711 3139 1715
rect 3143 1714 3144 1715
rect 3307 1715 3313 1716
rect 3307 1714 3308 1715
rect 3143 1712 3308 1714
rect 3143 1711 3144 1712
rect 3138 1710 3144 1711
rect 3307 1711 3308 1712
rect 3312 1711 3313 1715
rect 3307 1710 3313 1711
rect 3330 1715 3336 1716
rect 3330 1711 3331 1715
rect 3335 1714 3336 1715
rect 3499 1715 3505 1716
rect 3499 1714 3500 1715
rect 3335 1712 3500 1714
rect 3335 1711 3336 1712
rect 3330 1710 3336 1711
rect 3499 1711 3500 1712
rect 3504 1711 3505 1715
rect 3499 1710 3505 1711
rect 3699 1715 3705 1716
rect 3699 1711 3700 1715
rect 3704 1714 3705 1715
rect 3738 1715 3744 1716
rect 3738 1714 3739 1715
rect 3704 1712 3739 1714
rect 3704 1711 3705 1712
rect 3699 1710 3705 1711
rect 3738 1711 3739 1712
rect 3743 1711 3744 1715
rect 3738 1710 3744 1711
rect 3891 1715 3897 1716
rect 3891 1711 3892 1715
rect 3896 1714 3897 1715
rect 3914 1715 3920 1716
rect 3914 1714 3915 1715
rect 3896 1712 3915 1714
rect 3896 1711 3897 1712
rect 3891 1710 3897 1711
rect 3914 1711 3915 1712
rect 3919 1711 3920 1715
rect 3914 1710 3920 1711
rect 2123 1708 2129 1709
rect 1083 1706 1089 1707
rect 2124 1706 2126 1708
rect 2298 1707 2304 1708
rect 2298 1706 2299 1707
rect 2124 1704 2299 1706
rect 2298 1703 2299 1704
rect 2303 1703 2304 1707
rect 2298 1702 2304 1703
rect 187 1699 193 1700
rect 187 1695 188 1699
rect 192 1698 193 1699
rect 202 1699 208 1700
rect 202 1698 203 1699
rect 192 1696 203 1698
rect 192 1695 193 1696
rect 187 1694 193 1695
rect 202 1695 203 1696
rect 207 1695 208 1699
rect 202 1694 208 1695
rect 210 1699 216 1700
rect 210 1695 211 1699
rect 215 1698 216 1699
rect 315 1699 321 1700
rect 315 1698 316 1699
rect 215 1696 316 1698
rect 215 1695 216 1696
rect 210 1694 216 1695
rect 315 1695 316 1696
rect 320 1695 321 1699
rect 315 1694 321 1695
rect 338 1699 344 1700
rect 338 1695 339 1699
rect 343 1698 344 1699
rect 483 1699 489 1700
rect 483 1698 484 1699
rect 343 1696 484 1698
rect 343 1695 344 1696
rect 338 1694 344 1695
rect 483 1695 484 1696
rect 488 1695 489 1699
rect 483 1694 489 1695
rect 618 1699 624 1700
rect 618 1695 619 1699
rect 623 1698 624 1699
rect 659 1699 665 1700
rect 659 1698 660 1699
rect 623 1696 660 1698
rect 623 1695 624 1696
rect 618 1694 624 1695
rect 659 1695 660 1696
rect 664 1695 665 1699
rect 659 1694 665 1695
rect 682 1699 688 1700
rect 682 1695 683 1699
rect 687 1698 688 1699
rect 851 1699 857 1700
rect 851 1698 852 1699
rect 687 1696 852 1698
rect 687 1695 688 1696
rect 682 1694 688 1695
rect 851 1695 852 1696
rect 856 1695 857 1699
rect 1251 1699 1260 1700
rect 851 1694 857 1695
rect 1051 1697 1057 1698
rect 1051 1693 1052 1697
rect 1056 1693 1057 1697
rect 1251 1695 1252 1699
rect 1259 1695 1260 1699
rect 1251 1694 1260 1695
rect 1274 1699 1280 1700
rect 1274 1695 1275 1699
rect 1279 1698 1280 1699
rect 1459 1699 1465 1700
rect 1459 1698 1460 1699
rect 1279 1696 1460 1698
rect 1279 1695 1280 1696
rect 1274 1694 1280 1695
rect 1459 1695 1460 1696
rect 1464 1695 1465 1699
rect 1459 1694 1465 1695
rect 1675 1699 1681 1700
rect 1675 1695 1676 1699
rect 1680 1698 1681 1699
rect 1706 1699 1712 1700
rect 1706 1698 1707 1699
rect 1680 1696 1707 1698
rect 1680 1695 1681 1696
rect 1675 1694 1681 1695
rect 1706 1695 1707 1696
rect 1711 1695 1712 1699
rect 1706 1694 1712 1695
rect 1818 1699 1824 1700
rect 1818 1695 1819 1699
rect 1823 1698 1824 1699
rect 1891 1699 1897 1700
rect 1891 1698 1892 1699
rect 1823 1696 1892 1698
rect 1823 1695 1824 1696
rect 1818 1694 1824 1695
rect 1891 1695 1892 1696
rect 1896 1695 1897 1699
rect 1891 1694 1897 1695
rect 1051 1692 1057 1693
rect 2070 1692 2076 1693
rect 1052 1686 1054 1692
rect 2046 1689 2052 1690
rect 1302 1687 1308 1688
rect 1302 1686 1303 1687
rect 1052 1684 1303 1686
rect 1302 1683 1303 1684
rect 1307 1683 1308 1687
rect 2046 1685 2047 1689
rect 2051 1685 2052 1689
rect 2070 1688 2071 1692
rect 2075 1688 2076 1692
rect 2070 1687 2076 1688
rect 2190 1692 2196 1693
rect 2190 1688 2191 1692
rect 2195 1688 2196 1692
rect 2190 1687 2196 1688
rect 2342 1692 2348 1693
rect 2342 1688 2343 1692
rect 2347 1688 2348 1692
rect 2342 1687 2348 1688
rect 2510 1692 2516 1693
rect 2510 1688 2511 1692
rect 2515 1688 2516 1692
rect 2510 1687 2516 1688
rect 2686 1692 2692 1693
rect 2686 1688 2687 1692
rect 2691 1688 2692 1692
rect 2686 1687 2692 1688
rect 2870 1692 2876 1693
rect 2870 1688 2871 1692
rect 2875 1688 2876 1692
rect 2870 1687 2876 1688
rect 3062 1692 3068 1693
rect 3062 1688 3063 1692
rect 3067 1688 3068 1692
rect 3062 1687 3068 1688
rect 3254 1692 3260 1693
rect 3254 1688 3255 1692
rect 3259 1688 3260 1692
rect 3254 1687 3260 1688
rect 3446 1692 3452 1693
rect 3446 1688 3447 1692
rect 3451 1688 3452 1692
rect 3446 1687 3452 1688
rect 3646 1692 3652 1693
rect 3646 1688 3647 1692
rect 3651 1688 3652 1692
rect 3646 1687 3652 1688
rect 3838 1692 3844 1693
rect 3838 1688 3839 1692
rect 3843 1688 3844 1692
rect 3838 1687 3844 1688
rect 3942 1689 3948 1690
rect 2046 1684 2052 1685
rect 3942 1685 3943 1689
rect 3947 1685 3948 1689
rect 3942 1684 3948 1685
rect 1302 1682 1308 1683
rect 2146 1683 2152 1684
rect 2146 1679 2147 1683
rect 2151 1679 2152 1683
rect 2146 1678 2152 1679
rect 2266 1683 2272 1684
rect 2266 1679 2267 1683
rect 2271 1679 2272 1683
rect 2266 1678 2272 1679
rect 2418 1683 2424 1684
rect 2418 1679 2419 1683
rect 2423 1679 2424 1683
rect 2418 1678 2424 1679
rect 2578 1683 2584 1684
rect 2578 1679 2579 1683
rect 2583 1679 2584 1683
rect 2578 1678 2584 1679
rect 2654 1683 2660 1684
rect 2654 1679 2655 1683
rect 2659 1682 2660 1683
rect 2790 1683 2796 1684
rect 2659 1680 2729 1682
rect 2659 1679 2660 1680
rect 2654 1678 2660 1679
rect 2790 1679 2791 1683
rect 2795 1682 2796 1683
rect 3138 1683 3144 1684
rect 2795 1680 2913 1682
rect 2795 1679 2796 1680
rect 2790 1678 2796 1679
rect 3138 1679 3139 1683
rect 3143 1679 3144 1683
rect 3138 1678 3144 1679
rect 3330 1683 3336 1684
rect 3330 1679 3331 1683
rect 3335 1679 3336 1683
rect 3330 1678 3336 1679
rect 3514 1683 3520 1684
rect 3514 1679 3515 1683
rect 3519 1679 3520 1683
rect 3514 1678 3520 1679
rect 3614 1683 3620 1684
rect 3614 1679 3615 1683
rect 3619 1682 3620 1683
rect 3906 1683 3912 1684
rect 3619 1680 3689 1682
rect 3619 1679 3620 1680
rect 3614 1678 3620 1679
rect 3906 1679 3907 1683
rect 3911 1679 3912 1683
rect 3906 1678 3912 1679
rect 134 1676 140 1677
rect 110 1673 116 1674
rect 110 1669 111 1673
rect 115 1669 116 1673
rect 134 1672 135 1676
rect 139 1672 140 1676
rect 134 1671 140 1672
rect 262 1676 268 1677
rect 262 1672 263 1676
rect 267 1672 268 1676
rect 262 1671 268 1672
rect 430 1676 436 1677
rect 430 1672 431 1676
rect 435 1672 436 1676
rect 430 1671 436 1672
rect 606 1676 612 1677
rect 606 1672 607 1676
rect 611 1672 612 1676
rect 606 1671 612 1672
rect 798 1676 804 1677
rect 798 1672 799 1676
rect 803 1672 804 1676
rect 798 1671 804 1672
rect 998 1676 1004 1677
rect 998 1672 999 1676
rect 1003 1672 1004 1676
rect 998 1671 1004 1672
rect 1198 1676 1204 1677
rect 1198 1672 1199 1676
rect 1203 1672 1204 1676
rect 1198 1671 1204 1672
rect 1406 1676 1412 1677
rect 1406 1672 1407 1676
rect 1411 1672 1412 1676
rect 1406 1671 1412 1672
rect 1622 1676 1628 1677
rect 1622 1672 1623 1676
rect 1627 1672 1628 1676
rect 1622 1671 1628 1672
rect 1838 1676 1844 1677
rect 1838 1672 1839 1676
rect 1843 1672 1844 1676
rect 1838 1671 1844 1672
rect 2006 1673 2012 1674
rect 2070 1673 2076 1674
rect 110 1668 116 1669
rect 2006 1669 2007 1673
rect 2011 1669 2012 1673
rect 2006 1668 2012 1669
rect 2046 1672 2052 1673
rect 2046 1668 2047 1672
rect 2051 1668 2052 1672
rect 2070 1669 2071 1673
rect 2075 1669 2076 1673
rect 2070 1668 2076 1669
rect 2190 1673 2196 1674
rect 2190 1669 2191 1673
rect 2195 1669 2196 1673
rect 2190 1668 2196 1669
rect 2342 1673 2348 1674
rect 2342 1669 2343 1673
rect 2347 1669 2348 1673
rect 2342 1668 2348 1669
rect 2510 1673 2516 1674
rect 2510 1669 2511 1673
rect 2515 1669 2516 1673
rect 2510 1668 2516 1669
rect 2686 1673 2692 1674
rect 2686 1669 2687 1673
rect 2691 1669 2692 1673
rect 2686 1668 2692 1669
rect 2870 1673 2876 1674
rect 2870 1669 2871 1673
rect 2875 1669 2876 1673
rect 2870 1668 2876 1669
rect 3062 1673 3068 1674
rect 3062 1669 3063 1673
rect 3067 1669 3068 1673
rect 3062 1668 3068 1669
rect 3254 1673 3260 1674
rect 3254 1669 3255 1673
rect 3259 1669 3260 1673
rect 3254 1668 3260 1669
rect 3446 1673 3452 1674
rect 3446 1669 3447 1673
rect 3451 1669 3452 1673
rect 3446 1668 3452 1669
rect 3646 1673 3652 1674
rect 3646 1669 3647 1673
rect 3651 1669 3652 1673
rect 3646 1668 3652 1669
rect 3838 1673 3844 1674
rect 3838 1669 3839 1673
rect 3843 1669 3844 1673
rect 3838 1668 3844 1669
rect 3942 1672 3948 1673
rect 3942 1668 3943 1672
rect 3947 1668 3948 1672
rect 210 1667 216 1668
rect 210 1663 211 1667
rect 215 1663 216 1667
rect 210 1662 216 1663
rect 338 1667 344 1668
rect 338 1663 339 1667
rect 343 1663 344 1667
rect 338 1662 344 1663
rect 498 1667 504 1668
rect 498 1663 499 1667
rect 503 1663 504 1667
rect 498 1662 504 1663
rect 682 1667 688 1668
rect 682 1663 683 1667
rect 687 1663 688 1667
rect 682 1662 688 1663
rect 874 1667 880 1668
rect 874 1663 875 1667
rect 879 1663 880 1667
rect 874 1662 880 1663
rect 1074 1667 1080 1668
rect 1074 1663 1075 1667
rect 1079 1663 1080 1667
rect 1074 1662 1080 1663
rect 1274 1667 1280 1668
rect 1274 1663 1275 1667
rect 1279 1663 1280 1667
rect 1274 1662 1280 1663
rect 1302 1667 1308 1668
rect 1302 1663 1303 1667
rect 1307 1666 1308 1667
rect 1558 1667 1564 1668
rect 1307 1664 1449 1666
rect 1307 1663 1308 1664
rect 1302 1662 1308 1663
rect 1558 1663 1559 1667
rect 1563 1666 1564 1667
rect 1706 1667 1712 1668
rect 2046 1667 2052 1668
rect 3942 1667 3948 1668
rect 1563 1664 1665 1666
rect 1563 1663 1564 1664
rect 1558 1662 1564 1663
rect 1706 1663 1707 1667
rect 1711 1666 1712 1667
rect 1711 1664 1881 1666
rect 1711 1663 1712 1664
rect 1706 1662 1712 1663
rect 134 1657 140 1658
rect 110 1656 116 1657
rect 110 1652 111 1656
rect 115 1652 116 1656
rect 134 1653 135 1657
rect 139 1653 140 1657
rect 134 1652 140 1653
rect 262 1657 268 1658
rect 262 1653 263 1657
rect 267 1653 268 1657
rect 262 1652 268 1653
rect 430 1657 436 1658
rect 430 1653 431 1657
rect 435 1653 436 1657
rect 430 1652 436 1653
rect 606 1657 612 1658
rect 606 1653 607 1657
rect 611 1653 612 1657
rect 606 1652 612 1653
rect 798 1657 804 1658
rect 798 1653 799 1657
rect 803 1653 804 1657
rect 798 1652 804 1653
rect 998 1657 1004 1658
rect 998 1653 999 1657
rect 1003 1653 1004 1657
rect 998 1652 1004 1653
rect 1198 1657 1204 1658
rect 1198 1653 1199 1657
rect 1203 1653 1204 1657
rect 1198 1652 1204 1653
rect 1406 1657 1412 1658
rect 1406 1653 1407 1657
rect 1411 1653 1412 1657
rect 1406 1652 1412 1653
rect 1622 1657 1628 1658
rect 1622 1653 1623 1657
rect 1627 1653 1628 1657
rect 1622 1652 1628 1653
rect 1838 1657 1844 1658
rect 1838 1653 1839 1657
rect 1843 1653 1844 1657
rect 1838 1652 1844 1653
rect 2006 1656 2012 1657
rect 2006 1652 2007 1656
rect 2011 1652 2012 1656
rect 110 1651 116 1652
rect 2006 1651 2012 1652
rect 2046 1620 2052 1621
rect 3942 1620 3948 1621
rect 2046 1616 2047 1620
rect 2051 1616 2052 1620
rect 2046 1615 2052 1616
rect 2070 1619 2076 1620
rect 2070 1615 2071 1619
rect 2075 1615 2076 1619
rect 2070 1614 2076 1615
rect 2334 1619 2340 1620
rect 2334 1615 2335 1619
rect 2339 1615 2340 1619
rect 2334 1614 2340 1615
rect 2598 1619 2604 1620
rect 2598 1615 2599 1619
rect 2603 1615 2604 1619
rect 2598 1614 2604 1615
rect 2838 1619 2844 1620
rect 2838 1615 2839 1619
rect 2843 1615 2844 1619
rect 2838 1614 2844 1615
rect 3046 1619 3052 1620
rect 3046 1615 3047 1619
rect 3051 1615 3052 1619
rect 3046 1614 3052 1615
rect 3230 1619 3236 1620
rect 3230 1615 3231 1619
rect 3235 1615 3236 1619
rect 3230 1614 3236 1615
rect 3398 1619 3404 1620
rect 3398 1615 3399 1619
rect 3403 1615 3404 1619
rect 3398 1614 3404 1615
rect 3550 1619 3556 1620
rect 3550 1615 3551 1619
rect 3555 1615 3556 1619
rect 3550 1614 3556 1615
rect 3694 1619 3700 1620
rect 3694 1615 3695 1619
rect 3699 1615 3700 1619
rect 3694 1614 3700 1615
rect 3838 1619 3844 1620
rect 3838 1615 3839 1619
rect 3843 1615 3844 1619
rect 3942 1616 3943 1620
rect 3947 1616 3948 1620
rect 3942 1615 3948 1616
rect 3838 1614 3844 1615
rect 2298 1611 2304 1612
rect 2146 1607 2152 1608
rect 110 1604 116 1605
rect 2006 1604 2012 1605
rect 110 1600 111 1604
rect 115 1600 116 1604
rect 110 1599 116 1600
rect 134 1603 140 1604
rect 134 1599 135 1603
rect 139 1599 140 1603
rect 286 1603 292 1604
rect 134 1598 140 1599
rect 202 1599 208 1600
rect 202 1595 203 1599
rect 207 1598 208 1599
rect 286 1599 287 1603
rect 291 1599 292 1603
rect 286 1598 292 1599
rect 470 1603 476 1604
rect 470 1599 471 1603
rect 475 1599 476 1603
rect 470 1598 476 1599
rect 654 1603 660 1604
rect 654 1599 655 1603
rect 659 1599 660 1603
rect 654 1598 660 1599
rect 838 1603 844 1604
rect 838 1599 839 1603
rect 843 1599 844 1603
rect 838 1598 844 1599
rect 1014 1603 1020 1604
rect 1014 1599 1015 1603
rect 1019 1599 1020 1603
rect 1014 1598 1020 1599
rect 1182 1603 1188 1604
rect 1182 1599 1183 1603
rect 1187 1599 1188 1603
rect 1182 1598 1188 1599
rect 1342 1603 1348 1604
rect 1342 1599 1343 1603
rect 1347 1599 1348 1603
rect 1342 1598 1348 1599
rect 1494 1603 1500 1604
rect 1494 1599 1495 1603
rect 1499 1599 1500 1603
rect 1494 1598 1500 1599
rect 1638 1603 1644 1604
rect 1638 1599 1639 1603
rect 1643 1599 1644 1603
rect 1638 1598 1644 1599
rect 1782 1603 1788 1604
rect 1782 1599 1783 1603
rect 1787 1599 1788 1603
rect 1782 1598 1788 1599
rect 1902 1603 1908 1604
rect 1902 1599 1903 1603
rect 1907 1599 1908 1603
rect 2006 1600 2007 1604
rect 2011 1600 2012 1604
rect 2006 1599 2012 1600
rect 2046 1603 2052 1604
rect 2046 1599 2047 1603
rect 2051 1599 2052 1603
rect 2146 1603 2147 1607
rect 2151 1603 2152 1607
rect 2298 1607 2299 1611
rect 2303 1610 2304 1611
rect 3122 1611 3128 1612
rect 2303 1608 2377 1610
rect 2303 1607 2304 1608
rect 2298 1606 2304 1607
rect 2674 1607 2680 1608
rect 2146 1602 2152 1603
rect 2674 1603 2675 1607
rect 2679 1603 2680 1607
rect 2674 1602 2680 1603
rect 2914 1607 2920 1608
rect 2914 1603 2915 1607
rect 2919 1603 2920 1607
rect 3122 1607 3123 1611
rect 3127 1607 3128 1611
rect 3122 1606 3128 1607
rect 3130 1611 3136 1612
rect 3130 1607 3131 1611
rect 3135 1610 3136 1611
rect 3354 1611 3360 1612
rect 3135 1608 3273 1610
rect 3135 1607 3136 1608
rect 3130 1606 3136 1607
rect 3354 1607 3355 1611
rect 3359 1610 3360 1611
rect 3914 1611 3920 1612
rect 3359 1608 3441 1610
rect 3359 1607 3360 1608
rect 3354 1606 3360 1607
rect 3626 1607 3632 1608
rect 2914 1602 2920 1603
rect 3626 1603 3627 1607
rect 3631 1603 3632 1607
rect 3626 1602 3632 1603
rect 3770 1607 3776 1608
rect 3770 1603 3771 1607
rect 3775 1603 3776 1607
rect 3914 1607 3915 1611
rect 3919 1607 3920 1611
rect 3914 1606 3920 1607
rect 3770 1602 3776 1603
rect 3942 1603 3948 1604
rect 1902 1598 1908 1599
rect 2046 1598 2052 1599
rect 2070 1600 2076 1601
rect 207 1596 214 1598
rect 2070 1596 2071 1600
rect 2075 1596 2076 1600
rect 207 1595 208 1596
rect 202 1594 208 1595
rect 212 1593 214 1596
rect 222 1595 228 1596
rect 222 1591 223 1595
rect 227 1594 228 1595
rect 738 1595 744 1596
rect 227 1592 329 1594
rect 227 1591 228 1592
rect 222 1590 228 1591
rect 546 1591 552 1592
rect 110 1587 116 1588
rect 110 1583 111 1587
rect 115 1583 116 1587
rect 546 1587 547 1591
rect 551 1587 552 1591
rect 546 1586 552 1587
rect 730 1591 736 1592
rect 730 1587 731 1591
rect 735 1587 736 1591
rect 738 1591 739 1595
rect 743 1594 744 1595
rect 1258 1595 1264 1596
rect 743 1592 881 1594
rect 743 1591 744 1592
rect 738 1590 744 1591
rect 1118 1591 1124 1592
rect 1118 1590 1119 1591
rect 1093 1588 1119 1590
rect 730 1586 736 1587
rect 1118 1587 1119 1588
rect 1123 1587 1124 1591
rect 1258 1591 1259 1595
rect 1263 1591 1264 1595
rect 1258 1590 1264 1591
rect 1278 1595 1284 1596
rect 2070 1595 2076 1596
rect 2334 1600 2340 1601
rect 2334 1596 2335 1600
rect 2339 1596 2340 1600
rect 2334 1595 2340 1596
rect 2598 1600 2604 1601
rect 2598 1596 2599 1600
rect 2603 1596 2604 1600
rect 2598 1595 2604 1596
rect 2838 1600 2844 1601
rect 2838 1596 2839 1600
rect 2843 1596 2844 1600
rect 2838 1595 2844 1596
rect 3046 1600 3052 1601
rect 3046 1596 3047 1600
rect 3051 1596 3052 1600
rect 3046 1595 3052 1596
rect 3230 1600 3236 1601
rect 3230 1596 3231 1600
rect 3235 1596 3236 1600
rect 3230 1595 3236 1596
rect 3398 1600 3404 1601
rect 3398 1596 3399 1600
rect 3403 1596 3404 1600
rect 3398 1595 3404 1596
rect 3550 1600 3556 1601
rect 3550 1596 3551 1600
rect 3555 1596 3556 1600
rect 3550 1595 3556 1596
rect 3694 1600 3700 1601
rect 3694 1596 3695 1600
rect 3699 1596 3700 1600
rect 3694 1595 3700 1596
rect 3838 1600 3844 1601
rect 3838 1596 3839 1600
rect 3843 1596 3844 1600
rect 3942 1599 3943 1603
rect 3947 1599 3948 1603
rect 3942 1598 3948 1599
rect 3838 1595 3844 1596
rect 1278 1591 1279 1595
rect 1283 1594 1284 1595
rect 1283 1592 1385 1594
rect 1283 1591 1284 1592
rect 1278 1590 1284 1591
rect 1570 1591 1576 1592
rect 1118 1586 1124 1587
rect 1570 1587 1571 1591
rect 1575 1587 1576 1591
rect 1570 1586 1576 1587
rect 1714 1591 1720 1592
rect 1714 1587 1715 1591
rect 1719 1587 1720 1591
rect 1714 1586 1720 1587
rect 1858 1591 1864 1592
rect 1858 1587 1859 1591
rect 1863 1587 1864 1591
rect 1981 1588 2001 1590
rect 1858 1586 1864 1587
rect 110 1582 116 1583
rect 134 1584 140 1585
rect 134 1580 135 1584
rect 139 1580 140 1584
rect 134 1579 140 1580
rect 286 1584 292 1585
rect 286 1580 287 1584
rect 291 1580 292 1584
rect 286 1579 292 1580
rect 470 1584 476 1585
rect 470 1580 471 1584
rect 475 1580 476 1584
rect 470 1579 476 1580
rect 654 1584 660 1585
rect 654 1580 655 1584
rect 659 1580 660 1584
rect 654 1579 660 1580
rect 838 1584 844 1585
rect 838 1580 839 1584
rect 843 1580 844 1584
rect 838 1579 844 1580
rect 1014 1584 1020 1585
rect 1014 1580 1015 1584
rect 1019 1580 1020 1584
rect 1014 1579 1020 1580
rect 1182 1584 1188 1585
rect 1182 1580 1183 1584
rect 1187 1580 1188 1584
rect 1182 1579 1188 1580
rect 1342 1584 1348 1585
rect 1342 1580 1343 1584
rect 1347 1580 1348 1584
rect 1342 1579 1348 1580
rect 1494 1584 1500 1585
rect 1494 1580 1495 1584
rect 1499 1580 1500 1584
rect 1494 1579 1500 1580
rect 1638 1584 1644 1585
rect 1638 1580 1639 1584
rect 1643 1580 1644 1584
rect 1638 1579 1644 1580
rect 1782 1584 1788 1585
rect 1782 1580 1783 1584
rect 1787 1580 1788 1584
rect 1782 1579 1788 1580
rect 1902 1584 1908 1585
rect 1902 1580 1903 1584
rect 1907 1580 1908 1584
rect 1902 1579 1908 1580
rect 1999 1578 2001 1588
rect 2006 1587 2012 1588
rect 2006 1583 2007 1587
rect 2011 1583 2012 1587
rect 3130 1587 3136 1588
rect 3130 1586 3131 1587
rect 2006 1582 2012 1583
rect 2908 1584 3131 1586
rect 2123 1579 2129 1580
rect 2123 1578 2124 1579
rect 1999 1576 2124 1578
rect 2123 1575 2124 1576
rect 2128 1575 2129 1579
rect 2123 1574 2129 1575
rect 2146 1579 2152 1580
rect 2146 1575 2147 1579
rect 2151 1578 2152 1579
rect 2387 1579 2393 1580
rect 2387 1578 2388 1579
rect 2151 1576 2388 1578
rect 2151 1575 2152 1576
rect 2146 1574 2152 1575
rect 2387 1575 2388 1576
rect 2392 1575 2393 1579
rect 2387 1574 2393 1575
rect 2651 1579 2660 1580
rect 2651 1575 2652 1579
rect 2659 1575 2660 1579
rect 2651 1574 2660 1575
rect 2891 1579 2897 1580
rect 2891 1575 2892 1579
rect 2896 1578 2897 1579
rect 2908 1578 2910 1584
rect 3130 1583 3131 1584
rect 3135 1583 3136 1587
rect 3130 1582 3136 1583
rect 2896 1576 2910 1578
rect 2914 1579 2920 1580
rect 2896 1575 2897 1576
rect 2891 1574 2897 1575
rect 2914 1575 2915 1579
rect 2919 1578 2920 1579
rect 3099 1579 3105 1580
rect 3099 1578 3100 1579
rect 2919 1576 3100 1578
rect 2919 1575 2920 1576
rect 2914 1574 2920 1575
rect 3099 1575 3100 1576
rect 3104 1575 3105 1579
rect 3099 1574 3105 1575
rect 3283 1579 3289 1580
rect 3283 1575 3284 1579
rect 3288 1578 3289 1579
rect 3354 1579 3360 1580
rect 3354 1578 3355 1579
rect 3288 1576 3355 1578
rect 3288 1575 3289 1576
rect 3283 1574 3289 1575
rect 3354 1575 3355 1576
rect 3359 1575 3360 1579
rect 3603 1579 3609 1580
rect 3354 1574 3360 1575
rect 3450 1575 3457 1576
rect 738 1571 744 1572
rect 738 1570 739 1571
rect 540 1568 739 1570
rect 187 1563 193 1564
rect 187 1559 188 1563
rect 192 1562 193 1563
rect 222 1563 228 1564
rect 222 1562 223 1563
rect 192 1560 223 1562
rect 192 1559 193 1560
rect 187 1558 193 1559
rect 222 1559 223 1560
rect 227 1559 228 1563
rect 523 1563 529 1564
rect 222 1558 228 1559
rect 339 1559 345 1560
rect 339 1555 340 1559
rect 344 1558 345 1559
rect 390 1559 396 1560
rect 390 1558 391 1559
rect 344 1556 391 1558
rect 344 1555 345 1556
rect 339 1554 345 1555
rect 390 1555 391 1556
rect 395 1555 396 1559
rect 523 1559 524 1563
rect 528 1562 529 1563
rect 540 1562 542 1568
rect 738 1567 739 1568
rect 743 1567 744 1571
rect 1278 1571 1284 1572
rect 1278 1570 1279 1571
rect 738 1566 744 1567
rect 1159 1568 1279 1570
rect 1159 1566 1161 1568
rect 1278 1567 1279 1568
rect 1283 1567 1284 1571
rect 3450 1571 3451 1575
rect 3456 1571 3457 1575
rect 3603 1575 3604 1579
rect 3608 1578 3609 1579
rect 3614 1579 3620 1580
rect 3614 1578 3615 1579
rect 3608 1576 3615 1578
rect 3608 1575 3609 1576
rect 3603 1574 3609 1575
rect 3614 1575 3615 1576
rect 3619 1575 3620 1579
rect 3614 1574 3620 1575
rect 3626 1579 3632 1580
rect 3626 1575 3627 1579
rect 3631 1578 3632 1579
rect 3747 1579 3753 1580
rect 3747 1578 3748 1579
rect 3631 1576 3748 1578
rect 3631 1575 3632 1576
rect 3626 1574 3632 1575
rect 3747 1575 3748 1576
rect 3752 1575 3753 1579
rect 3747 1574 3753 1575
rect 3890 1575 3897 1576
rect 3450 1570 3457 1571
rect 3890 1571 3891 1575
rect 3896 1571 3897 1575
rect 3890 1570 3897 1571
rect 1278 1566 1284 1567
rect 1112 1564 1161 1566
rect 528 1560 542 1562
rect 546 1563 552 1564
rect 528 1559 529 1560
rect 523 1558 529 1559
rect 546 1559 547 1563
rect 551 1562 552 1563
rect 707 1563 713 1564
rect 707 1562 708 1563
rect 551 1560 708 1562
rect 551 1559 552 1560
rect 546 1558 552 1559
rect 707 1559 708 1560
rect 712 1559 713 1563
rect 707 1558 713 1559
rect 874 1563 880 1564
rect 874 1559 875 1563
rect 879 1562 880 1563
rect 891 1563 897 1564
rect 891 1562 892 1563
rect 879 1560 892 1562
rect 879 1559 880 1560
rect 874 1558 880 1559
rect 891 1559 892 1560
rect 896 1559 897 1563
rect 891 1558 897 1559
rect 1067 1563 1073 1564
rect 1067 1559 1068 1563
rect 1072 1562 1073 1563
rect 1112 1562 1114 1564
rect 1235 1563 1241 1564
rect 1235 1562 1236 1563
rect 1072 1560 1114 1562
rect 1159 1560 1236 1562
rect 1072 1559 1073 1560
rect 1067 1558 1073 1559
rect 1118 1559 1124 1560
rect 390 1554 396 1555
rect 1118 1555 1119 1559
rect 1123 1558 1124 1559
rect 1159 1558 1161 1560
rect 1235 1559 1236 1560
rect 1240 1559 1241 1563
rect 1547 1563 1553 1564
rect 1235 1558 1241 1559
rect 1350 1559 1356 1560
rect 1123 1556 1161 1558
rect 1123 1555 1124 1556
rect 1118 1554 1124 1555
rect 1350 1555 1351 1559
rect 1355 1558 1356 1559
rect 1395 1559 1401 1560
rect 1395 1558 1396 1559
rect 1355 1556 1396 1558
rect 1355 1555 1356 1556
rect 1350 1554 1356 1555
rect 1395 1555 1396 1556
rect 1400 1555 1401 1559
rect 1547 1559 1548 1563
rect 1552 1562 1553 1563
rect 1558 1563 1564 1564
rect 1558 1562 1559 1563
rect 1552 1560 1559 1562
rect 1552 1559 1553 1560
rect 1547 1558 1553 1559
rect 1558 1559 1559 1560
rect 1563 1559 1564 1563
rect 1558 1558 1564 1559
rect 1570 1563 1576 1564
rect 1570 1559 1571 1563
rect 1575 1562 1576 1563
rect 1691 1563 1697 1564
rect 1691 1562 1692 1563
rect 1575 1560 1692 1562
rect 1575 1559 1576 1560
rect 1570 1558 1576 1559
rect 1691 1559 1692 1560
rect 1696 1559 1697 1563
rect 1691 1558 1697 1559
rect 1714 1563 1720 1564
rect 1714 1559 1715 1563
rect 1719 1562 1720 1563
rect 1835 1563 1841 1564
rect 1835 1562 1836 1563
rect 1719 1560 1836 1562
rect 1719 1559 1720 1560
rect 1714 1558 1720 1559
rect 1835 1559 1836 1560
rect 1840 1559 1841 1563
rect 1835 1558 1841 1559
rect 1858 1563 1864 1564
rect 1858 1559 1859 1563
rect 1863 1562 1864 1563
rect 1955 1563 1961 1564
rect 1955 1562 1956 1563
rect 1863 1560 1956 1562
rect 1863 1559 1864 1560
rect 1858 1558 1864 1559
rect 1955 1559 1956 1560
rect 1960 1559 1961 1563
rect 1955 1558 1961 1559
rect 2635 1559 2641 1560
rect 1395 1554 1401 1555
rect 2635 1555 2636 1559
rect 2640 1558 2641 1559
rect 2674 1559 2680 1560
rect 2674 1558 2675 1559
rect 2640 1556 2675 1558
rect 2640 1555 2641 1556
rect 2635 1554 2641 1555
rect 2674 1555 2675 1556
rect 2679 1555 2680 1559
rect 2674 1554 2680 1555
rect 2710 1559 2716 1560
rect 2710 1555 2711 1559
rect 2715 1558 2716 1559
rect 2795 1559 2801 1560
rect 2795 1558 2796 1559
rect 2715 1556 2796 1558
rect 2715 1555 2716 1556
rect 2710 1554 2716 1555
rect 2795 1555 2796 1556
rect 2800 1555 2801 1559
rect 2795 1554 2801 1555
rect 2818 1559 2824 1560
rect 2818 1555 2819 1559
rect 2823 1558 2824 1559
rect 2955 1559 2961 1560
rect 2955 1558 2956 1559
rect 2823 1556 2956 1558
rect 2823 1555 2824 1556
rect 2818 1554 2824 1555
rect 2955 1555 2956 1556
rect 2960 1555 2961 1559
rect 2955 1554 2961 1555
rect 2978 1559 2984 1560
rect 2978 1555 2979 1559
rect 2983 1558 2984 1559
rect 3115 1559 3121 1560
rect 3115 1558 3116 1559
rect 2983 1556 3116 1558
rect 2983 1555 2984 1556
rect 2978 1554 2984 1555
rect 3115 1555 3116 1556
rect 3120 1555 3121 1559
rect 3298 1559 3304 1560
rect 3115 1554 3121 1555
rect 3275 1557 3281 1558
rect 3275 1553 3276 1557
rect 3280 1553 3281 1557
rect 3298 1555 3299 1559
rect 3303 1558 3304 1559
rect 3435 1559 3441 1560
rect 3435 1558 3436 1559
rect 3303 1556 3436 1558
rect 3303 1555 3304 1556
rect 3298 1554 3304 1555
rect 3435 1555 3436 1556
rect 3440 1555 3441 1559
rect 3435 1554 3441 1555
rect 3595 1559 3601 1560
rect 3595 1555 3596 1559
rect 3600 1558 3601 1559
rect 3638 1559 3644 1560
rect 3638 1558 3639 1559
rect 3600 1556 3639 1558
rect 3600 1555 3601 1556
rect 3595 1554 3601 1555
rect 3638 1555 3639 1556
rect 3643 1555 3644 1559
rect 3638 1554 3644 1555
rect 3755 1559 3761 1560
rect 3755 1555 3756 1559
rect 3760 1558 3761 1559
rect 3770 1559 3776 1560
rect 3770 1558 3771 1559
rect 3760 1556 3771 1558
rect 3760 1555 3761 1556
rect 3755 1554 3761 1555
rect 3770 1555 3771 1556
rect 3775 1555 3776 1559
rect 3770 1554 3776 1555
rect 3275 1552 3281 1553
rect 3276 1550 3278 1552
rect 3498 1551 3504 1552
rect 3498 1550 3499 1551
rect 3276 1548 3499 1550
rect 3498 1547 3499 1548
rect 3503 1547 3504 1551
rect 3498 1546 3504 1547
rect 187 1543 193 1544
rect 187 1539 188 1543
rect 192 1542 193 1543
rect 250 1543 256 1544
rect 250 1542 251 1543
rect 192 1540 251 1542
rect 192 1539 193 1540
rect 187 1538 193 1539
rect 250 1539 251 1540
rect 255 1539 256 1543
rect 250 1538 256 1539
rect 258 1543 264 1544
rect 258 1539 259 1543
rect 263 1542 264 1543
rect 347 1543 353 1544
rect 347 1542 348 1543
rect 263 1540 348 1542
rect 263 1539 264 1540
rect 258 1538 264 1539
rect 347 1539 348 1540
rect 352 1539 353 1543
rect 347 1538 353 1539
rect 370 1543 376 1544
rect 370 1539 371 1543
rect 375 1542 376 1543
rect 539 1543 545 1544
rect 539 1542 540 1543
rect 375 1540 540 1542
rect 375 1539 376 1540
rect 370 1538 376 1539
rect 539 1539 540 1540
rect 544 1539 545 1543
rect 539 1538 545 1539
rect 730 1543 736 1544
rect 730 1539 731 1543
rect 735 1542 736 1543
rect 739 1543 745 1544
rect 739 1542 740 1543
rect 735 1540 740 1542
rect 735 1539 736 1540
rect 730 1538 736 1539
rect 739 1539 740 1540
rect 744 1539 745 1543
rect 739 1538 745 1539
rect 762 1543 768 1544
rect 762 1539 763 1543
rect 767 1542 768 1543
rect 939 1543 945 1544
rect 939 1542 940 1543
rect 767 1540 940 1542
rect 767 1539 768 1540
rect 762 1538 768 1539
rect 939 1539 940 1540
rect 944 1539 945 1543
rect 1154 1543 1160 1544
rect 939 1538 945 1539
rect 1131 1541 1137 1542
rect 1131 1537 1132 1541
rect 1136 1537 1137 1541
rect 1154 1539 1155 1543
rect 1159 1542 1160 1543
rect 1315 1543 1321 1544
rect 1315 1542 1316 1543
rect 1159 1540 1316 1542
rect 1159 1539 1160 1540
rect 1154 1538 1160 1539
rect 1315 1539 1316 1540
rect 1320 1539 1321 1543
rect 1315 1538 1321 1539
rect 1499 1543 1505 1544
rect 1499 1539 1500 1543
rect 1504 1542 1505 1543
rect 1530 1543 1536 1544
rect 1530 1542 1531 1543
rect 1504 1540 1531 1542
rect 1504 1539 1505 1540
rect 1499 1538 1505 1539
rect 1530 1539 1531 1540
rect 1535 1539 1536 1543
rect 1530 1538 1536 1539
rect 1675 1543 1681 1544
rect 1675 1539 1676 1543
rect 1680 1542 1681 1543
rect 1706 1543 1712 1544
rect 1706 1542 1707 1543
rect 1680 1540 1707 1542
rect 1680 1539 1681 1540
rect 1675 1538 1681 1539
rect 1706 1539 1707 1540
rect 1711 1539 1712 1543
rect 1706 1538 1712 1539
rect 1859 1543 1868 1544
rect 1859 1539 1860 1543
rect 1867 1539 1868 1543
rect 1859 1538 1868 1539
rect 1131 1536 1137 1537
rect 2582 1536 2588 1537
rect 1132 1534 1134 1536
rect 1398 1535 1404 1536
rect 1398 1534 1399 1535
rect 1132 1532 1399 1534
rect 1398 1531 1399 1532
rect 1403 1531 1404 1535
rect 1398 1530 1404 1531
rect 2046 1533 2052 1534
rect 2046 1529 2047 1533
rect 2051 1529 2052 1533
rect 2582 1532 2583 1536
rect 2587 1532 2588 1536
rect 2582 1531 2588 1532
rect 2742 1536 2748 1537
rect 2742 1532 2743 1536
rect 2747 1532 2748 1536
rect 2742 1531 2748 1532
rect 2902 1536 2908 1537
rect 2902 1532 2903 1536
rect 2907 1532 2908 1536
rect 2902 1531 2908 1532
rect 3062 1536 3068 1537
rect 3062 1532 3063 1536
rect 3067 1532 3068 1536
rect 3062 1531 3068 1532
rect 3222 1536 3228 1537
rect 3222 1532 3223 1536
rect 3227 1532 3228 1536
rect 3222 1531 3228 1532
rect 3382 1536 3388 1537
rect 3382 1532 3383 1536
rect 3387 1532 3388 1536
rect 3382 1531 3388 1532
rect 3542 1536 3548 1537
rect 3542 1532 3543 1536
rect 3547 1532 3548 1536
rect 3542 1531 3548 1532
rect 3702 1536 3708 1537
rect 3702 1532 3703 1536
rect 3707 1532 3708 1536
rect 3702 1531 3708 1532
rect 3942 1533 3948 1534
rect 2046 1528 2052 1529
rect 3942 1529 3943 1533
rect 3947 1529 3948 1533
rect 3942 1528 3948 1529
rect 2710 1527 2716 1528
rect 2710 1526 2711 1527
rect 2661 1524 2711 1526
rect 2710 1523 2711 1524
rect 2715 1523 2716 1527
rect 2710 1522 2716 1523
rect 2818 1527 2824 1528
rect 2818 1523 2819 1527
rect 2823 1523 2824 1527
rect 2818 1522 2824 1523
rect 2978 1527 2984 1528
rect 2978 1523 2979 1527
rect 2983 1523 2984 1527
rect 2978 1522 2984 1523
rect 3018 1527 3024 1528
rect 3018 1523 3019 1527
rect 3023 1526 3024 1527
rect 3298 1527 3304 1528
rect 3023 1524 3105 1526
rect 3023 1523 3024 1524
rect 3018 1522 3024 1523
rect 3298 1523 3299 1527
rect 3303 1523 3304 1527
rect 3298 1522 3304 1523
rect 3450 1527 3456 1528
rect 3450 1523 3451 1527
rect 3455 1523 3456 1527
rect 3450 1522 3456 1523
rect 3498 1527 3504 1528
rect 3498 1523 3499 1527
rect 3503 1526 3504 1527
rect 3638 1527 3644 1528
rect 3503 1524 3585 1526
rect 3503 1523 3504 1524
rect 3498 1522 3504 1523
rect 3638 1523 3639 1527
rect 3643 1526 3644 1527
rect 3643 1524 3745 1526
rect 3643 1523 3644 1524
rect 3638 1522 3644 1523
rect 134 1520 140 1521
rect 110 1517 116 1518
rect 110 1513 111 1517
rect 115 1513 116 1517
rect 134 1516 135 1520
rect 139 1516 140 1520
rect 134 1515 140 1516
rect 294 1520 300 1521
rect 294 1516 295 1520
rect 299 1516 300 1520
rect 294 1515 300 1516
rect 486 1520 492 1521
rect 486 1516 487 1520
rect 491 1516 492 1520
rect 486 1515 492 1516
rect 686 1520 692 1521
rect 686 1516 687 1520
rect 691 1516 692 1520
rect 686 1515 692 1516
rect 886 1520 892 1521
rect 886 1516 887 1520
rect 891 1516 892 1520
rect 886 1515 892 1516
rect 1078 1520 1084 1521
rect 1078 1516 1079 1520
rect 1083 1516 1084 1520
rect 1078 1515 1084 1516
rect 1262 1520 1268 1521
rect 1262 1516 1263 1520
rect 1267 1516 1268 1520
rect 1262 1515 1268 1516
rect 1446 1520 1452 1521
rect 1446 1516 1447 1520
rect 1451 1516 1452 1520
rect 1446 1515 1452 1516
rect 1622 1520 1628 1521
rect 1622 1516 1623 1520
rect 1627 1516 1628 1520
rect 1622 1515 1628 1516
rect 1806 1520 1812 1521
rect 1806 1516 1807 1520
rect 1811 1516 1812 1520
rect 1806 1515 1812 1516
rect 2006 1517 2012 1518
rect 2582 1517 2588 1518
rect 110 1512 116 1513
rect 2006 1513 2007 1517
rect 2011 1513 2012 1517
rect 2006 1512 2012 1513
rect 2046 1516 2052 1517
rect 2046 1512 2047 1516
rect 2051 1512 2052 1516
rect 2582 1513 2583 1517
rect 2587 1513 2588 1517
rect 2582 1512 2588 1513
rect 2742 1517 2748 1518
rect 2742 1513 2743 1517
rect 2747 1513 2748 1517
rect 2742 1512 2748 1513
rect 2902 1517 2908 1518
rect 2902 1513 2903 1517
rect 2907 1513 2908 1517
rect 2902 1512 2908 1513
rect 3062 1517 3068 1518
rect 3062 1513 3063 1517
rect 3067 1513 3068 1517
rect 3062 1512 3068 1513
rect 3222 1517 3228 1518
rect 3222 1513 3223 1517
rect 3227 1513 3228 1517
rect 3222 1512 3228 1513
rect 3382 1517 3388 1518
rect 3382 1513 3383 1517
rect 3387 1513 3388 1517
rect 3382 1512 3388 1513
rect 3542 1517 3548 1518
rect 3542 1513 3543 1517
rect 3547 1513 3548 1517
rect 3542 1512 3548 1513
rect 3702 1517 3708 1518
rect 3702 1513 3703 1517
rect 3707 1513 3708 1517
rect 3702 1512 3708 1513
rect 3942 1516 3948 1517
rect 3942 1512 3943 1516
rect 3947 1512 3948 1516
rect 258 1511 264 1512
rect 258 1510 259 1511
rect 213 1508 259 1510
rect 258 1507 259 1508
rect 263 1507 264 1511
rect 258 1506 264 1507
rect 370 1511 376 1512
rect 370 1507 371 1511
rect 375 1507 376 1511
rect 370 1506 376 1507
rect 390 1511 396 1512
rect 390 1507 391 1511
rect 395 1510 396 1511
rect 762 1511 768 1512
rect 395 1508 529 1510
rect 395 1507 396 1508
rect 390 1506 396 1507
rect 762 1507 763 1511
rect 767 1507 768 1511
rect 762 1506 768 1507
rect 838 1511 844 1512
rect 838 1507 839 1511
rect 843 1510 844 1511
rect 1154 1511 1160 1512
rect 843 1508 929 1510
rect 843 1507 844 1508
rect 838 1506 844 1507
rect 1154 1507 1155 1511
rect 1159 1507 1160 1511
rect 1350 1511 1356 1512
rect 1350 1510 1351 1511
rect 1341 1508 1351 1510
rect 1154 1506 1160 1507
rect 1350 1507 1351 1508
rect 1355 1507 1356 1511
rect 1350 1506 1356 1507
rect 1398 1511 1404 1512
rect 1398 1507 1399 1511
rect 1403 1510 1404 1511
rect 1530 1511 1536 1512
rect 1403 1508 1489 1510
rect 1403 1507 1404 1508
rect 1398 1506 1404 1507
rect 1530 1507 1531 1511
rect 1535 1510 1536 1511
rect 1706 1511 1712 1512
rect 2046 1511 2052 1512
rect 3942 1511 3948 1512
rect 1535 1508 1665 1510
rect 1535 1507 1536 1508
rect 1530 1506 1536 1507
rect 1706 1507 1707 1511
rect 1711 1510 1712 1511
rect 1711 1508 1849 1510
rect 1711 1507 1712 1508
rect 1706 1506 1712 1507
rect 134 1501 140 1502
rect 110 1500 116 1501
rect 110 1496 111 1500
rect 115 1496 116 1500
rect 134 1497 135 1501
rect 139 1497 140 1501
rect 134 1496 140 1497
rect 294 1501 300 1502
rect 294 1497 295 1501
rect 299 1497 300 1501
rect 294 1496 300 1497
rect 486 1501 492 1502
rect 486 1497 487 1501
rect 491 1497 492 1501
rect 486 1496 492 1497
rect 686 1501 692 1502
rect 686 1497 687 1501
rect 691 1497 692 1501
rect 686 1496 692 1497
rect 886 1501 892 1502
rect 886 1497 887 1501
rect 891 1497 892 1501
rect 886 1496 892 1497
rect 1078 1501 1084 1502
rect 1078 1497 1079 1501
rect 1083 1497 1084 1501
rect 1078 1496 1084 1497
rect 1262 1501 1268 1502
rect 1262 1497 1263 1501
rect 1267 1497 1268 1501
rect 1262 1496 1268 1497
rect 1446 1501 1452 1502
rect 1446 1497 1447 1501
rect 1451 1497 1452 1501
rect 1446 1496 1452 1497
rect 1622 1501 1628 1502
rect 1622 1497 1623 1501
rect 1627 1497 1628 1501
rect 1622 1496 1628 1497
rect 1806 1501 1812 1502
rect 1806 1497 1807 1501
rect 1811 1497 1812 1501
rect 1806 1496 1812 1497
rect 2006 1500 2012 1501
rect 2006 1496 2007 1500
rect 2011 1496 2012 1500
rect 110 1495 116 1496
rect 2006 1495 2012 1496
rect 2046 1464 2052 1465
rect 3942 1464 3948 1465
rect 2046 1460 2047 1464
rect 2051 1460 2052 1464
rect 2046 1459 2052 1460
rect 2414 1463 2420 1464
rect 2414 1459 2415 1463
rect 2419 1459 2420 1463
rect 2414 1458 2420 1459
rect 2510 1463 2516 1464
rect 2510 1459 2511 1463
rect 2515 1459 2516 1463
rect 2510 1458 2516 1459
rect 2606 1463 2612 1464
rect 2606 1459 2607 1463
rect 2611 1459 2612 1463
rect 2606 1458 2612 1459
rect 2702 1463 2708 1464
rect 2702 1459 2703 1463
rect 2707 1459 2708 1463
rect 2702 1458 2708 1459
rect 2798 1463 2804 1464
rect 2798 1459 2799 1463
rect 2803 1459 2804 1463
rect 2798 1458 2804 1459
rect 2918 1463 2924 1464
rect 2918 1459 2919 1463
rect 2923 1459 2924 1463
rect 2918 1458 2924 1459
rect 3062 1463 3068 1464
rect 3062 1459 3063 1463
rect 3067 1459 3068 1463
rect 3062 1458 3068 1459
rect 3230 1463 3236 1464
rect 3230 1459 3231 1463
rect 3235 1459 3236 1463
rect 3230 1458 3236 1459
rect 3414 1463 3420 1464
rect 3414 1459 3415 1463
rect 3419 1459 3420 1463
rect 3414 1458 3420 1459
rect 3614 1463 3620 1464
rect 3614 1459 3615 1463
rect 3619 1459 3620 1463
rect 3614 1458 3620 1459
rect 3814 1463 3820 1464
rect 3814 1459 3815 1463
rect 3819 1459 3820 1463
rect 3942 1460 3943 1464
rect 3947 1460 3948 1464
rect 3942 1459 3948 1460
rect 3814 1458 3820 1459
rect 3558 1455 3564 1456
rect 2490 1451 2496 1452
rect 110 1448 116 1449
rect 2006 1448 2012 1449
rect 110 1444 111 1448
rect 115 1444 116 1448
rect 110 1443 116 1444
rect 174 1447 180 1448
rect 174 1443 175 1447
rect 179 1443 180 1447
rect 174 1442 180 1443
rect 358 1447 364 1448
rect 358 1443 359 1447
rect 363 1443 364 1447
rect 358 1442 364 1443
rect 566 1447 572 1448
rect 566 1443 567 1447
rect 571 1443 572 1447
rect 566 1442 572 1443
rect 782 1447 788 1448
rect 782 1443 783 1447
rect 787 1443 788 1447
rect 782 1442 788 1443
rect 1006 1447 1012 1448
rect 1006 1443 1007 1447
rect 1011 1443 1012 1447
rect 1006 1442 1012 1443
rect 1230 1447 1236 1448
rect 1230 1443 1231 1447
rect 1235 1443 1236 1447
rect 1230 1442 1236 1443
rect 1462 1447 1468 1448
rect 1462 1443 1463 1447
rect 1467 1443 1468 1447
rect 1462 1442 1468 1443
rect 1694 1447 1700 1448
rect 1694 1443 1695 1447
rect 1699 1443 1700 1447
rect 1694 1442 1700 1443
rect 1902 1447 1908 1448
rect 1902 1443 1903 1447
rect 1907 1443 1908 1447
rect 2006 1444 2007 1448
rect 2011 1444 2012 1448
rect 2006 1443 2012 1444
rect 2046 1447 2052 1448
rect 2046 1443 2047 1447
rect 2051 1443 2052 1447
rect 2490 1447 2491 1451
rect 2495 1447 2496 1451
rect 2490 1446 2496 1447
rect 2586 1451 2592 1452
rect 2586 1447 2587 1451
rect 2591 1447 2592 1451
rect 2586 1446 2592 1447
rect 2682 1451 2688 1452
rect 2682 1447 2683 1451
rect 2687 1447 2688 1451
rect 2682 1446 2688 1447
rect 2778 1451 2784 1452
rect 2778 1447 2779 1451
rect 2783 1447 2784 1451
rect 2778 1446 2784 1447
rect 2874 1451 2880 1452
rect 2874 1447 2875 1451
rect 2879 1447 2880 1451
rect 2874 1446 2880 1447
rect 2994 1451 3000 1452
rect 2994 1447 2995 1451
rect 2999 1447 3000 1451
rect 2994 1446 3000 1447
rect 3138 1451 3144 1452
rect 3138 1447 3139 1451
rect 3143 1447 3144 1451
rect 3138 1446 3144 1447
rect 3306 1451 3312 1452
rect 3306 1447 3307 1451
rect 3311 1447 3312 1451
rect 3306 1446 3312 1447
rect 3490 1451 3496 1452
rect 3490 1447 3491 1451
rect 3495 1447 3496 1451
rect 3558 1451 3559 1455
rect 3563 1454 3564 1455
rect 3890 1455 3896 1456
rect 3563 1452 3657 1454
rect 3563 1451 3564 1452
rect 3558 1450 3564 1451
rect 3890 1451 3891 1455
rect 3895 1451 3896 1455
rect 3890 1450 3896 1451
rect 3490 1446 3496 1447
rect 3942 1447 3948 1448
rect 1902 1442 1908 1443
rect 2046 1442 2052 1443
rect 2414 1444 2420 1445
rect 2414 1440 2415 1444
rect 2419 1440 2420 1444
rect 250 1439 256 1440
rect 250 1435 251 1439
rect 255 1435 256 1439
rect 250 1434 256 1435
rect 274 1439 280 1440
rect 274 1435 275 1439
rect 279 1438 280 1439
rect 442 1439 448 1440
rect 279 1436 401 1438
rect 279 1435 280 1436
rect 274 1434 280 1435
rect 442 1435 443 1439
rect 447 1438 448 1439
rect 655 1439 661 1440
rect 447 1436 609 1438
rect 447 1435 448 1436
rect 442 1434 448 1435
rect 655 1435 656 1439
rect 660 1438 661 1439
rect 1095 1439 1101 1440
rect 660 1436 825 1438
rect 660 1435 661 1436
rect 655 1434 661 1435
rect 1082 1435 1088 1436
rect 110 1431 116 1432
rect 110 1427 111 1431
rect 115 1427 116 1431
rect 1082 1431 1083 1435
rect 1087 1431 1088 1435
rect 1095 1435 1096 1439
rect 1100 1438 1101 1439
rect 1862 1439 1868 1440
rect 2414 1439 2420 1440
rect 2510 1444 2516 1445
rect 2510 1440 2511 1444
rect 2515 1440 2516 1444
rect 2510 1439 2516 1440
rect 2606 1444 2612 1445
rect 2606 1440 2607 1444
rect 2611 1440 2612 1444
rect 2606 1439 2612 1440
rect 2702 1444 2708 1445
rect 2702 1440 2703 1444
rect 2707 1440 2708 1444
rect 2702 1439 2708 1440
rect 2798 1444 2804 1445
rect 2798 1440 2799 1444
rect 2803 1440 2804 1444
rect 2798 1439 2804 1440
rect 2918 1444 2924 1445
rect 2918 1440 2919 1444
rect 2923 1440 2924 1444
rect 2918 1439 2924 1440
rect 3062 1444 3068 1445
rect 3062 1440 3063 1444
rect 3067 1440 3068 1444
rect 3062 1439 3068 1440
rect 3230 1444 3236 1445
rect 3230 1440 3231 1444
rect 3235 1440 3236 1444
rect 3230 1439 3236 1440
rect 3414 1444 3420 1445
rect 3414 1440 3415 1444
rect 3419 1440 3420 1444
rect 3414 1439 3420 1440
rect 3614 1444 3620 1445
rect 3614 1440 3615 1444
rect 3619 1440 3620 1444
rect 3614 1439 3620 1440
rect 3814 1444 3820 1445
rect 3814 1440 3815 1444
rect 3819 1440 3820 1444
rect 3942 1443 3943 1447
rect 3947 1443 3948 1447
rect 3942 1442 3948 1443
rect 3814 1439 3820 1440
rect 1100 1436 1273 1438
rect 1100 1435 1101 1436
rect 1095 1434 1101 1435
rect 1538 1435 1544 1436
rect 1082 1430 1088 1431
rect 1538 1431 1539 1435
rect 1543 1431 1544 1435
rect 1538 1430 1544 1431
rect 1770 1435 1776 1436
rect 1770 1431 1771 1435
rect 1775 1431 1776 1435
rect 1862 1435 1863 1439
rect 1867 1438 1868 1439
rect 1867 1436 1945 1438
rect 1867 1435 1868 1436
rect 1862 1434 1868 1435
rect 2626 1435 2632 1436
rect 1770 1430 1776 1431
rect 2006 1431 2012 1432
rect 110 1426 116 1427
rect 174 1428 180 1429
rect 174 1424 175 1428
rect 179 1424 180 1428
rect 174 1423 180 1424
rect 358 1428 364 1429
rect 358 1424 359 1428
rect 363 1424 364 1428
rect 358 1423 364 1424
rect 566 1428 572 1429
rect 566 1424 567 1428
rect 571 1424 572 1428
rect 566 1423 572 1424
rect 782 1428 788 1429
rect 782 1424 783 1428
rect 787 1424 788 1428
rect 782 1423 788 1424
rect 1006 1428 1012 1429
rect 1006 1424 1007 1428
rect 1011 1424 1012 1428
rect 1006 1423 1012 1424
rect 1230 1428 1236 1429
rect 1230 1424 1231 1428
rect 1235 1424 1236 1428
rect 1230 1423 1236 1424
rect 1462 1428 1468 1429
rect 1462 1424 1463 1428
rect 1467 1424 1468 1428
rect 1462 1423 1468 1424
rect 1694 1428 1700 1429
rect 1694 1424 1695 1428
rect 1699 1424 1700 1428
rect 1694 1423 1700 1424
rect 1902 1428 1908 1429
rect 1902 1424 1903 1428
rect 1907 1424 1908 1428
rect 2006 1427 2007 1431
rect 2011 1427 2012 1431
rect 2626 1431 2627 1435
rect 2631 1434 2632 1435
rect 3558 1435 3564 1436
rect 3558 1434 3559 1435
rect 2631 1432 3559 1434
rect 2631 1431 2632 1432
rect 2626 1430 2632 1431
rect 3558 1431 3559 1432
rect 3563 1431 3564 1435
rect 3558 1430 3564 1431
rect 2006 1426 2012 1427
rect 1902 1423 1908 1424
rect 2490 1423 2496 1424
rect 2467 1419 2473 1420
rect 2467 1415 2468 1419
rect 2472 1418 2473 1419
rect 2490 1419 2491 1423
rect 2495 1422 2496 1423
rect 2563 1423 2569 1424
rect 2563 1422 2564 1423
rect 2495 1420 2564 1422
rect 2495 1419 2496 1420
rect 2490 1418 2496 1419
rect 2563 1419 2564 1420
rect 2568 1419 2569 1423
rect 2563 1418 2569 1419
rect 2586 1423 2592 1424
rect 2586 1419 2587 1423
rect 2591 1422 2592 1423
rect 2659 1423 2665 1424
rect 2659 1422 2660 1423
rect 2591 1420 2660 1422
rect 2591 1419 2592 1420
rect 2586 1418 2592 1419
rect 2659 1419 2660 1420
rect 2664 1419 2665 1423
rect 2659 1418 2665 1419
rect 2682 1423 2688 1424
rect 2682 1419 2683 1423
rect 2687 1422 2688 1423
rect 2755 1423 2761 1424
rect 2755 1422 2756 1423
rect 2687 1420 2756 1422
rect 2687 1419 2688 1420
rect 2682 1418 2688 1419
rect 2755 1419 2756 1420
rect 2760 1419 2761 1423
rect 2755 1418 2761 1419
rect 2778 1423 2784 1424
rect 2778 1419 2779 1423
rect 2783 1422 2784 1423
rect 2851 1423 2857 1424
rect 2851 1422 2852 1423
rect 2783 1420 2852 1422
rect 2783 1419 2784 1420
rect 2778 1418 2784 1419
rect 2851 1419 2852 1420
rect 2856 1419 2857 1423
rect 2851 1418 2857 1419
rect 2874 1423 2880 1424
rect 2874 1419 2875 1423
rect 2879 1422 2880 1423
rect 2971 1423 2977 1424
rect 2971 1422 2972 1423
rect 2879 1420 2972 1422
rect 2879 1419 2880 1420
rect 2874 1418 2880 1419
rect 2971 1419 2972 1420
rect 2976 1419 2977 1423
rect 2971 1418 2977 1419
rect 2994 1423 3000 1424
rect 2994 1419 2995 1423
rect 2999 1422 3000 1423
rect 3115 1423 3121 1424
rect 3115 1422 3116 1423
rect 2999 1420 3116 1422
rect 2999 1419 3000 1420
rect 2994 1418 3000 1419
rect 3115 1419 3116 1420
rect 3120 1419 3121 1423
rect 3115 1418 3121 1419
rect 3138 1423 3144 1424
rect 3138 1419 3139 1423
rect 3143 1422 3144 1423
rect 3283 1423 3289 1424
rect 3283 1422 3284 1423
rect 3143 1420 3284 1422
rect 3143 1419 3144 1420
rect 3138 1418 3144 1419
rect 3283 1419 3284 1420
rect 3288 1419 3289 1423
rect 3283 1418 3289 1419
rect 3306 1423 3312 1424
rect 3306 1419 3307 1423
rect 3311 1422 3312 1423
rect 3467 1423 3473 1424
rect 3467 1422 3468 1423
rect 3311 1420 3468 1422
rect 3311 1419 3312 1420
rect 3306 1418 3312 1419
rect 3467 1419 3468 1420
rect 3472 1419 3473 1423
rect 3467 1418 3473 1419
rect 3490 1423 3496 1424
rect 3490 1419 3491 1423
rect 3495 1422 3496 1423
rect 3667 1423 3673 1424
rect 3667 1422 3668 1423
rect 3495 1420 3668 1422
rect 3495 1419 3496 1420
rect 3490 1418 3496 1419
rect 3667 1419 3668 1420
rect 3672 1419 3673 1423
rect 3667 1418 3673 1419
rect 3867 1419 3873 1420
rect 2472 1416 2486 1418
rect 2472 1415 2473 1416
rect 2467 1414 2473 1415
rect 2484 1414 2486 1416
rect 3018 1415 3024 1416
rect 3018 1414 3019 1415
rect 2484 1412 3019 1414
rect 3018 1411 3019 1412
rect 3023 1411 3024 1415
rect 3867 1415 3868 1419
rect 3872 1418 3873 1419
rect 3882 1419 3888 1420
rect 3882 1418 3883 1419
rect 3872 1416 3883 1418
rect 3872 1415 3873 1416
rect 3867 1414 3873 1415
rect 3882 1415 3883 1416
rect 3887 1415 3888 1419
rect 3882 1414 3888 1415
rect 3018 1410 3024 1411
rect 227 1407 233 1408
rect 227 1403 228 1407
rect 232 1406 233 1407
rect 274 1407 280 1408
rect 274 1406 275 1407
rect 232 1404 275 1406
rect 232 1403 233 1404
rect 227 1402 233 1403
rect 274 1403 275 1404
rect 279 1403 280 1407
rect 619 1407 625 1408
rect 274 1402 280 1403
rect 402 1403 408 1404
rect 402 1399 403 1403
rect 407 1402 408 1403
rect 411 1403 417 1404
rect 411 1402 412 1403
rect 407 1400 412 1402
rect 407 1399 408 1400
rect 402 1398 408 1399
rect 411 1399 412 1400
rect 416 1399 417 1403
rect 619 1403 620 1407
rect 624 1406 625 1407
rect 655 1407 661 1408
rect 655 1406 656 1407
rect 624 1404 656 1406
rect 624 1403 625 1404
rect 619 1402 625 1403
rect 655 1403 656 1404
rect 660 1403 661 1407
rect 655 1402 661 1403
rect 835 1407 844 1408
rect 835 1403 836 1407
rect 843 1403 844 1407
rect 1082 1407 1088 1408
rect 835 1402 844 1403
rect 930 1403 936 1404
rect 411 1398 417 1399
rect 930 1399 931 1403
rect 935 1402 936 1403
rect 1059 1403 1065 1404
rect 1059 1402 1060 1403
rect 935 1400 1060 1402
rect 935 1399 936 1400
rect 930 1398 936 1399
rect 1059 1399 1060 1400
rect 1064 1399 1065 1403
rect 1082 1403 1083 1407
rect 1087 1406 1088 1407
rect 1283 1407 1289 1408
rect 1283 1406 1284 1407
rect 1087 1404 1284 1406
rect 1087 1403 1088 1404
rect 1082 1402 1088 1403
rect 1283 1403 1284 1404
rect 1288 1403 1289 1407
rect 1538 1407 1544 1408
rect 1283 1402 1289 1403
rect 1515 1403 1521 1404
rect 1059 1398 1065 1399
rect 1515 1399 1516 1403
rect 1520 1402 1521 1403
rect 1538 1403 1539 1407
rect 1543 1406 1544 1407
rect 1747 1407 1753 1408
rect 1747 1406 1748 1407
rect 1543 1404 1748 1406
rect 1543 1403 1544 1404
rect 1538 1402 1544 1403
rect 1747 1403 1748 1404
rect 1752 1403 1753 1407
rect 1747 1402 1753 1403
rect 1770 1407 1776 1408
rect 1770 1403 1771 1407
rect 1775 1406 1776 1407
rect 1955 1407 1961 1408
rect 1955 1406 1956 1407
rect 1775 1404 1956 1406
rect 1775 1403 1776 1404
rect 1770 1402 1776 1403
rect 1955 1403 1956 1404
rect 1960 1403 1961 1407
rect 1955 1402 1961 1403
rect 1520 1400 1534 1402
rect 1520 1399 1521 1400
rect 1515 1398 1521 1399
rect 1532 1398 1534 1400
rect 1666 1399 1672 1400
rect 1666 1398 1667 1399
rect 1532 1396 1667 1398
rect 1666 1395 1667 1396
rect 1671 1395 1672 1399
rect 1666 1394 1672 1395
rect 379 1391 385 1392
rect 379 1387 380 1391
rect 384 1390 385 1391
rect 442 1391 448 1392
rect 442 1390 443 1391
rect 384 1388 443 1390
rect 384 1387 385 1388
rect 379 1386 385 1387
rect 442 1387 443 1388
rect 447 1387 448 1391
rect 442 1386 448 1387
rect 515 1391 524 1392
rect 515 1387 516 1391
rect 523 1387 524 1391
rect 515 1386 524 1387
rect 538 1391 544 1392
rect 538 1387 539 1391
rect 543 1390 544 1391
rect 651 1391 657 1392
rect 651 1390 652 1391
rect 543 1388 652 1390
rect 543 1387 544 1388
rect 538 1386 544 1387
rect 651 1387 652 1388
rect 656 1387 657 1391
rect 651 1386 657 1387
rect 674 1391 680 1392
rect 674 1387 675 1391
rect 679 1390 680 1391
rect 779 1391 785 1392
rect 779 1390 780 1391
rect 679 1388 780 1390
rect 679 1387 680 1388
rect 674 1386 680 1387
rect 779 1387 780 1388
rect 784 1387 785 1391
rect 779 1386 785 1387
rect 802 1391 808 1392
rect 802 1387 803 1391
rect 807 1390 808 1391
rect 907 1391 913 1392
rect 907 1390 908 1391
rect 807 1388 908 1390
rect 807 1387 808 1388
rect 802 1386 808 1387
rect 907 1387 908 1388
rect 912 1387 913 1391
rect 1058 1391 1064 1392
rect 907 1386 913 1387
rect 1035 1389 1041 1390
rect 1035 1385 1036 1389
rect 1040 1385 1041 1389
rect 1058 1387 1059 1391
rect 1063 1390 1064 1391
rect 1171 1391 1177 1392
rect 1171 1390 1172 1391
rect 1063 1388 1172 1390
rect 1063 1387 1064 1388
rect 1058 1386 1064 1387
rect 1171 1387 1172 1388
rect 1176 1387 1177 1391
rect 1171 1386 1177 1387
rect 1194 1391 1200 1392
rect 1194 1387 1195 1391
rect 1199 1390 1200 1391
rect 1315 1391 1321 1392
rect 1315 1390 1316 1391
rect 1199 1388 1316 1390
rect 1199 1387 1200 1388
rect 1194 1386 1200 1387
rect 1315 1387 1316 1388
rect 1320 1387 1321 1391
rect 1315 1386 1321 1387
rect 1338 1391 1344 1392
rect 1338 1387 1339 1391
rect 1343 1390 1344 1391
rect 1475 1391 1481 1392
rect 1475 1390 1476 1391
rect 1343 1388 1476 1390
rect 1343 1387 1344 1388
rect 1338 1386 1344 1387
rect 1475 1387 1476 1388
rect 1480 1387 1481 1391
rect 1803 1391 1809 1392
rect 1475 1386 1481 1387
rect 1635 1389 1641 1390
rect 1035 1384 1041 1385
rect 1635 1385 1636 1389
rect 1640 1385 1641 1389
rect 1803 1387 1804 1391
rect 1808 1390 1809 1391
rect 1834 1391 1840 1392
rect 1834 1390 1835 1391
rect 1808 1388 1835 1390
rect 1808 1387 1809 1388
rect 1803 1386 1809 1387
rect 1834 1387 1835 1388
rect 1839 1387 1840 1391
rect 1834 1386 1840 1387
rect 1955 1391 1961 1392
rect 1955 1387 1956 1391
rect 1960 1390 1961 1391
rect 1986 1391 1992 1392
rect 1986 1390 1987 1391
rect 1960 1388 1987 1390
rect 1960 1387 1961 1388
rect 1955 1386 1961 1387
rect 1986 1387 1987 1388
rect 1991 1387 1992 1391
rect 1986 1386 1992 1387
rect 2123 1387 2129 1388
rect 1635 1384 1641 1385
rect 1036 1382 1038 1384
rect 1095 1383 1101 1384
rect 1095 1382 1096 1383
rect 1036 1380 1096 1382
rect 1095 1379 1096 1380
rect 1100 1379 1101 1383
rect 1095 1378 1101 1379
rect 1402 1383 1408 1384
rect 1402 1379 1403 1383
rect 1407 1382 1408 1383
rect 1636 1382 1638 1384
rect 2123 1383 2124 1387
rect 2128 1386 2129 1387
rect 2154 1387 2160 1388
rect 2154 1386 2155 1387
rect 2128 1384 2155 1386
rect 2128 1383 2129 1384
rect 2123 1382 2129 1383
rect 2154 1383 2155 1384
rect 2159 1383 2160 1387
rect 2154 1382 2160 1383
rect 2310 1387 2316 1388
rect 2310 1383 2311 1387
rect 2315 1386 2316 1387
rect 2355 1387 2361 1388
rect 2355 1386 2356 1387
rect 2315 1384 2356 1386
rect 2315 1383 2316 1384
rect 2310 1382 2316 1383
rect 2355 1383 2356 1384
rect 2360 1383 2361 1387
rect 2355 1382 2361 1383
rect 2611 1387 2617 1388
rect 2611 1383 2612 1387
rect 2616 1386 2617 1387
rect 2626 1387 2632 1388
rect 2626 1386 2627 1387
rect 2616 1384 2627 1386
rect 2616 1383 2617 1384
rect 2611 1382 2617 1383
rect 2626 1383 2627 1384
rect 2631 1383 2632 1387
rect 2626 1382 2632 1383
rect 2634 1387 2640 1388
rect 2634 1383 2635 1387
rect 2639 1386 2640 1387
rect 2859 1387 2865 1388
rect 2859 1386 2860 1387
rect 2639 1384 2860 1386
rect 2639 1383 2640 1384
rect 2634 1382 2640 1383
rect 2859 1383 2860 1384
rect 2864 1383 2865 1387
rect 2859 1382 2865 1383
rect 2882 1387 2888 1388
rect 2882 1383 2883 1387
rect 2887 1386 2888 1387
rect 3107 1387 3113 1388
rect 3107 1386 3108 1387
rect 2887 1384 3108 1386
rect 2887 1383 2888 1384
rect 2882 1382 2888 1383
rect 3107 1383 3108 1384
rect 3112 1383 3113 1387
rect 3107 1382 3113 1383
rect 3130 1387 3136 1388
rect 3130 1383 3131 1387
rect 3135 1386 3136 1387
rect 3355 1387 3361 1388
rect 3355 1386 3356 1387
rect 3135 1384 3356 1386
rect 3135 1383 3136 1384
rect 3130 1382 3136 1383
rect 3355 1383 3356 1384
rect 3360 1383 3361 1387
rect 3355 1382 3361 1383
rect 3378 1387 3384 1388
rect 3378 1383 3379 1387
rect 3383 1386 3384 1387
rect 3611 1387 3617 1388
rect 3611 1386 3612 1387
rect 3383 1384 3612 1386
rect 3383 1383 3384 1384
rect 3378 1382 3384 1383
rect 3611 1383 3612 1384
rect 3616 1383 3617 1387
rect 3611 1382 3617 1383
rect 3867 1387 3873 1388
rect 3867 1383 3868 1387
rect 3872 1386 3873 1387
rect 3906 1387 3912 1388
rect 3906 1386 3907 1387
rect 3872 1384 3907 1386
rect 3872 1383 3873 1384
rect 3867 1382 3873 1383
rect 3906 1383 3907 1384
rect 3911 1383 3912 1387
rect 3906 1382 3912 1383
rect 1407 1380 1638 1382
rect 1407 1379 1408 1380
rect 1402 1378 1408 1379
rect 326 1368 332 1369
rect 110 1365 116 1366
rect 110 1361 111 1365
rect 115 1361 116 1365
rect 326 1364 327 1368
rect 331 1364 332 1368
rect 326 1363 332 1364
rect 462 1368 468 1369
rect 462 1364 463 1368
rect 467 1364 468 1368
rect 462 1363 468 1364
rect 598 1368 604 1369
rect 598 1364 599 1368
rect 603 1364 604 1368
rect 598 1363 604 1364
rect 726 1368 732 1369
rect 726 1364 727 1368
rect 731 1364 732 1368
rect 726 1363 732 1364
rect 854 1368 860 1369
rect 854 1364 855 1368
rect 859 1364 860 1368
rect 854 1363 860 1364
rect 982 1368 988 1369
rect 982 1364 983 1368
rect 987 1364 988 1368
rect 982 1363 988 1364
rect 1118 1368 1124 1369
rect 1118 1364 1119 1368
rect 1123 1364 1124 1368
rect 1118 1363 1124 1364
rect 1262 1368 1268 1369
rect 1262 1364 1263 1368
rect 1267 1364 1268 1368
rect 1262 1363 1268 1364
rect 1422 1368 1428 1369
rect 1422 1364 1423 1368
rect 1427 1364 1428 1368
rect 1422 1363 1428 1364
rect 1582 1368 1588 1369
rect 1582 1364 1583 1368
rect 1587 1364 1588 1368
rect 1582 1363 1588 1364
rect 1750 1368 1756 1369
rect 1750 1364 1751 1368
rect 1755 1364 1756 1368
rect 1750 1363 1756 1364
rect 1902 1368 1908 1369
rect 1902 1364 1903 1368
rect 1907 1364 1908 1368
rect 1902 1363 1908 1364
rect 2006 1365 2012 1366
rect 110 1360 116 1361
rect 2006 1361 2007 1365
rect 2011 1361 2012 1365
rect 2070 1364 2076 1365
rect 2006 1360 2012 1361
rect 2046 1361 2052 1362
rect 402 1359 408 1360
rect 402 1355 403 1359
rect 407 1355 408 1359
rect 402 1354 408 1355
rect 538 1359 544 1360
rect 538 1355 539 1359
rect 543 1355 544 1359
rect 538 1354 544 1355
rect 674 1359 680 1360
rect 674 1355 675 1359
rect 679 1355 680 1359
rect 674 1354 680 1355
rect 802 1359 808 1360
rect 802 1355 803 1359
rect 807 1355 808 1359
rect 802 1354 808 1355
rect 930 1359 936 1360
rect 930 1355 931 1359
rect 935 1355 936 1359
rect 930 1354 936 1355
rect 1058 1359 1064 1360
rect 1058 1355 1059 1359
rect 1063 1355 1064 1359
rect 1058 1354 1064 1355
rect 1194 1359 1200 1360
rect 1194 1355 1195 1359
rect 1199 1355 1200 1359
rect 1194 1354 1200 1355
rect 1338 1359 1344 1360
rect 1338 1355 1339 1359
rect 1343 1355 1344 1359
rect 1650 1359 1656 1360
rect 1338 1354 1344 1355
rect 1348 1356 1465 1358
rect 326 1349 332 1350
rect 110 1348 116 1349
rect 110 1344 111 1348
rect 115 1344 116 1348
rect 326 1345 327 1349
rect 331 1345 332 1349
rect 326 1344 332 1345
rect 462 1349 468 1350
rect 462 1345 463 1349
rect 467 1345 468 1349
rect 462 1344 468 1345
rect 598 1349 604 1350
rect 598 1345 599 1349
rect 603 1345 604 1349
rect 598 1344 604 1345
rect 726 1349 732 1350
rect 726 1345 727 1349
rect 731 1345 732 1349
rect 726 1344 732 1345
rect 854 1349 860 1350
rect 854 1345 855 1349
rect 859 1345 860 1349
rect 854 1344 860 1345
rect 982 1349 988 1350
rect 982 1345 983 1349
rect 987 1345 988 1349
rect 982 1344 988 1345
rect 1118 1349 1124 1350
rect 1118 1345 1119 1349
rect 1123 1345 1124 1349
rect 1118 1344 1124 1345
rect 1262 1349 1268 1350
rect 1262 1345 1263 1349
rect 1267 1345 1268 1349
rect 1262 1344 1268 1345
rect 110 1343 116 1344
rect 1178 1343 1184 1344
rect 1178 1339 1179 1343
rect 1183 1342 1184 1343
rect 1348 1342 1350 1356
rect 1650 1355 1651 1359
rect 1655 1355 1656 1359
rect 1650 1354 1656 1355
rect 1666 1359 1672 1360
rect 1666 1355 1667 1359
rect 1671 1358 1672 1359
rect 1834 1359 1840 1360
rect 1671 1356 1793 1358
rect 1671 1355 1672 1356
rect 1666 1354 1672 1355
rect 1834 1355 1835 1359
rect 1839 1358 1840 1359
rect 1839 1356 1945 1358
rect 2046 1357 2047 1361
rect 2051 1357 2052 1361
rect 2070 1360 2071 1364
rect 2075 1360 2076 1364
rect 2070 1359 2076 1360
rect 2302 1364 2308 1365
rect 2302 1360 2303 1364
rect 2307 1360 2308 1364
rect 2302 1359 2308 1360
rect 2558 1364 2564 1365
rect 2558 1360 2559 1364
rect 2563 1360 2564 1364
rect 2558 1359 2564 1360
rect 2806 1364 2812 1365
rect 2806 1360 2807 1364
rect 2811 1360 2812 1364
rect 2806 1359 2812 1360
rect 3054 1364 3060 1365
rect 3054 1360 3055 1364
rect 3059 1360 3060 1364
rect 3054 1359 3060 1360
rect 3302 1364 3308 1365
rect 3302 1360 3303 1364
rect 3307 1360 3308 1364
rect 3302 1359 3308 1360
rect 3558 1364 3564 1365
rect 3558 1360 3559 1364
rect 3563 1360 3564 1364
rect 3558 1359 3564 1360
rect 3814 1364 3820 1365
rect 3814 1360 3815 1364
rect 3819 1360 3820 1364
rect 3814 1359 3820 1360
rect 3942 1361 3948 1362
rect 2046 1356 2052 1357
rect 3942 1357 3943 1361
rect 3947 1357 3948 1361
rect 3942 1356 3948 1357
rect 1839 1355 1840 1356
rect 1834 1354 1840 1355
rect 1986 1355 1992 1356
rect 1986 1351 1987 1355
rect 1991 1354 1992 1355
rect 2154 1355 2160 1356
rect 1991 1352 2113 1354
rect 1991 1351 1992 1352
rect 1986 1350 1992 1351
rect 2154 1351 2155 1355
rect 2159 1354 2160 1355
rect 2634 1355 2640 1356
rect 2159 1352 2345 1354
rect 2159 1351 2160 1352
rect 2154 1350 2160 1351
rect 2634 1351 2635 1355
rect 2639 1351 2640 1355
rect 2634 1350 2640 1351
rect 2882 1355 2888 1356
rect 2882 1351 2883 1355
rect 2887 1351 2888 1355
rect 2882 1350 2888 1351
rect 3130 1355 3136 1356
rect 3130 1351 3131 1355
rect 3135 1351 3136 1355
rect 3130 1350 3136 1351
rect 3378 1355 3384 1356
rect 3378 1351 3379 1355
rect 3383 1351 3384 1355
rect 3378 1350 3384 1351
rect 3503 1355 3509 1356
rect 3503 1351 3504 1355
rect 3508 1354 3509 1355
rect 3882 1355 3888 1356
rect 3508 1352 3601 1354
rect 3508 1351 3509 1352
rect 3503 1350 3509 1351
rect 3882 1351 3883 1355
rect 3887 1351 3888 1355
rect 3882 1350 3888 1351
rect 1422 1349 1428 1350
rect 1422 1345 1423 1349
rect 1427 1345 1428 1349
rect 1422 1344 1428 1345
rect 1582 1349 1588 1350
rect 1582 1345 1583 1349
rect 1587 1345 1588 1349
rect 1582 1344 1588 1345
rect 1750 1349 1756 1350
rect 1750 1345 1751 1349
rect 1755 1345 1756 1349
rect 1750 1344 1756 1345
rect 1902 1349 1908 1350
rect 1902 1345 1903 1349
rect 1907 1345 1908 1349
rect 1902 1344 1908 1345
rect 2006 1348 2012 1349
rect 2006 1344 2007 1348
rect 2011 1344 2012 1348
rect 2070 1345 2076 1346
rect 2006 1343 2012 1344
rect 2046 1344 2052 1345
rect 1183 1340 1350 1342
rect 2046 1340 2047 1344
rect 2051 1340 2052 1344
rect 2070 1341 2071 1345
rect 2075 1341 2076 1345
rect 2070 1340 2076 1341
rect 2302 1345 2308 1346
rect 2302 1341 2303 1345
rect 2307 1341 2308 1345
rect 2302 1340 2308 1341
rect 2558 1345 2564 1346
rect 2558 1341 2559 1345
rect 2563 1341 2564 1345
rect 2558 1340 2564 1341
rect 2806 1345 2812 1346
rect 2806 1341 2807 1345
rect 2811 1341 2812 1345
rect 2806 1340 2812 1341
rect 3054 1345 3060 1346
rect 3054 1341 3055 1345
rect 3059 1341 3060 1345
rect 3054 1340 3060 1341
rect 3302 1345 3308 1346
rect 3302 1341 3303 1345
rect 3307 1341 3308 1345
rect 3302 1340 3308 1341
rect 3558 1345 3564 1346
rect 3558 1341 3559 1345
rect 3563 1341 3564 1345
rect 3558 1340 3564 1341
rect 3814 1345 3820 1346
rect 3814 1341 3815 1345
rect 3819 1341 3820 1345
rect 3814 1340 3820 1341
rect 3942 1344 3948 1345
rect 3942 1340 3943 1344
rect 3947 1340 3948 1344
rect 1183 1339 1184 1340
rect 2046 1339 2052 1340
rect 3942 1339 3948 1340
rect 1178 1338 1184 1339
rect 3054 1299 3060 1300
rect 3054 1295 3055 1299
rect 3059 1298 3060 1299
rect 3503 1299 3509 1300
rect 3503 1298 3504 1299
rect 3059 1296 3504 1298
rect 3059 1295 3060 1296
rect 3054 1294 3060 1295
rect 3503 1295 3504 1296
rect 3508 1295 3509 1299
rect 3503 1294 3509 1295
rect 110 1288 116 1289
rect 2006 1288 2012 1289
rect 110 1284 111 1288
rect 115 1284 116 1288
rect 110 1283 116 1284
rect 550 1287 556 1288
rect 550 1283 551 1287
rect 555 1283 556 1287
rect 550 1282 556 1283
rect 654 1287 660 1288
rect 654 1283 655 1287
rect 659 1283 660 1287
rect 654 1282 660 1283
rect 766 1287 772 1288
rect 766 1283 767 1287
rect 771 1283 772 1287
rect 766 1282 772 1283
rect 878 1287 884 1288
rect 878 1283 879 1287
rect 883 1283 884 1287
rect 878 1282 884 1283
rect 990 1287 996 1288
rect 990 1283 991 1287
rect 995 1283 996 1287
rect 990 1282 996 1283
rect 1102 1287 1108 1288
rect 1102 1283 1103 1287
rect 1107 1283 1108 1287
rect 1102 1282 1108 1283
rect 1214 1287 1220 1288
rect 1214 1283 1215 1287
rect 1219 1283 1220 1287
rect 1214 1282 1220 1283
rect 1326 1287 1332 1288
rect 1326 1283 1327 1287
rect 1331 1283 1332 1287
rect 1326 1282 1332 1283
rect 1438 1287 1444 1288
rect 1438 1283 1439 1287
rect 1443 1283 1444 1287
rect 1438 1282 1444 1283
rect 1558 1287 1564 1288
rect 1558 1283 1559 1287
rect 1563 1283 1564 1287
rect 2006 1284 2007 1288
rect 2011 1284 2012 1288
rect 2006 1283 2012 1284
rect 2046 1284 2052 1285
rect 3942 1284 3948 1285
rect 1558 1282 1564 1283
rect 2046 1280 2047 1284
rect 2051 1280 2052 1284
rect 962 1279 968 1280
rect 626 1275 632 1276
rect 110 1271 116 1272
rect 110 1267 111 1271
rect 115 1267 116 1271
rect 626 1271 627 1275
rect 631 1271 632 1275
rect 626 1270 632 1271
rect 730 1275 736 1276
rect 730 1271 731 1275
rect 735 1271 736 1275
rect 730 1270 736 1271
rect 842 1275 848 1276
rect 842 1271 843 1275
rect 847 1271 848 1275
rect 842 1270 848 1271
rect 954 1275 960 1276
rect 954 1271 955 1275
rect 959 1271 960 1275
rect 962 1275 963 1279
rect 967 1278 968 1279
rect 1086 1279 1092 1280
rect 967 1276 1033 1278
rect 967 1275 968 1276
rect 962 1274 968 1275
rect 1086 1275 1087 1279
rect 1091 1278 1092 1279
rect 1402 1279 1408 1280
rect 1091 1276 1145 1278
rect 1091 1275 1092 1276
rect 1086 1274 1092 1275
rect 1290 1275 1296 1276
rect 954 1270 960 1271
rect 1290 1271 1291 1275
rect 1295 1271 1296 1275
rect 1402 1275 1403 1279
rect 1407 1275 1408 1279
rect 1526 1279 1532 1280
rect 2046 1279 2052 1280
rect 2070 1283 2076 1284
rect 2070 1279 2071 1283
rect 2075 1279 2076 1283
rect 1402 1274 1408 1275
rect 1514 1275 1520 1276
rect 1290 1270 1296 1271
rect 1514 1271 1515 1275
rect 1519 1271 1520 1275
rect 1526 1275 1527 1279
rect 1531 1278 1532 1279
rect 2070 1278 2076 1279
rect 2222 1283 2228 1284
rect 2222 1279 2223 1283
rect 2227 1279 2228 1283
rect 2222 1278 2228 1279
rect 2414 1283 2420 1284
rect 2414 1279 2415 1283
rect 2419 1279 2420 1283
rect 2414 1278 2420 1279
rect 2614 1283 2620 1284
rect 2614 1279 2615 1283
rect 2619 1279 2620 1283
rect 2614 1278 2620 1279
rect 2814 1283 2820 1284
rect 2814 1279 2815 1283
rect 2819 1279 2820 1283
rect 2814 1278 2820 1279
rect 2998 1283 3004 1284
rect 2998 1279 2999 1283
rect 3003 1279 3004 1283
rect 2998 1278 3004 1279
rect 3174 1283 3180 1284
rect 3174 1279 3175 1283
rect 3179 1279 3180 1283
rect 3174 1278 3180 1279
rect 3342 1283 3348 1284
rect 3342 1279 3343 1283
rect 3347 1279 3348 1283
rect 3342 1278 3348 1279
rect 3502 1283 3508 1284
rect 3502 1279 3503 1283
rect 3507 1279 3508 1283
rect 3502 1278 3508 1279
rect 3662 1283 3668 1284
rect 3662 1279 3663 1283
rect 3667 1279 3668 1283
rect 3662 1278 3668 1279
rect 3830 1283 3836 1284
rect 3830 1279 3831 1283
rect 3835 1279 3836 1283
rect 3942 1280 3943 1284
rect 3947 1280 3948 1284
rect 3942 1279 3948 1280
rect 3830 1278 3836 1279
rect 1531 1276 1601 1278
rect 1531 1275 1532 1276
rect 1526 1274 1532 1275
rect 2310 1275 2316 1276
rect 2310 1274 2311 1275
rect 2301 1272 2311 1274
rect 1514 1270 1520 1271
rect 2006 1271 2012 1272
rect 110 1266 116 1267
rect 550 1268 556 1269
rect 550 1264 551 1268
rect 555 1264 556 1268
rect 550 1263 556 1264
rect 654 1268 660 1269
rect 654 1264 655 1268
rect 659 1264 660 1268
rect 654 1263 660 1264
rect 766 1268 772 1269
rect 766 1264 767 1268
rect 771 1264 772 1268
rect 766 1263 772 1264
rect 878 1268 884 1269
rect 878 1264 879 1268
rect 883 1264 884 1268
rect 878 1263 884 1264
rect 990 1268 996 1269
rect 990 1264 991 1268
rect 995 1264 996 1268
rect 990 1263 996 1264
rect 1102 1268 1108 1269
rect 1102 1264 1103 1268
rect 1107 1264 1108 1268
rect 1102 1263 1108 1264
rect 1214 1268 1220 1269
rect 1214 1264 1215 1268
rect 1219 1264 1220 1268
rect 1214 1263 1220 1264
rect 1326 1268 1332 1269
rect 1326 1264 1327 1268
rect 1331 1264 1332 1268
rect 1326 1263 1332 1264
rect 1438 1268 1444 1269
rect 1438 1264 1439 1268
rect 1443 1264 1444 1268
rect 1438 1263 1444 1264
rect 1558 1268 1564 1269
rect 1558 1264 1559 1268
rect 1563 1264 1564 1268
rect 2006 1267 2007 1271
rect 2011 1267 2012 1271
rect 2146 1271 2152 1272
rect 2006 1266 2012 1267
rect 2046 1267 2052 1268
rect 1558 1263 1564 1264
rect 2046 1263 2047 1267
rect 2051 1263 2052 1267
rect 2146 1267 2147 1271
rect 2151 1267 2152 1271
rect 2310 1271 2311 1272
rect 2315 1271 2316 1275
rect 2310 1270 2316 1271
rect 2358 1275 2364 1276
rect 2358 1271 2359 1275
rect 2363 1274 2364 1275
rect 2698 1275 2704 1276
rect 2363 1272 2457 1274
rect 2363 1271 2364 1272
rect 2358 1270 2364 1271
rect 2690 1271 2696 1272
rect 2146 1266 2152 1267
rect 2690 1267 2691 1271
rect 2695 1267 2696 1271
rect 2698 1271 2699 1275
rect 2703 1274 2704 1275
rect 3906 1275 3912 1276
rect 2703 1272 2857 1274
rect 2703 1271 2704 1272
rect 2698 1270 2704 1271
rect 3074 1271 3080 1272
rect 2690 1266 2696 1267
rect 3074 1267 3075 1271
rect 3079 1267 3080 1271
rect 3074 1266 3080 1267
rect 3250 1271 3256 1272
rect 3250 1267 3251 1271
rect 3255 1267 3256 1271
rect 3250 1266 3256 1267
rect 3418 1271 3424 1272
rect 3418 1267 3419 1271
rect 3423 1267 3424 1271
rect 3418 1266 3424 1267
rect 3578 1271 3584 1272
rect 3578 1267 3579 1271
rect 3583 1267 3584 1271
rect 3578 1266 3584 1267
rect 3738 1271 3744 1272
rect 3738 1267 3739 1271
rect 3743 1267 3744 1271
rect 3906 1271 3907 1275
rect 3911 1271 3912 1275
rect 3906 1270 3912 1271
rect 3738 1266 3744 1267
rect 3942 1267 3948 1268
rect 2046 1262 2052 1263
rect 2070 1264 2076 1265
rect 2070 1260 2071 1264
rect 2075 1260 2076 1264
rect 2070 1259 2076 1260
rect 2222 1264 2228 1265
rect 2222 1260 2223 1264
rect 2227 1260 2228 1264
rect 2222 1259 2228 1260
rect 2414 1264 2420 1265
rect 2414 1260 2415 1264
rect 2419 1260 2420 1264
rect 2414 1259 2420 1260
rect 2614 1264 2620 1265
rect 2614 1260 2615 1264
rect 2619 1260 2620 1264
rect 2614 1259 2620 1260
rect 2814 1264 2820 1265
rect 2814 1260 2815 1264
rect 2819 1260 2820 1264
rect 2814 1259 2820 1260
rect 2998 1264 3004 1265
rect 2998 1260 2999 1264
rect 3003 1260 3004 1264
rect 2998 1259 3004 1260
rect 3174 1264 3180 1265
rect 3174 1260 3175 1264
rect 3179 1260 3180 1264
rect 3174 1259 3180 1260
rect 3342 1264 3348 1265
rect 3342 1260 3343 1264
rect 3347 1260 3348 1264
rect 3342 1259 3348 1260
rect 3502 1264 3508 1265
rect 3502 1260 3503 1264
rect 3507 1260 3508 1264
rect 3502 1259 3508 1260
rect 3662 1264 3668 1265
rect 3662 1260 3663 1264
rect 3667 1260 3668 1264
rect 3662 1259 3668 1260
rect 3830 1264 3836 1265
rect 3830 1260 3831 1264
rect 3835 1260 3836 1264
rect 3942 1263 3943 1267
rect 3947 1263 3948 1267
rect 3942 1262 3948 1263
rect 3830 1259 3836 1260
rect 2358 1251 2364 1252
rect 2358 1250 2359 1251
rect 2140 1248 2359 1250
rect 626 1247 632 1248
rect 603 1243 609 1244
rect 603 1239 604 1243
rect 608 1242 609 1243
rect 626 1243 627 1247
rect 631 1246 632 1247
rect 707 1247 713 1248
rect 707 1246 708 1247
rect 631 1244 708 1246
rect 631 1243 632 1244
rect 626 1242 632 1243
rect 707 1243 708 1244
rect 712 1243 713 1247
rect 707 1242 713 1243
rect 730 1247 736 1248
rect 730 1243 731 1247
rect 735 1246 736 1247
rect 819 1247 825 1248
rect 819 1246 820 1247
rect 735 1244 820 1246
rect 735 1243 736 1244
rect 730 1242 736 1243
rect 819 1243 820 1244
rect 824 1243 825 1247
rect 819 1242 825 1243
rect 842 1247 848 1248
rect 842 1243 843 1247
rect 847 1246 848 1247
rect 931 1247 937 1248
rect 931 1246 932 1247
rect 847 1244 932 1246
rect 847 1243 848 1244
rect 842 1242 848 1243
rect 931 1243 932 1244
rect 936 1243 937 1247
rect 931 1242 937 1243
rect 954 1247 960 1248
rect 954 1243 955 1247
rect 959 1246 960 1247
rect 1043 1247 1049 1248
rect 1043 1246 1044 1247
rect 959 1244 1044 1246
rect 959 1243 960 1244
rect 954 1242 960 1243
rect 1043 1243 1044 1244
rect 1048 1243 1049 1247
rect 1043 1242 1049 1243
rect 1155 1247 1161 1248
rect 1155 1243 1156 1247
rect 1160 1246 1161 1247
rect 1178 1247 1184 1248
rect 1178 1246 1179 1247
rect 1160 1244 1179 1246
rect 1160 1243 1161 1244
rect 1155 1242 1161 1243
rect 1178 1243 1179 1244
rect 1183 1243 1184 1247
rect 1290 1247 1296 1248
rect 1178 1242 1184 1243
rect 1186 1243 1192 1244
rect 608 1240 622 1242
rect 608 1239 609 1240
rect 603 1238 609 1239
rect 620 1238 622 1240
rect 938 1239 944 1240
rect 938 1238 939 1239
rect 620 1236 939 1238
rect 938 1235 939 1236
rect 943 1235 944 1239
rect 1186 1239 1187 1243
rect 1191 1242 1192 1243
rect 1267 1243 1273 1244
rect 1267 1242 1268 1243
rect 1191 1240 1268 1242
rect 1191 1239 1192 1240
rect 1186 1238 1192 1239
rect 1267 1239 1268 1240
rect 1272 1239 1273 1243
rect 1290 1243 1291 1247
rect 1295 1246 1296 1247
rect 1379 1247 1385 1248
rect 1379 1246 1380 1247
rect 1295 1244 1380 1246
rect 1295 1243 1296 1244
rect 1290 1242 1296 1243
rect 1379 1243 1380 1244
rect 1384 1243 1385 1247
rect 1379 1242 1385 1243
rect 1491 1247 1497 1248
rect 1491 1243 1492 1247
rect 1496 1246 1497 1247
rect 1526 1247 1532 1248
rect 1526 1246 1527 1247
rect 1496 1244 1527 1246
rect 1496 1243 1497 1244
rect 1491 1242 1497 1243
rect 1526 1243 1527 1244
rect 1531 1243 1532 1247
rect 1526 1242 1532 1243
rect 1611 1247 1617 1248
rect 1611 1243 1612 1247
rect 1616 1246 1617 1247
rect 1650 1247 1656 1248
rect 1650 1246 1651 1247
rect 1616 1244 1651 1246
rect 1616 1243 1617 1244
rect 1611 1242 1617 1243
rect 1650 1243 1651 1244
rect 1655 1243 1656 1247
rect 1650 1242 1656 1243
rect 2123 1243 2129 1244
rect 1267 1238 1273 1239
rect 2123 1239 2124 1243
rect 2128 1242 2129 1243
rect 2140 1242 2142 1248
rect 2358 1247 2359 1248
rect 2363 1247 2364 1251
rect 2698 1251 2704 1252
rect 2698 1250 2699 1251
rect 2358 1246 2364 1247
rect 2548 1248 2699 1250
rect 2128 1240 2142 1242
rect 2146 1243 2152 1244
rect 2128 1239 2129 1240
rect 2123 1238 2129 1239
rect 2146 1239 2147 1243
rect 2151 1242 2152 1243
rect 2275 1243 2281 1244
rect 2275 1242 2276 1243
rect 2151 1240 2276 1242
rect 2151 1239 2152 1240
rect 2146 1238 2152 1239
rect 2275 1239 2276 1240
rect 2280 1239 2281 1243
rect 2275 1238 2281 1239
rect 2467 1243 2473 1244
rect 2467 1239 2468 1243
rect 2472 1242 2473 1243
rect 2548 1242 2550 1248
rect 2698 1247 2699 1248
rect 2703 1247 2704 1251
rect 2698 1246 2704 1247
rect 2472 1240 2550 1242
rect 2690 1243 2696 1244
rect 2472 1239 2473 1240
rect 2467 1238 2473 1239
rect 2578 1239 2584 1240
rect 938 1234 944 1235
rect 2578 1235 2579 1239
rect 2583 1238 2584 1239
rect 2667 1239 2673 1240
rect 2667 1238 2668 1239
rect 2583 1236 2668 1238
rect 2583 1235 2584 1236
rect 2578 1234 2584 1235
rect 2667 1235 2668 1236
rect 2672 1235 2673 1239
rect 2690 1239 2691 1243
rect 2695 1242 2696 1243
rect 2867 1243 2873 1244
rect 2867 1242 2868 1243
rect 2695 1240 2868 1242
rect 2695 1239 2696 1240
rect 2690 1238 2696 1239
rect 2867 1239 2868 1240
rect 2872 1239 2873 1243
rect 2867 1238 2873 1239
rect 3051 1243 3060 1244
rect 3051 1239 3052 1243
rect 3059 1239 3060 1243
rect 3051 1238 3060 1239
rect 3074 1243 3080 1244
rect 3074 1239 3075 1243
rect 3079 1242 3080 1243
rect 3227 1243 3233 1244
rect 3227 1242 3228 1243
rect 3079 1240 3228 1242
rect 3079 1239 3080 1240
rect 3074 1238 3080 1239
rect 3227 1239 3228 1240
rect 3232 1239 3233 1243
rect 3227 1238 3233 1239
rect 3250 1243 3256 1244
rect 3250 1239 3251 1243
rect 3255 1242 3256 1243
rect 3395 1243 3401 1244
rect 3395 1242 3396 1243
rect 3255 1240 3396 1242
rect 3255 1239 3256 1240
rect 3250 1238 3256 1239
rect 3395 1239 3396 1240
rect 3400 1239 3401 1243
rect 3395 1238 3401 1239
rect 3418 1243 3424 1244
rect 3418 1239 3419 1243
rect 3423 1242 3424 1243
rect 3555 1243 3561 1244
rect 3555 1242 3556 1243
rect 3423 1240 3556 1242
rect 3423 1239 3424 1240
rect 3418 1238 3424 1239
rect 3555 1239 3556 1240
rect 3560 1239 3561 1243
rect 3555 1238 3561 1239
rect 3578 1243 3584 1244
rect 3578 1239 3579 1243
rect 3583 1242 3584 1243
rect 3715 1243 3721 1244
rect 3715 1242 3716 1243
rect 3583 1240 3716 1242
rect 3583 1239 3584 1240
rect 3578 1238 3584 1239
rect 3715 1239 3716 1240
rect 3720 1239 3721 1243
rect 3715 1238 3721 1239
rect 3883 1239 3889 1240
rect 2667 1234 2673 1235
rect 3883 1235 3884 1239
rect 3888 1238 3889 1239
rect 3906 1239 3912 1240
rect 3906 1238 3907 1239
rect 3888 1236 3907 1238
rect 3888 1235 3889 1236
rect 3883 1234 3889 1235
rect 3906 1235 3907 1236
rect 3911 1235 3912 1239
rect 3906 1234 3912 1235
rect 466 1231 472 1232
rect 443 1229 449 1230
rect 443 1225 444 1229
rect 448 1225 449 1229
rect 466 1227 467 1231
rect 471 1230 472 1231
rect 571 1231 577 1232
rect 571 1230 572 1231
rect 471 1228 572 1230
rect 471 1227 472 1228
rect 466 1226 472 1227
rect 571 1227 572 1228
rect 576 1227 577 1231
rect 571 1226 577 1227
rect 594 1231 600 1232
rect 594 1227 595 1231
rect 599 1230 600 1231
rect 715 1231 721 1232
rect 715 1230 716 1231
rect 599 1228 716 1230
rect 599 1227 600 1228
rect 594 1226 600 1227
rect 715 1227 716 1228
rect 720 1227 721 1231
rect 715 1226 721 1227
rect 738 1231 744 1232
rect 738 1227 739 1231
rect 743 1230 744 1231
rect 859 1231 865 1232
rect 859 1230 860 1231
rect 743 1228 860 1230
rect 743 1227 744 1228
rect 738 1226 744 1227
rect 859 1227 860 1228
rect 864 1227 865 1231
rect 859 1226 865 1227
rect 927 1231 933 1232
rect 927 1227 928 1231
rect 932 1230 933 1231
rect 1011 1231 1017 1232
rect 1011 1230 1012 1231
rect 932 1228 1012 1230
rect 932 1227 933 1228
rect 927 1226 933 1227
rect 1011 1227 1012 1228
rect 1016 1227 1017 1231
rect 1011 1226 1017 1227
rect 1163 1231 1169 1232
rect 1163 1227 1164 1231
rect 1168 1230 1169 1231
rect 1194 1231 1200 1232
rect 1194 1230 1195 1231
rect 1168 1228 1195 1230
rect 1168 1227 1169 1228
rect 1163 1226 1169 1227
rect 1194 1227 1195 1228
rect 1199 1227 1200 1231
rect 1194 1226 1200 1227
rect 1282 1231 1288 1232
rect 1282 1227 1283 1231
rect 1287 1230 1288 1231
rect 1307 1231 1313 1232
rect 1307 1230 1308 1231
rect 1287 1228 1308 1230
rect 1287 1227 1288 1228
rect 1282 1226 1288 1227
rect 1307 1227 1308 1228
rect 1312 1227 1313 1231
rect 1307 1226 1313 1227
rect 1459 1231 1465 1232
rect 1459 1227 1460 1231
rect 1464 1230 1465 1231
rect 1514 1231 1520 1232
rect 1514 1230 1515 1231
rect 1464 1228 1515 1230
rect 1464 1227 1465 1228
rect 1459 1226 1465 1227
rect 1514 1227 1515 1228
rect 1519 1227 1520 1231
rect 1514 1226 1520 1227
rect 1527 1231 1533 1232
rect 1527 1227 1528 1231
rect 1532 1230 1533 1231
rect 1611 1231 1617 1232
rect 1611 1230 1612 1231
rect 1532 1228 1612 1230
rect 1532 1227 1533 1228
rect 1527 1226 1533 1227
rect 1611 1227 1612 1228
rect 1616 1227 1617 1231
rect 1611 1226 1617 1227
rect 1634 1231 1640 1232
rect 1634 1227 1635 1231
rect 1639 1230 1640 1231
rect 1763 1231 1769 1232
rect 1763 1230 1764 1231
rect 1639 1228 1764 1230
rect 1639 1227 1640 1228
rect 1634 1226 1640 1227
rect 1763 1227 1764 1228
rect 1768 1227 1769 1231
rect 1763 1226 1769 1227
rect 443 1224 449 1225
rect 444 1222 446 1224
rect 798 1223 804 1224
rect 798 1222 799 1223
rect 444 1220 799 1222
rect 798 1219 799 1220
rect 803 1219 804 1223
rect 798 1218 804 1219
rect 2210 1219 2216 1220
rect 2187 1217 2193 1218
rect 2187 1213 2188 1217
rect 2192 1213 2193 1217
rect 2210 1215 2211 1219
rect 2215 1218 2216 1219
rect 2363 1219 2369 1220
rect 2363 1218 2364 1219
rect 2215 1216 2364 1218
rect 2215 1215 2216 1216
rect 2210 1214 2216 1215
rect 2363 1215 2364 1216
rect 2368 1215 2369 1219
rect 2363 1214 2369 1215
rect 2386 1219 2392 1220
rect 2386 1215 2387 1219
rect 2391 1218 2392 1219
rect 2555 1219 2561 1220
rect 2555 1218 2556 1219
rect 2391 1216 2556 1218
rect 2391 1215 2392 1216
rect 2386 1214 2392 1215
rect 2555 1215 2556 1216
rect 2560 1215 2561 1219
rect 2555 1214 2561 1215
rect 2747 1219 2753 1220
rect 2747 1215 2748 1219
rect 2752 1218 2753 1219
rect 2791 1219 2797 1220
rect 2791 1218 2792 1219
rect 2752 1216 2792 1218
rect 2752 1215 2753 1216
rect 2747 1214 2753 1215
rect 2791 1215 2792 1216
rect 2796 1215 2797 1219
rect 2791 1214 2797 1215
rect 2914 1219 2920 1220
rect 2914 1215 2915 1219
rect 2919 1218 2920 1219
rect 2939 1219 2945 1220
rect 2939 1218 2940 1219
rect 2919 1216 2940 1218
rect 2919 1215 2920 1216
rect 2914 1214 2920 1215
rect 2939 1215 2940 1216
rect 2944 1215 2945 1219
rect 3146 1219 3152 1220
rect 2939 1214 2945 1215
rect 3123 1217 3129 1218
rect 2187 1212 2193 1213
rect 3123 1213 3124 1217
rect 3128 1213 3129 1217
rect 3146 1215 3147 1219
rect 3151 1218 3152 1219
rect 3291 1219 3297 1220
rect 3291 1218 3292 1219
rect 3151 1216 3292 1218
rect 3151 1215 3152 1216
rect 3146 1214 3152 1215
rect 3291 1215 3292 1216
rect 3296 1215 3297 1219
rect 3291 1214 3297 1215
rect 3314 1219 3320 1220
rect 3314 1215 3315 1219
rect 3319 1218 3320 1219
rect 3451 1219 3457 1220
rect 3451 1218 3452 1219
rect 3319 1216 3452 1218
rect 3319 1215 3320 1216
rect 3314 1214 3320 1215
rect 3451 1215 3452 1216
rect 3456 1215 3457 1219
rect 3451 1214 3457 1215
rect 3603 1219 3609 1220
rect 3603 1215 3604 1219
rect 3608 1218 3609 1219
rect 3639 1219 3645 1220
rect 3639 1218 3640 1219
rect 3608 1216 3640 1218
rect 3608 1215 3609 1216
rect 3603 1214 3609 1215
rect 3639 1215 3640 1216
rect 3644 1215 3645 1219
rect 3639 1214 3645 1215
rect 3738 1219 3744 1220
rect 3738 1215 3739 1219
rect 3743 1218 3744 1219
rect 3755 1219 3761 1220
rect 3755 1218 3756 1219
rect 3743 1216 3756 1218
rect 3743 1215 3744 1216
rect 3738 1214 3744 1215
rect 3755 1215 3756 1216
rect 3760 1215 3761 1219
rect 3755 1214 3761 1215
rect 3891 1219 3897 1220
rect 3891 1215 3892 1219
rect 3896 1218 3897 1219
rect 3914 1219 3920 1220
rect 3914 1218 3915 1219
rect 3896 1216 3915 1218
rect 3896 1215 3897 1216
rect 3891 1214 3897 1215
rect 3914 1215 3915 1216
rect 3919 1215 3920 1219
rect 3914 1214 3920 1215
rect 3123 1212 3129 1213
rect 2188 1210 2190 1212
rect 2658 1211 2664 1212
rect 2658 1210 2659 1211
rect 390 1208 396 1209
rect 110 1205 116 1206
rect 110 1201 111 1205
rect 115 1201 116 1205
rect 390 1204 391 1208
rect 395 1204 396 1208
rect 390 1203 396 1204
rect 518 1208 524 1209
rect 518 1204 519 1208
rect 523 1204 524 1208
rect 518 1203 524 1204
rect 662 1208 668 1209
rect 662 1204 663 1208
rect 667 1204 668 1208
rect 662 1203 668 1204
rect 806 1208 812 1209
rect 806 1204 807 1208
rect 811 1204 812 1208
rect 806 1203 812 1204
rect 958 1208 964 1209
rect 958 1204 959 1208
rect 963 1204 964 1208
rect 958 1203 964 1204
rect 1110 1208 1116 1209
rect 1110 1204 1111 1208
rect 1115 1204 1116 1208
rect 1110 1203 1116 1204
rect 1254 1208 1260 1209
rect 1254 1204 1255 1208
rect 1259 1204 1260 1208
rect 1254 1203 1260 1204
rect 1406 1208 1412 1209
rect 1406 1204 1407 1208
rect 1411 1204 1412 1208
rect 1406 1203 1412 1204
rect 1558 1208 1564 1209
rect 1558 1204 1559 1208
rect 1563 1204 1564 1208
rect 1558 1203 1564 1204
rect 1710 1208 1716 1209
rect 2188 1208 2659 1210
rect 1710 1204 1711 1208
rect 1715 1204 1716 1208
rect 2658 1207 2659 1208
rect 2663 1207 2664 1211
rect 3124 1210 3126 1212
rect 3498 1211 3504 1212
rect 3498 1210 3499 1211
rect 3124 1208 3499 1210
rect 2658 1206 2664 1207
rect 3498 1207 3499 1208
rect 3503 1207 3504 1211
rect 3498 1206 3504 1207
rect 1710 1203 1716 1204
rect 2006 1205 2012 1206
rect 110 1200 116 1201
rect 2006 1201 2007 1205
rect 2011 1201 2012 1205
rect 2006 1200 2012 1201
rect 466 1199 472 1200
rect 466 1195 467 1199
rect 471 1195 472 1199
rect 466 1194 472 1195
rect 594 1199 600 1200
rect 594 1195 595 1199
rect 599 1195 600 1199
rect 594 1194 600 1195
rect 738 1199 744 1200
rect 738 1195 739 1199
rect 743 1195 744 1199
rect 927 1199 933 1200
rect 927 1198 928 1199
rect 885 1196 928 1198
rect 738 1194 744 1195
rect 927 1195 928 1196
rect 932 1195 933 1199
rect 927 1194 933 1195
rect 938 1199 944 1200
rect 938 1195 939 1199
rect 943 1198 944 1199
rect 1186 1199 1192 1200
rect 943 1196 1001 1198
rect 943 1195 944 1196
rect 938 1194 944 1195
rect 1186 1195 1187 1199
rect 1191 1195 1192 1199
rect 1186 1194 1192 1195
rect 1194 1199 1200 1200
rect 1194 1195 1195 1199
rect 1199 1198 1200 1199
rect 1527 1199 1533 1200
rect 1527 1198 1528 1199
rect 1199 1196 1297 1198
rect 1485 1196 1528 1198
rect 1199 1195 1200 1196
rect 1194 1194 1200 1195
rect 1527 1195 1528 1196
rect 1532 1195 1533 1199
rect 1527 1194 1533 1195
rect 1634 1199 1640 1200
rect 1634 1195 1635 1199
rect 1639 1195 1640 1199
rect 1634 1194 1640 1195
rect 1662 1199 1668 1200
rect 1662 1195 1663 1199
rect 1667 1198 1668 1199
rect 1667 1196 1753 1198
rect 2134 1196 2140 1197
rect 1667 1195 1668 1196
rect 1662 1194 1668 1195
rect 2046 1193 2052 1194
rect 390 1189 396 1190
rect 110 1188 116 1189
rect 110 1184 111 1188
rect 115 1184 116 1188
rect 390 1185 391 1189
rect 395 1185 396 1189
rect 390 1184 396 1185
rect 518 1189 524 1190
rect 518 1185 519 1189
rect 523 1185 524 1189
rect 518 1184 524 1185
rect 662 1189 668 1190
rect 662 1185 663 1189
rect 667 1185 668 1189
rect 662 1184 668 1185
rect 806 1189 812 1190
rect 806 1185 807 1189
rect 811 1185 812 1189
rect 806 1184 812 1185
rect 958 1189 964 1190
rect 958 1185 959 1189
rect 963 1185 964 1189
rect 958 1184 964 1185
rect 1110 1189 1116 1190
rect 1110 1185 1111 1189
rect 1115 1185 1116 1189
rect 1110 1184 1116 1185
rect 1254 1189 1260 1190
rect 1254 1185 1255 1189
rect 1259 1185 1260 1189
rect 1254 1184 1260 1185
rect 1406 1189 1412 1190
rect 1406 1185 1407 1189
rect 1411 1185 1412 1189
rect 1406 1184 1412 1185
rect 1558 1189 1564 1190
rect 1558 1185 1559 1189
rect 1563 1185 1564 1189
rect 1558 1184 1564 1185
rect 1710 1189 1716 1190
rect 2046 1189 2047 1193
rect 2051 1189 2052 1193
rect 2134 1192 2135 1196
rect 2139 1192 2140 1196
rect 2134 1191 2140 1192
rect 2310 1196 2316 1197
rect 2310 1192 2311 1196
rect 2315 1192 2316 1196
rect 2310 1191 2316 1192
rect 2502 1196 2508 1197
rect 2502 1192 2503 1196
rect 2507 1192 2508 1196
rect 2502 1191 2508 1192
rect 2694 1196 2700 1197
rect 2694 1192 2695 1196
rect 2699 1192 2700 1196
rect 2694 1191 2700 1192
rect 2886 1196 2892 1197
rect 2886 1192 2887 1196
rect 2891 1192 2892 1196
rect 2886 1191 2892 1192
rect 3070 1196 3076 1197
rect 3070 1192 3071 1196
rect 3075 1192 3076 1196
rect 3070 1191 3076 1192
rect 3238 1196 3244 1197
rect 3238 1192 3239 1196
rect 3243 1192 3244 1196
rect 3238 1191 3244 1192
rect 3398 1196 3404 1197
rect 3398 1192 3399 1196
rect 3403 1192 3404 1196
rect 3398 1191 3404 1192
rect 3550 1196 3556 1197
rect 3550 1192 3551 1196
rect 3555 1192 3556 1196
rect 3550 1191 3556 1192
rect 3702 1196 3708 1197
rect 3702 1192 3703 1196
rect 3707 1192 3708 1196
rect 3702 1191 3708 1192
rect 3838 1196 3844 1197
rect 3838 1192 3839 1196
rect 3843 1192 3844 1196
rect 3838 1191 3844 1192
rect 3942 1193 3948 1194
rect 1710 1185 1711 1189
rect 1715 1185 1716 1189
rect 1710 1184 1716 1185
rect 2006 1188 2012 1189
rect 2046 1188 2052 1189
rect 3942 1189 3943 1193
rect 3947 1189 3948 1193
rect 3942 1188 3948 1189
rect 2006 1184 2007 1188
rect 2011 1184 2012 1188
rect 110 1183 116 1184
rect 2006 1183 2012 1184
rect 2210 1187 2216 1188
rect 2210 1183 2211 1187
rect 2215 1183 2216 1187
rect 2210 1182 2216 1183
rect 2386 1187 2392 1188
rect 2386 1183 2387 1187
rect 2391 1183 2392 1187
rect 2386 1182 2392 1183
rect 2578 1187 2584 1188
rect 2578 1183 2579 1187
rect 2583 1183 2584 1187
rect 2578 1182 2584 1183
rect 2658 1187 2664 1188
rect 2658 1183 2659 1187
rect 2663 1186 2664 1187
rect 2791 1187 2797 1188
rect 2663 1184 2737 1186
rect 2663 1183 2664 1184
rect 2658 1182 2664 1183
rect 2791 1183 2792 1187
rect 2796 1186 2797 1187
rect 3146 1187 3152 1188
rect 2796 1184 2929 1186
rect 2796 1183 2797 1184
rect 2791 1182 2797 1183
rect 3146 1183 3147 1187
rect 3151 1183 3152 1187
rect 3146 1182 3152 1183
rect 3314 1187 3320 1188
rect 3314 1183 3315 1187
rect 3319 1183 3320 1187
rect 3314 1182 3320 1183
rect 3474 1187 3480 1188
rect 3474 1183 3475 1187
rect 3479 1183 3480 1187
rect 3474 1182 3480 1183
rect 3498 1187 3504 1188
rect 3498 1183 3499 1187
rect 3503 1186 3504 1187
rect 3639 1187 3645 1188
rect 3503 1184 3593 1186
rect 3503 1183 3504 1184
rect 3498 1182 3504 1183
rect 3639 1183 3640 1187
rect 3644 1186 3645 1187
rect 3906 1187 3912 1188
rect 3644 1184 3745 1186
rect 3644 1183 3645 1184
rect 3639 1182 3645 1183
rect 3906 1183 3907 1187
rect 3911 1183 3912 1187
rect 3906 1182 3912 1183
rect 2134 1177 2140 1178
rect 2046 1176 2052 1177
rect 2046 1172 2047 1176
rect 2051 1172 2052 1176
rect 2134 1173 2135 1177
rect 2139 1173 2140 1177
rect 2134 1172 2140 1173
rect 2310 1177 2316 1178
rect 2310 1173 2311 1177
rect 2315 1173 2316 1177
rect 2310 1172 2316 1173
rect 2502 1177 2508 1178
rect 2502 1173 2503 1177
rect 2507 1173 2508 1177
rect 2502 1172 2508 1173
rect 2694 1177 2700 1178
rect 2694 1173 2695 1177
rect 2699 1173 2700 1177
rect 2694 1172 2700 1173
rect 2886 1177 2892 1178
rect 2886 1173 2887 1177
rect 2891 1173 2892 1177
rect 2886 1172 2892 1173
rect 3070 1177 3076 1178
rect 3070 1173 3071 1177
rect 3075 1173 3076 1177
rect 3070 1172 3076 1173
rect 3238 1177 3244 1178
rect 3238 1173 3239 1177
rect 3243 1173 3244 1177
rect 3238 1172 3244 1173
rect 3398 1177 3404 1178
rect 3398 1173 3399 1177
rect 3403 1173 3404 1177
rect 3398 1172 3404 1173
rect 3550 1177 3556 1178
rect 3550 1173 3551 1177
rect 3555 1173 3556 1177
rect 3550 1172 3556 1173
rect 3702 1177 3708 1178
rect 3702 1173 3703 1177
rect 3707 1173 3708 1177
rect 3702 1172 3708 1173
rect 3838 1177 3844 1178
rect 3838 1173 3839 1177
rect 3843 1173 3844 1177
rect 3838 1172 3844 1173
rect 3942 1176 3948 1177
rect 3942 1172 3943 1176
rect 3947 1172 3948 1176
rect 2046 1171 2052 1172
rect 3942 1171 3948 1172
rect 110 1132 116 1133
rect 2006 1132 2012 1133
rect 110 1128 111 1132
rect 115 1128 116 1132
rect 110 1127 116 1128
rect 174 1131 180 1132
rect 174 1127 175 1131
rect 179 1127 180 1131
rect 174 1126 180 1127
rect 326 1131 332 1132
rect 326 1127 327 1131
rect 331 1127 332 1131
rect 326 1126 332 1127
rect 494 1131 500 1132
rect 494 1127 495 1131
rect 499 1127 500 1131
rect 494 1126 500 1127
rect 670 1131 676 1132
rect 670 1127 671 1131
rect 675 1127 676 1131
rect 670 1126 676 1127
rect 846 1131 852 1132
rect 846 1127 847 1131
rect 851 1127 852 1131
rect 846 1126 852 1127
rect 1030 1131 1036 1132
rect 1030 1127 1031 1131
rect 1035 1127 1036 1131
rect 1030 1126 1036 1127
rect 1206 1131 1212 1132
rect 1206 1127 1207 1131
rect 1211 1127 1212 1131
rect 1206 1126 1212 1127
rect 1382 1131 1388 1132
rect 1382 1127 1383 1131
rect 1387 1127 1388 1131
rect 1382 1126 1388 1127
rect 1566 1131 1572 1132
rect 1566 1127 1567 1131
rect 1571 1127 1572 1131
rect 1566 1126 1572 1127
rect 1750 1131 1756 1132
rect 1750 1127 1751 1131
rect 1755 1127 1756 1131
rect 2006 1128 2007 1132
rect 2011 1128 2012 1132
rect 2006 1127 2012 1128
rect 1750 1126 1756 1127
rect 798 1123 804 1124
rect 250 1119 256 1120
rect 110 1115 116 1116
rect 110 1111 111 1115
rect 115 1111 116 1115
rect 250 1115 251 1119
rect 255 1115 256 1119
rect 250 1114 256 1115
rect 402 1119 408 1120
rect 402 1115 403 1119
rect 407 1115 408 1119
rect 402 1114 408 1115
rect 570 1119 576 1120
rect 570 1115 571 1119
rect 575 1115 576 1119
rect 570 1114 576 1115
rect 746 1119 752 1120
rect 746 1115 747 1119
rect 751 1115 752 1119
rect 798 1119 799 1123
rect 803 1122 804 1123
rect 1282 1123 1288 1124
rect 803 1120 889 1122
rect 803 1119 804 1120
rect 798 1118 804 1119
rect 1106 1119 1112 1120
rect 746 1114 752 1115
rect 1106 1115 1107 1119
rect 1111 1115 1112 1119
rect 1282 1119 1283 1123
rect 1287 1119 1288 1123
rect 1282 1118 1288 1119
rect 1326 1123 1332 1124
rect 1326 1119 1327 1123
rect 1331 1122 1332 1123
rect 1331 1120 1425 1122
rect 1331 1119 1332 1120
rect 1326 1118 1332 1119
rect 1703 1119 1709 1120
rect 1703 1118 1704 1119
rect 1645 1116 1704 1118
rect 1106 1114 1112 1115
rect 1703 1115 1704 1116
rect 1708 1115 1709 1119
rect 1838 1119 1844 1120
rect 1838 1118 1839 1119
rect 1829 1116 1839 1118
rect 1703 1114 1709 1115
rect 1838 1115 1839 1116
rect 1843 1115 1844 1119
rect 2046 1116 2052 1117
rect 3942 1116 3948 1117
rect 1838 1114 1844 1115
rect 2006 1115 2012 1116
rect 110 1110 116 1111
rect 174 1112 180 1113
rect 174 1108 175 1112
rect 179 1108 180 1112
rect 174 1107 180 1108
rect 326 1112 332 1113
rect 326 1108 327 1112
rect 331 1108 332 1112
rect 326 1107 332 1108
rect 494 1112 500 1113
rect 494 1108 495 1112
rect 499 1108 500 1112
rect 494 1107 500 1108
rect 670 1112 676 1113
rect 670 1108 671 1112
rect 675 1108 676 1112
rect 670 1107 676 1108
rect 846 1112 852 1113
rect 846 1108 847 1112
rect 851 1108 852 1112
rect 846 1107 852 1108
rect 1030 1112 1036 1113
rect 1030 1108 1031 1112
rect 1035 1108 1036 1112
rect 1030 1107 1036 1108
rect 1206 1112 1212 1113
rect 1206 1108 1207 1112
rect 1211 1108 1212 1112
rect 1206 1107 1212 1108
rect 1382 1112 1388 1113
rect 1382 1108 1383 1112
rect 1387 1108 1388 1112
rect 1382 1107 1388 1108
rect 1566 1112 1572 1113
rect 1566 1108 1567 1112
rect 1571 1108 1572 1112
rect 1566 1107 1572 1108
rect 1750 1112 1756 1113
rect 1750 1108 1751 1112
rect 1755 1108 1756 1112
rect 2006 1111 2007 1115
rect 2011 1111 2012 1115
rect 2046 1112 2047 1116
rect 2051 1112 2052 1116
rect 2046 1111 2052 1112
rect 2294 1115 2300 1116
rect 2294 1111 2295 1115
rect 2299 1111 2300 1115
rect 2006 1110 2012 1111
rect 2294 1110 2300 1111
rect 2422 1115 2428 1116
rect 2422 1111 2423 1115
rect 2427 1111 2428 1115
rect 2422 1110 2428 1111
rect 2558 1115 2564 1116
rect 2558 1111 2559 1115
rect 2563 1111 2564 1115
rect 2558 1110 2564 1111
rect 2694 1115 2700 1116
rect 2694 1111 2695 1115
rect 2699 1111 2700 1115
rect 2694 1110 2700 1111
rect 2838 1115 2844 1116
rect 2838 1111 2839 1115
rect 2843 1111 2844 1115
rect 2838 1110 2844 1111
rect 2990 1115 2996 1116
rect 2990 1111 2991 1115
rect 2995 1111 2996 1115
rect 2990 1110 2996 1111
rect 3150 1115 3156 1116
rect 3150 1111 3151 1115
rect 3155 1111 3156 1115
rect 3150 1110 3156 1111
rect 3318 1115 3324 1116
rect 3318 1111 3319 1115
rect 3323 1111 3324 1115
rect 3318 1110 3324 1111
rect 3494 1115 3500 1116
rect 3494 1111 3495 1115
rect 3499 1111 3500 1115
rect 3494 1110 3500 1111
rect 3678 1115 3684 1116
rect 3678 1111 3679 1115
rect 3683 1111 3684 1115
rect 3678 1110 3684 1111
rect 3838 1115 3844 1116
rect 3838 1111 3839 1115
rect 3843 1111 3844 1115
rect 3942 1112 3943 1116
rect 3947 1112 3948 1116
rect 3942 1111 3948 1112
rect 3838 1110 3844 1111
rect 1750 1107 1756 1108
rect 2914 1107 2920 1108
rect 2370 1103 2376 1104
rect 2046 1099 2052 1100
rect 2046 1095 2047 1099
rect 2051 1095 2052 1099
rect 2370 1099 2371 1103
rect 2375 1099 2376 1103
rect 2370 1098 2376 1099
rect 2498 1103 2504 1104
rect 2498 1099 2499 1103
rect 2503 1099 2504 1103
rect 2498 1098 2504 1099
rect 2634 1103 2640 1104
rect 2634 1099 2635 1103
rect 2639 1099 2640 1103
rect 2634 1098 2640 1099
rect 2770 1103 2776 1104
rect 2770 1099 2771 1103
rect 2775 1099 2776 1103
rect 2914 1103 2915 1107
rect 2919 1103 2920 1107
rect 3258 1107 3264 1108
rect 2914 1102 2920 1103
rect 3066 1103 3072 1104
rect 2770 1098 2776 1099
rect 3066 1099 3067 1103
rect 3071 1099 3072 1103
rect 3066 1098 3072 1099
rect 3226 1103 3232 1104
rect 3226 1099 3227 1103
rect 3231 1099 3232 1103
rect 3258 1103 3259 1107
rect 3263 1106 3264 1107
rect 3578 1107 3584 1108
rect 3263 1104 3361 1106
rect 3263 1103 3264 1104
rect 3258 1102 3264 1103
rect 3570 1103 3576 1104
rect 3226 1098 3232 1099
rect 3570 1099 3571 1103
rect 3575 1099 3576 1103
rect 3578 1103 3579 1107
rect 3583 1106 3584 1107
rect 3914 1107 3920 1108
rect 3583 1104 3721 1106
rect 3583 1103 3584 1104
rect 3578 1102 3584 1103
rect 3914 1103 3915 1107
rect 3919 1103 3920 1107
rect 3914 1102 3920 1103
rect 3570 1098 3576 1099
rect 3942 1099 3948 1100
rect 2046 1094 2052 1095
rect 2294 1096 2300 1097
rect 2294 1092 2295 1096
rect 2299 1092 2300 1096
rect 250 1091 256 1092
rect 227 1087 233 1088
rect 227 1083 228 1087
rect 232 1086 233 1087
rect 242 1087 248 1088
rect 242 1086 243 1087
rect 232 1084 243 1086
rect 232 1083 233 1084
rect 227 1082 233 1083
rect 242 1083 243 1084
rect 247 1083 248 1087
rect 250 1087 251 1091
rect 255 1090 256 1091
rect 379 1091 385 1092
rect 379 1090 380 1091
rect 255 1088 380 1090
rect 255 1087 256 1088
rect 250 1086 256 1087
rect 379 1087 380 1088
rect 384 1087 385 1091
rect 379 1086 385 1087
rect 402 1091 408 1092
rect 402 1087 403 1091
rect 407 1090 408 1091
rect 547 1091 553 1092
rect 547 1090 548 1091
rect 407 1088 548 1090
rect 407 1087 408 1088
rect 402 1086 408 1087
rect 547 1087 548 1088
rect 552 1087 553 1091
rect 547 1086 553 1087
rect 570 1091 576 1092
rect 570 1087 571 1091
rect 575 1090 576 1091
rect 723 1091 729 1092
rect 723 1090 724 1091
rect 575 1088 724 1090
rect 575 1087 576 1088
rect 570 1086 576 1087
rect 723 1087 724 1088
rect 728 1087 729 1091
rect 723 1086 729 1087
rect 746 1091 752 1092
rect 746 1087 747 1091
rect 751 1090 752 1091
rect 899 1091 905 1092
rect 899 1090 900 1091
rect 751 1088 900 1090
rect 751 1087 752 1088
rect 746 1086 752 1087
rect 899 1087 900 1088
rect 904 1087 905 1091
rect 899 1086 905 1087
rect 1083 1091 1092 1092
rect 1083 1087 1084 1091
rect 1091 1087 1092 1091
rect 1083 1086 1092 1087
rect 1259 1091 1265 1092
rect 1259 1087 1260 1091
rect 1264 1090 1265 1091
rect 1326 1091 1332 1092
rect 1326 1090 1327 1091
rect 1264 1088 1327 1090
rect 1264 1087 1265 1088
rect 1259 1086 1265 1087
rect 1326 1087 1327 1088
rect 1331 1087 1332 1091
rect 1619 1091 1625 1092
rect 1326 1086 1332 1087
rect 1435 1087 1441 1088
rect 242 1082 248 1083
rect 1435 1083 1436 1087
rect 1440 1086 1441 1087
rect 1455 1087 1461 1088
rect 1455 1086 1456 1087
rect 1440 1084 1456 1086
rect 1440 1083 1441 1084
rect 1435 1082 1441 1083
rect 1455 1083 1456 1084
rect 1460 1083 1461 1087
rect 1619 1087 1620 1091
rect 1624 1090 1625 1091
rect 1662 1091 1668 1092
rect 1662 1090 1663 1091
rect 1624 1088 1663 1090
rect 1624 1087 1625 1088
rect 1619 1086 1625 1087
rect 1662 1087 1663 1088
rect 1667 1087 1668 1091
rect 1662 1086 1668 1087
rect 1703 1091 1709 1092
rect 1703 1087 1704 1091
rect 1708 1090 1709 1091
rect 1803 1091 1809 1092
rect 2294 1091 2300 1092
rect 2422 1096 2428 1097
rect 2422 1092 2423 1096
rect 2427 1092 2428 1096
rect 2422 1091 2428 1092
rect 2558 1096 2564 1097
rect 2558 1092 2559 1096
rect 2563 1092 2564 1096
rect 2558 1091 2564 1092
rect 2694 1096 2700 1097
rect 2694 1092 2695 1096
rect 2699 1092 2700 1096
rect 2694 1091 2700 1092
rect 2838 1096 2844 1097
rect 2838 1092 2839 1096
rect 2843 1092 2844 1096
rect 2838 1091 2844 1092
rect 2990 1096 2996 1097
rect 2990 1092 2991 1096
rect 2995 1092 2996 1096
rect 2990 1091 2996 1092
rect 3150 1096 3156 1097
rect 3150 1092 3151 1096
rect 3155 1092 3156 1096
rect 3150 1091 3156 1092
rect 3318 1096 3324 1097
rect 3318 1092 3319 1096
rect 3323 1092 3324 1096
rect 3318 1091 3324 1092
rect 3494 1096 3500 1097
rect 3494 1092 3495 1096
rect 3499 1092 3500 1096
rect 3494 1091 3500 1092
rect 3678 1096 3684 1097
rect 3678 1092 3679 1096
rect 3683 1092 3684 1096
rect 3678 1091 3684 1092
rect 3838 1096 3844 1097
rect 3838 1092 3839 1096
rect 3843 1092 3844 1096
rect 3942 1095 3943 1099
rect 3947 1095 3948 1099
rect 3942 1094 3948 1095
rect 3838 1091 3844 1092
rect 1803 1090 1804 1091
rect 1708 1088 1804 1090
rect 1708 1087 1709 1088
rect 1703 1086 1709 1087
rect 1803 1087 1804 1088
rect 1808 1087 1809 1091
rect 1803 1086 1809 1087
rect 1455 1082 1461 1083
rect 3258 1083 3264 1084
rect 3258 1082 3259 1083
rect 3060 1080 3259 1082
rect 2370 1079 2376 1080
rect 2370 1075 2371 1079
rect 2375 1078 2376 1079
rect 2375 1076 2434 1078
rect 2375 1075 2376 1076
rect 2370 1074 2376 1075
rect 2432 1074 2434 1076
rect 2475 1075 2481 1076
rect 2475 1074 2476 1075
rect 2432 1072 2476 1074
rect 2347 1071 2353 1072
rect 187 1067 193 1068
rect 187 1063 188 1067
rect 192 1066 193 1067
rect 202 1067 208 1068
rect 202 1066 203 1067
rect 192 1064 203 1066
rect 192 1063 193 1064
rect 187 1062 193 1063
rect 202 1063 203 1064
rect 207 1063 208 1067
rect 202 1062 208 1063
rect 210 1067 216 1068
rect 210 1063 211 1067
rect 215 1066 216 1067
rect 283 1067 289 1068
rect 283 1066 284 1067
rect 215 1064 284 1066
rect 215 1063 216 1064
rect 210 1062 216 1063
rect 283 1063 284 1064
rect 288 1063 289 1067
rect 283 1062 289 1063
rect 306 1067 312 1068
rect 306 1063 307 1067
rect 311 1066 312 1067
rect 427 1067 433 1068
rect 427 1066 428 1067
rect 311 1064 428 1066
rect 311 1063 312 1064
rect 306 1062 312 1063
rect 427 1063 428 1064
rect 432 1063 433 1067
rect 427 1062 433 1063
rect 450 1067 456 1068
rect 450 1063 451 1067
rect 455 1066 456 1067
rect 595 1067 601 1068
rect 595 1066 596 1067
rect 455 1064 596 1066
rect 455 1063 456 1064
rect 450 1062 456 1063
rect 595 1063 596 1064
rect 600 1063 601 1067
rect 595 1062 601 1063
rect 618 1067 624 1068
rect 618 1063 619 1067
rect 623 1066 624 1067
rect 779 1067 785 1068
rect 779 1066 780 1067
rect 623 1064 780 1066
rect 623 1063 624 1064
rect 618 1062 624 1063
rect 779 1063 780 1064
rect 784 1063 785 1067
rect 779 1062 785 1063
rect 802 1067 808 1068
rect 802 1063 803 1067
rect 807 1066 808 1067
rect 963 1067 969 1068
rect 963 1066 964 1067
rect 807 1064 964 1066
rect 807 1063 808 1064
rect 802 1062 808 1063
rect 963 1063 964 1064
rect 968 1063 969 1067
rect 963 1062 969 1063
rect 1106 1067 1112 1068
rect 1106 1063 1107 1067
rect 1111 1066 1112 1067
rect 1147 1067 1153 1068
rect 1147 1066 1148 1067
rect 1111 1064 1148 1066
rect 1111 1063 1112 1064
rect 1106 1062 1112 1063
rect 1147 1063 1148 1064
rect 1152 1063 1153 1067
rect 1147 1062 1153 1063
rect 1326 1067 1337 1068
rect 1326 1063 1327 1067
rect 1331 1063 1332 1067
rect 1336 1063 1337 1067
rect 1326 1062 1337 1063
rect 1354 1067 1360 1068
rect 1354 1063 1355 1067
rect 1359 1066 1360 1067
rect 1515 1067 1521 1068
rect 1515 1066 1516 1067
rect 1359 1064 1516 1066
rect 1359 1063 1360 1064
rect 1354 1062 1360 1063
rect 1515 1063 1516 1064
rect 1520 1063 1521 1067
rect 1515 1062 1521 1063
rect 1699 1067 1705 1068
rect 1699 1063 1700 1067
rect 1704 1066 1705 1067
rect 1734 1067 1740 1068
rect 1734 1066 1735 1067
rect 1704 1064 1735 1066
rect 1704 1063 1705 1064
rect 1699 1062 1705 1063
rect 1734 1063 1735 1064
rect 1739 1063 1740 1067
rect 1734 1062 1740 1063
rect 1838 1067 1844 1068
rect 1838 1063 1839 1067
rect 1843 1066 1844 1067
rect 1883 1067 1889 1068
rect 1883 1066 1884 1067
rect 1843 1064 1884 1066
rect 1843 1063 1844 1064
rect 1838 1062 1844 1063
rect 1883 1063 1884 1064
rect 1888 1063 1889 1067
rect 2347 1067 2348 1071
rect 2352 1070 2353 1071
rect 2423 1071 2429 1072
rect 2423 1070 2424 1071
rect 2352 1068 2424 1070
rect 2352 1067 2353 1068
rect 2347 1066 2353 1067
rect 2423 1067 2424 1068
rect 2428 1067 2429 1071
rect 2475 1071 2476 1072
rect 2480 1071 2481 1075
rect 2475 1070 2481 1071
rect 2498 1075 2504 1076
rect 2498 1071 2499 1075
rect 2503 1074 2504 1075
rect 2611 1075 2617 1076
rect 2611 1074 2612 1075
rect 2503 1072 2612 1074
rect 2503 1071 2504 1072
rect 2498 1070 2504 1071
rect 2611 1071 2612 1072
rect 2616 1071 2617 1075
rect 2611 1070 2617 1071
rect 2634 1075 2640 1076
rect 2634 1071 2635 1075
rect 2639 1074 2640 1075
rect 2747 1075 2753 1076
rect 2747 1074 2748 1075
rect 2639 1072 2748 1074
rect 2639 1071 2640 1072
rect 2634 1070 2640 1071
rect 2747 1071 2748 1072
rect 2752 1071 2753 1075
rect 2747 1070 2753 1071
rect 2770 1075 2776 1076
rect 2770 1071 2771 1075
rect 2775 1074 2776 1075
rect 2891 1075 2897 1076
rect 2891 1074 2892 1075
rect 2775 1072 2892 1074
rect 2775 1071 2776 1072
rect 2770 1070 2776 1071
rect 2891 1071 2892 1072
rect 2896 1071 2897 1075
rect 2891 1070 2897 1071
rect 3043 1075 3049 1076
rect 3043 1071 3044 1075
rect 3048 1074 3049 1075
rect 3060 1074 3062 1080
rect 3258 1079 3259 1080
rect 3263 1079 3264 1083
rect 3578 1083 3584 1084
rect 3578 1082 3579 1083
rect 3258 1078 3264 1079
rect 3468 1080 3579 1082
rect 3048 1072 3062 1074
rect 3066 1075 3072 1076
rect 3048 1071 3049 1072
rect 3043 1070 3049 1071
rect 3066 1071 3067 1075
rect 3071 1074 3072 1075
rect 3203 1075 3209 1076
rect 3203 1074 3204 1075
rect 3071 1072 3204 1074
rect 3071 1071 3072 1072
rect 3066 1070 3072 1071
rect 3203 1071 3204 1072
rect 3208 1071 3209 1075
rect 3203 1070 3209 1071
rect 3371 1075 3377 1076
rect 3371 1071 3372 1075
rect 3376 1074 3377 1075
rect 3468 1074 3470 1080
rect 3578 1079 3579 1080
rect 3583 1079 3584 1083
rect 3578 1078 3584 1079
rect 3376 1072 3470 1074
rect 3474 1075 3480 1076
rect 3376 1071 3377 1072
rect 3371 1070 3377 1071
rect 3474 1071 3475 1075
rect 3479 1074 3480 1075
rect 3547 1075 3553 1076
rect 3547 1074 3548 1075
rect 3479 1072 3548 1074
rect 3479 1071 3480 1072
rect 3474 1070 3480 1071
rect 3547 1071 3548 1072
rect 3552 1071 3553 1075
rect 3547 1070 3553 1071
rect 3570 1075 3576 1076
rect 3570 1071 3571 1075
rect 3575 1074 3576 1075
rect 3731 1075 3737 1076
rect 3731 1074 3732 1075
rect 3575 1072 3732 1074
rect 3575 1071 3576 1072
rect 3570 1070 3576 1071
rect 3731 1071 3732 1072
rect 3736 1071 3737 1075
rect 3731 1070 3737 1071
rect 3891 1071 3897 1072
rect 2423 1066 2429 1067
rect 3891 1067 3892 1071
rect 3896 1070 3897 1071
rect 3906 1071 3912 1072
rect 3906 1070 3907 1071
rect 3896 1068 3907 1070
rect 3896 1067 3897 1068
rect 3891 1066 3897 1067
rect 3906 1067 3907 1068
rect 3911 1067 3912 1071
rect 3906 1066 3912 1067
rect 1883 1062 1889 1063
rect 2547 1055 2553 1056
rect 2547 1051 2548 1055
rect 2552 1054 2553 1055
rect 2578 1055 2584 1056
rect 2578 1054 2579 1055
rect 2552 1052 2579 1054
rect 2552 1051 2553 1052
rect 2547 1050 2553 1051
rect 2578 1051 2579 1052
rect 2583 1051 2584 1055
rect 2578 1050 2584 1051
rect 2651 1055 2657 1056
rect 2651 1051 2652 1055
rect 2656 1054 2657 1055
rect 2682 1055 2688 1056
rect 2682 1054 2683 1055
rect 2656 1052 2683 1054
rect 2656 1051 2657 1052
rect 2651 1050 2657 1051
rect 2682 1051 2683 1052
rect 2687 1051 2688 1055
rect 2682 1050 2688 1051
rect 2763 1055 2769 1056
rect 2763 1051 2764 1055
rect 2768 1054 2769 1055
rect 2799 1055 2805 1056
rect 2799 1054 2800 1055
rect 2768 1052 2800 1054
rect 2768 1051 2769 1052
rect 2763 1050 2769 1051
rect 2799 1051 2800 1052
rect 2804 1051 2805 1055
rect 2799 1050 2805 1051
rect 2899 1055 2905 1056
rect 2899 1051 2900 1055
rect 2904 1054 2905 1055
rect 2922 1055 2928 1056
rect 2922 1054 2923 1055
rect 2904 1052 2923 1054
rect 2904 1051 2905 1052
rect 2899 1050 2905 1051
rect 2922 1051 2923 1052
rect 2927 1051 2928 1055
rect 2922 1050 2928 1051
rect 3059 1055 3065 1056
rect 3059 1051 3060 1055
rect 3064 1054 3065 1055
rect 3190 1055 3196 1056
rect 3190 1054 3191 1055
rect 3064 1052 3191 1054
rect 3064 1051 3065 1052
rect 3059 1050 3065 1051
rect 3190 1051 3191 1052
rect 3195 1051 3196 1055
rect 3190 1050 3196 1051
rect 3226 1055 3232 1056
rect 3226 1051 3227 1055
rect 3231 1054 3232 1055
rect 3251 1055 3257 1056
rect 3251 1054 3252 1055
rect 3231 1052 3252 1054
rect 3231 1051 3232 1052
rect 3226 1050 3232 1051
rect 3251 1051 3252 1052
rect 3256 1051 3257 1055
rect 3251 1050 3257 1051
rect 3274 1055 3280 1056
rect 3274 1051 3275 1055
rect 3279 1054 3280 1055
rect 3459 1055 3465 1056
rect 3459 1054 3460 1055
rect 3279 1052 3460 1054
rect 3279 1051 3280 1052
rect 3274 1050 3280 1051
rect 3459 1051 3460 1052
rect 3464 1051 3465 1055
rect 3459 1050 3465 1051
rect 3482 1055 3488 1056
rect 3482 1051 3483 1055
rect 3487 1054 3488 1055
rect 3683 1055 3689 1056
rect 3683 1054 3684 1055
rect 3487 1052 3684 1054
rect 3487 1051 3488 1052
rect 3482 1050 3488 1051
rect 3683 1051 3684 1052
rect 3688 1051 3689 1055
rect 3683 1050 3689 1051
rect 3891 1055 3897 1056
rect 3891 1051 3892 1055
rect 3896 1054 3897 1055
rect 3914 1055 3920 1056
rect 3914 1054 3915 1055
rect 3896 1052 3915 1054
rect 3896 1051 3897 1052
rect 3891 1050 3897 1051
rect 3914 1051 3915 1052
rect 3919 1051 3920 1055
rect 3914 1050 3920 1051
rect 134 1044 140 1045
rect 110 1041 116 1042
rect 110 1037 111 1041
rect 115 1037 116 1041
rect 134 1040 135 1044
rect 139 1040 140 1044
rect 134 1039 140 1040
rect 230 1044 236 1045
rect 230 1040 231 1044
rect 235 1040 236 1044
rect 230 1039 236 1040
rect 374 1044 380 1045
rect 374 1040 375 1044
rect 379 1040 380 1044
rect 374 1039 380 1040
rect 542 1044 548 1045
rect 542 1040 543 1044
rect 547 1040 548 1044
rect 542 1039 548 1040
rect 726 1044 732 1045
rect 726 1040 727 1044
rect 731 1040 732 1044
rect 726 1039 732 1040
rect 910 1044 916 1045
rect 910 1040 911 1044
rect 915 1040 916 1044
rect 910 1039 916 1040
rect 1094 1044 1100 1045
rect 1094 1040 1095 1044
rect 1099 1040 1100 1044
rect 1094 1039 1100 1040
rect 1278 1044 1284 1045
rect 1278 1040 1279 1044
rect 1283 1040 1284 1044
rect 1278 1039 1284 1040
rect 1462 1044 1468 1045
rect 1462 1040 1463 1044
rect 1467 1040 1468 1044
rect 1462 1039 1468 1040
rect 1646 1044 1652 1045
rect 1646 1040 1647 1044
rect 1651 1040 1652 1044
rect 1646 1039 1652 1040
rect 1830 1044 1836 1045
rect 1830 1040 1831 1044
rect 1835 1040 1836 1044
rect 1830 1039 1836 1040
rect 2006 1041 2012 1042
rect 110 1036 116 1037
rect 2006 1037 2007 1041
rect 2011 1037 2012 1041
rect 2006 1036 2012 1037
rect 210 1035 216 1036
rect 210 1031 211 1035
rect 215 1031 216 1035
rect 210 1030 216 1031
rect 306 1035 312 1036
rect 306 1031 307 1035
rect 311 1031 312 1035
rect 306 1030 312 1031
rect 450 1035 456 1036
rect 450 1031 451 1035
rect 455 1031 456 1035
rect 450 1030 456 1031
rect 618 1035 624 1036
rect 618 1031 619 1035
rect 623 1031 624 1035
rect 618 1030 624 1031
rect 802 1035 808 1036
rect 802 1031 803 1035
rect 807 1031 808 1035
rect 802 1030 808 1031
rect 858 1035 864 1036
rect 858 1031 859 1035
rect 863 1034 864 1035
rect 1062 1035 1068 1036
rect 863 1032 953 1034
rect 863 1031 864 1032
rect 858 1030 864 1031
rect 1062 1031 1063 1035
rect 1067 1034 1068 1035
rect 1354 1035 1360 1036
rect 1067 1032 1137 1034
rect 1067 1031 1068 1032
rect 1062 1030 1068 1031
rect 1354 1031 1355 1035
rect 1359 1031 1360 1035
rect 1354 1030 1360 1031
rect 1455 1035 1461 1036
rect 1455 1031 1456 1035
rect 1460 1034 1461 1035
rect 1554 1035 1560 1036
rect 1460 1032 1505 1034
rect 1460 1031 1461 1032
rect 1455 1030 1461 1031
rect 1554 1031 1555 1035
rect 1559 1034 1560 1035
rect 1734 1035 1740 1036
rect 1559 1032 1689 1034
rect 1559 1031 1560 1032
rect 1554 1030 1560 1031
rect 1734 1031 1735 1035
rect 1739 1034 1740 1035
rect 1739 1032 1873 1034
rect 2494 1032 2500 1033
rect 1739 1031 1740 1032
rect 1734 1030 1740 1031
rect 2046 1029 2052 1030
rect 134 1025 140 1026
rect 110 1024 116 1025
rect 110 1020 111 1024
rect 115 1020 116 1024
rect 134 1021 135 1025
rect 139 1021 140 1025
rect 134 1020 140 1021
rect 230 1025 236 1026
rect 230 1021 231 1025
rect 235 1021 236 1025
rect 230 1020 236 1021
rect 374 1025 380 1026
rect 374 1021 375 1025
rect 379 1021 380 1025
rect 374 1020 380 1021
rect 542 1025 548 1026
rect 542 1021 543 1025
rect 547 1021 548 1025
rect 542 1020 548 1021
rect 726 1025 732 1026
rect 726 1021 727 1025
rect 731 1021 732 1025
rect 726 1020 732 1021
rect 910 1025 916 1026
rect 910 1021 911 1025
rect 915 1021 916 1025
rect 910 1020 916 1021
rect 1094 1025 1100 1026
rect 1094 1021 1095 1025
rect 1099 1021 1100 1025
rect 1094 1020 1100 1021
rect 1278 1025 1284 1026
rect 1278 1021 1279 1025
rect 1283 1021 1284 1025
rect 1278 1020 1284 1021
rect 1462 1025 1468 1026
rect 1462 1021 1463 1025
rect 1467 1021 1468 1025
rect 1462 1020 1468 1021
rect 1646 1025 1652 1026
rect 1646 1021 1647 1025
rect 1651 1021 1652 1025
rect 1646 1020 1652 1021
rect 1830 1025 1836 1026
rect 2046 1025 2047 1029
rect 2051 1025 2052 1029
rect 2494 1028 2495 1032
rect 2499 1028 2500 1032
rect 2494 1027 2500 1028
rect 2598 1032 2604 1033
rect 2598 1028 2599 1032
rect 2603 1028 2604 1032
rect 2598 1027 2604 1028
rect 2710 1032 2716 1033
rect 2710 1028 2711 1032
rect 2715 1028 2716 1032
rect 2710 1027 2716 1028
rect 2846 1032 2852 1033
rect 2846 1028 2847 1032
rect 2851 1028 2852 1032
rect 2846 1027 2852 1028
rect 3006 1032 3012 1033
rect 3006 1028 3007 1032
rect 3011 1028 3012 1032
rect 3006 1027 3012 1028
rect 3198 1032 3204 1033
rect 3198 1028 3199 1032
rect 3203 1028 3204 1032
rect 3198 1027 3204 1028
rect 3406 1032 3412 1033
rect 3406 1028 3407 1032
rect 3411 1028 3412 1032
rect 3406 1027 3412 1028
rect 3630 1032 3636 1033
rect 3630 1028 3631 1032
rect 3635 1028 3636 1032
rect 3630 1027 3636 1028
rect 3838 1032 3844 1033
rect 3838 1028 3839 1032
rect 3843 1028 3844 1032
rect 3838 1027 3844 1028
rect 3942 1029 3948 1030
rect 1830 1021 1831 1025
rect 1835 1021 1836 1025
rect 1830 1020 1836 1021
rect 2006 1024 2012 1025
rect 2046 1024 2052 1025
rect 3942 1025 3943 1029
rect 3947 1025 3948 1029
rect 3942 1024 3948 1025
rect 2006 1020 2007 1024
rect 2011 1020 2012 1024
rect 110 1019 116 1020
rect 2006 1019 2012 1020
rect 2423 1023 2429 1024
rect 2423 1019 2424 1023
rect 2428 1022 2429 1023
rect 2578 1023 2584 1024
rect 2428 1020 2537 1022
rect 2428 1019 2429 1020
rect 2423 1018 2429 1019
rect 2578 1019 2579 1023
rect 2583 1022 2584 1023
rect 2682 1023 2688 1024
rect 2583 1020 2641 1022
rect 2583 1019 2584 1020
rect 2578 1018 2584 1019
rect 2682 1019 2683 1023
rect 2687 1022 2688 1023
rect 2799 1023 2805 1024
rect 2687 1020 2753 1022
rect 2687 1019 2688 1020
rect 2682 1018 2688 1019
rect 2799 1019 2800 1023
rect 2804 1022 2805 1023
rect 3074 1023 3080 1024
rect 2804 1020 2889 1022
rect 2804 1019 2805 1020
rect 2799 1018 2805 1019
rect 3074 1019 3075 1023
rect 3079 1019 3080 1023
rect 3074 1018 3080 1019
rect 3274 1023 3280 1024
rect 3274 1019 3275 1023
rect 3279 1019 3280 1023
rect 3274 1018 3280 1019
rect 3482 1023 3488 1024
rect 3482 1019 3483 1023
rect 3487 1019 3488 1023
rect 3482 1018 3488 1019
rect 3558 1023 3564 1024
rect 3558 1019 3559 1023
rect 3563 1022 3564 1023
rect 3906 1023 3912 1024
rect 3563 1020 3673 1022
rect 3563 1019 3564 1020
rect 3558 1018 3564 1019
rect 3906 1019 3907 1023
rect 3911 1019 3912 1023
rect 3906 1018 3912 1019
rect 2494 1013 2500 1014
rect 2046 1012 2052 1013
rect 2046 1008 2047 1012
rect 2051 1008 2052 1012
rect 2494 1009 2495 1013
rect 2499 1009 2500 1013
rect 2494 1008 2500 1009
rect 2598 1013 2604 1014
rect 2598 1009 2599 1013
rect 2603 1009 2604 1013
rect 2598 1008 2604 1009
rect 2710 1013 2716 1014
rect 2710 1009 2711 1013
rect 2715 1009 2716 1013
rect 2710 1008 2716 1009
rect 2846 1013 2852 1014
rect 2846 1009 2847 1013
rect 2851 1009 2852 1013
rect 2846 1008 2852 1009
rect 3006 1013 3012 1014
rect 3006 1009 3007 1013
rect 3011 1009 3012 1013
rect 3006 1008 3012 1009
rect 3198 1013 3204 1014
rect 3198 1009 3199 1013
rect 3203 1009 3204 1013
rect 3198 1008 3204 1009
rect 3406 1013 3412 1014
rect 3406 1009 3407 1013
rect 3411 1009 3412 1013
rect 3406 1008 3412 1009
rect 3630 1013 3636 1014
rect 3630 1009 3631 1013
rect 3635 1009 3636 1013
rect 3630 1008 3636 1009
rect 3838 1013 3844 1014
rect 3838 1009 3839 1013
rect 3843 1009 3844 1013
rect 3838 1008 3844 1009
rect 3942 1012 3948 1013
rect 3942 1008 3943 1012
rect 3947 1008 3948 1012
rect 2046 1007 2052 1008
rect 3942 1007 3948 1008
rect 110 972 116 973
rect 2006 972 2012 973
rect 110 968 111 972
rect 115 968 116 972
rect 110 967 116 968
rect 134 971 140 972
rect 134 967 135 971
rect 139 967 140 971
rect 270 971 276 972
rect 134 966 140 967
rect 202 967 208 968
rect 202 963 203 967
rect 207 966 208 967
rect 270 967 271 971
rect 275 967 276 971
rect 270 966 276 967
rect 446 971 452 972
rect 446 967 447 971
rect 451 967 452 971
rect 446 966 452 967
rect 630 971 636 972
rect 630 967 631 971
rect 635 967 636 971
rect 630 966 636 967
rect 822 971 828 972
rect 822 967 823 971
rect 827 967 828 971
rect 822 966 828 967
rect 1006 971 1012 972
rect 1006 967 1007 971
rect 1011 967 1012 971
rect 1006 966 1012 967
rect 1174 971 1180 972
rect 1174 967 1175 971
rect 1179 967 1180 971
rect 1174 966 1180 967
rect 1334 971 1340 972
rect 1334 967 1335 971
rect 1339 967 1340 971
rect 1334 966 1340 967
rect 1486 971 1492 972
rect 1486 967 1487 971
rect 1491 967 1492 971
rect 1486 966 1492 967
rect 1630 971 1636 972
rect 1630 967 1631 971
rect 1635 967 1636 971
rect 1630 966 1636 967
rect 1774 971 1780 972
rect 1774 967 1775 971
rect 1779 967 1780 971
rect 1774 966 1780 967
rect 1902 971 1908 972
rect 1902 967 1903 971
rect 1907 967 1908 971
rect 2006 968 2007 972
rect 2011 968 2012 972
rect 2006 967 2012 968
rect 1902 966 1908 967
rect 207 964 214 966
rect 207 963 208 964
rect 202 962 208 963
rect 212 961 214 964
rect 250 963 256 964
rect 250 959 251 963
rect 255 962 256 963
rect 407 963 413 964
rect 255 960 313 962
rect 255 959 256 960
rect 250 958 256 959
rect 407 959 408 963
rect 412 962 413 963
rect 586 963 592 964
rect 412 960 489 962
rect 412 959 413 960
rect 407 958 413 959
rect 586 959 587 963
rect 591 962 592 963
rect 714 963 720 964
rect 591 960 673 962
rect 591 959 592 960
rect 586 958 592 959
rect 714 959 715 963
rect 719 962 720 963
rect 1326 963 1332 964
rect 719 960 865 962
rect 719 959 720 960
rect 714 958 720 959
rect 1082 959 1088 960
rect 110 955 116 956
rect 110 951 111 955
rect 115 951 116 955
rect 1082 955 1083 959
rect 1087 955 1088 959
rect 1082 954 1088 955
rect 1250 959 1256 960
rect 1250 955 1251 959
rect 1255 955 1256 959
rect 1326 959 1327 963
rect 1331 962 1332 963
rect 1870 963 1876 964
rect 1331 960 1377 962
rect 1331 959 1332 960
rect 1326 958 1332 959
rect 1562 959 1568 960
rect 1250 954 1256 955
rect 1562 955 1563 959
rect 1567 955 1568 959
rect 1562 954 1568 955
rect 1706 959 1712 960
rect 1706 955 1707 959
rect 1711 955 1712 959
rect 1706 954 1712 955
rect 1850 959 1856 960
rect 1850 955 1851 959
rect 1855 955 1856 959
rect 1870 959 1871 963
rect 1875 962 1876 963
rect 1875 960 1945 962
rect 2046 960 2052 961
rect 3942 960 3948 961
rect 1875 959 1876 960
rect 1870 958 1876 959
rect 2046 956 2047 960
rect 2051 956 2052 960
rect 1850 954 1856 955
rect 2006 955 2012 956
rect 2046 955 2052 956
rect 2646 959 2652 960
rect 2646 955 2647 959
rect 2651 955 2652 959
rect 110 950 116 951
rect 134 952 140 953
rect 134 948 135 952
rect 139 948 140 952
rect 134 947 140 948
rect 270 952 276 953
rect 270 948 271 952
rect 275 948 276 952
rect 270 947 276 948
rect 446 952 452 953
rect 446 948 447 952
rect 451 948 452 952
rect 446 947 452 948
rect 630 952 636 953
rect 630 948 631 952
rect 635 948 636 952
rect 630 947 636 948
rect 822 952 828 953
rect 822 948 823 952
rect 827 948 828 952
rect 822 947 828 948
rect 1006 952 1012 953
rect 1006 948 1007 952
rect 1011 948 1012 952
rect 1006 947 1012 948
rect 1174 952 1180 953
rect 1174 948 1175 952
rect 1179 948 1180 952
rect 1174 947 1180 948
rect 1334 952 1340 953
rect 1334 948 1335 952
rect 1339 948 1340 952
rect 1334 947 1340 948
rect 1486 952 1492 953
rect 1486 948 1487 952
rect 1491 948 1492 952
rect 1486 947 1492 948
rect 1630 952 1636 953
rect 1630 948 1631 952
rect 1635 948 1636 952
rect 1630 947 1636 948
rect 1774 952 1780 953
rect 1774 948 1775 952
rect 1779 948 1780 952
rect 1774 947 1780 948
rect 1902 952 1908 953
rect 1902 948 1903 952
rect 1907 948 1908 952
rect 2006 951 2007 955
rect 2011 951 2012 955
rect 2646 954 2652 955
rect 2742 959 2748 960
rect 2742 955 2743 959
rect 2747 955 2748 959
rect 2742 954 2748 955
rect 2846 959 2852 960
rect 2846 955 2847 959
rect 2851 955 2852 959
rect 2846 954 2852 955
rect 2966 959 2972 960
rect 2966 955 2967 959
rect 2971 955 2972 959
rect 2966 954 2972 955
rect 3110 959 3116 960
rect 3110 955 3111 959
rect 3115 955 3116 959
rect 3110 954 3116 955
rect 3278 959 3284 960
rect 3278 955 3279 959
rect 3283 955 3284 959
rect 3278 954 3284 955
rect 3462 959 3468 960
rect 3462 955 3463 959
rect 3467 955 3468 959
rect 3462 954 3468 955
rect 3662 959 3668 960
rect 3662 955 3663 959
rect 3667 955 3668 959
rect 3662 954 3668 955
rect 3838 959 3844 960
rect 3838 955 3839 959
rect 3843 955 3844 959
rect 3942 956 3943 960
rect 3947 956 3948 960
rect 3942 955 3948 956
rect 3838 954 3844 955
rect 2006 950 2012 951
rect 2922 951 2928 952
rect 1902 947 1908 948
rect 2722 947 2728 948
rect 2046 943 2052 944
rect 2046 939 2047 943
rect 2051 939 2052 943
rect 2722 943 2723 947
rect 2727 943 2728 947
rect 2722 942 2728 943
rect 2818 947 2824 948
rect 2818 943 2819 947
rect 2823 943 2824 947
rect 2922 947 2923 951
rect 2927 947 2928 951
rect 3622 951 3628 952
rect 2922 946 2928 947
rect 3086 947 3092 948
rect 3086 946 3087 947
rect 3045 944 3087 946
rect 2818 942 2824 943
rect 3086 943 3087 944
rect 3091 943 3092 947
rect 3086 942 3092 943
rect 3186 947 3192 948
rect 3186 943 3187 947
rect 3191 943 3192 947
rect 3186 942 3192 943
rect 3354 947 3360 948
rect 3354 943 3355 947
rect 3359 943 3360 947
rect 3354 942 3360 943
rect 3538 947 3544 948
rect 3538 943 3539 947
rect 3543 943 3544 947
rect 3622 947 3623 951
rect 3627 950 3628 951
rect 3914 951 3920 952
rect 3627 948 3705 950
rect 3627 947 3628 948
rect 3622 946 3628 947
rect 3914 947 3915 951
rect 3919 947 3920 951
rect 3914 946 3920 947
rect 3538 942 3544 943
rect 3942 943 3948 944
rect 2046 938 2052 939
rect 2646 940 2652 941
rect 2646 936 2647 940
rect 2651 936 2652 940
rect 2646 935 2652 936
rect 2742 940 2748 941
rect 2742 936 2743 940
rect 2747 936 2748 940
rect 2742 935 2748 936
rect 2846 940 2852 941
rect 2846 936 2847 940
rect 2851 936 2852 940
rect 2846 935 2852 936
rect 2966 940 2972 941
rect 2966 936 2967 940
rect 2971 936 2972 940
rect 2966 935 2972 936
rect 3110 940 3116 941
rect 3110 936 3111 940
rect 3115 936 3116 940
rect 3110 935 3116 936
rect 3278 940 3284 941
rect 3278 936 3279 940
rect 3283 936 3284 940
rect 3278 935 3284 936
rect 3462 940 3468 941
rect 3462 936 3463 940
rect 3467 936 3468 940
rect 3462 935 3468 936
rect 3662 940 3668 941
rect 3662 936 3663 940
rect 3667 936 3668 940
rect 3662 935 3668 936
rect 3838 940 3844 941
rect 3838 936 3839 940
rect 3843 936 3844 940
rect 3942 939 3943 943
rect 3947 939 3948 943
rect 3942 938 3948 939
rect 3838 935 3844 936
rect 187 931 193 932
rect 187 927 188 931
rect 192 930 193 931
rect 250 931 256 932
rect 250 930 251 931
rect 192 928 251 930
rect 192 927 193 928
rect 187 926 193 927
rect 250 927 251 928
rect 255 927 256 931
rect 250 926 256 927
rect 323 931 329 932
rect 323 927 324 931
rect 328 930 329 931
rect 407 931 413 932
rect 407 930 408 931
rect 328 928 408 930
rect 328 927 329 928
rect 323 926 329 927
rect 407 927 408 928
rect 412 927 413 931
rect 407 926 413 927
rect 499 931 505 932
rect 499 927 500 931
rect 504 930 505 931
rect 586 931 592 932
rect 586 930 587 931
rect 504 928 587 930
rect 504 927 505 928
rect 499 926 505 927
rect 586 927 587 928
rect 591 927 592 931
rect 586 926 592 927
rect 683 931 689 932
rect 683 927 684 931
rect 688 930 689 931
rect 714 931 720 932
rect 714 930 715 931
rect 688 928 715 930
rect 688 927 689 928
rect 683 926 689 927
rect 714 927 715 928
rect 719 927 720 931
rect 1059 931 1068 932
rect 714 926 720 927
rect 875 927 881 928
rect 875 923 876 927
rect 880 926 881 927
rect 922 927 928 928
rect 922 926 923 927
rect 880 924 923 926
rect 880 923 881 924
rect 875 922 881 923
rect 922 923 923 924
rect 927 923 928 927
rect 1059 927 1060 931
rect 1067 927 1068 931
rect 1250 931 1256 932
rect 1059 926 1068 927
rect 1227 927 1236 928
rect 922 922 928 923
rect 1227 923 1228 927
rect 1235 923 1236 927
rect 1250 927 1251 931
rect 1255 930 1256 931
rect 1387 931 1393 932
rect 1387 930 1388 931
rect 1255 928 1388 930
rect 1255 927 1256 928
rect 1250 926 1256 927
rect 1387 927 1388 928
rect 1392 927 1393 931
rect 1387 926 1393 927
rect 1539 931 1545 932
rect 1539 927 1540 931
rect 1544 930 1545 931
rect 1554 931 1560 932
rect 1554 930 1555 931
rect 1544 928 1555 930
rect 1544 927 1545 928
rect 1539 926 1545 927
rect 1554 927 1555 928
rect 1559 927 1560 931
rect 1554 926 1560 927
rect 1562 931 1568 932
rect 1562 927 1563 931
rect 1567 930 1568 931
rect 1683 931 1689 932
rect 1683 930 1684 931
rect 1567 928 1684 930
rect 1567 927 1568 928
rect 1562 926 1568 927
rect 1683 927 1684 928
rect 1688 927 1689 931
rect 1683 926 1689 927
rect 1706 931 1712 932
rect 1706 927 1707 931
rect 1711 930 1712 931
rect 1827 931 1833 932
rect 1827 930 1828 931
rect 1711 928 1828 930
rect 1711 927 1712 928
rect 1706 926 1712 927
rect 1827 927 1828 928
rect 1832 927 1833 931
rect 1827 926 1833 927
rect 1850 931 1856 932
rect 1850 927 1851 931
rect 1855 930 1856 931
rect 1955 931 1961 932
rect 1955 930 1956 931
rect 1855 928 1956 930
rect 1855 927 1856 928
rect 1850 926 1856 927
rect 1955 927 1956 928
rect 1960 927 1961 931
rect 1955 926 1961 927
rect 1227 922 1236 923
rect 1870 923 1876 924
rect 1870 922 1871 923
rect 1804 920 1871 922
rect 1804 918 1806 920
rect 1870 919 1871 920
rect 1875 919 1876 923
rect 1870 918 1876 919
rect 2722 923 2728 924
rect 2722 919 2723 923
rect 2727 922 2728 923
rect 2727 920 2762 922
rect 2727 919 2728 920
rect 2722 918 2728 919
rect 2760 918 2762 920
rect 2795 919 2801 920
rect 2795 918 2796 919
rect 1803 917 1809 918
rect 187 915 196 916
rect 187 911 188 915
rect 195 911 196 915
rect 187 910 196 911
rect 210 915 216 916
rect 210 911 211 915
rect 215 914 216 915
rect 323 915 329 916
rect 323 914 324 915
rect 215 912 324 914
rect 215 911 216 912
rect 210 910 216 911
rect 323 911 324 912
rect 328 911 329 915
rect 323 910 329 911
rect 346 915 352 916
rect 346 911 347 915
rect 351 914 352 915
rect 507 915 513 916
rect 507 914 508 915
rect 351 912 508 914
rect 351 911 352 912
rect 346 910 352 911
rect 507 911 508 912
rect 512 911 513 915
rect 507 910 513 911
rect 530 915 536 916
rect 530 911 531 915
rect 535 914 536 915
rect 707 915 713 916
rect 707 914 708 915
rect 535 912 708 914
rect 535 911 536 912
rect 530 910 536 911
rect 707 911 708 912
rect 712 911 713 915
rect 707 910 713 911
rect 730 915 736 916
rect 730 911 731 915
rect 735 914 736 915
rect 907 915 913 916
rect 907 914 908 915
rect 735 912 908 914
rect 735 911 736 912
rect 730 910 736 911
rect 907 911 908 912
rect 912 911 913 915
rect 907 910 913 911
rect 1082 915 1088 916
rect 1082 911 1083 915
rect 1087 914 1088 915
rect 1107 915 1113 916
rect 1107 914 1108 915
rect 1087 912 1108 914
rect 1087 911 1088 912
rect 1082 910 1088 911
rect 1107 911 1108 912
rect 1112 911 1113 915
rect 1107 910 1113 911
rect 1291 915 1297 916
rect 1291 911 1292 915
rect 1296 914 1297 915
rect 1322 915 1328 916
rect 1322 914 1323 915
rect 1296 912 1323 914
rect 1296 911 1297 912
rect 1291 910 1297 911
rect 1322 911 1323 912
rect 1327 911 1328 915
rect 1322 910 1328 911
rect 1467 915 1473 916
rect 1467 911 1468 915
rect 1472 914 1473 915
rect 1498 915 1504 916
rect 1498 914 1499 915
rect 1472 912 1499 914
rect 1472 911 1473 912
rect 1467 910 1473 911
rect 1498 911 1499 912
rect 1503 911 1504 915
rect 1498 910 1504 911
rect 1610 915 1616 916
rect 1610 911 1611 915
rect 1615 914 1616 915
rect 1635 915 1641 916
rect 1635 914 1636 915
rect 1615 912 1636 914
rect 1615 911 1616 912
rect 1610 910 1616 911
rect 1635 911 1636 912
rect 1640 911 1641 915
rect 1803 913 1804 917
rect 1808 913 1809 917
rect 2760 916 2796 918
rect 1803 912 1809 913
rect 1826 915 1832 916
rect 1635 910 1641 911
rect 1826 911 1827 915
rect 1831 914 1832 915
rect 1955 915 1961 916
rect 1955 914 1956 915
rect 1831 912 1956 914
rect 1831 911 1832 912
rect 1826 910 1832 911
rect 1955 911 1956 912
rect 1960 911 1961 915
rect 1955 910 1961 911
rect 2699 915 2705 916
rect 2699 911 2700 915
rect 2704 914 2705 915
rect 2750 915 2756 916
rect 2750 914 2751 915
rect 2704 912 2751 914
rect 2704 911 2705 912
rect 2699 910 2705 911
rect 2750 911 2751 912
rect 2755 911 2756 915
rect 2795 915 2796 916
rect 2800 915 2801 919
rect 2795 914 2801 915
rect 2818 919 2824 920
rect 2818 915 2819 919
rect 2823 918 2824 919
rect 2899 919 2905 920
rect 2899 918 2900 919
rect 2823 916 2900 918
rect 2823 915 2824 916
rect 2818 914 2824 915
rect 2899 915 2900 916
rect 2904 915 2905 919
rect 2899 914 2905 915
rect 3019 919 3025 920
rect 3019 915 3020 919
rect 3024 918 3025 919
rect 3074 919 3080 920
rect 3074 918 3075 919
rect 3024 916 3075 918
rect 3024 915 3025 916
rect 3019 914 3025 915
rect 3074 915 3075 916
rect 3079 915 3080 919
rect 3074 914 3080 915
rect 3086 919 3092 920
rect 3086 915 3087 919
rect 3091 918 3092 919
rect 3163 919 3169 920
rect 3163 918 3164 919
rect 3091 916 3164 918
rect 3091 915 3092 916
rect 3086 914 3092 915
rect 3163 915 3164 916
rect 3168 915 3169 919
rect 3163 914 3169 915
rect 3186 919 3192 920
rect 3186 915 3187 919
rect 3191 918 3192 919
rect 3331 919 3337 920
rect 3331 918 3332 919
rect 3191 916 3332 918
rect 3191 915 3192 916
rect 3186 914 3192 915
rect 3331 915 3332 916
rect 3336 915 3337 919
rect 3331 914 3337 915
rect 3354 919 3360 920
rect 3354 915 3355 919
rect 3359 918 3360 919
rect 3515 919 3521 920
rect 3515 918 3516 919
rect 3359 916 3516 918
rect 3359 915 3360 916
rect 3354 914 3360 915
rect 3515 915 3516 916
rect 3520 915 3521 919
rect 3515 914 3521 915
rect 3538 919 3544 920
rect 3538 915 3539 919
rect 3543 918 3544 919
rect 3715 919 3721 920
rect 3715 918 3716 919
rect 3543 916 3716 918
rect 3543 915 3544 916
rect 3538 914 3544 915
rect 3715 915 3716 916
rect 3720 915 3721 919
rect 3715 914 3721 915
rect 3891 915 3897 916
rect 2750 910 2756 911
rect 3891 911 3892 915
rect 3896 914 3897 915
rect 3906 915 3912 916
rect 3906 914 3907 915
rect 3896 912 3907 914
rect 3896 911 3897 912
rect 3891 910 3897 911
rect 3906 911 3907 912
rect 3911 911 3912 915
rect 3906 910 3912 911
rect 3622 899 3628 900
rect 3622 898 3623 899
rect 3180 896 3623 898
rect 3180 894 3182 896
rect 3622 895 3623 896
rect 3627 895 3628 899
rect 3622 894 3628 895
rect 3179 893 3185 894
rect 134 892 140 893
rect 110 889 116 890
rect 110 885 111 889
rect 115 885 116 889
rect 134 888 135 892
rect 139 888 140 892
rect 134 887 140 888
rect 270 892 276 893
rect 270 888 271 892
rect 275 888 276 892
rect 270 887 276 888
rect 454 892 460 893
rect 454 888 455 892
rect 459 888 460 892
rect 454 887 460 888
rect 654 892 660 893
rect 654 888 655 892
rect 659 888 660 892
rect 654 887 660 888
rect 854 892 860 893
rect 854 888 855 892
rect 859 888 860 892
rect 854 887 860 888
rect 1054 892 1060 893
rect 1054 888 1055 892
rect 1059 888 1060 892
rect 1054 887 1060 888
rect 1238 892 1244 893
rect 1238 888 1239 892
rect 1243 888 1244 892
rect 1238 887 1244 888
rect 1414 892 1420 893
rect 1414 888 1415 892
rect 1419 888 1420 892
rect 1414 887 1420 888
rect 1582 892 1588 893
rect 1582 888 1583 892
rect 1587 888 1588 892
rect 1582 887 1588 888
rect 1750 892 1756 893
rect 1750 888 1751 892
rect 1755 888 1756 892
rect 1750 887 1756 888
rect 1902 892 1908 893
rect 1902 888 1903 892
rect 1907 888 1908 892
rect 2146 891 2152 892
rect 1902 887 1908 888
rect 2006 889 2012 890
rect 110 884 116 885
rect 2006 885 2007 889
rect 2011 885 2012 889
rect 2006 884 2012 885
rect 2123 889 2129 890
rect 2123 885 2124 889
rect 2128 885 2129 889
rect 2146 887 2147 891
rect 2151 890 2152 891
rect 2307 891 2313 892
rect 2307 890 2308 891
rect 2151 888 2308 890
rect 2151 887 2152 888
rect 2146 886 2152 887
rect 2307 887 2308 888
rect 2312 887 2313 891
rect 2307 886 2313 887
rect 2330 891 2336 892
rect 2330 887 2331 891
rect 2335 890 2336 891
rect 2515 891 2521 892
rect 2515 890 2516 891
rect 2335 888 2516 890
rect 2335 887 2336 888
rect 2330 886 2336 887
rect 2515 887 2516 888
rect 2520 887 2521 891
rect 2515 886 2521 887
rect 2731 891 2737 892
rect 2731 887 2732 891
rect 2736 890 2737 891
rect 2783 891 2789 892
rect 2783 890 2784 891
rect 2736 888 2784 890
rect 2736 887 2737 888
rect 2731 886 2737 887
rect 2783 887 2784 888
rect 2788 887 2789 891
rect 2783 886 2789 887
rect 2947 889 2953 890
rect 2123 884 2129 885
rect 2947 885 2948 889
rect 2952 886 2953 889
rect 3179 889 3180 893
rect 3184 889 3185 893
rect 3179 888 3185 889
rect 3202 891 3208 892
rect 2970 887 2976 888
rect 2970 886 2971 887
rect 2952 885 2971 886
rect 2947 884 2971 885
rect 210 883 216 884
rect 210 879 211 883
rect 215 879 216 883
rect 210 878 216 879
rect 346 883 352 884
rect 346 879 347 883
rect 351 879 352 883
rect 346 878 352 879
rect 530 883 536 884
rect 530 879 531 883
rect 535 879 536 883
rect 530 878 536 879
rect 730 883 736 884
rect 730 879 731 883
rect 735 879 736 883
rect 730 878 736 879
rect 922 883 928 884
rect 922 879 923 883
rect 927 879 928 883
rect 1166 883 1172 884
rect 1166 882 1167 883
rect 1133 880 1167 882
rect 922 878 928 879
rect 1166 879 1167 880
rect 1171 879 1172 883
rect 1166 878 1172 879
rect 1230 883 1236 884
rect 1230 879 1231 883
rect 1235 882 1236 883
rect 1322 883 1328 884
rect 1235 880 1281 882
rect 1235 879 1236 880
rect 1230 878 1236 879
rect 1322 879 1323 883
rect 1327 882 1328 883
rect 1498 883 1504 884
rect 1327 880 1457 882
rect 1327 879 1328 880
rect 1322 878 1328 879
rect 1498 879 1499 883
rect 1503 882 1504 883
rect 1826 883 1832 884
rect 1503 880 1625 882
rect 1503 879 1504 880
rect 1498 878 1504 879
rect 1826 879 1827 883
rect 1831 879 1832 883
rect 2124 882 2126 884
rect 2970 883 2971 884
rect 2975 883 2976 887
rect 3202 887 3203 891
rect 3207 890 3208 891
rect 3419 891 3425 892
rect 3419 890 3420 891
rect 3207 888 3420 890
rect 3207 887 3208 888
rect 3202 886 3208 887
rect 3419 887 3420 888
rect 3424 887 3425 891
rect 3419 886 3425 887
rect 3442 891 3448 892
rect 3442 887 3443 891
rect 3447 890 3448 891
rect 3667 891 3673 892
rect 3667 890 3668 891
rect 3447 888 3668 890
rect 3447 887 3448 888
rect 3442 886 3448 887
rect 3667 887 3668 888
rect 3672 887 3673 891
rect 3667 886 3673 887
rect 3891 891 3897 892
rect 3891 887 3892 891
rect 3896 890 3897 891
rect 3914 891 3920 892
rect 3914 890 3915 891
rect 3896 888 3915 890
rect 3896 887 3897 888
rect 3891 886 3897 887
rect 3914 887 3915 888
rect 3919 887 3920 891
rect 3914 886 3920 887
rect 2970 882 2976 883
rect 1981 880 2126 882
rect 1826 878 1832 879
rect 134 873 140 874
rect 110 872 116 873
rect 110 868 111 872
rect 115 868 116 872
rect 134 869 135 873
rect 139 869 140 873
rect 134 868 140 869
rect 270 873 276 874
rect 270 869 271 873
rect 275 869 276 873
rect 270 868 276 869
rect 454 873 460 874
rect 454 869 455 873
rect 459 869 460 873
rect 454 868 460 869
rect 654 873 660 874
rect 654 869 655 873
rect 659 869 660 873
rect 654 868 660 869
rect 854 873 860 874
rect 854 869 855 873
rect 859 869 860 873
rect 854 868 860 869
rect 1054 873 1060 874
rect 1054 869 1055 873
rect 1059 869 1060 873
rect 1054 868 1060 869
rect 1238 873 1244 874
rect 1238 869 1239 873
rect 1243 869 1244 873
rect 1238 868 1244 869
rect 1414 873 1420 874
rect 1414 869 1415 873
rect 1419 869 1420 873
rect 1414 868 1420 869
rect 1582 873 1588 874
rect 1582 869 1583 873
rect 1587 869 1588 873
rect 1582 868 1588 869
rect 1750 873 1756 874
rect 1750 869 1751 873
rect 1755 869 1756 873
rect 1750 868 1756 869
rect 1902 873 1908 874
rect 1902 869 1903 873
rect 1907 869 1908 873
rect 1902 868 1908 869
rect 2006 872 2012 873
rect 2006 868 2007 872
rect 2011 868 2012 872
rect 110 867 116 868
rect 2006 867 2012 868
rect 2070 868 2076 869
rect 2046 865 2052 866
rect 2046 861 2047 865
rect 2051 861 2052 865
rect 2070 864 2071 868
rect 2075 864 2076 868
rect 2070 863 2076 864
rect 2254 868 2260 869
rect 2254 864 2255 868
rect 2259 864 2260 868
rect 2254 863 2260 864
rect 2462 868 2468 869
rect 2462 864 2463 868
rect 2467 864 2468 868
rect 2462 863 2468 864
rect 2678 868 2684 869
rect 2678 864 2679 868
rect 2683 864 2684 868
rect 2678 863 2684 864
rect 2894 868 2900 869
rect 2894 864 2895 868
rect 2899 864 2900 868
rect 2894 863 2900 864
rect 3126 868 3132 869
rect 3126 864 3127 868
rect 3131 864 3132 868
rect 3126 863 3132 864
rect 3366 868 3372 869
rect 3366 864 3367 868
rect 3371 864 3372 868
rect 3366 863 3372 864
rect 3614 868 3620 869
rect 3614 864 3615 868
rect 3619 864 3620 868
rect 3614 863 3620 864
rect 3838 868 3844 869
rect 3838 864 3839 868
rect 3843 864 3844 868
rect 3838 863 3844 864
rect 3942 865 3948 866
rect 2046 860 2052 861
rect 3942 861 3943 865
rect 3947 861 3948 865
rect 3942 860 3948 861
rect 2146 859 2152 860
rect 2146 855 2147 859
rect 2151 855 2152 859
rect 2146 854 2152 855
rect 2330 859 2336 860
rect 2330 855 2331 859
rect 2335 855 2336 859
rect 2330 854 2336 855
rect 2350 859 2356 860
rect 2350 855 2351 859
rect 2355 858 2356 859
rect 2750 859 2756 860
rect 2355 856 2505 858
rect 2355 855 2356 856
rect 2350 854 2356 855
rect 2750 855 2751 859
rect 2755 855 2756 859
rect 2750 854 2756 855
rect 2783 859 2789 860
rect 2783 855 2784 859
rect 2788 858 2789 859
rect 3202 859 3208 860
rect 2788 856 2937 858
rect 2788 855 2789 856
rect 2783 854 2789 855
rect 3202 855 3203 859
rect 3207 855 3208 859
rect 3202 854 3208 855
rect 3442 859 3448 860
rect 3442 855 3443 859
rect 3447 855 3448 859
rect 3442 854 3448 855
rect 3690 859 3696 860
rect 3690 855 3691 859
rect 3695 855 3696 859
rect 3690 854 3696 855
rect 3906 859 3912 860
rect 3906 855 3907 859
rect 3911 855 3912 859
rect 3906 854 3912 855
rect 2070 849 2076 850
rect 2046 848 2052 849
rect 2046 844 2047 848
rect 2051 844 2052 848
rect 2070 845 2071 849
rect 2075 845 2076 849
rect 2070 844 2076 845
rect 2254 849 2260 850
rect 2254 845 2255 849
rect 2259 845 2260 849
rect 2254 844 2260 845
rect 2462 849 2468 850
rect 2462 845 2463 849
rect 2467 845 2468 849
rect 2462 844 2468 845
rect 2678 849 2684 850
rect 2678 845 2679 849
rect 2683 845 2684 849
rect 2678 844 2684 845
rect 2894 849 2900 850
rect 2894 845 2895 849
rect 2899 845 2900 849
rect 2894 844 2900 845
rect 3126 849 3132 850
rect 3126 845 3127 849
rect 3131 845 3132 849
rect 3126 844 3132 845
rect 3366 849 3372 850
rect 3366 845 3367 849
rect 3371 845 3372 849
rect 3366 844 3372 845
rect 3614 849 3620 850
rect 3614 845 3615 849
rect 3619 845 3620 849
rect 3614 844 3620 845
rect 3838 849 3844 850
rect 3838 845 3839 849
rect 3843 845 3844 849
rect 3838 844 3844 845
rect 3942 848 3948 849
rect 3942 844 3943 848
rect 3947 844 3948 848
rect 2046 843 2052 844
rect 3942 843 3948 844
rect 110 820 116 821
rect 2006 820 2012 821
rect 110 816 111 820
rect 115 816 116 820
rect 110 815 116 816
rect 214 819 220 820
rect 214 815 215 819
rect 219 815 220 819
rect 214 814 220 815
rect 342 819 348 820
rect 342 815 343 819
rect 347 815 348 819
rect 342 814 348 815
rect 494 819 500 820
rect 494 815 495 819
rect 499 815 500 819
rect 494 814 500 815
rect 654 819 660 820
rect 654 815 655 819
rect 659 815 660 819
rect 654 814 660 815
rect 830 819 836 820
rect 830 815 831 819
rect 835 815 836 819
rect 830 814 836 815
rect 1006 819 1012 820
rect 1006 815 1007 819
rect 1011 815 1012 819
rect 1006 814 1012 815
rect 1182 819 1188 820
rect 1182 815 1183 819
rect 1187 815 1188 819
rect 1182 814 1188 815
rect 1358 819 1364 820
rect 1358 815 1359 819
rect 1363 815 1364 819
rect 1358 814 1364 815
rect 1534 819 1540 820
rect 1534 815 1535 819
rect 1539 815 1540 819
rect 1534 814 1540 815
rect 1718 819 1724 820
rect 1718 815 1719 819
rect 1723 815 1724 819
rect 2006 816 2007 820
rect 2011 816 2012 820
rect 2006 815 2012 816
rect 1718 814 1724 815
rect 190 811 196 812
rect 190 807 191 811
rect 195 810 196 811
rect 330 811 336 812
rect 195 808 257 810
rect 195 807 196 808
rect 190 806 196 807
rect 330 807 331 811
rect 335 810 336 811
rect 431 811 437 812
rect 335 808 385 810
rect 335 807 336 808
rect 330 806 336 807
rect 431 807 432 811
rect 436 810 437 811
rect 614 811 620 812
rect 436 808 537 810
rect 436 807 437 808
rect 431 806 437 807
rect 614 807 615 811
rect 619 810 620 811
rect 791 811 797 812
rect 619 808 697 810
rect 619 807 620 808
rect 614 806 620 807
rect 791 807 792 811
rect 796 810 797 811
rect 1094 811 1100 812
rect 796 808 873 810
rect 796 807 797 808
rect 791 806 797 807
rect 1082 807 1088 808
rect 110 803 116 804
rect 110 799 111 803
rect 115 799 116 803
rect 1082 803 1083 807
rect 1087 803 1088 807
rect 1094 807 1095 811
rect 1099 810 1100 811
rect 1610 811 1616 812
rect 1099 808 1225 810
rect 1099 807 1100 808
rect 1094 806 1100 807
rect 1462 807 1468 808
rect 1462 806 1463 807
rect 1437 804 1463 806
rect 1082 802 1088 803
rect 1462 803 1463 804
rect 1467 803 1468 807
rect 1610 807 1611 811
rect 1615 807 1616 811
rect 1610 806 1616 807
rect 1638 811 1644 812
rect 1638 807 1639 811
rect 1643 810 1644 811
rect 1643 808 1761 810
rect 1643 807 1644 808
rect 1638 806 1644 807
rect 1462 802 1468 803
rect 2006 803 2012 804
rect 110 798 116 799
rect 214 800 220 801
rect 214 796 215 800
rect 219 796 220 800
rect 214 795 220 796
rect 342 800 348 801
rect 342 796 343 800
rect 347 796 348 800
rect 342 795 348 796
rect 494 800 500 801
rect 494 796 495 800
rect 499 796 500 800
rect 494 795 500 796
rect 654 800 660 801
rect 654 796 655 800
rect 659 796 660 800
rect 654 795 660 796
rect 830 800 836 801
rect 830 796 831 800
rect 835 796 836 800
rect 830 795 836 796
rect 1006 800 1012 801
rect 1006 796 1007 800
rect 1011 796 1012 800
rect 1006 795 1012 796
rect 1182 800 1188 801
rect 1182 796 1183 800
rect 1187 796 1188 800
rect 1182 795 1188 796
rect 1358 800 1364 801
rect 1358 796 1359 800
rect 1363 796 1364 800
rect 1358 795 1364 796
rect 1534 800 1540 801
rect 1534 796 1535 800
rect 1539 796 1540 800
rect 1534 795 1540 796
rect 1718 800 1724 801
rect 1718 796 1719 800
rect 1723 796 1724 800
rect 2006 799 2007 803
rect 2011 799 2012 803
rect 2006 798 2012 799
rect 1718 795 1724 796
rect 2046 796 2052 797
rect 3942 796 3948 797
rect 2046 792 2047 796
rect 2051 792 2052 796
rect 2046 791 2052 792
rect 2214 795 2220 796
rect 2214 791 2215 795
rect 2219 791 2220 795
rect 2214 790 2220 791
rect 2326 795 2332 796
rect 2326 791 2327 795
rect 2331 791 2332 795
rect 2326 790 2332 791
rect 2446 795 2452 796
rect 2446 791 2447 795
rect 2451 791 2452 795
rect 2446 790 2452 791
rect 2582 795 2588 796
rect 2582 791 2583 795
rect 2587 791 2588 795
rect 2582 790 2588 791
rect 2734 795 2740 796
rect 2734 791 2735 795
rect 2739 791 2740 795
rect 2734 790 2740 791
rect 2894 795 2900 796
rect 2894 791 2895 795
rect 2899 791 2900 795
rect 2894 790 2900 791
rect 3062 795 3068 796
rect 3062 791 3063 795
rect 3067 791 3068 795
rect 3062 790 3068 791
rect 3246 795 3252 796
rect 3246 791 3247 795
rect 3251 791 3252 795
rect 3246 790 3252 791
rect 3446 795 3452 796
rect 3446 791 3447 795
rect 3451 791 3452 795
rect 3446 790 3452 791
rect 3654 795 3660 796
rect 3654 791 3655 795
rect 3659 791 3660 795
rect 3654 790 3660 791
rect 3838 795 3844 796
rect 3838 791 3839 795
rect 3843 791 3844 795
rect 3942 792 3943 796
rect 3947 792 3948 796
rect 3942 791 3948 792
rect 3838 790 3844 791
rect 1638 787 1644 788
rect 1638 786 1639 787
rect 1519 784 1639 786
rect 1519 782 1521 784
rect 1638 783 1639 784
rect 1643 783 1644 787
rect 2970 787 2976 788
rect 1638 782 1644 783
rect 2290 783 2296 784
rect 1456 780 1521 782
rect 267 779 273 780
rect 267 775 268 779
rect 272 778 273 779
rect 330 779 336 780
rect 330 778 331 779
rect 272 776 331 778
rect 272 775 273 776
rect 267 774 273 775
rect 330 775 331 776
rect 335 775 336 779
rect 330 774 336 775
rect 395 779 401 780
rect 395 775 396 779
rect 400 778 401 779
rect 431 779 437 780
rect 431 778 432 779
rect 400 776 432 778
rect 400 775 401 776
rect 395 774 401 775
rect 431 775 432 776
rect 436 775 437 779
rect 431 774 437 775
rect 547 779 553 780
rect 547 775 548 779
rect 552 778 553 779
rect 614 779 620 780
rect 614 778 615 779
rect 552 776 615 778
rect 552 775 553 776
rect 547 774 553 775
rect 614 775 615 776
rect 619 775 620 779
rect 614 774 620 775
rect 707 779 713 780
rect 707 775 708 779
rect 712 778 713 779
rect 791 779 797 780
rect 791 778 792 779
rect 712 776 792 778
rect 712 775 713 776
rect 707 774 713 775
rect 791 775 792 776
rect 796 775 797 779
rect 1059 779 1065 780
rect 791 774 797 775
rect 878 775 889 776
rect 878 771 879 775
rect 883 771 884 775
rect 888 771 889 775
rect 1059 775 1060 779
rect 1064 778 1065 779
rect 1094 779 1100 780
rect 1094 778 1095 779
rect 1064 776 1095 778
rect 1064 775 1065 776
rect 1059 774 1065 775
rect 1094 775 1095 776
rect 1099 775 1100 779
rect 1094 774 1100 775
rect 1166 779 1172 780
rect 1166 775 1167 779
rect 1171 778 1172 779
rect 1235 779 1241 780
rect 1235 778 1236 779
rect 1171 776 1236 778
rect 1171 775 1172 776
rect 1166 774 1172 775
rect 1235 775 1236 776
rect 1240 775 1241 779
rect 1235 774 1241 775
rect 1411 779 1417 780
rect 1411 775 1412 779
rect 1416 778 1417 779
rect 1456 778 1458 780
rect 1587 779 1593 780
rect 1587 778 1588 779
rect 1416 776 1458 778
rect 1519 776 1588 778
rect 1416 775 1417 776
rect 1411 774 1417 775
rect 1462 775 1468 776
rect 878 770 889 771
rect 1462 771 1463 775
rect 1467 774 1468 775
rect 1519 774 1521 776
rect 1587 775 1588 776
rect 1592 775 1593 779
rect 2046 779 2052 780
rect 1587 774 1593 775
rect 1674 775 1680 776
rect 1467 772 1521 774
rect 1467 771 1468 772
rect 1462 770 1468 771
rect 1674 771 1675 775
rect 1679 774 1680 775
rect 1771 775 1777 776
rect 1771 774 1772 775
rect 1679 772 1772 774
rect 1679 771 1680 772
rect 1674 770 1680 771
rect 1771 771 1772 772
rect 1776 771 1777 775
rect 2046 775 2047 779
rect 2051 775 2052 779
rect 2290 779 2291 783
rect 2295 779 2296 783
rect 2290 778 2296 779
rect 2402 783 2408 784
rect 2402 779 2403 783
rect 2407 779 2408 783
rect 2402 778 2408 779
rect 2522 783 2528 784
rect 2522 779 2523 783
rect 2527 779 2528 783
rect 2522 778 2528 779
rect 2658 783 2664 784
rect 2658 779 2659 783
rect 2663 779 2664 783
rect 2658 778 2664 779
rect 2810 783 2816 784
rect 2810 779 2811 783
rect 2815 779 2816 783
rect 2970 783 2971 787
rect 2975 783 2976 787
rect 2970 782 2976 783
rect 3023 787 3029 788
rect 3023 783 3024 787
rect 3028 786 3029 787
rect 3330 787 3336 788
rect 3028 784 3105 786
rect 3028 783 3029 784
rect 3023 782 3029 783
rect 3322 783 3328 784
rect 2810 778 2816 779
rect 3322 779 3323 783
rect 3327 779 3328 783
rect 3330 783 3331 787
rect 3335 786 3336 787
rect 3530 787 3536 788
rect 3335 784 3489 786
rect 3335 783 3336 784
rect 3330 782 3336 783
rect 3530 783 3531 787
rect 3535 786 3536 787
rect 3914 787 3920 788
rect 3535 784 3697 786
rect 3535 783 3536 784
rect 3530 782 3536 783
rect 3914 783 3915 787
rect 3919 783 3920 787
rect 3914 782 3920 783
rect 3322 778 3328 779
rect 3942 779 3948 780
rect 2046 774 2052 775
rect 2214 776 2220 777
rect 2214 772 2215 776
rect 2219 772 2220 776
rect 2214 771 2220 772
rect 2326 776 2332 777
rect 2326 772 2327 776
rect 2331 772 2332 776
rect 2326 771 2332 772
rect 2446 776 2452 777
rect 2446 772 2447 776
rect 2451 772 2452 776
rect 2446 771 2452 772
rect 2582 776 2588 777
rect 2582 772 2583 776
rect 2587 772 2588 776
rect 2582 771 2588 772
rect 2734 776 2740 777
rect 2734 772 2735 776
rect 2739 772 2740 776
rect 2734 771 2740 772
rect 2894 776 2900 777
rect 2894 772 2895 776
rect 2899 772 2900 776
rect 2894 771 2900 772
rect 3062 776 3068 777
rect 3062 772 3063 776
rect 3067 772 3068 776
rect 3062 771 3068 772
rect 3246 776 3252 777
rect 3246 772 3247 776
rect 3251 772 3252 776
rect 3246 771 3252 772
rect 3446 776 3452 777
rect 3446 772 3447 776
rect 3451 772 3452 776
rect 3446 771 3452 772
rect 3654 776 3660 777
rect 3654 772 3655 776
rect 3659 772 3660 776
rect 3654 771 3660 772
rect 3838 776 3844 777
rect 3838 772 3839 776
rect 3843 772 3844 776
rect 3942 775 3943 779
rect 3947 775 3948 779
rect 3942 774 3948 775
rect 3838 771 3844 772
rect 1771 770 1777 771
rect 450 763 456 764
rect 427 761 433 762
rect 427 757 428 761
rect 432 757 433 761
rect 450 759 451 763
rect 455 762 456 763
rect 547 763 553 764
rect 547 762 548 763
rect 455 760 548 762
rect 455 759 456 760
rect 450 758 456 759
rect 547 759 548 760
rect 552 759 553 763
rect 547 758 553 759
rect 570 763 576 764
rect 570 759 571 763
rect 575 762 576 763
rect 675 763 681 764
rect 675 762 676 763
rect 575 760 676 762
rect 575 759 576 760
rect 570 758 576 759
rect 675 759 676 760
rect 680 759 681 763
rect 675 758 681 759
rect 803 763 809 764
rect 803 759 804 763
rect 808 762 809 763
rect 818 763 824 764
rect 818 762 819 763
rect 808 760 819 762
rect 808 759 809 760
rect 803 758 809 759
rect 818 759 819 760
rect 823 759 824 763
rect 1075 763 1084 764
rect 818 758 824 759
rect 939 761 945 762
rect 427 756 433 757
rect 939 757 940 761
rect 944 757 945 761
rect 1075 759 1076 763
rect 1083 759 1084 763
rect 1075 758 1084 759
rect 1098 763 1104 764
rect 1098 759 1099 763
rect 1103 762 1104 763
rect 1219 763 1225 764
rect 1219 762 1220 763
rect 1103 760 1220 762
rect 1103 759 1104 760
rect 1098 758 1104 759
rect 1219 759 1220 760
rect 1224 759 1225 763
rect 1219 758 1225 759
rect 1363 763 1372 764
rect 1363 759 1364 763
rect 1371 759 1372 763
rect 1363 758 1372 759
rect 1386 763 1392 764
rect 1386 759 1387 763
rect 1391 762 1392 763
rect 1507 763 1513 764
rect 1507 762 1508 763
rect 1391 760 1508 762
rect 1391 759 1392 760
rect 1386 758 1392 759
rect 1507 759 1508 760
rect 1512 759 1513 763
rect 1507 758 1513 759
rect 1591 763 1597 764
rect 1591 759 1592 763
rect 1596 762 1597 763
rect 1651 763 1657 764
rect 1651 762 1652 763
rect 1596 760 1652 762
rect 1596 759 1597 760
rect 1591 758 1597 759
rect 1651 759 1652 760
rect 1656 759 1657 763
rect 2350 763 2356 764
rect 2350 762 2351 763
rect 1651 758 1657 759
rect 2284 760 2351 762
rect 939 756 945 757
rect 428 746 430 756
rect 698 755 704 756
rect 698 751 699 755
rect 703 754 704 755
rect 940 754 942 756
rect 703 752 942 754
rect 2267 755 2273 756
rect 703 751 704 752
rect 698 750 704 751
rect 2267 751 2268 755
rect 2272 754 2273 755
rect 2284 754 2286 760
rect 2350 759 2351 760
rect 2355 759 2356 763
rect 2350 758 2356 759
rect 2272 752 2286 754
rect 2290 755 2296 756
rect 2272 751 2273 752
rect 2267 750 2273 751
rect 2290 751 2291 755
rect 2295 754 2296 755
rect 2379 755 2385 756
rect 2379 754 2380 755
rect 2295 752 2380 754
rect 2295 751 2296 752
rect 2290 750 2296 751
rect 2379 751 2380 752
rect 2384 751 2385 755
rect 2379 750 2385 751
rect 2402 755 2408 756
rect 2402 751 2403 755
rect 2407 754 2408 755
rect 2499 755 2505 756
rect 2499 754 2500 755
rect 2407 752 2500 754
rect 2407 751 2408 752
rect 2402 750 2408 751
rect 2499 751 2500 752
rect 2504 751 2505 755
rect 2499 750 2505 751
rect 2522 755 2528 756
rect 2522 751 2523 755
rect 2527 754 2528 755
rect 2635 755 2641 756
rect 2635 754 2636 755
rect 2527 752 2636 754
rect 2527 751 2528 752
rect 2522 750 2528 751
rect 2635 751 2636 752
rect 2640 751 2641 755
rect 2635 750 2641 751
rect 2658 755 2664 756
rect 2658 751 2659 755
rect 2663 754 2664 755
rect 2787 755 2793 756
rect 2787 754 2788 755
rect 2663 752 2788 754
rect 2663 751 2664 752
rect 2658 750 2664 751
rect 2787 751 2788 752
rect 2792 751 2793 755
rect 2787 750 2793 751
rect 2947 755 2953 756
rect 2947 751 2948 755
rect 2952 754 2953 755
rect 3023 755 3029 756
rect 3023 754 3024 755
rect 2952 752 3024 754
rect 2952 751 2953 752
rect 2947 750 2953 751
rect 3023 751 3024 752
rect 3028 751 3029 755
rect 3299 755 3305 756
rect 3023 750 3029 751
rect 3115 751 3121 752
rect 3115 747 3116 751
rect 3120 750 3121 751
rect 3130 751 3136 752
rect 3130 750 3131 751
rect 3120 748 3131 750
rect 3120 747 3121 748
rect 3115 746 3121 747
rect 3130 747 3131 748
rect 3135 747 3136 751
rect 3299 751 3300 755
rect 3304 754 3305 755
rect 3330 755 3336 756
rect 3330 754 3331 755
rect 3304 752 3331 754
rect 3304 751 3305 752
rect 3299 750 3305 751
rect 3330 751 3331 752
rect 3335 751 3336 755
rect 3330 750 3336 751
rect 3499 755 3505 756
rect 3499 751 3500 755
rect 3504 754 3505 755
rect 3530 755 3536 756
rect 3530 754 3531 755
rect 3504 752 3531 754
rect 3504 751 3505 752
rect 3499 750 3505 751
rect 3530 751 3531 752
rect 3535 751 3536 755
rect 3530 750 3536 751
rect 3690 755 3696 756
rect 3690 751 3691 755
rect 3695 754 3696 755
rect 3707 755 3713 756
rect 3707 754 3708 755
rect 3695 752 3708 754
rect 3695 751 3696 752
rect 3690 750 3696 751
rect 3707 751 3708 752
rect 3712 751 3713 755
rect 3707 750 3713 751
rect 3891 751 3897 752
rect 3130 746 3136 747
rect 3891 747 3892 751
rect 3896 750 3897 751
rect 3906 751 3912 752
rect 3906 750 3907 751
rect 3896 748 3907 750
rect 3896 747 3897 748
rect 3891 746 3897 747
rect 3906 747 3907 748
rect 3911 747 3912 751
rect 3906 746 3912 747
rect 428 744 710 746
rect 374 740 380 741
rect 110 737 116 738
rect 110 733 111 737
rect 115 733 116 737
rect 374 736 375 740
rect 379 736 380 740
rect 374 735 380 736
rect 494 740 500 741
rect 494 736 495 740
rect 499 736 500 740
rect 494 735 500 736
rect 622 740 628 741
rect 622 736 623 740
rect 627 736 628 740
rect 622 735 628 736
rect 110 732 116 733
rect 450 731 456 732
rect 450 727 451 731
rect 455 727 456 731
rect 450 726 456 727
rect 570 731 576 732
rect 570 727 571 731
rect 575 727 576 731
rect 570 726 576 727
rect 698 731 704 732
rect 698 727 699 731
rect 703 727 704 731
rect 708 730 710 744
rect 750 740 756 741
rect 750 736 751 740
rect 755 736 756 740
rect 750 735 756 736
rect 886 740 892 741
rect 886 736 887 740
rect 891 736 892 740
rect 886 735 892 736
rect 1022 740 1028 741
rect 1022 736 1023 740
rect 1027 736 1028 740
rect 1022 735 1028 736
rect 1166 740 1172 741
rect 1166 736 1167 740
rect 1171 736 1172 740
rect 1166 735 1172 736
rect 1310 740 1316 741
rect 1310 736 1311 740
rect 1315 736 1316 740
rect 1310 735 1316 736
rect 1454 740 1460 741
rect 1454 736 1455 740
rect 1459 736 1460 740
rect 1454 735 1460 736
rect 1598 740 1604 741
rect 1598 736 1599 740
rect 1603 736 1604 740
rect 1598 735 1604 736
rect 2006 737 2012 738
rect 2006 733 2007 737
rect 2011 733 2012 737
rect 2466 735 2472 736
rect 2006 732 2012 733
rect 2427 733 2433 734
rect 878 731 884 732
rect 708 728 793 730
rect 698 726 704 727
rect 878 727 879 731
rect 883 730 884 731
rect 1098 731 1104 732
rect 883 728 929 730
rect 883 727 884 728
rect 878 726 884 727
rect 1098 727 1099 731
rect 1103 727 1104 731
rect 1098 726 1104 727
rect 1234 731 1240 732
rect 1234 727 1235 731
rect 1239 727 1240 731
rect 1234 726 1240 727
rect 1386 731 1392 732
rect 1386 727 1387 731
rect 1391 727 1392 731
rect 1591 731 1597 732
rect 1591 730 1592 731
rect 1533 728 1592 730
rect 1386 726 1392 727
rect 1591 727 1592 728
rect 1596 727 1597 731
rect 1591 726 1597 727
rect 1674 731 1680 732
rect 1674 727 1675 731
rect 1679 727 1680 731
rect 2427 729 2428 733
rect 2432 729 2433 733
rect 2466 731 2467 735
rect 2471 734 2472 735
rect 2547 735 2553 736
rect 2547 734 2548 735
rect 2471 732 2548 734
rect 2471 731 2472 732
rect 2466 730 2472 731
rect 2547 731 2548 732
rect 2552 731 2553 735
rect 2810 735 2816 736
rect 2547 730 2553 731
rect 2675 733 2681 734
rect 2427 728 2433 729
rect 2675 729 2676 733
rect 2680 729 2681 733
rect 2810 731 2811 735
rect 2815 734 2816 735
rect 2819 735 2825 736
rect 2819 734 2820 735
rect 2815 732 2820 734
rect 2815 731 2816 732
rect 2810 730 2816 731
rect 2819 731 2820 732
rect 2824 731 2825 735
rect 2819 730 2825 731
rect 2842 735 2848 736
rect 2842 731 2843 735
rect 2847 734 2848 735
rect 2963 735 2969 736
rect 2963 734 2964 735
rect 2847 732 2964 734
rect 2847 731 2848 732
rect 2842 730 2848 731
rect 2963 731 2964 732
rect 2968 731 2969 735
rect 2963 730 2969 731
rect 3115 735 3124 736
rect 3115 731 3116 735
rect 3123 731 3124 735
rect 3115 730 3124 731
rect 3267 735 3273 736
rect 3267 731 3268 735
rect 3272 734 3273 735
rect 3322 735 3328 736
rect 3322 734 3323 735
rect 3272 732 3323 734
rect 3272 731 3273 732
rect 3267 730 3273 731
rect 3322 731 3323 732
rect 3327 731 3328 735
rect 3322 730 3328 731
rect 3335 735 3341 736
rect 3335 731 3336 735
rect 3340 734 3341 735
rect 3419 735 3425 736
rect 3419 734 3420 735
rect 3340 732 3420 734
rect 3340 731 3341 732
rect 3335 730 3341 731
rect 3419 731 3420 732
rect 3424 731 3425 735
rect 3419 730 3425 731
rect 3487 735 3493 736
rect 3487 731 3488 735
rect 3492 734 3493 735
rect 3571 735 3577 736
rect 3571 734 3572 735
rect 3492 732 3572 734
rect 3492 731 3493 732
rect 3487 730 3493 731
rect 3571 731 3572 732
rect 3576 731 3577 735
rect 3571 730 3577 731
rect 3594 735 3600 736
rect 3594 731 3595 735
rect 3599 734 3600 735
rect 3731 735 3737 736
rect 3731 734 3732 735
rect 3599 732 3732 734
rect 3599 731 3600 732
rect 3594 730 3600 731
rect 3731 731 3732 732
rect 3736 731 3737 735
rect 3731 730 3737 731
rect 3891 735 3900 736
rect 3891 731 3892 735
rect 3899 731 3900 735
rect 3891 730 3900 731
rect 2675 728 2681 729
rect 1674 726 1680 727
rect 2428 726 2430 728
rect 2590 727 2596 728
rect 2590 726 2591 727
rect 2428 724 2591 726
rect 2590 723 2591 724
rect 2595 723 2596 727
rect 2676 726 2678 728
rect 2882 727 2888 728
rect 2882 726 2883 727
rect 2676 724 2883 726
rect 2590 722 2596 723
rect 2882 723 2883 724
rect 2887 723 2888 727
rect 2882 722 2888 723
rect 374 721 380 722
rect 110 720 116 721
rect 110 716 111 720
rect 115 716 116 720
rect 374 717 375 721
rect 379 717 380 721
rect 374 716 380 717
rect 494 721 500 722
rect 494 717 495 721
rect 499 717 500 721
rect 494 716 500 717
rect 622 721 628 722
rect 622 717 623 721
rect 627 717 628 721
rect 622 716 628 717
rect 750 721 756 722
rect 750 717 751 721
rect 755 717 756 721
rect 750 716 756 717
rect 886 721 892 722
rect 886 717 887 721
rect 891 717 892 721
rect 886 716 892 717
rect 1022 721 1028 722
rect 1022 717 1023 721
rect 1027 717 1028 721
rect 1022 716 1028 717
rect 1166 721 1172 722
rect 1166 717 1167 721
rect 1171 717 1172 721
rect 1166 716 1172 717
rect 1310 721 1316 722
rect 1310 717 1311 721
rect 1315 717 1316 721
rect 1310 716 1316 717
rect 1454 721 1460 722
rect 1454 717 1455 721
rect 1459 717 1460 721
rect 1454 716 1460 717
rect 1598 721 1604 722
rect 1598 717 1599 721
rect 1603 717 1604 721
rect 1598 716 1604 717
rect 2006 720 2012 721
rect 2006 716 2007 720
rect 2011 716 2012 720
rect 110 715 116 716
rect 2006 715 2012 716
rect 2374 712 2380 713
rect 2046 709 2052 710
rect 2046 705 2047 709
rect 2051 705 2052 709
rect 2374 708 2375 712
rect 2379 708 2380 712
rect 2374 707 2380 708
rect 2494 712 2500 713
rect 2494 708 2495 712
rect 2499 708 2500 712
rect 2494 707 2500 708
rect 2622 712 2628 713
rect 2622 708 2623 712
rect 2627 708 2628 712
rect 2622 707 2628 708
rect 2766 712 2772 713
rect 2766 708 2767 712
rect 2771 708 2772 712
rect 2766 707 2772 708
rect 2910 712 2916 713
rect 2910 708 2911 712
rect 2915 708 2916 712
rect 2910 707 2916 708
rect 3062 712 3068 713
rect 3062 708 3063 712
rect 3067 708 3068 712
rect 3062 707 3068 708
rect 3214 712 3220 713
rect 3214 708 3215 712
rect 3219 708 3220 712
rect 3214 707 3220 708
rect 3366 712 3372 713
rect 3366 708 3367 712
rect 3371 708 3372 712
rect 3366 707 3372 708
rect 3518 712 3524 713
rect 3518 708 3519 712
rect 3523 708 3524 712
rect 3518 707 3524 708
rect 3678 712 3684 713
rect 3678 708 3679 712
rect 3683 708 3684 712
rect 3678 707 3684 708
rect 3838 712 3844 713
rect 3838 708 3839 712
rect 3843 708 3844 712
rect 3838 707 3844 708
rect 3942 709 3948 710
rect 2046 704 2052 705
rect 3942 705 3943 709
rect 3947 705 3948 709
rect 3942 704 3948 705
rect 2466 703 2472 704
rect 2466 702 2467 703
rect 2453 700 2467 702
rect 2466 699 2467 700
rect 2471 699 2472 703
rect 2582 703 2588 704
rect 2582 702 2583 703
rect 2573 700 2583 702
rect 2466 698 2472 699
rect 2582 699 2583 700
rect 2587 699 2588 703
rect 2582 698 2588 699
rect 2590 703 2596 704
rect 2590 699 2591 703
rect 2595 702 2596 703
rect 2842 703 2848 704
rect 2595 700 2665 702
rect 2595 699 2596 700
rect 2590 698 2596 699
rect 2842 699 2843 703
rect 2847 699 2848 703
rect 2842 698 2848 699
rect 2882 703 2888 704
rect 2882 699 2883 703
rect 2887 702 2888 703
rect 3130 703 3136 704
rect 2887 700 2953 702
rect 2887 699 2888 700
rect 2882 698 2888 699
rect 3130 699 3131 703
rect 3135 699 3136 703
rect 3335 703 3341 704
rect 3335 702 3336 703
rect 3293 700 3336 702
rect 3130 698 3136 699
rect 3335 699 3336 700
rect 3340 699 3341 703
rect 3487 703 3493 704
rect 3487 702 3488 703
rect 3445 700 3488 702
rect 3335 698 3341 699
rect 3487 699 3488 700
rect 3492 699 3493 703
rect 3487 698 3493 699
rect 3594 703 3600 704
rect 3594 699 3595 703
rect 3599 699 3600 703
rect 3594 698 3600 699
rect 3746 703 3752 704
rect 3746 699 3747 703
rect 3751 699 3752 703
rect 3746 698 3752 699
rect 3906 703 3912 704
rect 3906 699 3907 703
rect 3911 699 3912 703
rect 3906 698 3912 699
rect 2374 693 2380 694
rect 2046 692 2052 693
rect 2046 688 2047 692
rect 2051 688 2052 692
rect 2374 689 2375 693
rect 2379 689 2380 693
rect 2374 688 2380 689
rect 2494 693 2500 694
rect 2494 689 2495 693
rect 2499 689 2500 693
rect 2494 688 2500 689
rect 2622 693 2628 694
rect 2622 689 2623 693
rect 2627 689 2628 693
rect 2622 688 2628 689
rect 2766 693 2772 694
rect 2766 689 2767 693
rect 2771 689 2772 693
rect 2766 688 2772 689
rect 2910 693 2916 694
rect 2910 689 2911 693
rect 2915 689 2916 693
rect 2910 688 2916 689
rect 3062 693 3068 694
rect 3062 689 3063 693
rect 3067 689 3068 693
rect 3062 688 3068 689
rect 3214 693 3220 694
rect 3214 689 3215 693
rect 3219 689 3220 693
rect 3214 688 3220 689
rect 3366 693 3372 694
rect 3366 689 3367 693
rect 3371 689 3372 693
rect 3366 688 3372 689
rect 3518 693 3524 694
rect 3518 689 3519 693
rect 3523 689 3524 693
rect 3518 688 3524 689
rect 3678 693 3684 694
rect 3678 689 3679 693
rect 3683 689 3684 693
rect 3678 688 3684 689
rect 3838 693 3844 694
rect 3838 689 3839 693
rect 3843 689 3844 693
rect 3838 688 3844 689
rect 3942 692 3948 693
rect 3942 688 3943 692
rect 3947 688 3948 692
rect 2046 687 2052 688
rect 3942 687 3948 688
rect 110 668 116 669
rect 2006 668 2012 669
rect 110 664 111 668
rect 115 664 116 668
rect 110 663 116 664
rect 526 667 532 668
rect 526 663 527 667
rect 531 663 532 667
rect 526 662 532 663
rect 630 667 636 668
rect 630 663 631 667
rect 635 663 636 667
rect 630 662 636 663
rect 742 667 748 668
rect 742 663 743 667
rect 747 663 748 667
rect 742 662 748 663
rect 854 667 860 668
rect 854 663 855 667
rect 859 663 860 667
rect 854 662 860 663
rect 966 667 972 668
rect 966 663 967 667
rect 971 663 972 667
rect 966 662 972 663
rect 1070 667 1076 668
rect 1070 663 1071 667
rect 1075 663 1076 667
rect 1070 662 1076 663
rect 1182 667 1188 668
rect 1182 663 1183 667
rect 1187 663 1188 667
rect 1182 662 1188 663
rect 1294 667 1300 668
rect 1294 663 1295 667
rect 1299 663 1300 667
rect 1294 662 1300 663
rect 1406 667 1412 668
rect 1406 663 1407 667
rect 1411 663 1412 667
rect 1406 662 1412 663
rect 1518 667 1524 668
rect 1518 663 1519 667
rect 1523 663 1524 667
rect 2006 664 2007 668
rect 2011 664 2012 668
rect 2006 663 2012 664
rect 1518 662 1524 663
rect 818 659 824 660
rect 602 655 608 656
rect 110 651 116 652
rect 110 647 111 651
rect 115 647 116 651
rect 602 651 603 655
rect 607 651 608 655
rect 602 650 608 651
rect 706 655 712 656
rect 706 651 707 655
rect 711 651 712 655
rect 818 655 819 659
rect 823 655 824 659
rect 818 654 824 655
rect 826 659 832 660
rect 826 655 827 659
rect 831 658 832 659
rect 959 659 965 660
rect 831 656 897 658
rect 831 655 832 656
rect 826 654 832 655
rect 959 655 960 659
rect 964 658 965 659
rect 1159 659 1165 660
rect 964 656 1009 658
rect 964 655 965 656
rect 959 654 965 655
rect 1146 655 1152 656
rect 706 650 712 651
rect 1146 651 1147 655
rect 1151 651 1152 655
rect 1159 655 1160 659
rect 1164 658 1165 659
rect 1370 659 1376 660
rect 1164 656 1225 658
rect 1164 655 1165 656
rect 1159 654 1165 655
rect 1370 655 1371 659
rect 1375 655 1376 659
rect 1370 654 1376 655
rect 1382 659 1388 660
rect 1382 655 1383 659
rect 1387 658 1388 659
rect 1490 659 1496 660
rect 1387 656 1449 658
rect 1387 655 1388 656
rect 1382 654 1388 655
rect 1490 655 1491 659
rect 1495 658 1496 659
rect 1495 656 1561 658
rect 1495 655 1496 656
rect 1490 654 1496 655
rect 1146 650 1152 651
rect 2006 651 2012 652
rect 110 646 116 647
rect 526 648 532 649
rect 526 644 527 648
rect 531 644 532 648
rect 526 643 532 644
rect 630 648 636 649
rect 630 644 631 648
rect 635 644 636 648
rect 630 643 636 644
rect 742 648 748 649
rect 742 644 743 648
rect 747 644 748 648
rect 742 643 748 644
rect 854 648 860 649
rect 854 644 855 648
rect 859 644 860 648
rect 854 643 860 644
rect 966 648 972 649
rect 966 644 967 648
rect 971 644 972 648
rect 966 643 972 644
rect 1070 648 1076 649
rect 1070 644 1071 648
rect 1075 644 1076 648
rect 1070 643 1076 644
rect 1182 648 1188 649
rect 1182 644 1183 648
rect 1187 644 1188 648
rect 1182 643 1188 644
rect 1294 648 1300 649
rect 1294 644 1295 648
rect 1299 644 1300 648
rect 1294 643 1300 644
rect 1406 648 1412 649
rect 1406 644 1407 648
rect 1411 644 1412 648
rect 1406 643 1412 644
rect 1518 648 1524 649
rect 1518 644 1519 648
rect 1523 644 1524 648
rect 2006 647 2007 651
rect 2011 647 2012 651
rect 2006 646 2012 647
rect 1518 643 1524 644
rect 826 635 832 636
rect 826 634 827 635
rect 596 632 827 634
rect 579 627 585 628
rect 579 623 580 627
rect 584 626 585 627
rect 596 626 598 632
rect 826 631 827 632
rect 831 631 832 635
rect 826 630 832 631
rect 2046 632 2052 633
rect 3942 632 3948 633
rect 2046 628 2047 632
rect 2051 628 2052 632
rect 584 624 598 626
rect 602 627 608 628
rect 584 623 585 624
rect 579 622 585 623
rect 602 623 603 627
rect 607 626 608 627
rect 683 627 689 628
rect 683 626 684 627
rect 607 624 684 626
rect 607 623 608 624
rect 602 622 608 623
rect 683 623 684 624
rect 688 623 689 627
rect 683 622 689 623
rect 706 627 712 628
rect 706 623 707 627
rect 711 626 712 627
rect 795 627 801 628
rect 795 626 796 627
rect 711 624 796 626
rect 711 623 712 624
rect 706 622 712 623
rect 795 623 796 624
rect 800 623 801 627
rect 795 622 801 623
rect 907 627 913 628
rect 907 623 908 627
rect 912 626 913 627
rect 959 627 965 628
rect 959 626 960 627
rect 912 624 960 626
rect 912 623 913 624
rect 907 622 913 623
rect 959 623 960 624
rect 964 623 965 627
rect 1123 627 1129 628
rect 959 622 965 623
rect 967 623 973 624
rect 967 619 968 623
rect 972 622 973 623
rect 1019 623 1025 624
rect 1019 622 1020 623
rect 972 620 1020 622
rect 972 619 973 620
rect 967 618 973 619
rect 1019 619 1020 620
rect 1024 619 1025 623
rect 1123 623 1124 627
rect 1128 626 1129 627
rect 1159 627 1165 628
rect 1159 626 1160 627
rect 1128 624 1160 626
rect 1128 623 1129 624
rect 1123 622 1129 623
rect 1159 623 1160 624
rect 1164 623 1165 627
rect 1159 622 1165 623
rect 1234 627 1241 628
rect 1234 623 1235 627
rect 1240 623 1241 627
rect 1234 622 1241 623
rect 1347 627 1353 628
rect 1347 623 1348 627
rect 1352 626 1353 627
rect 1382 627 1388 628
rect 1382 626 1383 627
rect 1352 624 1383 626
rect 1352 623 1353 624
rect 1347 622 1353 623
rect 1382 623 1383 624
rect 1387 623 1388 627
rect 1382 622 1388 623
rect 1459 627 1465 628
rect 1459 623 1460 627
rect 1464 626 1465 627
rect 1490 627 1496 628
rect 2046 627 2052 628
rect 2110 631 2116 632
rect 2110 627 2111 631
rect 2115 627 2116 631
rect 1490 626 1491 627
rect 1464 624 1491 626
rect 1464 623 1465 624
rect 1459 622 1465 623
rect 1490 623 1491 624
rect 1495 623 1496 627
rect 2110 626 2116 627
rect 2246 631 2252 632
rect 2246 627 2247 631
rect 2251 627 2252 631
rect 2246 626 2252 627
rect 2398 631 2404 632
rect 2398 627 2399 631
rect 2403 627 2404 631
rect 2398 626 2404 627
rect 2574 631 2580 632
rect 2574 627 2575 631
rect 2579 627 2580 631
rect 2574 626 2580 627
rect 2758 631 2764 632
rect 2758 627 2759 631
rect 2763 627 2764 631
rect 2758 626 2764 627
rect 2942 631 2948 632
rect 2942 627 2943 631
rect 2947 627 2948 631
rect 2942 626 2948 627
rect 3126 631 3132 632
rect 3126 627 3127 631
rect 3131 627 3132 631
rect 3126 626 3132 627
rect 3302 631 3308 632
rect 3302 627 3303 631
rect 3307 627 3308 631
rect 3302 626 3308 627
rect 3478 631 3484 632
rect 3478 627 3479 631
rect 3483 627 3484 631
rect 3478 626 3484 627
rect 3654 631 3660 632
rect 3654 627 3655 631
rect 3659 627 3660 631
rect 3654 626 3660 627
rect 3830 631 3836 632
rect 3830 627 3831 631
rect 3835 627 3836 631
rect 3942 628 3943 632
rect 3947 628 3948 632
rect 3830 626 3836 627
rect 3898 627 3904 628
rect 3942 627 3948 628
rect 1490 622 1496 623
rect 1530 623 1536 624
rect 1019 618 1025 619
rect 1530 619 1531 623
rect 1535 622 1536 623
rect 1571 623 1577 624
rect 1571 622 1572 623
rect 1535 620 1572 622
rect 1535 619 1536 620
rect 1530 618 1536 619
rect 1571 619 1572 620
rect 1576 619 1577 623
rect 1571 618 1577 619
rect 2103 623 2109 624
rect 2103 619 2104 623
rect 2108 622 2109 623
rect 2194 623 2200 624
rect 2108 620 2153 622
rect 2108 619 2109 620
rect 2103 618 2109 619
rect 2194 619 2195 623
rect 2199 622 2200 623
rect 2359 623 2365 624
rect 2199 620 2289 622
rect 2199 619 2200 620
rect 2194 618 2200 619
rect 2359 619 2360 623
rect 2364 622 2365 623
rect 2658 623 2664 624
rect 2364 620 2441 622
rect 2364 619 2365 620
rect 2359 618 2365 619
rect 2650 619 2656 620
rect 2046 615 2052 616
rect 762 611 768 612
rect 739 609 745 610
rect 739 605 740 609
rect 744 605 745 609
rect 762 607 763 611
rect 767 610 768 611
rect 835 611 841 612
rect 835 610 836 611
rect 767 608 836 610
rect 767 607 768 608
rect 762 606 768 607
rect 835 607 836 608
rect 840 607 841 611
rect 835 606 841 607
rect 871 611 877 612
rect 871 607 872 611
rect 876 610 877 611
rect 931 611 937 612
rect 931 610 932 611
rect 876 608 932 610
rect 876 607 877 608
rect 871 606 877 607
rect 931 607 932 608
rect 936 607 937 611
rect 931 606 937 607
rect 1027 611 1033 612
rect 1027 607 1028 611
rect 1032 610 1033 611
rect 1058 611 1064 612
rect 1058 610 1059 611
rect 1032 608 1059 610
rect 1032 607 1033 608
rect 1027 606 1033 607
rect 1058 607 1059 608
rect 1063 607 1064 611
rect 1146 611 1152 612
rect 1058 606 1064 607
rect 1123 609 1129 610
rect 739 604 745 605
rect 1123 605 1124 609
rect 1128 605 1129 609
rect 1146 607 1147 611
rect 1151 610 1152 611
rect 1219 611 1225 612
rect 1219 610 1220 611
rect 1151 608 1220 610
rect 1151 607 1152 608
rect 1146 606 1152 607
rect 1219 607 1220 608
rect 1224 607 1225 611
rect 1219 606 1225 607
rect 1242 611 1248 612
rect 1242 607 1243 611
rect 1247 610 1248 611
rect 1315 611 1321 612
rect 1315 610 1316 611
rect 1247 608 1316 610
rect 1247 607 1248 608
rect 1242 606 1248 607
rect 1315 607 1316 608
rect 1320 607 1321 611
rect 1315 606 1321 607
rect 1338 611 1344 612
rect 1338 607 1339 611
rect 1343 610 1344 611
rect 1411 611 1417 612
rect 1411 610 1412 611
rect 1343 608 1412 610
rect 1343 607 1344 608
rect 1338 606 1344 607
rect 1411 607 1412 608
rect 1416 607 1417 611
rect 1411 606 1417 607
rect 1434 611 1440 612
rect 1434 607 1435 611
rect 1439 610 1440 611
rect 1507 611 1513 612
rect 1507 610 1508 611
rect 1439 608 1508 610
rect 1439 607 1440 608
rect 1434 606 1440 607
rect 1507 607 1508 608
rect 1512 607 1513 611
rect 2046 611 2047 615
rect 2051 611 2052 615
rect 2650 615 2651 619
rect 2655 615 2656 619
rect 2658 619 2659 623
rect 2663 622 2664 623
rect 3118 623 3124 624
rect 2663 620 2801 622
rect 2663 619 2664 620
rect 2658 618 2664 619
rect 3018 619 3024 620
rect 2650 614 2656 615
rect 3018 615 3019 619
rect 3023 615 3024 619
rect 3118 619 3119 623
rect 3123 622 3124 623
rect 3390 623 3396 624
rect 3123 620 3169 622
rect 3123 619 3124 620
rect 3118 618 3124 619
rect 3378 619 3384 620
rect 3018 614 3024 615
rect 3378 615 3379 619
rect 3383 615 3384 619
rect 3390 619 3391 623
rect 3395 622 3396 623
rect 3598 623 3604 624
rect 3395 620 3521 622
rect 3395 619 3396 620
rect 3390 618 3396 619
rect 3598 619 3599 623
rect 3603 622 3604 623
rect 3898 623 3899 627
rect 3903 626 3904 627
rect 3903 624 3910 626
rect 3903 623 3904 624
rect 3898 622 3904 623
rect 3603 620 3697 622
rect 3908 621 3910 624
rect 3603 619 3604 620
rect 3598 618 3604 619
rect 3378 614 3384 615
rect 3942 615 3948 616
rect 2046 610 2052 611
rect 2110 612 2116 613
rect 2110 608 2111 612
rect 2115 608 2116 612
rect 2110 607 2116 608
rect 2246 612 2252 613
rect 2246 608 2247 612
rect 2251 608 2252 612
rect 2246 607 2252 608
rect 2398 612 2404 613
rect 2398 608 2399 612
rect 2403 608 2404 612
rect 2398 607 2404 608
rect 2574 612 2580 613
rect 2574 608 2575 612
rect 2579 608 2580 612
rect 2574 607 2580 608
rect 2758 612 2764 613
rect 2758 608 2759 612
rect 2763 608 2764 612
rect 2758 607 2764 608
rect 2942 612 2948 613
rect 2942 608 2943 612
rect 2947 608 2948 612
rect 2942 607 2948 608
rect 3126 612 3132 613
rect 3126 608 3127 612
rect 3131 608 3132 612
rect 3126 607 3132 608
rect 3302 612 3308 613
rect 3302 608 3303 612
rect 3307 608 3308 612
rect 3302 607 3308 608
rect 3478 612 3484 613
rect 3478 608 3479 612
rect 3483 608 3484 612
rect 3478 607 3484 608
rect 3654 612 3660 613
rect 3654 608 3655 612
rect 3659 608 3660 612
rect 3654 607 3660 608
rect 3830 612 3836 613
rect 3830 608 3831 612
rect 3835 608 3836 612
rect 3942 611 3943 615
rect 3947 611 3948 615
rect 3942 610 3948 611
rect 3830 607 3836 608
rect 1507 606 1513 607
rect 1123 604 1129 605
rect 740 602 742 604
rect 1042 603 1048 604
rect 1042 602 1043 603
rect 740 600 1043 602
rect 1042 599 1043 600
rect 1047 599 1048 603
rect 1124 602 1126 604
rect 1330 603 1336 604
rect 1330 602 1331 603
rect 1124 600 1331 602
rect 1042 598 1048 599
rect 1330 599 1331 600
rect 1335 599 1336 603
rect 1330 598 1336 599
rect 2658 599 2664 600
rect 2658 598 2659 599
rect 2476 596 2659 598
rect 2163 591 2169 592
rect 686 588 692 589
rect 110 585 116 586
rect 110 581 111 585
rect 115 581 116 585
rect 686 584 687 588
rect 691 584 692 588
rect 686 583 692 584
rect 782 588 788 589
rect 782 584 783 588
rect 787 584 788 588
rect 782 583 788 584
rect 878 588 884 589
rect 878 584 879 588
rect 883 584 884 588
rect 878 583 884 584
rect 974 588 980 589
rect 974 584 975 588
rect 979 584 980 588
rect 974 583 980 584
rect 1070 588 1076 589
rect 1070 584 1071 588
rect 1075 584 1076 588
rect 1070 583 1076 584
rect 1166 588 1172 589
rect 1166 584 1167 588
rect 1171 584 1172 588
rect 1166 583 1172 584
rect 1262 588 1268 589
rect 1262 584 1263 588
rect 1267 584 1268 588
rect 1262 583 1268 584
rect 1358 588 1364 589
rect 1358 584 1359 588
rect 1363 584 1364 588
rect 1358 583 1364 584
rect 1454 588 1460 589
rect 1454 584 1455 588
rect 1459 584 1460 588
rect 2163 587 2164 591
rect 2168 590 2169 591
rect 2194 591 2200 592
rect 2194 590 2195 591
rect 2168 588 2195 590
rect 2168 587 2169 588
rect 2163 586 2169 587
rect 2194 587 2195 588
rect 2199 587 2200 591
rect 2194 586 2200 587
rect 2299 591 2305 592
rect 2299 587 2300 591
rect 2304 590 2305 591
rect 2359 591 2365 592
rect 2359 590 2360 591
rect 2304 588 2360 590
rect 2304 587 2305 588
rect 2299 586 2305 587
rect 2359 587 2360 588
rect 2364 587 2365 591
rect 2359 586 2365 587
rect 2451 591 2457 592
rect 2451 587 2452 591
rect 2456 590 2457 591
rect 2476 590 2478 596
rect 2658 595 2659 596
rect 2663 595 2664 599
rect 2658 594 2664 595
rect 2456 588 2478 590
rect 2582 591 2588 592
rect 2456 587 2457 588
rect 2451 586 2457 587
rect 2582 587 2583 591
rect 2587 590 2588 591
rect 2627 591 2633 592
rect 2627 590 2628 591
rect 2587 588 2628 590
rect 2587 587 2588 588
rect 2582 586 2588 587
rect 2627 587 2628 588
rect 2632 587 2633 591
rect 2627 586 2633 587
rect 2650 591 2656 592
rect 2650 587 2651 591
rect 2655 590 2656 591
rect 2811 591 2817 592
rect 2811 590 2812 591
rect 2655 588 2812 590
rect 2655 587 2656 588
rect 2650 586 2656 587
rect 2811 587 2812 588
rect 2816 587 2817 591
rect 3018 591 3024 592
rect 2811 586 2817 587
rect 2954 587 2960 588
rect 1454 583 1460 584
rect 2006 585 2012 586
rect 110 580 116 581
rect 2006 581 2007 585
rect 2011 581 2012 585
rect 2954 583 2955 587
rect 2959 586 2960 587
rect 2995 587 3001 588
rect 2995 586 2996 587
rect 2959 584 2996 586
rect 2959 583 2960 584
rect 2954 582 2960 583
rect 2995 583 2996 584
rect 3000 583 3001 587
rect 3018 587 3019 591
rect 3023 590 3024 591
rect 3179 591 3185 592
rect 3179 590 3180 591
rect 3023 588 3180 590
rect 3023 587 3024 588
rect 3018 586 3024 587
rect 3179 587 3180 588
rect 3184 587 3185 591
rect 3179 586 3185 587
rect 3355 591 3361 592
rect 3355 587 3356 591
rect 3360 590 3361 591
rect 3390 591 3396 592
rect 3390 590 3391 591
rect 3360 588 3391 590
rect 3360 587 3361 588
rect 3355 586 3361 587
rect 3390 587 3391 588
rect 3395 587 3396 591
rect 3390 586 3396 587
rect 3531 591 3537 592
rect 3531 587 3532 591
rect 3536 590 3537 591
rect 3598 591 3604 592
rect 3598 590 3599 591
rect 3536 588 3599 590
rect 3536 587 3537 588
rect 3531 586 3537 587
rect 3598 587 3599 588
rect 3603 587 3604 591
rect 3598 586 3604 587
rect 3707 591 3713 592
rect 3707 587 3708 591
rect 3712 590 3713 591
rect 3746 591 3752 592
rect 3746 590 3747 591
rect 3712 588 3747 590
rect 3712 587 3713 588
rect 3707 586 3713 587
rect 3746 587 3747 588
rect 3751 587 3752 591
rect 3746 586 3752 587
rect 3883 587 3889 588
rect 2995 582 3001 583
rect 3883 583 3884 587
rect 3888 586 3889 587
rect 3906 587 3912 588
rect 3906 586 3907 587
rect 3888 584 3907 586
rect 3888 583 3889 584
rect 3883 582 3889 583
rect 3906 583 3907 584
rect 3911 583 3912 587
rect 3906 582 3912 583
rect 2006 580 2012 581
rect 762 579 768 580
rect 762 575 763 579
rect 767 575 768 579
rect 871 579 877 580
rect 871 578 872 579
rect 861 576 872 578
rect 762 574 768 575
rect 871 575 872 576
rect 876 575 877 579
rect 967 579 973 580
rect 967 578 968 579
rect 957 576 968 578
rect 871 574 877 575
rect 967 575 968 576
rect 972 575 973 579
rect 967 574 973 575
rect 1042 579 1048 580
rect 1042 575 1043 579
rect 1047 575 1048 579
rect 1042 574 1048 575
rect 1058 579 1064 580
rect 1058 575 1059 579
rect 1063 578 1064 579
rect 1242 579 1248 580
rect 1063 576 1113 578
rect 1063 575 1064 576
rect 1058 574 1064 575
rect 1242 575 1243 579
rect 1247 575 1248 579
rect 1242 574 1248 575
rect 1338 579 1344 580
rect 1338 575 1339 579
rect 1343 575 1344 579
rect 1338 574 1344 575
rect 1434 579 1440 580
rect 1434 575 1435 579
rect 1439 575 1440 579
rect 1434 574 1440 575
rect 1530 579 1536 580
rect 1530 575 1531 579
rect 1535 575 1536 579
rect 1530 574 1536 575
rect 2103 571 2109 572
rect 686 569 692 570
rect 110 568 116 569
rect 110 564 111 568
rect 115 564 116 568
rect 686 565 687 569
rect 691 565 692 569
rect 686 564 692 565
rect 782 569 788 570
rect 782 565 783 569
rect 787 565 788 569
rect 782 564 788 565
rect 878 569 884 570
rect 878 565 879 569
rect 883 565 884 569
rect 878 564 884 565
rect 974 569 980 570
rect 974 565 975 569
rect 979 565 980 569
rect 974 564 980 565
rect 1070 569 1076 570
rect 1070 565 1071 569
rect 1075 565 1076 569
rect 1070 564 1076 565
rect 1166 569 1172 570
rect 1166 565 1167 569
rect 1171 565 1172 569
rect 1166 564 1172 565
rect 1262 569 1268 570
rect 1262 565 1263 569
rect 1267 565 1268 569
rect 1262 564 1268 565
rect 1358 569 1364 570
rect 1358 565 1359 569
rect 1363 565 1364 569
rect 1358 564 1364 565
rect 1454 569 1460 570
rect 1454 565 1455 569
rect 1459 565 1460 569
rect 1454 564 1460 565
rect 2006 568 2012 569
rect 2006 564 2007 568
rect 2011 564 2012 568
rect 2103 567 2104 571
rect 2108 570 2109 571
rect 2123 571 2129 572
rect 2123 570 2124 571
rect 2108 568 2124 570
rect 2108 567 2109 568
rect 2103 566 2109 567
rect 2123 567 2124 568
rect 2128 567 2129 571
rect 2123 566 2129 567
rect 2146 571 2152 572
rect 2146 567 2147 571
rect 2151 570 2152 571
rect 2235 571 2241 572
rect 2235 570 2236 571
rect 2151 568 2236 570
rect 2151 567 2152 568
rect 2146 566 2152 567
rect 2235 567 2236 568
rect 2240 567 2241 571
rect 2235 566 2241 567
rect 2258 571 2264 572
rect 2258 567 2259 571
rect 2263 570 2264 571
rect 2387 571 2393 572
rect 2387 570 2388 571
rect 2263 568 2388 570
rect 2263 567 2264 568
rect 2258 566 2264 567
rect 2387 567 2388 568
rect 2392 567 2393 571
rect 2387 566 2393 567
rect 2410 571 2416 572
rect 2410 567 2411 571
rect 2415 570 2416 571
rect 2555 571 2561 572
rect 2555 570 2556 571
rect 2415 568 2556 570
rect 2415 567 2416 568
rect 2410 566 2416 567
rect 2555 567 2556 568
rect 2560 567 2561 571
rect 2555 566 2561 567
rect 2639 571 2645 572
rect 2639 567 2640 571
rect 2644 570 2645 571
rect 2739 571 2745 572
rect 2739 570 2740 571
rect 2644 568 2740 570
rect 2644 567 2645 568
rect 2639 566 2645 567
rect 2739 567 2740 568
rect 2744 567 2745 571
rect 2739 566 2745 567
rect 2931 571 2937 572
rect 2931 567 2932 571
rect 2936 570 2937 571
rect 2962 571 2968 572
rect 2962 570 2963 571
rect 2936 568 2963 570
rect 2936 567 2937 568
rect 2931 566 2937 567
rect 2962 567 2963 568
rect 2967 567 2968 571
rect 2962 566 2968 567
rect 3123 571 3129 572
rect 3123 567 3124 571
rect 3128 570 3129 571
rect 3174 571 3180 572
rect 3174 570 3175 571
rect 3128 568 3175 570
rect 3128 567 3129 568
rect 3123 566 3129 567
rect 3174 567 3175 568
rect 3179 567 3180 571
rect 3174 566 3180 567
rect 3234 571 3240 572
rect 3234 567 3235 571
rect 3239 570 3240 571
rect 3315 571 3321 572
rect 3315 570 3316 571
rect 3239 568 3316 570
rect 3239 567 3240 568
rect 3234 566 3240 567
rect 3315 567 3316 568
rect 3320 567 3321 571
rect 3315 566 3321 567
rect 3378 571 3384 572
rect 3378 567 3379 571
rect 3383 570 3384 571
rect 3507 571 3513 572
rect 3507 570 3508 571
rect 3383 568 3508 570
rect 3383 567 3384 568
rect 3378 566 3384 567
rect 3507 567 3508 568
rect 3512 567 3513 571
rect 3507 566 3513 567
rect 3530 571 3536 572
rect 3530 567 3531 571
rect 3535 570 3536 571
rect 3699 571 3705 572
rect 3699 570 3700 571
rect 3535 568 3700 570
rect 3535 567 3536 568
rect 3530 566 3536 567
rect 3699 567 3700 568
rect 3704 567 3705 571
rect 3699 566 3705 567
rect 3722 571 3728 572
rect 3722 567 3723 571
rect 3727 570 3728 571
rect 3891 571 3897 572
rect 3891 570 3892 571
rect 3727 568 3892 570
rect 3727 567 3728 568
rect 3722 566 3728 567
rect 3891 567 3892 568
rect 3896 567 3897 571
rect 3891 566 3897 567
rect 110 563 116 564
rect 2006 563 2012 564
rect 2070 548 2076 549
rect 2046 545 2052 546
rect 2046 541 2047 545
rect 2051 541 2052 545
rect 2070 544 2071 548
rect 2075 544 2076 548
rect 2070 543 2076 544
rect 2182 548 2188 549
rect 2182 544 2183 548
rect 2187 544 2188 548
rect 2182 543 2188 544
rect 2334 548 2340 549
rect 2334 544 2335 548
rect 2339 544 2340 548
rect 2334 543 2340 544
rect 2502 548 2508 549
rect 2502 544 2503 548
rect 2507 544 2508 548
rect 2502 543 2508 544
rect 2686 548 2692 549
rect 2686 544 2687 548
rect 2691 544 2692 548
rect 2686 543 2692 544
rect 2878 548 2884 549
rect 2878 544 2879 548
rect 2883 544 2884 548
rect 2878 543 2884 544
rect 3070 548 3076 549
rect 3070 544 3071 548
rect 3075 544 3076 548
rect 3070 543 3076 544
rect 3262 548 3268 549
rect 3262 544 3263 548
rect 3267 544 3268 548
rect 3262 543 3268 544
rect 3454 548 3460 549
rect 3454 544 3455 548
rect 3459 544 3460 548
rect 3454 543 3460 544
rect 3646 548 3652 549
rect 3646 544 3647 548
rect 3651 544 3652 548
rect 3646 543 3652 544
rect 3838 548 3844 549
rect 3838 544 3839 548
rect 3843 544 3844 548
rect 3838 543 3844 544
rect 3942 545 3948 546
rect 2046 540 2052 541
rect 3942 541 3943 545
rect 3947 541 3948 545
rect 3942 540 3948 541
rect 2146 539 2152 540
rect 2146 535 2147 539
rect 2151 535 2152 539
rect 2146 534 2152 535
rect 2258 539 2264 540
rect 2258 535 2259 539
rect 2263 535 2264 539
rect 2258 534 2264 535
rect 2410 539 2416 540
rect 2410 535 2411 539
rect 2415 535 2416 539
rect 2639 539 2645 540
rect 2639 538 2640 539
rect 2581 536 2640 538
rect 2410 534 2416 535
rect 2639 535 2640 536
rect 2644 535 2645 539
rect 2639 534 2645 535
rect 2658 539 2664 540
rect 2658 535 2659 539
rect 2663 538 2664 539
rect 2954 539 2960 540
rect 2663 536 2729 538
rect 2663 535 2664 536
rect 2658 534 2664 535
rect 2954 535 2955 539
rect 2959 535 2960 539
rect 2954 534 2960 535
rect 2962 539 2968 540
rect 2962 535 2963 539
rect 2967 538 2968 539
rect 3174 539 3180 540
rect 2967 536 3113 538
rect 2967 535 2968 536
rect 2962 534 2968 535
rect 3174 535 3175 539
rect 3179 538 3180 539
rect 3530 539 3536 540
rect 3179 536 3305 538
rect 3179 535 3180 536
rect 3174 534 3180 535
rect 3530 535 3531 539
rect 3535 535 3536 539
rect 3530 534 3536 535
rect 3722 539 3728 540
rect 3722 535 3723 539
rect 3727 535 3728 539
rect 3722 534 3728 535
rect 3906 539 3912 540
rect 3906 535 3907 539
rect 3911 535 3912 539
rect 3906 534 3912 535
rect 2070 529 2076 530
rect 2046 528 2052 529
rect 2046 524 2047 528
rect 2051 524 2052 528
rect 2070 525 2071 529
rect 2075 525 2076 529
rect 2070 524 2076 525
rect 2182 529 2188 530
rect 2182 525 2183 529
rect 2187 525 2188 529
rect 2182 524 2188 525
rect 2334 529 2340 530
rect 2334 525 2335 529
rect 2339 525 2340 529
rect 2334 524 2340 525
rect 2502 529 2508 530
rect 2502 525 2503 529
rect 2507 525 2508 529
rect 2502 524 2508 525
rect 2686 529 2692 530
rect 2686 525 2687 529
rect 2691 525 2692 529
rect 2686 524 2692 525
rect 2878 529 2884 530
rect 2878 525 2879 529
rect 2883 525 2884 529
rect 2878 524 2884 525
rect 3070 529 3076 530
rect 3070 525 3071 529
rect 3075 525 3076 529
rect 3070 524 3076 525
rect 3262 529 3268 530
rect 3262 525 3263 529
rect 3267 525 3268 529
rect 3262 524 3268 525
rect 3454 529 3460 530
rect 3454 525 3455 529
rect 3459 525 3460 529
rect 3454 524 3460 525
rect 3646 529 3652 530
rect 3646 525 3647 529
rect 3651 525 3652 529
rect 3646 524 3652 525
rect 3838 529 3844 530
rect 3838 525 3839 529
rect 3843 525 3844 529
rect 3838 524 3844 525
rect 3942 528 3948 529
rect 3942 524 3943 528
rect 3947 524 3948 528
rect 2046 523 2052 524
rect 3942 523 3948 524
rect 110 496 116 497
rect 2006 496 2012 497
rect 110 492 111 496
rect 115 492 116 496
rect 110 491 116 492
rect 382 495 388 496
rect 382 491 383 495
rect 387 491 388 495
rect 382 490 388 491
rect 478 495 484 496
rect 478 491 479 495
rect 483 491 484 495
rect 478 490 484 491
rect 574 495 580 496
rect 574 491 575 495
rect 579 491 580 495
rect 574 490 580 491
rect 670 495 676 496
rect 670 491 671 495
rect 675 491 676 495
rect 670 490 676 491
rect 766 495 772 496
rect 766 491 767 495
rect 771 491 772 495
rect 766 490 772 491
rect 862 495 868 496
rect 862 491 863 495
rect 867 491 868 495
rect 862 490 868 491
rect 958 495 964 496
rect 958 491 959 495
rect 963 491 964 495
rect 958 490 964 491
rect 1054 495 1060 496
rect 1054 491 1055 495
rect 1059 491 1060 495
rect 1054 490 1060 491
rect 1150 495 1156 496
rect 1150 491 1151 495
rect 1155 491 1156 495
rect 1150 490 1156 491
rect 1246 495 1252 496
rect 1246 491 1247 495
rect 1251 491 1252 495
rect 1246 490 1252 491
rect 1342 495 1348 496
rect 1342 491 1343 495
rect 1347 491 1348 495
rect 1342 490 1348 491
rect 1438 495 1444 496
rect 1438 491 1439 495
rect 1443 491 1444 495
rect 1438 490 1444 491
rect 1534 495 1540 496
rect 1534 491 1535 495
rect 1539 491 1540 495
rect 2006 492 2007 496
rect 2011 492 2012 496
rect 2006 491 2012 492
rect 1534 490 1540 491
rect 1239 487 1245 488
rect 458 483 464 484
rect 110 479 116 480
rect 110 475 111 479
rect 115 475 116 479
rect 458 479 459 483
rect 463 479 464 483
rect 458 478 464 479
rect 554 483 560 484
rect 554 479 555 483
rect 559 479 560 483
rect 554 478 560 479
rect 650 483 656 484
rect 650 479 651 483
rect 655 479 656 483
rect 650 478 656 479
rect 746 483 752 484
rect 746 479 747 483
rect 751 479 752 483
rect 746 478 752 479
rect 842 483 848 484
rect 842 479 843 483
rect 847 479 848 483
rect 842 478 848 479
rect 938 483 944 484
rect 938 479 939 483
rect 943 479 944 483
rect 938 478 944 479
rect 1034 483 1040 484
rect 1034 479 1035 483
rect 1039 479 1040 483
rect 1034 478 1040 479
rect 1130 483 1136 484
rect 1130 479 1131 483
rect 1135 479 1136 483
rect 1130 478 1136 479
rect 1226 483 1232 484
rect 1226 479 1227 483
rect 1231 479 1232 483
rect 1239 483 1240 487
rect 1244 486 1245 487
rect 1330 487 1336 488
rect 1244 484 1289 486
rect 1244 483 1245 484
rect 1239 482 1245 483
rect 1330 483 1331 487
rect 1335 486 1336 487
rect 1527 487 1533 488
rect 1335 484 1385 486
rect 1335 483 1336 484
rect 1330 482 1336 483
rect 1514 483 1520 484
rect 1226 478 1232 479
rect 1514 479 1515 483
rect 1519 479 1520 483
rect 1527 483 1528 487
rect 1532 486 1533 487
rect 1532 484 1577 486
rect 1532 483 1533 484
rect 1527 482 1533 483
rect 1514 478 1520 479
rect 2006 479 2012 480
rect 110 474 116 475
rect 382 476 388 477
rect 382 472 383 476
rect 387 472 388 476
rect 382 471 388 472
rect 478 476 484 477
rect 478 472 479 476
rect 483 472 484 476
rect 478 471 484 472
rect 574 476 580 477
rect 574 472 575 476
rect 579 472 580 476
rect 574 471 580 472
rect 670 476 676 477
rect 670 472 671 476
rect 675 472 676 476
rect 670 471 676 472
rect 766 476 772 477
rect 766 472 767 476
rect 771 472 772 476
rect 766 471 772 472
rect 862 476 868 477
rect 862 472 863 476
rect 867 472 868 476
rect 862 471 868 472
rect 958 476 964 477
rect 958 472 959 476
rect 963 472 964 476
rect 958 471 964 472
rect 1054 476 1060 477
rect 1054 472 1055 476
rect 1059 472 1060 476
rect 1054 471 1060 472
rect 1150 476 1156 477
rect 1150 472 1151 476
rect 1155 472 1156 476
rect 1150 471 1156 472
rect 1246 476 1252 477
rect 1246 472 1247 476
rect 1251 472 1252 476
rect 1246 471 1252 472
rect 1342 476 1348 477
rect 1342 472 1343 476
rect 1347 472 1348 476
rect 1342 471 1348 472
rect 1438 476 1444 477
rect 1438 472 1439 476
rect 1443 472 1444 476
rect 1438 471 1444 472
rect 1534 476 1540 477
rect 1534 472 1535 476
rect 1539 472 1540 476
rect 2006 475 2007 479
rect 2011 475 2012 479
rect 2006 474 2012 475
rect 2046 476 2052 477
rect 3942 476 3948 477
rect 1534 471 1540 472
rect 2046 472 2047 476
rect 2051 472 2052 476
rect 2046 471 2052 472
rect 2182 475 2188 476
rect 2182 471 2183 475
rect 2187 471 2188 475
rect 2182 470 2188 471
rect 2318 475 2324 476
rect 2318 471 2319 475
rect 2323 471 2324 475
rect 2318 470 2324 471
rect 2462 475 2468 476
rect 2462 471 2463 475
rect 2467 471 2468 475
rect 2462 470 2468 471
rect 2614 475 2620 476
rect 2614 471 2615 475
rect 2619 471 2620 475
rect 2614 470 2620 471
rect 2774 475 2780 476
rect 2774 471 2775 475
rect 2779 471 2780 475
rect 2774 470 2780 471
rect 2958 475 2964 476
rect 2958 471 2959 475
rect 2963 471 2964 475
rect 2958 470 2964 471
rect 3158 475 3164 476
rect 3158 471 3159 475
rect 3163 471 3164 475
rect 3158 470 3164 471
rect 3366 475 3372 476
rect 3366 471 3367 475
rect 3371 471 3372 475
rect 3366 470 3372 471
rect 3582 475 3588 476
rect 3582 471 3583 475
rect 3587 471 3588 475
rect 3582 470 3588 471
rect 3806 475 3812 476
rect 3806 471 3807 475
rect 3811 471 3812 475
rect 3942 472 3943 476
rect 3947 472 3948 476
rect 3942 471 3948 472
rect 3806 470 3812 471
rect 2698 467 2704 468
rect 1527 463 1533 464
rect 1527 462 1528 463
rect 1460 460 1528 462
rect 458 455 464 456
rect 435 451 441 452
rect 435 447 436 451
rect 440 450 441 451
rect 458 451 459 455
rect 463 454 464 455
rect 531 455 537 456
rect 531 454 532 455
rect 463 452 532 454
rect 463 451 464 452
rect 458 450 464 451
rect 531 451 532 452
rect 536 451 537 455
rect 531 450 537 451
rect 554 455 560 456
rect 554 451 555 455
rect 559 454 560 455
rect 627 455 633 456
rect 627 454 628 455
rect 559 452 628 454
rect 559 451 560 452
rect 554 450 560 451
rect 627 451 628 452
rect 632 451 633 455
rect 627 450 633 451
rect 650 455 656 456
rect 650 451 651 455
rect 655 454 656 455
rect 723 455 729 456
rect 723 454 724 455
rect 655 452 724 454
rect 655 451 656 452
rect 650 450 656 451
rect 723 451 724 452
rect 728 451 729 455
rect 723 450 729 451
rect 746 455 752 456
rect 746 451 747 455
rect 751 454 752 455
rect 819 455 825 456
rect 819 454 820 455
rect 751 452 820 454
rect 751 451 752 452
rect 746 450 752 451
rect 819 451 820 452
rect 824 451 825 455
rect 819 450 825 451
rect 842 455 848 456
rect 842 451 843 455
rect 847 454 848 455
rect 915 455 921 456
rect 915 454 916 455
rect 847 452 916 454
rect 847 451 848 452
rect 842 450 848 451
rect 915 451 916 452
rect 920 451 921 455
rect 915 450 921 451
rect 938 455 944 456
rect 938 451 939 455
rect 943 454 944 455
rect 1011 455 1017 456
rect 1011 454 1012 455
rect 943 452 1012 454
rect 943 451 944 452
rect 938 450 944 451
rect 1011 451 1012 452
rect 1016 451 1017 455
rect 1011 450 1017 451
rect 1034 455 1040 456
rect 1034 451 1035 455
rect 1039 454 1040 455
rect 1107 455 1113 456
rect 1107 454 1108 455
rect 1039 452 1108 454
rect 1039 451 1040 452
rect 1034 450 1040 451
rect 1107 451 1108 452
rect 1112 451 1113 455
rect 1107 450 1113 451
rect 1130 455 1136 456
rect 1130 451 1131 455
rect 1135 454 1136 455
rect 1203 455 1209 456
rect 1203 454 1204 455
rect 1135 452 1204 454
rect 1135 451 1136 452
rect 1130 450 1136 451
rect 1203 451 1204 452
rect 1208 451 1209 455
rect 1203 450 1209 451
rect 1226 455 1232 456
rect 1226 451 1227 455
rect 1231 454 1232 455
rect 1299 455 1305 456
rect 1299 454 1300 455
rect 1231 452 1300 454
rect 1231 451 1232 452
rect 1226 450 1232 451
rect 1299 451 1300 452
rect 1304 451 1305 455
rect 1299 450 1305 451
rect 1395 455 1401 456
rect 1395 451 1396 455
rect 1400 454 1401 455
rect 1460 454 1462 460
rect 1527 459 1528 460
rect 1532 459 1533 463
rect 2258 463 2264 464
rect 1527 458 1533 459
rect 2046 459 2052 460
rect 1400 452 1462 454
rect 1514 455 1520 456
rect 1400 451 1401 452
rect 1395 450 1401 451
rect 1491 451 1500 452
rect 440 448 454 450
rect 440 447 441 448
rect 435 446 441 447
rect 452 446 454 448
rect 966 447 972 448
rect 966 446 967 447
rect 452 444 967 446
rect 966 443 967 444
rect 971 443 972 447
rect 1491 447 1492 451
rect 1499 447 1500 451
rect 1514 451 1515 455
rect 1519 454 1520 455
rect 1587 455 1593 456
rect 1587 454 1588 455
rect 1519 452 1588 454
rect 1519 451 1520 452
rect 1514 450 1520 451
rect 1587 451 1588 452
rect 1592 451 1593 455
rect 2046 455 2047 459
rect 2051 455 2052 459
rect 2258 459 2259 463
rect 2263 459 2264 463
rect 2258 458 2264 459
rect 2394 463 2400 464
rect 2394 459 2395 463
rect 2399 459 2400 463
rect 2394 458 2400 459
rect 2538 463 2544 464
rect 2538 459 2539 463
rect 2543 459 2544 463
rect 2538 458 2544 459
rect 2690 463 2696 464
rect 2690 459 2691 463
rect 2695 459 2696 463
rect 2698 463 2699 467
rect 2703 466 2704 467
rect 3234 467 3240 468
rect 2703 464 2817 466
rect 2703 463 2704 464
rect 2698 462 2704 463
rect 3034 463 3040 464
rect 2690 458 2696 459
rect 3034 459 3035 463
rect 3039 459 3040 463
rect 3234 463 3235 467
rect 3239 463 3240 467
rect 3234 462 3240 463
rect 3242 467 3248 468
rect 3242 463 3243 467
rect 3247 466 3248 467
rect 3455 467 3461 468
rect 3247 464 3409 466
rect 3247 463 3248 464
rect 3242 462 3248 463
rect 3455 463 3456 467
rect 3460 466 3461 467
rect 3766 467 3772 468
rect 3460 464 3625 466
rect 3460 463 3461 464
rect 3455 462 3461 463
rect 3766 463 3767 467
rect 3771 466 3772 467
rect 3771 464 3849 466
rect 3771 463 3772 464
rect 3766 462 3772 463
rect 3034 458 3040 459
rect 3942 459 3948 460
rect 2046 454 2052 455
rect 2182 456 2188 457
rect 2182 452 2183 456
rect 2187 452 2188 456
rect 2182 451 2188 452
rect 2318 456 2324 457
rect 2318 452 2319 456
rect 2323 452 2324 456
rect 2318 451 2324 452
rect 2462 456 2468 457
rect 2462 452 2463 456
rect 2467 452 2468 456
rect 2462 451 2468 452
rect 2614 456 2620 457
rect 2614 452 2615 456
rect 2619 452 2620 456
rect 2614 451 2620 452
rect 2774 456 2780 457
rect 2774 452 2775 456
rect 2779 452 2780 456
rect 2774 451 2780 452
rect 2958 456 2964 457
rect 2958 452 2959 456
rect 2963 452 2964 456
rect 2958 451 2964 452
rect 3158 456 3164 457
rect 3158 452 3159 456
rect 3163 452 3164 456
rect 3158 451 3164 452
rect 3366 456 3372 457
rect 3366 452 3367 456
rect 3371 452 3372 456
rect 3366 451 3372 452
rect 3582 456 3588 457
rect 3582 452 3583 456
rect 3587 452 3588 456
rect 3582 451 3588 452
rect 3806 456 3812 457
rect 3806 452 3807 456
rect 3811 452 3812 456
rect 3942 455 3943 459
rect 3947 455 3948 459
rect 3942 454 3948 455
rect 3806 451 3812 452
rect 1587 450 1593 451
rect 1491 446 1500 447
rect 966 442 972 443
rect 2658 443 2664 444
rect 2658 442 2659 443
rect 2252 440 2659 442
rect 2235 435 2241 436
rect 2235 431 2236 435
rect 2240 434 2241 435
rect 2252 434 2254 440
rect 2658 439 2659 440
rect 2663 439 2664 443
rect 3242 443 3248 444
rect 3242 442 3243 443
rect 2658 438 2664 439
rect 3028 440 3243 442
rect 2240 432 2254 434
rect 2258 435 2264 436
rect 2240 431 2241 432
rect 2235 430 2241 431
rect 2258 431 2259 435
rect 2263 434 2264 435
rect 2371 435 2377 436
rect 2371 434 2372 435
rect 2263 432 2372 434
rect 2263 431 2264 432
rect 2258 430 2264 431
rect 2371 431 2372 432
rect 2376 431 2377 435
rect 2371 430 2377 431
rect 2394 435 2400 436
rect 2394 431 2395 435
rect 2399 434 2400 435
rect 2515 435 2521 436
rect 2515 434 2516 435
rect 2399 432 2516 434
rect 2399 431 2400 432
rect 2394 430 2400 431
rect 2515 431 2516 432
rect 2520 431 2521 435
rect 2515 430 2521 431
rect 2538 435 2544 436
rect 2538 431 2539 435
rect 2543 434 2544 435
rect 2667 435 2673 436
rect 2667 434 2668 435
rect 2543 432 2668 434
rect 2543 431 2544 432
rect 2538 430 2544 431
rect 2667 431 2668 432
rect 2672 431 2673 435
rect 2667 430 2673 431
rect 2690 435 2696 436
rect 2690 431 2691 435
rect 2695 434 2696 435
rect 2827 435 2833 436
rect 2827 434 2828 435
rect 2695 432 2828 434
rect 2695 431 2696 432
rect 2690 430 2696 431
rect 2827 431 2828 432
rect 2832 431 2833 435
rect 2827 430 2833 431
rect 3011 435 3017 436
rect 3011 431 3012 435
rect 3016 434 3017 435
rect 3028 434 3030 440
rect 3242 439 3243 440
rect 3247 439 3248 443
rect 3242 438 3248 439
rect 3016 432 3030 434
rect 3034 435 3040 436
rect 3016 431 3017 432
rect 3011 430 3017 431
rect 3034 431 3035 435
rect 3039 434 3040 435
rect 3211 435 3217 436
rect 3211 434 3212 435
rect 3039 432 3212 434
rect 3039 431 3040 432
rect 3034 430 3040 431
rect 3211 431 3212 432
rect 3216 431 3217 435
rect 3211 430 3217 431
rect 3419 435 3425 436
rect 3419 431 3420 435
rect 3424 434 3425 435
rect 3455 435 3461 436
rect 3455 434 3456 435
rect 3424 432 3456 434
rect 3424 431 3425 432
rect 3419 430 3425 431
rect 3455 431 3456 432
rect 3460 431 3461 435
rect 3455 430 3461 431
rect 3490 431 3496 432
rect 562 427 568 428
rect 539 425 545 426
rect 539 424 540 425
rect 538 423 540 424
rect 538 419 539 423
rect 544 421 545 425
rect 562 423 563 427
rect 567 426 568 427
rect 635 427 641 428
rect 635 426 636 427
rect 567 424 636 426
rect 567 423 568 424
rect 562 422 568 423
rect 635 423 636 424
rect 640 423 641 427
rect 635 422 641 423
rect 658 427 664 428
rect 658 423 659 427
rect 663 426 664 427
rect 739 427 745 428
rect 739 426 740 427
rect 663 424 740 426
rect 663 423 664 424
rect 658 422 664 423
rect 739 423 740 424
rect 744 423 745 427
rect 739 422 745 423
rect 783 427 789 428
rect 783 423 784 427
rect 788 426 789 427
rect 843 427 849 428
rect 843 426 844 427
rect 788 424 844 426
rect 788 423 789 424
rect 783 422 789 423
rect 843 423 844 424
rect 848 423 849 427
rect 843 422 849 423
rect 887 427 893 428
rect 887 423 888 427
rect 892 426 893 427
rect 947 427 953 428
rect 947 426 948 427
rect 892 424 948 426
rect 892 423 893 424
rect 887 422 893 423
rect 947 423 948 424
rect 952 423 953 427
rect 947 422 953 423
rect 1051 427 1057 428
rect 1051 423 1052 427
rect 1056 426 1057 427
rect 1095 427 1101 428
rect 1095 426 1096 427
rect 1056 424 1096 426
rect 1056 423 1057 424
rect 1051 422 1057 423
rect 1095 423 1096 424
rect 1100 423 1101 427
rect 1095 422 1101 423
rect 1155 427 1161 428
rect 1155 423 1156 427
rect 1160 426 1161 427
rect 1186 427 1192 428
rect 1186 426 1187 427
rect 1160 424 1187 426
rect 1160 423 1161 424
rect 1155 422 1161 423
rect 1186 423 1187 424
rect 1191 423 1192 427
rect 1186 422 1192 423
rect 1239 427 1245 428
rect 1239 423 1240 427
rect 1244 426 1245 427
rect 1259 427 1265 428
rect 1259 426 1260 427
rect 1244 424 1260 426
rect 1244 423 1245 424
rect 1239 422 1245 423
rect 1259 423 1260 424
rect 1264 423 1265 427
rect 1259 422 1265 423
rect 1371 427 1377 428
rect 1371 423 1372 427
rect 1376 426 1377 427
rect 1418 427 1424 428
rect 1418 426 1419 427
rect 1376 424 1419 426
rect 1376 423 1377 424
rect 1371 422 1377 423
rect 1418 423 1419 424
rect 1423 423 1424 427
rect 2698 427 2704 428
rect 2698 426 2699 427
rect 1418 422 1424 423
rect 1483 425 1489 426
rect 543 420 545 421
rect 1483 421 1484 425
rect 1488 421 1489 425
rect 2396 424 2699 426
rect 2396 422 2398 424
rect 2698 423 2699 424
rect 2703 423 2704 427
rect 3490 427 3491 431
rect 3495 430 3496 431
rect 3635 431 3641 432
rect 3635 430 3636 431
rect 3495 428 3636 430
rect 3495 427 3496 428
rect 3490 426 3496 427
rect 3635 427 3636 428
rect 3640 427 3641 431
rect 3635 426 3641 427
rect 3859 431 3865 432
rect 3859 427 3860 431
rect 3864 430 3865 431
rect 3906 431 3912 432
rect 3906 430 3907 431
rect 3864 428 3907 430
rect 3864 427 3865 428
rect 3859 426 3865 427
rect 3906 427 3907 428
rect 3911 427 3912 431
rect 3906 426 3912 427
rect 2698 422 2704 423
rect 1483 420 1489 421
rect 2395 421 2401 422
rect 543 419 544 420
rect 538 418 544 419
rect 1394 419 1400 420
rect 1394 415 1395 419
rect 1399 418 1400 419
rect 1484 418 1486 420
rect 1399 416 1486 418
rect 2395 417 2396 421
rect 2400 417 2401 421
rect 2395 416 2401 417
rect 2418 419 2424 420
rect 1399 415 1400 416
rect 1394 414 1400 415
rect 2418 415 2419 419
rect 2423 418 2424 419
rect 2539 419 2545 420
rect 2539 418 2540 419
rect 2423 416 2540 418
rect 2423 415 2424 416
rect 2418 414 2424 415
rect 2539 415 2540 416
rect 2544 415 2545 419
rect 2539 414 2545 415
rect 2562 419 2568 420
rect 2562 415 2563 419
rect 2567 418 2568 419
rect 2691 419 2697 420
rect 2691 418 2692 419
rect 2567 416 2692 418
rect 2567 415 2568 416
rect 2562 414 2568 415
rect 2691 415 2692 416
rect 2696 415 2697 419
rect 2691 414 2697 415
rect 2714 419 2720 420
rect 2714 415 2715 419
rect 2719 418 2720 419
rect 2851 419 2857 420
rect 2851 418 2852 419
rect 2719 416 2852 418
rect 2719 415 2720 416
rect 2714 414 2720 415
rect 2851 415 2852 416
rect 2856 415 2857 419
rect 2851 414 2857 415
rect 2874 419 2880 420
rect 2874 415 2875 419
rect 2879 418 2880 419
rect 3011 419 3017 420
rect 3011 418 3012 419
rect 2879 416 3012 418
rect 2879 415 2880 416
rect 2874 414 2880 415
rect 3011 415 3012 416
rect 3016 415 3017 419
rect 3186 419 3192 420
rect 3011 414 3017 415
rect 3163 417 3169 418
rect 3163 413 3164 417
rect 3168 413 3169 417
rect 3186 415 3187 419
rect 3191 418 3192 419
rect 3315 419 3321 420
rect 3315 418 3316 419
rect 3191 416 3316 418
rect 3191 415 3192 416
rect 3186 414 3192 415
rect 3315 415 3316 416
rect 3320 415 3321 419
rect 3315 414 3321 415
rect 3338 419 3344 420
rect 3338 415 3339 419
rect 3343 418 3344 419
rect 3467 419 3473 420
rect 3467 418 3468 419
rect 3343 416 3468 418
rect 3343 415 3344 416
rect 3338 414 3344 415
rect 3467 415 3468 416
rect 3472 415 3473 419
rect 3467 414 3473 415
rect 3611 419 3617 420
rect 3611 415 3612 419
rect 3616 418 3617 419
rect 3646 419 3652 420
rect 3646 418 3647 419
rect 3616 416 3647 418
rect 3616 415 3617 416
rect 3611 414 3617 415
rect 3646 415 3647 416
rect 3651 415 3652 419
rect 3646 414 3652 415
rect 3763 419 3769 420
rect 3763 415 3764 419
rect 3768 418 3769 419
rect 3786 419 3792 420
rect 3786 418 3787 419
rect 3768 416 3787 418
rect 3768 415 3769 416
rect 3763 414 3769 415
rect 3786 415 3787 416
rect 3791 415 3792 419
rect 3786 414 3792 415
rect 3891 419 3897 420
rect 3891 415 3892 419
rect 3896 418 3897 419
rect 3914 419 3920 420
rect 3914 418 3915 419
rect 3896 416 3915 418
rect 3896 415 3897 416
rect 3891 414 3897 415
rect 3914 415 3915 416
rect 3919 415 3920 419
rect 3914 414 3920 415
rect 3163 412 3169 413
rect 3164 410 3166 412
rect 3498 411 3504 412
rect 3498 410 3499 411
rect 3164 408 3499 410
rect 3498 407 3499 408
rect 3503 407 3504 411
rect 3498 406 3504 407
rect 486 404 492 405
rect 110 401 116 402
rect 110 397 111 401
rect 115 397 116 401
rect 486 400 487 404
rect 491 400 492 404
rect 486 399 492 400
rect 582 404 588 405
rect 582 400 583 404
rect 587 400 588 404
rect 582 399 588 400
rect 686 404 692 405
rect 686 400 687 404
rect 691 400 692 404
rect 686 399 692 400
rect 790 404 796 405
rect 790 400 791 404
rect 795 400 796 404
rect 790 399 796 400
rect 894 404 900 405
rect 894 400 895 404
rect 899 400 900 404
rect 894 399 900 400
rect 998 404 1004 405
rect 998 400 999 404
rect 1003 400 1004 404
rect 998 399 1004 400
rect 1102 404 1108 405
rect 1102 400 1103 404
rect 1107 400 1108 404
rect 1102 399 1108 400
rect 1206 404 1212 405
rect 1206 400 1207 404
rect 1211 400 1212 404
rect 1206 399 1212 400
rect 1318 404 1324 405
rect 1318 400 1319 404
rect 1323 400 1324 404
rect 1318 399 1324 400
rect 1430 404 1436 405
rect 1430 400 1431 404
rect 1435 400 1436 404
rect 1430 399 1436 400
rect 2006 401 2012 402
rect 110 396 116 397
rect 2006 397 2007 401
rect 2011 397 2012 401
rect 2006 396 2012 397
rect 2342 396 2348 397
rect 562 395 568 396
rect 562 391 563 395
rect 567 391 568 395
rect 562 390 568 391
rect 658 395 664 396
rect 658 391 659 395
rect 663 391 664 395
rect 783 395 789 396
rect 783 394 784 395
rect 765 392 784 394
rect 658 390 664 391
rect 783 391 784 392
rect 788 391 789 395
rect 887 395 893 396
rect 887 394 888 395
rect 869 392 888 394
rect 783 390 789 391
rect 887 391 888 392
rect 892 391 893 395
rect 887 390 893 391
rect 966 395 972 396
rect 966 391 967 395
rect 971 391 972 395
rect 966 390 972 391
rect 1074 395 1080 396
rect 1074 391 1075 395
rect 1079 391 1080 395
rect 1074 390 1080 391
rect 1095 395 1101 396
rect 1095 391 1096 395
rect 1100 394 1101 395
rect 1186 395 1192 396
rect 1100 392 1145 394
rect 1100 391 1101 392
rect 1095 390 1101 391
rect 1186 391 1187 395
rect 1191 394 1192 395
rect 1394 395 1400 396
rect 1191 392 1249 394
rect 1191 391 1192 392
rect 1186 390 1192 391
rect 1394 391 1395 395
rect 1399 391 1400 395
rect 1394 390 1400 391
rect 1498 395 1504 396
rect 1498 391 1499 395
rect 1503 391 1504 395
rect 1498 390 1504 391
rect 2046 393 2052 394
rect 2046 389 2047 393
rect 2051 389 2052 393
rect 2342 392 2343 396
rect 2347 392 2348 396
rect 2342 391 2348 392
rect 2486 396 2492 397
rect 2486 392 2487 396
rect 2491 392 2492 396
rect 2486 391 2492 392
rect 2638 396 2644 397
rect 2638 392 2639 396
rect 2643 392 2644 396
rect 2638 391 2644 392
rect 2798 396 2804 397
rect 2798 392 2799 396
rect 2803 392 2804 396
rect 2798 391 2804 392
rect 2958 396 2964 397
rect 2958 392 2959 396
rect 2963 392 2964 396
rect 2958 391 2964 392
rect 3110 396 3116 397
rect 3110 392 3111 396
rect 3115 392 3116 396
rect 3110 391 3116 392
rect 3262 396 3268 397
rect 3262 392 3263 396
rect 3267 392 3268 396
rect 3262 391 3268 392
rect 3414 396 3420 397
rect 3414 392 3415 396
rect 3419 392 3420 396
rect 3414 391 3420 392
rect 3558 396 3564 397
rect 3558 392 3559 396
rect 3563 392 3564 396
rect 3558 391 3564 392
rect 3710 396 3716 397
rect 3710 392 3711 396
rect 3715 392 3716 396
rect 3710 391 3716 392
rect 3838 396 3844 397
rect 3838 392 3839 396
rect 3843 392 3844 396
rect 3838 391 3844 392
rect 3942 393 3948 394
rect 2046 388 2052 389
rect 3942 389 3943 393
rect 3947 389 3948 393
rect 3942 388 3948 389
rect 2418 387 2424 388
rect 486 385 492 386
rect 110 384 116 385
rect 110 380 111 384
rect 115 380 116 384
rect 486 381 487 385
rect 491 381 492 385
rect 486 380 492 381
rect 582 385 588 386
rect 582 381 583 385
rect 587 381 588 385
rect 582 380 588 381
rect 686 385 692 386
rect 686 381 687 385
rect 691 381 692 385
rect 686 380 692 381
rect 790 385 796 386
rect 790 381 791 385
rect 795 381 796 385
rect 790 380 796 381
rect 894 385 900 386
rect 894 381 895 385
rect 899 381 900 385
rect 894 380 900 381
rect 998 385 1004 386
rect 998 381 999 385
rect 1003 381 1004 385
rect 998 380 1004 381
rect 1102 385 1108 386
rect 1102 381 1103 385
rect 1107 381 1108 385
rect 1102 380 1108 381
rect 1206 385 1212 386
rect 1206 381 1207 385
rect 1211 381 1212 385
rect 1206 380 1212 381
rect 1318 385 1324 386
rect 1318 381 1319 385
rect 1323 381 1324 385
rect 1318 380 1324 381
rect 1430 385 1436 386
rect 1430 381 1431 385
rect 1435 381 1436 385
rect 1430 380 1436 381
rect 2006 384 2012 385
rect 2006 380 2007 384
rect 2011 380 2012 384
rect 2418 383 2419 387
rect 2423 383 2424 387
rect 2418 382 2424 383
rect 2562 387 2568 388
rect 2562 383 2563 387
rect 2567 383 2568 387
rect 2562 382 2568 383
rect 2714 387 2720 388
rect 2714 383 2715 387
rect 2719 383 2720 387
rect 2714 382 2720 383
rect 2874 387 2880 388
rect 2874 383 2875 387
rect 2879 383 2880 387
rect 2874 382 2880 383
rect 2898 387 2904 388
rect 2898 383 2899 387
rect 2903 386 2904 387
rect 3186 387 3192 388
rect 2903 384 3001 386
rect 2903 383 2904 384
rect 2898 382 2904 383
rect 3186 383 3187 387
rect 3191 383 3192 387
rect 3186 382 3192 383
rect 3338 387 3344 388
rect 3338 383 3339 387
rect 3343 383 3344 387
rect 3338 382 3344 383
rect 3490 387 3496 388
rect 3490 383 3491 387
rect 3495 383 3496 387
rect 3490 382 3496 383
rect 3498 387 3504 388
rect 3498 383 3499 387
rect 3503 386 3504 387
rect 3646 387 3652 388
rect 3503 384 3601 386
rect 3503 383 3504 384
rect 3498 382 3504 383
rect 3646 383 3647 387
rect 3651 386 3652 387
rect 3906 387 3912 388
rect 3651 384 3753 386
rect 3651 383 3652 384
rect 3646 382 3652 383
rect 3906 383 3907 387
rect 3911 383 3912 387
rect 3906 382 3912 383
rect 110 379 116 380
rect 2006 379 2012 380
rect 2342 377 2348 378
rect 2046 376 2052 377
rect 2046 372 2047 376
rect 2051 372 2052 376
rect 2342 373 2343 377
rect 2347 373 2348 377
rect 2342 372 2348 373
rect 2486 377 2492 378
rect 2486 373 2487 377
rect 2491 373 2492 377
rect 2486 372 2492 373
rect 2638 377 2644 378
rect 2638 373 2639 377
rect 2643 373 2644 377
rect 2638 372 2644 373
rect 2798 377 2804 378
rect 2798 373 2799 377
rect 2803 373 2804 377
rect 2798 372 2804 373
rect 2958 377 2964 378
rect 2958 373 2959 377
rect 2963 373 2964 377
rect 2958 372 2964 373
rect 3110 377 3116 378
rect 3110 373 3111 377
rect 3115 373 3116 377
rect 3110 372 3116 373
rect 3262 377 3268 378
rect 3262 373 3263 377
rect 3267 373 3268 377
rect 3262 372 3268 373
rect 3414 377 3420 378
rect 3414 373 3415 377
rect 3419 373 3420 377
rect 3414 372 3420 373
rect 3558 377 3564 378
rect 3558 373 3559 377
rect 3563 373 3564 377
rect 3558 372 3564 373
rect 3710 377 3716 378
rect 3710 373 3711 377
rect 3715 373 3716 377
rect 3710 372 3716 373
rect 3838 377 3844 378
rect 3838 373 3839 377
rect 3843 373 3844 377
rect 3838 372 3844 373
rect 3942 376 3948 377
rect 3942 372 3943 376
rect 3947 372 3948 376
rect 2046 371 2052 372
rect 3942 371 3948 372
rect 110 328 116 329
rect 2006 328 2012 329
rect 110 324 111 328
rect 115 324 116 328
rect 110 323 116 324
rect 326 327 332 328
rect 326 323 327 327
rect 331 323 332 327
rect 326 322 332 323
rect 462 327 468 328
rect 462 323 463 327
rect 467 323 468 327
rect 462 322 468 323
rect 614 327 620 328
rect 614 323 615 327
rect 619 323 620 327
rect 614 322 620 323
rect 766 327 772 328
rect 766 323 767 327
rect 771 323 772 327
rect 766 322 772 323
rect 918 327 924 328
rect 918 323 919 327
rect 923 323 924 327
rect 918 322 924 323
rect 1062 327 1068 328
rect 1062 323 1063 327
rect 1067 323 1068 327
rect 1062 322 1068 323
rect 1206 327 1212 328
rect 1206 323 1207 327
rect 1211 323 1212 327
rect 1206 322 1212 323
rect 1350 327 1356 328
rect 1350 323 1351 327
rect 1355 323 1356 327
rect 1494 327 1500 328
rect 1350 322 1356 323
rect 1418 323 1424 324
rect 858 319 864 320
rect 402 315 408 316
rect 110 311 116 312
rect 110 307 111 311
rect 115 307 116 311
rect 402 311 403 315
rect 407 311 408 315
rect 402 310 408 311
rect 538 315 544 316
rect 538 311 539 315
rect 543 311 544 315
rect 538 310 544 311
rect 690 315 696 316
rect 690 311 691 315
rect 695 311 696 315
rect 690 310 696 311
rect 842 315 848 316
rect 842 311 843 315
rect 847 311 848 315
rect 858 315 859 319
rect 863 318 864 319
rect 1418 319 1419 323
rect 1423 322 1424 323
rect 1494 323 1495 327
rect 1499 323 1500 327
rect 1494 322 1500 323
rect 1638 327 1644 328
rect 1638 323 1639 327
rect 1643 323 1644 327
rect 2006 324 2007 328
rect 2011 324 2012 328
rect 2006 323 2012 324
rect 1638 322 1644 323
rect 1423 320 1430 322
rect 2046 320 2052 321
rect 3942 320 3948 321
rect 1423 319 1424 320
rect 1418 318 1424 319
rect 863 316 961 318
rect 1428 317 1430 320
rect 1434 319 1440 320
rect 863 315 864 316
rect 858 314 864 315
rect 1138 315 1144 316
rect 842 310 848 311
rect 1138 311 1139 315
rect 1143 311 1144 315
rect 1138 310 1144 311
rect 1282 315 1288 316
rect 1282 311 1283 315
rect 1287 311 1288 315
rect 1434 315 1435 319
rect 1439 318 1440 319
rect 1578 319 1584 320
rect 1439 316 1537 318
rect 1439 315 1440 316
rect 1434 314 1440 315
rect 1578 315 1579 319
rect 1583 318 1584 319
rect 1583 316 1681 318
rect 2046 316 2047 320
rect 2051 316 2052 320
rect 1583 315 1584 316
rect 2046 315 2052 316
rect 2494 319 2500 320
rect 2494 315 2495 319
rect 2499 315 2500 319
rect 1578 314 1584 315
rect 2494 314 2500 315
rect 2638 319 2644 320
rect 2638 315 2639 319
rect 2643 315 2644 319
rect 2638 314 2644 315
rect 2798 319 2804 320
rect 2798 315 2799 319
rect 2803 315 2804 319
rect 2798 314 2804 315
rect 2958 319 2964 320
rect 2958 315 2959 319
rect 2963 315 2964 319
rect 2958 314 2964 315
rect 3118 319 3124 320
rect 3118 315 3119 319
rect 3123 315 3124 319
rect 3118 314 3124 315
rect 3270 319 3276 320
rect 3270 315 3271 319
rect 3275 315 3276 319
rect 3270 314 3276 315
rect 3422 319 3428 320
rect 3422 315 3423 319
rect 3427 315 3428 319
rect 3422 314 3428 315
rect 3566 319 3572 320
rect 3566 315 3567 319
rect 3571 315 3572 319
rect 3566 314 3572 315
rect 3710 319 3716 320
rect 3710 315 3711 319
rect 3715 315 3716 319
rect 3710 314 3716 315
rect 3838 319 3844 320
rect 3838 315 3839 319
rect 3843 315 3844 319
rect 3942 316 3943 320
rect 3947 316 3948 320
rect 3942 315 3948 316
rect 3838 314 3844 315
rect 1282 310 1288 311
rect 2006 311 2012 312
rect 110 306 116 307
rect 326 308 332 309
rect 326 304 327 308
rect 331 304 332 308
rect 326 303 332 304
rect 462 308 468 309
rect 462 304 463 308
rect 467 304 468 308
rect 462 303 468 304
rect 614 308 620 309
rect 614 304 615 308
rect 619 304 620 308
rect 614 303 620 304
rect 766 308 772 309
rect 766 304 767 308
rect 771 304 772 308
rect 766 303 772 304
rect 918 308 924 309
rect 918 304 919 308
rect 923 304 924 308
rect 918 303 924 304
rect 1062 308 1068 309
rect 1062 304 1063 308
rect 1067 304 1068 308
rect 1062 303 1068 304
rect 1206 308 1212 309
rect 1206 304 1207 308
rect 1211 304 1212 308
rect 1206 303 1212 304
rect 1350 308 1356 309
rect 1350 304 1351 308
rect 1355 304 1356 308
rect 1350 303 1356 304
rect 1494 308 1500 309
rect 1494 304 1495 308
rect 1499 304 1500 308
rect 1494 303 1500 304
rect 1638 308 1644 309
rect 1638 304 1639 308
rect 1643 304 1644 308
rect 2006 307 2007 311
rect 2011 307 2012 311
rect 3042 311 3048 312
rect 2006 306 2012 307
rect 2570 307 2576 308
rect 1638 303 1644 304
rect 2046 303 2052 304
rect 2046 299 2047 303
rect 2051 299 2052 303
rect 2570 303 2571 307
rect 2575 303 2576 307
rect 2570 302 2576 303
rect 2714 307 2720 308
rect 2714 303 2715 307
rect 2719 303 2720 307
rect 2714 302 2720 303
rect 2874 307 2880 308
rect 2874 303 2875 307
rect 2879 303 2880 307
rect 2874 302 2880 303
rect 3034 307 3040 308
rect 3034 303 3035 307
rect 3039 303 3040 307
rect 3042 307 3043 311
rect 3047 310 3048 311
rect 3786 311 3792 312
rect 3047 308 3161 310
rect 3047 307 3048 308
rect 3042 306 3048 307
rect 3346 307 3352 308
rect 3034 302 3040 303
rect 3346 303 3347 307
rect 3351 303 3352 307
rect 3346 302 3352 303
rect 3498 307 3504 308
rect 3498 303 3499 307
rect 3503 303 3504 307
rect 3498 302 3504 303
rect 3642 307 3648 308
rect 3642 303 3643 307
rect 3647 303 3648 307
rect 3786 307 3787 311
rect 3791 307 3792 311
rect 3786 306 3792 307
rect 3914 311 3920 312
rect 3914 307 3915 311
rect 3919 307 3920 311
rect 3914 306 3920 307
rect 3642 302 3648 303
rect 3942 303 3948 304
rect 2046 298 2052 299
rect 2494 300 2500 301
rect 2494 296 2495 300
rect 2499 296 2500 300
rect 2494 295 2500 296
rect 2638 300 2644 301
rect 2638 296 2639 300
rect 2643 296 2644 300
rect 2638 295 2644 296
rect 2798 300 2804 301
rect 2798 296 2799 300
rect 2803 296 2804 300
rect 2798 295 2804 296
rect 2958 300 2964 301
rect 2958 296 2959 300
rect 2963 296 2964 300
rect 2958 295 2964 296
rect 3118 300 3124 301
rect 3118 296 3119 300
rect 3123 296 3124 300
rect 3118 295 3124 296
rect 3270 300 3276 301
rect 3270 296 3271 300
rect 3275 296 3276 300
rect 3270 295 3276 296
rect 3422 300 3428 301
rect 3422 296 3423 300
rect 3427 296 3428 300
rect 3422 295 3428 296
rect 3566 300 3572 301
rect 3566 296 3567 300
rect 3571 296 3572 300
rect 3566 295 3572 296
rect 3710 300 3716 301
rect 3710 296 3711 300
rect 3715 296 3716 300
rect 3710 295 3716 296
rect 3838 300 3844 301
rect 3838 296 3839 300
rect 3843 296 3844 300
rect 3942 299 3943 303
rect 3947 299 3948 303
rect 3942 298 3948 299
rect 3838 295 3844 296
rect 402 287 408 288
rect 379 283 385 284
rect 379 279 380 283
rect 384 282 385 283
rect 402 283 403 287
rect 407 286 408 287
rect 515 287 521 288
rect 515 286 516 287
rect 407 284 516 286
rect 407 283 408 284
rect 402 282 408 283
rect 515 283 516 284
rect 520 283 521 287
rect 515 282 521 283
rect 538 287 544 288
rect 538 283 539 287
rect 543 286 544 287
rect 667 287 673 288
rect 667 286 668 287
rect 543 284 668 286
rect 543 283 544 284
rect 538 282 544 283
rect 667 283 668 284
rect 672 283 673 287
rect 667 282 673 283
rect 690 287 696 288
rect 690 283 691 287
rect 695 286 696 287
rect 819 287 825 288
rect 819 286 820 287
rect 695 284 820 286
rect 695 283 696 284
rect 690 282 696 283
rect 819 283 820 284
rect 824 283 825 287
rect 819 282 825 283
rect 842 287 848 288
rect 842 283 843 287
rect 847 286 848 287
rect 971 287 977 288
rect 971 286 972 287
rect 847 284 972 286
rect 847 283 848 284
rect 842 282 848 283
rect 971 283 972 284
rect 976 283 977 287
rect 971 282 977 283
rect 1074 287 1080 288
rect 1074 283 1075 287
rect 1079 286 1080 287
rect 1115 287 1121 288
rect 1115 286 1116 287
rect 1079 284 1116 286
rect 1079 283 1080 284
rect 1074 282 1080 283
rect 1115 283 1116 284
rect 1120 283 1121 287
rect 1115 282 1121 283
rect 1138 287 1144 288
rect 1138 283 1139 287
rect 1143 286 1144 287
rect 1259 287 1265 288
rect 1259 286 1260 287
rect 1143 284 1260 286
rect 1143 283 1144 284
rect 1138 282 1144 283
rect 1259 283 1260 284
rect 1264 283 1265 287
rect 1259 282 1265 283
rect 1403 287 1409 288
rect 1403 283 1404 287
rect 1408 286 1409 287
rect 1434 287 1440 288
rect 1434 286 1435 287
rect 1408 284 1435 286
rect 1408 283 1409 284
rect 1403 282 1409 283
rect 1434 283 1435 284
rect 1439 283 1440 287
rect 1434 282 1440 283
rect 1547 287 1553 288
rect 1547 283 1548 287
rect 1552 286 1553 287
rect 1578 287 1584 288
rect 1578 286 1579 287
rect 1552 284 1579 286
rect 1552 283 1553 284
rect 1547 282 1553 283
rect 1578 283 1579 284
rect 1583 283 1584 287
rect 1578 282 1584 283
rect 1586 283 1592 284
rect 384 280 398 282
rect 384 279 385 280
rect 379 278 385 279
rect 396 278 398 280
rect 831 279 837 280
rect 831 278 832 279
rect 396 276 832 278
rect 831 275 832 276
rect 836 275 837 279
rect 1586 279 1587 283
rect 1591 282 1592 283
rect 1691 283 1697 284
rect 1691 282 1692 283
rect 1591 280 1692 282
rect 1591 279 1592 280
rect 1586 278 1592 279
rect 1691 279 1692 280
rect 1696 279 1697 283
rect 1691 278 1697 279
rect 2547 279 2556 280
rect 831 274 837 275
rect 2547 275 2548 279
rect 2555 275 2556 279
rect 2547 274 2556 275
rect 2570 279 2576 280
rect 2570 275 2571 279
rect 2575 278 2576 279
rect 2691 279 2697 280
rect 2691 278 2692 279
rect 2575 276 2692 278
rect 2575 275 2576 276
rect 2570 274 2576 275
rect 2691 275 2692 276
rect 2696 275 2697 279
rect 2691 274 2697 275
rect 2714 279 2720 280
rect 2714 275 2715 279
rect 2719 278 2720 279
rect 2851 279 2857 280
rect 2851 278 2852 279
rect 2719 276 2852 278
rect 2719 275 2720 276
rect 2714 274 2720 275
rect 2851 275 2852 276
rect 2856 275 2857 279
rect 2851 274 2857 275
rect 2874 279 2880 280
rect 2874 275 2875 279
rect 2879 278 2880 279
rect 3011 279 3017 280
rect 3011 278 3012 279
rect 2879 276 3012 278
rect 2879 275 2880 276
rect 2874 274 2880 275
rect 3011 275 3012 276
rect 3016 275 3017 279
rect 3011 274 3017 275
rect 3034 279 3040 280
rect 3034 275 3035 279
rect 3039 278 3040 279
rect 3171 279 3177 280
rect 3171 278 3172 279
rect 3039 276 3172 278
rect 3039 275 3040 276
rect 3034 274 3040 275
rect 3171 275 3172 276
rect 3176 275 3177 279
rect 3346 279 3352 280
rect 3171 274 3177 275
rect 3323 275 3329 276
rect 3323 271 3324 275
rect 3328 274 3329 275
rect 3346 275 3347 279
rect 3351 278 3352 279
rect 3475 279 3481 280
rect 3475 278 3476 279
rect 3351 276 3476 278
rect 3351 275 3352 276
rect 3346 274 3352 275
rect 3475 275 3476 276
rect 3480 275 3481 279
rect 3475 274 3481 275
rect 3498 279 3504 280
rect 3498 275 3499 279
rect 3503 278 3504 279
rect 3619 279 3625 280
rect 3619 278 3620 279
rect 3503 276 3620 278
rect 3503 275 3504 276
rect 3498 274 3504 275
rect 3619 275 3620 276
rect 3624 275 3625 279
rect 3619 274 3625 275
rect 3763 279 3772 280
rect 3763 275 3764 279
rect 3771 275 3772 279
rect 3763 274 3772 275
rect 3891 275 3897 276
rect 3328 272 3342 274
rect 3328 271 3329 272
rect 3323 270 3329 271
rect 3340 270 3342 272
rect 3618 271 3624 272
rect 3618 270 3619 271
rect 3340 268 3619 270
rect 3618 267 3619 268
rect 3623 267 3624 271
rect 3891 271 3892 275
rect 3896 274 3897 275
rect 3906 275 3912 276
rect 3906 274 3907 275
rect 3896 272 3907 274
rect 3896 271 3897 272
rect 3891 270 3897 271
rect 3906 271 3907 272
rect 3911 271 3912 275
rect 3906 270 3912 271
rect 3618 266 3624 267
rect 242 263 248 264
rect 219 261 225 262
rect 219 257 220 261
rect 224 257 225 261
rect 242 259 243 263
rect 247 262 248 263
rect 379 263 385 264
rect 379 262 380 263
rect 247 260 380 262
rect 247 259 248 260
rect 242 258 248 259
rect 379 259 380 260
rect 384 259 385 263
rect 379 258 385 259
rect 402 263 408 264
rect 402 259 403 263
rect 407 262 408 263
rect 555 263 561 264
rect 555 262 556 263
rect 407 260 556 262
rect 407 259 408 260
rect 402 258 408 259
rect 555 259 556 260
rect 560 259 561 263
rect 555 258 561 259
rect 578 263 584 264
rect 578 259 579 263
rect 583 262 584 263
rect 739 263 745 264
rect 739 262 740 263
rect 583 260 740 262
rect 583 259 584 260
rect 578 258 584 259
rect 739 259 740 260
rect 744 259 745 263
rect 739 258 745 259
rect 823 263 829 264
rect 823 259 824 263
rect 828 262 829 263
rect 923 263 929 264
rect 923 262 924 263
rect 828 260 924 262
rect 828 259 829 260
rect 823 258 829 259
rect 923 259 924 260
rect 928 259 929 263
rect 1267 263 1273 264
rect 923 258 929 259
rect 1099 261 1105 262
rect 219 256 225 257
rect 1099 257 1100 261
rect 1104 257 1105 261
rect 1267 259 1268 263
rect 1272 262 1273 263
rect 1282 263 1288 264
rect 1282 262 1283 263
rect 1272 260 1283 262
rect 1272 259 1273 260
rect 1267 258 1273 259
rect 1282 259 1283 260
rect 1287 259 1288 263
rect 1282 258 1288 259
rect 1290 263 1296 264
rect 1290 259 1291 263
rect 1295 262 1296 263
rect 1419 263 1425 264
rect 1419 262 1420 263
rect 1295 260 1420 262
rect 1295 259 1296 260
rect 1290 258 1296 259
rect 1419 259 1420 260
rect 1424 259 1425 263
rect 1419 258 1425 259
rect 1563 263 1569 264
rect 1563 259 1564 263
rect 1568 262 1569 263
rect 1594 263 1600 264
rect 1594 262 1595 263
rect 1568 260 1595 262
rect 1568 259 1569 260
rect 1563 258 1569 259
rect 1594 259 1595 260
rect 1599 259 1600 263
rect 1594 258 1600 259
rect 1699 263 1705 264
rect 1699 259 1700 263
rect 1704 262 1705 263
rect 1730 263 1736 264
rect 1730 262 1731 263
rect 1704 260 1731 262
rect 1704 259 1705 260
rect 1699 258 1705 259
rect 1730 259 1731 260
rect 1735 259 1736 263
rect 1730 258 1736 259
rect 1835 263 1841 264
rect 1835 259 1836 263
rect 1840 262 1841 263
rect 1866 263 1872 264
rect 1866 262 1867 263
rect 1840 260 1867 262
rect 1840 259 1841 260
rect 1835 258 1841 259
rect 1866 259 1867 260
rect 1871 259 1872 263
rect 1866 258 1872 259
rect 1955 263 1961 264
rect 1955 259 1956 263
rect 1960 262 1961 263
rect 1986 263 1992 264
rect 1986 262 1987 263
rect 1960 260 1987 262
rect 1960 259 1961 260
rect 1955 258 1961 259
rect 1986 259 1987 260
rect 1991 259 1992 263
rect 1986 258 1992 259
rect 2123 263 2129 264
rect 2123 259 2124 263
rect 2128 262 2129 263
rect 2154 263 2160 264
rect 2154 262 2155 263
rect 2128 260 2155 262
rect 2128 259 2129 260
rect 2123 258 2129 259
rect 2154 259 2155 260
rect 2159 259 2160 263
rect 2154 258 2160 259
rect 2323 263 2329 264
rect 2323 259 2324 263
rect 2328 262 2329 263
rect 2538 263 2544 264
rect 2538 262 2539 263
rect 2328 260 2539 262
rect 2328 259 2329 260
rect 2323 258 2329 259
rect 2538 259 2539 260
rect 2543 259 2544 263
rect 2538 258 2544 259
rect 2547 263 2553 264
rect 2547 259 2548 263
rect 2552 262 2553 263
rect 2578 263 2584 264
rect 2578 262 2579 263
rect 2552 260 2579 262
rect 2552 259 2553 260
rect 2547 258 2553 259
rect 2578 259 2579 260
rect 2583 259 2584 263
rect 2578 258 2584 259
rect 2755 263 2761 264
rect 2755 259 2756 263
rect 2760 262 2761 263
rect 2799 263 2805 264
rect 2799 262 2800 263
rect 2760 260 2800 262
rect 2760 259 2761 260
rect 2755 258 2761 259
rect 2799 259 2800 260
rect 2804 259 2805 263
rect 2799 258 2805 259
rect 2955 263 2961 264
rect 2955 259 2956 263
rect 2960 262 2961 263
rect 3042 263 3048 264
rect 3042 262 3043 263
rect 2960 260 3043 262
rect 2960 259 2961 260
rect 2955 258 2961 259
rect 3042 259 3043 260
rect 3047 259 3048 263
rect 3170 263 3176 264
rect 3042 258 3048 259
rect 3147 261 3153 262
rect 1099 256 1105 257
rect 3147 257 3148 261
rect 3152 257 3153 261
rect 3170 259 3171 263
rect 3175 262 3176 263
rect 3339 263 3345 264
rect 3339 262 3340 263
rect 3175 260 3340 262
rect 3175 259 3176 260
rect 3170 258 3176 259
rect 3339 259 3340 260
rect 3344 259 3345 263
rect 3339 258 3345 259
rect 3362 263 3368 264
rect 3362 259 3363 263
rect 3367 262 3368 263
rect 3531 263 3537 264
rect 3531 262 3532 263
rect 3367 260 3532 262
rect 3367 259 3368 260
rect 3362 258 3368 259
rect 3531 259 3532 260
rect 3536 259 3537 263
rect 3531 258 3537 259
rect 3554 263 3560 264
rect 3554 259 3555 263
rect 3559 262 3560 263
rect 3723 263 3729 264
rect 3723 262 3724 263
rect 3559 260 3724 262
rect 3559 259 3560 260
rect 3554 258 3560 259
rect 3723 259 3724 260
rect 3728 259 3729 263
rect 3723 258 3729 259
rect 3891 263 3897 264
rect 3891 259 3892 263
rect 3896 262 3897 263
rect 3914 263 3920 264
rect 3914 262 3915 263
rect 3896 260 3915 262
rect 3896 259 3897 260
rect 3891 258 3897 259
rect 3914 259 3915 260
rect 3919 259 3920 263
rect 3914 258 3920 259
rect 3147 256 3153 257
rect 220 250 222 256
rect 1100 254 1102 256
rect 1338 255 1344 256
rect 1338 254 1339 255
rect 1100 252 1339 254
rect 858 251 864 252
rect 858 250 859 251
rect 220 248 859 250
rect 858 247 859 248
rect 863 247 864 251
rect 1338 251 1339 252
rect 1343 251 1344 255
rect 3148 254 3150 256
rect 3498 255 3504 256
rect 3498 254 3499 255
rect 3148 252 3499 254
rect 1338 250 1344 251
rect 3498 251 3499 252
rect 3503 251 3504 255
rect 3498 250 3504 251
rect 858 246 864 247
rect 166 240 172 241
rect 110 237 116 238
rect 110 233 111 237
rect 115 233 116 237
rect 166 236 167 240
rect 171 236 172 240
rect 166 235 172 236
rect 326 240 332 241
rect 326 236 327 240
rect 331 236 332 240
rect 326 235 332 236
rect 502 240 508 241
rect 502 236 503 240
rect 507 236 508 240
rect 502 235 508 236
rect 686 240 692 241
rect 686 236 687 240
rect 691 236 692 240
rect 686 235 692 236
rect 870 240 876 241
rect 870 236 871 240
rect 875 236 876 240
rect 870 235 876 236
rect 1046 240 1052 241
rect 1046 236 1047 240
rect 1051 236 1052 240
rect 1046 235 1052 236
rect 1214 240 1220 241
rect 1214 236 1215 240
rect 1219 236 1220 240
rect 1214 235 1220 236
rect 1366 240 1372 241
rect 1366 236 1367 240
rect 1371 236 1372 240
rect 1366 235 1372 236
rect 1510 240 1516 241
rect 1510 236 1511 240
rect 1515 236 1516 240
rect 1510 235 1516 236
rect 1646 240 1652 241
rect 1646 236 1647 240
rect 1651 236 1652 240
rect 1646 235 1652 236
rect 1782 240 1788 241
rect 1782 236 1783 240
rect 1787 236 1788 240
rect 1782 235 1788 236
rect 1902 240 1908 241
rect 1902 236 1903 240
rect 1907 236 1908 240
rect 2070 240 2076 241
rect 1902 235 1908 236
rect 2006 237 2012 238
rect 110 232 116 233
rect 2006 233 2007 237
rect 2011 233 2012 237
rect 2006 232 2012 233
rect 2046 237 2052 238
rect 2046 233 2047 237
rect 2051 233 2052 237
rect 2070 236 2071 240
rect 2075 236 2076 240
rect 2070 235 2076 236
rect 2270 240 2276 241
rect 2270 236 2271 240
rect 2275 236 2276 240
rect 2270 235 2276 236
rect 2494 240 2500 241
rect 2494 236 2495 240
rect 2499 236 2500 240
rect 2494 235 2500 236
rect 2702 240 2708 241
rect 2702 236 2703 240
rect 2707 236 2708 240
rect 2702 235 2708 236
rect 2902 240 2908 241
rect 2902 236 2903 240
rect 2907 236 2908 240
rect 2902 235 2908 236
rect 3094 240 3100 241
rect 3094 236 3095 240
rect 3099 236 3100 240
rect 3094 235 3100 236
rect 3286 240 3292 241
rect 3286 236 3287 240
rect 3291 236 3292 240
rect 3286 235 3292 236
rect 3478 240 3484 241
rect 3478 236 3479 240
rect 3483 236 3484 240
rect 3478 235 3484 236
rect 3670 240 3676 241
rect 3670 236 3671 240
rect 3675 236 3676 240
rect 3670 235 3676 236
rect 3838 240 3844 241
rect 3838 236 3839 240
rect 3843 236 3844 240
rect 3838 235 3844 236
rect 3942 237 3948 238
rect 2046 232 2052 233
rect 3942 233 3943 237
rect 3947 233 3948 237
rect 3942 232 3948 233
rect 242 231 248 232
rect 242 227 243 231
rect 247 227 248 231
rect 242 226 248 227
rect 402 231 408 232
rect 402 227 403 231
rect 407 227 408 231
rect 402 226 408 227
rect 578 231 584 232
rect 578 227 579 231
rect 583 227 584 231
rect 823 231 829 232
rect 823 230 824 231
rect 765 228 824 230
rect 578 226 584 227
rect 823 227 824 228
rect 828 227 829 231
rect 823 226 829 227
rect 831 231 837 232
rect 831 227 832 231
rect 836 230 837 231
rect 1114 231 1120 232
rect 836 228 913 230
rect 836 227 837 228
rect 831 226 837 227
rect 1114 227 1115 231
rect 1119 227 1120 231
rect 1114 226 1120 227
rect 1290 231 1296 232
rect 1290 227 1291 231
rect 1295 227 1296 231
rect 1290 226 1296 227
rect 1338 231 1344 232
rect 1338 227 1339 231
rect 1343 230 1344 231
rect 1586 231 1592 232
rect 1343 228 1409 230
rect 1343 227 1344 228
rect 1338 226 1344 227
rect 1586 227 1587 231
rect 1591 227 1592 231
rect 1586 226 1592 227
rect 1594 231 1600 232
rect 1594 227 1595 231
rect 1599 230 1600 231
rect 1730 231 1736 232
rect 1599 228 1689 230
rect 1599 227 1600 228
rect 1594 226 1600 227
rect 1730 227 1731 231
rect 1735 230 1736 231
rect 1866 231 1872 232
rect 1735 228 1825 230
rect 1735 227 1736 228
rect 1730 226 1736 227
rect 1866 227 1867 231
rect 1871 230 1872 231
rect 1986 231 1992 232
rect 1871 228 1945 230
rect 1871 227 1872 228
rect 1866 226 1872 227
rect 1986 227 1987 231
rect 1991 230 1992 231
rect 2154 231 2160 232
rect 1991 228 2113 230
rect 1991 227 1992 228
rect 1986 226 1992 227
rect 2154 227 2155 231
rect 2159 230 2160 231
rect 2578 231 2584 232
rect 2159 228 2313 230
rect 2159 227 2160 228
rect 2154 226 2160 227
rect 2572 222 2574 229
rect 2578 227 2579 231
rect 2583 230 2584 231
rect 2799 231 2805 232
rect 2583 228 2745 230
rect 2583 227 2584 228
rect 2578 226 2584 227
rect 2799 227 2800 231
rect 2804 230 2805 231
rect 3170 231 3176 232
rect 2804 228 2945 230
rect 2804 227 2805 228
rect 2799 226 2805 227
rect 3170 227 3171 231
rect 3175 227 3176 231
rect 3170 226 3176 227
rect 3362 231 3368 232
rect 3362 227 3363 231
rect 3367 227 3368 231
rect 3362 226 3368 227
rect 3554 231 3560 232
rect 3554 227 3555 231
rect 3559 227 3560 231
rect 3554 226 3560 227
rect 3618 231 3624 232
rect 3618 227 3619 231
rect 3623 230 3624 231
rect 3906 231 3912 232
rect 3623 228 3713 230
rect 3623 227 3624 228
rect 3618 226 3624 227
rect 3906 227 3907 231
rect 3911 227 3912 231
rect 3906 226 3912 227
rect 2614 223 2620 224
rect 2614 222 2615 223
rect 166 221 172 222
rect 110 220 116 221
rect 110 216 111 220
rect 115 216 116 220
rect 166 217 167 221
rect 171 217 172 221
rect 166 216 172 217
rect 326 221 332 222
rect 326 217 327 221
rect 331 217 332 221
rect 326 216 332 217
rect 502 221 508 222
rect 502 217 503 221
rect 507 217 508 221
rect 502 216 508 217
rect 686 221 692 222
rect 686 217 687 221
rect 691 217 692 221
rect 686 216 692 217
rect 870 221 876 222
rect 870 217 871 221
rect 875 217 876 221
rect 870 216 876 217
rect 1046 221 1052 222
rect 1046 217 1047 221
rect 1051 217 1052 221
rect 1046 216 1052 217
rect 1214 221 1220 222
rect 1214 217 1215 221
rect 1219 217 1220 221
rect 1214 216 1220 217
rect 1366 221 1372 222
rect 1366 217 1367 221
rect 1371 217 1372 221
rect 1366 216 1372 217
rect 1510 221 1516 222
rect 1510 217 1511 221
rect 1515 217 1516 221
rect 1510 216 1516 217
rect 1646 221 1652 222
rect 1646 217 1647 221
rect 1651 217 1652 221
rect 1646 216 1652 217
rect 1782 221 1788 222
rect 1782 217 1783 221
rect 1787 217 1788 221
rect 1782 216 1788 217
rect 1902 221 1908 222
rect 2070 221 2076 222
rect 1902 217 1903 221
rect 1907 217 1908 221
rect 1902 216 1908 217
rect 2006 220 2012 221
rect 2006 216 2007 220
rect 2011 216 2012 220
rect 110 215 116 216
rect 2006 215 2012 216
rect 2046 220 2052 221
rect 2046 216 2047 220
rect 2051 216 2052 220
rect 2070 217 2071 221
rect 2075 217 2076 221
rect 2070 216 2076 217
rect 2270 221 2276 222
rect 2270 217 2271 221
rect 2275 217 2276 221
rect 2270 216 2276 217
rect 2494 221 2500 222
rect 2494 217 2495 221
rect 2499 217 2500 221
rect 2572 220 2615 222
rect 2614 219 2615 220
rect 2619 219 2620 223
rect 2614 218 2620 219
rect 2702 221 2708 222
rect 2494 216 2500 217
rect 2702 217 2703 221
rect 2707 217 2708 221
rect 2702 216 2708 217
rect 2902 221 2908 222
rect 2902 217 2903 221
rect 2907 217 2908 221
rect 2902 216 2908 217
rect 3094 221 3100 222
rect 3094 217 3095 221
rect 3099 217 3100 221
rect 3094 216 3100 217
rect 3286 221 3292 222
rect 3286 217 3287 221
rect 3291 217 3292 221
rect 3286 216 3292 217
rect 3478 221 3484 222
rect 3478 217 3479 221
rect 3483 217 3484 221
rect 3478 216 3484 217
rect 3670 221 3676 222
rect 3670 217 3671 221
rect 3675 217 3676 221
rect 3670 216 3676 217
rect 3838 221 3844 222
rect 3838 217 3839 221
rect 3843 217 3844 221
rect 3838 216 3844 217
rect 3942 220 3948 221
rect 3942 216 3943 220
rect 3947 216 3948 220
rect 2046 215 2052 216
rect 3942 215 3948 216
rect 2046 144 2052 145
rect 3942 144 3948 145
rect 110 140 116 141
rect 2006 140 2012 141
rect 110 136 111 140
rect 115 136 116 140
rect 110 135 116 136
rect 134 139 140 140
rect 134 135 135 139
rect 139 135 140 139
rect 134 134 140 135
rect 230 139 236 140
rect 230 135 231 139
rect 235 135 236 139
rect 230 134 236 135
rect 326 139 332 140
rect 326 135 327 139
rect 331 135 332 139
rect 326 134 332 135
rect 422 139 428 140
rect 422 135 423 139
rect 427 135 428 139
rect 422 134 428 135
rect 526 139 532 140
rect 526 135 527 139
rect 531 135 532 139
rect 526 134 532 135
rect 646 139 652 140
rect 646 135 647 139
rect 651 135 652 139
rect 646 134 652 135
rect 774 139 780 140
rect 774 135 775 139
rect 779 135 780 139
rect 774 134 780 135
rect 902 139 908 140
rect 902 135 903 139
rect 907 135 908 139
rect 902 134 908 135
rect 1030 139 1036 140
rect 1030 135 1031 139
rect 1035 135 1036 139
rect 1030 134 1036 135
rect 1150 139 1156 140
rect 1150 135 1151 139
rect 1155 135 1156 139
rect 1150 134 1156 135
rect 1270 139 1276 140
rect 1270 135 1271 139
rect 1275 135 1276 139
rect 1270 134 1276 135
rect 1382 139 1388 140
rect 1382 135 1383 139
rect 1387 135 1388 139
rect 1382 134 1388 135
rect 1486 139 1492 140
rect 1486 135 1487 139
rect 1491 135 1492 139
rect 1486 134 1492 135
rect 1590 139 1596 140
rect 1590 135 1591 139
rect 1595 135 1596 139
rect 1590 134 1596 135
rect 1702 139 1708 140
rect 1702 135 1703 139
rect 1707 135 1708 139
rect 1702 134 1708 135
rect 1806 139 1812 140
rect 1806 135 1807 139
rect 1811 135 1812 139
rect 1806 134 1812 135
rect 1902 139 1908 140
rect 1902 135 1903 139
rect 1907 135 1908 139
rect 2006 136 2007 140
rect 2011 136 2012 140
rect 2046 140 2047 144
rect 2051 140 2052 144
rect 2046 139 2052 140
rect 2070 143 2076 144
rect 2070 139 2071 143
rect 2075 139 2076 143
rect 2070 138 2076 139
rect 2166 143 2172 144
rect 2166 139 2167 143
rect 2171 139 2172 143
rect 2166 138 2172 139
rect 2262 143 2268 144
rect 2262 139 2263 143
rect 2267 139 2268 143
rect 2262 138 2268 139
rect 2358 143 2364 144
rect 2358 139 2359 143
rect 2363 139 2364 143
rect 2358 138 2364 139
rect 2454 143 2460 144
rect 2454 139 2455 143
rect 2459 139 2460 143
rect 2454 138 2460 139
rect 2550 143 2556 144
rect 2550 139 2551 143
rect 2555 139 2556 143
rect 2550 138 2556 139
rect 2654 143 2660 144
rect 2654 139 2655 143
rect 2659 139 2660 143
rect 2654 138 2660 139
rect 2758 143 2764 144
rect 2758 139 2759 143
rect 2763 139 2764 143
rect 2758 138 2764 139
rect 2862 143 2868 144
rect 2862 139 2863 143
rect 2867 139 2868 143
rect 2862 138 2868 139
rect 2974 143 2980 144
rect 2974 139 2975 143
rect 2979 139 2980 143
rect 2974 138 2980 139
rect 3102 143 3108 144
rect 3102 139 3103 143
rect 3107 139 3108 143
rect 3102 138 3108 139
rect 3238 143 3244 144
rect 3238 139 3239 143
rect 3243 139 3244 143
rect 3238 138 3244 139
rect 3382 143 3388 144
rect 3382 139 3383 143
rect 3387 139 3388 143
rect 3382 138 3388 139
rect 3534 143 3540 144
rect 3534 139 3535 143
rect 3539 139 3540 143
rect 3534 138 3540 139
rect 3694 143 3700 144
rect 3694 139 3695 143
rect 3699 139 3700 143
rect 3694 138 3700 139
rect 3838 143 3844 144
rect 3838 139 3839 143
rect 3843 139 3844 143
rect 3942 140 3943 144
rect 3947 140 3948 144
rect 3942 139 3948 140
rect 3838 138 3844 139
rect 2006 135 2012 136
rect 2538 135 2544 136
rect 1902 134 1908 135
rect 858 131 864 132
rect 210 127 216 128
rect 110 123 116 124
rect 110 119 111 123
rect 115 119 116 123
rect 210 123 211 127
rect 215 123 216 127
rect 210 122 216 123
rect 306 127 312 128
rect 306 123 307 127
rect 311 123 312 127
rect 306 122 312 123
rect 402 127 408 128
rect 402 123 403 127
rect 407 123 408 127
rect 402 122 408 123
rect 498 127 504 128
rect 498 123 499 127
rect 503 123 504 127
rect 498 122 504 123
rect 602 127 608 128
rect 602 123 603 127
rect 607 123 608 127
rect 602 122 608 123
rect 722 127 728 128
rect 722 123 723 127
rect 727 123 728 127
rect 722 122 728 123
rect 850 127 856 128
rect 850 123 851 127
rect 855 123 856 127
rect 858 127 859 131
rect 863 130 864 131
rect 2146 131 2152 132
rect 863 128 945 130
rect 863 127 864 128
rect 858 126 864 127
rect 1122 127 1128 128
rect 1122 126 1123 127
rect 1109 124 1123 126
rect 850 122 856 123
rect 1122 123 1123 124
rect 1127 123 1128 127
rect 1122 122 1128 123
rect 1226 127 1232 128
rect 1226 123 1227 127
rect 1231 123 1232 127
rect 1226 122 1232 123
rect 1346 127 1352 128
rect 1346 123 1347 127
rect 1351 123 1352 127
rect 1346 122 1352 123
rect 1458 127 1464 128
rect 1458 123 1459 127
rect 1463 123 1464 127
rect 1458 122 1464 123
rect 1562 127 1568 128
rect 1562 123 1563 127
rect 1567 123 1568 127
rect 1562 122 1568 123
rect 1666 127 1672 128
rect 1666 123 1667 127
rect 1671 123 1672 127
rect 1666 122 1672 123
rect 1778 127 1784 128
rect 1778 123 1779 127
rect 1783 123 1784 127
rect 1778 122 1784 123
rect 1882 127 1888 128
rect 1882 123 1883 127
rect 1887 123 1888 127
rect 1882 122 1888 123
rect 1978 127 1984 128
rect 1978 123 1979 127
rect 1983 123 1984 127
rect 2046 127 2052 128
rect 1978 122 1984 123
rect 2006 123 2012 124
rect 110 118 116 119
rect 134 120 140 121
rect 134 116 135 120
rect 139 116 140 120
rect 134 115 140 116
rect 230 120 236 121
rect 230 116 231 120
rect 235 116 236 120
rect 230 115 236 116
rect 326 120 332 121
rect 326 116 327 120
rect 331 116 332 120
rect 326 115 332 116
rect 422 120 428 121
rect 422 116 423 120
rect 427 116 428 120
rect 422 115 428 116
rect 526 120 532 121
rect 526 116 527 120
rect 531 116 532 120
rect 526 115 532 116
rect 646 120 652 121
rect 646 116 647 120
rect 651 116 652 120
rect 646 115 652 116
rect 774 120 780 121
rect 774 116 775 120
rect 779 116 780 120
rect 774 115 780 116
rect 902 120 908 121
rect 902 116 903 120
rect 907 116 908 120
rect 902 115 908 116
rect 1030 120 1036 121
rect 1030 116 1031 120
rect 1035 116 1036 120
rect 1030 115 1036 116
rect 1150 120 1156 121
rect 1150 116 1151 120
rect 1155 116 1156 120
rect 1150 115 1156 116
rect 1270 120 1276 121
rect 1270 116 1271 120
rect 1275 116 1276 120
rect 1270 115 1276 116
rect 1382 120 1388 121
rect 1382 116 1383 120
rect 1387 116 1388 120
rect 1382 115 1388 116
rect 1486 120 1492 121
rect 1486 116 1487 120
rect 1491 116 1492 120
rect 1486 115 1492 116
rect 1590 120 1596 121
rect 1590 116 1591 120
rect 1595 116 1596 120
rect 1590 115 1596 116
rect 1702 120 1708 121
rect 1702 116 1703 120
rect 1707 116 1708 120
rect 1702 115 1708 116
rect 1806 120 1812 121
rect 1806 116 1807 120
rect 1811 116 1812 120
rect 1806 115 1812 116
rect 1902 120 1908 121
rect 1902 116 1903 120
rect 1907 116 1908 120
rect 2006 119 2007 123
rect 2011 119 2012 123
rect 2046 123 2047 127
rect 2051 123 2052 127
rect 2146 127 2147 131
rect 2151 127 2152 131
rect 2146 126 2152 127
rect 2242 131 2248 132
rect 2242 127 2243 131
rect 2247 127 2248 131
rect 2242 126 2248 127
rect 2338 131 2344 132
rect 2338 127 2339 131
rect 2343 127 2344 131
rect 2338 126 2344 127
rect 2434 131 2440 132
rect 2434 127 2435 131
rect 2439 127 2440 131
rect 2434 126 2440 127
rect 2530 131 2536 132
rect 2530 127 2531 131
rect 2535 127 2536 131
rect 2538 131 2539 135
rect 2543 134 2544 135
rect 3498 135 3504 136
rect 2543 132 2593 134
rect 2543 131 2544 132
rect 2538 130 2544 131
rect 2730 131 2736 132
rect 2530 126 2536 127
rect 2730 127 2731 131
rect 2735 127 2736 131
rect 2730 126 2736 127
rect 2834 131 2840 132
rect 2834 127 2835 131
rect 2839 127 2840 131
rect 2834 126 2840 127
rect 2938 131 2944 132
rect 2938 127 2939 131
rect 2943 127 2944 131
rect 2938 126 2944 127
rect 3050 131 3056 132
rect 3050 127 3051 131
rect 3055 127 3056 131
rect 3050 126 3056 127
rect 3178 131 3184 132
rect 3178 127 3179 131
rect 3183 127 3184 131
rect 3178 126 3184 127
rect 3314 131 3320 132
rect 3314 127 3315 131
rect 3319 127 3320 131
rect 3314 126 3320 127
rect 3458 131 3464 132
rect 3458 127 3459 131
rect 3463 127 3464 131
rect 3498 131 3499 135
rect 3503 134 3504 135
rect 3914 135 3920 136
rect 3503 132 3577 134
rect 3503 131 3504 132
rect 3498 130 3504 131
rect 3770 131 3776 132
rect 3458 126 3464 127
rect 3770 127 3771 131
rect 3775 127 3776 131
rect 3914 131 3915 135
rect 3919 131 3920 135
rect 3914 130 3920 131
rect 3770 126 3776 127
rect 3942 127 3948 128
rect 2046 122 2052 123
rect 2070 124 2076 125
rect 2070 120 2071 124
rect 2075 120 2076 124
rect 2070 119 2076 120
rect 2166 124 2172 125
rect 2166 120 2167 124
rect 2171 120 2172 124
rect 2166 119 2172 120
rect 2262 124 2268 125
rect 2262 120 2263 124
rect 2267 120 2268 124
rect 2262 119 2268 120
rect 2358 124 2364 125
rect 2358 120 2359 124
rect 2363 120 2364 124
rect 2358 119 2364 120
rect 2454 124 2460 125
rect 2454 120 2455 124
rect 2459 120 2460 124
rect 2454 119 2460 120
rect 2550 124 2556 125
rect 2550 120 2551 124
rect 2555 120 2556 124
rect 2550 119 2556 120
rect 2654 124 2660 125
rect 2654 120 2655 124
rect 2659 120 2660 124
rect 2654 119 2660 120
rect 2758 124 2764 125
rect 2758 120 2759 124
rect 2763 120 2764 124
rect 2758 119 2764 120
rect 2862 124 2868 125
rect 2862 120 2863 124
rect 2867 120 2868 124
rect 2862 119 2868 120
rect 2974 124 2980 125
rect 2974 120 2975 124
rect 2979 120 2980 124
rect 2974 119 2980 120
rect 3102 124 3108 125
rect 3102 120 3103 124
rect 3107 120 3108 124
rect 3102 119 3108 120
rect 3238 124 3244 125
rect 3238 120 3239 124
rect 3243 120 3244 124
rect 3238 119 3244 120
rect 3382 124 3388 125
rect 3382 120 3383 124
rect 3387 120 3388 124
rect 3382 119 3388 120
rect 3534 124 3540 125
rect 3534 120 3535 124
rect 3539 120 3540 124
rect 3534 119 3540 120
rect 3694 124 3700 125
rect 3694 120 3695 124
rect 3699 120 3700 124
rect 3694 119 3700 120
rect 3838 124 3844 125
rect 3838 120 3839 124
rect 3843 120 3844 124
rect 3942 123 3943 127
rect 3947 123 3948 127
rect 3942 122 3948 123
rect 3838 119 3844 120
rect 2006 118 2012 119
rect 1902 115 1908 116
rect 1978 103 1984 104
rect 210 99 216 100
rect 210 95 211 99
rect 215 98 216 99
rect 283 99 289 100
rect 283 98 284 99
rect 215 96 284 98
rect 215 95 216 96
rect 210 94 216 95
rect 283 95 284 96
rect 288 95 289 99
rect 283 94 289 95
rect 306 99 312 100
rect 306 95 307 99
rect 311 98 312 99
rect 379 99 385 100
rect 379 98 380 99
rect 311 96 380 98
rect 311 95 312 96
rect 306 94 312 95
rect 379 95 380 96
rect 384 95 385 99
rect 379 94 385 95
rect 402 99 408 100
rect 402 95 403 99
rect 407 98 408 99
rect 475 99 481 100
rect 475 98 476 99
rect 407 96 476 98
rect 407 95 408 96
rect 402 94 408 95
rect 475 95 476 96
rect 480 95 481 99
rect 475 94 481 95
rect 498 99 504 100
rect 498 95 499 99
rect 503 98 504 99
rect 579 99 585 100
rect 579 98 580 99
rect 503 96 580 98
rect 503 95 504 96
rect 498 94 504 95
rect 579 95 580 96
rect 584 95 585 99
rect 579 94 585 95
rect 602 99 608 100
rect 602 95 603 99
rect 607 98 608 99
rect 699 99 705 100
rect 699 98 700 99
rect 607 96 700 98
rect 607 95 608 96
rect 602 94 608 95
rect 699 95 700 96
rect 704 95 705 99
rect 699 94 705 95
rect 722 99 728 100
rect 722 95 723 99
rect 727 98 728 99
rect 827 99 833 100
rect 827 98 828 99
rect 727 96 828 98
rect 727 95 728 96
rect 722 94 728 95
rect 827 95 828 96
rect 832 95 833 99
rect 827 94 833 95
rect 850 99 856 100
rect 850 95 851 99
rect 855 98 856 99
rect 955 99 961 100
rect 955 98 956 99
rect 855 96 956 98
rect 855 95 856 96
rect 850 94 856 95
rect 955 95 956 96
rect 960 95 961 99
rect 955 94 961 95
rect 1083 99 1089 100
rect 1083 95 1084 99
rect 1088 98 1089 99
rect 1114 99 1120 100
rect 1114 98 1115 99
rect 1088 96 1115 98
rect 1088 95 1089 96
rect 1083 94 1089 95
rect 1114 95 1115 96
rect 1119 95 1120 99
rect 1114 94 1120 95
rect 1122 99 1128 100
rect 1122 95 1123 99
rect 1127 98 1128 99
rect 1203 99 1209 100
rect 1203 98 1204 99
rect 1127 96 1204 98
rect 1127 95 1128 96
rect 1122 94 1128 95
rect 1203 95 1204 96
rect 1208 95 1209 99
rect 1203 94 1209 95
rect 1226 99 1232 100
rect 1226 95 1227 99
rect 1231 98 1232 99
rect 1323 99 1329 100
rect 1323 98 1324 99
rect 1231 96 1324 98
rect 1231 95 1232 96
rect 1226 94 1232 95
rect 1323 95 1324 96
rect 1328 95 1329 99
rect 1323 94 1329 95
rect 1346 99 1352 100
rect 1346 95 1347 99
rect 1351 98 1352 99
rect 1435 99 1441 100
rect 1435 98 1436 99
rect 1351 96 1436 98
rect 1351 95 1352 96
rect 1346 94 1352 95
rect 1435 95 1436 96
rect 1440 95 1441 99
rect 1435 94 1441 95
rect 1458 99 1464 100
rect 1458 95 1459 99
rect 1463 98 1464 99
rect 1539 99 1545 100
rect 1539 98 1540 99
rect 1463 96 1540 98
rect 1463 95 1464 96
rect 1458 94 1464 95
rect 1539 95 1540 96
rect 1544 95 1545 99
rect 1539 94 1545 95
rect 1562 99 1568 100
rect 1562 95 1563 99
rect 1567 98 1568 99
rect 1643 99 1649 100
rect 1643 98 1644 99
rect 1567 96 1644 98
rect 1567 95 1568 96
rect 1562 94 1568 95
rect 1643 95 1644 96
rect 1648 95 1649 99
rect 1643 94 1649 95
rect 1666 99 1672 100
rect 1666 95 1667 99
rect 1671 98 1672 99
rect 1755 99 1761 100
rect 1755 98 1756 99
rect 1671 96 1756 98
rect 1671 95 1672 96
rect 1666 94 1672 95
rect 1755 95 1756 96
rect 1760 95 1761 99
rect 1755 94 1761 95
rect 1778 99 1784 100
rect 1778 95 1779 99
rect 1783 98 1784 99
rect 1859 99 1865 100
rect 1859 98 1860 99
rect 1783 96 1860 98
rect 1783 95 1784 96
rect 1778 94 1784 95
rect 1859 95 1860 96
rect 1864 95 1865 99
rect 1859 94 1865 95
rect 1882 99 1888 100
rect 1882 95 1883 99
rect 1887 98 1888 99
rect 1955 99 1961 100
rect 1955 98 1956 99
rect 1887 96 1956 98
rect 1887 95 1888 96
rect 1882 94 1888 95
rect 1955 95 1956 96
rect 1960 95 1961 99
rect 1978 99 1979 103
rect 1983 102 1984 103
rect 2123 103 2129 104
rect 2123 102 2124 103
rect 1983 100 2124 102
rect 1983 99 1984 100
rect 1978 98 1984 99
rect 2123 99 2124 100
rect 2128 99 2129 103
rect 2123 98 2129 99
rect 2146 103 2152 104
rect 2146 99 2147 103
rect 2151 102 2152 103
rect 2219 103 2225 104
rect 2219 102 2220 103
rect 2151 100 2220 102
rect 2151 99 2152 100
rect 2146 98 2152 99
rect 2219 99 2220 100
rect 2224 99 2225 103
rect 2219 98 2225 99
rect 2242 103 2248 104
rect 2242 99 2243 103
rect 2247 102 2248 103
rect 2315 103 2321 104
rect 2315 102 2316 103
rect 2247 100 2316 102
rect 2247 99 2248 100
rect 2242 98 2248 99
rect 2315 99 2316 100
rect 2320 99 2321 103
rect 2315 98 2321 99
rect 2338 103 2344 104
rect 2338 99 2339 103
rect 2343 102 2344 103
rect 2411 103 2417 104
rect 2411 102 2412 103
rect 2343 100 2412 102
rect 2343 99 2344 100
rect 2338 98 2344 99
rect 2411 99 2412 100
rect 2416 99 2417 103
rect 2411 98 2417 99
rect 2434 103 2440 104
rect 2434 99 2435 103
rect 2439 102 2440 103
rect 2507 103 2513 104
rect 2507 102 2508 103
rect 2439 100 2508 102
rect 2439 99 2440 100
rect 2434 98 2440 99
rect 2507 99 2508 100
rect 2512 99 2513 103
rect 2507 98 2513 99
rect 2530 103 2536 104
rect 2530 99 2531 103
rect 2535 102 2536 103
rect 2603 103 2609 104
rect 2603 102 2604 103
rect 2535 100 2604 102
rect 2535 99 2536 100
rect 2530 98 2536 99
rect 2603 99 2604 100
rect 2608 99 2609 103
rect 2603 98 2609 99
rect 2614 103 2620 104
rect 2614 99 2615 103
rect 2619 102 2620 103
rect 2707 103 2713 104
rect 2707 102 2708 103
rect 2619 100 2708 102
rect 2619 99 2620 100
rect 2614 98 2620 99
rect 2707 99 2708 100
rect 2712 99 2713 103
rect 2707 98 2713 99
rect 2730 103 2736 104
rect 2730 99 2731 103
rect 2735 102 2736 103
rect 2811 103 2817 104
rect 2811 102 2812 103
rect 2735 100 2812 102
rect 2735 99 2736 100
rect 2730 98 2736 99
rect 2811 99 2812 100
rect 2816 99 2817 103
rect 2811 98 2817 99
rect 2834 103 2840 104
rect 2834 99 2835 103
rect 2839 102 2840 103
rect 2915 103 2921 104
rect 2915 102 2916 103
rect 2839 100 2916 102
rect 2839 99 2840 100
rect 2834 98 2840 99
rect 2915 99 2916 100
rect 2920 99 2921 103
rect 2915 98 2921 99
rect 2938 103 2944 104
rect 2938 99 2939 103
rect 2943 102 2944 103
rect 3027 103 3033 104
rect 3027 102 3028 103
rect 2943 100 3028 102
rect 2943 99 2944 100
rect 2938 98 2944 99
rect 3027 99 3028 100
rect 3032 99 3033 103
rect 3027 98 3033 99
rect 3050 103 3056 104
rect 3050 99 3051 103
rect 3055 102 3056 103
rect 3155 103 3161 104
rect 3155 102 3156 103
rect 3055 100 3156 102
rect 3055 99 3056 100
rect 3050 98 3056 99
rect 3155 99 3156 100
rect 3160 99 3161 103
rect 3155 98 3161 99
rect 3178 103 3184 104
rect 3178 99 3179 103
rect 3183 102 3184 103
rect 3291 103 3297 104
rect 3291 102 3292 103
rect 3183 100 3292 102
rect 3183 99 3184 100
rect 3178 98 3184 99
rect 3291 99 3292 100
rect 3296 99 3297 103
rect 3291 98 3297 99
rect 3314 103 3320 104
rect 3314 99 3315 103
rect 3319 102 3320 103
rect 3435 103 3441 104
rect 3435 102 3436 103
rect 3319 100 3436 102
rect 3319 99 3320 100
rect 3314 98 3320 99
rect 3435 99 3436 100
rect 3440 99 3441 103
rect 3435 98 3441 99
rect 3458 103 3464 104
rect 3458 99 3459 103
rect 3463 102 3464 103
rect 3587 103 3593 104
rect 3587 102 3588 103
rect 3463 100 3588 102
rect 3463 99 3464 100
rect 3458 98 3464 99
rect 3587 99 3588 100
rect 3592 99 3593 103
rect 3587 98 3593 99
rect 3642 103 3648 104
rect 3642 99 3643 103
rect 3647 102 3648 103
rect 3747 103 3753 104
rect 3747 102 3748 103
rect 3647 100 3748 102
rect 3647 99 3648 100
rect 3642 98 3648 99
rect 3747 99 3748 100
rect 3752 99 3753 103
rect 3747 98 3753 99
rect 3770 103 3776 104
rect 3770 99 3771 103
rect 3775 102 3776 103
rect 3891 103 3897 104
rect 3891 102 3892 103
rect 3775 100 3892 102
rect 3775 99 3776 100
rect 3770 98 3776 99
rect 3891 99 3892 100
rect 3896 99 3897 103
rect 3891 98 3897 99
rect 1955 94 1961 95
<< m3c >>
rect 2147 4007 2151 4011
rect 2243 4007 2247 4011
rect 111 4000 115 4004
rect 1519 3999 1523 4003
rect 1615 3999 1619 4003
rect 1711 3999 1715 4003
rect 1807 3999 1811 4003
rect 1903 3999 1907 4003
rect 2007 4000 2011 4004
rect 111 3983 115 3987
rect 1691 3987 1695 3991
rect 1787 3987 1791 3991
rect 1883 3987 1887 3991
rect 1519 3980 1523 3984
rect 1615 3980 1619 3984
rect 1711 3980 1715 3984
rect 1807 3980 1811 3984
rect 1903 3980 1907 3984
rect 2007 3983 2011 3987
rect 2047 3981 2051 3985
rect 2071 3984 2075 3988
rect 2167 3984 2171 3988
rect 2263 3984 2267 3988
rect 3943 3981 3947 3985
rect 2147 3975 2151 3979
rect 2243 3975 2247 3979
rect 2047 3964 2051 3968
rect 2071 3965 2075 3969
rect 2167 3965 2171 3969
rect 2263 3965 2267 3969
rect 3943 3964 3947 3968
rect 1691 3959 1695 3963
rect 1787 3959 1791 3963
rect 1883 3959 1887 3963
rect 267 3943 271 3947
rect 275 3943 279 3947
rect 371 3943 375 3947
rect 467 3943 471 3947
rect 571 3943 575 3947
rect 691 3943 695 3947
rect 819 3943 823 3947
rect 947 3943 951 3947
rect 1179 3943 1180 3947
rect 1180 3943 1183 3947
rect 1203 3943 1207 3947
rect 1331 3943 1335 3947
rect 1459 3943 1463 3947
rect 1587 3943 1591 3947
rect 111 3917 115 3921
rect 199 3920 203 3924
rect 295 3920 299 3924
rect 391 3920 395 3924
rect 495 3920 499 3924
rect 615 3920 619 3924
rect 743 3920 747 3924
rect 871 3920 875 3924
rect 999 3920 1003 3924
rect 1127 3920 1131 3924
rect 1255 3920 1259 3924
rect 1383 3920 1387 3924
rect 1511 3920 1515 3924
rect 1647 3920 1651 3924
rect 2007 3917 2011 3921
rect 275 3911 279 3915
rect 371 3911 375 3915
rect 467 3911 471 3915
rect 571 3911 575 3915
rect 691 3911 695 3915
rect 819 3911 823 3915
rect 947 3911 951 3915
rect 955 3911 959 3915
rect 1203 3911 1207 3915
rect 1331 3911 1335 3915
rect 1459 3911 1463 3915
rect 1587 3911 1591 3915
rect 2047 3912 2051 3916
rect 2159 3911 2163 3915
rect 2287 3911 2291 3915
rect 2415 3911 2419 3915
rect 2551 3911 2555 3915
rect 2687 3911 2691 3915
rect 2823 3911 2827 3915
rect 2951 3911 2955 3915
rect 3071 3911 3075 3915
rect 3191 3911 3195 3915
rect 3303 3911 3307 3915
rect 3407 3911 3411 3915
rect 3519 3911 3523 3915
rect 3631 3911 3635 3915
rect 3743 3911 3747 3915
rect 3943 3912 3947 3916
rect 111 3900 115 3904
rect 199 3901 203 3905
rect 295 3901 299 3905
rect 391 3901 395 3905
rect 495 3901 499 3905
rect 615 3901 619 3905
rect 743 3901 747 3905
rect 871 3901 875 3905
rect 999 3901 1003 3905
rect 1127 3901 1131 3905
rect 1255 3901 1259 3905
rect 1383 3901 1387 3905
rect 1511 3901 1515 3905
rect 1647 3901 1651 3905
rect 2007 3900 2011 3904
rect 2047 3895 2051 3899
rect 2271 3899 2275 3903
rect 2363 3899 2367 3903
rect 2491 3899 2495 3903
rect 2627 3899 2631 3903
rect 2783 3899 2787 3903
rect 2899 3899 2903 3903
rect 3027 3899 3031 3903
rect 3147 3899 3151 3903
rect 3267 3899 3271 3903
rect 3379 3899 3383 3903
rect 3483 3899 3487 3903
rect 3595 3899 3599 3903
rect 3707 3899 3711 3903
rect 3715 3903 3719 3907
rect 2159 3892 2163 3896
rect 2287 3892 2291 3896
rect 2415 3892 2419 3896
rect 2551 3892 2555 3896
rect 2687 3892 2691 3896
rect 2823 3892 2827 3896
rect 2951 3892 2955 3896
rect 3071 3892 3075 3896
rect 3191 3892 3195 3896
rect 3303 3892 3307 3896
rect 3407 3892 3411 3896
rect 3519 3892 3523 3896
rect 3631 3892 3635 3896
rect 3743 3892 3747 3896
rect 3943 3895 3947 3899
rect 2271 3871 2275 3875
rect 2363 3871 2367 3875
rect 2491 3871 2495 3875
rect 2627 3871 2631 3875
rect 2899 3871 2903 3875
rect 3027 3871 3031 3875
rect 3147 3871 3151 3875
rect 3267 3871 3271 3875
rect 3379 3871 3383 3875
rect 3483 3871 3487 3875
rect 3595 3871 3599 3875
rect 3707 3871 3711 3875
rect 111 3848 115 3852
rect 335 3847 339 3851
rect 455 3847 459 3851
rect 583 3847 587 3851
rect 719 3847 723 3851
rect 847 3847 851 3851
rect 975 3847 979 3851
rect 1103 3847 1107 3851
rect 1231 3847 1235 3851
rect 1359 3847 1363 3851
rect 1487 3847 1491 3851
rect 2007 3848 2011 3852
rect 2295 3847 2299 3851
rect 2427 3847 2431 3851
rect 2571 3847 2575 3851
rect 2783 3847 2787 3851
rect 3099 3847 3103 3851
rect 3311 3847 3315 3851
rect 3395 3847 3399 3851
rect 3711 3847 3712 3851
rect 3712 3847 3715 3851
rect 267 3839 271 3843
rect 111 3831 115 3835
rect 795 3835 799 3839
rect 923 3835 927 3839
rect 1051 3835 1055 3839
rect 1179 3839 1183 3843
rect 1215 3839 1219 3843
rect 1343 3839 1347 3843
rect 335 3828 339 3832
rect 455 3828 459 3832
rect 583 3828 587 3832
rect 719 3828 723 3832
rect 847 3828 851 3832
rect 975 3828 979 3832
rect 1103 3828 1107 3832
rect 1231 3828 1235 3832
rect 1359 3828 1363 3832
rect 1487 3828 1491 3832
rect 2007 3831 2011 3835
rect 2047 3821 2051 3825
rect 2207 3824 2211 3828
rect 2343 3824 2347 3828
rect 2487 3824 2491 3828
rect 2647 3824 2651 3828
rect 2823 3824 2827 3828
rect 3015 3824 3019 3828
rect 3223 3824 3227 3828
rect 3439 3824 3443 3828
rect 3655 3824 3659 3828
rect 3943 3821 3947 3825
rect 575 3799 579 3803
rect 955 3815 959 3819
rect 2275 3815 2279 3819
rect 2295 3815 2299 3819
rect 2427 3815 2431 3819
rect 2571 3815 2575 3819
rect 3099 3815 3103 3819
rect 3311 3815 3315 3819
rect 3731 3815 3735 3819
rect 795 3807 799 3811
rect 923 3807 927 3811
rect 1215 3807 1219 3811
rect 1343 3807 1347 3811
rect 1507 3803 1511 3807
rect 2047 3804 2051 3808
rect 2207 3805 2211 3809
rect 2343 3805 2347 3809
rect 2487 3805 2491 3809
rect 2647 3805 2651 3809
rect 2823 3805 2827 3809
rect 3015 3805 3019 3809
rect 3223 3805 3227 3809
rect 3439 3805 3443 3809
rect 3655 3805 3659 3809
rect 3943 3804 3947 3808
rect 591 3787 595 3791
rect 699 3787 703 3791
rect 819 3787 823 3791
rect 903 3787 907 3791
rect 1051 3787 1052 3791
rect 1052 3787 1055 3791
rect 1075 3787 1079 3791
rect 1407 3787 1411 3791
rect 1571 3787 1575 3791
rect 1515 3779 1519 3783
rect 111 3761 115 3765
rect 503 3764 507 3768
rect 615 3764 619 3768
rect 735 3764 739 3768
rect 863 3764 867 3768
rect 999 3764 1003 3768
rect 1143 3764 1147 3768
rect 1287 3764 1291 3768
rect 1431 3764 1435 3768
rect 1583 3764 1587 3768
rect 2007 3761 2011 3765
rect 575 3755 579 3759
rect 591 3755 595 3759
rect 699 3755 703 3759
rect 819 3755 823 3759
rect 1075 3755 1079 3759
rect 1219 3755 1223 3759
rect 1407 3755 1411 3759
rect 1507 3755 1511 3759
rect 1515 3755 1519 3759
rect 2047 3752 2051 3756
rect 2191 3751 2195 3755
rect 2375 3751 2379 3755
rect 2559 3751 2563 3755
rect 2743 3751 2747 3755
rect 2935 3751 2939 3755
rect 3127 3751 3131 3755
rect 3319 3751 3323 3755
rect 3511 3751 3515 3755
rect 3711 3751 3715 3755
rect 3943 3752 3947 3756
rect 111 3744 115 3748
rect 503 3745 507 3749
rect 615 3745 619 3749
rect 735 3745 739 3749
rect 863 3745 867 3749
rect 999 3745 1003 3749
rect 1143 3745 1147 3749
rect 1287 3745 1291 3749
rect 1431 3745 1435 3749
rect 1583 3745 1587 3749
rect 2007 3744 2011 3748
rect 2047 3735 2051 3739
rect 2451 3739 2455 3743
rect 2635 3739 2639 3743
rect 2827 3739 2831 3743
rect 3011 3739 3015 3743
rect 3203 3739 3207 3743
rect 3395 3743 3399 3747
rect 3439 3743 3443 3747
rect 3787 3739 3791 3743
rect 2191 3732 2195 3736
rect 2375 3732 2379 3736
rect 2559 3732 2563 3736
rect 2743 3732 2747 3736
rect 2935 3732 2939 3736
rect 3127 3732 3131 3736
rect 3319 3732 3323 3736
rect 3511 3732 3515 3736
rect 3711 3732 3715 3736
rect 3943 3735 3947 3739
rect 2275 3711 2279 3715
rect 2451 3711 2455 3715
rect 2635 3711 2639 3715
rect 3439 3719 3443 3723
rect 3011 3711 3015 3715
rect 3203 3711 3207 3715
rect 3579 3707 3583 3711
rect 3731 3711 3735 3715
rect 2435 3691 2439 3695
rect 2667 3691 2671 3695
rect 2827 3691 2831 3695
rect 3143 3691 3147 3695
rect 3355 3691 3359 3695
rect 3787 3691 3791 3695
rect 111 3684 115 3688
rect 495 3683 499 3687
rect 591 3683 595 3687
rect 687 3683 691 3687
rect 791 3683 795 3687
rect 911 3683 915 3687
rect 1039 3683 1043 3687
rect 1183 3683 1187 3687
rect 1335 3683 1339 3687
rect 1495 3683 1499 3687
rect 1655 3683 1659 3687
rect 2007 3684 2011 3688
rect 3379 3683 3383 3687
rect 111 3667 115 3671
rect 571 3671 575 3675
rect 667 3671 671 3675
rect 763 3671 767 3675
rect 867 3671 871 3675
rect 903 3675 907 3679
rect 1115 3671 1119 3675
rect 1259 3671 1263 3675
rect 1267 3675 1271 3679
rect 1571 3675 1575 3679
rect 1615 3675 1619 3679
rect 495 3664 499 3668
rect 591 3664 595 3668
rect 687 3664 691 3668
rect 791 3664 795 3668
rect 911 3664 915 3668
rect 1039 3664 1043 3668
rect 1183 3664 1187 3668
rect 1335 3664 1339 3668
rect 1495 3664 1499 3668
rect 1655 3664 1659 3668
rect 2007 3667 2011 3671
rect 2047 3665 2051 3669
rect 2127 3668 2131 3672
rect 2351 3668 2355 3672
rect 2583 3668 2587 3672
rect 2815 3668 2819 3672
rect 3047 3668 3051 3672
rect 3279 3668 3283 3672
rect 3511 3668 3515 3672
rect 3751 3668 3755 3672
rect 3943 3665 3947 3669
rect 2203 3659 2207 3663
rect 2435 3659 2439 3663
rect 2667 3659 2671 3663
rect 3143 3659 3147 3663
rect 3355 3659 3359 3663
rect 3579 3659 3583 3663
rect 3827 3659 3831 3663
rect 571 3643 575 3647
rect 667 3643 671 3647
rect 763 3643 767 3647
rect 867 3643 871 3647
rect 1267 3651 1271 3655
rect 2047 3648 2051 3652
rect 2127 3649 2131 3653
rect 2351 3649 2355 3653
rect 2583 3649 2587 3653
rect 2815 3649 2819 3653
rect 3047 3649 3051 3653
rect 3279 3649 3283 3653
rect 3511 3649 3515 3653
rect 3751 3649 3755 3653
rect 3943 3648 3947 3652
rect 1219 3643 1223 3647
rect 1259 3643 1263 3647
rect 1615 3643 1619 3647
rect 859 3635 863 3639
rect 1691 3639 1695 3643
rect 411 3619 415 3623
rect 539 3619 543 3623
rect 835 3619 839 3623
rect 1115 3619 1119 3623
rect 1171 3619 1175 3623
rect 1515 3619 1519 3623
rect 1847 3619 1848 3623
rect 1848 3619 1851 3623
rect 739 3611 743 3615
rect 1759 3611 1763 3615
rect 111 3593 115 3597
rect 335 3596 339 3600
rect 463 3596 467 3600
rect 607 3596 611 3600
rect 759 3596 763 3600
rect 927 3596 931 3600
rect 1095 3596 1099 3600
rect 1263 3596 1267 3600
rect 1439 3596 1443 3600
rect 1615 3596 1619 3600
rect 1791 3596 1795 3600
rect 2007 3593 2011 3597
rect 411 3587 415 3591
rect 539 3587 543 3591
rect 835 3587 839 3591
rect 859 3587 863 3591
rect 1171 3587 1175 3591
rect 1339 3587 1343 3591
rect 1515 3587 1519 3591
rect 1691 3587 1695 3591
rect 1759 3587 1763 3591
rect 2047 3588 2051 3592
rect 2191 3587 2195 3591
rect 2327 3587 2331 3591
rect 2455 3587 2459 3591
rect 2583 3587 2587 3591
rect 2719 3587 2723 3591
rect 2855 3587 2859 3591
rect 2999 3587 3003 3591
rect 3143 3587 3147 3591
rect 3295 3587 3299 3591
rect 3455 3587 3459 3591
rect 3623 3587 3627 3591
rect 3943 3588 3947 3592
rect 111 3576 115 3580
rect 335 3577 339 3581
rect 463 3577 467 3581
rect 607 3577 611 3581
rect 759 3577 763 3581
rect 927 3577 931 3581
rect 1095 3577 1099 3581
rect 1263 3577 1267 3581
rect 1439 3577 1443 3581
rect 1615 3577 1619 3581
rect 1791 3577 1795 3581
rect 2007 3576 2011 3580
rect 2047 3571 2051 3575
rect 2279 3575 2283 3579
rect 2531 3575 2535 3579
rect 2659 3575 2663 3579
rect 2795 3575 2799 3579
rect 2931 3575 2935 3579
rect 3075 3575 3079 3579
rect 3219 3575 3223 3579
rect 3259 3579 3263 3583
rect 3379 3579 3383 3583
rect 3587 3579 3591 3583
rect 2191 3568 2195 3572
rect 2327 3568 2331 3572
rect 2455 3568 2459 3572
rect 2583 3568 2587 3572
rect 2719 3568 2723 3572
rect 2855 3568 2859 3572
rect 2999 3568 3003 3572
rect 3143 3568 3147 3572
rect 3295 3568 3299 3572
rect 3455 3568 3459 3572
rect 3623 3568 3627 3572
rect 3943 3571 3947 3575
rect 2203 3547 2207 3551
rect 2531 3547 2535 3551
rect 2659 3547 2663 3551
rect 2795 3547 2799 3551
rect 2931 3547 2935 3551
rect 3075 3547 3079 3551
rect 3219 3547 3223 3551
rect 3587 3547 3591 3551
rect 3259 3539 3263 3543
rect 3595 3543 3599 3547
rect 2279 3531 2283 3535
rect 2531 3531 2535 3535
rect 2779 3531 2783 3535
rect 3075 3531 3079 3535
rect 3399 3531 3403 3535
rect 3427 3531 3431 3535
rect 3771 3531 3775 3535
rect 3915 3531 3919 3535
rect 111 3512 115 3516
rect 159 3511 163 3515
rect 303 3511 307 3515
rect 463 3511 467 3515
rect 639 3511 643 3515
rect 815 3511 819 3515
rect 999 3511 1003 3515
rect 1175 3511 1179 3515
rect 1351 3511 1355 3515
rect 1527 3511 1531 3515
rect 1703 3511 1707 3515
rect 1879 3511 1883 3515
rect 2007 3512 2011 3516
rect 111 3495 115 3499
rect 235 3499 239 3503
rect 379 3499 383 3503
rect 539 3499 543 3503
rect 715 3499 719 3503
rect 739 3503 743 3507
rect 1075 3499 1079 3503
rect 1083 3503 1087 3507
rect 1663 3499 1667 3503
rect 1779 3499 1783 3503
rect 1847 3503 1851 3507
rect 2047 3505 2051 3509
rect 2103 3508 2107 3512
rect 2271 3508 2275 3512
rect 2447 3508 2451 3512
rect 2631 3508 2635 3512
rect 2815 3508 2819 3512
rect 2999 3508 3003 3512
rect 3175 3508 3179 3512
rect 3351 3508 3355 3512
rect 3519 3508 3523 3512
rect 3687 3508 3691 3512
rect 3839 3508 3843 3512
rect 3943 3505 3947 3509
rect 159 3492 163 3496
rect 303 3492 307 3496
rect 463 3492 467 3496
rect 639 3492 643 3496
rect 815 3492 819 3496
rect 999 3492 1003 3496
rect 1175 3492 1179 3496
rect 1351 3492 1355 3496
rect 1527 3492 1531 3496
rect 1703 3492 1707 3496
rect 1879 3492 1883 3496
rect 2007 3495 2011 3499
rect 2179 3499 2183 3503
rect 2531 3499 2535 3503
rect 3075 3499 3079 3503
rect 3251 3499 3255 3503
rect 3427 3499 3431 3503
rect 3595 3499 3599 3503
rect 3771 3499 3775 3503
rect 2047 3488 2051 3492
rect 2103 3489 2107 3493
rect 2271 3489 2275 3493
rect 2447 3489 2451 3493
rect 2631 3489 2635 3493
rect 2815 3489 2819 3493
rect 2999 3489 3003 3493
rect 3175 3489 3179 3493
rect 3351 3489 3355 3493
rect 3519 3489 3523 3493
rect 3687 3489 3691 3493
rect 3839 3489 3843 3493
rect 3943 3488 3947 3492
rect 235 3475 239 3479
rect 379 3471 383 3475
rect 539 3471 543 3475
rect 715 3471 719 3475
rect 1083 3471 1087 3475
rect 1339 3471 1343 3475
rect 679 3463 683 3467
rect 1603 3467 1607 3471
rect 1663 3471 1667 3475
rect 1779 3471 1783 3475
rect 255 3447 259 3451
rect 263 3447 267 3451
rect 395 3447 399 3451
rect 611 3447 615 3451
rect 1075 3447 1079 3451
rect 1083 3447 1087 3451
rect 1235 3447 1239 3451
rect 1619 3447 1623 3451
rect 1803 3447 1807 3451
rect 1947 3447 1951 3451
rect 2047 3432 2051 3436
rect 2127 3431 2131 3435
rect 2311 3431 2315 3435
rect 2495 3431 2499 3435
rect 2679 3431 2683 3435
rect 2863 3431 2867 3435
rect 3047 3431 3051 3435
rect 3223 3431 3227 3435
rect 3407 3431 3411 3435
rect 3591 3431 3595 3435
rect 3775 3431 3779 3435
rect 3943 3432 3947 3436
rect 111 3421 115 3425
rect 135 3424 139 3428
rect 319 3424 323 3428
rect 535 3424 539 3428
rect 751 3424 755 3428
rect 959 3424 963 3428
rect 1159 3424 1163 3428
rect 1351 3424 1355 3428
rect 1535 3424 1539 3428
rect 1719 3424 1723 3428
rect 1903 3424 1907 3428
rect 2007 3421 2011 3425
rect 263 3415 267 3419
rect 395 3415 399 3419
rect 611 3415 615 3419
rect 679 3415 683 3419
rect 1083 3415 1087 3419
rect 1235 3415 1239 3419
rect 1427 3415 1431 3419
rect 1603 3415 1607 3419
rect 1619 3415 1623 3419
rect 1803 3415 1807 3419
rect 2047 3415 2051 3419
rect 2203 3419 2207 3423
rect 2387 3419 2391 3423
rect 2571 3419 2575 3423
rect 2779 3423 2783 3427
rect 2947 3419 2951 3423
rect 3175 3423 3179 3427
rect 3399 3423 3403 3427
rect 3547 3423 3551 3427
rect 3851 3419 3855 3423
rect 2127 3412 2131 3416
rect 2311 3412 2315 3416
rect 2495 3412 2499 3416
rect 2679 3412 2683 3416
rect 2863 3412 2867 3416
rect 3047 3412 3051 3416
rect 3223 3412 3227 3416
rect 3407 3412 3411 3416
rect 3591 3412 3595 3416
rect 3775 3412 3779 3416
rect 3943 3415 3947 3419
rect 111 3404 115 3408
rect 135 3405 139 3409
rect 319 3405 323 3409
rect 535 3405 539 3409
rect 751 3405 755 3409
rect 959 3405 963 3409
rect 1159 3405 1163 3409
rect 1351 3405 1355 3409
rect 1535 3405 1539 3409
rect 1719 3405 1723 3409
rect 1903 3405 1907 3409
rect 2007 3404 2011 3408
rect 2179 3391 2180 3395
rect 2180 3391 2183 3395
rect 2387 3391 2391 3395
rect 2571 3391 2575 3395
rect 3175 3391 3179 3395
rect 3251 3391 3255 3395
rect 3547 3391 3551 3395
rect 3659 3387 3663 3391
rect 3827 3391 3828 3395
rect 3828 3391 3831 3395
rect 2155 3359 2159 3363
rect 2203 3359 2207 3363
rect 2443 3359 2447 3363
rect 2595 3359 2599 3363
rect 2775 3359 2779 3363
rect 2871 3359 2875 3363
rect 2947 3359 2951 3363
rect 3011 3359 3015 3363
rect 3155 3359 3159 3363
rect 3499 3359 3503 3363
rect 3507 3359 3511 3363
rect 3611 3359 3615 3363
rect 3907 3359 3911 3363
rect 111 3352 115 3356
rect 135 3351 139 3355
rect 231 3351 235 3355
rect 375 3351 379 3355
rect 535 3351 539 3355
rect 703 3351 707 3355
rect 871 3351 875 3355
rect 1047 3351 1051 3355
rect 1215 3351 1219 3355
rect 1383 3351 1387 3355
rect 1543 3351 1547 3355
rect 1703 3351 1707 3355
rect 1871 3351 1875 3355
rect 2007 3352 2011 3356
rect 111 3335 115 3339
rect 211 3339 215 3343
rect 307 3339 311 3343
rect 451 3339 455 3343
rect 611 3339 615 3343
rect 779 3339 783 3343
rect 799 3343 803 3347
rect 1123 3339 1127 3343
rect 1167 3343 1171 3347
rect 1343 3343 1347 3347
rect 1619 3339 1623 3343
rect 1779 3339 1783 3343
rect 1947 3343 1951 3347
rect 135 3332 139 3336
rect 231 3332 235 3336
rect 375 3332 379 3336
rect 535 3332 539 3336
rect 703 3332 707 3336
rect 871 3332 875 3336
rect 1047 3332 1051 3336
rect 1215 3332 1219 3336
rect 1383 3332 1387 3336
rect 1543 3332 1547 3336
rect 1703 3332 1707 3336
rect 1871 3332 1875 3336
rect 2007 3335 2011 3339
rect 2047 3333 2051 3337
rect 2071 3336 2075 3340
rect 2215 3336 2219 3340
rect 2359 3336 2363 3340
rect 2511 3336 2515 3340
rect 2655 3336 2659 3340
rect 2799 3336 2803 3340
rect 2935 3336 2939 3340
rect 3079 3336 3083 3340
rect 3223 3336 3227 3340
rect 3375 3336 3379 3340
rect 3535 3336 3539 3340
rect 3695 3336 3699 3340
rect 3839 3336 3843 3340
rect 3943 3333 3947 3337
rect 2147 3327 2151 3331
rect 2155 3327 2159 3331
rect 2443 3327 2447 3331
rect 2595 3327 2599 3331
rect 2775 3327 2779 3331
rect 3011 3327 3015 3331
rect 3155 3327 3159 3331
rect 3299 3327 3303 3331
rect 3507 3327 3511 3331
rect 3611 3327 3615 3331
rect 3659 3327 3663 3331
rect 3915 3327 3919 3331
rect 2047 3316 2051 3320
rect 2071 3317 2075 3321
rect 2215 3317 2219 3321
rect 2359 3317 2363 3321
rect 2511 3317 2515 3321
rect 2655 3317 2659 3321
rect 2799 3317 2803 3321
rect 2935 3317 2939 3321
rect 3079 3317 3083 3321
rect 3223 3317 3227 3321
rect 3375 3317 3379 3321
rect 3535 3317 3539 3321
rect 3695 3317 3699 3321
rect 3839 3317 3843 3321
rect 3943 3316 3947 3320
rect 203 3307 207 3311
rect 211 3311 215 3315
rect 307 3311 311 3315
rect 451 3311 455 3315
rect 611 3311 615 3315
rect 779 3311 783 3315
rect 1167 3311 1171 3315
rect 1343 3311 1347 3315
rect 1427 3311 1431 3315
rect 1595 3307 1596 3311
rect 1596 3307 1599 3311
rect 1619 3311 1623 3315
rect 1779 3311 1783 3315
rect 255 3295 259 3299
rect 519 3295 520 3299
rect 520 3295 523 3299
rect 739 3295 743 3299
rect 1123 3295 1127 3299
rect 1155 3295 1159 3299
rect 1603 3295 1607 3299
rect 1771 3295 1775 3299
rect 799 3283 803 3287
rect 111 3269 115 3273
rect 135 3272 139 3276
rect 279 3272 283 3276
rect 463 3272 467 3276
rect 663 3272 667 3276
rect 871 3272 875 3276
rect 1079 3272 1083 3276
rect 1295 3272 1299 3276
rect 1519 3272 1523 3276
rect 1743 3272 1747 3276
rect 2007 3269 2011 3273
rect 203 3263 207 3267
rect 255 3263 259 3267
rect 739 3263 743 3267
rect 799 3263 803 3267
rect 1155 3263 1159 3267
rect 1371 3263 1375 3267
rect 1595 3263 1599 3267
rect 1603 3263 1607 3267
rect 111 3252 115 3256
rect 135 3253 139 3257
rect 279 3253 283 3257
rect 463 3253 467 3257
rect 663 3253 667 3257
rect 871 3253 875 3257
rect 1079 3253 1083 3257
rect 1295 3253 1299 3257
rect 1519 3253 1523 3257
rect 1743 3253 1747 3257
rect 2007 3252 2011 3256
rect 2047 3256 2051 3260
rect 2111 3255 2115 3259
rect 2247 3255 2251 3259
rect 2399 3255 2403 3259
rect 2575 3255 2579 3259
rect 2783 3255 2787 3259
rect 2871 3251 2875 3255
rect 3015 3255 3019 3259
rect 3263 3255 3267 3259
rect 3527 3255 3531 3259
rect 3791 3255 3795 3259
rect 3943 3256 3947 3260
rect 2047 3239 2051 3243
rect 2187 3243 2191 3247
rect 2475 3243 2479 3247
rect 2651 3243 2655 3247
rect 2859 3243 2863 3247
rect 3339 3243 3343 3247
rect 3499 3247 3503 3251
rect 3867 3243 3871 3247
rect 2111 3236 2115 3240
rect 2247 3236 2251 3240
rect 2399 3236 2403 3240
rect 2575 3236 2579 3240
rect 2783 3236 2787 3240
rect 3015 3236 3019 3240
rect 3263 3236 3267 3240
rect 3527 3236 3531 3240
rect 3791 3236 3795 3240
rect 3943 3239 3947 3243
rect 2147 3215 2151 3219
rect 2331 3211 2335 3215
rect 2475 3215 2479 3219
rect 2651 3215 2655 3219
rect 2859 3215 2863 3219
rect 3311 3211 3315 3215
rect 3507 3215 3511 3219
rect 3847 3215 3848 3219
rect 3848 3215 3851 3219
rect 111 3200 115 3204
rect 135 3199 139 3203
rect 287 3199 291 3203
rect 447 3199 451 3203
rect 615 3199 619 3203
rect 791 3199 795 3203
rect 967 3199 971 3203
rect 1143 3199 1147 3203
rect 1327 3199 1331 3203
rect 1511 3199 1515 3203
rect 1695 3199 1699 3203
rect 2007 3200 2011 3204
rect 2187 3199 2191 3203
rect 2347 3199 2351 3203
rect 2443 3199 2447 3203
rect 2539 3199 2543 3203
rect 2635 3199 2639 3203
rect 2731 3199 2735 3203
rect 2827 3199 2831 3203
rect 2923 3199 2927 3203
rect 3023 3199 3027 3203
rect 3115 3199 3119 3203
rect 3211 3199 3215 3203
rect 3339 3199 3343 3203
rect 3403 3199 3407 3203
rect 3587 3199 3591 3203
rect 3651 3199 3655 3203
rect 3915 3199 3919 3203
rect 111 3183 115 3187
rect 259 3187 263 3191
rect 363 3187 367 3191
rect 523 3191 527 3195
rect 559 3191 563 3195
rect 751 3191 755 3195
rect 1043 3187 1047 3191
rect 1091 3191 1095 3195
rect 1587 3187 1591 3191
rect 1771 3191 1775 3195
rect 2147 3191 2151 3195
rect 3659 3191 3663 3195
rect 135 3180 139 3184
rect 287 3180 291 3184
rect 447 3180 451 3184
rect 615 3180 619 3184
rect 791 3180 795 3184
rect 967 3180 971 3184
rect 1143 3180 1147 3184
rect 1327 3180 1331 3184
rect 1511 3180 1515 3184
rect 1695 3180 1699 3184
rect 2007 3183 2011 3187
rect 2047 3173 2051 3177
rect 2071 3176 2075 3180
rect 2167 3176 2171 3180
rect 2263 3176 2267 3180
rect 2359 3176 2363 3180
rect 2455 3176 2459 3180
rect 2551 3176 2555 3180
rect 2647 3176 2651 3180
rect 2743 3176 2747 3180
rect 2839 3176 2843 3180
rect 2935 3176 2939 3180
rect 3031 3176 3035 3180
rect 3127 3176 3131 3180
rect 3223 3176 3227 3180
rect 3319 3176 3323 3180
rect 3439 3176 3443 3180
rect 3575 3176 3579 3180
rect 3719 3176 3723 3180
rect 3839 3176 3843 3180
rect 3943 3173 3947 3177
rect 559 3167 563 3171
rect 2147 3167 2151 3171
rect 259 3155 263 3159
rect 363 3159 367 3163
rect 751 3159 755 3163
rect 1091 3159 1095 3163
rect 1371 3159 1375 3163
rect 1467 3155 1471 3159
rect 1587 3159 1591 3163
rect 2047 3156 2051 3160
rect 2071 3157 2075 3161
rect 2167 3157 2171 3161
rect 2331 3167 2335 3171
rect 2347 3167 2351 3171
rect 2443 3167 2447 3171
rect 2539 3167 2543 3171
rect 2635 3167 2639 3171
rect 2731 3167 2735 3171
rect 2827 3167 2831 3171
rect 2923 3167 2927 3171
rect 3023 3167 3027 3171
rect 3115 3167 3119 3171
rect 3211 3167 3215 3171
rect 3311 3167 3315 3171
rect 3403 3167 3407 3171
rect 3651 3167 3655 3171
rect 3659 3167 3663 3171
rect 3907 3167 3911 3171
rect 2263 3157 2267 3161
rect 2359 3157 2363 3161
rect 2455 3157 2459 3161
rect 2551 3157 2555 3161
rect 2647 3157 2651 3161
rect 2743 3157 2747 3161
rect 2839 3157 2843 3161
rect 2935 3157 2939 3161
rect 3031 3157 3035 3161
rect 3127 3157 3131 3161
rect 3223 3157 3227 3161
rect 3319 3157 3323 3161
rect 3439 3157 3443 3161
rect 3575 3157 3579 3161
rect 3719 3157 3723 3161
rect 3839 3157 3843 3161
rect 3943 3156 3947 3160
rect 2299 3151 2303 3155
rect 367 3139 368 3143
rect 368 3139 371 3143
rect 387 3139 391 3143
rect 515 3139 519 3143
rect 659 3139 663 3143
rect 819 3139 823 3143
rect 1043 3139 1047 3143
rect 1475 3139 1479 3143
rect 1643 3139 1647 3143
rect 1795 3139 1799 3143
rect 111 3113 115 3117
rect 311 3116 315 3120
rect 439 3116 443 3120
rect 583 3116 587 3120
rect 743 3116 747 3120
rect 903 3116 907 3120
rect 1063 3116 1067 3120
rect 1223 3116 1227 3120
rect 1391 3116 1395 3120
rect 1559 3116 1563 3120
rect 1727 3116 1731 3120
rect 2007 3113 2011 3117
rect 387 3107 391 3111
rect 515 3107 519 3111
rect 659 3107 663 3111
rect 819 3107 823 3111
rect 1351 3107 1355 3111
rect 1467 3107 1471 3111
rect 1475 3107 1479 3111
rect 1643 3107 1647 3111
rect 111 3096 115 3100
rect 311 3097 315 3101
rect 439 3097 443 3101
rect 583 3097 587 3101
rect 743 3097 747 3101
rect 903 3097 907 3101
rect 1063 3097 1067 3101
rect 1223 3097 1227 3101
rect 1391 3097 1395 3101
rect 1559 3097 1563 3101
rect 1727 3097 1731 3101
rect 2007 3096 2011 3100
rect 2047 3092 2051 3096
rect 2071 3091 2075 3095
rect 2335 3091 2339 3095
rect 2623 3091 2627 3095
rect 2911 3091 2915 3095
rect 3207 3091 3211 3095
rect 3503 3091 3507 3095
rect 3799 3091 3803 3095
rect 3943 3092 3947 3096
rect 2047 3075 2051 3079
rect 2147 3079 2151 3083
rect 2183 3083 2187 3087
rect 2699 3079 2703 3083
rect 2987 3079 2991 3083
rect 3283 3079 3287 3083
rect 3587 3083 3591 3087
rect 3875 3079 3879 3083
rect 2071 3072 2075 3076
rect 2335 3072 2339 3076
rect 2623 3072 2627 3076
rect 2911 3072 2915 3076
rect 3207 3072 3211 3076
rect 3503 3072 3507 3076
rect 3799 3072 3803 3076
rect 3943 3075 3947 3079
rect 2183 3051 2187 3055
rect 2299 3051 2303 3055
rect 2675 3047 2676 3051
rect 2676 3047 2679 3051
rect 2699 3051 2703 3055
rect 2987 3051 2991 3055
rect 3283 3051 3287 3055
rect 3867 3051 3871 3055
rect 111 3036 115 3040
rect 503 3035 507 3039
rect 599 3035 603 3039
rect 703 3035 707 3039
rect 815 3035 819 3039
rect 935 3035 939 3039
rect 1071 3035 1075 3039
rect 1223 3035 1227 3039
rect 1383 3035 1387 3039
rect 1551 3035 1555 3039
rect 1719 3035 1723 3039
rect 2007 3036 2011 3040
rect 2147 3035 2151 3039
rect 2959 3035 2963 3039
rect 3259 3035 3263 3039
rect 3371 3035 3375 3039
rect 3923 3035 3927 3039
rect 367 3027 371 3031
rect 587 3027 591 3031
rect 683 3027 687 3031
rect 807 3027 811 3031
rect 903 3027 907 3031
rect 111 3019 115 3023
rect 1147 3023 1151 3027
rect 1343 3027 1347 3031
rect 1627 3023 1631 3027
rect 1795 3027 1799 3031
rect 503 3016 507 3020
rect 599 3016 603 3020
rect 703 3016 707 3020
rect 815 3016 819 3020
rect 935 3016 939 3020
rect 1071 3016 1075 3020
rect 1223 3016 1227 3020
rect 1383 3016 1387 3020
rect 1551 3016 1555 3020
rect 1719 3016 1723 3020
rect 2007 3019 2011 3023
rect 2047 3009 2051 3013
rect 2071 3012 2075 3016
rect 2383 3012 2387 3016
rect 2703 3012 2707 3016
rect 2999 3012 3003 3016
rect 3287 3012 3291 3016
rect 3575 3012 3579 3016
rect 3839 3012 3843 3016
rect 3943 3009 3947 3013
rect 2451 3003 2455 3007
rect 2675 3003 2679 3007
rect 2959 3003 2963 3007
rect 3259 3003 3263 3007
rect 3371 3003 3375 3007
rect 3915 3003 3919 3007
rect 587 2995 591 2999
rect 683 2995 687 2999
rect 807 2995 811 2999
rect 903 2995 907 2999
rect 991 2991 992 2995
rect 992 2991 995 2995
rect 1343 2995 1347 2999
rect 1351 2995 1355 2999
rect 1563 2991 1567 2995
rect 1627 2995 1631 2999
rect 2047 2992 2051 2996
rect 2071 2993 2075 2997
rect 2383 2993 2387 2997
rect 2703 2993 2707 2997
rect 2999 2993 3003 2997
rect 3287 2993 3291 2997
rect 3575 2993 3579 2997
rect 3839 2993 3843 2997
rect 3943 2992 3947 2996
rect 627 2975 631 2979
rect 723 2975 727 2979
rect 835 2975 839 2979
rect 963 2975 967 2979
rect 1147 2975 1151 2979
rect 1251 2975 1255 2979
rect 1571 2975 1575 2979
rect 1739 2975 1743 2979
rect 1923 2975 1927 2979
rect 923 2967 927 2971
rect 111 2949 115 2953
rect 551 2952 555 2956
rect 647 2952 651 2956
rect 759 2952 763 2956
rect 887 2952 891 2956
rect 1023 2952 1027 2956
rect 1175 2952 1179 2956
rect 1327 2952 1331 2956
rect 1487 2952 1491 2956
rect 1655 2952 1659 2956
rect 1823 2952 1827 2956
rect 2007 2949 2011 2953
rect 627 2943 631 2947
rect 723 2943 727 2947
rect 835 2943 839 2947
rect 963 2943 967 2947
rect 991 2943 995 2947
rect 1251 2943 1255 2947
rect 1563 2943 1567 2947
rect 1571 2943 1575 2947
rect 1739 2943 1743 2947
rect 111 2932 115 2936
rect 551 2933 555 2937
rect 647 2933 651 2937
rect 759 2933 763 2937
rect 887 2933 891 2937
rect 1023 2933 1027 2937
rect 1175 2933 1179 2937
rect 1327 2933 1331 2937
rect 1487 2933 1491 2937
rect 1655 2933 1659 2937
rect 1823 2933 1827 2937
rect 2007 2932 2011 2936
rect 2047 2936 2051 2940
rect 2071 2935 2075 2939
rect 2391 2935 2395 2939
rect 2703 2935 2707 2939
rect 2975 2935 2979 2939
rect 3215 2935 3219 2939
rect 3439 2935 3443 2939
rect 3647 2935 3651 2939
rect 3839 2935 3843 2939
rect 3943 2936 3947 2940
rect 2047 2919 2051 2923
rect 2147 2923 2151 2927
rect 2779 2923 2783 2927
rect 3051 2923 3055 2927
rect 3291 2923 3295 2927
rect 3515 2923 3519 2927
rect 3723 2923 3727 2927
rect 2071 2916 2075 2920
rect 2391 2916 2395 2920
rect 2703 2916 2707 2920
rect 2975 2916 2979 2920
rect 3215 2916 3219 2920
rect 3439 2916 3443 2920
rect 3647 2916 3651 2920
rect 3839 2916 3843 2920
rect 3943 2919 3947 2923
rect 2447 2895 2448 2899
rect 2448 2895 2451 2899
rect 3619 2903 3623 2907
rect 2779 2887 2783 2891
rect 3051 2895 3055 2899
rect 3291 2895 3295 2899
rect 3515 2895 3519 2899
rect 3723 2895 3727 2899
rect 2147 2879 2151 2883
rect 2231 2879 2235 2883
rect 2371 2879 2375 2883
rect 2611 2879 2615 2883
rect 3067 2879 3071 2883
rect 3291 2879 3295 2883
rect 3507 2879 3511 2883
rect 3907 2879 3911 2883
rect 111 2872 115 2876
rect 471 2871 475 2875
rect 575 2871 579 2875
rect 695 2871 699 2875
rect 839 2871 843 2875
rect 991 2871 995 2875
rect 1151 2871 1155 2875
rect 1319 2871 1323 2875
rect 1495 2871 1499 2875
rect 1671 2871 1675 2875
rect 1847 2871 1851 2875
rect 2007 2872 2011 2876
rect 3439 2871 3443 2875
rect 111 2855 115 2859
rect 567 2859 571 2863
rect 651 2859 655 2863
rect 771 2859 775 2863
rect 915 2859 919 2863
rect 923 2863 927 2867
rect 1227 2859 1231 2863
rect 1395 2859 1399 2863
rect 1631 2859 1635 2863
rect 1747 2859 1751 2863
rect 1923 2863 1927 2867
rect 471 2852 475 2856
rect 575 2852 579 2856
rect 695 2852 699 2856
rect 839 2852 843 2856
rect 991 2852 995 2856
rect 1151 2852 1155 2856
rect 1319 2852 1323 2856
rect 1495 2852 1499 2856
rect 1671 2852 1675 2856
rect 1847 2852 1851 2856
rect 2007 2855 2011 2859
rect 2047 2853 2051 2857
rect 2071 2856 2075 2860
rect 2295 2856 2299 2860
rect 2535 2856 2539 2860
rect 2767 2856 2771 2860
rect 2991 2856 2995 2860
rect 3215 2856 3219 2860
rect 3431 2856 3435 2860
rect 3647 2856 3651 2860
rect 3839 2856 3843 2860
rect 3943 2853 3947 2857
rect 2231 2847 2235 2851
rect 2371 2847 2375 2851
rect 2611 2847 2615 2851
rect 2719 2847 2723 2851
rect 3067 2847 3071 2851
rect 3291 2847 3295 2851
rect 3507 2847 3511 2851
rect 3619 2847 3623 2851
rect 3923 2847 3927 2851
rect 547 2827 551 2831
rect 567 2831 571 2835
rect 651 2831 655 2835
rect 771 2831 775 2835
rect 915 2831 919 2835
rect 2047 2836 2051 2840
rect 2071 2837 2075 2841
rect 2295 2837 2299 2841
rect 2535 2837 2539 2841
rect 2767 2837 2771 2841
rect 2991 2837 2995 2841
rect 3215 2837 3219 2841
rect 3431 2837 3435 2841
rect 3647 2837 3651 2841
rect 3839 2837 3843 2841
rect 3943 2836 3947 2840
rect 1227 2831 1231 2835
rect 1551 2827 1552 2831
rect 1552 2827 1555 2831
rect 1631 2831 1635 2835
rect 1747 2831 1751 2835
rect 563 2811 567 2815
rect 659 2811 663 2815
rect 763 2811 767 2815
rect 883 2811 887 2815
rect 999 2811 1003 2815
rect 1191 2811 1195 2815
rect 1327 2811 1331 2815
rect 1395 2811 1399 2815
rect 1683 2811 1687 2815
rect 1859 2811 1863 2815
rect 111 2785 115 2789
rect 479 2788 483 2792
rect 575 2788 579 2792
rect 679 2788 683 2792
rect 799 2788 803 2792
rect 935 2788 939 2792
rect 1079 2788 1083 2792
rect 1239 2788 1243 2792
rect 1415 2788 1419 2792
rect 1599 2788 1603 2792
rect 1783 2788 1787 2792
rect 2007 2785 2011 2789
rect 547 2779 551 2783
rect 563 2779 567 2783
rect 659 2779 663 2783
rect 763 2779 767 2783
rect 883 2779 887 2783
rect 1151 2779 1155 2783
rect 1191 2779 1195 2783
rect 1327 2779 1331 2783
rect 1551 2779 1555 2783
rect 1683 2779 1687 2783
rect 2047 2780 2051 2784
rect 2071 2779 2075 2783
rect 2199 2779 2203 2783
rect 2367 2779 2371 2783
rect 2551 2779 2555 2783
rect 2735 2779 2739 2783
rect 2927 2779 2931 2783
rect 3111 2779 3115 2783
rect 3295 2779 3299 2783
rect 3479 2779 3483 2783
rect 3671 2779 3675 2783
rect 3839 2779 3843 2783
rect 3943 2780 3947 2784
rect 111 2768 115 2772
rect 479 2769 483 2773
rect 575 2769 579 2773
rect 679 2769 683 2773
rect 799 2769 803 2773
rect 935 2769 939 2773
rect 1079 2769 1083 2773
rect 1239 2769 1243 2773
rect 1415 2769 1419 2773
rect 1599 2769 1603 2773
rect 1783 2769 1787 2773
rect 2007 2768 2011 2772
rect 2047 2763 2051 2767
rect 2147 2767 2151 2771
rect 2275 2767 2279 2771
rect 2443 2767 2447 2771
rect 2627 2767 2631 2771
rect 2659 2771 2663 2775
rect 3003 2767 3007 2771
rect 3187 2767 3191 2771
rect 3371 2767 3375 2771
rect 3439 2771 3443 2775
rect 3907 2775 3911 2779
rect 3747 2767 3751 2771
rect 2071 2760 2075 2764
rect 2199 2760 2203 2764
rect 2367 2760 2371 2764
rect 2551 2760 2555 2764
rect 2735 2760 2739 2764
rect 2927 2760 2931 2764
rect 3111 2760 3115 2764
rect 3295 2760 3299 2764
rect 3479 2760 3483 2764
rect 3671 2760 3675 2764
rect 3839 2760 3843 2764
rect 3943 2763 3947 2767
rect 2719 2747 2723 2751
rect 2147 2739 2151 2743
rect 2275 2739 2279 2743
rect 2443 2739 2447 2743
rect 2627 2739 2631 2743
rect 3003 2739 3007 2743
rect 3187 2739 3191 2743
rect 3371 2739 3375 2743
rect 3875 2739 3879 2743
rect 2659 2727 2663 2731
rect 3379 2731 3383 2735
rect 3907 2735 3911 2739
rect 2147 2719 2151 2723
rect 2267 2719 2271 2723
rect 2395 2719 2399 2723
rect 2523 2719 2527 2723
rect 2783 2719 2784 2723
rect 2784 2719 2787 2723
rect 2803 2719 2807 2723
rect 2963 2719 2967 2723
rect 3139 2719 3143 2723
rect 3331 2719 3335 2723
rect 3747 2719 3751 2723
rect 111 2712 115 2716
rect 511 2711 515 2715
rect 623 2711 627 2715
rect 743 2711 747 2715
rect 879 2711 883 2715
rect 1015 2711 1019 2715
rect 1159 2711 1163 2715
rect 1311 2711 1315 2715
rect 1463 2711 1467 2715
rect 1623 2711 1627 2715
rect 1783 2711 1787 2715
rect 2007 2712 2011 2716
rect 111 2695 115 2699
rect 587 2699 591 2703
rect 699 2699 703 2703
rect 819 2699 823 2703
rect 955 2699 959 2703
rect 999 2703 1003 2707
rect 1235 2699 1239 2703
rect 1387 2699 1391 2703
rect 1539 2699 1543 2703
rect 1699 2699 1703 2703
rect 1859 2703 1863 2707
rect 511 2692 515 2696
rect 623 2692 627 2696
rect 743 2692 747 2696
rect 879 2692 883 2696
rect 1015 2692 1019 2696
rect 1159 2692 1163 2696
rect 1311 2692 1315 2696
rect 1463 2692 1467 2696
rect 1623 2692 1627 2696
rect 1783 2692 1787 2696
rect 2007 2695 2011 2699
rect 2047 2693 2051 2697
rect 2071 2696 2075 2700
rect 2191 2696 2195 2700
rect 2319 2696 2323 2700
rect 2447 2696 2451 2700
rect 2583 2696 2587 2700
rect 2727 2696 2731 2700
rect 2887 2696 2891 2700
rect 3063 2696 3067 2700
rect 3255 2696 3259 2700
rect 3455 2696 3459 2700
rect 3655 2696 3659 2700
rect 3839 2696 3843 2700
rect 3943 2693 3947 2697
rect 2147 2687 2151 2691
rect 2267 2687 2271 2691
rect 2395 2687 2399 2691
rect 2523 2687 2527 2691
rect 2539 2687 2543 2691
rect 2803 2687 2807 2691
rect 2963 2687 2967 2691
rect 3139 2687 3143 2691
rect 3331 2687 3335 2691
rect 3379 2687 3383 2691
rect 3907 2687 3911 2691
rect 2047 2676 2051 2680
rect 2071 2677 2075 2681
rect 2191 2677 2195 2681
rect 2319 2677 2323 2681
rect 2447 2677 2451 2681
rect 2583 2677 2587 2681
rect 2727 2677 2731 2681
rect 2887 2677 2891 2681
rect 3063 2677 3067 2681
rect 3255 2677 3259 2681
rect 3455 2677 3459 2681
rect 3655 2677 3659 2681
rect 3839 2677 3843 2681
rect 3943 2676 3947 2680
rect 587 2671 591 2675
rect 699 2671 703 2675
rect 819 2671 823 2675
rect 955 2671 959 2675
rect 1151 2671 1155 2675
rect 1235 2671 1239 2675
rect 859 2663 863 2667
rect 1507 2667 1511 2671
rect 1539 2671 1543 2675
rect 1699 2671 1703 2675
rect 443 2651 447 2655
rect 563 2651 567 2655
rect 691 2651 695 2655
rect 827 2651 831 2655
rect 1251 2651 1255 2655
rect 1387 2651 1391 2655
rect 1515 2651 1519 2655
rect 1651 2651 1655 2655
rect 1803 2651 1807 2655
rect 739 2643 743 2647
rect 111 2625 115 2629
rect 367 2628 371 2632
rect 487 2628 491 2632
rect 615 2628 619 2632
rect 751 2628 755 2632
rect 895 2628 899 2632
rect 1031 2628 1035 2632
rect 1167 2628 1171 2632
rect 1303 2628 1307 2632
rect 1431 2628 1435 2632
rect 1567 2628 1571 2632
rect 1703 2628 1707 2632
rect 2007 2625 2011 2629
rect 443 2619 447 2623
rect 563 2619 567 2623
rect 691 2619 695 2623
rect 827 2619 831 2623
rect 859 2619 863 2623
rect 979 2619 983 2623
rect 1251 2619 1255 2623
rect 1507 2619 1511 2623
rect 1515 2619 1519 2623
rect 1651 2619 1655 2623
rect 2047 2616 2051 2620
rect 2231 2615 2235 2619
rect 2335 2615 2339 2619
rect 2447 2615 2451 2619
rect 2559 2615 2563 2619
rect 2671 2615 2675 2619
rect 2791 2615 2795 2619
rect 2911 2615 2915 2619
rect 3031 2615 3035 2619
rect 3151 2615 3155 2619
rect 3943 2616 3947 2620
rect 111 2608 115 2612
rect 367 2609 371 2613
rect 487 2609 491 2613
rect 615 2609 619 2613
rect 751 2609 755 2613
rect 895 2609 899 2613
rect 1031 2609 1035 2613
rect 1167 2609 1171 2613
rect 1303 2609 1307 2613
rect 1431 2609 1435 2613
rect 1567 2609 1571 2613
rect 1703 2609 1707 2613
rect 2007 2608 2011 2612
rect 2047 2599 2051 2603
rect 2307 2603 2311 2607
rect 2411 2603 2415 2607
rect 2523 2603 2527 2607
rect 2635 2603 2639 2607
rect 2643 2607 2647 2611
rect 2783 2607 2787 2611
rect 3107 2603 3111 2607
rect 3115 2607 3119 2611
rect 2231 2596 2235 2600
rect 2335 2596 2339 2600
rect 2447 2596 2451 2600
rect 2559 2596 2563 2600
rect 2671 2596 2675 2600
rect 2791 2596 2795 2600
rect 2911 2596 2915 2600
rect 3031 2596 3035 2600
rect 3151 2596 3155 2600
rect 3943 2599 3947 2603
rect 2539 2583 2543 2587
rect 2307 2575 2311 2579
rect 2411 2575 2415 2579
rect 2523 2575 2527 2579
rect 2635 2575 2639 2579
rect 3115 2583 3119 2587
rect 3067 2571 3071 2575
rect 3107 2575 3111 2579
rect 2643 2563 2647 2567
rect 111 2556 115 2560
rect 135 2555 139 2559
rect 287 2555 291 2559
rect 447 2555 451 2559
rect 607 2555 611 2559
rect 767 2555 771 2559
rect 919 2555 923 2559
rect 1063 2555 1067 2559
rect 1199 2555 1203 2559
rect 1335 2555 1339 2559
rect 1463 2555 1467 2559
rect 1591 2555 1595 2559
rect 1727 2555 1731 2559
rect 2007 2556 2011 2560
rect 2459 2555 2463 2559
rect 2571 2555 2575 2559
rect 2691 2555 2695 2559
rect 2819 2555 2823 2559
rect 3075 2555 3079 2559
rect 3195 2555 3199 2559
rect 3315 2555 3319 2559
rect 3443 2555 3447 2559
rect 111 2539 115 2543
rect 211 2543 215 2547
rect 363 2543 367 2547
rect 523 2543 527 2547
rect 683 2543 687 2547
rect 739 2547 743 2551
rect 995 2543 999 2547
rect 1139 2543 1143 2547
rect 1275 2543 1279 2547
rect 1411 2543 1415 2547
rect 1539 2543 1543 2547
rect 1667 2543 1671 2547
rect 1803 2547 1807 2551
rect 3435 2547 3439 2551
rect 135 2536 139 2540
rect 287 2536 291 2540
rect 447 2536 451 2540
rect 607 2536 611 2540
rect 767 2536 771 2540
rect 919 2536 923 2540
rect 1063 2536 1067 2540
rect 1199 2536 1203 2540
rect 1335 2536 1339 2540
rect 1463 2536 1467 2540
rect 1591 2536 1595 2540
rect 1727 2536 1731 2540
rect 2007 2539 2011 2543
rect 2047 2529 2051 2533
rect 2383 2532 2387 2536
rect 2495 2532 2499 2536
rect 2615 2532 2619 2536
rect 2743 2532 2747 2536
rect 2871 2532 2875 2536
rect 2991 2532 2995 2536
rect 3111 2532 3115 2536
rect 3231 2532 3235 2536
rect 3359 2532 3363 2536
rect 3487 2532 3491 2536
rect 3943 2529 3947 2533
rect 211 2519 215 2523
rect 2459 2523 2463 2527
rect 2571 2523 2575 2527
rect 2691 2523 2695 2527
rect 2819 2523 2823 2527
rect 2827 2523 2831 2527
rect 3067 2523 3071 2527
rect 3075 2523 3079 2527
rect 3195 2523 3199 2527
rect 3315 2523 3319 2527
rect 3443 2523 3447 2527
rect 363 2515 367 2519
rect 523 2515 527 2519
rect 683 2515 687 2519
rect 975 2515 976 2519
rect 976 2515 979 2519
rect 995 2515 999 2519
rect 1139 2515 1143 2519
rect 1275 2515 1279 2519
rect 1411 2515 1415 2519
rect 1539 2515 1543 2519
rect 1667 2515 1671 2519
rect 2047 2512 2051 2516
rect 2383 2513 2387 2517
rect 2495 2513 2499 2517
rect 2615 2513 2619 2517
rect 2743 2513 2747 2517
rect 2871 2513 2875 2517
rect 2991 2513 2995 2517
rect 3111 2513 3115 2517
rect 3231 2513 3235 2517
rect 3359 2513 3363 2517
rect 3487 2513 3491 2517
rect 3943 2512 3947 2516
rect 507 2507 511 2511
rect 203 2483 207 2487
rect 211 2483 215 2487
rect 307 2483 311 2487
rect 403 2483 407 2487
rect 499 2483 503 2487
rect 111 2457 115 2461
rect 135 2460 139 2464
rect 231 2460 235 2464
rect 327 2460 331 2464
rect 423 2460 427 2464
rect 519 2460 523 2464
rect 2007 2457 2011 2461
rect 2047 2456 2051 2460
rect 211 2451 215 2455
rect 307 2451 311 2455
rect 403 2451 407 2455
rect 499 2451 503 2455
rect 2535 2455 2539 2459
rect 507 2451 511 2455
rect 2711 2455 2715 2459
rect 2879 2455 2883 2459
rect 3047 2455 3051 2459
rect 3207 2455 3211 2459
rect 3359 2455 3363 2459
rect 3503 2455 3507 2459
rect 3655 2455 3659 2459
rect 3807 2455 3811 2459
rect 3943 2456 3947 2460
rect 111 2440 115 2444
rect 135 2441 139 2445
rect 231 2441 235 2445
rect 327 2441 331 2445
rect 423 2441 427 2445
rect 519 2441 523 2445
rect 2007 2440 2011 2444
rect 2047 2439 2051 2443
rect 2611 2443 2615 2447
rect 2787 2443 2791 2447
rect 2955 2443 2959 2447
rect 3123 2443 3127 2447
rect 3283 2443 3287 2447
rect 3435 2447 3439 2451
rect 3443 2447 3447 2451
rect 3587 2447 3591 2451
rect 2535 2436 2539 2440
rect 2711 2436 2715 2440
rect 2879 2436 2883 2440
rect 3047 2436 3051 2440
rect 3207 2436 3211 2440
rect 3359 2436 3363 2440
rect 3503 2436 3507 2440
rect 3655 2436 3659 2440
rect 3807 2436 3811 2440
rect 3943 2439 3947 2443
rect 2827 2423 2831 2427
rect 2611 2415 2615 2419
rect 2787 2415 2791 2419
rect 2955 2415 2959 2419
rect 3443 2423 3447 2427
rect 3283 2415 3287 2419
rect 3587 2415 3591 2419
rect 3907 2411 3911 2415
rect 2683 2387 2687 2391
rect 3123 2387 3127 2391
rect 3267 2387 3271 2391
rect 3435 2387 3439 2391
rect 3595 2387 3599 2391
rect 3755 2387 3759 2391
rect 2943 2379 2947 2383
rect 3619 2379 3623 2383
rect 111 2372 115 2376
rect 135 2371 139 2375
rect 203 2367 207 2371
rect 255 2371 259 2375
rect 415 2371 419 2375
rect 575 2371 579 2375
rect 735 2371 739 2375
rect 887 2371 891 2375
rect 1039 2371 1043 2375
rect 1183 2371 1187 2375
rect 1327 2371 1331 2375
rect 1479 2371 1483 2375
rect 2007 2372 2011 2376
rect 219 2363 223 2367
rect 359 2363 363 2367
rect 511 2363 515 2367
rect 703 2363 707 2367
rect 111 2355 115 2359
rect 963 2359 967 2363
rect 971 2363 975 2367
rect 1123 2363 1127 2367
rect 1267 2363 1271 2367
rect 1415 2363 1419 2367
rect 2047 2361 2051 2365
rect 2607 2364 2611 2368
rect 2815 2364 2819 2368
rect 3007 2364 3011 2368
rect 3191 2364 3195 2368
rect 3359 2364 3363 2368
rect 3519 2364 3523 2368
rect 3679 2364 3683 2368
rect 3839 2364 3843 2368
rect 3943 2361 3947 2365
rect 135 2352 139 2356
rect 255 2352 259 2356
rect 415 2352 419 2356
rect 575 2352 579 2356
rect 735 2352 739 2356
rect 887 2352 891 2356
rect 1039 2352 1043 2356
rect 1183 2352 1187 2356
rect 1327 2352 1331 2356
rect 1479 2352 1483 2356
rect 2007 2355 2011 2359
rect 2683 2355 2687 2359
rect 2891 2355 2895 2359
rect 2943 2355 2947 2359
rect 3267 2355 3271 2359
rect 3435 2355 3439 2359
rect 3595 2355 3599 2359
rect 3755 2355 3759 2359
rect 3907 2355 3911 2359
rect 2047 2344 2051 2348
rect 2607 2345 2611 2349
rect 2815 2345 2819 2349
rect 3007 2345 3011 2349
rect 3191 2345 3195 2349
rect 3359 2345 3363 2349
rect 3519 2345 3523 2349
rect 3679 2345 3683 2349
rect 3839 2345 3843 2349
rect 3943 2344 3947 2348
rect 219 2331 223 2335
rect 359 2331 363 2335
rect 511 2331 515 2335
rect 703 2331 707 2335
rect 811 2327 815 2331
rect 971 2331 975 2335
rect 1123 2331 1127 2335
rect 1267 2331 1271 2335
rect 1415 2331 1419 2335
rect 1571 2327 1575 2331
rect 191 2315 192 2319
rect 192 2315 195 2319
rect 211 2315 215 2319
rect 339 2315 343 2319
rect 499 2315 503 2319
rect 659 2315 663 2319
rect 963 2315 967 2319
rect 971 2315 975 2319
rect 1255 2315 1256 2319
rect 1256 2315 1259 2319
rect 1275 2315 1279 2319
rect 1427 2315 1431 2319
rect 111 2289 115 2293
rect 135 2292 139 2296
rect 263 2292 267 2296
rect 423 2292 427 2296
rect 583 2292 587 2296
rect 743 2292 747 2296
rect 895 2292 899 2296
rect 1047 2292 1051 2296
rect 1199 2292 1203 2296
rect 1351 2292 1355 2296
rect 1503 2292 1507 2296
rect 2007 2289 2011 2293
rect 211 2283 215 2287
rect 339 2283 343 2287
rect 499 2283 503 2287
rect 659 2283 663 2287
rect 811 2283 815 2287
rect 971 2283 975 2287
rect 1015 2283 1019 2287
rect 1275 2283 1279 2287
rect 1427 2283 1431 2287
rect 1571 2283 1575 2287
rect 111 2272 115 2276
rect 135 2273 139 2277
rect 263 2273 267 2277
rect 423 2273 427 2277
rect 583 2273 587 2277
rect 743 2273 747 2277
rect 895 2273 899 2277
rect 1047 2273 1051 2277
rect 1199 2273 1203 2277
rect 1351 2273 1355 2277
rect 1503 2273 1507 2277
rect 2007 2272 2011 2276
rect 2047 2276 2051 2280
rect 2071 2275 2075 2279
rect 2167 2275 2171 2279
rect 2271 2275 2275 2279
rect 2415 2275 2419 2279
rect 2575 2275 2579 2279
rect 2743 2275 2747 2279
rect 2911 2275 2915 2279
rect 3071 2275 3075 2279
rect 3231 2275 3235 2279
rect 3383 2275 3387 2279
rect 3535 2275 3539 2279
rect 3695 2275 3699 2279
rect 3943 2276 3947 2280
rect 2047 2259 2051 2263
rect 2147 2263 2151 2267
rect 2243 2263 2247 2267
rect 2251 2267 2255 2271
rect 2359 2267 2363 2271
rect 2535 2267 2539 2271
rect 2659 2267 2663 2271
rect 2871 2267 2875 2271
rect 3147 2263 3151 2267
rect 3307 2263 3311 2267
rect 3459 2263 3463 2267
rect 3611 2263 3615 2267
rect 3619 2267 3623 2271
rect 2071 2256 2075 2260
rect 2167 2256 2171 2260
rect 2271 2256 2275 2260
rect 2415 2256 2419 2260
rect 2575 2256 2579 2260
rect 2743 2256 2747 2260
rect 2911 2256 2915 2260
rect 3071 2256 3075 2260
rect 3231 2256 3235 2260
rect 3383 2256 3387 2260
rect 3535 2256 3539 2260
rect 3695 2256 3699 2260
rect 3943 2259 3947 2263
rect 2251 2243 2255 2247
rect 2147 2235 2151 2239
rect 2359 2235 2363 2239
rect 2535 2235 2539 2239
rect 2659 2235 2663 2239
rect 2699 2231 2703 2235
rect 2891 2235 2895 2239
rect 3451 2243 3455 2247
rect 3147 2235 3151 2239
rect 3307 2235 3311 2239
rect 3459 2235 3463 2239
rect 3611 2235 3615 2239
rect 111 2216 115 2220
rect 223 2215 227 2219
rect 351 2215 355 2219
rect 495 2215 499 2219
rect 647 2215 651 2219
rect 799 2215 803 2219
rect 959 2215 963 2219
rect 1119 2215 1123 2219
rect 1279 2215 1283 2219
rect 1439 2215 1443 2219
rect 1599 2215 1603 2219
rect 2007 2216 2011 2220
rect 2155 2219 2159 2223
rect 2243 2219 2247 2223
rect 2355 2219 2359 2223
rect 2395 2219 2399 2223
rect 2547 2219 2551 2223
rect 2871 2219 2875 2223
rect 2991 2219 2992 2223
rect 2992 2219 2995 2223
rect 3011 2219 3015 2223
rect 3155 2219 3159 2223
rect 3299 2219 3303 2223
rect 3443 2219 3447 2223
rect 191 2207 195 2211
rect 307 2207 311 2211
rect 111 2199 115 2203
rect 1035 2203 1039 2207
rect 1195 2203 1199 2207
rect 1255 2207 1259 2211
rect 223 2196 227 2200
rect 351 2196 355 2200
rect 495 2196 499 2200
rect 647 2196 651 2200
rect 799 2196 803 2200
rect 959 2196 963 2200
rect 1119 2196 1123 2200
rect 1279 2196 1283 2200
rect 1439 2196 1443 2200
rect 1599 2196 1603 2200
rect 2007 2199 2011 2203
rect 2047 2193 2051 2197
rect 2071 2196 2075 2200
rect 2175 2196 2179 2200
rect 2319 2196 2323 2200
rect 2471 2196 2475 2200
rect 2623 2196 2627 2200
rect 2783 2196 2787 2200
rect 2935 2196 2939 2200
rect 3079 2196 3083 2200
rect 3223 2196 3227 2200
rect 3367 2196 3371 2200
rect 3519 2196 3523 2200
rect 3943 2193 3947 2197
rect 2155 2187 2159 2191
rect 2395 2187 2399 2191
rect 2547 2187 2551 2191
rect 2699 2187 2703 2191
rect 2851 2187 2855 2191
rect 3011 2187 3015 2191
rect 3155 2187 3159 2191
rect 3299 2187 3303 2191
rect 3443 2187 3447 2191
rect 3451 2187 3455 2191
rect 307 2175 311 2179
rect 1015 2175 1016 2179
rect 1016 2175 1019 2179
rect 1035 2175 1039 2179
rect 2047 2176 2051 2180
rect 2071 2177 2075 2181
rect 2175 2177 2179 2181
rect 2319 2177 2323 2181
rect 2471 2177 2475 2181
rect 2623 2177 2627 2181
rect 2783 2177 2787 2181
rect 2935 2177 2939 2181
rect 3079 2177 3083 2181
rect 3223 2177 3227 2181
rect 3367 2177 3371 2181
rect 3519 2177 3523 2181
rect 3943 2176 3947 2180
rect 1579 2171 1583 2175
rect 547 2159 551 2163
rect 671 2159 675 2163
rect 891 2159 895 2163
rect 1195 2159 1199 2163
rect 1731 2159 1735 2163
rect 1867 2159 1871 2163
rect 1587 2151 1591 2155
rect 111 2133 115 2137
rect 471 2136 475 2140
rect 567 2136 571 2140
rect 679 2136 683 2140
rect 807 2136 811 2140
rect 943 2136 947 2140
rect 1079 2136 1083 2140
rect 1223 2136 1227 2140
rect 1367 2136 1371 2140
rect 1503 2136 1507 2140
rect 1639 2136 1643 2140
rect 1783 2136 1787 2140
rect 1903 2136 1907 2140
rect 2007 2133 2011 2137
rect 547 2127 551 2131
rect 671 2127 675 2131
rect 891 2127 895 2131
rect 1299 2127 1303 2131
rect 1579 2127 1583 2131
rect 1587 2127 1591 2131
rect 1851 2127 1855 2131
rect 1867 2127 1871 2131
rect 111 2116 115 2120
rect 471 2117 475 2121
rect 567 2117 571 2121
rect 679 2117 683 2121
rect 807 2117 811 2121
rect 943 2117 947 2121
rect 1079 2117 1083 2121
rect 1223 2117 1227 2121
rect 1367 2117 1371 2121
rect 1503 2117 1507 2121
rect 1639 2117 1643 2121
rect 1783 2117 1787 2121
rect 1903 2117 1907 2121
rect 2007 2116 2011 2120
rect 2991 2111 2995 2115
rect 2047 2104 2051 2108
rect 2279 2103 2283 2107
rect 2391 2103 2395 2107
rect 2511 2103 2515 2107
rect 2631 2103 2635 2107
rect 2759 2103 2763 2107
rect 2895 2103 2899 2107
rect 3039 2103 3043 2107
rect 3191 2103 3195 2107
rect 3351 2103 3355 2107
rect 2355 2095 2359 2099
rect 2383 2095 2387 2099
rect 2499 2095 2503 2099
rect 2047 2087 2051 2091
rect 2707 2091 2711 2095
rect 3519 2103 3523 2107
rect 3687 2103 3691 2107
rect 3839 2103 3843 2107
rect 3943 2104 3947 2108
rect 2971 2091 2975 2095
rect 3115 2091 3119 2095
rect 3267 2091 3271 2095
rect 3427 2091 3431 2095
rect 3763 2091 3767 2095
rect 3831 2095 3835 2099
rect 2279 2084 2283 2088
rect 2391 2084 2395 2088
rect 2511 2084 2515 2088
rect 2631 2084 2635 2088
rect 2759 2084 2763 2088
rect 2895 2084 2899 2088
rect 3039 2084 3043 2088
rect 3191 2084 3195 2088
rect 3351 2084 3355 2088
rect 3519 2084 3523 2088
rect 3687 2084 3691 2088
rect 3839 2084 3843 2088
rect 3943 2087 3947 2091
rect 111 2064 115 2068
rect 623 2063 627 2067
rect 735 2063 739 2067
rect 855 2063 859 2067
rect 983 2063 987 2067
rect 1119 2063 1123 2067
rect 1255 2063 1259 2067
rect 1391 2063 1395 2067
rect 1527 2063 1531 2067
rect 1655 2063 1659 2067
rect 1791 2063 1795 2067
rect 1903 2063 1907 2067
rect 2007 2064 2011 2068
rect 2383 2063 2387 2067
rect 2499 2063 2503 2067
rect 111 2047 115 2051
rect 699 2051 703 2055
rect 811 2051 815 2055
rect 931 2051 935 2055
rect 1059 2051 1063 2055
rect 1331 2051 1335 2055
rect 1603 2051 1607 2055
rect 1731 2055 1735 2059
rect 2519 2059 2523 2063
rect 2851 2063 2855 2067
rect 2971 2063 2975 2067
rect 3115 2063 3119 2067
rect 3267 2063 3271 2067
rect 3427 2063 3431 2067
rect 1867 2051 1871 2055
rect 1979 2051 1983 2055
rect 3379 2055 3383 2059
rect 3731 2059 3735 2063
rect 3763 2063 3767 2067
rect 623 2044 627 2048
rect 735 2044 739 2048
rect 855 2044 859 2048
rect 983 2044 987 2048
rect 1119 2044 1123 2048
rect 1255 2044 1259 2048
rect 1391 2044 1395 2048
rect 1527 2044 1531 2048
rect 1655 2044 1659 2048
rect 1791 2044 1795 2048
rect 1903 2044 1907 2048
rect 2007 2047 2011 2051
rect 2403 2039 2407 2043
rect 2619 2039 2623 2043
rect 2703 2039 2704 2043
rect 2704 2039 2707 2043
rect 2843 2039 2847 2043
rect 2851 2039 2855 2043
rect 2995 2039 2999 2043
rect 3155 2039 3159 2043
rect 3339 2039 3343 2043
rect 3739 2039 3743 2043
rect 3907 2039 3911 2043
rect 2527 2031 2531 2035
rect 699 2023 703 2027
rect 811 2023 815 2027
rect 931 2023 935 2027
rect 1059 2023 1063 2027
rect 1299 2023 1303 2027
rect 811 2015 815 2019
rect 1467 2019 1471 2023
rect 1603 2023 1607 2027
rect 1847 2023 1848 2027
rect 1848 2023 1851 2027
rect 1867 2023 1871 2027
rect 2047 2013 2051 2017
rect 2327 2016 2331 2020
rect 2431 2016 2435 2020
rect 2535 2016 2539 2020
rect 2647 2016 2651 2020
rect 2775 2016 2779 2020
rect 2919 2016 2923 2020
rect 3079 2016 3083 2020
rect 3263 2016 3267 2020
rect 3455 2016 3459 2020
rect 3655 2016 3659 2020
rect 3839 2016 3843 2020
rect 3943 2013 3947 2017
rect 515 2003 519 2007
rect 523 2003 527 2007
rect 651 2003 655 2007
rect 803 2003 807 2007
rect 1107 2003 1108 2007
rect 1108 2003 1111 2007
rect 1331 2003 1335 2007
rect 1487 2003 1491 2007
rect 1663 2003 1667 2007
rect 1835 2003 1839 2007
rect 1979 2003 1983 2007
rect 2403 2007 2407 2011
rect 2519 2007 2523 2011
rect 2527 2007 2531 2011
rect 2715 2007 2719 2011
rect 2851 2007 2855 2011
rect 2995 2007 2999 2011
rect 3155 2007 3159 2011
rect 3339 2007 3343 2011
rect 3379 2007 3383 2011
rect 3731 2007 3735 2011
rect 3739 2007 3743 2011
rect 2047 1996 2051 2000
rect 2327 1997 2331 2001
rect 2431 1997 2435 2001
rect 2535 1997 2539 2001
rect 2647 1997 2651 2001
rect 2775 1997 2779 2001
rect 2919 1997 2923 2001
rect 3079 1997 3083 2001
rect 3263 1997 3267 2001
rect 3455 1997 3459 2001
rect 3655 1997 3659 2001
rect 3839 1997 3843 2001
rect 3943 1996 3947 2000
rect 111 1977 115 1981
rect 447 1980 451 1984
rect 575 1980 579 1984
rect 727 1980 731 1984
rect 887 1980 891 1984
rect 1055 1980 1059 1984
rect 1231 1980 1235 1984
rect 1399 1980 1403 1984
rect 1575 1980 1579 1984
rect 1751 1980 1755 1984
rect 1903 1980 1907 1984
rect 2007 1977 2011 1981
rect 523 1971 527 1975
rect 651 1971 655 1975
rect 803 1971 807 1975
rect 811 1971 815 1975
rect 1123 1971 1127 1975
rect 1203 1971 1207 1975
rect 1467 1971 1471 1975
rect 1487 1971 1491 1975
rect 1663 1971 1667 1975
rect 1835 1971 1839 1975
rect 111 1960 115 1964
rect 447 1961 451 1965
rect 575 1961 579 1965
rect 727 1961 731 1965
rect 887 1961 891 1965
rect 1055 1961 1059 1965
rect 1231 1961 1235 1965
rect 1399 1961 1403 1965
rect 1575 1961 1579 1965
rect 1751 1961 1755 1965
rect 1903 1961 1907 1965
rect 2007 1960 2011 1964
rect 2047 1940 2051 1944
rect 2255 1939 2259 1943
rect 2351 1939 2355 1943
rect 2447 1939 2451 1943
rect 2543 1939 2547 1943
rect 2647 1939 2651 1943
rect 2767 1939 2771 1943
rect 2919 1939 2923 1943
rect 3103 1939 3107 1943
rect 3319 1939 3323 1943
rect 3543 1939 3547 1943
rect 3775 1939 3779 1943
rect 3943 1940 3947 1944
rect 2047 1923 2051 1927
rect 2331 1927 2335 1931
rect 2427 1927 2431 1931
rect 2523 1927 2527 1931
rect 2619 1931 2623 1935
rect 2639 1931 2643 1935
rect 2843 1931 2847 1935
rect 2859 1931 2863 1935
rect 3007 1931 3011 1935
rect 3187 1931 3191 1935
rect 3403 1931 3407 1935
rect 3751 1931 3755 1935
rect 2255 1920 2259 1924
rect 2351 1920 2355 1924
rect 2447 1920 2451 1924
rect 2543 1920 2547 1924
rect 2647 1920 2651 1924
rect 2767 1920 2771 1924
rect 2919 1920 2923 1924
rect 3103 1920 3107 1924
rect 3319 1920 3323 1924
rect 3543 1920 3547 1924
rect 3775 1920 3779 1924
rect 3943 1923 3947 1927
rect 111 1908 115 1912
rect 655 1907 659 1911
rect 751 1907 755 1911
rect 847 1907 851 1911
rect 943 1907 947 1911
rect 1039 1907 1043 1911
rect 739 1899 743 1903
rect 931 1899 935 1903
rect 1107 1903 1111 1907
rect 1135 1907 1139 1911
rect 1231 1907 1235 1911
rect 1327 1907 1331 1911
rect 1423 1907 1427 1911
rect 2007 1908 2011 1912
rect 111 1891 115 1895
rect 1307 1895 1311 1899
rect 1403 1895 1407 1899
rect 1499 1895 1503 1899
rect 655 1888 659 1892
rect 751 1888 755 1892
rect 847 1888 851 1892
rect 943 1888 947 1892
rect 1039 1888 1043 1892
rect 1135 1888 1139 1892
rect 1231 1888 1235 1892
rect 1327 1888 1331 1892
rect 1423 1888 1427 1892
rect 2007 1891 2011 1895
rect 2331 1899 2335 1903
rect 2427 1899 2431 1903
rect 2523 1899 2527 1903
rect 2715 1899 2719 1903
rect 2859 1899 2863 1903
rect 3007 1899 3011 1903
rect 3187 1899 3191 1903
rect 3403 1899 3407 1903
rect 2467 1891 2471 1895
rect 3831 1899 3832 1903
rect 3832 1899 3835 1903
rect 739 1867 743 1871
rect 931 1867 935 1871
rect 1123 1867 1127 1871
rect 1203 1867 1207 1871
rect 1307 1871 1311 1875
rect 1335 1863 1339 1867
rect 1403 1867 1407 1871
rect 2203 1871 2207 1875
rect 2459 1871 2463 1875
rect 2639 1871 2643 1875
rect 2667 1871 2671 1875
rect 2871 1871 2875 1875
rect 2907 1871 2911 1875
rect 3067 1871 3071 1875
rect 3259 1871 3263 1875
rect 3475 1871 3479 1875
rect 3907 1871 3911 1875
rect 331 1851 335 1855
rect 395 1851 399 1855
rect 795 1851 799 1855
rect 1067 1851 1071 1855
rect 1203 1851 1207 1855
rect 1483 1851 1487 1855
rect 1499 1851 1503 1855
rect 1171 1843 1175 1847
rect 2047 1845 2051 1849
rect 2183 1848 2187 1852
rect 2279 1848 2283 1852
rect 2383 1848 2387 1852
rect 2487 1848 2491 1852
rect 2591 1848 2595 1852
rect 2703 1848 2707 1852
rect 2831 1848 2835 1852
rect 2991 1848 2995 1852
rect 3183 1848 3187 1852
rect 3399 1848 3403 1852
rect 3631 1848 3635 1852
rect 3839 1848 3843 1852
rect 3943 1845 3947 1849
rect 2459 1839 2463 1843
rect 2467 1839 2471 1843
rect 2667 1839 2671 1843
rect 2771 1839 2775 1843
rect 2907 1839 2911 1843
rect 3067 1839 3071 1843
rect 3259 1839 3263 1843
rect 3475 1839 3479 1843
rect 3915 1839 3919 1843
rect 111 1825 115 1829
rect 319 1828 323 1832
rect 447 1828 451 1832
rect 583 1828 587 1832
rect 719 1828 723 1832
rect 855 1828 859 1832
rect 991 1828 995 1832
rect 1127 1828 1131 1832
rect 1263 1828 1267 1832
rect 1399 1828 1403 1832
rect 1535 1828 1539 1832
rect 2007 1825 2011 1829
rect 2047 1828 2051 1832
rect 2183 1829 2187 1833
rect 2279 1829 2283 1833
rect 2383 1829 2387 1833
rect 2487 1829 2491 1833
rect 2591 1829 2595 1833
rect 2703 1829 2707 1833
rect 2831 1829 2835 1833
rect 2991 1829 2995 1833
rect 3183 1829 3187 1833
rect 3399 1829 3403 1833
rect 3631 1829 3635 1833
rect 3839 1829 3843 1833
rect 3943 1828 3947 1832
rect 395 1819 399 1823
rect 515 1819 519 1823
rect 795 1819 799 1823
rect 923 1819 927 1823
rect 1067 1819 1071 1823
rect 1203 1819 1207 1823
rect 1335 1819 1339 1823
rect 1467 1819 1471 1823
rect 1483 1819 1487 1823
rect 111 1808 115 1812
rect 319 1809 323 1813
rect 447 1809 451 1813
rect 583 1809 587 1813
rect 719 1809 723 1813
rect 855 1809 859 1813
rect 991 1809 995 1813
rect 1127 1809 1131 1813
rect 1263 1809 1267 1813
rect 1399 1809 1403 1813
rect 1535 1809 1539 1813
rect 2007 1808 2011 1812
rect 2047 1772 2051 1776
rect 2127 1771 2131 1775
rect 2311 1771 2315 1775
rect 2495 1771 2499 1775
rect 2687 1771 2691 1775
rect 2879 1771 2883 1775
rect 3071 1771 3075 1775
rect 3263 1771 3267 1775
rect 3463 1771 3467 1775
rect 3663 1771 3667 1775
rect 3839 1771 3843 1775
rect 3943 1772 3947 1776
rect 2203 1763 2207 1767
rect 111 1752 115 1756
rect 255 1751 259 1755
rect 391 1751 395 1755
rect 535 1751 539 1755
rect 695 1751 699 1755
rect 863 1751 867 1755
rect 1031 1751 1035 1755
rect 1207 1751 1211 1755
rect 1383 1751 1387 1755
rect 1559 1751 1563 1755
rect 1743 1751 1747 1755
rect 2007 1752 2011 1756
rect 2047 1755 2051 1759
rect 2799 1759 2803 1763
rect 2871 1763 2875 1767
rect 3159 1763 3163 1767
rect 3347 1763 3351 1767
rect 3907 1767 3911 1771
rect 3739 1759 3743 1763
rect 2127 1752 2131 1756
rect 2311 1752 2315 1756
rect 2495 1752 2499 1756
rect 2687 1752 2691 1756
rect 2879 1752 2883 1756
rect 3071 1752 3075 1756
rect 3263 1752 3267 1756
rect 3463 1752 3467 1756
rect 3663 1752 3667 1756
rect 3839 1752 3843 1756
rect 3943 1755 3947 1759
rect 331 1743 335 1747
rect 343 1743 347 1747
rect 111 1735 115 1739
rect 619 1739 623 1743
rect 663 1743 667 1747
rect 815 1743 819 1747
rect 1107 1739 1111 1743
rect 1171 1743 1175 1747
rect 1519 1739 1523 1743
rect 1635 1739 1639 1743
rect 1819 1739 1823 1743
rect 255 1732 259 1736
rect 391 1732 395 1736
rect 535 1732 539 1736
rect 695 1732 699 1736
rect 863 1732 867 1736
rect 1031 1732 1035 1736
rect 1207 1732 1211 1736
rect 1383 1732 1387 1736
rect 1559 1732 1563 1736
rect 1743 1732 1747 1736
rect 2007 1735 2011 1739
rect 2579 1727 2583 1731
rect 2771 1731 2775 1735
rect 3159 1731 3163 1735
rect 3347 1731 3351 1735
rect 3515 1727 3516 1731
rect 3516 1727 3519 1731
rect 3751 1731 3755 1735
rect 3907 1727 3911 1731
rect 343 1711 347 1715
rect 499 1707 503 1711
rect 663 1711 667 1715
rect 815 1711 819 1715
rect 919 1711 920 1715
rect 920 1711 923 1715
rect 1075 1707 1079 1711
rect 1107 1711 1111 1715
rect 1467 1711 1471 1715
rect 1519 1711 1523 1715
rect 1635 1711 1639 1715
rect 2147 1711 2151 1715
rect 2267 1711 2271 1715
rect 2419 1711 2423 1715
rect 2791 1711 2795 1715
rect 2799 1711 2803 1715
rect 3119 1711 3120 1715
rect 3120 1711 3123 1715
rect 3139 1711 3143 1715
rect 3331 1711 3335 1715
rect 3739 1711 3743 1715
rect 3915 1711 3919 1715
rect 2299 1703 2303 1707
rect 203 1695 207 1699
rect 211 1695 215 1699
rect 339 1695 343 1699
rect 619 1695 623 1699
rect 683 1695 687 1699
rect 1255 1695 1256 1699
rect 1256 1695 1259 1699
rect 1275 1695 1279 1699
rect 1707 1695 1711 1699
rect 1819 1695 1823 1699
rect 1303 1683 1307 1687
rect 2047 1685 2051 1689
rect 2071 1688 2075 1692
rect 2191 1688 2195 1692
rect 2343 1688 2347 1692
rect 2511 1688 2515 1692
rect 2687 1688 2691 1692
rect 2871 1688 2875 1692
rect 3063 1688 3067 1692
rect 3255 1688 3259 1692
rect 3447 1688 3451 1692
rect 3647 1688 3651 1692
rect 3839 1688 3843 1692
rect 3943 1685 3947 1689
rect 2147 1679 2151 1683
rect 2267 1679 2271 1683
rect 2419 1679 2423 1683
rect 2579 1679 2583 1683
rect 2655 1679 2659 1683
rect 2791 1679 2795 1683
rect 3139 1679 3143 1683
rect 3331 1679 3335 1683
rect 3515 1679 3519 1683
rect 3615 1679 3619 1683
rect 3907 1679 3911 1683
rect 111 1669 115 1673
rect 135 1672 139 1676
rect 263 1672 267 1676
rect 431 1672 435 1676
rect 607 1672 611 1676
rect 799 1672 803 1676
rect 999 1672 1003 1676
rect 1199 1672 1203 1676
rect 1407 1672 1411 1676
rect 1623 1672 1627 1676
rect 1839 1672 1843 1676
rect 2007 1669 2011 1673
rect 2047 1668 2051 1672
rect 2071 1669 2075 1673
rect 2191 1669 2195 1673
rect 2343 1669 2347 1673
rect 2511 1669 2515 1673
rect 2687 1669 2691 1673
rect 2871 1669 2875 1673
rect 3063 1669 3067 1673
rect 3255 1669 3259 1673
rect 3447 1669 3451 1673
rect 3647 1669 3651 1673
rect 3839 1669 3843 1673
rect 3943 1668 3947 1672
rect 211 1663 215 1667
rect 339 1663 343 1667
rect 499 1663 503 1667
rect 683 1663 687 1667
rect 875 1663 879 1667
rect 1075 1663 1079 1667
rect 1275 1663 1279 1667
rect 1303 1663 1307 1667
rect 1559 1663 1563 1667
rect 1707 1663 1711 1667
rect 111 1652 115 1656
rect 135 1653 139 1657
rect 263 1653 267 1657
rect 431 1653 435 1657
rect 607 1653 611 1657
rect 799 1653 803 1657
rect 999 1653 1003 1657
rect 1199 1653 1203 1657
rect 1407 1653 1411 1657
rect 1623 1653 1627 1657
rect 1839 1653 1843 1657
rect 2007 1652 2011 1656
rect 2047 1616 2051 1620
rect 2071 1615 2075 1619
rect 2335 1615 2339 1619
rect 2599 1615 2603 1619
rect 2839 1615 2843 1619
rect 3047 1615 3051 1619
rect 3231 1615 3235 1619
rect 3399 1615 3403 1619
rect 3551 1615 3555 1619
rect 3695 1615 3699 1619
rect 3839 1615 3843 1619
rect 3943 1616 3947 1620
rect 111 1600 115 1604
rect 135 1599 139 1603
rect 203 1595 207 1599
rect 287 1599 291 1603
rect 471 1599 475 1603
rect 655 1599 659 1603
rect 839 1599 843 1603
rect 1015 1599 1019 1603
rect 1183 1599 1187 1603
rect 1343 1599 1347 1603
rect 1495 1599 1499 1603
rect 1639 1599 1643 1603
rect 1783 1599 1787 1603
rect 1903 1599 1907 1603
rect 2007 1600 2011 1604
rect 2047 1599 2051 1603
rect 2147 1603 2151 1607
rect 2299 1607 2303 1611
rect 2675 1603 2679 1607
rect 2915 1603 2919 1607
rect 3123 1607 3127 1611
rect 3131 1607 3135 1611
rect 3355 1607 3359 1611
rect 3627 1603 3631 1607
rect 3771 1603 3775 1607
rect 3915 1607 3919 1611
rect 2071 1596 2075 1600
rect 223 1591 227 1595
rect 111 1583 115 1587
rect 547 1587 551 1591
rect 731 1587 735 1591
rect 739 1591 743 1595
rect 1119 1587 1123 1591
rect 1259 1591 1263 1595
rect 2335 1596 2339 1600
rect 2599 1596 2603 1600
rect 2839 1596 2843 1600
rect 3047 1596 3051 1600
rect 3231 1596 3235 1600
rect 3399 1596 3403 1600
rect 3551 1596 3555 1600
rect 3695 1596 3699 1600
rect 3839 1596 3843 1600
rect 3943 1599 3947 1603
rect 1279 1591 1283 1595
rect 1571 1587 1575 1591
rect 1715 1587 1719 1591
rect 1859 1587 1863 1591
rect 135 1580 139 1584
rect 287 1580 291 1584
rect 471 1580 475 1584
rect 655 1580 659 1584
rect 839 1580 843 1584
rect 1015 1580 1019 1584
rect 1183 1580 1187 1584
rect 1343 1580 1347 1584
rect 1495 1580 1499 1584
rect 1639 1580 1643 1584
rect 1783 1580 1787 1584
rect 1903 1580 1907 1584
rect 2007 1583 2011 1587
rect 2147 1575 2151 1579
rect 2655 1575 2656 1579
rect 2656 1575 2659 1579
rect 3131 1583 3135 1587
rect 2915 1575 2919 1579
rect 3355 1575 3359 1579
rect 223 1559 227 1563
rect 391 1555 395 1559
rect 739 1567 743 1571
rect 1279 1567 1283 1571
rect 3451 1571 3452 1575
rect 3452 1571 3455 1575
rect 3615 1575 3619 1579
rect 3627 1575 3631 1579
rect 3891 1571 3892 1575
rect 3892 1571 3895 1575
rect 547 1559 551 1563
rect 875 1559 879 1563
rect 1119 1555 1123 1559
rect 1351 1555 1355 1559
rect 1559 1559 1563 1563
rect 1571 1559 1575 1563
rect 1715 1559 1719 1563
rect 1859 1559 1863 1563
rect 2675 1555 2679 1559
rect 2711 1555 2715 1559
rect 2819 1555 2823 1559
rect 2979 1555 2983 1559
rect 3299 1555 3303 1559
rect 3639 1555 3643 1559
rect 3771 1555 3775 1559
rect 3499 1547 3503 1551
rect 251 1539 255 1543
rect 259 1539 263 1543
rect 371 1539 375 1543
rect 731 1539 735 1543
rect 763 1539 767 1543
rect 1155 1539 1159 1543
rect 1531 1539 1535 1543
rect 1707 1539 1711 1543
rect 1863 1539 1864 1543
rect 1864 1539 1867 1543
rect 1399 1531 1403 1535
rect 2047 1529 2051 1533
rect 2583 1532 2587 1536
rect 2743 1532 2747 1536
rect 2903 1532 2907 1536
rect 3063 1532 3067 1536
rect 3223 1532 3227 1536
rect 3383 1532 3387 1536
rect 3543 1532 3547 1536
rect 3703 1532 3707 1536
rect 3943 1529 3947 1533
rect 2711 1523 2715 1527
rect 2819 1523 2823 1527
rect 2979 1523 2983 1527
rect 3019 1523 3023 1527
rect 3299 1523 3303 1527
rect 3451 1523 3455 1527
rect 3499 1523 3503 1527
rect 3639 1523 3643 1527
rect 111 1513 115 1517
rect 135 1516 139 1520
rect 295 1516 299 1520
rect 487 1516 491 1520
rect 687 1516 691 1520
rect 887 1516 891 1520
rect 1079 1516 1083 1520
rect 1263 1516 1267 1520
rect 1447 1516 1451 1520
rect 1623 1516 1627 1520
rect 1807 1516 1811 1520
rect 2007 1513 2011 1517
rect 2047 1512 2051 1516
rect 2583 1513 2587 1517
rect 2743 1513 2747 1517
rect 2903 1513 2907 1517
rect 3063 1513 3067 1517
rect 3223 1513 3227 1517
rect 3383 1513 3387 1517
rect 3543 1513 3547 1517
rect 3703 1513 3707 1517
rect 3943 1512 3947 1516
rect 259 1507 263 1511
rect 371 1507 375 1511
rect 391 1507 395 1511
rect 763 1507 767 1511
rect 839 1507 843 1511
rect 1155 1507 1159 1511
rect 1351 1507 1355 1511
rect 1399 1507 1403 1511
rect 1531 1507 1535 1511
rect 1707 1507 1711 1511
rect 111 1496 115 1500
rect 135 1497 139 1501
rect 295 1497 299 1501
rect 487 1497 491 1501
rect 687 1497 691 1501
rect 887 1497 891 1501
rect 1079 1497 1083 1501
rect 1263 1497 1267 1501
rect 1447 1497 1451 1501
rect 1623 1497 1627 1501
rect 1807 1497 1811 1501
rect 2007 1496 2011 1500
rect 2047 1460 2051 1464
rect 2415 1459 2419 1463
rect 2511 1459 2515 1463
rect 2607 1459 2611 1463
rect 2703 1459 2707 1463
rect 2799 1459 2803 1463
rect 2919 1459 2923 1463
rect 3063 1459 3067 1463
rect 3231 1459 3235 1463
rect 3415 1459 3419 1463
rect 3615 1459 3619 1463
rect 3815 1459 3819 1463
rect 3943 1460 3947 1464
rect 111 1444 115 1448
rect 175 1443 179 1447
rect 359 1443 363 1447
rect 567 1443 571 1447
rect 783 1443 787 1447
rect 1007 1443 1011 1447
rect 1231 1443 1235 1447
rect 1463 1443 1467 1447
rect 1695 1443 1699 1447
rect 1903 1443 1907 1447
rect 2007 1444 2011 1448
rect 2047 1443 2051 1447
rect 2491 1447 2495 1451
rect 2587 1447 2591 1451
rect 2683 1447 2687 1451
rect 2779 1447 2783 1451
rect 2875 1447 2879 1451
rect 2995 1447 2999 1451
rect 3139 1447 3143 1451
rect 3307 1447 3311 1451
rect 3491 1447 3495 1451
rect 3559 1451 3563 1455
rect 3891 1451 3895 1455
rect 2415 1440 2419 1444
rect 251 1435 255 1439
rect 275 1435 279 1439
rect 443 1435 447 1439
rect 111 1427 115 1431
rect 1083 1431 1087 1435
rect 2511 1440 2515 1444
rect 2607 1440 2611 1444
rect 2703 1440 2707 1444
rect 2799 1440 2803 1444
rect 2919 1440 2923 1444
rect 3063 1440 3067 1444
rect 3231 1440 3235 1444
rect 3415 1440 3419 1444
rect 3615 1440 3619 1444
rect 3815 1440 3819 1444
rect 3943 1443 3947 1447
rect 1539 1431 1543 1435
rect 1771 1431 1775 1435
rect 1863 1435 1867 1439
rect 175 1424 179 1428
rect 359 1424 363 1428
rect 567 1424 571 1428
rect 783 1424 787 1428
rect 1007 1424 1011 1428
rect 1231 1424 1235 1428
rect 1463 1424 1467 1428
rect 1695 1424 1699 1428
rect 1903 1424 1907 1428
rect 2007 1427 2011 1431
rect 2627 1431 2631 1435
rect 3559 1431 3563 1435
rect 2491 1419 2495 1423
rect 2587 1419 2591 1423
rect 2683 1419 2687 1423
rect 2779 1419 2783 1423
rect 2875 1419 2879 1423
rect 2995 1419 2999 1423
rect 3139 1419 3143 1423
rect 3307 1419 3311 1423
rect 3491 1419 3495 1423
rect 3019 1411 3023 1415
rect 3883 1415 3887 1419
rect 275 1403 279 1407
rect 403 1399 407 1403
rect 839 1403 840 1407
rect 840 1403 843 1407
rect 931 1399 935 1403
rect 1083 1403 1087 1407
rect 1539 1403 1543 1407
rect 1771 1403 1775 1407
rect 1667 1395 1671 1399
rect 443 1387 447 1391
rect 519 1387 520 1391
rect 520 1387 523 1391
rect 539 1387 543 1391
rect 675 1387 679 1391
rect 803 1387 807 1391
rect 1059 1387 1063 1391
rect 1195 1387 1199 1391
rect 1339 1387 1343 1391
rect 1835 1387 1839 1391
rect 1987 1387 1991 1391
rect 1403 1379 1407 1383
rect 2155 1383 2159 1387
rect 2311 1383 2315 1387
rect 2627 1383 2631 1387
rect 2635 1383 2639 1387
rect 2883 1383 2887 1387
rect 3131 1383 3135 1387
rect 3379 1383 3383 1387
rect 3907 1383 3911 1387
rect 111 1361 115 1365
rect 327 1364 331 1368
rect 463 1364 467 1368
rect 599 1364 603 1368
rect 727 1364 731 1368
rect 855 1364 859 1368
rect 983 1364 987 1368
rect 1119 1364 1123 1368
rect 1263 1364 1267 1368
rect 1423 1364 1427 1368
rect 1583 1364 1587 1368
rect 1751 1364 1755 1368
rect 1903 1364 1907 1368
rect 2007 1361 2011 1365
rect 403 1355 407 1359
rect 539 1355 543 1359
rect 675 1355 679 1359
rect 803 1355 807 1359
rect 931 1355 935 1359
rect 1059 1355 1063 1359
rect 1195 1355 1199 1359
rect 1339 1355 1343 1359
rect 111 1344 115 1348
rect 327 1345 331 1349
rect 463 1345 467 1349
rect 599 1345 603 1349
rect 727 1345 731 1349
rect 855 1345 859 1349
rect 983 1345 987 1349
rect 1119 1345 1123 1349
rect 1263 1345 1267 1349
rect 1179 1339 1183 1343
rect 1651 1355 1655 1359
rect 1667 1355 1671 1359
rect 1835 1355 1839 1359
rect 2047 1357 2051 1361
rect 2071 1360 2075 1364
rect 2303 1360 2307 1364
rect 2559 1360 2563 1364
rect 2807 1360 2811 1364
rect 3055 1360 3059 1364
rect 3303 1360 3307 1364
rect 3559 1360 3563 1364
rect 3815 1360 3819 1364
rect 3943 1357 3947 1361
rect 1987 1351 1991 1355
rect 2155 1351 2159 1355
rect 2635 1351 2639 1355
rect 2883 1351 2887 1355
rect 3131 1351 3135 1355
rect 3379 1351 3383 1355
rect 3883 1351 3887 1355
rect 1423 1345 1427 1349
rect 1583 1345 1587 1349
rect 1751 1345 1755 1349
rect 1903 1345 1907 1349
rect 2007 1344 2011 1348
rect 2047 1340 2051 1344
rect 2071 1341 2075 1345
rect 2303 1341 2307 1345
rect 2559 1341 2563 1345
rect 2807 1341 2811 1345
rect 3055 1341 3059 1345
rect 3303 1341 3307 1345
rect 3559 1341 3563 1345
rect 3815 1341 3819 1345
rect 3943 1340 3947 1344
rect 3055 1295 3059 1299
rect 111 1284 115 1288
rect 551 1283 555 1287
rect 655 1283 659 1287
rect 767 1283 771 1287
rect 879 1283 883 1287
rect 991 1283 995 1287
rect 1103 1283 1107 1287
rect 1215 1283 1219 1287
rect 1327 1283 1331 1287
rect 1439 1283 1443 1287
rect 1559 1283 1563 1287
rect 2007 1284 2011 1288
rect 2047 1280 2051 1284
rect 111 1267 115 1271
rect 627 1271 631 1275
rect 731 1271 735 1275
rect 843 1271 847 1275
rect 955 1271 959 1275
rect 963 1275 967 1279
rect 1087 1275 1091 1279
rect 1291 1271 1295 1275
rect 1403 1275 1407 1279
rect 2071 1279 2075 1283
rect 1515 1271 1519 1275
rect 1527 1275 1531 1279
rect 2223 1279 2227 1283
rect 2415 1279 2419 1283
rect 2615 1279 2619 1283
rect 2815 1279 2819 1283
rect 2999 1279 3003 1283
rect 3175 1279 3179 1283
rect 3343 1279 3347 1283
rect 3503 1279 3507 1283
rect 3663 1279 3667 1283
rect 3831 1279 3835 1283
rect 3943 1280 3947 1284
rect 551 1264 555 1268
rect 655 1264 659 1268
rect 767 1264 771 1268
rect 879 1264 883 1268
rect 991 1264 995 1268
rect 1103 1264 1107 1268
rect 1215 1264 1219 1268
rect 1327 1264 1331 1268
rect 1439 1264 1443 1268
rect 1559 1264 1563 1268
rect 2007 1267 2011 1271
rect 2047 1263 2051 1267
rect 2147 1267 2151 1271
rect 2311 1271 2315 1275
rect 2359 1271 2363 1275
rect 2691 1267 2695 1271
rect 2699 1271 2703 1275
rect 3075 1267 3079 1271
rect 3251 1267 3255 1271
rect 3419 1267 3423 1271
rect 3579 1267 3583 1271
rect 3739 1267 3743 1271
rect 3907 1271 3911 1275
rect 2071 1260 2075 1264
rect 2223 1260 2227 1264
rect 2415 1260 2419 1264
rect 2615 1260 2619 1264
rect 2815 1260 2819 1264
rect 2999 1260 3003 1264
rect 3175 1260 3179 1264
rect 3343 1260 3347 1264
rect 3503 1260 3507 1264
rect 3663 1260 3667 1264
rect 3831 1260 3835 1264
rect 3943 1263 3947 1267
rect 627 1243 631 1247
rect 731 1243 735 1247
rect 843 1243 847 1247
rect 955 1243 959 1247
rect 1179 1243 1183 1247
rect 939 1235 943 1239
rect 1187 1239 1191 1243
rect 1291 1243 1295 1247
rect 1527 1243 1531 1247
rect 1651 1243 1655 1247
rect 2359 1247 2363 1251
rect 2147 1239 2151 1243
rect 2699 1247 2703 1251
rect 2579 1235 2583 1239
rect 2691 1239 2695 1243
rect 3055 1239 3056 1243
rect 3056 1239 3059 1243
rect 3075 1239 3079 1243
rect 3251 1239 3255 1243
rect 3419 1239 3423 1243
rect 3579 1239 3583 1243
rect 3907 1235 3911 1239
rect 467 1227 471 1231
rect 595 1227 599 1231
rect 739 1227 743 1231
rect 1195 1227 1199 1231
rect 1283 1227 1287 1231
rect 1515 1227 1519 1231
rect 1635 1227 1639 1231
rect 799 1219 803 1223
rect 2211 1215 2215 1219
rect 2387 1215 2391 1219
rect 2915 1215 2919 1219
rect 3147 1215 3151 1219
rect 3315 1215 3319 1219
rect 3739 1215 3743 1219
rect 3915 1215 3919 1219
rect 111 1201 115 1205
rect 391 1204 395 1208
rect 519 1204 523 1208
rect 663 1204 667 1208
rect 807 1204 811 1208
rect 959 1204 963 1208
rect 1111 1204 1115 1208
rect 1255 1204 1259 1208
rect 1407 1204 1411 1208
rect 1559 1204 1563 1208
rect 1711 1204 1715 1208
rect 2659 1207 2663 1211
rect 3499 1207 3503 1211
rect 2007 1201 2011 1205
rect 467 1195 471 1199
rect 595 1195 599 1199
rect 739 1195 743 1199
rect 939 1195 943 1199
rect 1187 1195 1191 1199
rect 1195 1195 1199 1199
rect 1635 1195 1639 1199
rect 1663 1195 1667 1199
rect 111 1184 115 1188
rect 391 1185 395 1189
rect 519 1185 523 1189
rect 663 1185 667 1189
rect 807 1185 811 1189
rect 959 1185 963 1189
rect 1111 1185 1115 1189
rect 1255 1185 1259 1189
rect 1407 1185 1411 1189
rect 1559 1185 1563 1189
rect 2047 1189 2051 1193
rect 2135 1192 2139 1196
rect 2311 1192 2315 1196
rect 2503 1192 2507 1196
rect 2695 1192 2699 1196
rect 2887 1192 2891 1196
rect 3071 1192 3075 1196
rect 3239 1192 3243 1196
rect 3399 1192 3403 1196
rect 3551 1192 3555 1196
rect 3703 1192 3707 1196
rect 3839 1192 3843 1196
rect 1711 1185 1715 1189
rect 3943 1189 3947 1193
rect 2007 1184 2011 1188
rect 2211 1183 2215 1187
rect 2387 1183 2391 1187
rect 2579 1183 2583 1187
rect 2659 1183 2663 1187
rect 3147 1183 3151 1187
rect 3315 1183 3319 1187
rect 3475 1183 3479 1187
rect 3499 1183 3503 1187
rect 3907 1183 3911 1187
rect 2047 1172 2051 1176
rect 2135 1173 2139 1177
rect 2311 1173 2315 1177
rect 2503 1173 2507 1177
rect 2695 1173 2699 1177
rect 2887 1173 2891 1177
rect 3071 1173 3075 1177
rect 3239 1173 3243 1177
rect 3399 1173 3403 1177
rect 3551 1173 3555 1177
rect 3703 1173 3707 1177
rect 3839 1173 3843 1177
rect 3943 1172 3947 1176
rect 111 1128 115 1132
rect 175 1127 179 1131
rect 327 1127 331 1131
rect 495 1127 499 1131
rect 671 1127 675 1131
rect 847 1127 851 1131
rect 1031 1127 1035 1131
rect 1207 1127 1211 1131
rect 1383 1127 1387 1131
rect 1567 1127 1571 1131
rect 1751 1127 1755 1131
rect 2007 1128 2011 1132
rect 111 1111 115 1115
rect 251 1115 255 1119
rect 403 1115 407 1119
rect 571 1115 575 1119
rect 747 1115 751 1119
rect 799 1119 803 1123
rect 1107 1115 1111 1119
rect 1283 1119 1287 1123
rect 1327 1119 1331 1123
rect 1839 1115 1843 1119
rect 175 1108 179 1112
rect 327 1108 331 1112
rect 495 1108 499 1112
rect 671 1108 675 1112
rect 847 1108 851 1112
rect 1031 1108 1035 1112
rect 1207 1108 1211 1112
rect 1383 1108 1387 1112
rect 1567 1108 1571 1112
rect 1751 1108 1755 1112
rect 2007 1111 2011 1115
rect 2047 1112 2051 1116
rect 2295 1111 2299 1115
rect 2423 1111 2427 1115
rect 2559 1111 2563 1115
rect 2695 1111 2699 1115
rect 2839 1111 2843 1115
rect 2991 1111 2995 1115
rect 3151 1111 3155 1115
rect 3319 1111 3323 1115
rect 3495 1111 3499 1115
rect 3679 1111 3683 1115
rect 3839 1111 3843 1115
rect 3943 1112 3947 1116
rect 2047 1095 2051 1099
rect 2371 1099 2375 1103
rect 2499 1099 2503 1103
rect 2635 1099 2639 1103
rect 2771 1099 2775 1103
rect 2915 1103 2919 1107
rect 3067 1099 3071 1103
rect 3227 1099 3231 1103
rect 3259 1103 3263 1107
rect 3571 1099 3575 1103
rect 3579 1103 3583 1107
rect 3915 1103 3919 1107
rect 2295 1092 2299 1096
rect 243 1083 247 1087
rect 251 1087 255 1091
rect 403 1087 407 1091
rect 571 1087 575 1091
rect 747 1087 751 1091
rect 1087 1087 1088 1091
rect 1088 1087 1091 1091
rect 1327 1087 1331 1091
rect 1663 1087 1667 1091
rect 2423 1092 2427 1096
rect 2559 1092 2563 1096
rect 2695 1092 2699 1096
rect 2839 1092 2843 1096
rect 2991 1092 2995 1096
rect 3151 1092 3155 1096
rect 3319 1092 3323 1096
rect 3495 1092 3499 1096
rect 3679 1092 3683 1096
rect 3839 1092 3843 1096
rect 3943 1095 3947 1099
rect 2371 1075 2375 1079
rect 203 1063 207 1067
rect 211 1063 215 1067
rect 307 1063 311 1067
rect 451 1063 455 1067
rect 619 1063 623 1067
rect 803 1063 807 1067
rect 1107 1063 1111 1067
rect 1327 1063 1331 1067
rect 1355 1063 1359 1067
rect 1735 1063 1739 1067
rect 1839 1063 1843 1067
rect 2499 1071 2503 1075
rect 2635 1071 2639 1075
rect 2771 1071 2775 1075
rect 3259 1079 3263 1083
rect 3067 1071 3071 1075
rect 3579 1079 3583 1083
rect 3475 1071 3479 1075
rect 3571 1071 3575 1075
rect 3907 1067 3911 1071
rect 2579 1051 2583 1055
rect 2683 1051 2687 1055
rect 2923 1051 2927 1055
rect 3191 1051 3195 1055
rect 3227 1051 3231 1055
rect 3275 1051 3279 1055
rect 3483 1051 3487 1055
rect 3915 1051 3919 1055
rect 111 1037 115 1041
rect 135 1040 139 1044
rect 231 1040 235 1044
rect 375 1040 379 1044
rect 543 1040 547 1044
rect 727 1040 731 1044
rect 911 1040 915 1044
rect 1095 1040 1099 1044
rect 1279 1040 1283 1044
rect 1463 1040 1467 1044
rect 1647 1040 1651 1044
rect 1831 1040 1835 1044
rect 2007 1037 2011 1041
rect 211 1031 215 1035
rect 307 1031 311 1035
rect 451 1031 455 1035
rect 619 1031 623 1035
rect 803 1031 807 1035
rect 859 1031 863 1035
rect 1063 1031 1067 1035
rect 1355 1031 1359 1035
rect 1555 1031 1559 1035
rect 1735 1031 1739 1035
rect 111 1020 115 1024
rect 135 1021 139 1025
rect 231 1021 235 1025
rect 375 1021 379 1025
rect 543 1021 547 1025
rect 727 1021 731 1025
rect 911 1021 915 1025
rect 1095 1021 1099 1025
rect 1279 1021 1283 1025
rect 1463 1021 1467 1025
rect 1647 1021 1651 1025
rect 2047 1025 2051 1029
rect 2495 1028 2499 1032
rect 2599 1028 2603 1032
rect 2711 1028 2715 1032
rect 2847 1028 2851 1032
rect 3007 1028 3011 1032
rect 3199 1028 3203 1032
rect 3407 1028 3411 1032
rect 3631 1028 3635 1032
rect 3839 1028 3843 1032
rect 1831 1021 1835 1025
rect 3943 1025 3947 1029
rect 2007 1020 2011 1024
rect 2579 1019 2583 1023
rect 2683 1019 2687 1023
rect 3075 1019 3079 1023
rect 3275 1019 3279 1023
rect 3483 1019 3487 1023
rect 3559 1019 3563 1023
rect 3907 1019 3911 1023
rect 2047 1008 2051 1012
rect 2495 1009 2499 1013
rect 2599 1009 2603 1013
rect 2711 1009 2715 1013
rect 2847 1009 2851 1013
rect 3007 1009 3011 1013
rect 3199 1009 3203 1013
rect 3407 1009 3411 1013
rect 3631 1009 3635 1013
rect 3839 1009 3843 1013
rect 3943 1008 3947 1012
rect 111 968 115 972
rect 135 967 139 971
rect 203 963 207 967
rect 271 967 275 971
rect 447 967 451 971
rect 631 967 635 971
rect 823 967 827 971
rect 1007 967 1011 971
rect 1175 967 1179 971
rect 1335 967 1339 971
rect 1487 967 1491 971
rect 1631 967 1635 971
rect 1775 967 1779 971
rect 1903 967 1907 971
rect 2007 968 2011 972
rect 251 959 255 963
rect 587 959 591 963
rect 715 959 719 963
rect 111 951 115 955
rect 1083 955 1087 959
rect 1251 955 1255 959
rect 1327 959 1331 963
rect 1563 955 1567 959
rect 1707 955 1711 959
rect 1851 955 1855 959
rect 1871 959 1875 963
rect 2047 956 2051 960
rect 2647 955 2651 959
rect 135 948 139 952
rect 271 948 275 952
rect 447 948 451 952
rect 631 948 635 952
rect 823 948 827 952
rect 1007 948 1011 952
rect 1175 948 1179 952
rect 1335 948 1339 952
rect 1487 948 1491 952
rect 1631 948 1635 952
rect 1775 948 1779 952
rect 1903 948 1907 952
rect 2007 951 2011 955
rect 2743 955 2747 959
rect 2847 955 2851 959
rect 2967 955 2971 959
rect 3111 955 3115 959
rect 3279 955 3283 959
rect 3463 955 3467 959
rect 3663 955 3667 959
rect 3839 955 3843 959
rect 3943 956 3947 960
rect 2047 939 2051 943
rect 2723 943 2727 947
rect 2819 943 2823 947
rect 2923 947 2927 951
rect 3087 943 3091 947
rect 3187 943 3191 947
rect 3355 943 3359 947
rect 3539 943 3543 947
rect 3623 947 3627 951
rect 3915 947 3919 951
rect 2647 936 2651 940
rect 2743 936 2747 940
rect 2847 936 2851 940
rect 2967 936 2971 940
rect 3111 936 3115 940
rect 3279 936 3283 940
rect 3463 936 3467 940
rect 3663 936 3667 940
rect 3839 936 3843 940
rect 3943 939 3947 943
rect 251 927 255 931
rect 587 927 591 931
rect 715 927 719 931
rect 923 923 927 927
rect 1063 927 1064 931
rect 1064 927 1067 931
rect 1231 923 1232 927
rect 1232 923 1235 927
rect 1251 927 1255 931
rect 1555 927 1559 931
rect 1563 927 1567 931
rect 1707 927 1711 931
rect 1851 927 1855 931
rect 1871 919 1875 923
rect 2723 919 2727 923
rect 191 911 192 915
rect 192 911 195 915
rect 211 911 215 915
rect 347 911 351 915
rect 531 911 535 915
rect 731 911 735 915
rect 1083 911 1087 915
rect 1323 911 1327 915
rect 1499 911 1503 915
rect 1611 911 1615 915
rect 1827 911 1831 915
rect 2751 911 2755 915
rect 2819 915 2823 919
rect 3075 915 3079 919
rect 3087 915 3091 919
rect 3187 915 3191 919
rect 3355 915 3359 919
rect 3539 915 3543 919
rect 3907 911 3911 915
rect 3623 895 3627 899
rect 111 885 115 889
rect 135 888 139 892
rect 271 888 275 892
rect 455 888 459 892
rect 655 888 659 892
rect 855 888 859 892
rect 1055 888 1059 892
rect 1239 888 1243 892
rect 1415 888 1419 892
rect 1583 888 1587 892
rect 1751 888 1755 892
rect 1903 888 1907 892
rect 2007 885 2011 889
rect 2147 887 2151 891
rect 2331 887 2335 891
rect 211 879 215 883
rect 347 879 351 883
rect 531 879 535 883
rect 731 879 735 883
rect 923 879 927 883
rect 1167 879 1171 883
rect 1231 879 1235 883
rect 1323 879 1327 883
rect 1499 879 1503 883
rect 1827 879 1831 883
rect 2971 883 2975 887
rect 3203 887 3207 891
rect 3443 887 3447 891
rect 3915 887 3919 891
rect 111 868 115 872
rect 135 869 139 873
rect 271 869 275 873
rect 455 869 459 873
rect 655 869 659 873
rect 855 869 859 873
rect 1055 869 1059 873
rect 1239 869 1243 873
rect 1415 869 1419 873
rect 1583 869 1587 873
rect 1751 869 1755 873
rect 1903 869 1907 873
rect 2007 868 2011 872
rect 2047 861 2051 865
rect 2071 864 2075 868
rect 2255 864 2259 868
rect 2463 864 2467 868
rect 2679 864 2683 868
rect 2895 864 2899 868
rect 3127 864 3131 868
rect 3367 864 3371 868
rect 3615 864 3619 868
rect 3839 864 3843 868
rect 3943 861 3947 865
rect 2147 855 2151 859
rect 2331 855 2335 859
rect 2351 855 2355 859
rect 2751 855 2755 859
rect 3203 855 3207 859
rect 3443 855 3447 859
rect 3691 855 3695 859
rect 3907 855 3911 859
rect 2047 844 2051 848
rect 2071 845 2075 849
rect 2255 845 2259 849
rect 2463 845 2467 849
rect 2679 845 2683 849
rect 2895 845 2899 849
rect 3127 845 3131 849
rect 3367 845 3371 849
rect 3615 845 3619 849
rect 3839 845 3843 849
rect 3943 844 3947 848
rect 111 816 115 820
rect 215 815 219 819
rect 343 815 347 819
rect 495 815 499 819
rect 655 815 659 819
rect 831 815 835 819
rect 1007 815 1011 819
rect 1183 815 1187 819
rect 1359 815 1363 819
rect 1535 815 1539 819
rect 1719 815 1723 819
rect 2007 816 2011 820
rect 191 807 195 811
rect 331 807 335 811
rect 615 807 619 811
rect 111 799 115 803
rect 1083 803 1087 807
rect 1095 807 1099 811
rect 1463 803 1467 807
rect 1611 807 1615 811
rect 1639 807 1643 811
rect 215 796 219 800
rect 343 796 347 800
rect 495 796 499 800
rect 655 796 659 800
rect 831 796 835 800
rect 1007 796 1011 800
rect 1183 796 1187 800
rect 1359 796 1363 800
rect 1535 796 1539 800
rect 1719 796 1723 800
rect 2007 799 2011 803
rect 2047 792 2051 796
rect 2215 791 2219 795
rect 2327 791 2331 795
rect 2447 791 2451 795
rect 2583 791 2587 795
rect 2735 791 2739 795
rect 2895 791 2899 795
rect 3063 791 3067 795
rect 3247 791 3251 795
rect 3447 791 3451 795
rect 3655 791 3659 795
rect 3839 791 3843 795
rect 3943 792 3947 796
rect 1639 783 1643 787
rect 331 775 335 779
rect 615 775 619 779
rect 879 771 883 775
rect 1095 775 1099 779
rect 1167 775 1171 779
rect 1463 771 1467 775
rect 1675 771 1679 775
rect 2047 775 2051 779
rect 2291 779 2295 783
rect 2403 779 2407 783
rect 2523 779 2527 783
rect 2659 779 2663 783
rect 2811 779 2815 783
rect 2971 783 2975 787
rect 3323 779 3327 783
rect 3331 783 3335 787
rect 3531 783 3535 787
rect 3915 783 3919 787
rect 2215 772 2219 776
rect 2327 772 2331 776
rect 2447 772 2451 776
rect 2583 772 2587 776
rect 2735 772 2739 776
rect 2895 772 2899 776
rect 3063 772 3067 776
rect 3247 772 3251 776
rect 3447 772 3451 776
rect 3655 772 3659 776
rect 3839 772 3843 776
rect 3943 775 3947 779
rect 451 759 455 763
rect 571 759 575 763
rect 819 759 823 763
rect 1079 759 1080 763
rect 1080 759 1083 763
rect 1099 759 1103 763
rect 1367 759 1368 763
rect 1368 759 1371 763
rect 1387 759 1391 763
rect 699 751 703 755
rect 2351 759 2355 763
rect 2291 751 2295 755
rect 2403 751 2407 755
rect 2523 751 2527 755
rect 2659 751 2663 755
rect 3131 747 3135 751
rect 3331 751 3335 755
rect 3531 751 3535 755
rect 3691 751 3695 755
rect 3907 747 3911 751
rect 111 733 115 737
rect 375 736 379 740
rect 495 736 499 740
rect 623 736 627 740
rect 451 727 455 731
rect 571 727 575 731
rect 699 727 703 731
rect 751 736 755 740
rect 887 736 891 740
rect 1023 736 1027 740
rect 1167 736 1171 740
rect 1311 736 1315 740
rect 1455 736 1459 740
rect 1599 736 1603 740
rect 2007 733 2011 737
rect 879 727 883 731
rect 1099 727 1103 731
rect 1235 727 1239 731
rect 1387 727 1391 731
rect 1675 727 1679 731
rect 2467 731 2471 735
rect 2811 731 2815 735
rect 2843 731 2847 735
rect 3119 731 3120 735
rect 3120 731 3123 735
rect 3323 731 3327 735
rect 3595 731 3599 735
rect 3895 731 3896 735
rect 3896 731 3899 735
rect 2591 723 2595 727
rect 2883 723 2887 727
rect 111 716 115 720
rect 375 717 379 721
rect 495 717 499 721
rect 623 717 627 721
rect 751 717 755 721
rect 887 717 891 721
rect 1023 717 1027 721
rect 1167 717 1171 721
rect 1311 717 1315 721
rect 1455 717 1459 721
rect 1599 717 1603 721
rect 2007 716 2011 720
rect 2047 705 2051 709
rect 2375 708 2379 712
rect 2495 708 2499 712
rect 2623 708 2627 712
rect 2767 708 2771 712
rect 2911 708 2915 712
rect 3063 708 3067 712
rect 3215 708 3219 712
rect 3367 708 3371 712
rect 3519 708 3523 712
rect 3679 708 3683 712
rect 3839 708 3843 712
rect 3943 705 3947 709
rect 2467 699 2471 703
rect 2583 699 2587 703
rect 2591 699 2595 703
rect 2843 699 2847 703
rect 2883 699 2887 703
rect 3131 699 3135 703
rect 3595 699 3599 703
rect 3747 699 3751 703
rect 3907 699 3911 703
rect 2047 688 2051 692
rect 2375 689 2379 693
rect 2495 689 2499 693
rect 2623 689 2627 693
rect 2767 689 2771 693
rect 2911 689 2915 693
rect 3063 689 3067 693
rect 3215 689 3219 693
rect 3367 689 3371 693
rect 3519 689 3523 693
rect 3679 689 3683 693
rect 3839 689 3843 693
rect 3943 688 3947 692
rect 111 664 115 668
rect 527 663 531 667
rect 631 663 635 667
rect 743 663 747 667
rect 855 663 859 667
rect 967 663 971 667
rect 1071 663 1075 667
rect 1183 663 1187 667
rect 1295 663 1299 667
rect 1407 663 1411 667
rect 1519 663 1523 667
rect 2007 664 2011 668
rect 111 647 115 651
rect 603 651 607 655
rect 707 651 711 655
rect 819 655 823 659
rect 827 655 831 659
rect 1147 651 1151 655
rect 1371 655 1375 659
rect 1383 655 1387 659
rect 1491 655 1495 659
rect 527 644 531 648
rect 631 644 635 648
rect 743 644 747 648
rect 855 644 859 648
rect 967 644 971 648
rect 1071 644 1075 648
rect 1183 644 1187 648
rect 1295 644 1299 648
rect 1407 644 1411 648
rect 1519 644 1523 648
rect 2007 647 2011 651
rect 827 631 831 635
rect 2047 628 2051 632
rect 603 623 607 627
rect 707 623 711 627
rect 1235 623 1236 627
rect 1236 623 1239 627
rect 1383 623 1387 627
rect 2111 627 2115 631
rect 1491 623 1495 627
rect 2247 627 2251 631
rect 2399 627 2403 631
rect 2575 627 2579 631
rect 2759 627 2763 631
rect 2943 627 2947 631
rect 3127 627 3131 631
rect 3303 627 3307 631
rect 3479 627 3483 631
rect 3655 627 3659 631
rect 3831 627 3835 631
rect 3943 628 3947 632
rect 1531 619 1535 623
rect 2195 619 2199 623
rect 763 607 767 611
rect 1059 607 1063 611
rect 1147 607 1151 611
rect 1243 607 1247 611
rect 1339 607 1343 611
rect 1435 607 1439 611
rect 2047 611 2051 615
rect 2651 615 2655 619
rect 2659 619 2663 623
rect 3019 615 3023 619
rect 3119 619 3123 623
rect 3379 615 3383 619
rect 3391 619 3395 623
rect 3599 619 3603 623
rect 3899 623 3903 627
rect 2111 608 2115 612
rect 2247 608 2251 612
rect 2399 608 2403 612
rect 2575 608 2579 612
rect 2759 608 2763 612
rect 2943 608 2947 612
rect 3127 608 3131 612
rect 3303 608 3307 612
rect 3479 608 3483 612
rect 3655 608 3659 612
rect 3831 608 3835 612
rect 3943 611 3947 615
rect 1043 599 1047 603
rect 1331 599 1335 603
rect 111 581 115 585
rect 687 584 691 588
rect 783 584 787 588
rect 879 584 883 588
rect 975 584 979 588
rect 1071 584 1075 588
rect 1167 584 1171 588
rect 1263 584 1267 588
rect 1359 584 1363 588
rect 1455 584 1459 588
rect 2195 587 2199 591
rect 2659 595 2663 599
rect 2583 587 2587 591
rect 2651 587 2655 591
rect 2007 581 2011 585
rect 2955 583 2959 587
rect 3019 587 3023 591
rect 3391 587 3395 591
rect 3599 587 3603 591
rect 3747 587 3751 591
rect 3907 583 3911 587
rect 763 575 767 579
rect 1043 575 1047 579
rect 1059 575 1063 579
rect 1243 575 1247 579
rect 1339 575 1343 579
rect 1435 575 1439 579
rect 1531 575 1535 579
rect 111 564 115 568
rect 687 565 691 569
rect 783 565 787 569
rect 879 565 883 569
rect 975 565 979 569
rect 1071 565 1075 569
rect 1167 565 1171 569
rect 1263 565 1267 569
rect 1359 565 1363 569
rect 1455 565 1459 569
rect 2007 564 2011 568
rect 2147 567 2151 571
rect 2259 567 2263 571
rect 2411 567 2415 571
rect 2963 567 2967 571
rect 3175 567 3179 571
rect 3235 567 3239 571
rect 3379 567 3383 571
rect 3531 567 3535 571
rect 3723 567 3727 571
rect 2047 541 2051 545
rect 2071 544 2075 548
rect 2183 544 2187 548
rect 2335 544 2339 548
rect 2503 544 2507 548
rect 2687 544 2691 548
rect 2879 544 2883 548
rect 3071 544 3075 548
rect 3263 544 3267 548
rect 3455 544 3459 548
rect 3647 544 3651 548
rect 3839 544 3843 548
rect 3943 541 3947 545
rect 2147 535 2151 539
rect 2259 535 2263 539
rect 2411 535 2415 539
rect 2659 535 2663 539
rect 2955 535 2959 539
rect 2963 535 2967 539
rect 3175 535 3179 539
rect 3531 535 3535 539
rect 3723 535 3727 539
rect 3907 535 3911 539
rect 2047 524 2051 528
rect 2071 525 2075 529
rect 2183 525 2187 529
rect 2335 525 2339 529
rect 2503 525 2507 529
rect 2687 525 2691 529
rect 2879 525 2883 529
rect 3071 525 3075 529
rect 3263 525 3267 529
rect 3455 525 3459 529
rect 3647 525 3651 529
rect 3839 525 3843 529
rect 3943 524 3947 528
rect 111 492 115 496
rect 383 491 387 495
rect 479 491 483 495
rect 575 491 579 495
rect 671 491 675 495
rect 767 491 771 495
rect 863 491 867 495
rect 959 491 963 495
rect 1055 491 1059 495
rect 1151 491 1155 495
rect 1247 491 1251 495
rect 1343 491 1347 495
rect 1439 491 1443 495
rect 1535 491 1539 495
rect 2007 492 2011 496
rect 111 475 115 479
rect 459 479 463 483
rect 555 479 559 483
rect 651 479 655 483
rect 747 479 751 483
rect 843 479 847 483
rect 939 479 943 483
rect 1035 479 1039 483
rect 1131 479 1135 483
rect 1227 479 1231 483
rect 1331 483 1335 487
rect 1515 479 1519 483
rect 383 472 387 476
rect 479 472 483 476
rect 575 472 579 476
rect 671 472 675 476
rect 767 472 771 476
rect 863 472 867 476
rect 959 472 963 476
rect 1055 472 1059 476
rect 1151 472 1155 476
rect 1247 472 1251 476
rect 1343 472 1347 476
rect 1439 472 1443 476
rect 1535 472 1539 476
rect 2007 475 2011 479
rect 2047 472 2051 476
rect 2183 471 2187 475
rect 2319 471 2323 475
rect 2463 471 2467 475
rect 2615 471 2619 475
rect 2775 471 2779 475
rect 2959 471 2963 475
rect 3159 471 3163 475
rect 3367 471 3371 475
rect 3583 471 3587 475
rect 3807 471 3811 475
rect 3943 472 3947 476
rect 459 451 463 455
rect 555 451 559 455
rect 651 451 655 455
rect 747 451 751 455
rect 843 451 847 455
rect 939 451 943 455
rect 1035 451 1039 455
rect 1131 451 1135 455
rect 1227 451 1231 455
rect 967 443 971 447
rect 1495 447 1496 451
rect 1496 447 1499 451
rect 1515 451 1519 455
rect 2047 455 2051 459
rect 2259 459 2263 463
rect 2395 459 2399 463
rect 2539 459 2543 463
rect 2691 459 2695 463
rect 2699 463 2703 467
rect 3035 459 3039 463
rect 3235 463 3239 467
rect 3243 463 3247 467
rect 3767 463 3771 467
rect 2183 452 2187 456
rect 2319 452 2323 456
rect 2463 452 2467 456
rect 2615 452 2619 456
rect 2775 452 2779 456
rect 2959 452 2963 456
rect 3159 452 3163 456
rect 3367 452 3371 456
rect 3583 452 3587 456
rect 3807 452 3811 456
rect 3943 455 3947 459
rect 2659 439 2663 443
rect 2259 431 2263 435
rect 2395 431 2399 435
rect 2539 431 2543 435
rect 2691 431 2695 435
rect 3243 439 3247 443
rect 3035 431 3039 435
rect 539 421 540 423
rect 540 421 543 423
rect 563 423 567 427
rect 659 423 663 427
rect 1187 423 1191 427
rect 1419 423 1423 427
rect 539 419 543 421
rect 2699 423 2703 427
rect 3491 427 3495 431
rect 3907 427 3911 431
rect 1395 415 1399 419
rect 2419 415 2423 419
rect 2563 415 2567 419
rect 2715 415 2719 419
rect 2875 415 2879 419
rect 3187 415 3191 419
rect 3339 415 3343 419
rect 3647 415 3651 419
rect 3787 415 3791 419
rect 3915 415 3919 419
rect 3499 407 3503 411
rect 111 397 115 401
rect 487 400 491 404
rect 583 400 587 404
rect 687 400 691 404
rect 791 400 795 404
rect 895 400 899 404
rect 999 400 1003 404
rect 1103 400 1107 404
rect 1207 400 1211 404
rect 1319 400 1323 404
rect 1431 400 1435 404
rect 2007 397 2011 401
rect 563 391 567 395
rect 659 391 663 395
rect 967 391 971 395
rect 1075 391 1079 395
rect 1187 391 1191 395
rect 1395 391 1399 395
rect 1499 391 1503 395
rect 2047 389 2051 393
rect 2343 392 2347 396
rect 2487 392 2491 396
rect 2639 392 2643 396
rect 2799 392 2803 396
rect 2959 392 2963 396
rect 3111 392 3115 396
rect 3263 392 3267 396
rect 3415 392 3419 396
rect 3559 392 3563 396
rect 3711 392 3715 396
rect 3839 392 3843 396
rect 3943 389 3947 393
rect 111 380 115 384
rect 487 381 491 385
rect 583 381 587 385
rect 687 381 691 385
rect 791 381 795 385
rect 895 381 899 385
rect 999 381 1003 385
rect 1103 381 1107 385
rect 1207 381 1211 385
rect 1319 381 1323 385
rect 1431 381 1435 385
rect 2007 380 2011 384
rect 2419 383 2423 387
rect 2563 383 2567 387
rect 2715 383 2719 387
rect 2875 383 2879 387
rect 2899 383 2903 387
rect 3187 383 3191 387
rect 3339 383 3343 387
rect 3491 383 3495 387
rect 3499 383 3503 387
rect 3647 383 3651 387
rect 3907 383 3911 387
rect 2047 372 2051 376
rect 2343 373 2347 377
rect 2487 373 2491 377
rect 2639 373 2643 377
rect 2799 373 2803 377
rect 2959 373 2963 377
rect 3111 373 3115 377
rect 3263 373 3267 377
rect 3415 373 3419 377
rect 3559 373 3563 377
rect 3711 373 3715 377
rect 3839 373 3843 377
rect 3943 372 3947 376
rect 111 324 115 328
rect 327 323 331 327
rect 463 323 467 327
rect 615 323 619 327
rect 767 323 771 327
rect 919 323 923 327
rect 1063 323 1067 327
rect 1207 323 1211 327
rect 1351 323 1355 327
rect 111 307 115 311
rect 403 311 407 315
rect 539 311 543 315
rect 691 311 695 315
rect 843 311 847 315
rect 859 315 863 319
rect 1419 319 1423 323
rect 1495 323 1499 327
rect 1639 323 1643 327
rect 2007 324 2011 328
rect 1139 311 1143 315
rect 1283 311 1287 315
rect 1435 315 1439 319
rect 1579 315 1583 319
rect 2047 316 2051 320
rect 2495 315 2499 319
rect 2639 315 2643 319
rect 2799 315 2803 319
rect 2959 315 2963 319
rect 3119 315 3123 319
rect 3271 315 3275 319
rect 3423 315 3427 319
rect 3567 315 3571 319
rect 3711 315 3715 319
rect 3839 315 3843 319
rect 3943 316 3947 320
rect 327 304 331 308
rect 463 304 467 308
rect 615 304 619 308
rect 767 304 771 308
rect 919 304 923 308
rect 1063 304 1067 308
rect 1207 304 1211 308
rect 1351 304 1355 308
rect 1495 304 1499 308
rect 1639 304 1643 308
rect 2007 307 2011 311
rect 2047 299 2051 303
rect 2571 303 2575 307
rect 2715 303 2719 307
rect 2875 303 2879 307
rect 3035 303 3039 307
rect 3043 307 3047 311
rect 3347 303 3351 307
rect 3499 303 3503 307
rect 3643 303 3647 307
rect 3787 307 3791 311
rect 3915 307 3919 311
rect 2495 296 2499 300
rect 2639 296 2643 300
rect 2799 296 2803 300
rect 2959 296 2963 300
rect 3119 296 3123 300
rect 3271 296 3275 300
rect 3423 296 3427 300
rect 3567 296 3571 300
rect 3711 296 3715 300
rect 3839 296 3843 300
rect 3943 299 3947 303
rect 403 283 407 287
rect 539 283 543 287
rect 691 283 695 287
rect 843 283 847 287
rect 1075 283 1079 287
rect 1139 283 1143 287
rect 1435 283 1439 287
rect 1579 283 1583 287
rect 1587 279 1591 283
rect 2551 275 2552 279
rect 2552 275 2555 279
rect 2571 275 2575 279
rect 2715 275 2719 279
rect 2875 275 2879 279
rect 3035 275 3039 279
rect 3347 275 3351 279
rect 3499 275 3503 279
rect 3767 275 3768 279
rect 3768 275 3771 279
rect 3619 267 3623 271
rect 3907 271 3911 275
rect 243 259 247 263
rect 403 259 407 263
rect 579 259 583 263
rect 1283 259 1287 263
rect 1291 259 1295 263
rect 1595 259 1599 263
rect 1731 259 1735 263
rect 1867 259 1871 263
rect 1987 259 1991 263
rect 2155 259 2159 263
rect 2539 259 2543 263
rect 2579 259 2583 263
rect 3043 259 3047 263
rect 3171 259 3175 263
rect 3363 259 3367 263
rect 3555 259 3559 263
rect 3915 259 3919 263
rect 859 247 863 251
rect 1339 251 1343 255
rect 3499 251 3503 255
rect 111 233 115 237
rect 167 236 171 240
rect 327 236 331 240
rect 503 236 507 240
rect 687 236 691 240
rect 871 236 875 240
rect 1047 236 1051 240
rect 1215 236 1219 240
rect 1367 236 1371 240
rect 1511 236 1515 240
rect 1647 236 1651 240
rect 1783 236 1787 240
rect 1903 236 1907 240
rect 2007 233 2011 237
rect 2047 233 2051 237
rect 2071 236 2075 240
rect 2271 236 2275 240
rect 2495 236 2499 240
rect 2703 236 2707 240
rect 2903 236 2907 240
rect 3095 236 3099 240
rect 3287 236 3291 240
rect 3479 236 3483 240
rect 3671 236 3675 240
rect 3839 236 3843 240
rect 3943 233 3947 237
rect 243 227 247 231
rect 403 227 407 231
rect 579 227 583 231
rect 1115 227 1119 231
rect 1291 227 1295 231
rect 1339 227 1343 231
rect 1587 227 1591 231
rect 1595 227 1599 231
rect 1731 227 1735 231
rect 1867 227 1871 231
rect 1987 227 1991 231
rect 2155 227 2159 231
rect 2579 227 2583 231
rect 3171 227 3175 231
rect 3363 227 3367 231
rect 3555 227 3559 231
rect 3619 227 3623 231
rect 3907 227 3911 231
rect 111 216 115 220
rect 167 217 171 221
rect 327 217 331 221
rect 503 217 507 221
rect 687 217 691 221
rect 871 217 875 221
rect 1047 217 1051 221
rect 1215 217 1219 221
rect 1367 217 1371 221
rect 1511 217 1515 221
rect 1647 217 1651 221
rect 1783 217 1787 221
rect 1903 217 1907 221
rect 2007 216 2011 220
rect 2047 216 2051 220
rect 2071 217 2075 221
rect 2271 217 2275 221
rect 2495 217 2499 221
rect 2615 219 2619 223
rect 2703 217 2707 221
rect 2903 217 2907 221
rect 3095 217 3099 221
rect 3287 217 3291 221
rect 3479 217 3483 221
rect 3671 217 3675 221
rect 3839 217 3843 221
rect 3943 216 3947 220
rect 111 136 115 140
rect 135 135 139 139
rect 231 135 235 139
rect 327 135 331 139
rect 423 135 427 139
rect 527 135 531 139
rect 647 135 651 139
rect 775 135 779 139
rect 903 135 907 139
rect 1031 135 1035 139
rect 1151 135 1155 139
rect 1271 135 1275 139
rect 1383 135 1387 139
rect 1487 135 1491 139
rect 1591 135 1595 139
rect 1703 135 1707 139
rect 1807 135 1811 139
rect 1903 135 1907 139
rect 2007 136 2011 140
rect 2047 140 2051 144
rect 2071 139 2075 143
rect 2167 139 2171 143
rect 2263 139 2267 143
rect 2359 139 2363 143
rect 2455 139 2459 143
rect 2551 139 2555 143
rect 2655 139 2659 143
rect 2759 139 2763 143
rect 2863 139 2867 143
rect 2975 139 2979 143
rect 3103 139 3107 143
rect 3239 139 3243 143
rect 3383 139 3387 143
rect 3535 139 3539 143
rect 3695 139 3699 143
rect 3839 139 3843 143
rect 3943 140 3947 144
rect 111 119 115 123
rect 211 123 215 127
rect 307 123 311 127
rect 403 123 407 127
rect 499 123 503 127
rect 603 123 607 127
rect 723 123 727 127
rect 851 123 855 127
rect 859 127 863 131
rect 1123 123 1127 127
rect 1227 123 1231 127
rect 1347 123 1351 127
rect 1459 123 1463 127
rect 1563 123 1567 127
rect 1667 123 1671 127
rect 1779 123 1783 127
rect 1883 123 1887 127
rect 1979 123 1983 127
rect 135 116 139 120
rect 231 116 235 120
rect 327 116 331 120
rect 423 116 427 120
rect 527 116 531 120
rect 647 116 651 120
rect 775 116 779 120
rect 903 116 907 120
rect 1031 116 1035 120
rect 1151 116 1155 120
rect 1271 116 1275 120
rect 1383 116 1387 120
rect 1487 116 1491 120
rect 1591 116 1595 120
rect 1703 116 1707 120
rect 1807 116 1811 120
rect 1903 116 1907 120
rect 2007 119 2011 123
rect 2047 123 2051 127
rect 2147 127 2151 131
rect 2243 127 2247 131
rect 2339 127 2343 131
rect 2435 127 2439 131
rect 2531 127 2535 131
rect 2539 131 2543 135
rect 2731 127 2735 131
rect 2835 127 2839 131
rect 2939 127 2943 131
rect 3051 127 3055 131
rect 3179 127 3183 131
rect 3315 127 3319 131
rect 3459 127 3463 131
rect 3499 131 3503 135
rect 3771 127 3775 131
rect 3915 131 3919 135
rect 2071 120 2075 124
rect 2167 120 2171 124
rect 2263 120 2267 124
rect 2359 120 2363 124
rect 2455 120 2459 124
rect 2551 120 2555 124
rect 2655 120 2659 124
rect 2759 120 2763 124
rect 2863 120 2867 124
rect 2975 120 2979 124
rect 3103 120 3107 124
rect 3239 120 3243 124
rect 3383 120 3387 124
rect 3535 120 3539 124
rect 3695 120 3699 124
rect 3839 120 3843 124
rect 3943 123 3947 127
rect 211 95 215 99
rect 307 95 311 99
rect 403 95 407 99
rect 499 95 503 99
rect 603 95 607 99
rect 723 95 727 99
rect 851 95 855 99
rect 1115 95 1119 99
rect 1123 95 1127 99
rect 1227 95 1231 99
rect 1347 95 1351 99
rect 1459 95 1463 99
rect 1563 95 1567 99
rect 1667 95 1671 99
rect 1779 95 1783 99
rect 1883 95 1887 99
rect 1979 99 1983 103
rect 2147 99 2151 103
rect 2243 99 2247 103
rect 2339 99 2343 103
rect 2435 99 2439 103
rect 2531 99 2535 103
rect 2615 99 2619 103
rect 2731 99 2735 103
rect 2835 99 2839 103
rect 2939 99 2943 103
rect 3051 99 3055 103
rect 3179 99 3183 103
rect 3315 99 3319 103
rect 3459 99 3463 103
rect 3643 99 3647 103
rect 3771 99 3775 103
<< m3 >>
rect 111 4030 115 4031
rect 111 4025 115 4026
rect 1519 4030 1523 4031
rect 1519 4025 1523 4026
rect 1615 4030 1619 4031
rect 1615 4025 1619 4026
rect 1711 4030 1715 4031
rect 1711 4025 1715 4026
rect 1807 4030 1811 4031
rect 1807 4025 1811 4026
rect 1903 4030 1907 4031
rect 1903 4025 1907 4026
rect 2007 4030 2011 4031
rect 2007 4025 2011 4026
rect 112 4005 114 4025
rect 110 4004 116 4005
rect 1520 4004 1522 4025
rect 1616 4004 1618 4025
rect 1712 4004 1714 4025
rect 1808 4004 1810 4025
rect 1904 4004 1906 4025
rect 2008 4005 2010 4025
rect 2047 4018 2051 4019
rect 2047 4013 2051 4014
rect 2071 4018 2075 4019
rect 2071 4013 2075 4014
rect 2167 4018 2171 4019
rect 2167 4013 2171 4014
rect 2263 4018 2267 4019
rect 2263 4013 2267 4014
rect 3943 4018 3947 4019
rect 3943 4013 3947 4014
rect 2006 4004 2012 4005
rect 110 4000 111 4004
rect 115 4000 116 4004
rect 110 3999 116 4000
rect 1518 4003 1524 4004
rect 1518 3999 1519 4003
rect 1523 3999 1524 4003
rect 1518 3998 1524 3999
rect 1614 4003 1620 4004
rect 1614 3999 1615 4003
rect 1619 3999 1620 4003
rect 1614 3998 1620 3999
rect 1710 4003 1716 4004
rect 1710 3999 1711 4003
rect 1715 3999 1716 4003
rect 1710 3998 1716 3999
rect 1806 4003 1812 4004
rect 1806 3999 1807 4003
rect 1811 3999 1812 4003
rect 1806 3998 1812 3999
rect 1902 4003 1908 4004
rect 1902 3999 1903 4003
rect 1907 3999 1908 4003
rect 2006 4000 2007 4004
rect 2011 4000 2012 4004
rect 2006 3999 2012 4000
rect 1902 3998 1908 3999
rect 1690 3991 1696 3992
rect 110 3987 116 3988
rect 110 3983 111 3987
rect 115 3983 116 3987
rect 1690 3987 1691 3991
rect 1695 3987 1696 3991
rect 1690 3986 1696 3987
rect 1786 3991 1792 3992
rect 1786 3987 1787 3991
rect 1791 3987 1792 3991
rect 1786 3986 1792 3987
rect 1882 3991 1888 3992
rect 1882 3987 1883 3991
rect 1887 3987 1888 3991
rect 1882 3986 1888 3987
rect 2006 3987 2012 3988
rect 110 3982 116 3983
rect 1518 3984 1524 3985
rect 112 3955 114 3982
rect 1518 3980 1519 3984
rect 1523 3980 1524 3984
rect 1518 3979 1524 3980
rect 1614 3984 1620 3985
rect 1614 3980 1615 3984
rect 1619 3980 1620 3984
rect 1614 3979 1620 3980
rect 1520 3955 1522 3979
rect 1616 3955 1618 3979
rect 1692 3964 1694 3986
rect 1710 3984 1716 3985
rect 1710 3980 1711 3984
rect 1715 3980 1716 3984
rect 1710 3979 1716 3980
rect 1690 3963 1696 3964
rect 1690 3959 1691 3963
rect 1695 3959 1696 3963
rect 1690 3958 1696 3959
rect 1712 3955 1714 3979
rect 1788 3964 1790 3986
rect 1806 3984 1812 3985
rect 1806 3980 1807 3984
rect 1811 3980 1812 3984
rect 1806 3979 1812 3980
rect 1786 3963 1792 3964
rect 1786 3959 1787 3963
rect 1791 3959 1792 3963
rect 1786 3958 1792 3959
rect 1808 3955 1810 3979
rect 1884 3964 1886 3986
rect 1902 3984 1908 3985
rect 1902 3980 1903 3984
rect 1907 3980 1908 3984
rect 2006 3983 2007 3987
rect 2011 3983 2012 3987
rect 2048 3986 2050 4013
rect 2072 3989 2074 4013
rect 2146 4011 2152 4012
rect 2146 4007 2147 4011
rect 2151 4007 2152 4011
rect 2146 4006 2152 4007
rect 2070 3988 2076 3989
rect 2006 3982 2012 3983
rect 2046 3985 2052 3986
rect 1902 3979 1908 3980
rect 1882 3963 1888 3964
rect 1882 3959 1883 3963
rect 1887 3959 1888 3963
rect 1882 3958 1888 3959
rect 1904 3955 1906 3979
rect 2008 3955 2010 3982
rect 2046 3981 2047 3985
rect 2051 3981 2052 3985
rect 2070 3984 2071 3988
rect 2075 3984 2076 3988
rect 2070 3983 2076 3984
rect 2046 3980 2052 3981
rect 2148 3980 2150 4006
rect 2168 3989 2170 4013
rect 2242 4011 2248 4012
rect 2242 4007 2243 4011
rect 2247 4007 2248 4011
rect 2242 4006 2248 4007
rect 2166 3988 2172 3989
rect 2166 3984 2167 3988
rect 2171 3984 2172 3988
rect 2166 3983 2172 3984
rect 2244 3980 2246 4006
rect 2264 3989 2266 4013
rect 2262 3988 2268 3989
rect 2262 3984 2263 3988
rect 2267 3984 2268 3988
rect 3944 3986 3946 4013
rect 2262 3983 2268 3984
rect 3942 3985 3948 3986
rect 3942 3981 3943 3985
rect 3947 3981 3948 3985
rect 3942 3980 3948 3981
rect 2146 3979 2152 3980
rect 2146 3975 2147 3979
rect 2151 3975 2152 3979
rect 2146 3974 2152 3975
rect 2242 3979 2248 3980
rect 2242 3975 2243 3979
rect 2247 3975 2248 3979
rect 2242 3974 2248 3975
rect 2070 3969 2076 3970
rect 2046 3968 2052 3969
rect 2046 3964 2047 3968
rect 2051 3964 2052 3968
rect 2070 3965 2071 3969
rect 2075 3965 2076 3969
rect 2070 3964 2076 3965
rect 2166 3969 2172 3970
rect 2166 3965 2167 3969
rect 2171 3965 2172 3969
rect 2166 3964 2172 3965
rect 2262 3969 2268 3970
rect 2262 3965 2263 3969
rect 2267 3965 2268 3969
rect 2262 3964 2268 3965
rect 3942 3968 3948 3969
rect 3942 3964 3943 3968
rect 3947 3964 3948 3968
rect 2046 3963 2052 3964
rect 111 3954 115 3955
rect 111 3949 115 3950
rect 199 3954 203 3955
rect 199 3949 203 3950
rect 295 3954 299 3955
rect 295 3949 299 3950
rect 391 3954 395 3955
rect 391 3949 395 3950
rect 495 3954 499 3955
rect 495 3949 499 3950
rect 615 3954 619 3955
rect 615 3949 619 3950
rect 743 3954 747 3955
rect 743 3949 747 3950
rect 871 3954 875 3955
rect 871 3949 875 3950
rect 999 3954 1003 3955
rect 999 3949 1003 3950
rect 1127 3954 1131 3955
rect 1127 3949 1131 3950
rect 1255 3954 1259 3955
rect 1255 3949 1259 3950
rect 1383 3954 1387 3955
rect 1383 3949 1387 3950
rect 1511 3954 1515 3955
rect 1511 3949 1515 3950
rect 1519 3954 1523 3955
rect 1519 3949 1523 3950
rect 1615 3954 1619 3955
rect 1615 3949 1619 3950
rect 1647 3954 1651 3955
rect 1647 3949 1651 3950
rect 1711 3954 1715 3955
rect 1711 3949 1715 3950
rect 1807 3954 1811 3955
rect 1807 3949 1811 3950
rect 1903 3954 1907 3955
rect 1903 3949 1907 3950
rect 2007 3954 2011 3955
rect 2007 3949 2011 3950
rect 112 3922 114 3949
rect 200 3925 202 3949
rect 266 3947 272 3948
rect 266 3943 267 3947
rect 271 3943 272 3947
rect 266 3942 272 3943
rect 274 3947 280 3948
rect 274 3943 275 3947
rect 279 3943 280 3947
rect 274 3942 280 3943
rect 198 3924 204 3925
rect 110 3921 116 3922
rect 110 3917 111 3921
rect 115 3917 116 3921
rect 198 3920 199 3924
rect 203 3920 204 3924
rect 198 3919 204 3920
rect 110 3916 116 3917
rect 198 3905 204 3906
rect 110 3904 116 3905
rect 110 3900 111 3904
rect 115 3900 116 3904
rect 198 3901 199 3905
rect 203 3901 204 3905
rect 198 3900 204 3901
rect 110 3899 116 3900
rect 112 3879 114 3899
rect 200 3879 202 3900
rect 111 3878 115 3879
rect 111 3873 115 3874
rect 199 3878 203 3879
rect 199 3873 203 3874
rect 112 3853 114 3873
rect 110 3852 116 3853
rect 110 3848 111 3852
rect 115 3848 116 3852
rect 110 3847 116 3848
rect 268 3844 270 3942
rect 276 3916 278 3942
rect 296 3925 298 3949
rect 370 3947 376 3948
rect 370 3943 371 3947
rect 375 3943 376 3947
rect 370 3942 376 3943
rect 294 3924 300 3925
rect 294 3920 295 3924
rect 299 3920 300 3924
rect 294 3919 300 3920
rect 372 3916 374 3942
rect 392 3925 394 3949
rect 466 3947 472 3948
rect 466 3943 467 3947
rect 471 3943 472 3947
rect 466 3942 472 3943
rect 390 3924 396 3925
rect 390 3920 391 3924
rect 395 3920 396 3924
rect 390 3919 396 3920
rect 468 3916 470 3942
rect 496 3925 498 3949
rect 570 3947 576 3948
rect 570 3943 571 3947
rect 575 3943 576 3947
rect 570 3942 576 3943
rect 494 3924 500 3925
rect 494 3920 495 3924
rect 499 3920 500 3924
rect 494 3919 500 3920
rect 572 3916 574 3942
rect 616 3925 618 3949
rect 690 3947 696 3948
rect 690 3943 691 3947
rect 695 3943 696 3947
rect 690 3942 696 3943
rect 614 3924 620 3925
rect 614 3920 615 3924
rect 619 3920 620 3924
rect 614 3919 620 3920
rect 692 3916 694 3942
rect 744 3925 746 3949
rect 818 3947 824 3948
rect 818 3943 819 3947
rect 823 3943 824 3947
rect 818 3942 824 3943
rect 742 3924 748 3925
rect 742 3920 743 3924
rect 747 3920 748 3924
rect 742 3919 748 3920
rect 820 3916 822 3942
rect 872 3925 874 3949
rect 946 3947 952 3948
rect 946 3943 947 3947
rect 951 3943 952 3947
rect 946 3942 952 3943
rect 870 3924 876 3925
rect 870 3920 871 3924
rect 875 3920 876 3924
rect 870 3919 876 3920
rect 948 3916 950 3942
rect 1000 3925 1002 3949
rect 1128 3925 1130 3949
rect 1178 3947 1184 3948
rect 1178 3943 1179 3947
rect 1183 3943 1184 3947
rect 1178 3942 1184 3943
rect 1202 3947 1208 3948
rect 1202 3943 1203 3947
rect 1207 3943 1208 3947
rect 1202 3942 1208 3943
rect 998 3924 1004 3925
rect 998 3920 999 3924
rect 1003 3920 1004 3924
rect 998 3919 1004 3920
rect 1126 3924 1132 3925
rect 1126 3920 1127 3924
rect 1131 3920 1132 3924
rect 1126 3919 1132 3920
rect 274 3915 280 3916
rect 274 3911 275 3915
rect 279 3911 280 3915
rect 274 3910 280 3911
rect 370 3915 376 3916
rect 370 3911 371 3915
rect 375 3911 376 3915
rect 370 3910 376 3911
rect 466 3915 472 3916
rect 466 3911 467 3915
rect 471 3911 472 3915
rect 466 3910 472 3911
rect 570 3915 576 3916
rect 570 3911 571 3915
rect 575 3911 576 3915
rect 570 3910 576 3911
rect 690 3915 696 3916
rect 690 3911 691 3915
rect 695 3911 696 3915
rect 690 3910 696 3911
rect 818 3915 824 3916
rect 818 3911 819 3915
rect 823 3911 824 3915
rect 818 3910 824 3911
rect 946 3915 952 3916
rect 946 3911 947 3915
rect 951 3911 952 3915
rect 946 3910 952 3911
rect 954 3915 960 3916
rect 954 3911 955 3915
rect 959 3911 960 3915
rect 954 3910 960 3911
rect 294 3905 300 3906
rect 294 3901 295 3905
rect 299 3901 300 3905
rect 294 3900 300 3901
rect 390 3905 396 3906
rect 390 3901 391 3905
rect 395 3901 396 3905
rect 390 3900 396 3901
rect 494 3905 500 3906
rect 494 3901 495 3905
rect 499 3901 500 3905
rect 494 3900 500 3901
rect 614 3905 620 3906
rect 614 3901 615 3905
rect 619 3901 620 3905
rect 614 3900 620 3901
rect 742 3905 748 3906
rect 742 3901 743 3905
rect 747 3901 748 3905
rect 742 3900 748 3901
rect 870 3905 876 3906
rect 870 3901 871 3905
rect 875 3901 876 3905
rect 870 3900 876 3901
rect 296 3879 298 3900
rect 392 3879 394 3900
rect 496 3879 498 3900
rect 616 3879 618 3900
rect 744 3879 746 3900
rect 872 3879 874 3900
rect 295 3878 299 3879
rect 295 3873 299 3874
rect 335 3878 339 3879
rect 335 3873 339 3874
rect 391 3878 395 3879
rect 391 3873 395 3874
rect 455 3878 459 3879
rect 455 3873 459 3874
rect 495 3878 499 3879
rect 495 3873 499 3874
rect 583 3878 587 3879
rect 583 3873 587 3874
rect 615 3878 619 3879
rect 615 3873 619 3874
rect 719 3878 723 3879
rect 719 3873 723 3874
rect 743 3878 747 3879
rect 743 3873 747 3874
rect 847 3878 851 3879
rect 847 3873 851 3874
rect 871 3878 875 3879
rect 871 3873 875 3874
rect 336 3852 338 3873
rect 456 3852 458 3873
rect 584 3852 586 3873
rect 720 3852 722 3873
rect 848 3852 850 3873
rect 334 3851 340 3852
rect 334 3847 335 3851
rect 339 3847 340 3851
rect 334 3846 340 3847
rect 454 3851 460 3852
rect 454 3847 455 3851
rect 459 3847 460 3851
rect 454 3846 460 3847
rect 582 3851 588 3852
rect 582 3847 583 3851
rect 587 3847 588 3851
rect 582 3846 588 3847
rect 718 3851 724 3852
rect 718 3847 719 3851
rect 723 3847 724 3851
rect 718 3846 724 3847
rect 846 3851 852 3852
rect 846 3847 847 3851
rect 851 3847 852 3851
rect 846 3846 852 3847
rect 266 3843 272 3844
rect 266 3839 267 3843
rect 271 3839 272 3843
rect 266 3838 272 3839
rect 794 3839 800 3840
rect 110 3835 116 3836
rect 110 3831 111 3835
rect 115 3831 116 3835
rect 794 3835 795 3839
rect 799 3835 800 3839
rect 794 3834 800 3835
rect 922 3839 928 3840
rect 922 3835 923 3839
rect 927 3835 928 3839
rect 922 3834 928 3835
rect 110 3830 116 3831
rect 334 3832 340 3833
rect 112 3799 114 3830
rect 334 3828 335 3832
rect 339 3828 340 3832
rect 334 3827 340 3828
rect 454 3832 460 3833
rect 454 3828 455 3832
rect 459 3828 460 3832
rect 454 3827 460 3828
rect 582 3832 588 3833
rect 582 3828 583 3832
rect 587 3828 588 3832
rect 582 3827 588 3828
rect 718 3832 724 3833
rect 718 3828 719 3832
rect 723 3828 724 3832
rect 718 3827 724 3828
rect 336 3799 338 3827
rect 456 3799 458 3827
rect 574 3803 580 3804
rect 574 3799 575 3803
rect 579 3799 580 3803
rect 584 3799 586 3827
rect 720 3799 722 3827
rect 796 3812 798 3834
rect 846 3832 852 3833
rect 846 3828 847 3832
rect 851 3828 852 3832
rect 846 3827 852 3828
rect 794 3811 800 3812
rect 794 3807 795 3811
rect 799 3807 800 3811
rect 794 3806 800 3807
rect 848 3799 850 3827
rect 924 3812 926 3834
rect 956 3820 958 3910
rect 998 3905 1004 3906
rect 998 3901 999 3905
rect 1003 3901 1004 3905
rect 998 3900 1004 3901
rect 1126 3905 1132 3906
rect 1126 3901 1127 3905
rect 1131 3901 1132 3905
rect 1126 3900 1132 3901
rect 1000 3879 1002 3900
rect 1128 3879 1130 3900
rect 975 3878 979 3879
rect 975 3873 979 3874
rect 999 3878 1003 3879
rect 999 3873 1003 3874
rect 1103 3878 1107 3879
rect 1103 3873 1107 3874
rect 1127 3878 1131 3879
rect 1127 3873 1131 3874
rect 976 3852 978 3873
rect 1104 3852 1106 3873
rect 974 3851 980 3852
rect 974 3847 975 3851
rect 979 3847 980 3851
rect 974 3846 980 3847
rect 1102 3851 1108 3852
rect 1102 3847 1103 3851
rect 1107 3847 1108 3851
rect 1102 3846 1108 3847
rect 1180 3844 1182 3942
rect 1204 3916 1206 3942
rect 1256 3925 1258 3949
rect 1330 3947 1336 3948
rect 1330 3943 1331 3947
rect 1335 3943 1336 3947
rect 1330 3942 1336 3943
rect 1254 3924 1260 3925
rect 1254 3920 1255 3924
rect 1259 3920 1260 3924
rect 1254 3919 1260 3920
rect 1332 3916 1334 3942
rect 1384 3925 1386 3949
rect 1458 3947 1464 3948
rect 1458 3943 1459 3947
rect 1463 3943 1464 3947
rect 1458 3942 1464 3943
rect 1382 3924 1388 3925
rect 1382 3920 1383 3924
rect 1387 3920 1388 3924
rect 1382 3919 1388 3920
rect 1460 3916 1462 3942
rect 1512 3925 1514 3949
rect 1586 3947 1592 3948
rect 1586 3943 1587 3947
rect 1591 3943 1592 3947
rect 1586 3942 1592 3943
rect 1510 3924 1516 3925
rect 1510 3920 1511 3924
rect 1515 3920 1516 3924
rect 1510 3919 1516 3920
rect 1588 3916 1590 3942
rect 1648 3925 1650 3949
rect 1646 3924 1652 3925
rect 1646 3920 1647 3924
rect 1651 3920 1652 3924
rect 2008 3922 2010 3949
rect 2048 3943 2050 3963
rect 2072 3943 2074 3964
rect 2168 3943 2170 3964
rect 2264 3943 2266 3964
rect 3942 3963 3948 3964
rect 3944 3943 3946 3963
rect 2047 3942 2051 3943
rect 2047 3937 2051 3938
rect 2071 3942 2075 3943
rect 2071 3937 2075 3938
rect 2159 3942 2163 3943
rect 2159 3937 2163 3938
rect 2167 3942 2171 3943
rect 2167 3937 2171 3938
rect 2263 3942 2267 3943
rect 2263 3937 2267 3938
rect 2287 3942 2291 3943
rect 2287 3937 2291 3938
rect 2415 3942 2419 3943
rect 2415 3937 2419 3938
rect 2551 3942 2555 3943
rect 2551 3937 2555 3938
rect 2687 3942 2691 3943
rect 2687 3937 2691 3938
rect 2823 3942 2827 3943
rect 2823 3937 2827 3938
rect 2951 3942 2955 3943
rect 2951 3937 2955 3938
rect 3071 3942 3075 3943
rect 3071 3937 3075 3938
rect 3191 3942 3195 3943
rect 3191 3937 3195 3938
rect 3303 3942 3307 3943
rect 3303 3937 3307 3938
rect 3407 3942 3411 3943
rect 3407 3937 3411 3938
rect 3519 3942 3523 3943
rect 3519 3937 3523 3938
rect 3631 3942 3635 3943
rect 3631 3937 3635 3938
rect 3743 3942 3747 3943
rect 3743 3937 3747 3938
rect 3943 3942 3947 3943
rect 3943 3937 3947 3938
rect 1646 3919 1652 3920
rect 2006 3921 2012 3922
rect 2006 3917 2007 3921
rect 2011 3917 2012 3921
rect 2048 3917 2050 3937
rect 2006 3916 2012 3917
rect 2046 3916 2052 3917
rect 2160 3916 2162 3937
rect 2288 3916 2290 3937
rect 2416 3916 2418 3937
rect 2552 3916 2554 3937
rect 2688 3916 2690 3937
rect 2824 3916 2826 3937
rect 2952 3916 2954 3937
rect 3072 3916 3074 3937
rect 3192 3916 3194 3937
rect 3304 3916 3306 3937
rect 3408 3916 3410 3937
rect 3520 3916 3522 3937
rect 3632 3916 3634 3937
rect 3744 3916 3746 3937
rect 3944 3917 3946 3937
rect 3942 3916 3948 3917
rect 1202 3915 1208 3916
rect 1202 3911 1203 3915
rect 1207 3911 1208 3915
rect 1202 3910 1208 3911
rect 1330 3915 1336 3916
rect 1330 3911 1331 3915
rect 1335 3911 1336 3915
rect 1330 3910 1336 3911
rect 1458 3915 1464 3916
rect 1458 3911 1459 3915
rect 1463 3911 1464 3915
rect 1458 3910 1464 3911
rect 1586 3915 1592 3916
rect 1586 3911 1587 3915
rect 1591 3911 1592 3915
rect 2046 3912 2047 3916
rect 2051 3912 2052 3916
rect 2046 3911 2052 3912
rect 2158 3915 2164 3916
rect 2158 3911 2159 3915
rect 2163 3911 2164 3915
rect 1586 3910 1592 3911
rect 2158 3910 2164 3911
rect 2286 3915 2292 3916
rect 2286 3911 2287 3915
rect 2291 3911 2292 3915
rect 2286 3910 2292 3911
rect 2414 3915 2420 3916
rect 2414 3911 2415 3915
rect 2419 3911 2420 3915
rect 2414 3910 2420 3911
rect 2550 3915 2556 3916
rect 2550 3911 2551 3915
rect 2555 3911 2556 3915
rect 2550 3910 2556 3911
rect 2686 3915 2692 3916
rect 2686 3911 2687 3915
rect 2691 3911 2692 3915
rect 2686 3910 2692 3911
rect 2822 3915 2828 3916
rect 2822 3911 2823 3915
rect 2827 3911 2828 3915
rect 2822 3910 2828 3911
rect 2950 3915 2956 3916
rect 2950 3911 2951 3915
rect 2955 3911 2956 3915
rect 2950 3910 2956 3911
rect 3070 3915 3076 3916
rect 3070 3911 3071 3915
rect 3075 3911 3076 3915
rect 3070 3910 3076 3911
rect 3190 3915 3196 3916
rect 3190 3911 3191 3915
rect 3195 3911 3196 3915
rect 3190 3910 3196 3911
rect 3302 3915 3308 3916
rect 3302 3911 3303 3915
rect 3307 3911 3308 3915
rect 3302 3910 3308 3911
rect 3406 3915 3412 3916
rect 3406 3911 3407 3915
rect 3411 3911 3412 3915
rect 3406 3910 3412 3911
rect 3518 3915 3524 3916
rect 3518 3911 3519 3915
rect 3523 3911 3524 3915
rect 3518 3910 3524 3911
rect 3630 3915 3636 3916
rect 3630 3911 3631 3915
rect 3635 3911 3636 3915
rect 3630 3910 3636 3911
rect 3742 3915 3748 3916
rect 3742 3911 3743 3915
rect 3747 3911 3748 3915
rect 3942 3912 3943 3916
rect 3947 3912 3948 3916
rect 3942 3911 3948 3912
rect 3742 3910 3748 3911
rect 3714 3907 3720 3908
rect 1254 3905 1260 3906
rect 1254 3901 1255 3905
rect 1259 3901 1260 3905
rect 1254 3900 1260 3901
rect 1382 3905 1388 3906
rect 1382 3901 1383 3905
rect 1387 3901 1388 3905
rect 1382 3900 1388 3901
rect 1510 3905 1516 3906
rect 1510 3901 1511 3905
rect 1515 3901 1516 3905
rect 1510 3900 1516 3901
rect 1646 3905 1652 3906
rect 1646 3901 1647 3905
rect 1651 3901 1652 3905
rect 1646 3900 1652 3901
rect 2006 3904 2012 3905
rect 2006 3900 2007 3904
rect 2011 3900 2012 3904
rect 2270 3903 2276 3904
rect 1256 3879 1258 3900
rect 1384 3879 1386 3900
rect 1512 3879 1514 3900
rect 1648 3879 1650 3900
rect 2006 3899 2012 3900
rect 2046 3899 2052 3900
rect 2008 3879 2010 3899
rect 2046 3895 2047 3899
rect 2051 3895 2052 3899
rect 2270 3899 2271 3903
rect 2275 3899 2276 3903
rect 2270 3898 2276 3899
rect 2362 3903 2368 3904
rect 2362 3899 2363 3903
rect 2367 3899 2368 3903
rect 2362 3898 2368 3899
rect 2490 3903 2496 3904
rect 2490 3899 2491 3903
rect 2495 3899 2496 3903
rect 2490 3898 2496 3899
rect 2626 3903 2632 3904
rect 2626 3899 2627 3903
rect 2631 3899 2632 3903
rect 2626 3898 2632 3899
rect 2782 3903 2788 3904
rect 2782 3899 2783 3903
rect 2787 3899 2788 3903
rect 2782 3898 2788 3899
rect 2898 3903 2904 3904
rect 2898 3899 2899 3903
rect 2903 3899 2904 3903
rect 2898 3898 2904 3899
rect 3026 3903 3032 3904
rect 3026 3899 3027 3903
rect 3031 3899 3032 3903
rect 3026 3898 3032 3899
rect 3146 3903 3152 3904
rect 3146 3899 3147 3903
rect 3151 3899 3152 3903
rect 3146 3898 3152 3899
rect 3266 3903 3272 3904
rect 3266 3899 3267 3903
rect 3271 3899 3272 3903
rect 3266 3898 3272 3899
rect 3378 3903 3384 3904
rect 3378 3899 3379 3903
rect 3383 3899 3384 3903
rect 3378 3898 3384 3899
rect 3482 3903 3488 3904
rect 3482 3899 3483 3903
rect 3487 3899 3488 3903
rect 3482 3898 3488 3899
rect 3594 3903 3600 3904
rect 3594 3899 3595 3903
rect 3599 3899 3600 3903
rect 3594 3898 3600 3899
rect 3706 3903 3712 3904
rect 3706 3899 3707 3903
rect 3711 3899 3712 3903
rect 3714 3903 3715 3907
rect 3719 3903 3720 3907
rect 3714 3902 3720 3903
rect 3706 3898 3712 3899
rect 2046 3894 2052 3895
rect 2158 3896 2164 3897
rect 1231 3878 1235 3879
rect 1231 3873 1235 3874
rect 1255 3878 1259 3879
rect 1255 3873 1259 3874
rect 1359 3878 1363 3879
rect 1359 3873 1363 3874
rect 1383 3878 1387 3879
rect 1383 3873 1387 3874
rect 1487 3878 1491 3879
rect 1487 3873 1491 3874
rect 1511 3878 1515 3879
rect 1511 3873 1515 3874
rect 1647 3878 1651 3879
rect 1647 3873 1651 3874
rect 2007 3878 2011 3879
rect 2007 3873 2011 3874
rect 1232 3852 1234 3873
rect 1360 3852 1362 3873
rect 1488 3852 1490 3873
rect 2008 3853 2010 3873
rect 2048 3859 2050 3894
rect 2158 3892 2159 3896
rect 2163 3892 2164 3896
rect 2158 3891 2164 3892
rect 2160 3859 2162 3891
rect 2272 3876 2274 3898
rect 2286 3896 2292 3897
rect 2286 3892 2287 3896
rect 2291 3892 2292 3896
rect 2286 3891 2292 3892
rect 2270 3875 2276 3876
rect 2270 3871 2271 3875
rect 2275 3871 2276 3875
rect 2270 3870 2276 3871
rect 2288 3859 2290 3891
rect 2364 3876 2366 3898
rect 2414 3896 2420 3897
rect 2414 3892 2415 3896
rect 2419 3892 2420 3896
rect 2414 3891 2420 3892
rect 2362 3875 2368 3876
rect 2362 3871 2363 3875
rect 2367 3871 2368 3875
rect 2362 3870 2368 3871
rect 2416 3859 2418 3891
rect 2492 3876 2494 3898
rect 2550 3896 2556 3897
rect 2550 3892 2551 3896
rect 2555 3892 2556 3896
rect 2550 3891 2556 3892
rect 2490 3875 2496 3876
rect 2490 3871 2491 3875
rect 2495 3871 2496 3875
rect 2490 3870 2496 3871
rect 2552 3859 2554 3891
rect 2628 3876 2630 3898
rect 2686 3896 2692 3897
rect 2686 3892 2687 3896
rect 2691 3892 2692 3896
rect 2686 3891 2692 3892
rect 2626 3875 2632 3876
rect 2626 3871 2627 3875
rect 2631 3871 2632 3875
rect 2626 3870 2632 3871
rect 2688 3859 2690 3891
rect 2047 3858 2051 3859
rect 2047 3853 2051 3854
rect 2159 3858 2163 3859
rect 2159 3853 2163 3854
rect 2207 3858 2211 3859
rect 2207 3853 2211 3854
rect 2287 3858 2291 3859
rect 2287 3853 2291 3854
rect 2343 3858 2347 3859
rect 2343 3853 2347 3854
rect 2415 3858 2419 3859
rect 2415 3853 2419 3854
rect 2487 3858 2491 3859
rect 2487 3853 2491 3854
rect 2551 3858 2555 3859
rect 2551 3853 2555 3854
rect 2647 3858 2651 3859
rect 2647 3853 2651 3854
rect 2687 3858 2691 3859
rect 2687 3853 2691 3854
rect 2006 3852 2012 3853
rect 1230 3851 1236 3852
rect 1230 3847 1231 3851
rect 1235 3847 1236 3851
rect 1230 3846 1236 3847
rect 1358 3851 1364 3852
rect 1358 3847 1359 3851
rect 1363 3847 1364 3851
rect 1358 3846 1364 3847
rect 1486 3851 1492 3852
rect 1486 3847 1487 3851
rect 1491 3847 1492 3851
rect 2006 3848 2007 3852
rect 2011 3848 2012 3852
rect 2006 3847 2012 3848
rect 1486 3846 1492 3847
rect 1178 3843 1184 3844
rect 1050 3839 1056 3840
rect 1050 3835 1051 3839
rect 1055 3835 1056 3839
rect 1178 3839 1179 3843
rect 1183 3839 1184 3843
rect 1178 3838 1184 3839
rect 1214 3843 1220 3844
rect 1214 3839 1215 3843
rect 1219 3839 1220 3843
rect 1214 3838 1220 3839
rect 1342 3843 1348 3844
rect 1342 3839 1343 3843
rect 1347 3839 1348 3843
rect 1342 3838 1348 3839
rect 1050 3834 1056 3835
rect 974 3832 980 3833
rect 974 3828 975 3832
rect 979 3828 980 3832
rect 974 3827 980 3828
rect 954 3819 960 3820
rect 954 3815 955 3819
rect 959 3815 960 3819
rect 954 3814 960 3815
rect 922 3811 928 3812
rect 922 3807 923 3811
rect 927 3807 928 3811
rect 922 3806 928 3807
rect 976 3799 978 3827
rect 111 3798 115 3799
rect 111 3793 115 3794
rect 335 3798 339 3799
rect 335 3793 339 3794
rect 455 3798 459 3799
rect 455 3793 459 3794
rect 503 3798 507 3799
rect 574 3798 580 3799
rect 583 3798 587 3799
rect 503 3793 507 3794
rect 112 3766 114 3793
rect 504 3769 506 3793
rect 502 3768 508 3769
rect 110 3765 116 3766
rect 110 3761 111 3765
rect 115 3761 116 3765
rect 502 3764 503 3768
rect 507 3764 508 3768
rect 502 3763 508 3764
rect 110 3760 116 3761
rect 576 3760 578 3798
rect 583 3793 587 3794
rect 615 3798 619 3799
rect 615 3793 619 3794
rect 719 3798 723 3799
rect 719 3793 723 3794
rect 735 3798 739 3799
rect 735 3793 739 3794
rect 847 3798 851 3799
rect 847 3793 851 3794
rect 863 3798 867 3799
rect 863 3793 867 3794
rect 975 3798 979 3799
rect 975 3793 979 3794
rect 999 3798 1003 3799
rect 999 3793 1003 3794
rect 590 3791 596 3792
rect 590 3787 591 3791
rect 595 3787 596 3791
rect 590 3786 596 3787
rect 592 3760 594 3786
rect 616 3769 618 3793
rect 698 3791 704 3792
rect 698 3787 699 3791
rect 703 3787 704 3791
rect 698 3786 704 3787
rect 614 3768 620 3769
rect 614 3764 615 3768
rect 619 3764 620 3768
rect 614 3763 620 3764
rect 700 3760 702 3786
rect 736 3769 738 3793
rect 818 3791 824 3792
rect 818 3787 819 3791
rect 823 3787 824 3791
rect 818 3786 824 3787
rect 734 3768 740 3769
rect 734 3764 735 3768
rect 739 3764 740 3768
rect 734 3763 740 3764
rect 820 3760 822 3786
rect 864 3769 866 3793
rect 902 3791 908 3792
rect 902 3787 903 3791
rect 907 3787 908 3791
rect 902 3786 908 3787
rect 862 3768 868 3769
rect 862 3764 863 3768
rect 867 3764 868 3768
rect 862 3763 868 3764
rect 574 3759 580 3760
rect 574 3755 575 3759
rect 579 3755 580 3759
rect 574 3754 580 3755
rect 590 3759 596 3760
rect 590 3755 591 3759
rect 595 3755 596 3759
rect 590 3754 596 3755
rect 698 3759 704 3760
rect 698 3755 699 3759
rect 703 3755 704 3759
rect 698 3754 704 3755
rect 818 3759 824 3760
rect 818 3755 819 3759
rect 823 3755 824 3759
rect 818 3754 824 3755
rect 502 3749 508 3750
rect 110 3748 116 3749
rect 110 3744 111 3748
rect 115 3744 116 3748
rect 502 3745 503 3749
rect 507 3745 508 3749
rect 502 3744 508 3745
rect 614 3749 620 3750
rect 614 3745 615 3749
rect 619 3745 620 3749
rect 614 3744 620 3745
rect 734 3749 740 3750
rect 734 3745 735 3749
rect 739 3745 740 3749
rect 734 3744 740 3745
rect 862 3749 868 3750
rect 862 3745 863 3749
rect 867 3745 868 3749
rect 862 3744 868 3745
rect 110 3743 116 3744
rect 112 3715 114 3743
rect 504 3715 506 3744
rect 616 3715 618 3744
rect 736 3715 738 3744
rect 864 3715 866 3744
rect 111 3714 115 3715
rect 111 3709 115 3710
rect 495 3714 499 3715
rect 495 3709 499 3710
rect 503 3714 507 3715
rect 503 3709 507 3710
rect 591 3714 595 3715
rect 591 3709 595 3710
rect 615 3714 619 3715
rect 615 3709 619 3710
rect 687 3714 691 3715
rect 687 3709 691 3710
rect 735 3714 739 3715
rect 735 3709 739 3710
rect 791 3714 795 3715
rect 791 3709 795 3710
rect 863 3714 867 3715
rect 863 3709 867 3710
rect 112 3689 114 3709
rect 110 3688 116 3689
rect 496 3688 498 3709
rect 592 3688 594 3709
rect 688 3688 690 3709
rect 792 3688 794 3709
rect 110 3684 111 3688
rect 115 3684 116 3688
rect 110 3683 116 3684
rect 494 3687 500 3688
rect 494 3683 495 3687
rect 499 3683 500 3687
rect 494 3682 500 3683
rect 590 3687 596 3688
rect 590 3683 591 3687
rect 595 3683 596 3687
rect 590 3682 596 3683
rect 686 3687 692 3688
rect 686 3683 687 3687
rect 691 3683 692 3687
rect 686 3682 692 3683
rect 790 3687 796 3688
rect 790 3683 791 3687
rect 795 3683 796 3687
rect 790 3682 796 3683
rect 904 3680 906 3786
rect 1000 3769 1002 3793
rect 1052 3792 1054 3834
rect 1102 3832 1108 3833
rect 1102 3828 1103 3832
rect 1107 3828 1108 3832
rect 1102 3827 1108 3828
rect 1104 3799 1106 3827
rect 1216 3812 1218 3838
rect 1230 3832 1236 3833
rect 1230 3828 1231 3832
rect 1235 3828 1236 3832
rect 1230 3827 1236 3828
rect 1214 3811 1220 3812
rect 1214 3807 1215 3811
rect 1219 3807 1220 3811
rect 1214 3806 1220 3807
rect 1232 3799 1234 3827
rect 1344 3812 1346 3838
rect 2006 3835 2012 3836
rect 1358 3832 1364 3833
rect 1358 3828 1359 3832
rect 1363 3828 1364 3832
rect 1358 3827 1364 3828
rect 1486 3832 1492 3833
rect 1486 3828 1487 3832
rect 1491 3828 1492 3832
rect 2006 3831 2007 3835
rect 2011 3831 2012 3835
rect 2006 3830 2012 3831
rect 1486 3827 1492 3828
rect 1342 3811 1348 3812
rect 1342 3807 1343 3811
rect 1347 3807 1348 3811
rect 1342 3806 1348 3807
rect 1360 3799 1362 3827
rect 1488 3799 1490 3827
rect 1506 3807 1512 3808
rect 1506 3803 1507 3807
rect 1511 3803 1512 3807
rect 1506 3802 1512 3803
rect 1103 3798 1107 3799
rect 1103 3793 1107 3794
rect 1143 3798 1147 3799
rect 1143 3793 1147 3794
rect 1231 3798 1235 3799
rect 1231 3793 1235 3794
rect 1287 3798 1291 3799
rect 1287 3793 1291 3794
rect 1359 3798 1363 3799
rect 1359 3793 1363 3794
rect 1431 3798 1435 3799
rect 1431 3793 1435 3794
rect 1487 3798 1491 3799
rect 1487 3793 1491 3794
rect 1050 3791 1056 3792
rect 1050 3787 1051 3791
rect 1055 3787 1056 3791
rect 1050 3786 1056 3787
rect 1074 3791 1080 3792
rect 1074 3787 1075 3791
rect 1079 3787 1080 3791
rect 1074 3786 1080 3787
rect 998 3768 1004 3769
rect 998 3764 999 3768
rect 1003 3764 1004 3768
rect 998 3763 1004 3764
rect 1076 3760 1078 3786
rect 1144 3769 1146 3793
rect 1288 3769 1290 3793
rect 1406 3791 1412 3792
rect 1406 3787 1407 3791
rect 1411 3787 1412 3791
rect 1406 3786 1412 3787
rect 1142 3768 1148 3769
rect 1142 3764 1143 3768
rect 1147 3764 1148 3768
rect 1142 3763 1148 3764
rect 1286 3768 1292 3769
rect 1286 3764 1287 3768
rect 1291 3764 1292 3768
rect 1286 3763 1292 3764
rect 1408 3760 1410 3786
rect 1432 3769 1434 3793
rect 1430 3768 1436 3769
rect 1430 3764 1431 3768
rect 1435 3764 1436 3768
rect 1430 3763 1436 3764
rect 1508 3760 1510 3802
rect 2008 3799 2010 3830
rect 2048 3826 2050 3853
rect 2208 3829 2210 3853
rect 2294 3851 2300 3852
rect 2294 3847 2295 3851
rect 2299 3847 2300 3851
rect 2294 3846 2300 3847
rect 2206 3828 2212 3829
rect 2046 3825 2052 3826
rect 2046 3821 2047 3825
rect 2051 3821 2052 3825
rect 2206 3824 2207 3828
rect 2211 3824 2212 3828
rect 2206 3823 2212 3824
rect 2046 3820 2052 3821
rect 2296 3820 2298 3846
rect 2344 3829 2346 3853
rect 2426 3851 2432 3852
rect 2426 3847 2427 3851
rect 2431 3847 2432 3851
rect 2426 3846 2432 3847
rect 2342 3828 2348 3829
rect 2342 3824 2343 3828
rect 2347 3824 2348 3828
rect 2342 3823 2348 3824
rect 2428 3820 2430 3846
rect 2488 3829 2490 3853
rect 2570 3851 2576 3852
rect 2570 3847 2571 3851
rect 2575 3847 2576 3851
rect 2570 3846 2576 3847
rect 2486 3828 2492 3829
rect 2486 3824 2487 3828
rect 2491 3824 2492 3828
rect 2486 3823 2492 3824
rect 2572 3820 2574 3846
rect 2648 3829 2650 3853
rect 2784 3852 2786 3898
rect 2822 3896 2828 3897
rect 2822 3892 2823 3896
rect 2827 3892 2828 3896
rect 2822 3891 2828 3892
rect 2824 3859 2826 3891
rect 2900 3876 2902 3898
rect 2950 3896 2956 3897
rect 2950 3892 2951 3896
rect 2955 3892 2956 3896
rect 2950 3891 2956 3892
rect 2898 3875 2904 3876
rect 2898 3871 2899 3875
rect 2903 3871 2904 3875
rect 2898 3870 2904 3871
rect 2952 3859 2954 3891
rect 3028 3876 3030 3898
rect 3070 3896 3076 3897
rect 3070 3892 3071 3896
rect 3075 3892 3076 3896
rect 3070 3891 3076 3892
rect 3026 3875 3032 3876
rect 3026 3871 3027 3875
rect 3031 3871 3032 3875
rect 3026 3870 3032 3871
rect 3072 3859 3074 3891
rect 3148 3876 3150 3898
rect 3190 3896 3196 3897
rect 3190 3892 3191 3896
rect 3195 3892 3196 3896
rect 3190 3891 3196 3892
rect 3146 3875 3152 3876
rect 3146 3871 3147 3875
rect 3151 3871 3152 3875
rect 3146 3870 3152 3871
rect 3192 3859 3194 3891
rect 3268 3876 3270 3898
rect 3302 3896 3308 3897
rect 3302 3892 3303 3896
rect 3307 3892 3308 3896
rect 3302 3891 3308 3892
rect 3266 3875 3272 3876
rect 3266 3871 3267 3875
rect 3271 3871 3272 3875
rect 3266 3870 3272 3871
rect 3304 3859 3306 3891
rect 3380 3876 3382 3898
rect 3406 3896 3412 3897
rect 3406 3892 3407 3896
rect 3411 3892 3412 3896
rect 3406 3891 3412 3892
rect 3378 3875 3384 3876
rect 3378 3871 3379 3875
rect 3383 3871 3384 3875
rect 3378 3870 3384 3871
rect 3408 3859 3410 3891
rect 3484 3876 3486 3898
rect 3518 3896 3524 3897
rect 3518 3892 3519 3896
rect 3523 3892 3524 3896
rect 3518 3891 3524 3892
rect 3482 3875 3488 3876
rect 3482 3871 3483 3875
rect 3487 3871 3488 3875
rect 3482 3870 3488 3871
rect 3520 3859 3522 3891
rect 3596 3876 3598 3898
rect 3630 3896 3636 3897
rect 3630 3892 3631 3896
rect 3635 3892 3636 3896
rect 3630 3891 3636 3892
rect 3594 3875 3600 3876
rect 3594 3871 3595 3875
rect 3599 3871 3600 3875
rect 3594 3870 3600 3871
rect 3632 3859 3634 3891
rect 3708 3876 3710 3898
rect 3706 3875 3712 3876
rect 3706 3871 3707 3875
rect 3711 3871 3712 3875
rect 3706 3870 3712 3871
rect 3716 3859 3718 3902
rect 3942 3899 3948 3900
rect 3742 3896 3748 3897
rect 3742 3892 3743 3896
rect 3747 3892 3748 3896
rect 3942 3895 3943 3899
rect 3947 3895 3948 3899
rect 3942 3894 3948 3895
rect 3742 3891 3748 3892
rect 3744 3859 3746 3891
rect 3944 3859 3946 3894
rect 2823 3858 2827 3859
rect 2823 3853 2827 3854
rect 2951 3858 2955 3859
rect 2951 3853 2955 3854
rect 3015 3858 3019 3859
rect 3015 3853 3019 3854
rect 3071 3858 3075 3859
rect 3071 3853 3075 3854
rect 3191 3858 3195 3859
rect 3191 3853 3195 3854
rect 3223 3858 3227 3859
rect 3223 3853 3227 3854
rect 3303 3858 3307 3859
rect 3303 3853 3307 3854
rect 3407 3858 3411 3859
rect 3407 3853 3411 3854
rect 3439 3858 3443 3859
rect 3439 3853 3443 3854
rect 3519 3858 3523 3859
rect 3519 3853 3523 3854
rect 3631 3858 3635 3859
rect 3631 3853 3635 3854
rect 3655 3858 3659 3859
rect 3655 3853 3659 3854
rect 3712 3857 3718 3859
rect 3743 3858 3747 3859
rect 2782 3851 2788 3852
rect 2782 3847 2783 3851
rect 2787 3847 2788 3851
rect 2782 3846 2788 3847
rect 2824 3829 2826 3853
rect 3016 3829 3018 3853
rect 3098 3851 3104 3852
rect 3098 3847 3099 3851
rect 3103 3847 3104 3851
rect 3098 3846 3104 3847
rect 2646 3828 2652 3829
rect 2646 3824 2647 3828
rect 2651 3824 2652 3828
rect 2646 3823 2652 3824
rect 2822 3828 2828 3829
rect 2822 3824 2823 3828
rect 2827 3824 2828 3828
rect 2822 3823 2828 3824
rect 3014 3828 3020 3829
rect 3014 3824 3015 3828
rect 3019 3824 3020 3828
rect 3014 3823 3020 3824
rect 3100 3820 3102 3846
rect 3224 3829 3226 3853
rect 3310 3851 3316 3852
rect 3310 3847 3311 3851
rect 3315 3847 3316 3851
rect 3310 3846 3316 3847
rect 3394 3851 3400 3852
rect 3394 3847 3395 3851
rect 3399 3847 3400 3851
rect 3394 3846 3400 3847
rect 3222 3828 3228 3829
rect 3222 3824 3223 3828
rect 3227 3824 3228 3828
rect 3222 3823 3228 3824
rect 3312 3820 3314 3846
rect 2274 3819 2280 3820
rect 2274 3815 2275 3819
rect 2279 3815 2280 3819
rect 2274 3814 2280 3815
rect 2294 3819 2300 3820
rect 2294 3815 2295 3819
rect 2299 3815 2300 3819
rect 2294 3814 2300 3815
rect 2426 3819 2432 3820
rect 2426 3815 2427 3819
rect 2431 3815 2432 3819
rect 2426 3814 2432 3815
rect 2570 3819 2576 3820
rect 2570 3815 2571 3819
rect 2575 3815 2576 3819
rect 2570 3814 2576 3815
rect 3098 3819 3104 3820
rect 3098 3815 3099 3819
rect 3103 3815 3104 3819
rect 3098 3814 3104 3815
rect 3310 3819 3316 3820
rect 3310 3815 3311 3819
rect 3315 3815 3316 3819
rect 3310 3814 3316 3815
rect 2206 3809 2212 3810
rect 2046 3808 2052 3809
rect 2046 3804 2047 3808
rect 2051 3804 2052 3808
rect 2206 3805 2207 3809
rect 2211 3805 2212 3809
rect 2206 3804 2212 3805
rect 2046 3803 2052 3804
rect 1583 3798 1587 3799
rect 1583 3793 1587 3794
rect 2007 3798 2011 3799
rect 2007 3793 2011 3794
rect 1570 3791 1576 3792
rect 1570 3787 1571 3791
rect 1575 3787 1576 3791
rect 1570 3786 1576 3787
rect 1514 3783 1520 3784
rect 1514 3779 1515 3783
rect 1519 3779 1520 3783
rect 1514 3778 1520 3779
rect 1516 3760 1518 3778
rect 1074 3759 1080 3760
rect 1074 3755 1075 3759
rect 1079 3755 1080 3759
rect 1074 3754 1080 3755
rect 1218 3759 1224 3760
rect 1218 3755 1219 3759
rect 1223 3755 1224 3759
rect 1218 3754 1224 3755
rect 1406 3759 1412 3760
rect 1406 3755 1407 3759
rect 1411 3755 1412 3759
rect 1406 3754 1412 3755
rect 1506 3759 1512 3760
rect 1506 3755 1507 3759
rect 1511 3755 1512 3759
rect 1506 3754 1512 3755
rect 1514 3759 1520 3760
rect 1514 3755 1515 3759
rect 1519 3755 1520 3759
rect 1514 3754 1520 3755
rect 998 3749 1004 3750
rect 998 3745 999 3749
rect 1003 3745 1004 3749
rect 998 3744 1004 3745
rect 1142 3749 1148 3750
rect 1142 3745 1143 3749
rect 1147 3745 1148 3749
rect 1142 3744 1148 3745
rect 1000 3715 1002 3744
rect 1144 3715 1146 3744
rect 911 3714 915 3715
rect 911 3709 915 3710
rect 999 3714 1003 3715
rect 999 3709 1003 3710
rect 1039 3714 1043 3715
rect 1039 3709 1043 3710
rect 1143 3714 1147 3715
rect 1143 3709 1147 3710
rect 1183 3714 1187 3715
rect 1183 3709 1187 3710
rect 912 3688 914 3709
rect 1040 3688 1042 3709
rect 1184 3688 1186 3709
rect 910 3687 916 3688
rect 910 3683 911 3687
rect 915 3683 916 3687
rect 910 3682 916 3683
rect 1038 3687 1044 3688
rect 1038 3683 1039 3687
rect 1043 3683 1044 3687
rect 1038 3682 1044 3683
rect 1182 3687 1188 3688
rect 1182 3683 1183 3687
rect 1187 3683 1188 3687
rect 1182 3682 1188 3683
rect 902 3679 908 3680
rect 570 3675 576 3676
rect 110 3671 116 3672
rect 110 3667 111 3671
rect 115 3667 116 3671
rect 570 3671 571 3675
rect 575 3671 576 3675
rect 570 3670 576 3671
rect 666 3675 672 3676
rect 666 3671 667 3675
rect 671 3671 672 3675
rect 666 3670 672 3671
rect 762 3675 768 3676
rect 762 3671 763 3675
rect 767 3671 768 3675
rect 762 3670 768 3671
rect 866 3675 872 3676
rect 866 3671 867 3675
rect 871 3671 872 3675
rect 902 3675 903 3679
rect 907 3675 908 3679
rect 902 3674 908 3675
rect 1114 3675 1120 3676
rect 866 3670 872 3671
rect 1114 3671 1115 3675
rect 1119 3671 1120 3675
rect 1114 3670 1120 3671
rect 110 3666 116 3667
rect 494 3668 500 3669
rect 112 3631 114 3666
rect 494 3664 495 3668
rect 499 3664 500 3668
rect 494 3663 500 3664
rect 496 3631 498 3663
rect 572 3648 574 3670
rect 590 3668 596 3669
rect 590 3664 591 3668
rect 595 3664 596 3668
rect 590 3663 596 3664
rect 570 3647 576 3648
rect 570 3643 571 3647
rect 575 3643 576 3647
rect 570 3642 576 3643
rect 592 3631 594 3663
rect 668 3648 670 3670
rect 686 3668 692 3669
rect 686 3664 687 3668
rect 691 3664 692 3668
rect 686 3663 692 3664
rect 666 3647 672 3648
rect 666 3643 667 3647
rect 671 3643 672 3647
rect 666 3642 672 3643
rect 688 3631 690 3663
rect 764 3648 766 3670
rect 790 3668 796 3669
rect 790 3664 791 3668
rect 795 3664 796 3668
rect 790 3663 796 3664
rect 762 3647 768 3648
rect 762 3643 763 3647
rect 767 3643 768 3647
rect 762 3642 768 3643
rect 792 3631 794 3663
rect 868 3648 870 3670
rect 910 3668 916 3669
rect 910 3664 911 3668
rect 915 3664 916 3668
rect 910 3663 916 3664
rect 1038 3668 1044 3669
rect 1038 3664 1039 3668
rect 1043 3664 1044 3668
rect 1038 3663 1044 3664
rect 866 3647 872 3648
rect 866 3643 867 3647
rect 871 3643 872 3647
rect 866 3642 872 3643
rect 858 3639 864 3640
rect 858 3635 859 3639
rect 863 3635 864 3639
rect 858 3634 864 3635
rect 111 3630 115 3631
rect 111 3625 115 3626
rect 335 3630 339 3631
rect 335 3625 339 3626
rect 463 3630 467 3631
rect 463 3625 467 3626
rect 495 3630 499 3631
rect 495 3625 499 3626
rect 591 3630 595 3631
rect 591 3625 595 3626
rect 607 3630 611 3631
rect 607 3625 611 3626
rect 687 3630 691 3631
rect 687 3625 691 3626
rect 759 3630 763 3631
rect 759 3625 763 3626
rect 791 3630 795 3631
rect 791 3625 795 3626
rect 112 3598 114 3625
rect 336 3601 338 3625
rect 410 3623 416 3624
rect 410 3619 411 3623
rect 415 3619 416 3623
rect 410 3618 416 3619
rect 334 3600 340 3601
rect 110 3597 116 3598
rect 110 3593 111 3597
rect 115 3593 116 3597
rect 334 3596 335 3600
rect 339 3596 340 3600
rect 334 3595 340 3596
rect 110 3592 116 3593
rect 412 3592 414 3618
rect 464 3601 466 3625
rect 538 3623 544 3624
rect 538 3619 539 3623
rect 543 3619 544 3623
rect 538 3618 544 3619
rect 462 3600 468 3601
rect 462 3596 463 3600
rect 467 3596 468 3600
rect 462 3595 468 3596
rect 540 3592 542 3618
rect 608 3601 610 3625
rect 738 3615 744 3616
rect 738 3611 739 3615
rect 743 3611 744 3615
rect 738 3610 744 3611
rect 606 3600 612 3601
rect 606 3596 607 3600
rect 611 3596 612 3600
rect 606 3595 612 3596
rect 410 3591 416 3592
rect 410 3587 411 3591
rect 415 3587 416 3591
rect 410 3586 416 3587
rect 538 3591 544 3592
rect 538 3587 539 3591
rect 543 3587 544 3591
rect 538 3586 544 3587
rect 334 3581 340 3582
rect 110 3580 116 3581
rect 110 3576 111 3580
rect 115 3576 116 3580
rect 334 3577 335 3581
rect 339 3577 340 3581
rect 334 3576 340 3577
rect 462 3581 468 3582
rect 462 3577 463 3581
rect 467 3577 468 3581
rect 462 3576 468 3577
rect 606 3581 612 3582
rect 606 3577 607 3581
rect 611 3577 612 3581
rect 606 3576 612 3577
rect 110 3575 116 3576
rect 112 3543 114 3575
rect 336 3543 338 3576
rect 464 3543 466 3576
rect 608 3543 610 3576
rect 111 3542 115 3543
rect 111 3537 115 3538
rect 159 3542 163 3543
rect 159 3537 163 3538
rect 303 3542 307 3543
rect 303 3537 307 3538
rect 335 3542 339 3543
rect 335 3537 339 3538
rect 463 3542 467 3543
rect 463 3537 467 3538
rect 607 3542 611 3543
rect 607 3537 611 3538
rect 639 3542 643 3543
rect 639 3537 643 3538
rect 112 3517 114 3537
rect 110 3516 116 3517
rect 160 3516 162 3537
rect 304 3516 306 3537
rect 464 3516 466 3537
rect 640 3516 642 3537
rect 110 3512 111 3516
rect 115 3512 116 3516
rect 110 3511 116 3512
rect 158 3515 164 3516
rect 158 3511 159 3515
rect 163 3511 164 3515
rect 158 3510 164 3511
rect 302 3515 308 3516
rect 302 3511 303 3515
rect 307 3511 308 3515
rect 302 3510 308 3511
rect 462 3515 468 3516
rect 462 3511 463 3515
rect 467 3511 468 3515
rect 462 3510 468 3511
rect 638 3515 644 3516
rect 638 3511 639 3515
rect 643 3511 644 3515
rect 638 3510 644 3511
rect 740 3508 742 3610
rect 760 3601 762 3625
rect 834 3623 840 3624
rect 834 3619 835 3623
rect 839 3619 840 3623
rect 834 3618 840 3619
rect 758 3600 764 3601
rect 758 3596 759 3600
rect 763 3596 764 3600
rect 758 3595 764 3596
rect 836 3592 838 3618
rect 860 3592 862 3634
rect 912 3631 914 3663
rect 1040 3631 1042 3663
rect 911 3630 915 3631
rect 911 3625 915 3626
rect 927 3630 931 3631
rect 927 3625 931 3626
rect 1039 3630 1043 3631
rect 1039 3625 1043 3626
rect 1095 3630 1099 3631
rect 1095 3625 1099 3626
rect 928 3601 930 3625
rect 1096 3601 1098 3625
rect 1116 3624 1118 3670
rect 1182 3668 1188 3669
rect 1182 3664 1183 3668
rect 1187 3664 1188 3668
rect 1182 3663 1188 3664
rect 1184 3631 1186 3663
rect 1220 3648 1222 3754
rect 1286 3749 1292 3750
rect 1286 3745 1287 3749
rect 1291 3745 1292 3749
rect 1286 3744 1292 3745
rect 1430 3749 1436 3750
rect 1430 3745 1431 3749
rect 1435 3745 1436 3749
rect 1430 3744 1436 3745
rect 1288 3715 1290 3744
rect 1432 3715 1434 3744
rect 1287 3714 1291 3715
rect 1287 3709 1291 3710
rect 1335 3714 1339 3715
rect 1335 3709 1339 3710
rect 1431 3714 1435 3715
rect 1431 3709 1435 3710
rect 1495 3714 1499 3715
rect 1495 3709 1499 3710
rect 1336 3688 1338 3709
rect 1496 3688 1498 3709
rect 1334 3687 1340 3688
rect 1334 3683 1335 3687
rect 1339 3683 1340 3687
rect 1334 3682 1340 3683
rect 1494 3687 1500 3688
rect 1494 3683 1495 3687
rect 1499 3683 1500 3687
rect 1494 3682 1500 3683
rect 1572 3680 1574 3786
rect 1584 3769 1586 3793
rect 1582 3768 1588 3769
rect 1582 3764 1583 3768
rect 1587 3764 1588 3768
rect 2008 3766 2010 3793
rect 2048 3783 2050 3803
rect 2208 3783 2210 3804
rect 2047 3782 2051 3783
rect 2047 3777 2051 3778
rect 2191 3782 2195 3783
rect 2191 3777 2195 3778
rect 2207 3782 2211 3783
rect 2207 3777 2211 3778
rect 1582 3763 1588 3764
rect 2006 3765 2012 3766
rect 2006 3761 2007 3765
rect 2011 3761 2012 3765
rect 2006 3760 2012 3761
rect 2048 3757 2050 3777
rect 2046 3756 2052 3757
rect 2192 3756 2194 3777
rect 2046 3752 2047 3756
rect 2051 3752 2052 3756
rect 2046 3751 2052 3752
rect 2190 3755 2196 3756
rect 2190 3751 2191 3755
rect 2195 3751 2196 3755
rect 2190 3750 2196 3751
rect 1582 3749 1588 3750
rect 1582 3745 1583 3749
rect 1587 3745 1588 3749
rect 1582 3744 1588 3745
rect 2006 3748 2012 3749
rect 2006 3744 2007 3748
rect 2011 3744 2012 3748
rect 1584 3715 1586 3744
rect 2006 3743 2012 3744
rect 2008 3715 2010 3743
rect 2046 3739 2052 3740
rect 2046 3735 2047 3739
rect 2051 3735 2052 3739
rect 2046 3734 2052 3735
rect 2190 3736 2196 3737
rect 1583 3714 1587 3715
rect 1583 3709 1587 3710
rect 1655 3714 1659 3715
rect 1655 3709 1659 3710
rect 2007 3714 2011 3715
rect 2007 3709 2011 3710
rect 1656 3688 1658 3709
rect 2008 3689 2010 3709
rect 2048 3703 2050 3734
rect 2190 3732 2191 3736
rect 2195 3732 2196 3736
rect 2190 3731 2196 3732
rect 2192 3703 2194 3731
rect 2276 3716 2278 3814
rect 2342 3809 2348 3810
rect 2342 3805 2343 3809
rect 2347 3805 2348 3809
rect 2342 3804 2348 3805
rect 2486 3809 2492 3810
rect 2486 3805 2487 3809
rect 2491 3805 2492 3809
rect 2486 3804 2492 3805
rect 2646 3809 2652 3810
rect 2646 3805 2647 3809
rect 2651 3805 2652 3809
rect 2646 3804 2652 3805
rect 2822 3809 2828 3810
rect 2822 3805 2823 3809
rect 2827 3805 2828 3809
rect 2822 3804 2828 3805
rect 3014 3809 3020 3810
rect 3014 3805 3015 3809
rect 3019 3805 3020 3809
rect 3014 3804 3020 3805
rect 3222 3809 3228 3810
rect 3222 3805 3223 3809
rect 3227 3805 3228 3809
rect 3222 3804 3228 3805
rect 2344 3783 2346 3804
rect 2488 3783 2490 3804
rect 2648 3783 2650 3804
rect 2824 3783 2826 3804
rect 3016 3783 3018 3804
rect 3224 3783 3226 3804
rect 2343 3782 2347 3783
rect 2343 3777 2347 3778
rect 2375 3782 2379 3783
rect 2375 3777 2379 3778
rect 2487 3782 2491 3783
rect 2487 3777 2491 3778
rect 2559 3782 2563 3783
rect 2559 3777 2563 3778
rect 2647 3782 2651 3783
rect 2647 3777 2651 3778
rect 2743 3782 2747 3783
rect 2743 3777 2747 3778
rect 2823 3782 2827 3783
rect 2823 3777 2827 3778
rect 2935 3782 2939 3783
rect 2935 3777 2939 3778
rect 3015 3782 3019 3783
rect 3015 3777 3019 3778
rect 3127 3782 3131 3783
rect 3127 3777 3131 3778
rect 3223 3782 3227 3783
rect 3223 3777 3227 3778
rect 3319 3782 3323 3783
rect 3319 3777 3323 3778
rect 2376 3756 2378 3777
rect 2560 3756 2562 3777
rect 2744 3756 2746 3777
rect 2936 3756 2938 3777
rect 3128 3756 3130 3777
rect 3320 3756 3322 3777
rect 2374 3755 2380 3756
rect 2374 3751 2375 3755
rect 2379 3751 2380 3755
rect 2374 3750 2380 3751
rect 2558 3755 2564 3756
rect 2558 3751 2559 3755
rect 2563 3751 2564 3755
rect 2558 3750 2564 3751
rect 2742 3755 2748 3756
rect 2742 3751 2743 3755
rect 2747 3751 2748 3755
rect 2742 3750 2748 3751
rect 2934 3755 2940 3756
rect 2934 3751 2935 3755
rect 2939 3751 2940 3755
rect 2934 3750 2940 3751
rect 3126 3755 3132 3756
rect 3126 3751 3127 3755
rect 3131 3751 3132 3755
rect 3126 3750 3132 3751
rect 3318 3755 3324 3756
rect 3318 3751 3319 3755
rect 3323 3751 3324 3755
rect 3318 3750 3324 3751
rect 3396 3748 3398 3846
rect 3440 3829 3442 3853
rect 3656 3829 3658 3853
rect 3712 3852 3714 3857
rect 3743 3853 3747 3854
rect 3943 3858 3947 3859
rect 3943 3853 3947 3854
rect 3710 3851 3716 3852
rect 3710 3847 3711 3851
rect 3715 3847 3716 3851
rect 3710 3846 3716 3847
rect 3438 3828 3444 3829
rect 3438 3824 3439 3828
rect 3443 3824 3444 3828
rect 3438 3823 3444 3824
rect 3654 3828 3660 3829
rect 3654 3824 3655 3828
rect 3659 3824 3660 3828
rect 3944 3826 3946 3853
rect 3654 3823 3660 3824
rect 3942 3825 3948 3826
rect 3942 3821 3943 3825
rect 3947 3821 3948 3825
rect 3942 3820 3948 3821
rect 3730 3819 3736 3820
rect 3730 3815 3731 3819
rect 3735 3815 3736 3819
rect 3730 3814 3736 3815
rect 3438 3809 3444 3810
rect 3438 3805 3439 3809
rect 3443 3805 3444 3809
rect 3438 3804 3444 3805
rect 3654 3809 3660 3810
rect 3654 3805 3655 3809
rect 3659 3805 3660 3809
rect 3654 3804 3660 3805
rect 3440 3783 3442 3804
rect 3656 3783 3658 3804
rect 3439 3782 3443 3783
rect 3439 3777 3443 3778
rect 3511 3782 3515 3783
rect 3511 3777 3515 3778
rect 3655 3782 3659 3783
rect 3655 3777 3659 3778
rect 3711 3782 3715 3783
rect 3711 3777 3715 3778
rect 3512 3756 3514 3777
rect 3712 3756 3714 3777
rect 3510 3755 3516 3756
rect 3510 3751 3511 3755
rect 3515 3751 3516 3755
rect 3510 3750 3516 3751
rect 3710 3755 3716 3756
rect 3710 3751 3711 3755
rect 3715 3751 3716 3755
rect 3710 3750 3716 3751
rect 3394 3747 3400 3748
rect 2450 3743 2456 3744
rect 2450 3739 2451 3743
rect 2455 3739 2456 3743
rect 2450 3738 2456 3739
rect 2634 3743 2640 3744
rect 2634 3739 2635 3743
rect 2639 3739 2640 3743
rect 2634 3738 2640 3739
rect 2826 3743 2832 3744
rect 2826 3739 2827 3743
rect 2831 3739 2832 3743
rect 2826 3738 2832 3739
rect 3010 3743 3016 3744
rect 3010 3739 3011 3743
rect 3015 3739 3016 3743
rect 3010 3738 3016 3739
rect 3202 3743 3208 3744
rect 3202 3739 3203 3743
rect 3207 3739 3208 3743
rect 3394 3743 3395 3747
rect 3399 3743 3400 3747
rect 3394 3742 3400 3743
rect 3438 3747 3444 3748
rect 3438 3743 3439 3747
rect 3443 3743 3444 3747
rect 3438 3742 3444 3743
rect 3202 3738 3208 3739
rect 2374 3736 2380 3737
rect 2374 3732 2375 3736
rect 2379 3732 2380 3736
rect 2374 3731 2380 3732
rect 2274 3715 2280 3716
rect 2274 3711 2275 3715
rect 2279 3711 2280 3715
rect 2274 3710 2280 3711
rect 2376 3703 2378 3731
rect 2452 3716 2454 3738
rect 2558 3736 2564 3737
rect 2558 3732 2559 3736
rect 2563 3732 2564 3736
rect 2558 3731 2564 3732
rect 2450 3715 2456 3716
rect 2450 3711 2451 3715
rect 2455 3711 2456 3715
rect 2450 3710 2456 3711
rect 2560 3703 2562 3731
rect 2636 3716 2638 3738
rect 2742 3736 2748 3737
rect 2742 3732 2743 3736
rect 2747 3732 2748 3736
rect 2742 3731 2748 3732
rect 2634 3715 2640 3716
rect 2634 3711 2635 3715
rect 2639 3711 2640 3715
rect 2634 3710 2640 3711
rect 2744 3703 2746 3731
rect 2047 3702 2051 3703
rect 2047 3697 2051 3698
rect 2127 3702 2131 3703
rect 2127 3697 2131 3698
rect 2191 3702 2195 3703
rect 2191 3697 2195 3698
rect 2351 3702 2355 3703
rect 2351 3697 2355 3698
rect 2375 3702 2379 3703
rect 2375 3697 2379 3698
rect 2559 3702 2563 3703
rect 2559 3697 2563 3698
rect 2583 3702 2587 3703
rect 2583 3697 2587 3698
rect 2743 3702 2747 3703
rect 2743 3697 2747 3698
rect 2815 3702 2819 3703
rect 2815 3697 2819 3698
rect 2006 3688 2012 3689
rect 1654 3687 1660 3688
rect 1654 3683 1655 3687
rect 1659 3683 1660 3687
rect 2006 3684 2007 3688
rect 2011 3684 2012 3688
rect 2006 3683 2012 3684
rect 1654 3682 1660 3683
rect 1266 3679 1272 3680
rect 1258 3675 1264 3676
rect 1258 3671 1259 3675
rect 1263 3671 1264 3675
rect 1266 3675 1267 3679
rect 1271 3675 1272 3679
rect 1266 3674 1272 3675
rect 1570 3679 1576 3680
rect 1570 3675 1571 3679
rect 1575 3675 1576 3679
rect 1570 3674 1576 3675
rect 1614 3679 1620 3680
rect 1614 3675 1615 3679
rect 1619 3675 1620 3679
rect 1614 3674 1620 3675
rect 1258 3670 1264 3671
rect 1260 3648 1262 3670
rect 1268 3656 1270 3674
rect 1334 3668 1340 3669
rect 1334 3664 1335 3668
rect 1339 3664 1340 3668
rect 1334 3663 1340 3664
rect 1494 3668 1500 3669
rect 1494 3664 1495 3668
rect 1499 3664 1500 3668
rect 1494 3663 1500 3664
rect 1266 3655 1272 3656
rect 1266 3651 1267 3655
rect 1271 3651 1272 3655
rect 1266 3650 1272 3651
rect 1218 3647 1224 3648
rect 1218 3643 1219 3647
rect 1223 3643 1224 3647
rect 1218 3642 1224 3643
rect 1258 3647 1264 3648
rect 1258 3643 1259 3647
rect 1263 3643 1264 3647
rect 1258 3642 1264 3643
rect 1336 3631 1338 3663
rect 1496 3631 1498 3663
rect 1616 3648 1618 3674
rect 2006 3671 2012 3672
rect 1654 3668 1660 3669
rect 1654 3664 1655 3668
rect 1659 3664 1660 3668
rect 2006 3667 2007 3671
rect 2011 3667 2012 3671
rect 2048 3670 2050 3697
rect 2128 3673 2130 3697
rect 2352 3673 2354 3697
rect 2434 3695 2440 3696
rect 2434 3691 2435 3695
rect 2439 3691 2440 3695
rect 2434 3690 2440 3691
rect 2126 3672 2132 3673
rect 2006 3666 2012 3667
rect 2046 3669 2052 3670
rect 1654 3663 1660 3664
rect 1614 3647 1620 3648
rect 1614 3643 1615 3647
rect 1619 3643 1620 3647
rect 1614 3642 1620 3643
rect 1656 3631 1658 3663
rect 1690 3643 1696 3644
rect 1690 3639 1691 3643
rect 1695 3639 1696 3643
rect 1690 3638 1696 3639
rect 1183 3630 1187 3631
rect 1183 3625 1187 3626
rect 1263 3630 1267 3631
rect 1263 3625 1267 3626
rect 1335 3630 1339 3631
rect 1335 3625 1339 3626
rect 1439 3630 1443 3631
rect 1439 3625 1443 3626
rect 1495 3630 1499 3631
rect 1495 3625 1499 3626
rect 1615 3630 1619 3631
rect 1615 3625 1619 3626
rect 1655 3630 1659 3631
rect 1655 3625 1659 3626
rect 1114 3623 1120 3624
rect 1114 3619 1115 3623
rect 1119 3619 1120 3623
rect 1114 3618 1120 3619
rect 1170 3623 1176 3624
rect 1170 3619 1171 3623
rect 1175 3619 1176 3623
rect 1170 3618 1176 3619
rect 926 3600 932 3601
rect 926 3596 927 3600
rect 931 3596 932 3600
rect 926 3595 932 3596
rect 1094 3600 1100 3601
rect 1094 3596 1095 3600
rect 1099 3596 1100 3600
rect 1094 3595 1100 3596
rect 1172 3592 1174 3618
rect 1264 3601 1266 3625
rect 1440 3601 1442 3625
rect 1514 3623 1520 3624
rect 1514 3619 1515 3623
rect 1519 3619 1520 3623
rect 1514 3618 1520 3619
rect 1262 3600 1268 3601
rect 1262 3596 1263 3600
rect 1267 3596 1268 3600
rect 1262 3595 1268 3596
rect 1438 3600 1444 3601
rect 1438 3596 1439 3600
rect 1443 3596 1444 3600
rect 1438 3595 1444 3596
rect 1516 3592 1518 3618
rect 1616 3601 1618 3625
rect 1614 3600 1620 3601
rect 1614 3596 1615 3600
rect 1619 3596 1620 3600
rect 1614 3595 1620 3596
rect 1692 3592 1694 3638
rect 2008 3631 2010 3666
rect 2046 3665 2047 3669
rect 2051 3665 2052 3669
rect 2126 3668 2127 3672
rect 2131 3668 2132 3672
rect 2126 3667 2132 3668
rect 2350 3672 2356 3673
rect 2350 3668 2351 3672
rect 2355 3668 2356 3672
rect 2350 3667 2356 3668
rect 2046 3664 2052 3665
rect 2436 3664 2438 3690
rect 2584 3673 2586 3697
rect 2666 3695 2672 3696
rect 2666 3691 2667 3695
rect 2671 3691 2672 3695
rect 2666 3690 2672 3691
rect 2582 3672 2588 3673
rect 2582 3668 2583 3672
rect 2587 3668 2588 3672
rect 2582 3667 2588 3668
rect 2668 3664 2670 3690
rect 2816 3673 2818 3697
rect 2828 3696 2830 3738
rect 2934 3736 2940 3737
rect 2934 3732 2935 3736
rect 2939 3732 2940 3736
rect 2934 3731 2940 3732
rect 2936 3703 2938 3731
rect 3012 3716 3014 3738
rect 3126 3736 3132 3737
rect 3126 3732 3127 3736
rect 3131 3732 3132 3736
rect 3126 3731 3132 3732
rect 3010 3715 3016 3716
rect 3010 3711 3011 3715
rect 3015 3711 3016 3715
rect 3010 3710 3016 3711
rect 3128 3703 3130 3731
rect 3204 3716 3206 3738
rect 3318 3736 3324 3737
rect 3318 3732 3319 3736
rect 3323 3732 3324 3736
rect 3318 3731 3324 3732
rect 3202 3715 3208 3716
rect 3202 3711 3203 3715
rect 3207 3711 3208 3715
rect 3202 3710 3208 3711
rect 3320 3703 3322 3731
rect 3440 3724 3442 3742
rect 3510 3736 3516 3737
rect 3510 3732 3511 3736
rect 3515 3732 3516 3736
rect 3510 3731 3516 3732
rect 3710 3736 3716 3737
rect 3710 3732 3711 3736
rect 3715 3732 3716 3736
rect 3710 3731 3716 3732
rect 3438 3723 3444 3724
rect 3438 3719 3439 3723
rect 3443 3719 3444 3723
rect 3438 3718 3444 3719
rect 3512 3703 3514 3731
rect 3578 3711 3584 3712
rect 3578 3707 3579 3711
rect 3583 3707 3584 3711
rect 3578 3706 3584 3707
rect 2935 3702 2939 3703
rect 2935 3697 2939 3698
rect 3047 3702 3051 3703
rect 3047 3697 3051 3698
rect 3127 3702 3131 3703
rect 3127 3697 3131 3698
rect 3279 3702 3283 3703
rect 3279 3697 3283 3698
rect 3319 3702 3323 3703
rect 3319 3697 3323 3698
rect 3511 3702 3515 3703
rect 3511 3697 3515 3698
rect 2826 3695 2832 3696
rect 2826 3691 2827 3695
rect 2831 3691 2832 3695
rect 2826 3690 2832 3691
rect 3048 3673 3050 3697
rect 3142 3695 3148 3696
rect 3142 3691 3143 3695
rect 3147 3691 3148 3695
rect 3142 3690 3148 3691
rect 2814 3672 2820 3673
rect 2814 3668 2815 3672
rect 2819 3668 2820 3672
rect 2814 3667 2820 3668
rect 3046 3672 3052 3673
rect 3046 3668 3047 3672
rect 3051 3668 3052 3672
rect 3046 3667 3052 3668
rect 3144 3664 3146 3690
rect 3280 3673 3282 3697
rect 3354 3695 3360 3696
rect 3354 3691 3355 3695
rect 3359 3691 3360 3695
rect 3354 3690 3360 3691
rect 3278 3672 3284 3673
rect 3278 3668 3279 3672
rect 3283 3668 3284 3672
rect 3278 3667 3284 3668
rect 3356 3664 3358 3690
rect 3378 3687 3384 3688
rect 3378 3683 3379 3687
rect 3383 3683 3384 3687
rect 3378 3682 3384 3683
rect 2202 3663 2208 3664
rect 2202 3659 2203 3663
rect 2207 3659 2208 3663
rect 2202 3658 2208 3659
rect 2434 3663 2440 3664
rect 2434 3659 2435 3663
rect 2439 3659 2440 3663
rect 2434 3658 2440 3659
rect 2666 3663 2672 3664
rect 2666 3659 2667 3663
rect 2671 3659 2672 3663
rect 2666 3658 2672 3659
rect 3142 3663 3148 3664
rect 3142 3659 3143 3663
rect 3147 3659 3148 3663
rect 3142 3658 3148 3659
rect 3354 3663 3360 3664
rect 3354 3659 3355 3663
rect 3359 3659 3360 3663
rect 3354 3658 3360 3659
rect 2126 3653 2132 3654
rect 2046 3652 2052 3653
rect 2046 3648 2047 3652
rect 2051 3648 2052 3652
rect 2126 3649 2127 3653
rect 2131 3649 2132 3653
rect 2126 3648 2132 3649
rect 2046 3647 2052 3648
rect 1791 3630 1795 3631
rect 1791 3625 1795 3626
rect 2007 3630 2011 3631
rect 2007 3625 2011 3626
rect 1758 3615 1764 3616
rect 1758 3611 1759 3615
rect 1763 3611 1764 3615
rect 1758 3610 1764 3611
rect 1760 3592 1762 3610
rect 1792 3601 1794 3625
rect 1846 3623 1852 3624
rect 1846 3619 1847 3623
rect 1851 3619 1852 3623
rect 1846 3618 1852 3619
rect 1790 3600 1796 3601
rect 1790 3596 1791 3600
rect 1795 3596 1796 3600
rect 1790 3595 1796 3596
rect 834 3591 840 3592
rect 834 3587 835 3591
rect 839 3587 840 3591
rect 834 3586 840 3587
rect 858 3591 864 3592
rect 858 3587 859 3591
rect 863 3587 864 3591
rect 858 3586 864 3587
rect 1170 3591 1176 3592
rect 1170 3587 1171 3591
rect 1175 3587 1176 3591
rect 1170 3586 1176 3587
rect 1338 3591 1344 3592
rect 1338 3587 1339 3591
rect 1343 3587 1344 3591
rect 1338 3586 1344 3587
rect 1514 3591 1520 3592
rect 1514 3587 1515 3591
rect 1519 3587 1520 3591
rect 1514 3586 1520 3587
rect 1690 3591 1696 3592
rect 1690 3587 1691 3591
rect 1695 3587 1696 3591
rect 1690 3586 1696 3587
rect 1758 3591 1764 3592
rect 1758 3587 1759 3591
rect 1763 3587 1764 3591
rect 1758 3586 1764 3587
rect 758 3581 764 3582
rect 758 3577 759 3581
rect 763 3577 764 3581
rect 758 3576 764 3577
rect 926 3581 932 3582
rect 926 3577 927 3581
rect 931 3577 932 3581
rect 926 3576 932 3577
rect 1094 3581 1100 3582
rect 1094 3577 1095 3581
rect 1099 3577 1100 3581
rect 1094 3576 1100 3577
rect 1262 3581 1268 3582
rect 1262 3577 1263 3581
rect 1267 3577 1268 3581
rect 1262 3576 1268 3577
rect 760 3543 762 3576
rect 928 3543 930 3576
rect 1096 3543 1098 3576
rect 1264 3543 1266 3576
rect 759 3542 763 3543
rect 759 3537 763 3538
rect 815 3542 819 3543
rect 815 3537 819 3538
rect 927 3542 931 3543
rect 927 3537 931 3538
rect 999 3542 1003 3543
rect 999 3537 1003 3538
rect 1095 3542 1099 3543
rect 1095 3537 1099 3538
rect 1175 3542 1179 3543
rect 1175 3537 1179 3538
rect 1263 3542 1267 3543
rect 1263 3537 1267 3538
rect 816 3516 818 3537
rect 1000 3516 1002 3537
rect 1176 3516 1178 3537
rect 814 3515 820 3516
rect 814 3511 815 3515
rect 819 3511 820 3515
rect 814 3510 820 3511
rect 998 3515 1004 3516
rect 998 3511 999 3515
rect 1003 3511 1004 3515
rect 998 3510 1004 3511
rect 1174 3515 1180 3516
rect 1174 3511 1175 3515
rect 1179 3511 1180 3515
rect 1174 3510 1180 3511
rect 738 3507 744 3508
rect 234 3503 240 3504
rect 110 3499 116 3500
rect 110 3495 111 3499
rect 115 3495 116 3499
rect 234 3499 235 3503
rect 239 3499 240 3503
rect 234 3498 240 3499
rect 378 3503 384 3504
rect 378 3499 379 3503
rect 383 3499 384 3503
rect 378 3498 384 3499
rect 538 3503 544 3504
rect 538 3499 539 3503
rect 543 3499 544 3503
rect 538 3498 544 3499
rect 714 3503 720 3504
rect 714 3499 715 3503
rect 719 3499 720 3503
rect 738 3503 739 3507
rect 743 3503 744 3507
rect 1082 3507 1088 3508
rect 738 3502 744 3503
rect 1074 3503 1080 3504
rect 714 3498 720 3499
rect 1074 3499 1075 3503
rect 1079 3499 1080 3503
rect 1082 3503 1083 3507
rect 1087 3503 1088 3507
rect 1082 3502 1088 3503
rect 1074 3498 1080 3499
rect 110 3494 116 3495
rect 158 3496 164 3497
rect 112 3459 114 3494
rect 158 3492 159 3496
rect 163 3492 164 3496
rect 158 3491 164 3492
rect 160 3459 162 3491
rect 236 3480 238 3498
rect 302 3496 308 3497
rect 302 3492 303 3496
rect 307 3492 308 3496
rect 302 3491 308 3492
rect 234 3479 240 3480
rect 234 3475 235 3479
rect 239 3475 240 3479
rect 234 3474 240 3475
rect 304 3459 306 3491
rect 380 3476 382 3498
rect 462 3496 468 3497
rect 462 3492 463 3496
rect 467 3492 468 3496
rect 462 3491 468 3492
rect 378 3475 384 3476
rect 378 3471 379 3475
rect 383 3471 384 3475
rect 378 3470 384 3471
rect 464 3459 466 3491
rect 540 3476 542 3498
rect 638 3496 644 3497
rect 638 3492 639 3496
rect 643 3492 644 3496
rect 638 3491 644 3492
rect 538 3475 544 3476
rect 538 3471 539 3475
rect 543 3471 544 3475
rect 538 3470 544 3471
rect 640 3459 642 3491
rect 716 3476 718 3498
rect 814 3496 820 3497
rect 814 3492 815 3496
rect 819 3492 820 3496
rect 814 3491 820 3492
rect 998 3496 1004 3497
rect 998 3492 999 3496
rect 1003 3492 1004 3496
rect 998 3491 1004 3492
rect 714 3475 720 3476
rect 714 3471 715 3475
rect 719 3471 720 3475
rect 714 3470 720 3471
rect 678 3467 684 3468
rect 678 3463 679 3467
rect 683 3463 684 3467
rect 678 3462 684 3463
rect 111 3458 115 3459
rect 111 3453 115 3454
rect 135 3458 139 3459
rect 135 3453 139 3454
rect 159 3458 163 3459
rect 159 3453 163 3454
rect 303 3458 307 3459
rect 303 3453 307 3454
rect 319 3458 323 3459
rect 319 3453 323 3454
rect 463 3458 467 3459
rect 463 3453 467 3454
rect 535 3458 539 3459
rect 535 3453 539 3454
rect 639 3458 643 3459
rect 639 3453 643 3454
rect 112 3426 114 3453
rect 136 3429 138 3453
rect 254 3451 260 3452
rect 254 3447 255 3451
rect 259 3447 260 3451
rect 254 3446 260 3447
rect 262 3451 268 3452
rect 262 3447 263 3451
rect 267 3447 268 3451
rect 262 3446 268 3447
rect 256 3429 258 3446
rect 134 3428 140 3429
rect 110 3425 116 3426
rect 110 3421 111 3425
rect 115 3421 116 3425
rect 134 3424 135 3428
rect 139 3424 140 3428
rect 134 3423 140 3424
rect 255 3428 259 3429
rect 255 3423 259 3424
rect 110 3420 116 3421
rect 264 3420 266 3446
rect 320 3429 322 3453
rect 394 3451 400 3452
rect 394 3447 395 3451
rect 399 3447 400 3451
rect 394 3446 400 3447
rect 318 3428 324 3429
rect 318 3424 319 3428
rect 323 3424 324 3428
rect 318 3423 324 3424
rect 396 3420 398 3446
rect 536 3429 538 3453
rect 610 3451 616 3452
rect 610 3447 611 3451
rect 615 3447 616 3451
rect 610 3446 616 3447
rect 534 3428 540 3429
rect 534 3424 535 3428
rect 539 3424 540 3428
rect 534 3423 540 3424
rect 612 3420 614 3446
rect 680 3420 682 3462
rect 816 3459 818 3491
rect 1000 3459 1002 3491
rect 751 3458 755 3459
rect 751 3453 755 3454
rect 815 3458 819 3459
rect 815 3453 819 3454
rect 959 3458 963 3459
rect 959 3453 963 3454
rect 999 3458 1003 3459
rect 999 3453 1003 3454
rect 752 3429 754 3453
rect 960 3429 962 3453
rect 1076 3452 1078 3498
rect 1084 3476 1086 3502
rect 1174 3496 1180 3497
rect 1174 3492 1175 3496
rect 1179 3492 1180 3496
rect 1174 3491 1180 3492
rect 1082 3475 1088 3476
rect 1082 3471 1083 3475
rect 1087 3471 1088 3475
rect 1082 3470 1088 3471
rect 1176 3459 1178 3491
rect 1340 3476 1342 3586
rect 1438 3581 1444 3582
rect 1438 3577 1439 3581
rect 1443 3577 1444 3581
rect 1438 3576 1444 3577
rect 1614 3581 1620 3582
rect 1614 3577 1615 3581
rect 1619 3577 1620 3581
rect 1614 3576 1620 3577
rect 1790 3581 1796 3582
rect 1790 3577 1791 3581
rect 1795 3577 1796 3581
rect 1790 3576 1796 3577
rect 1440 3543 1442 3576
rect 1616 3543 1618 3576
rect 1792 3543 1794 3576
rect 1351 3542 1355 3543
rect 1351 3537 1355 3538
rect 1439 3542 1443 3543
rect 1439 3537 1443 3538
rect 1527 3542 1531 3543
rect 1527 3537 1531 3538
rect 1615 3542 1619 3543
rect 1615 3537 1619 3538
rect 1703 3542 1707 3543
rect 1703 3537 1707 3538
rect 1791 3542 1795 3543
rect 1791 3537 1795 3538
rect 1352 3516 1354 3537
rect 1528 3516 1530 3537
rect 1704 3516 1706 3537
rect 1350 3515 1356 3516
rect 1350 3511 1351 3515
rect 1355 3511 1356 3515
rect 1350 3510 1356 3511
rect 1526 3515 1532 3516
rect 1526 3511 1527 3515
rect 1531 3511 1532 3515
rect 1526 3510 1532 3511
rect 1702 3515 1708 3516
rect 1702 3511 1703 3515
rect 1707 3511 1708 3515
rect 1702 3510 1708 3511
rect 1848 3508 1850 3618
rect 2008 3598 2010 3625
rect 2048 3619 2050 3647
rect 2128 3619 2130 3648
rect 2047 3618 2051 3619
rect 2047 3613 2051 3614
rect 2127 3618 2131 3619
rect 2127 3613 2131 3614
rect 2191 3618 2195 3619
rect 2191 3613 2195 3614
rect 2006 3597 2012 3598
rect 2006 3593 2007 3597
rect 2011 3593 2012 3597
rect 2048 3593 2050 3613
rect 2006 3592 2012 3593
rect 2046 3592 2052 3593
rect 2192 3592 2194 3613
rect 2046 3588 2047 3592
rect 2051 3588 2052 3592
rect 2046 3587 2052 3588
rect 2190 3591 2196 3592
rect 2190 3587 2191 3591
rect 2195 3587 2196 3591
rect 2190 3586 2196 3587
rect 2006 3580 2012 3581
rect 2006 3576 2007 3580
rect 2011 3576 2012 3580
rect 2006 3575 2012 3576
rect 2046 3575 2052 3576
rect 2008 3543 2010 3575
rect 2046 3571 2047 3575
rect 2051 3571 2052 3575
rect 2046 3570 2052 3571
rect 2190 3572 2196 3573
rect 2048 3543 2050 3570
rect 2190 3568 2191 3572
rect 2195 3568 2196 3572
rect 2190 3567 2196 3568
rect 2192 3543 2194 3567
rect 2204 3552 2206 3658
rect 2350 3653 2356 3654
rect 2350 3649 2351 3653
rect 2355 3649 2356 3653
rect 2350 3648 2356 3649
rect 2582 3653 2588 3654
rect 2582 3649 2583 3653
rect 2587 3649 2588 3653
rect 2582 3648 2588 3649
rect 2814 3653 2820 3654
rect 2814 3649 2815 3653
rect 2819 3649 2820 3653
rect 2814 3648 2820 3649
rect 3046 3653 3052 3654
rect 3046 3649 3047 3653
rect 3051 3649 3052 3653
rect 3046 3648 3052 3649
rect 3278 3653 3284 3654
rect 3278 3649 3279 3653
rect 3283 3649 3284 3653
rect 3278 3648 3284 3649
rect 2352 3619 2354 3648
rect 2584 3619 2586 3648
rect 2816 3619 2818 3648
rect 3048 3619 3050 3648
rect 3280 3619 3282 3648
rect 2327 3618 2331 3619
rect 2327 3613 2331 3614
rect 2351 3618 2355 3619
rect 2351 3613 2355 3614
rect 2455 3618 2459 3619
rect 2455 3613 2459 3614
rect 2583 3618 2587 3619
rect 2583 3613 2587 3614
rect 2719 3618 2723 3619
rect 2719 3613 2723 3614
rect 2815 3618 2819 3619
rect 2815 3613 2819 3614
rect 2855 3618 2859 3619
rect 2855 3613 2859 3614
rect 2999 3618 3003 3619
rect 2999 3613 3003 3614
rect 3047 3618 3051 3619
rect 3047 3613 3051 3614
rect 3143 3618 3147 3619
rect 3143 3613 3147 3614
rect 3279 3618 3283 3619
rect 3279 3613 3283 3614
rect 3295 3618 3299 3619
rect 3295 3613 3299 3614
rect 2328 3592 2330 3613
rect 2456 3592 2458 3613
rect 2584 3592 2586 3613
rect 2720 3592 2722 3613
rect 2856 3592 2858 3613
rect 3000 3592 3002 3613
rect 3144 3592 3146 3613
rect 3296 3592 3298 3613
rect 2326 3591 2332 3592
rect 2326 3587 2327 3591
rect 2331 3587 2332 3591
rect 2326 3586 2332 3587
rect 2454 3591 2460 3592
rect 2454 3587 2455 3591
rect 2459 3587 2460 3591
rect 2454 3586 2460 3587
rect 2582 3591 2588 3592
rect 2582 3587 2583 3591
rect 2587 3587 2588 3591
rect 2582 3586 2588 3587
rect 2718 3591 2724 3592
rect 2718 3587 2719 3591
rect 2723 3587 2724 3591
rect 2718 3586 2724 3587
rect 2854 3591 2860 3592
rect 2854 3587 2855 3591
rect 2859 3587 2860 3591
rect 2854 3586 2860 3587
rect 2998 3591 3004 3592
rect 2998 3587 2999 3591
rect 3003 3587 3004 3591
rect 2998 3586 3004 3587
rect 3142 3591 3148 3592
rect 3142 3587 3143 3591
rect 3147 3587 3148 3591
rect 3142 3586 3148 3587
rect 3294 3591 3300 3592
rect 3294 3587 3295 3591
rect 3299 3587 3300 3591
rect 3294 3586 3300 3587
rect 3380 3584 3382 3682
rect 3512 3673 3514 3697
rect 3510 3672 3516 3673
rect 3510 3668 3511 3672
rect 3515 3668 3516 3672
rect 3510 3667 3516 3668
rect 3580 3664 3582 3706
rect 3712 3703 3714 3731
rect 3732 3716 3734 3814
rect 3942 3808 3948 3809
rect 3942 3804 3943 3808
rect 3947 3804 3948 3808
rect 3942 3803 3948 3804
rect 3944 3783 3946 3803
rect 3943 3782 3947 3783
rect 3943 3777 3947 3778
rect 3944 3757 3946 3777
rect 3942 3756 3948 3757
rect 3942 3752 3943 3756
rect 3947 3752 3948 3756
rect 3942 3751 3948 3752
rect 3786 3743 3792 3744
rect 3786 3739 3787 3743
rect 3791 3739 3792 3743
rect 3786 3738 3792 3739
rect 3942 3739 3948 3740
rect 3730 3715 3736 3716
rect 3730 3711 3731 3715
rect 3735 3711 3736 3715
rect 3730 3710 3736 3711
rect 3711 3702 3715 3703
rect 3711 3697 3715 3698
rect 3751 3702 3755 3703
rect 3751 3697 3755 3698
rect 3752 3673 3754 3697
rect 3788 3696 3790 3738
rect 3942 3735 3943 3739
rect 3947 3735 3948 3739
rect 3942 3734 3948 3735
rect 3944 3703 3946 3734
rect 3943 3702 3947 3703
rect 3943 3697 3947 3698
rect 3786 3695 3792 3696
rect 3786 3691 3787 3695
rect 3791 3691 3792 3695
rect 3786 3690 3792 3691
rect 3750 3672 3756 3673
rect 3750 3668 3751 3672
rect 3755 3668 3756 3672
rect 3944 3670 3946 3697
rect 3750 3667 3756 3668
rect 3942 3669 3948 3670
rect 3942 3665 3943 3669
rect 3947 3665 3948 3669
rect 3942 3664 3948 3665
rect 3578 3663 3584 3664
rect 3578 3659 3579 3663
rect 3583 3659 3584 3663
rect 3578 3658 3584 3659
rect 3826 3663 3832 3664
rect 3826 3659 3827 3663
rect 3831 3659 3832 3663
rect 3826 3658 3832 3659
rect 3510 3653 3516 3654
rect 3510 3649 3511 3653
rect 3515 3649 3516 3653
rect 3510 3648 3516 3649
rect 3750 3653 3756 3654
rect 3750 3649 3751 3653
rect 3755 3649 3756 3653
rect 3750 3648 3756 3649
rect 3512 3619 3514 3648
rect 3752 3619 3754 3648
rect 3455 3618 3459 3619
rect 3455 3613 3459 3614
rect 3511 3618 3515 3619
rect 3511 3613 3515 3614
rect 3623 3618 3627 3619
rect 3623 3613 3627 3614
rect 3751 3618 3755 3619
rect 3751 3613 3755 3614
rect 3456 3592 3458 3613
rect 3624 3592 3626 3613
rect 3454 3591 3460 3592
rect 3454 3587 3455 3591
rect 3459 3587 3460 3591
rect 3454 3586 3460 3587
rect 3622 3591 3628 3592
rect 3622 3587 3623 3591
rect 3627 3587 3628 3591
rect 3622 3586 3628 3587
rect 3258 3583 3264 3584
rect 2278 3579 2284 3580
rect 2278 3575 2279 3579
rect 2283 3575 2284 3579
rect 2278 3574 2284 3575
rect 2530 3579 2536 3580
rect 2530 3575 2531 3579
rect 2535 3575 2536 3579
rect 2530 3574 2536 3575
rect 2658 3579 2664 3580
rect 2658 3575 2659 3579
rect 2663 3575 2664 3579
rect 2658 3574 2664 3575
rect 2794 3579 2800 3580
rect 2794 3575 2795 3579
rect 2799 3575 2800 3579
rect 2794 3574 2800 3575
rect 2930 3579 2936 3580
rect 2930 3575 2931 3579
rect 2935 3575 2936 3579
rect 2930 3574 2936 3575
rect 3074 3579 3080 3580
rect 3074 3575 3075 3579
rect 3079 3575 3080 3579
rect 3074 3574 3080 3575
rect 3218 3579 3224 3580
rect 3218 3575 3219 3579
rect 3223 3575 3224 3579
rect 3258 3579 3259 3583
rect 3263 3579 3264 3583
rect 3258 3578 3264 3579
rect 3378 3583 3384 3584
rect 3378 3579 3379 3583
rect 3383 3579 3384 3583
rect 3378 3578 3384 3579
rect 3586 3583 3592 3584
rect 3586 3579 3587 3583
rect 3591 3579 3592 3583
rect 3586 3578 3592 3579
rect 3218 3574 3224 3575
rect 2202 3551 2208 3552
rect 2202 3547 2203 3551
rect 2207 3547 2208 3551
rect 2202 3546 2208 3547
rect 1879 3542 1883 3543
rect 1879 3537 1883 3538
rect 2007 3542 2011 3543
rect 2007 3537 2011 3538
rect 2047 3542 2051 3543
rect 2047 3537 2051 3538
rect 2103 3542 2107 3543
rect 2103 3537 2107 3538
rect 2191 3542 2195 3543
rect 2191 3537 2195 3538
rect 2271 3542 2275 3543
rect 2271 3537 2275 3538
rect 1880 3516 1882 3537
rect 2008 3517 2010 3537
rect 2006 3516 2012 3517
rect 1878 3515 1884 3516
rect 1878 3511 1879 3515
rect 1883 3511 1884 3515
rect 2006 3512 2007 3516
rect 2011 3512 2012 3516
rect 2006 3511 2012 3512
rect 1878 3510 1884 3511
rect 2048 3510 2050 3537
rect 2104 3513 2106 3537
rect 2272 3513 2274 3537
rect 2280 3536 2282 3574
rect 2326 3572 2332 3573
rect 2326 3568 2327 3572
rect 2331 3568 2332 3572
rect 2326 3567 2332 3568
rect 2454 3572 2460 3573
rect 2454 3568 2455 3572
rect 2459 3568 2460 3572
rect 2454 3567 2460 3568
rect 2328 3543 2330 3567
rect 2456 3543 2458 3567
rect 2532 3552 2534 3574
rect 2582 3572 2588 3573
rect 2582 3568 2583 3572
rect 2587 3568 2588 3572
rect 2582 3567 2588 3568
rect 2530 3551 2536 3552
rect 2530 3547 2531 3551
rect 2535 3547 2536 3551
rect 2530 3546 2536 3547
rect 2584 3543 2586 3567
rect 2660 3552 2662 3574
rect 2718 3572 2724 3573
rect 2718 3568 2719 3572
rect 2723 3568 2724 3572
rect 2718 3567 2724 3568
rect 2658 3551 2664 3552
rect 2658 3547 2659 3551
rect 2663 3547 2664 3551
rect 2658 3546 2664 3547
rect 2720 3543 2722 3567
rect 2796 3552 2798 3574
rect 2854 3572 2860 3573
rect 2854 3568 2855 3572
rect 2859 3568 2860 3572
rect 2854 3567 2860 3568
rect 2794 3551 2800 3552
rect 2794 3547 2795 3551
rect 2799 3547 2800 3551
rect 2794 3546 2800 3547
rect 2856 3543 2858 3567
rect 2932 3552 2934 3574
rect 2998 3572 3004 3573
rect 2998 3568 2999 3572
rect 3003 3568 3004 3572
rect 2998 3567 3004 3568
rect 2930 3551 2936 3552
rect 2930 3547 2931 3551
rect 2935 3547 2936 3551
rect 2930 3546 2936 3547
rect 3000 3543 3002 3567
rect 3076 3552 3078 3574
rect 3142 3572 3148 3573
rect 3142 3568 3143 3572
rect 3147 3568 3148 3572
rect 3142 3567 3148 3568
rect 3074 3551 3080 3552
rect 3074 3547 3075 3551
rect 3079 3547 3080 3551
rect 3074 3546 3080 3547
rect 3144 3543 3146 3567
rect 3220 3552 3222 3574
rect 3218 3551 3224 3552
rect 3218 3547 3219 3551
rect 3223 3547 3224 3551
rect 3218 3546 3224 3547
rect 3260 3544 3262 3578
rect 3294 3572 3300 3573
rect 3294 3568 3295 3572
rect 3299 3568 3300 3572
rect 3294 3567 3300 3568
rect 3454 3572 3460 3573
rect 3454 3568 3455 3572
rect 3459 3568 3460 3572
rect 3454 3567 3460 3568
rect 3258 3543 3264 3544
rect 3296 3543 3298 3567
rect 3456 3543 3458 3567
rect 3588 3552 3590 3578
rect 3622 3572 3628 3573
rect 3622 3568 3623 3572
rect 3627 3568 3628 3572
rect 3622 3567 3628 3568
rect 3586 3551 3592 3552
rect 3586 3547 3587 3551
rect 3591 3547 3592 3551
rect 3586 3546 3592 3547
rect 3594 3547 3600 3548
rect 3594 3543 3595 3547
rect 3599 3543 3600 3547
rect 3624 3543 3626 3567
rect 2327 3542 2331 3543
rect 2327 3537 2331 3538
rect 2447 3542 2451 3543
rect 2447 3537 2451 3538
rect 2455 3542 2459 3543
rect 2455 3537 2459 3538
rect 2583 3542 2587 3543
rect 2583 3537 2587 3538
rect 2631 3542 2635 3543
rect 2631 3537 2635 3538
rect 2719 3542 2723 3543
rect 2719 3537 2723 3538
rect 2815 3542 2819 3543
rect 2815 3537 2819 3538
rect 2855 3542 2859 3543
rect 2855 3537 2859 3538
rect 2999 3542 3003 3543
rect 2999 3537 3003 3538
rect 3143 3542 3147 3543
rect 3143 3537 3147 3538
rect 3175 3542 3179 3543
rect 3258 3539 3259 3543
rect 3263 3539 3264 3543
rect 3258 3538 3264 3539
rect 3295 3542 3299 3543
rect 3175 3537 3179 3538
rect 3295 3537 3299 3538
rect 3351 3542 3355 3543
rect 3351 3537 3355 3538
rect 3455 3542 3459 3543
rect 3455 3537 3459 3538
rect 3519 3542 3523 3543
rect 3594 3542 3600 3543
rect 3623 3542 3627 3543
rect 3519 3537 3523 3538
rect 2278 3535 2284 3536
rect 2278 3531 2279 3535
rect 2283 3531 2284 3535
rect 2278 3530 2284 3531
rect 2448 3513 2450 3537
rect 2530 3535 2536 3536
rect 2530 3531 2531 3535
rect 2535 3531 2536 3535
rect 2530 3530 2536 3531
rect 2102 3512 2108 3513
rect 2046 3509 2052 3510
rect 1846 3507 1852 3508
rect 1662 3503 1668 3504
rect 1662 3499 1663 3503
rect 1667 3499 1668 3503
rect 1662 3498 1668 3499
rect 1778 3503 1784 3504
rect 1778 3499 1779 3503
rect 1783 3499 1784 3503
rect 1846 3503 1847 3507
rect 1851 3503 1852 3507
rect 2046 3505 2047 3509
rect 2051 3505 2052 3509
rect 2102 3508 2103 3512
rect 2107 3508 2108 3512
rect 2102 3507 2108 3508
rect 2270 3512 2276 3513
rect 2270 3508 2271 3512
rect 2275 3508 2276 3512
rect 2270 3507 2276 3508
rect 2446 3512 2452 3513
rect 2446 3508 2447 3512
rect 2451 3508 2452 3512
rect 2446 3507 2452 3508
rect 2046 3504 2052 3505
rect 2532 3504 2534 3530
rect 2632 3513 2634 3537
rect 2778 3535 2784 3536
rect 2778 3531 2779 3535
rect 2783 3531 2784 3535
rect 2778 3530 2784 3531
rect 2630 3512 2636 3513
rect 2630 3508 2631 3512
rect 2635 3508 2636 3512
rect 2630 3507 2636 3508
rect 1846 3502 1852 3503
rect 2178 3503 2184 3504
rect 1778 3498 1784 3499
rect 2006 3499 2012 3500
rect 1350 3496 1356 3497
rect 1350 3492 1351 3496
rect 1355 3492 1356 3496
rect 1350 3491 1356 3492
rect 1526 3496 1532 3497
rect 1526 3492 1527 3496
rect 1531 3492 1532 3496
rect 1526 3491 1532 3492
rect 1338 3475 1344 3476
rect 1338 3471 1339 3475
rect 1343 3471 1344 3475
rect 1338 3470 1344 3471
rect 1352 3459 1354 3491
rect 1528 3459 1530 3491
rect 1664 3476 1666 3498
rect 1702 3496 1708 3497
rect 1702 3492 1703 3496
rect 1707 3492 1708 3496
rect 1702 3491 1708 3492
rect 1662 3475 1668 3476
rect 1602 3471 1608 3472
rect 1602 3467 1603 3471
rect 1607 3467 1608 3471
rect 1662 3471 1663 3475
rect 1667 3471 1668 3475
rect 1662 3470 1668 3471
rect 1602 3466 1608 3467
rect 1159 3458 1163 3459
rect 1159 3453 1163 3454
rect 1175 3458 1179 3459
rect 1175 3453 1179 3454
rect 1351 3458 1355 3459
rect 1351 3453 1355 3454
rect 1527 3458 1531 3459
rect 1527 3453 1531 3454
rect 1535 3458 1539 3459
rect 1535 3453 1539 3454
rect 1074 3451 1080 3452
rect 1074 3447 1075 3451
rect 1079 3447 1080 3451
rect 1074 3446 1080 3447
rect 1082 3451 1088 3452
rect 1082 3447 1083 3451
rect 1087 3447 1088 3451
rect 1082 3446 1088 3447
rect 750 3428 756 3429
rect 750 3424 751 3428
rect 755 3424 756 3428
rect 750 3423 756 3424
rect 799 3428 803 3429
rect 799 3423 803 3424
rect 958 3428 964 3429
rect 958 3424 959 3428
rect 963 3424 964 3428
rect 958 3423 964 3424
rect 262 3419 268 3420
rect 262 3415 263 3419
rect 267 3415 268 3419
rect 262 3414 268 3415
rect 394 3419 400 3420
rect 394 3415 395 3419
rect 399 3415 400 3419
rect 394 3414 400 3415
rect 610 3419 616 3420
rect 610 3415 611 3419
rect 615 3415 616 3419
rect 610 3414 616 3415
rect 678 3419 684 3420
rect 678 3415 679 3419
rect 683 3415 684 3419
rect 678 3414 684 3415
rect 134 3409 140 3410
rect 110 3408 116 3409
rect 110 3404 111 3408
rect 115 3404 116 3408
rect 134 3405 135 3409
rect 139 3405 140 3409
rect 134 3404 140 3405
rect 318 3409 324 3410
rect 318 3405 319 3409
rect 323 3405 324 3409
rect 318 3404 324 3405
rect 534 3409 540 3410
rect 534 3405 535 3409
rect 539 3405 540 3409
rect 534 3404 540 3405
rect 750 3409 756 3410
rect 750 3405 751 3409
rect 755 3405 756 3409
rect 750 3404 756 3405
rect 110 3403 116 3404
rect 112 3383 114 3403
rect 136 3383 138 3404
rect 320 3383 322 3404
rect 536 3383 538 3404
rect 752 3383 754 3404
rect 111 3382 115 3383
rect 111 3377 115 3378
rect 135 3382 139 3383
rect 135 3377 139 3378
rect 231 3382 235 3383
rect 231 3377 235 3378
rect 319 3382 323 3383
rect 319 3377 323 3378
rect 375 3382 379 3383
rect 375 3377 379 3378
rect 535 3382 539 3383
rect 535 3377 539 3378
rect 703 3382 707 3383
rect 703 3377 707 3378
rect 751 3382 755 3383
rect 751 3377 755 3378
rect 112 3357 114 3377
rect 110 3356 116 3357
rect 136 3356 138 3377
rect 232 3356 234 3377
rect 376 3356 378 3377
rect 536 3356 538 3377
rect 704 3356 706 3377
rect 110 3352 111 3356
rect 115 3352 116 3356
rect 110 3351 116 3352
rect 134 3355 140 3356
rect 134 3351 135 3355
rect 139 3351 140 3355
rect 134 3350 140 3351
rect 230 3355 236 3356
rect 230 3351 231 3355
rect 235 3351 236 3355
rect 230 3350 236 3351
rect 374 3355 380 3356
rect 374 3351 375 3355
rect 379 3351 380 3355
rect 374 3350 380 3351
rect 534 3355 540 3356
rect 534 3351 535 3355
rect 539 3351 540 3355
rect 534 3350 540 3351
rect 702 3355 708 3356
rect 702 3351 703 3355
rect 707 3351 708 3355
rect 702 3350 708 3351
rect 800 3348 802 3423
rect 1084 3420 1086 3446
rect 1160 3429 1162 3453
rect 1234 3451 1240 3452
rect 1234 3447 1235 3451
rect 1239 3447 1240 3451
rect 1234 3446 1240 3447
rect 1158 3428 1164 3429
rect 1158 3424 1159 3428
rect 1163 3424 1164 3428
rect 1158 3423 1164 3424
rect 1236 3420 1238 3446
rect 1352 3429 1354 3453
rect 1536 3429 1538 3453
rect 1350 3428 1356 3429
rect 1350 3424 1351 3428
rect 1355 3424 1356 3428
rect 1350 3423 1356 3424
rect 1534 3428 1540 3429
rect 1534 3424 1535 3428
rect 1539 3424 1540 3428
rect 1534 3423 1540 3424
rect 1604 3420 1606 3466
rect 1704 3459 1706 3491
rect 1780 3476 1782 3498
rect 1878 3496 1884 3497
rect 1878 3492 1879 3496
rect 1883 3492 1884 3496
rect 2006 3495 2007 3499
rect 2011 3495 2012 3499
rect 2178 3499 2179 3503
rect 2183 3499 2184 3503
rect 2178 3498 2184 3499
rect 2530 3503 2536 3504
rect 2530 3499 2531 3503
rect 2535 3499 2536 3503
rect 2530 3498 2536 3499
rect 2006 3494 2012 3495
rect 1878 3491 1884 3492
rect 1778 3475 1784 3476
rect 1778 3471 1779 3475
rect 1783 3471 1784 3475
rect 1778 3470 1784 3471
rect 1880 3459 1882 3491
rect 2008 3459 2010 3494
rect 2102 3493 2108 3494
rect 2046 3492 2052 3493
rect 2046 3488 2047 3492
rect 2051 3488 2052 3492
rect 2102 3489 2103 3493
rect 2107 3489 2108 3493
rect 2102 3488 2108 3489
rect 2046 3487 2052 3488
rect 2048 3463 2050 3487
rect 2104 3463 2106 3488
rect 2047 3462 2051 3463
rect 1703 3458 1707 3459
rect 1703 3453 1707 3454
rect 1719 3458 1723 3459
rect 1719 3453 1723 3454
rect 1879 3458 1883 3459
rect 1879 3453 1883 3454
rect 1903 3458 1907 3459
rect 1903 3453 1907 3454
rect 2007 3458 2011 3459
rect 2047 3457 2051 3458
rect 2103 3462 2107 3463
rect 2103 3457 2107 3458
rect 2127 3462 2131 3463
rect 2127 3457 2131 3458
rect 2007 3453 2011 3454
rect 1618 3451 1624 3452
rect 1618 3447 1619 3451
rect 1623 3447 1624 3451
rect 1618 3446 1624 3447
rect 1620 3420 1622 3446
rect 1720 3429 1722 3453
rect 1802 3451 1808 3452
rect 1802 3447 1803 3451
rect 1807 3447 1808 3451
rect 1802 3446 1808 3447
rect 1718 3428 1724 3429
rect 1718 3424 1719 3428
rect 1723 3424 1724 3428
rect 1718 3423 1724 3424
rect 1804 3420 1806 3446
rect 1904 3429 1906 3453
rect 1946 3451 1952 3452
rect 1946 3447 1947 3451
rect 1951 3447 1952 3451
rect 1946 3446 1952 3447
rect 1902 3428 1908 3429
rect 1902 3424 1903 3428
rect 1907 3424 1908 3428
rect 1902 3423 1908 3424
rect 1082 3419 1088 3420
rect 1082 3415 1083 3419
rect 1087 3415 1088 3419
rect 1082 3414 1088 3415
rect 1234 3419 1240 3420
rect 1234 3415 1235 3419
rect 1239 3415 1240 3419
rect 1234 3414 1240 3415
rect 1426 3419 1432 3420
rect 1426 3415 1427 3419
rect 1431 3415 1432 3419
rect 1426 3414 1432 3415
rect 1602 3419 1608 3420
rect 1602 3415 1603 3419
rect 1607 3415 1608 3419
rect 1602 3414 1608 3415
rect 1618 3419 1624 3420
rect 1618 3415 1619 3419
rect 1623 3415 1624 3419
rect 1618 3414 1624 3415
rect 1802 3419 1808 3420
rect 1802 3415 1803 3419
rect 1807 3415 1808 3419
rect 1802 3414 1808 3415
rect 958 3409 964 3410
rect 958 3405 959 3409
rect 963 3405 964 3409
rect 958 3404 964 3405
rect 1158 3409 1164 3410
rect 1158 3405 1159 3409
rect 1163 3405 1164 3409
rect 1158 3404 1164 3405
rect 1350 3409 1356 3410
rect 1350 3405 1351 3409
rect 1355 3405 1356 3409
rect 1350 3404 1356 3405
rect 960 3383 962 3404
rect 1160 3383 1162 3404
rect 1352 3383 1354 3404
rect 871 3382 875 3383
rect 871 3377 875 3378
rect 959 3382 963 3383
rect 959 3377 963 3378
rect 1047 3382 1051 3383
rect 1047 3377 1051 3378
rect 1159 3382 1163 3383
rect 1159 3377 1163 3378
rect 1215 3382 1219 3383
rect 1215 3377 1219 3378
rect 1351 3382 1355 3383
rect 1351 3377 1355 3378
rect 1383 3382 1387 3383
rect 1383 3377 1387 3378
rect 872 3356 874 3377
rect 1048 3356 1050 3377
rect 1216 3356 1218 3377
rect 1384 3356 1386 3377
rect 870 3355 876 3356
rect 870 3351 871 3355
rect 875 3351 876 3355
rect 870 3350 876 3351
rect 1046 3355 1052 3356
rect 1046 3351 1047 3355
rect 1051 3351 1052 3355
rect 1046 3350 1052 3351
rect 1214 3355 1220 3356
rect 1214 3351 1215 3355
rect 1219 3351 1220 3355
rect 1214 3350 1220 3351
rect 1382 3355 1388 3356
rect 1382 3351 1383 3355
rect 1387 3351 1388 3355
rect 1382 3350 1388 3351
rect 798 3347 804 3348
rect 210 3343 216 3344
rect 110 3339 116 3340
rect 110 3335 111 3339
rect 115 3335 116 3339
rect 210 3339 211 3343
rect 215 3339 216 3343
rect 210 3338 216 3339
rect 306 3343 312 3344
rect 306 3339 307 3343
rect 311 3339 312 3343
rect 306 3338 312 3339
rect 450 3343 456 3344
rect 450 3339 451 3343
rect 455 3339 456 3343
rect 450 3338 456 3339
rect 610 3343 616 3344
rect 610 3339 611 3343
rect 615 3339 616 3343
rect 610 3338 616 3339
rect 778 3343 784 3344
rect 778 3339 779 3343
rect 783 3339 784 3343
rect 798 3343 799 3347
rect 803 3343 804 3347
rect 1166 3347 1172 3348
rect 798 3342 804 3343
rect 1122 3343 1128 3344
rect 778 3338 784 3339
rect 1122 3339 1123 3343
rect 1127 3339 1128 3343
rect 1166 3343 1167 3347
rect 1171 3343 1172 3347
rect 1166 3342 1172 3343
rect 1342 3347 1348 3348
rect 1342 3343 1343 3347
rect 1347 3343 1348 3347
rect 1342 3342 1348 3343
rect 1122 3338 1128 3339
rect 110 3334 116 3335
rect 134 3336 140 3337
rect 112 3307 114 3334
rect 134 3332 135 3336
rect 139 3332 140 3336
rect 134 3331 140 3332
rect 136 3307 138 3331
rect 212 3316 214 3338
rect 230 3336 236 3337
rect 230 3332 231 3336
rect 235 3332 236 3336
rect 230 3331 236 3332
rect 210 3315 216 3316
rect 202 3311 208 3312
rect 202 3307 203 3311
rect 207 3307 208 3311
rect 210 3311 211 3315
rect 215 3311 216 3315
rect 210 3310 216 3311
rect 232 3307 234 3331
rect 308 3316 310 3338
rect 374 3336 380 3337
rect 374 3332 375 3336
rect 379 3332 380 3336
rect 374 3331 380 3332
rect 306 3315 312 3316
rect 306 3311 307 3315
rect 311 3311 312 3315
rect 306 3310 312 3311
rect 376 3307 378 3331
rect 452 3316 454 3338
rect 534 3336 540 3337
rect 534 3332 535 3336
rect 539 3332 540 3336
rect 534 3331 540 3332
rect 450 3315 456 3316
rect 450 3311 451 3315
rect 455 3311 456 3315
rect 450 3310 456 3311
rect 536 3307 538 3331
rect 612 3316 614 3338
rect 702 3336 708 3337
rect 702 3332 703 3336
rect 707 3332 708 3336
rect 702 3331 708 3332
rect 610 3315 616 3316
rect 610 3311 611 3315
rect 615 3311 616 3315
rect 610 3310 616 3311
rect 704 3307 706 3331
rect 780 3316 782 3338
rect 870 3336 876 3337
rect 870 3332 871 3336
rect 875 3332 876 3336
rect 870 3331 876 3332
rect 1046 3336 1052 3337
rect 1046 3332 1047 3336
rect 1051 3332 1052 3336
rect 1046 3331 1052 3332
rect 778 3315 784 3316
rect 778 3311 779 3315
rect 783 3311 784 3315
rect 778 3310 784 3311
rect 872 3307 874 3331
rect 1048 3307 1050 3331
rect 111 3306 115 3307
rect 111 3301 115 3302
rect 135 3306 139 3307
rect 202 3306 208 3307
rect 231 3306 235 3307
rect 135 3301 139 3302
rect 112 3274 114 3301
rect 136 3277 138 3301
rect 134 3276 140 3277
rect 110 3273 116 3274
rect 110 3269 111 3273
rect 115 3269 116 3273
rect 134 3272 135 3276
rect 139 3272 140 3276
rect 134 3271 140 3272
rect 110 3268 116 3269
rect 204 3268 206 3306
rect 231 3301 235 3302
rect 279 3306 283 3307
rect 279 3301 283 3302
rect 375 3306 379 3307
rect 375 3301 379 3302
rect 463 3306 467 3307
rect 463 3301 467 3302
rect 535 3306 539 3307
rect 535 3301 539 3302
rect 663 3306 667 3307
rect 663 3301 667 3302
rect 703 3306 707 3307
rect 703 3301 707 3302
rect 871 3306 875 3307
rect 871 3301 875 3302
rect 1047 3306 1051 3307
rect 1047 3301 1051 3302
rect 1079 3306 1083 3307
rect 1079 3301 1083 3302
rect 254 3299 260 3300
rect 254 3295 255 3299
rect 259 3295 260 3299
rect 254 3294 260 3295
rect 256 3268 258 3294
rect 280 3277 282 3301
rect 464 3277 466 3301
rect 518 3299 524 3300
rect 518 3295 519 3299
rect 523 3298 524 3299
rect 523 3295 526 3298
rect 518 3294 526 3295
rect 278 3276 284 3277
rect 278 3272 279 3276
rect 283 3272 284 3276
rect 278 3271 284 3272
rect 462 3276 468 3277
rect 462 3272 463 3276
rect 467 3272 468 3276
rect 462 3271 468 3272
rect 202 3267 208 3268
rect 202 3263 203 3267
rect 207 3263 208 3267
rect 202 3262 208 3263
rect 254 3267 260 3268
rect 254 3263 255 3267
rect 259 3263 260 3267
rect 254 3262 260 3263
rect 134 3257 140 3258
rect 110 3256 116 3257
rect 110 3252 111 3256
rect 115 3252 116 3256
rect 134 3253 135 3257
rect 139 3253 140 3257
rect 134 3252 140 3253
rect 278 3257 284 3258
rect 278 3253 279 3257
rect 283 3253 284 3257
rect 278 3252 284 3253
rect 462 3257 468 3258
rect 462 3253 463 3257
rect 467 3253 468 3257
rect 462 3252 468 3253
rect 110 3251 116 3252
rect 112 3231 114 3251
rect 136 3231 138 3252
rect 280 3231 282 3252
rect 464 3231 466 3252
rect 111 3230 115 3231
rect 111 3225 115 3226
rect 135 3230 139 3231
rect 135 3225 139 3226
rect 279 3230 283 3231
rect 279 3225 283 3226
rect 287 3230 291 3231
rect 287 3225 291 3226
rect 447 3230 451 3231
rect 447 3225 451 3226
rect 463 3230 467 3231
rect 463 3225 467 3226
rect 112 3205 114 3225
rect 110 3204 116 3205
rect 136 3204 138 3225
rect 288 3204 290 3225
rect 448 3204 450 3225
rect 110 3200 111 3204
rect 115 3200 116 3204
rect 110 3199 116 3200
rect 134 3203 140 3204
rect 134 3199 135 3203
rect 139 3199 140 3203
rect 134 3198 140 3199
rect 286 3203 292 3204
rect 286 3199 287 3203
rect 291 3199 292 3203
rect 286 3198 292 3199
rect 446 3203 452 3204
rect 446 3199 447 3203
rect 451 3199 452 3203
rect 446 3198 452 3199
rect 524 3196 526 3294
rect 664 3277 666 3301
rect 738 3299 744 3300
rect 738 3295 739 3299
rect 743 3295 744 3299
rect 738 3294 744 3295
rect 662 3276 668 3277
rect 662 3272 663 3276
rect 667 3272 668 3276
rect 662 3271 668 3272
rect 740 3268 742 3294
rect 798 3287 804 3288
rect 798 3283 799 3287
rect 803 3283 804 3287
rect 798 3282 804 3283
rect 800 3268 802 3282
rect 872 3277 874 3301
rect 1080 3277 1082 3301
rect 1124 3300 1126 3338
rect 1168 3316 1170 3342
rect 1214 3336 1220 3337
rect 1214 3332 1215 3336
rect 1219 3332 1220 3336
rect 1214 3331 1220 3332
rect 1166 3315 1172 3316
rect 1166 3311 1167 3315
rect 1171 3311 1172 3315
rect 1166 3310 1172 3311
rect 1216 3307 1218 3331
rect 1344 3316 1346 3342
rect 1382 3336 1388 3337
rect 1382 3332 1383 3336
rect 1387 3332 1388 3336
rect 1382 3331 1388 3332
rect 1342 3315 1348 3316
rect 1342 3311 1343 3315
rect 1347 3311 1348 3315
rect 1342 3310 1348 3311
rect 1384 3307 1386 3331
rect 1428 3316 1430 3414
rect 1534 3409 1540 3410
rect 1534 3405 1535 3409
rect 1539 3405 1540 3409
rect 1534 3404 1540 3405
rect 1718 3409 1724 3410
rect 1718 3405 1719 3409
rect 1723 3405 1724 3409
rect 1718 3404 1724 3405
rect 1902 3409 1908 3410
rect 1902 3405 1903 3409
rect 1907 3405 1908 3409
rect 1902 3404 1908 3405
rect 1536 3383 1538 3404
rect 1720 3383 1722 3404
rect 1904 3383 1906 3404
rect 1535 3382 1539 3383
rect 1535 3377 1539 3378
rect 1543 3382 1547 3383
rect 1543 3377 1547 3378
rect 1703 3382 1707 3383
rect 1703 3377 1707 3378
rect 1719 3382 1723 3383
rect 1719 3377 1723 3378
rect 1871 3382 1875 3383
rect 1871 3377 1875 3378
rect 1903 3382 1907 3383
rect 1903 3377 1907 3378
rect 1544 3356 1546 3377
rect 1704 3356 1706 3377
rect 1872 3356 1874 3377
rect 1542 3355 1548 3356
rect 1542 3351 1543 3355
rect 1547 3351 1548 3355
rect 1542 3350 1548 3351
rect 1702 3355 1708 3356
rect 1702 3351 1703 3355
rect 1707 3351 1708 3355
rect 1702 3350 1708 3351
rect 1870 3355 1876 3356
rect 1870 3351 1871 3355
rect 1875 3351 1876 3355
rect 1870 3350 1876 3351
rect 1948 3348 1950 3446
rect 2008 3426 2010 3453
rect 2048 3437 2050 3457
rect 2046 3436 2052 3437
rect 2128 3436 2130 3457
rect 2046 3432 2047 3436
rect 2051 3432 2052 3436
rect 2046 3431 2052 3432
rect 2126 3435 2132 3436
rect 2126 3431 2127 3435
rect 2131 3431 2132 3435
rect 2126 3430 2132 3431
rect 2006 3425 2012 3426
rect 2006 3421 2007 3425
rect 2011 3421 2012 3425
rect 2006 3420 2012 3421
rect 2046 3419 2052 3420
rect 2046 3415 2047 3419
rect 2051 3415 2052 3419
rect 2046 3414 2052 3415
rect 2126 3416 2132 3417
rect 2006 3408 2012 3409
rect 2006 3404 2007 3408
rect 2011 3404 2012 3408
rect 2006 3403 2012 3404
rect 2008 3383 2010 3403
rect 2007 3382 2011 3383
rect 2007 3377 2011 3378
rect 2008 3357 2010 3377
rect 2048 3371 2050 3414
rect 2126 3412 2127 3416
rect 2131 3412 2132 3416
rect 2126 3411 2132 3412
rect 2128 3371 2130 3411
rect 2180 3396 2182 3498
rect 2270 3493 2276 3494
rect 2270 3489 2271 3493
rect 2275 3489 2276 3493
rect 2270 3488 2276 3489
rect 2446 3493 2452 3494
rect 2446 3489 2447 3493
rect 2451 3489 2452 3493
rect 2446 3488 2452 3489
rect 2630 3493 2636 3494
rect 2630 3489 2631 3493
rect 2635 3489 2636 3493
rect 2630 3488 2636 3489
rect 2272 3463 2274 3488
rect 2448 3463 2450 3488
rect 2632 3463 2634 3488
rect 2271 3462 2275 3463
rect 2271 3457 2275 3458
rect 2311 3462 2315 3463
rect 2311 3457 2315 3458
rect 2447 3462 2451 3463
rect 2447 3457 2451 3458
rect 2495 3462 2499 3463
rect 2495 3457 2499 3458
rect 2631 3462 2635 3463
rect 2631 3457 2635 3458
rect 2679 3462 2683 3463
rect 2679 3457 2683 3458
rect 2312 3436 2314 3457
rect 2496 3436 2498 3457
rect 2680 3436 2682 3457
rect 2310 3435 2316 3436
rect 2310 3431 2311 3435
rect 2315 3431 2316 3435
rect 2310 3430 2316 3431
rect 2494 3435 2500 3436
rect 2494 3431 2495 3435
rect 2499 3431 2500 3435
rect 2494 3430 2500 3431
rect 2678 3435 2684 3436
rect 2678 3431 2679 3435
rect 2683 3431 2684 3435
rect 2678 3430 2684 3431
rect 2780 3428 2782 3530
rect 2816 3513 2818 3537
rect 3000 3513 3002 3537
rect 3074 3535 3080 3536
rect 3074 3531 3075 3535
rect 3079 3531 3080 3535
rect 3074 3530 3080 3531
rect 2814 3512 2820 3513
rect 2814 3508 2815 3512
rect 2819 3508 2820 3512
rect 2814 3507 2820 3508
rect 2998 3512 3004 3513
rect 2998 3508 2999 3512
rect 3003 3508 3004 3512
rect 2998 3507 3004 3508
rect 3076 3504 3078 3530
rect 3176 3513 3178 3537
rect 3352 3513 3354 3537
rect 3398 3535 3404 3536
rect 3398 3531 3399 3535
rect 3403 3531 3404 3535
rect 3398 3530 3404 3531
rect 3426 3535 3432 3536
rect 3426 3531 3427 3535
rect 3431 3531 3432 3535
rect 3426 3530 3432 3531
rect 3174 3512 3180 3513
rect 3174 3508 3175 3512
rect 3179 3508 3180 3512
rect 3174 3507 3180 3508
rect 3350 3512 3356 3513
rect 3350 3508 3351 3512
rect 3355 3508 3356 3512
rect 3350 3507 3356 3508
rect 3074 3503 3080 3504
rect 3074 3499 3075 3503
rect 3079 3499 3080 3503
rect 3074 3498 3080 3499
rect 3250 3503 3256 3504
rect 3250 3499 3251 3503
rect 3255 3499 3256 3503
rect 3250 3498 3256 3499
rect 2814 3493 2820 3494
rect 2814 3489 2815 3493
rect 2819 3489 2820 3493
rect 2814 3488 2820 3489
rect 2998 3493 3004 3494
rect 2998 3489 2999 3493
rect 3003 3489 3004 3493
rect 2998 3488 3004 3489
rect 3174 3493 3180 3494
rect 3174 3489 3175 3493
rect 3179 3489 3180 3493
rect 3174 3488 3180 3489
rect 2816 3463 2818 3488
rect 3000 3463 3002 3488
rect 3176 3463 3178 3488
rect 2815 3462 2819 3463
rect 2815 3457 2819 3458
rect 2863 3462 2867 3463
rect 2863 3457 2867 3458
rect 2999 3462 3003 3463
rect 2999 3457 3003 3458
rect 3047 3462 3051 3463
rect 3047 3457 3051 3458
rect 3175 3462 3179 3463
rect 3175 3457 3179 3458
rect 3223 3462 3227 3463
rect 3223 3457 3227 3458
rect 2864 3436 2866 3457
rect 3048 3436 3050 3457
rect 3224 3436 3226 3457
rect 2862 3435 2868 3436
rect 2862 3431 2863 3435
rect 2867 3431 2868 3435
rect 2862 3430 2868 3431
rect 3046 3435 3052 3436
rect 3046 3431 3047 3435
rect 3051 3431 3052 3435
rect 3046 3430 3052 3431
rect 3222 3435 3228 3436
rect 3222 3431 3223 3435
rect 3227 3431 3228 3435
rect 3222 3430 3228 3431
rect 2778 3427 2784 3428
rect 2202 3423 2208 3424
rect 2202 3419 2203 3423
rect 2207 3419 2208 3423
rect 2202 3418 2208 3419
rect 2386 3423 2392 3424
rect 2386 3419 2387 3423
rect 2391 3419 2392 3423
rect 2386 3418 2392 3419
rect 2570 3423 2576 3424
rect 2570 3419 2571 3423
rect 2575 3419 2576 3423
rect 2778 3423 2779 3427
rect 2783 3423 2784 3427
rect 3174 3427 3180 3428
rect 2778 3422 2784 3423
rect 2946 3423 2952 3424
rect 2570 3418 2576 3419
rect 2946 3419 2947 3423
rect 2951 3419 2952 3423
rect 3174 3423 3175 3427
rect 3179 3423 3180 3427
rect 3174 3422 3180 3423
rect 2946 3418 2952 3419
rect 2178 3395 2184 3396
rect 2178 3391 2179 3395
rect 2183 3391 2184 3395
rect 2178 3390 2184 3391
rect 2047 3370 2051 3371
rect 2047 3365 2051 3366
rect 2071 3370 2075 3371
rect 2071 3365 2075 3366
rect 2127 3370 2131 3371
rect 2127 3365 2131 3366
rect 2006 3356 2012 3357
rect 2006 3352 2007 3356
rect 2011 3352 2012 3356
rect 2006 3351 2012 3352
rect 1946 3347 1952 3348
rect 1618 3343 1624 3344
rect 1618 3339 1619 3343
rect 1623 3339 1624 3343
rect 1618 3338 1624 3339
rect 1778 3343 1784 3344
rect 1778 3339 1779 3343
rect 1783 3339 1784 3343
rect 1946 3343 1947 3347
rect 1951 3343 1952 3347
rect 1946 3342 1952 3343
rect 1778 3338 1784 3339
rect 2006 3339 2012 3340
rect 1542 3336 1548 3337
rect 1542 3332 1543 3336
rect 1547 3332 1548 3336
rect 1542 3331 1548 3332
rect 1426 3315 1432 3316
rect 1426 3311 1427 3315
rect 1431 3311 1432 3315
rect 1426 3310 1432 3311
rect 1544 3307 1546 3331
rect 1620 3316 1622 3338
rect 1702 3336 1708 3337
rect 1702 3332 1703 3336
rect 1707 3332 1708 3336
rect 1702 3331 1708 3332
rect 1618 3315 1624 3316
rect 1594 3311 1600 3312
rect 1594 3307 1595 3311
rect 1599 3307 1600 3311
rect 1618 3311 1619 3315
rect 1623 3311 1624 3315
rect 1618 3310 1624 3311
rect 1704 3307 1706 3331
rect 1780 3316 1782 3338
rect 1870 3336 1876 3337
rect 1870 3332 1871 3336
rect 1875 3332 1876 3336
rect 2006 3335 2007 3339
rect 2011 3335 2012 3339
rect 2048 3338 2050 3365
rect 2072 3341 2074 3365
rect 2204 3364 2206 3418
rect 2310 3416 2316 3417
rect 2310 3412 2311 3416
rect 2315 3412 2316 3416
rect 2310 3411 2316 3412
rect 2312 3371 2314 3411
rect 2388 3396 2390 3418
rect 2494 3416 2500 3417
rect 2494 3412 2495 3416
rect 2499 3412 2500 3416
rect 2494 3411 2500 3412
rect 2386 3395 2392 3396
rect 2386 3391 2387 3395
rect 2391 3391 2392 3395
rect 2386 3390 2392 3391
rect 2496 3371 2498 3411
rect 2572 3396 2574 3418
rect 2678 3416 2684 3417
rect 2678 3412 2679 3416
rect 2683 3412 2684 3416
rect 2678 3411 2684 3412
rect 2862 3416 2868 3417
rect 2862 3412 2863 3416
rect 2867 3412 2868 3416
rect 2862 3411 2868 3412
rect 2570 3395 2576 3396
rect 2570 3391 2571 3395
rect 2575 3391 2576 3395
rect 2570 3390 2576 3391
rect 2680 3371 2682 3411
rect 2864 3371 2866 3411
rect 2215 3370 2219 3371
rect 2215 3365 2219 3366
rect 2311 3370 2315 3371
rect 2311 3365 2315 3366
rect 2359 3370 2363 3371
rect 2359 3365 2363 3366
rect 2495 3370 2499 3371
rect 2495 3365 2499 3366
rect 2511 3370 2515 3371
rect 2511 3365 2515 3366
rect 2655 3370 2659 3371
rect 2655 3365 2659 3366
rect 2679 3370 2683 3371
rect 2679 3365 2683 3366
rect 2799 3370 2803 3371
rect 2799 3365 2803 3366
rect 2863 3370 2867 3371
rect 2863 3365 2867 3366
rect 2935 3370 2939 3371
rect 2935 3365 2939 3366
rect 2154 3363 2160 3364
rect 2154 3359 2155 3363
rect 2159 3359 2160 3363
rect 2154 3358 2160 3359
rect 2202 3363 2208 3364
rect 2202 3359 2203 3363
rect 2207 3359 2208 3363
rect 2202 3358 2208 3359
rect 2070 3340 2076 3341
rect 2006 3334 2012 3335
rect 2046 3337 2052 3338
rect 1870 3331 1876 3332
rect 1778 3315 1784 3316
rect 1778 3311 1779 3315
rect 1783 3311 1784 3315
rect 1778 3310 1784 3311
rect 1872 3307 1874 3331
rect 2008 3307 2010 3334
rect 2046 3333 2047 3337
rect 2051 3333 2052 3337
rect 2070 3336 2071 3340
rect 2075 3336 2076 3340
rect 2070 3335 2076 3336
rect 2046 3332 2052 3333
rect 2156 3332 2158 3358
rect 2216 3341 2218 3365
rect 2360 3341 2362 3365
rect 2442 3363 2448 3364
rect 2442 3359 2443 3363
rect 2447 3359 2448 3363
rect 2442 3358 2448 3359
rect 2214 3340 2220 3341
rect 2214 3336 2215 3340
rect 2219 3336 2220 3340
rect 2214 3335 2220 3336
rect 2358 3340 2364 3341
rect 2358 3336 2359 3340
rect 2363 3336 2364 3340
rect 2358 3335 2364 3336
rect 2444 3332 2446 3358
rect 2512 3341 2514 3365
rect 2594 3363 2600 3364
rect 2594 3359 2595 3363
rect 2599 3359 2600 3363
rect 2594 3358 2600 3359
rect 2510 3340 2516 3341
rect 2510 3336 2511 3340
rect 2515 3336 2516 3340
rect 2510 3335 2516 3336
rect 2596 3332 2598 3358
rect 2656 3341 2658 3365
rect 2774 3363 2780 3364
rect 2774 3359 2775 3363
rect 2779 3359 2780 3363
rect 2774 3358 2780 3359
rect 2654 3340 2660 3341
rect 2654 3336 2655 3340
rect 2659 3336 2660 3340
rect 2654 3335 2660 3336
rect 2776 3332 2778 3358
rect 2800 3341 2802 3365
rect 2870 3363 2876 3364
rect 2870 3359 2871 3363
rect 2875 3359 2876 3363
rect 2870 3358 2876 3359
rect 2798 3340 2804 3341
rect 2798 3336 2799 3340
rect 2803 3336 2804 3340
rect 2798 3335 2804 3336
rect 2146 3331 2152 3332
rect 2146 3327 2147 3331
rect 2151 3327 2152 3331
rect 2146 3326 2152 3327
rect 2154 3331 2160 3332
rect 2154 3327 2155 3331
rect 2159 3327 2160 3331
rect 2154 3326 2160 3327
rect 2442 3331 2448 3332
rect 2442 3327 2443 3331
rect 2447 3327 2448 3331
rect 2442 3326 2448 3327
rect 2594 3331 2600 3332
rect 2594 3327 2595 3331
rect 2599 3327 2600 3331
rect 2594 3326 2600 3327
rect 2774 3331 2780 3332
rect 2774 3327 2775 3331
rect 2779 3327 2780 3331
rect 2774 3326 2780 3327
rect 2070 3321 2076 3322
rect 2046 3320 2052 3321
rect 2046 3316 2047 3320
rect 2051 3316 2052 3320
rect 2070 3317 2071 3321
rect 2075 3317 2076 3321
rect 2070 3316 2076 3317
rect 2046 3315 2052 3316
rect 1215 3306 1219 3307
rect 1215 3301 1219 3302
rect 1295 3306 1299 3307
rect 1295 3301 1299 3302
rect 1383 3306 1387 3307
rect 1383 3301 1387 3302
rect 1519 3306 1523 3307
rect 1519 3301 1523 3302
rect 1543 3306 1547 3307
rect 1594 3306 1600 3307
rect 1703 3306 1707 3307
rect 1543 3301 1547 3302
rect 1122 3299 1128 3300
rect 1122 3295 1123 3299
rect 1127 3295 1128 3299
rect 1122 3294 1128 3295
rect 1154 3299 1160 3300
rect 1154 3295 1155 3299
rect 1159 3295 1160 3299
rect 1154 3294 1160 3295
rect 870 3276 876 3277
rect 870 3272 871 3276
rect 875 3272 876 3276
rect 870 3271 876 3272
rect 1078 3276 1084 3277
rect 1078 3272 1079 3276
rect 1083 3272 1084 3276
rect 1078 3271 1084 3272
rect 1156 3268 1158 3294
rect 1296 3277 1298 3301
rect 1520 3277 1522 3301
rect 1294 3276 1300 3277
rect 1294 3272 1295 3276
rect 1299 3272 1300 3276
rect 1294 3271 1300 3272
rect 1518 3276 1524 3277
rect 1518 3272 1519 3276
rect 1523 3272 1524 3276
rect 1518 3271 1524 3272
rect 1596 3268 1598 3306
rect 1703 3301 1707 3302
rect 1743 3306 1747 3307
rect 1743 3301 1747 3302
rect 1871 3306 1875 3307
rect 1871 3301 1875 3302
rect 2007 3306 2011 3307
rect 2007 3301 2011 3302
rect 1602 3299 1608 3300
rect 1602 3295 1603 3299
rect 1607 3295 1608 3299
rect 1602 3294 1608 3295
rect 1604 3268 1606 3294
rect 1744 3277 1746 3301
rect 1770 3299 1776 3300
rect 1770 3295 1771 3299
rect 1775 3295 1776 3299
rect 1770 3294 1776 3295
rect 1742 3276 1748 3277
rect 1742 3272 1743 3276
rect 1747 3272 1748 3276
rect 1742 3271 1748 3272
rect 738 3267 744 3268
rect 738 3263 739 3267
rect 743 3263 744 3267
rect 738 3262 744 3263
rect 798 3267 804 3268
rect 798 3263 799 3267
rect 803 3263 804 3267
rect 798 3262 804 3263
rect 1154 3267 1160 3268
rect 1154 3263 1155 3267
rect 1159 3263 1160 3267
rect 1154 3262 1160 3263
rect 1370 3267 1376 3268
rect 1370 3263 1371 3267
rect 1375 3263 1376 3267
rect 1370 3262 1376 3263
rect 1594 3267 1600 3268
rect 1594 3263 1595 3267
rect 1599 3263 1600 3267
rect 1594 3262 1600 3263
rect 1602 3267 1608 3268
rect 1602 3263 1603 3267
rect 1607 3263 1608 3267
rect 1602 3262 1608 3263
rect 662 3257 668 3258
rect 662 3253 663 3257
rect 667 3253 668 3257
rect 662 3252 668 3253
rect 870 3257 876 3258
rect 870 3253 871 3257
rect 875 3253 876 3257
rect 870 3252 876 3253
rect 1078 3257 1084 3258
rect 1078 3253 1079 3257
rect 1083 3253 1084 3257
rect 1078 3252 1084 3253
rect 1294 3257 1300 3258
rect 1294 3253 1295 3257
rect 1299 3253 1300 3257
rect 1294 3252 1300 3253
rect 664 3231 666 3252
rect 872 3231 874 3252
rect 1080 3231 1082 3252
rect 1296 3231 1298 3252
rect 615 3230 619 3231
rect 615 3225 619 3226
rect 663 3230 667 3231
rect 663 3225 667 3226
rect 791 3230 795 3231
rect 791 3225 795 3226
rect 871 3230 875 3231
rect 871 3225 875 3226
rect 967 3230 971 3231
rect 967 3225 971 3226
rect 1079 3230 1083 3231
rect 1079 3225 1083 3226
rect 1143 3230 1147 3231
rect 1143 3225 1147 3226
rect 1295 3230 1299 3231
rect 1295 3225 1299 3226
rect 1327 3230 1331 3231
rect 1327 3225 1331 3226
rect 616 3204 618 3225
rect 792 3204 794 3225
rect 968 3204 970 3225
rect 1144 3204 1146 3225
rect 1328 3204 1330 3225
rect 614 3203 620 3204
rect 614 3199 615 3203
rect 619 3199 620 3203
rect 614 3198 620 3199
rect 790 3203 796 3204
rect 790 3199 791 3203
rect 795 3199 796 3203
rect 790 3198 796 3199
rect 966 3203 972 3204
rect 966 3199 967 3203
rect 971 3199 972 3203
rect 966 3198 972 3199
rect 1142 3203 1148 3204
rect 1142 3199 1143 3203
rect 1147 3199 1148 3203
rect 1142 3198 1148 3199
rect 1326 3203 1332 3204
rect 1326 3199 1327 3203
rect 1331 3199 1332 3203
rect 1326 3198 1332 3199
rect 522 3195 528 3196
rect 258 3191 264 3192
rect 110 3187 116 3188
rect 110 3183 111 3187
rect 115 3183 116 3187
rect 258 3187 259 3191
rect 263 3187 264 3191
rect 258 3186 264 3187
rect 362 3191 368 3192
rect 362 3187 363 3191
rect 367 3187 368 3191
rect 522 3191 523 3195
rect 527 3191 528 3195
rect 522 3190 528 3191
rect 558 3195 564 3196
rect 558 3191 559 3195
rect 563 3191 564 3195
rect 558 3190 564 3191
rect 750 3195 756 3196
rect 750 3191 751 3195
rect 755 3191 756 3195
rect 1090 3195 1096 3196
rect 750 3190 756 3191
rect 1042 3191 1048 3192
rect 362 3186 368 3187
rect 110 3182 116 3183
rect 134 3184 140 3185
rect 112 3151 114 3182
rect 134 3180 135 3184
rect 139 3180 140 3184
rect 134 3179 140 3180
rect 136 3151 138 3179
rect 260 3160 262 3186
rect 286 3184 292 3185
rect 286 3180 287 3184
rect 291 3180 292 3184
rect 286 3179 292 3180
rect 258 3159 264 3160
rect 258 3155 259 3159
rect 263 3155 264 3159
rect 258 3154 264 3155
rect 288 3151 290 3179
rect 364 3164 366 3186
rect 446 3184 452 3185
rect 446 3180 447 3184
rect 451 3180 452 3184
rect 446 3179 452 3180
rect 362 3163 368 3164
rect 362 3159 363 3163
rect 367 3159 368 3163
rect 362 3158 368 3159
rect 448 3151 450 3179
rect 560 3172 562 3190
rect 614 3184 620 3185
rect 614 3180 615 3184
rect 619 3180 620 3184
rect 614 3179 620 3180
rect 558 3171 564 3172
rect 558 3167 559 3171
rect 563 3167 564 3171
rect 558 3166 564 3167
rect 616 3151 618 3179
rect 752 3164 754 3190
rect 1042 3187 1043 3191
rect 1047 3187 1048 3191
rect 1090 3191 1091 3195
rect 1095 3191 1096 3195
rect 1090 3190 1096 3191
rect 1042 3186 1048 3187
rect 790 3184 796 3185
rect 790 3180 791 3184
rect 795 3180 796 3184
rect 790 3179 796 3180
rect 966 3184 972 3185
rect 966 3180 967 3184
rect 971 3180 972 3184
rect 966 3179 972 3180
rect 750 3163 756 3164
rect 750 3159 751 3163
rect 755 3159 756 3163
rect 750 3158 756 3159
rect 792 3151 794 3179
rect 968 3151 970 3179
rect 111 3150 115 3151
rect 111 3145 115 3146
rect 135 3150 139 3151
rect 135 3145 139 3146
rect 287 3150 291 3151
rect 287 3145 291 3146
rect 311 3150 315 3151
rect 311 3145 315 3146
rect 439 3150 443 3151
rect 439 3145 443 3146
rect 447 3150 451 3151
rect 447 3145 451 3146
rect 583 3150 587 3151
rect 583 3145 587 3146
rect 615 3150 619 3151
rect 615 3145 619 3146
rect 743 3150 747 3151
rect 743 3145 747 3146
rect 791 3150 795 3151
rect 791 3145 795 3146
rect 903 3150 907 3151
rect 903 3145 907 3146
rect 967 3150 971 3151
rect 967 3145 971 3146
rect 112 3118 114 3145
rect 312 3121 314 3145
rect 366 3143 372 3144
rect 366 3139 367 3143
rect 371 3139 372 3143
rect 366 3138 372 3139
rect 386 3143 392 3144
rect 386 3139 387 3143
rect 391 3139 392 3143
rect 386 3138 392 3139
rect 310 3120 316 3121
rect 110 3117 116 3118
rect 110 3113 111 3117
rect 115 3113 116 3117
rect 310 3116 311 3120
rect 315 3116 316 3120
rect 310 3115 316 3116
rect 110 3112 116 3113
rect 310 3101 316 3102
rect 110 3100 116 3101
rect 110 3096 111 3100
rect 115 3096 116 3100
rect 310 3097 311 3101
rect 315 3097 316 3101
rect 310 3096 316 3097
rect 110 3095 116 3096
rect 112 3067 114 3095
rect 312 3067 314 3096
rect 111 3066 115 3067
rect 111 3061 115 3062
rect 311 3066 315 3067
rect 311 3061 315 3062
rect 112 3041 114 3061
rect 110 3040 116 3041
rect 110 3036 111 3040
rect 115 3036 116 3040
rect 110 3035 116 3036
rect 368 3032 370 3138
rect 388 3112 390 3138
rect 440 3121 442 3145
rect 514 3143 520 3144
rect 514 3139 515 3143
rect 519 3139 520 3143
rect 514 3138 520 3139
rect 438 3120 444 3121
rect 438 3116 439 3120
rect 443 3116 444 3120
rect 438 3115 444 3116
rect 516 3112 518 3138
rect 584 3121 586 3145
rect 658 3143 664 3144
rect 658 3139 659 3143
rect 663 3139 664 3143
rect 658 3138 664 3139
rect 582 3120 588 3121
rect 582 3116 583 3120
rect 587 3116 588 3120
rect 582 3115 588 3116
rect 660 3112 662 3138
rect 744 3121 746 3145
rect 818 3143 824 3144
rect 818 3139 819 3143
rect 823 3139 824 3143
rect 818 3138 824 3139
rect 742 3120 748 3121
rect 742 3116 743 3120
rect 747 3116 748 3120
rect 742 3115 748 3116
rect 820 3112 822 3138
rect 904 3121 906 3145
rect 1044 3144 1046 3186
rect 1092 3164 1094 3190
rect 1142 3184 1148 3185
rect 1142 3180 1143 3184
rect 1147 3180 1148 3184
rect 1142 3179 1148 3180
rect 1326 3184 1332 3185
rect 1326 3180 1327 3184
rect 1331 3180 1332 3184
rect 1326 3179 1332 3180
rect 1090 3163 1096 3164
rect 1090 3159 1091 3163
rect 1095 3159 1096 3163
rect 1090 3158 1096 3159
rect 1144 3151 1146 3179
rect 1328 3151 1330 3179
rect 1372 3164 1374 3262
rect 1518 3257 1524 3258
rect 1518 3253 1519 3257
rect 1523 3253 1524 3257
rect 1518 3252 1524 3253
rect 1742 3257 1748 3258
rect 1742 3253 1743 3257
rect 1747 3253 1748 3257
rect 1742 3252 1748 3253
rect 1520 3231 1522 3252
rect 1744 3231 1746 3252
rect 1511 3230 1515 3231
rect 1511 3225 1515 3226
rect 1519 3230 1523 3231
rect 1519 3225 1523 3226
rect 1695 3230 1699 3231
rect 1695 3225 1699 3226
rect 1743 3230 1747 3231
rect 1743 3225 1747 3226
rect 1512 3204 1514 3225
rect 1696 3204 1698 3225
rect 1510 3203 1516 3204
rect 1510 3199 1511 3203
rect 1515 3199 1516 3203
rect 1510 3198 1516 3199
rect 1694 3203 1700 3204
rect 1694 3199 1695 3203
rect 1699 3199 1700 3203
rect 1694 3198 1700 3199
rect 1772 3196 1774 3294
rect 2008 3274 2010 3301
rect 2048 3287 2050 3315
rect 2072 3287 2074 3316
rect 2047 3286 2051 3287
rect 2047 3281 2051 3282
rect 2071 3286 2075 3287
rect 2071 3281 2075 3282
rect 2111 3286 2115 3287
rect 2111 3281 2115 3282
rect 2006 3273 2012 3274
rect 2006 3269 2007 3273
rect 2011 3269 2012 3273
rect 2006 3268 2012 3269
rect 2048 3261 2050 3281
rect 2046 3260 2052 3261
rect 2112 3260 2114 3281
rect 2006 3256 2012 3257
rect 2006 3252 2007 3256
rect 2011 3252 2012 3256
rect 2046 3256 2047 3260
rect 2051 3256 2052 3260
rect 2046 3255 2052 3256
rect 2110 3259 2116 3260
rect 2110 3255 2111 3259
rect 2115 3255 2116 3259
rect 2110 3254 2116 3255
rect 2006 3251 2012 3252
rect 2008 3231 2010 3251
rect 2046 3243 2052 3244
rect 2046 3239 2047 3243
rect 2051 3239 2052 3243
rect 2046 3238 2052 3239
rect 2110 3240 2116 3241
rect 2007 3230 2011 3231
rect 2007 3225 2011 3226
rect 2008 3205 2010 3225
rect 2048 3211 2050 3238
rect 2110 3236 2111 3240
rect 2115 3236 2116 3240
rect 2110 3235 2116 3236
rect 2112 3211 2114 3235
rect 2148 3220 2150 3326
rect 2214 3321 2220 3322
rect 2214 3317 2215 3321
rect 2219 3317 2220 3321
rect 2214 3316 2220 3317
rect 2358 3321 2364 3322
rect 2358 3317 2359 3321
rect 2363 3317 2364 3321
rect 2358 3316 2364 3317
rect 2510 3321 2516 3322
rect 2510 3317 2511 3321
rect 2515 3317 2516 3321
rect 2510 3316 2516 3317
rect 2654 3321 2660 3322
rect 2654 3317 2655 3321
rect 2659 3317 2660 3321
rect 2654 3316 2660 3317
rect 2798 3321 2804 3322
rect 2798 3317 2799 3321
rect 2803 3317 2804 3321
rect 2798 3316 2804 3317
rect 2216 3287 2218 3316
rect 2360 3287 2362 3316
rect 2512 3287 2514 3316
rect 2656 3287 2658 3316
rect 2800 3287 2802 3316
rect 2215 3286 2219 3287
rect 2215 3281 2219 3282
rect 2247 3286 2251 3287
rect 2247 3281 2251 3282
rect 2359 3286 2363 3287
rect 2359 3281 2363 3282
rect 2399 3286 2403 3287
rect 2399 3281 2403 3282
rect 2511 3286 2515 3287
rect 2511 3281 2515 3282
rect 2575 3286 2579 3287
rect 2575 3281 2579 3282
rect 2655 3286 2659 3287
rect 2655 3281 2659 3282
rect 2783 3286 2787 3287
rect 2783 3281 2787 3282
rect 2799 3286 2803 3287
rect 2799 3281 2803 3282
rect 2248 3260 2250 3281
rect 2400 3260 2402 3281
rect 2576 3260 2578 3281
rect 2784 3260 2786 3281
rect 2246 3259 2252 3260
rect 2246 3255 2247 3259
rect 2251 3255 2252 3259
rect 2246 3254 2252 3255
rect 2398 3259 2404 3260
rect 2398 3255 2399 3259
rect 2403 3255 2404 3259
rect 2398 3254 2404 3255
rect 2574 3259 2580 3260
rect 2574 3255 2575 3259
rect 2579 3255 2580 3259
rect 2574 3254 2580 3255
rect 2782 3259 2788 3260
rect 2782 3255 2783 3259
rect 2787 3255 2788 3259
rect 2872 3256 2874 3358
rect 2936 3341 2938 3365
rect 2948 3364 2950 3418
rect 3046 3416 3052 3417
rect 3046 3412 3047 3416
rect 3051 3412 3052 3416
rect 3046 3411 3052 3412
rect 3048 3371 3050 3411
rect 3176 3396 3178 3422
rect 3222 3416 3228 3417
rect 3222 3412 3223 3416
rect 3227 3412 3228 3416
rect 3222 3411 3228 3412
rect 3174 3395 3180 3396
rect 3174 3391 3175 3395
rect 3179 3391 3180 3395
rect 3174 3390 3180 3391
rect 3224 3371 3226 3411
rect 3252 3396 3254 3498
rect 3350 3493 3356 3494
rect 3350 3489 3351 3493
rect 3355 3489 3356 3493
rect 3350 3488 3356 3489
rect 3352 3463 3354 3488
rect 3351 3462 3355 3463
rect 3351 3457 3355 3458
rect 3400 3428 3402 3530
rect 3428 3504 3430 3530
rect 3520 3513 3522 3537
rect 3518 3512 3524 3513
rect 3518 3508 3519 3512
rect 3523 3508 3524 3512
rect 3518 3507 3524 3508
rect 3596 3504 3598 3542
rect 3623 3537 3627 3538
rect 3687 3542 3691 3543
rect 3687 3537 3691 3538
rect 3688 3513 3690 3537
rect 3770 3535 3776 3536
rect 3770 3531 3771 3535
rect 3775 3531 3776 3535
rect 3770 3530 3776 3531
rect 3686 3512 3692 3513
rect 3686 3508 3687 3512
rect 3691 3508 3692 3512
rect 3686 3507 3692 3508
rect 3772 3504 3774 3530
rect 3426 3503 3432 3504
rect 3426 3499 3427 3503
rect 3431 3499 3432 3503
rect 3426 3498 3432 3499
rect 3594 3503 3600 3504
rect 3594 3499 3595 3503
rect 3599 3499 3600 3503
rect 3594 3498 3600 3499
rect 3770 3503 3776 3504
rect 3770 3499 3771 3503
rect 3775 3499 3776 3503
rect 3770 3498 3776 3499
rect 3518 3493 3524 3494
rect 3518 3489 3519 3493
rect 3523 3489 3524 3493
rect 3518 3488 3524 3489
rect 3686 3493 3692 3494
rect 3686 3489 3687 3493
rect 3691 3489 3692 3493
rect 3686 3488 3692 3489
rect 3520 3463 3522 3488
rect 3688 3463 3690 3488
rect 3407 3462 3411 3463
rect 3407 3457 3411 3458
rect 3519 3462 3523 3463
rect 3519 3457 3523 3458
rect 3591 3462 3595 3463
rect 3591 3457 3595 3458
rect 3687 3462 3691 3463
rect 3687 3457 3691 3458
rect 3775 3462 3779 3463
rect 3775 3457 3779 3458
rect 3408 3436 3410 3457
rect 3592 3436 3594 3457
rect 3776 3436 3778 3457
rect 3406 3435 3412 3436
rect 3406 3431 3407 3435
rect 3411 3431 3412 3435
rect 3406 3430 3412 3431
rect 3590 3435 3596 3436
rect 3590 3431 3591 3435
rect 3595 3431 3596 3435
rect 3590 3430 3596 3431
rect 3774 3435 3780 3436
rect 3774 3431 3775 3435
rect 3779 3431 3780 3435
rect 3774 3430 3780 3431
rect 3398 3427 3404 3428
rect 3398 3423 3399 3427
rect 3403 3423 3404 3427
rect 3398 3422 3404 3423
rect 3546 3427 3552 3428
rect 3546 3423 3547 3427
rect 3551 3423 3552 3427
rect 3546 3422 3552 3423
rect 3406 3416 3412 3417
rect 3406 3412 3407 3416
rect 3411 3412 3412 3416
rect 3406 3411 3412 3412
rect 3250 3395 3256 3396
rect 3250 3391 3251 3395
rect 3255 3391 3256 3395
rect 3250 3390 3256 3391
rect 3408 3371 3410 3411
rect 3548 3396 3550 3422
rect 3590 3416 3596 3417
rect 3590 3412 3591 3416
rect 3595 3412 3596 3416
rect 3590 3411 3596 3412
rect 3774 3416 3780 3417
rect 3774 3412 3775 3416
rect 3779 3412 3780 3416
rect 3774 3411 3780 3412
rect 3546 3395 3552 3396
rect 3546 3391 3547 3395
rect 3551 3391 3552 3395
rect 3546 3390 3552 3391
rect 3592 3371 3594 3411
rect 3658 3391 3664 3392
rect 3658 3387 3659 3391
rect 3663 3387 3664 3391
rect 3658 3386 3664 3387
rect 3047 3370 3051 3371
rect 3047 3365 3051 3366
rect 3079 3370 3083 3371
rect 3079 3365 3083 3366
rect 3223 3370 3227 3371
rect 3223 3365 3227 3366
rect 3375 3370 3379 3371
rect 3375 3365 3379 3366
rect 3407 3370 3411 3371
rect 3407 3365 3411 3366
rect 3535 3370 3539 3371
rect 3535 3365 3539 3366
rect 3591 3370 3595 3371
rect 3591 3365 3595 3366
rect 2946 3363 2952 3364
rect 2946 3359 2947 3363
rect 2951 3359 2952 3363
rect 2946 3358 2952 3359
rect 3010 3363 3016 3364
rect 3010 3359 3011 3363
rect 3015 3359 3016 3363
rect 3010 3358 3016 3359
rect 2934 3340 2940 3341
rect 2934 3336 2935 3340
rect 2939 3336 2940 3340
rect 2934 3335 2940 3336
rect 3012 3332 3014 3358
rect 3080 3341 3082 3365
rect 3154 3363 3160 3364
rect 3154 3359 3155 3363
rect 3159 3359 3160 3363
rect 3154 3358 3160 3359
rect 3078 3340 3084 3341
rect 3078 3336 3079 3340
rect 3083 3336 3084 3340
rect 3078 3335 3084 3336
rect 3156 3332 3158 3358
rect 3224 3341 3226 3365
rect 3376 3341 3378 3365
rect 3498 3363 3504 3364
rect 3498 3359 3499 3363
rect 3503 3359 3504 3363
rect 3498 3358 3504 3359
rect 3506 3363 3512 3364
rect 3506 3359 3507 3363
rect 3511 3359 3512 3363
rect 3506 3358 3512 3359
rect 3222 3340 3228 3341
rect 3222 3336 3223 3340
rect 3227 3336 3228 3340
rect 3222 3335 3228 3336
rect 3374 3340 3380 3341
rect 3374 3336 3375 3340
rect 3379 3336 3380 3340
rect 3374 3335 3380 3336
rect 3010 3331 3016 3332
rect 3010 3327 3011 3331
rect 3015 3327 3016 3331
rect 3010 3326 3016 3327
rect 3154 3331 3160 3332
rect 3154 3327 3155 3331
rect 3159 3327 3160 3331
rect 3154 3326 3160 3327
rect 3298 3331 3304 3332
rect 3298 3327 3299 3331
rect 3303 3327 3304 3331
rect 3298 3326 3304 3327
rect 2934 3321 2940 3322
rect 2934 3317 2935 3321
rect 2939 3317 2940 3321
rect 2934 3316 2940 3317
rect 3078 3321 3084 3322
rect 3078 3317 3079 3321
rect 3083 3317 3084 3321
rect 3078 3316 3084 3317
rect 3222 3321 3228 3322
rect 3222 3317 3223 3321
rect 3227 3317 3228 3321
rect 3222 3316 3228 3317
rect 2936 3287 2938 3316
rect 3080 3287 3082 3316
rect 3224 3287 3226 3316
rect 3300 3309 3302 3326
rect 3374 3321 3380 3322
rect 3374 3317 3375 3321
rect 3379 3317 3380 3321
rect 3374 3316 3380 3317
rect 3299 3308 3303 3309
rect 3299 3303 3303 3304
rect 3376 3287 3378 3316
rect 2935 3286 2939 3287
rect 2935 3281 2939 3282
rect 3015 3286 3019 3287
rect 3015 3281 3019 3282
rect 3079 3286 3083 3287
rect 3079 3281 3083 3282
rect 3223 3286 3227 3287
rect 3223 3281 3227 3282
rect 3263 3286 3267 3287
rect 3263 3281 3267 3282
rect 3375 3286 3379 3287
rect 3375 3281 3379 3282
rect 3016 3260 3018 3281
rect 3264 3260 3266 3281
rect 3014 3259 3020 3260
rect 2782 3254 2788 3255
rect 2870 3255 2876 3256
rect 2870 3251 2871 3255
rect 2875 3251 2876 3255
rect 3014 3255 3015 3259
rect 3019 3255 3020 3259
rect 3014 3254 3020 3255
rect 3262 3259 3268 3260
rect 3262 3255 3263 3259
rect 3267 3255 3268 3259
rect 3262 3254 3268 3255
rect 3500 3252 3502 3358
rect 3508 3332 3510 3358
rect 3536 3341 3538 3365
rect 3610 3363 3616 3364
rect 3610 3359 3611 3363
rect 3615 3359 3616 3363
rect 3610 3358 3616 3359
rect 3534 3340 3540 3341
rect 3534 3336 3535 3340
rect 3539 3336 3540 3340
rect 3534 3335 3540 3336
rect 3612 3332 3614 3358
rect 3660 3332 3662 3386
rect 3776 3371 3778 3411
rect 3828 3396 3830 3658
rect 3942 3652 3948 3653
rect 3942 3648 3943 3652
rect 3947 3648 3948 3652
rect 3942 3647 3948 3648
rect 3944 3619 3946 3647
rect 3943 3618 3947 3619
rect 3943 3613 3947 3614
rect 3944 3593 3946 3613
rect 3942 3592 3948 3593
rect 3942 3588 3943 3592
rect 3947 3588 3948 3592
rect 3942 3587 3948 3588
rect 3942 3575 3948 3576
rect 3942 3571 3943 3575
rect 3947 3571 3948 3575
rect 3942 3570 3948 3571
rect 3944 3543 3946 3570
rect 3839 3542 3843 3543
rect 3839 3537 3843 3538
rect 3943 3542 3947 3543
rect 3943 3537 3947 3538
rect 3840 3513 3842 3537
rect 3914 3535 3920 3536
rect 3914 3531 3915 3535
rect 3919 3531 3920 3535
rect 3914 3530 3920 3531
rect 3838 3512 3844 3513
rect 3838 3508 3839 3512
rect 3843 3508 3844 3512
rect 3838 3507 3844 3508
rect 3838 3493 3844 3494
rect 3838 3489 3839 3493
rect 3843 3489 3844 3493
rect 3838 3488 3844 3489
rect 3840 3463 3842 3488
rect 3839 3462 3843 3463
rect 3839 3457 3843 3458
rect 3850 3423 3856 3424
rect 3850 3419 3851 3423
rect 3855 3419 3856 3423
rect 3850 3418 3856 3419
rect 3826 3395 3832 3396
rect 3826 3391 3827 3395
rect 3831 3391 3832 3395
rect 3826 3390 3832 3391
rect 3695 3370 3699 3371
rect 3695 3365 3699 3366
rect 3775 3370 3779 3371
rect 3775 3365 3779 3366
rect 3839 3370 3843 3371
rect 3839 3365 3843 3366
rect 3696 3341 3698 3365
rect 3840 3341 3842 3365
rect 3694 3340 3700 3341
rect 3694 3336 3695 3340
rect 3699 3336 3700 3340
rect 3694 3335 3700 3336
rect 3838 3340 3844 3341
rect 3838 3336 3839 3340
rect 3843 3336 3844 3340
rect 3838 3335 3844 3336
rect 3506 3331 3512 3332
rect 3506 3327 3507 3331
rect 3511 3327 3512 3331
rect 3506 3326 3512 3327
rect 3610 3331 3616 3332
rect 3610 3327 3611 3331
rect 3615 3327 3616 3331
rect 3610 3326 3616 3327
rect 3658 3331 3664 3332
rect 3658 3327 3659 3331
rect 3663 3327 3664 3331
rect 3658 3326 3664 3327
rect 3534 3321 3540 3322
rect 3534 3317 3535 3321
rect 3539 3317 3540 3321
rect 3534 3316 3540 3317
rect 3694 3321 3700 3322
rect 3694 3317 3695 3321
rect 3699 3317 3700 3321
rect 3694 3316 3700 3317
rect 3838 3321 3844 3322
rect 3838 3317 3839 3321
rect 3843 3317 3844 3321
rect 3838 3316 3844 3317
rect 3507 3308 3511 3309
rect 3507 3303 3511 3304
rect 2870 3250 2876 3251
rect 3498 3251 3504 3252
rect 2186 3247 2192 3248
rect 2186 3243 2187 3247
rect 2191 3243 2192 3247
rect 2186 3242 2192 3243
rect 2474 3247 2480 3248
rect 2474 3243 2475 3247
rect 2479 3243 2480 3247
rect 2474 3242 2480 3243
rect 2650 3247 2656 3248
rect 2650 3243 2651 3247
rect 2655 3243 2656 3247
rect 2650 3242 2656 3243
rect 2858 3247 2864 3248
rect 2858 3243 2859 3247
rect 2863 3243 2864 3247
rect 2858 3242 2864 3243
rect 3338 3247 3344 3248
rect 3338 3243 3339 3247
rect 3343 3243 3344 3247
rect 3498 3247 3499 3251
rect 3503 3247 3504 3251
rect 3498 3246 3504 3247
rect 3338 3242 3344 3243
rect 2146 3219 2152 3220
rect 2146 3215 2147 3219
rect 2151 3215 2152 3219
rect 2146 3214 2152 3215
rect 2047 3210 2051 3211
rect 2047 3205 2051 3206
rect 2071 3210 2075 3211
rect 2071 3205 2075 3206
rect 2111 3210 2115 3211
rect 2111 3205 2115 3206
rect 2167 3210 2171 3211
rect 2167 3205 2171 3206
rect 2006 3204 2012 3205
rect 2006 3200 2007 3204
rect 2011 3200 2012 3204
rect 2006 3199 2012 3200
rect 1770 3195 1776 3196
rect 1586 3191 1592 3192
rect 1586 3187 1587 3191
rect 1591 3187 1592 3191
rect 1770 3191 1771 3195
rect 1775 3191 1776 3195
rect 1770 3190 1776 3191
rect 1586 3186 1592 3187
rect 2006 3187 2012 3188
rect 1510 3184 1516 3185
rect 1510 3180 1511 3184
rect 1515 3180 1516 3184
rect 1510 3179 1516 3180
rect 1370 3163 1376 3164
rect 1370 3159 1371 3163
rect 1375 3159 1376 3163
rect 1370 3158 1376 3159
rect 1466 3159 1472 3160
rect 1466 3155 1467 3159
rect 1471 3155 1472 3159
rect 1466 3154 1472 3155
rect 1063 3150 1067 3151
rect 1063 3145 1067 3146
rect 1143 3150 1147 3151
rect 1143 3145 1147 3146
rect 1223 3150 1227 3151
rect 1223 3145 1227 3146
rect 1327 3150 1331 3151
rect 1327 3145 1331 3146
rect 1391 3150 1395 3151
rect 1391 3145 1395 3146
rect 1042 3143 1048 3144
rect 1042 3139 1043 3143
rect 1047 3139 1048 3143
rect 1042 3138 1048 3139
rect 1064 3121 1066 3145
rect 1224 3121 1226 3145
rect 1392 3121 1394 3145
rect 902 3120 908 3121
rect 902 3116 903 3120
rect 907 3116 908 3120
rect 902 3115 908 3116
rect 1062 3120 1068 3121
rect 1062 3116 1063 3120
rect 1067 3116 1068 3120
rect 1062 3115 1068 3116
rect 1222 3120 1228 3121
rect 1222 3116 1223 3120
rect 1227 3116 1228 3120
rect 1222 3115 1228 3116
rect 1390 3120 1396 3121
rect 1390 3116 1391 3120
rect 1395 3116 1396 3120
rect 1390 3115 1396 3116
rect 1468 3112 1470 3154
rect 1512 3151 1514 3179
rect 1588 3164 1590 3186
rect 1694 3184 1700 3185
rect 1694 3180 1695 3184
rect 1699 3180 1700 3184
rect 2006 3183 2007 3187
rect 2011 3183 2012 3187
rect 2006 3182 2012 3183
rect 1694 3179 1700 3180
rect 1586 3163 1592 3164
rect 1586 3159 1587 3163
rect 1591 3159 1592 3163
rect 1586 3158 1592 3159
rect 1696 3151 1698 3179
rect 2008 3151 2010 3182
rect 2048 3178 2050 3205
rect 2072 3181 2074 3205
rect 2146 3195 2152 3196
rect 2146 3191 2147 3195
rect 2151 3191 2152 3195
rect 2146 3190 2152 3191
rect 2070 3180 2076 3181
rect 2046 3177 2052 3178
rect 2046 3173 2047 3177
rect 2051 3173 2052 3177
rect 2070 3176 2071 3180
rect 2075 3176 2076 3180
rect 2070 3175 2076 3176
rect 2046 3172 2052 3173
rect 2148 3172 2150 3190
rect 2168 3181 2170 3205
rect 2188 3204 2190 3242
rect 2246 3240 2252 3241
rect 2246 3236 2247 3240
rect 2251 3236 2252 3240
rect 2246 3235 2252 3236
rect 2398 3240 2404 3241
rect 2398 3236 2399 3240
rect 2403 3236 2404 3240
rect 2398 3235 2404 3236
rect 2248 3211 2250 3235
rect 2330 3215 2336 3216
rect 2330 3211 2331 3215
rect 2335 3211 2336 3215
rect 2400 3211 2402 3235
rect 2476 3220 2478 3242
rect 2574 3240 2580 3241
rect 2574 3236 2575 3240
rect 2579 3236 2580 3240
rect 2574 3235 2580 3236
rect 2474 3219 2480 3220
rect 2474 3215 2475 3219
rect 2479 3215 2480 3219
rect 2474 3214 2480 3215
rect 2576 3211 2578 3235
rect 2652 3220 2654 3242
rect 2782 3240 2788 3241
rect 2782 3236 2783 3240
rect 2787 3236 2788 3240
rect 2782 3235 2788 3236
rect 2650 3219 2656 3220
rect 2650 3215 2651 3219
rect 2655 3215 2656 3219
rect 2650 3214 2656 3215
rect 2784 3211 2786 3235
rect 2860 3220 2862 3242
rect 3014 3240 3020 3241
rect 3014 3236 3015 3240
rect 3019 3236 3020 3240
rect 3014 3235 3020 3236
rect 3262 3240 3268 3241
rect 3262 3236 3263 3240
rect 3267 3236 3268 3240
rect 3262 3235 3268 3236
rect 2858 3219 2864 3220
rect 2858 3215 2859 3219
rect 2863 3215 2864 3219
rect 2858 3214 2864 3215
rect 3016 3211 3018 3235
rect 3264 3211 3266 3235
rect 3310 3215 3316 3216
rect 3310 3211 3311 3215
rect 3315 3211 3316 3215
rect 2247 3210 2251 3211
rect 2247 3205 2251 3206
rect 2263 3210 2267 3211
rect 2330 3210 2336 3211
rect 2359 3210 2363 3211
rect 2263 3205 2267 3206
rect 2186 3203 2192 3204
rect 2186 3199 2187 3203
rect 2191 3199 2192 3203
rect 2186 3198 2192 3199
rect 2264 3181 2266 3205
rect 2166 3180 2172 3181
rect 2166 3176 2167 3180
rect 2171 3176 2172 3180
rect 2166 3175 2172 3176
rect 2262 3180 2268 3181
rect 2262 3176 2263 3180
rect 2267 3176 2268 3180
rect 2262 3175 2268 3176
rect 2332 3172 2334 3210
rect 2359 3205 2363 3206
rect 2399 3210 2403 3211
rect 2399 3205 2403 3206
rect 2455 3210 2459 3211
rect 2455 3205 2459 3206
rect 2551 3210 2555 3211
rect 2551 3205 2555 3206
rect 2575 3210 2579 3211
rect 2575 3205 2579 3206
rect 2647 3210 2651 3211
rect 2647 3205 2651 3206
rect 2743 3210 2747 3211
rect 2743 3205 2747 3206
rect 2783 3210 2787 3211
rect 2783 3205 2787 3206
rect 2839 3210 2843 3211
rect 2839 3205 2843 3206
rect 2935 3210 2939 3211
rect 2935 3205 2939 3206
rect 3015 3210 3019 3211
rect 3015 3205 3019 3206
rect 3031 3210 3035 3211
rect 3031 3205 3035 3206
rect 3127 3210 3131 3211
rect 3127 3205 3131 3206
rect 3223 3210 3227 3211
rect 3223 3205 3227 3206
rect 3263 3210 3267 3211
rect 3310 3210 3316 3211
rect 3319 3210 3323 3211
rect 3263 3205 3267 3206
rect 2346 3203 2352 3204
rect 2346 3199 2347 3203
rect 2351 3199 2352 3203
rect 2346 3198 2352 3199
rect 2348 3172 2350 3198
rect 2360 3181 2362 3205
rect 2442 3203 2448 3204
rect 2442 3199 2443 3203
rect 2447 3199 2448 3203
rect 2442 3198 2448 3199
rect 2358 3180 2364 3181
rect 2358 3176 2359 3180
rect 2363 3176 2364 3180
rect 2358 3175 2364 3176
rect 2444 3172 2446 3198
rect 2456 3181 2458 3205
rect 2538 3203 2544 3204
rect 2538 3199 2539 3203
rect 2543 3199 2544 3203
rect 2538 3198 2544 3199
rect 2454 3180 2460 3181
rect 2454 3176 2455 3180
rect 2459 3176 2460 3180
rect 2454 3175 2460 3176
rect 2540 3172 2542 3198
rect 2552 3181 2554 3205
rect 2634 3203 2640 3204
rect 2634 3199 2635 3203
rect 2639 3199 2640 3203
rect 2634 3198 2640 3199
rect 2550 3180 2556 3181
rect 2550 3176 2551 3180
rect 2555 3176 2556 3180
rect 2550 3175 2556 3176
rect 2636 3172 2638 3198
rect 2648 3181 2650 3205
rect 2730 3203 2736 3204
rect 2730 3199 2731 3203
rect 2735 3199 2736 3203
rect 2730 3198 2736 3199
rect 2646 3180 2652 3181
rect 2646 3176 2647 3180
rect 2651 3176 2652 3180
rect 2646 3175 2652 3176
rect 2732 3172 2734 3198
rect 2744 3181 2746 3205
rect 2826 3203 2832 3204
rect 2826 3199 2827 3203
rect 2831 3199 2832 3203
rect 2826 3198 2832 3199
rect 2742 3180 2748 3181
rect 2742 3176 2743 3180
rect 2747 3176 2748 3180
rect 2742 3175 2748 3176
rect 2828 3172 2830 3198
rect 2840 3181 2842 3205
rect 2922 3203 2928 3204
rect 2922 3199 2923 3203
rect 2927 3199 2928 3203
rect 2922 3198 2928 3199
rect 2838 3180 2844 3181
rect 2838 3176 2839 3180
rect 2843 3176 2844 3180
rect 2838 3175 2844 3176
rect 2924 3172 2926 3198
rect 2936 3181 2938 3205
rect 3022 3203 3028 3204
rect 3022 3199 3023 3203
rect 3027 3199 3028 3203
rect 3022 3198 3028 3199
rect 2934 3180 2940 3181
rect 2934 3176 2935 3180
rect 2939 3176 2940 3180
rect 2934 3175 2940 3176
rect 3024 3172 3026 3198
rect 3032 3181 3034 3205
rect 3114 3203 3120 3204
rect 3114 3199 3115 3203
rect 3119 3199 3120 3203
rect 3114 3198 3120 3199
rect 3030 3180 3036 3181
rect 3030 3176 3031 3180
rect 3035 3176 3036 3180
rect 3030 3175 3036 3176
rect 3116 3172 3118 3198
rect 3128 3181 3130 3205
rect 3210 3203 3216 3204
rect 3210 3199 3211 3203
rect 3215 3199 3216 3203
rect 3210 3198 3216 3199
rect 3126 3180 3132 3181
rect 3126 3176 3127 3180
rect 3131 3176 3132 3180
rect 3126 3175 3132 3176
rect 3212 3172 3214 3198
rect 3224 3181 3226 3205
rect 3222 3180 3228 3181
rect 3222 3176 3223 3180
rect 3227 3176 3228 3180
rect 3222 3175 3228 3176
rect 3312 3172 3314 3210
rect 3319 3205 3323 3206
rect 3320 3181 3322 3205
rect 3340 3204 3342 3242
rect 3508 3220 3510 3303
rect 3536 3287 3538 3316
rect 3696 3287 3698 3316
rect 3840 3287 3842 3316
rect 3527 3286 3531 3287
rect 3527 3281 3531 3282
rect 3535 3286 3539 3287
rect 3535 3281 3539 3282
rect 3695 3286 3699 3287
rect 3695 3281 3699 3282
rect 3791 3286 3795 3287
rect 3791 3281 3795 3282
rect 3839 3286 3843 3287
rect 3839 3281 3843 3282
rect 3528 3260 3530 3281
rect 3792 3260 3794 3281
rect 3526 3259 3532 3260
rect 3526 3255 3527 3259
rect 3531 3255 3532 3259
rect 3526 3254 3532 3255
rect 3790 3259 3796 3260
rect 3790 3255 3791 3259
rect 3795 3255 3796 3259
rect 3790 3254 3796 3255
rect 3526 3240 3532 3241
rect 3526 3236 3527 3240
rect 3531 3236 3532 3240
rect 3526 3235 3532 3236
rect 3790 3240 3796 3241
rect 3790 3236 3791 3240
rect 3795 3236 3796 3240
rect 3790 3235 3796 3236
rect 3506 3219 3512 3220
rect 3506 3215 3507 3219
rect 3511 3215 3512 3219
rect 3506 3214 3512 3215
rect 3528 3211 3530 3235
rect 3792 3211 3794 3235
rect 3852 3220 3854 3418
rect 3906 3363 3912 3364
rect 3906 3359 3907 3363
rect 3911 3359 3912 3363
rect 3906 3358 3912 3359
rect 3866 3247 3872 3248
rect 3866 3243 3867 3247
rect 3871 3243 3872 3247
rect 3866 3242 3872 3243
rect 3846 3219 3854 3220
rect 3846 3215 3847 3219
rect 3851 3217 3854 3219
rect 3851 3215 3852 3217
rect 3846 3214 3852 3215
rect 3439 3210 3443 3211
rect 3439 3205 3443 3206
rect 3527 3210 3531 3211
rect 3527 3205 3531 3206
rect 3575 3210 3579 3211
rect 3575 3205 3579 3206
rect 3719 3210 3723 3211
rect 3719 3205 3723 3206
rect 3791 3210 3795 3211
rect 3791 3205 3795 3206
rect 3839 3210 3843 3211
rect 3839 3205 3843 3206
rect 3338 3203 3344 3204
rect 3338 3199 3339 3203
rect 3343 3199 3344 3203
rect 3338 3198 3344 3199
rect 3402 3203 3408 3204
rect 3402 3199 3403 3203
rect 3407 3199 3408 3203
rect 3402 3198 3408 3199
rect 3318 3180 3324 3181
rect 3318 3176 3319 3180
rect 3323 3176 3324 3180
rect 3318 3175 3324 3176
rect 3404 3172 3406 3198
rect 3440 3181 3442 3205
rect 3576 3181 3578 3205
rect 3586 3203 3592 3204
rect 3586 3199 3587 3203
rect 3591 3199 3592 3203
rect 3586 3198 3592 3199
rect 3650 3203 3656 3204
rect 3650 3199 3651 3203
rect 3655 3199 3656 3203
rect 3650 3198 3656 3199
rect 3438 3180 3444 3181
rect 3438 3176 3439 3180
rect 3443 3176 3444 3180
rect 3438 3175 3444 3176
rect 3574 3180 3580 3181
rect 3574 3176 3575 3180
rect 3579 3176 3580 3180
rect 3574 3175 3580 3176
rect 2146 3171 2152 3172
rect 2146 3167 2147 3171
rect 2151 3167 2152 3171
rect 2146 3166 2152 3167
rect 2330 3171 2336 3172
rect 2330 3167 2331 3171
rect 2335 3167 2336 3171
rect 2330 3166 2336 3167
rect 2346 3171 2352 3172
rect 2346 3167 2347 3171
rect 2351 3167 2352 3171
rect 2346 3166 2352 3167
rect 2442 3171 2448 3172
rect 2442 3167 2443 3171
rect 2447 3167 2448 3171
rect 2442 3166 2448 3167
rect 2538 3171 2544 3172
rect 2538 3167 2539 3171
rect 2543 3167 2544 3171
rect 2538 3166 2544 3167
rect 2634 3171 2640 3172
rect 2634 3167 2635 3171
rect 2639 3167 2640 3171
rect 2634 3166 2640 3167
rect 2730 3171 2736 3172
rect 2730 3167 2731 3171
rect 2735 3167 2736 3171
rect 2730 3166 2736 3167
rect 2826 3171 2832 3172
rect 2826 3167 2827 3171
rect 2831 3167 2832 3171
rect 2826 3166 2832 3167
rect 2922 3171 2928 3172
rect 2922 3167 2923 3171
rect 2927 3167 2928 3171
rect 2922 3166 2928 3167
rect 3022 3171 3028 3172
rect 3022 3167 3023 3171
rect 3027 3167 3028 3171
rect 3022 3166 3028 3167
rect 3114 3171 3120 3172
rect 3114 3167 3115 3171
rect 3119 3167 3120 3171
rect 3114 3166 3120 3167
rect 3210 3171 3216 3172
rect 3210 3167 3211 3171
rect 3215 3167 3216 3171
rect 3210 3166 3216 3167
rect 3310 3171 3316 3172
rect 3310 3167 3311 3171
rect 3315 3167 3316 3171
rect 3310 3166 3316 3167
rect 3402 3171 3408 3172
rect 3402 3167 3403 3171
rect 3407 3167 3408 3171
rect 3402 3166 3408 3167
rect 2070 3161 2076 3162
rect 2046 3160 2052 3161
rect 2046 3156 2047 3160
rect 2051 3156 2052 3160
rect 2070 3157 2071 3161
rect 2075 3157 2076 3161
rect 2070 3156 2076 3157
rect 2166 3161 2172 3162
rect 2166 3157 2167 3161
rect 2171 3157 2172 3161
rect 2166 3156 2172 3157
rect 2262 3161 2268 3162
rect 2262 3157 2263 3161
rect 2267 3157 2268 3161
rect 2262 3156 2268 3157
rect 2358 3161 2364 3162
rect 2358 3157 2359 3161
rect 2363 3157 2364 3161
rect 2358 3156 2364 3157
rect 2454 3161 2460 3162
rect 2454 3157 2455 3161
rect 2459 3157 2460 3161
rect 2454 3156 2460 3157
rect 2550 3161 2556 3162
rect 2550 3157 2551 3161
rect 2555 3157 2556 3161
rect 2550 3156 2556 3157
rect 2646 3161 2652 3162
rect 2646 3157 2647 3161
rect 2651 3157 2652 3161
rect 2646 3156 2652 3157
rect 2742 3161 2748 3162
rect 2742 3157 2743 3161
rect 2747 3157 2748 3161
rect 2742 3156 2748 3157
rect 2838 3161 2844 3162
rect 2838 3157 2839 3161
rect 2843 3157 2844 3161
rect 2838 3156 2844 3157
rect 2934 3161 2940 3162
rect 2934 3157 2935 3161
rect 2939 3157 2940 3161
rect 2934 3156 2940 3157
rect 3030 3161 3036 3162
rect 3030 3157 3031 3161
rect 3035 3157 3036 3161
rect 3030 3156 3036 3157
rect 3126 3161 3132 3162
rect 3126 3157 3127 3161
rect 3131 3157 3132 3161
rect 3126 3156 3132 3157
rect 3222 3161 3228 3162
rect 3222 3157 3223 3161
rect 3227 3157 3228 3161
rect 3222 3156 3228 3157
rect 3318 3161 3324 3162
rect 3318 3157 3319 3161
rect 3323 3157 3324 3161
rect 3318 3156 3324 3157
rect 3438 3161 3444 3162
rect 3438 3157 3439 3161
rect 3443 3157 3444 3161
rect 3438 3156 3444 3157
rect 3574 3161 3580 3162
rect 3574 3157 3575 3161
rect 3579 3157 3580 3161
rect 3574 3156 3580 3157
rect 2046 3155 2052 3156
rect 1511 3150 1515 3151
rect 1511 3145 1515 3146
rect 1559 3150 1563 3151
rect 1559 3145 1563 3146
rect 1695 3150 1699 3151
rect 1695 3145 1699 3146
rect 1727 3150 1731 3151
rect 1727 3145 1731 3146
rect 2007 3150 2011 3151
rect 2007 3145 2011 3146
rect 1474 3143 1480 3144
rect 1474 3139 1475 3143
rect 1479 3139 1480 3143
rect 1474 3138 1480 3139
rect 1476 3112 1478 3138
rect 1560 3121 1562 3145
rect 1642 3143 1648 3144
rect 1642 3139 1643 3143
rect 1647 3139 1648 3143
rect 1642 3138 1648 3139
rect 1558 3120 1564 3121
rect 1558 3116 1559 3120
rect 1563 3116 1564 3120
rect 1558 3115 1564 3116
rect 1644 3112 1646 3138
rect 1728 3121 1730 3145
rect 1794 3143 1800 3144
rect 1794 3139 1795 3143
rect 1799 3139 1800 3143
rect 1794 3138 1800 3139
rect 1726 3120 1732 3121
rect 1726 3116 1727 3120
rect 1731 3116 1732 3120
rect 1726 3115 1732 3116
rect 386 3111 392 3112
rect 386 3107 387 3111
rect 391 3107 392 3111
rect 386 3106 392 3107
rect 514 3111 520 3112
rect 514 3107 515 3111
rect 519 3107 520 3111
rect 514 3106 520 3107
rect 658 3111 664 3112
rect 658 3107 659 3111
rect 663 3107 664 3111
rect 658 3106 664 3107
rect 818 3111 824 3112
rect 818 3107 819 3111
rect 823 3107 824 3111
rect 818 3106 824 3107
rect 1350 3111 1356 3112
rect 1350 3107 1351 3111
rect 1355 3107 1356 3111
rect 1350 3106 1356 3107
rect 1466 3111 1472 3112
rect 1466 3107 1467 3111
rect 1471 3107 1472 3111
rect 1466 3106 1472 3107
rect 1474 3111 1480 3112
rect 1474 3107 1475 3111
rect 1479 3107 1480 3111
rect 1474 3106 1480 3107
rect 1642 3111 1648 3112
rect 1642 3107 1643 3111
rect 1647 3107 1648 3111
rect 1642 3106 1648 3107
rect 438 3101 444 3102
rect 438 3097 439 3101
rect 443 3097 444 3101
rect 438 3096 444 3097
rect 582 3101 588 3102
rect 582 3097 583 3101
rect 587 3097 588 3101
rect 582 3096 588 3097
rect 742 3101 748 3102
rect 742 3097 743 3101
rect 747 3097 748 3101
rect 742 3096 748 3097
rect 902 3101 908 3102
rect 902 3097 903 3101
rect 907 3097 908 3101
rect 902 3096 908 3097
rect 1062 3101 1068 3102
rect 1062 3097 1063 3101
rect 1067 3097 1068 3101
rect 1062 3096 1068 3097
rect 1222 3101 1228 3102
rect 1222 3097 1223 3101
rect 1227 3097 1228 3101
rect 1222 3096 1228 3097
rect 440 3067 442 3096
rect 584 3067 586 3096
rect 744 3067 746 3096
rect 904 3067 906 3096
rect 1064 3067 1066 3096
rect 1224 3067 1226 3096
rect 439 3066 443 3067
rect 439 3061 443 3062
rect 503 3066 507 3067
rect 503 3061 507 3062
rect 583 3066 587 3067
rect 583 3061 587 3062
rect 599 3066 603 3067
rect 599 3061 603 3062
rect 703 3066 707 3067
rect 703 3061 707 3062
rect 743 3066 747 3067
rect 743 3061 747 3062
rect 815 3066 819 3067
rect 815 3061 819 3062
rect 903 3066 907 3067
rect 903 3061 907 3062
rect 935 3066 939 3067
rect 935 3061 939 3062
rect 1063 3066 1067 3067
rect 1063 3061 1067 3062
rect 1071 3066 1075 3067
rect 1071 3061 1075 3062
rect 1223 3066 1227 3067
rect 1223 3061 1227 3062
rect 504 3040 506 3061
rect 600 3040 602 3061
rect 704 3040 706 3061
rect 816 3040 818 3061
rect 936 3040 938 3061
rect 1072 3040 1074 3061
rect 1224 3040 1226 3061
rect 502 3039 508 3040
rect 502 3035 503 3039
rect 507 3035 508 3039
rect 502 3034 508 3035
rect 598 3039 604 3040
rect 598 3035 599 3039
rect 603 3035 604 3039
rect 598 3034 604 3035
rect 702 3039 708 3040
rect 702 3035 703 3039
rect 707 3035 708 3039
rect 702 3034 708 3035
rect 814 3039 820 3040
rect 814 3035 815 3039
rect 819 3035 820 3039
rect 814 3034 820 3035
rect 934 3039 940 3040
rect 934 3035 935 3039
rect 939 3035 940 3039
rect 934 3034 940 3035
rect 1070 3039 1076 3040
rect 1070 3035 1071 3039
rect 1075 3035 1076 3039
rect 1070 3034 1076 3035
rect 1222 3039 1228 3040
rect 1222 3035 1223 3039
rect 1227 3035 1228 3039
rect 1222 3034 1228 3035
rect 366 3031 372 3032
rect 366 3027 367 3031
rect 371 3027 372 3031
rect 366 3026 372 3027
rect 586 3031 592 3032
rect 586 3027 587 3031
rect 591 3027 592 3031
rect 586 3026 592 3027
rect 682 3031 688 3032
rect 682 3027 683 3031
rect 687 3027 688 3031
rect 682 3026 688 3027
rect 806 3031 812 3032
rect 806 3027 807 3031
rect 811 3027 812 3031
rect 806 3026 812 3027
rect 902 3031 908 3032
rect 902 3027 903 3031
rect 907 3027 908 3031
rect 1342 3031 1348 3032
rect 902 3026 908 3027
rect 1146 3027 1152 3028
rect 110 3023 116 3024
rect 110 3019 111 3023
rect 115 3019 116 3023
rect 110 3018 116 3019
rect 502 3020 508 3021
rect 112 2987 114 3018
rect 502 3016 503 3020
rect 507 3016 508 3020
rect 502 3015 508 3016
rect 504 2987 506 3015
rect 588 3000 590 3026
rect 598 3020 604 3021
rect 598 3016 599 3020
rect 603 3016 604 3020
rect 598 3015 604 3016
rect 586 2999 592 3000
rect 586 2995 587 2999
rect 591 2995 592 2999
rect 586 2994 592 2995
rect 600 2987 602 3015
rect 684 3000 686 3026
rect 702 3020 708 3021
rect 702 3016 703 3020
rect 707 3016 708 3020
rect 702 3015 708 3016
rect 682 2999 688 3000
rect 682 2995 683 2999
rect 687 2995 688 2999
rect 682 2994 688 2995
rect 704 2987 706 3015
rect 808 3000 810 3026
rect 814 3020 820 3021
rect 814 3016 815 3020
rect 819 3016 820 3020
rect 814 3015 820 3016
rect 806 2999 812 3000
rect 806 2995 807 2999
rect 811 2995 812 2999
rect 806 2994 812 2995
rect 816 2987 818 3015
rect 904 3000 906 3026
rect 1146 3023 1147 3027
rect 1151 3023 1152 3027
rect 1342 3027 1343 3031
rect 1347 3027 1348 3031
rect 1342 3026 1348 3027
rect 1146 3022 1152 3023
rect 934 3020 940 3021
rect 934 3016 935 3020
rect 939 3016 940 3020
rect 934 3015 940 3016
rect 1070 3020 1076 3021
rect 1070 3016 1071 3020
rect 1075 3016 1076 3020
rect 1070 3015 1076 3016
rect 902 2999 908 3000
rect 902 2995 903 2999
rect 907 2995 908 2999
rect 902 2994 908 2995
rect 936 2987 938 3015
rect 990 2995 996 2996
rect 990 2991 991 2995
rect 995 2991 996 2995
rect 990 2990 996 2991
rect 111 2986 115 2987
rect 111 2981 115 2982
rect 503 2986 507 2987
rect 503 2981 507 2982
rect 551 2986 555 2987
rect 551 2981 555 2982
rect 599 2986 603 2987
rect 599 2981 603 2982
rect 647 2986 651 2987
rect 647 2981 651 2982
rect 703 2986 707 2987
rect 703 2981 707 2982
rect 759 2986 763 2987
rect 759 2981 763 2982
rect 815 2986 819 2987
rect 815 2981 819 2982
rect 887 2986 891 2987
rect 887 2981 891 2982
rect 935 2986 939 2987
rect 935 2981 939 2982
rect 112 2954 114 2981
rect 552 2957 554 2981
rect 626 2979 632 2980
rect 626 2975 627 2979
rect 631 2975 632 2979
rect 626 2974 632 2975
rect 550 2956 556 2957
rect 110 2953 116 2954
rect 110 2949 111 2953
rect 115 2949 116 2953
rect 550 2952 551 2956
rect 555 2952 556 2956
rect 550 2951 556 2952
rect 110 2948 116 2949
rect 628 2948 630 2974
rect 648 2957 650 2981
rect 722 2979 728 2980
rect 722 2975 723 2979
rect 727 2975 728 2979
rect 722 2974 728 2975
rect 646 2956 652 2957
rect 646 2952 647 2956
rect 651 2952 652 2956
rect 646 2951 652 2952
rect 724 2948 726 2974
rect 760 2957 762 2981
rect 834 2979 840 2980
rect 834 2975 835 2979
rect 839 2975 840 2979
rect 834 2974 840 2975
rect 758 2956 764 2957
rect 758 2952 759 2956
rect 763 2952 764 2956
rect 758 2951 764 2952
rect 836 2948 838 2974
rect 888 2957 890 2981
rect 962 2979 968 2980
rect 962 2975 963 2979
rect 967 2975 968 2979
rect 962 2974 968 2975
rect 922 2971 928 2972
rect 922 2967 923 2971
rect 927 2967 928 2971
rect 922 2966 928 2967
rect 886 2956 892 2957
rect 886 2952 887 2956
rect 891 2952 892 2956
rect 886 2951 892 2952
rect 626 2947 632 2948
rect 626 2943 627 2947
rect 631 2943 632 2947
rect 626 2942 632 2943
rect 722 2947 728 2948
rect 722 2943 723 2947
rect 727 2943 728 2947
rect 722 2942 728 2943
rect 834 2947 840 2948
rect 834 2943 835 2947
rect 839 2943 840 2947
rect 834 2942 840 2943
rect 550 2937 556 2938
rect 110 2936 116 2937
rect 110 2932 111 2936
rect 115 2932 116 2936
rect 550 2933 551 2937
rect 555 2933 556 2937
rect 550 2932 556 2933
rect 646 2937 652 2938
rect 646 2933 647 2937
rect 651 2933 652 2937
rect 646 2932 652 2933
rect 758 2937 764 2938
rect 758 2933 759 2937
rect 763 2933 764 2937
rect 758 2932 764 2933
rect 886 2937 892 2938
rect 886 2933 887 2937
rect 891 2933 892 2937
rect 886 2932 892 2933
rect 110 2931 116 2932
rect 112 2903 114 2931
rect 552 2903 554 2932
rect 648 2903 650 2932
rect 760 2903 762 2932
rect 888 2903 890 2932
rect 111 2902 115 2903
rect 111 2897 115 2898
rect 471 2902 475 2903
rect 471 2897 475 2898
rect 551 2902 555 2903
rect 551 2897 555 2898
rect 575 2902 579 2903
rect 575 2897 579 2898
rect 647 2902 651 2903
rect 647 2897 651 2898
rect 695 2902 699 2903
rect 695 2897 699 2898
rect 759 2902 763 2903
rect 759 2897 763 2898
rect 839 2902 843 2903
rect 839 2897 843 2898
rect 887 2902 891 2903
rect 887 2897 891 2898
rect 112 2877 114 2897
rect 110 2876 116 2877
rect 472 2876 474 2897
rect 576 2876 578 2897
rect 696 2876 698 2897
rect 840 2876 842 2897
rect 110 2872 111 2876
rect 115 2872 116 2876
rect 110 2871 116 2872
rect 470 2875 476 2876
rect 470 2871 471 2875
rect 475 2871 476 2875
rect 470 2870 476 2871
rect 574 2875 580 2876
rect 574 2871 575 2875
rect 579 2871 580 2875
rect 574 2870 580 2871
rect 694 2875 700 2876
rect 694 2871 695 2875
rect 699 2871 700 2875
rect 694 2870 700 2871
rect 838 2875 844 2876
rect 838 2871 839 2875
rect 843 2871 844 2875
rect 838 2870 844 2871
rect 924 2868 926 2966
rect 964 2948 966 2974
rect 992 2948 994 2990
rect 1072 2987 1074 3015
rect 1023 2986 1027 2987
rect 1023 2981 1027 2982
rect 1071 2986 1075 2987
rect 1071 2981 1075 2982
rect 1024 2957 1026 2981
rect 1148 2980 1150 3022
rect 1222 3020 1228 3021
rect 1222 3016 1223 3020
rect 1227 3016 1228 3020
rect 1222 3015 1228 3016
rect 1224 2987 1226 3015
rect 1344 3000 1346 3026
rect 1352 3000 1354 3106
rect 1390 3101 1396 3102
rect 1390 3097 1391 3101
rect 1395 3097 1396 3101
rect 1390 3096 1396 3097
rect 1558 3101 1564 3102
rect 1558 3097 1559 3101
rect 1563 3097 1564 3101
rect 1558 3096 1564 3097
rect 1726 3101 1732 3102
rect 1726 3097 1727 3101
rect 1731 3097 1732 3101
rect 1726 3096 1732 3097
rect 1392 3067 1394 3096
rect 1560 3067 1562 3096
rect 1728 3067 1730 3096
rect 1383 3066 1387 3067
rect 1383 3061 1387 3062
rect 1391 3066 1395 3067
rect 1391 3061 1395 3062
rect 1551 3066 1555 3067
rect 1551 3061 1555 3062
rect 1559 3066 1563 3067
rect 1559 3061 1563 3062
rect 1719 3066 1723 3067
rect 1719 3061 1723 3062
rect 1727 3066 1731 3067
rect 1727 3061 1731 3062
rect 1384 3040 1386 3061
rect 1552 3040 1554 3061
rect 1720 3040 1722 3061
rect 1382 3039 1388 3040
rect 1382 3035 1383 3039
rect 1387 3035 1388 3039
rect 1382 3034 1388 3035
rect 1550 3039 1556 3040
rect 1550 3035 1551 3039
rect 1555 3035 1556 3039
rect 1550 3034 1556 3035
rect 1718 3039 1724 3040
rect 1718 3035 1719 3039
rect 1723 3035 1724 3039
rect 1718 3034 1724 3035
rect 1796 3032 1798 3138
rect 2008 3118 2010 3145
rect 2048 3123 2050 3155
rect 2072 3123 2074 3156
rect 2168 3123 2170 3156
rect 2264 3123 2266 3156
rect 2298 3155 2304 3156
rect 2298 3151 2299 3155
rect 2303 3151 2304 3155
rect 2298 3150 2304 3151
rect 2047 3122 2051 3123
rect 2006 3117 2012 3118
rect 2047 3117 2051 3118
rect 2071 3122 2075 3123
rect 2071 3117 2075 3118
rect 2167 3122 2171 3123
rect 2167 3117 2171 3118
rect 2263 3122 2267 3123
rect 2263 3117 2267 3118
rect 2006 3113 2007 3117
rect 2011 3113 2012 3117
rect 2006 3112 2012 3113
rect 2006 3100 2012 3101
rect 2006 3096 2007 3100
rect 2011 3096 2012 3100
rect 2048 3097 2050 3117
rect 2006 3095 2012 3096
rect 2046 3096 2052 3097
rect 2072 3096 2074 3117
rect 2008 3067 2010 3095
rect 2046 3092 2047 3096
rect 2051 3092 2052 3096
rect 2046 3091 2052 3092
rect 2070 3095 2076 3096
rect 2070 3091 2071 3095
rect 2075 3091 2076 3095
rect 2070 3090 2076 3091
rect 2182 3087 2188 3088
rect 2146 3083 2152 3084
rect 2046 3079 2052 3080
rect 2046 3075 2047 3079
rect 2051 3075 2052 3079
rect 2146 3079 2147 3083
rect 2151 3079 2152 3083
rect 2182 3083 2183 3087
rect 2187 3083 2188 3087
rect 2182 3082 2188 3083
rect 2146 3078 2152 3079
rect 2046 3074 2052 3075
rect 2070 3076 2076 3077
rect 2007 3066 2011 3067
rect 2007 3061 2011 3062
rect 2008 3041 2010 3061
rect 2048 3047 2050 3074
rect 2070 3072 2071 3076
rect 2075 3072 2076 3076
rect 2070 3071 2076 3072
rect 2072 3047 2074 3071
rect 2047 3046 2051 3047
rect 2047 3041 2051 3042
rect 2071 3046 2075 3047
rect 2071 3041 2075 3042
rect 2006 3040 2012 3041
rect 2006 3036 2007 3040
rect 2011 3036 2012 3040
rect 2006 3035 2012 3036
rect 1794 3031 1800 3032
rect 1626 3027 1632 3028
rect 1626 3023 1627 3027
rect 1631 3023 1632 3027
rect 1794 3027 1795 3031
rect 1799 3027 1800 3031
rect 1794 3026 1800 3027
rect 1626 3022 1632 3023
rect 2006 3023 2012 3024
rect 1382 3020 1388 3021
rect 1382 3016 1383 3020
rect 1387 3016 1388 3020
rect 1382 3015 1388 3016
rect 1550 3020 1556 3021
rect 1550 3016 1551 3020
rect 1555 3016 1556 3020
rect 1550 3015 1556 3016
rect 1342 2999 1348 3000
rect 1342 2995 1343 2999
rect 1347 2995 1348 2999
rect 1342 2994 1348 2995
rect 1350 2999 1356 3000
rect 1350 2995 1351 2999
rect 1355 2995 1356 2999
rect 1350 2994 1356 2995
rect 1384 2987 1386 3015
rect 1552 2987 1554 3015
rect 1628 3000 1630 3022
rect 1718 3020 1724 3021
rect 1718 3016 1719 3020
rect 1723 3016 1724 3020
rect 2006 3019 2007 3023
rect 2011 3019 2012 3023
rect 2006 3018 2012 3019
rect 1718 3015 1724 3016
rect 1626 2999 1632 3000
rect 1562 2995 1568 2996
rect 1562 2991 1563 2995
rect 1567 2991 1568 2995
rect 1626 2995 1627 2999
rect 1631 2995 1632 2999
rect 1626 2994 1632 2995
rect 1562 2990 1568 2991
rect 1175 2986 1179 2987
rect 1175 2981 1179 2982
rect 1223 2986 1227 2987
rect 1223 2981 1227 2982
rect 1327 2986 1331 2987
rect 1327 2981 1331 2982
rect 1383 2986 1387 2987
rect 1383 2981 1387 2982
rect 1487 2986 1491 2987
rect 1487 2981 1491 2982
rect 1551 2986 1555 2987
rect 1551 2981 1555 2982
rect 1146 2979 1152 2980
rect 1146 2975 1147 2979
rect 1151 2975 1152 2979
rect 1146 2974 1152 2975
rect 1176 2957 1178 2981
rect 1250 2979 1256 2980
rect 1250 2975 1251 2979
rect 1255 2975 1256 2979
rect 1250 2974 1256 2975
rect 1022 2956 1028 2957
rect 1022 2952 1023 2956
rect 1027 2952 1028 2956
rect 1022 2951 1028 2952
rect 1174 2956 1180 2957
rect 1174 2952 1175 2956
rect 1179 2952 1180 2956
rect 1174 2951 1180 2952
rect 1252 2948 1254 2974
rect 1328 2957 1330 2981
rect 1488 2957 1490 2981
rect 1326 2956 1332 2957
rect 1326 2952 1327 2956
rect 1331 2952 1332 2956
rect 1326 2951 1332 2952
rect 1486 2956 1492 2957
rect 1486 2952 1487 2956
rect 1491 2952 1492 2956
rect 1486 2951 1492 2952
rect 1564 2948 1566 2990
rect 1720 2987 1722 3015
rect 2008 2987 2010 3018
rect 2048 3014 2050 3041
rect 2072 3017 2074 3041
rect 2148 3040 2150 3078
rect 2184 3056 2186 3082
rect 2300 3056 2302 3150
rect 2360 3123 2362 3156
rect 2456 3123 2458 3156
rect 2552 3123 2554 3156
rect 2648 3123 2650 3156
rect 2744 3123 2746 3156
rect 2840 3123 2842 3156
rect 2936 3123 2938 3156
rect 3032 3123 3034 3156
rect 3128 3123 3130 3156
rect 3224 3123 3226 3156
rect 3320 3123 3322 3156
rect 3440 3123 3442 3156
rect 3576 3123 3578 3156
rect 2335 3122 2339 3123
rect 2335 3117 2339 3118
rect 2359 3122 2363 3123
rect 2359 3117 2363 3118
rect 2455 3122 2459 3123
rect 2455 3117 2459 3118
rect 2551 3122 2555 3123
rect 2551 3117 2555 3118
rect 2623 3122 2627 3123
rect 2623 3117 2627 3118
rect 2647 3122 2651 3123
rect 2647 3117 2651 3118
rect 2743 3122 2747 3123
rect 2743 3117 2747 3118
rect 2839 3122 2843 3123
rect 2839 3117 2843 3118
rect 2911 3122 2915 3123
rect 2911 3117 2915 3118
rect 2935 3122 2939 3123
rect 2935 3117 2939 3118
rect 3031 3122 3035 3123
rect 3031 3117 3035 3118
rect 3127 3122 3131 3123
rect 3127 3117 3131 3118
rect 3207 3122 3211 3123
rect 3207 3117 3211 3118
rect 3223 3122 3227 3123
rect 3223 3117 3227 3118
rect 3319 3122 3323 3123
rect 3319 3117 3323 3118
rect 3439 3122 3443 3123
rect 3439 3117 3443 3118
rect 3503 3122 3507 3123
rect 3503 3117 3507 3118
rect 3575 3122 3579 3123
rect 3575 3117 3579 3118
rect 2336 3096 2338 3117
rect 2624 3096 2626 3117
rect 2912 3096 2914 3117
rect 3208 3096 3210 3117
rect 3504 3096 3506 3117
rect 2334 3095 2340 3096
rect 2334 3091 2335 3095
rect 2339 3091 2340 3095
rect 2334 3090 2340 3091
rect 2622 3095 2628 3096
rect 2622 3091 2623 3095
rect 2627 3091 2628 3095
rect 2622 3090 2628 3091
rect 2910 3095 2916 3096
rect 2910 3091 2911 3095
rect 2915 3091 2916 3095
rect 2910 3090 2916 3091
rect 3206 3095 3212 3096
rect 3206 3091 3207 3095
rect 3211 3091 3212 3095
rect 3206 3090 3212 3091
rect 3502 3095 3508 3096
rect 3502 3091 3503 3095
rect 3507 3091 3508 3095
rect 3502 3090 3508 3091
rect 3588 3088 3590 3198
rect 3652 3172 3654 3198
rect 3658 3195 3664 3196
rect 3658 3191 3659 3195
rect 3663 3191 3664 3195
rect 3658 3190 3664 3191
rect 3660 3172 3662 3190
rect 3720 3181 3722 3205
rect 3840 3181 3842 3205
rect 3718 3180 3724 3181
rect 3718 3176 3719 3180
rect 3723 3176 3724 3180
rect 3718 3175 3724 3176
rect 3838 3180 3844 3181
rect 3838 3176 3839 3180
rect 3843 3176 3844 3180
rect 3838 3175 3844 3176
rect 3650 3171 3656 3172
rect 3650 3167 3651 3171
rect 3655 3167 3656 3171
rect 3650 3166 3656 3167
rect 3658 3171 3664 3172
rect 3658 3167 3659 3171
rect 3663 3167 3664 3171
rect 3658 3166 3664 3167
rect 3718 3161 3724 3162
rect 3718 3157 3719 3161
rect 3723 3157 3724 3161
rect 3718 3156 3724 3157
rect 3838 3161 3844 3162
rect 3838 3157 3839 3161
rect 3843 3157 3844 3161
rect 3838 3156 3844 3157
rect 3720 3123 3722 3156
rect 3840 3123 3842 3156
rect 3719 3122 3723 3123
rect 3719 3117 3723 3118
rect 3799 3122 3803 3123
rect 3799 3117 3803 3118
rect 3839 3122 3843 3123
rect 3839 3117 3843 3118
rect 3800 3096 3802 3117
rect 3798 3095 3804 3096
rect 3798 3091 3799 3095
rect 3803 3091 3804 3095
rect 3798 3090 3804 3091
rect 3586 3087 3592 3088
rect 2698 3083 2704 3084
rect 2698 3079 2699 3083
rect 2703 3079 2704 3083
rect 2698 3078 2704 3079
rect 2986 3083 2992 3084
rect 2986 3079 2987 3083
rect 2991 3079 2992 3083
rect 2986 3078 2992 3079
rect 3282 3083 3288 3084
rect 3282 3079 3283 3083
rect 3287 3079 3288 3083
rect 3586 3083 3587 3087
rect 3591 3083 3592 3087
rect 3586 3082 3592 3083
rect 3282 3078 3288 3079
rect 2334 3076 2340 3077
rect 2334 3072 2335 3076
rect 2339 3072 2340 3076
rect 2334 3071 2340 3072
rect 2622 3076 2628 3077
rect 2622 3072 2623 3076
rect 2627 3072 2628 3076
rect 2622 3071 2628 3072
rect 2182 3055 2188 3056
rect 2182 3051 2183 3055
rect 2187 3051 2188 3055
rect 2182 3050 2188 3051
rect 2298 3055 2304 3056
rect 2298 3051 2299 3055
rect 2303 3051 2304 3055
rect 2298 3050 2304 3051
rect 2336 3047 2338 3071
rect 2624 3047 2626 3071
rect 2700 3056 2702 3078
rect 2910 3076 2916 3077
rect 2910 3072 2911 3076
rect 2915 3072 2916 3076
rect 2910 3071 2916 3072
rect 2698 3055 2704 3056
rect 2674 3051 2680 3052
rect 2674 3047 2675 3051
rect 2679 3047 2680 3051
rect 2698 3051 2699 3055
rect 2703 3051 2704 3055
rect 2698 3050 2704 3051
rect 2912 3047 2914 3071
rect 2988 3056 2990 3078
rect 3206 3076 3212 3077
rect 3206 3072 3207 3076
rect 3211 3072 3212 3076
rect 3206 3071 3212 3072
rect 2986 3055 2992 3056
rect 2986 3051 2987 3055
rect 2991 3051 2992 3055
rect 2986 3050 2992 3051
rect 3208 3047 3210 3071
rect 3284 3056 3286 3078
rect 3502 3076 3508 3077
rect 3502 3072 3503 3076
rect 3507 3072 3508 3076
rect 3502 3071 3508 3072
rect 3798 3076 3804 3077
rect 3798 3072 3799 3076
rect 3803 3072 3804 3076
rect 3798 3071 3804 3072
rect 3282 3055 3288 3056
rect 3282 3051 3283 3055
rect 3287 3051 3288 3055
rect 3282 3050 3288 3051
rect 3504 3047 3506 3071
rect 3800 3047 3802 3071
rect 3868 3056 3870 3242
rect 3908 3172 3910 3358
rect 3916 3332 3918 3530
rect 3944 3510 3946 3537
rect 3942 3509 3948 3510
rect 3942 3505 3943 3509
rect 3947 3505 3948 3509
rect 3942 3504 3948 3505
rect 3942 3492 3948 3493
rect 3942 3488 3943 3492
rect 3947 3488 3948 3492
rect 3942 3487 3948 3488
rect 3944 3463 3946 3487
rect 3943 3462 3947 3463
rect 3943 3457 3947 3458
rect 3944 3437 3946 3457
rect 3942 3436 3948 3437
rect 3942 3432 3943 3436
rect 3947 3432 3948 3436
rect 3942 3431 3948 3432
rect 3942 3419 3948 3420
rect 3942 3415 3943 3419
rect 3947 3415 3948 3419
rect 3942 3414 3948 3415
rect 3944 3371 3946 3414
rect 3943 3370 3947 3371
rect 3943 3365 3947 3366
rect 3944 3338 3946 3365
rect 3942 3337 3948 3338
rect 3942 3333 3943 3337
rect 3947 3333 3948 3337
rect 3942 3332 3948 3333
rect 3914 3331 3920 3332
rect 3914 3327 3915 3331
rect 3919 3327 3920 3331
rect 3914 3326 3920 3327
rect 3942 3320 3948 3321
rect 3942 3316 3943 3320
rect 3947 3316 3948 3320
rect 3942 3315 3948 3316
rect 3944 3287 3946 3315
rect 3943 3286 3947 3287
rect 3943 3281 3947 3282
rect 3944 3261 3946 3281
rect 3942 3260 3948 3261
rect 3942 3256 3943 3260
rect 3947 3256 3948 3260
rect 3942 3255 3948 3256
rect 3942 3243 3948 3244
rect 3942 3239 3943 3243
rect 3947 3239 3948 3243
rect 3942 3238 3948 3239
rect 3944 3211 3946 3238
rect 3943 3210 3947 3211
rect 3943 3205 3947 3206
rect 3914 3203 3920 3204
rect 3914 3199 3915 3203
rect 3919 3199 3920 3203
rect 3914 3198 3920 3199
rect 3906 3171 3912 3172
rect 3906 3167 3907 3171
rect 3911 3167 3912 3171
rect 3906 3166 3912 3167
rect 3874 3083 3880 3084
rect 3874 3079 3875 3083
rect 3879 3079 3880 3083
rect 3874 3078 3880 3079
rect 3866 3055 3872 3056
rect 3866 3051 3867 3055
rect 3871 3051 3872 3055
rect 3866 3050 3872 3051
rect 2335 3046 2339 3047
rect 2335 3041 2339 3042
rect 2383 3046 2387 3047
rect 2383 3041 2387 3042
rect 2623 3046 2627 3047
rect 2674 3046 2680 3047
rect 2703 3046 2707 3047
rect 2623 3041 2627 3042
rect 2146 3039 2152 3040
rect 2146 3035 2147 3039
rect 2151 3035 2152 3039
rect 2146 3034 2152 3035
rect 2384 3017 2386 3041
rect 2070 3016 2076 3017
rect 2046 3013 2052 3014
rect 2046 3009 2047 3013
rect 2051 3009 2052 3013
rect 2070 3012 2071 3016
rect 2075 3012 2076 3016
rect 2070 3011 2076 3012
rect 2382 3016 2388 3017
rect 2382 3012 2383 3016
rect 2387 3012 2388 3016
rect 2382 3011 2388 3012
rect 2046 3008 2052 3009
rect 2676 3008 2678 3046
rect 2703 3041 2707 3042
rect 2911 3046 2915 3047
rect 2911 3041 2915 3042
rect 2999 3046 3003 3047
rect 2999 3041 3003 3042
rect 3207 3046 3211 3047
rect 3207 3041 3211 3042
rect 3287 3046 3291 3047
rect 3287 3041 3291 3042
rect 3503 3046 3507 3047
rect 3503 3041 3507 3042
rect 3575 3046 3579 3047
rect 3575 3041 3579 3042
rect 3799 3046 3803 3047
rect 3799 3041 3803 3042
rect 3839 3046 3843 3047
rect 3839 3041 3843 3042
rect 2704 3017 2706 3041
rect 2958 3039 2964 3040
rect 2958 3035 2959 3039
rect 2963 3035 2964 3039
rect 2958 3034 2964 3035
rect 2702 3016 2708 3017
rect 2702 3012 2703 3016
rect 2707 3012 2708 3016
rect 2702 3011 2708 3012
rect 2960 3008 2962 3034
rect 3000 3017 3002 3041
rect 3258 3039 3264 3040
rect 3258 3035 3259 3039
rect 3263 3035 3264 3039
rect 3258 3034 3264 3035
rect 2998 3016 3004 3017
rect 2998 3012 2999 3016
rect 3003 3012 3004 3016
rect 2998 3011 3004 3012
rect 3260 3008 3262 3034
rect 3288 3017 3290 3041
rect 3370 3039 3376 3040
rect 3370 3035 3371 3039
rect 3375 3035 3376 3039
rect 3370 3034 3376 3035
rect 3286 3016 3292 3017
rect 3286 3012 3287 3016
rect 3291 3012 3292 3016
rect 3286 3011 3292 3012
rect 3372 3008 3374 3034
rect 3576 3017 3578 3041
rect 3840 3017 3842 3041
rect 3574 3016 3580 3017
rect 3574 3012 3575 3016
rect 3579 3012 3580 3016
rect 3574 3011 3580 3012
rect 3838 3016 3844 3017
rect 3838 3012 3839 3016
rect 3843 3012 3844 3016
rect 3838 3011 3844 3012
rect 2450 3007 2456 3008
rect 2450 3003 2451 3007
rect 2455 3003 2456 3007
rect 2450 3002 2456 3003
rect 2674 3007 2680 3008
rect 2674 3003 2675 3007
rect 2679 3003 2680 3007
rect 2674 3002 2680 3003
rect 2958 3007 2964 3008
rect 2958 3003 2959 3007
rect 2963 3003 2964 3007
rect 2958 3002 2964 3003
rect 3258 3007 3264 3008
rect 3258 3003 3259 3007
rect 3263 3003 3264 3007
rect 3258 3002 3264 3003
rect 3370 3007 3376 3008
rect 3370 3003 3371 3007
rect 3375 3003 3376 3007
rect 3370 3002 3376 3003
rect 2070 2997 2076 2998
rect 2046 2996 2052 2997
rect 2046 2992 2047 2996
rect 2051 2992 2052 2996
rect 2070 2993 2071 2997
rect 2075 2993 2076 2997
rect 2070 2992 2076 2993
rect 2382 2997 2388 2998
rect 2382 2993 2383 2997
rect 2387 2993 2388 2997
rect 2382 2992 2388 2993
rect 2046 2991 2052 2992
rect 1655 2986 1659 2987
rect 1655 2981 1659 2982
rect 1719 2986 1723 2987
rect 1719 2981 1723 2982
rect 1823 2986 1827 2987
rect 1823 2981 1827 2982
rect 2007 2986 2011 2987
rect 2007 2981 2011 2982
rect 1570 2979 1576 2980
rect 1570 2975 1571 2979
rect 1575 2975 1576 2979
rect 1570 2974 1576 2975
rect 1572 2948 1574 2974
rect 1656 2957 1658 2981
rect 1738 2979 1744 2980
rect 1738 2975 1739 2979
rect 1743 2975 1744 2979
rect 1738 2974 1744 2975
rect 1654 2956 1660 2957
rect 1654 2952 1655 2956
rect 1659 2952 1660 2956
rect 1654 2951 1660 2952
rect 1740 2948 1742 2974
rect 1824 2957 1826 2981
rect 1922 2979 1928 2980
rect 1922 2975 1923 2979
rect 1927 2975 1928 2979
rect 1922 2974 1928 2975
rect 1822 2956 1828 2957
rect 1822 2952 1823 2956
rect 1827 2952 1828 2956
rect 1822 2951 1828 2952
rect 962 2947 968 2948
rect 962 2943 963 2947
rect 967 2943 968 2947
rect 962 2942 968 2943
rect 990 2947 996 2948
rect 990 2943 991 2947
rect 995 2943 996 2947
rect 990 2942 996 2943
rect 1250 2947 1256 2948
rect 1250 2943 1251 2947
rect 1255 2943 1256 2947
rect 1250 2942 1256 2943
rect 1562 2947 1568 2948
rect 1562 2943 1563 2947
rect 1567 2943 1568 2947
rect 1562 2942 1568 2943
rect 1570 2947 1576 2948
rect 1570 2943 1571 2947
rect 1575 2943 1576 2947
rect 1570 2942 1576 2943
rect 1738 2947 1744 2948
rect 1738 2943 1739 2947
rect 1743 2943 1744 2947
rect 1738 2942 1744 2943
rect 1022 2937 1028 2938
rect 1022 2933 1023 2937
rect 1027 2933 1028 2937
rect 1022 2932 1028 2933
rect 1174 2937 1180 2938
rect 1174 2933 1175 2937
rect 1179 2933 1180 2937
rect 1174 2932 1180 2933
rect 1326 2937 1332 2938
rect 1326 2933 1327 2937
rect 1331 2933 1332 2937
rect 1326 2932 1332 2933
rect 1486 2937 1492 2938
rect 1486 2933 1487 2937
rect 1491 2933 1492 2937
rect 1486 2932 1492 2933
rect 1654 2937 1660 2938
rect 1654 2933 1655 2937
rect 1659 2933 1660 2937
rect 1654 2932 1660 2933
rect 1822 2937 1828 2938
rect 1822 2933 1823 2937
rect 1827 2933 1828 2937
rect 1822 2932 1828 2933
rect 1024 2903 1026 2932
rect 1176 2903 1178 2932
rect 1328 2903 1330 2932
rect 1488 2903 1490 2932
rect 1656 2903 1658 2932
rect 1824 2903 1826 2932
rect 991 2902 995 2903
rect 991 2897 995 2898
rect 1023 2902 1027 2903
rect 1023 2897 1027 2898
rect 1151 2902 1155 2903
rect 1151 2897 1155 2898
rect 1175 2902 1179 2903
rect 1175 2897 1179 2898
rect 1319 2902 1323 2903
rect 1319 2897 1323 2898
rect 1327 2902 1331 2903
rect 1327 2897 1331 2898
rect 1487 2902 1491 2903
rect 1487 2897 1491 2898
rect 1495 2902 1499 2903
rect 1495 2897 1499 2898
rect 1655 2902 1659 2903
rect 1655 2897 1659 2898
rect 1671 2902 1675 2903
rect 1671 2897 1675 2898
rect 1823 2902 1827 2903
rect 1823 2897 1827 2898
rect 1847 2902 1851 2903
rect 1847 2897 1851 2898
rect 992 2876 994 2897
rect 1152 2876 1154 2897
rect 1320 2876 1322 2897
rect 1496 2876 1498 2897
rect 1672 2876 1674 2897
rect 1848 2876 1850 2897
rect 990 2875 996 2876
rect 990 2871 991 2875
rect 995 2871 996 2875
rect 990 2870 996 2871
rect 1150 2875 1156 2876
rect 1150 2871 1151 2875
rect 1155 2871 1156 2875
rect 1150 2870 1156 2871
rect 1318 2875 1324 2876
rect 1318 2871 1319 2875
rect 1323 2871 1324 2875
rect 1318 2870 1324 2871
rect 1494 2875 1500 2876
rect 1494 2871 1495 2875
rect 1499 2871 1500 2875
rect 1494 2870 1500 2871
rect 1670 2875 1676 2876
rect 1670 2871 1671 2875
rect 1675 2871 1676 2875
rect 1670 2870 1676 2871
rect 1846 2875 1852 2876
rect 1846 2871 1847 2875
rect 1851 2871 1852 2875
rect 1846 2870 1852 2871
rect 1924 2868 1926 2974
rect 2008 2954 2010 2981
rect 2048 2967 2050 2991
rect 2072 2967 2074 2992
rect 2384 2967 2386 2992
rect 2047 2966 2051 2967
rect 2047 2961 2051 2962
rect 2071 2966 2075 2967
rect 2071 2961 2075 2962
rect 2383 2966 2387 2967
rect 2383 2961 2387 2962
rect 2391 2966 2395 2967
rect 2391 2961 2395 2962
rect 2006 2953 2012 2954
rect 2006 2949 2007 2953
rect 2011 2949 2012 2953
rect 2006 2948 2012 2949
rect 2048 2941 2050 2961
rect 2046 2940 2052 2941
rect 2072 2940 2074 2961
rect 2392 2940 2394 2961
rect 2006 2936 2012 2937
rect 2006 2932 2007 2936
rect 2011 2932 2012 2936
rect 2046 2936 2047 2940
rect 2051 2936 2052 2940
rect 2046 2935 2052 2936
rect 2070 2939 2076 2940
rect 2070 2935 2071 2939
rect 2075 2935 2076 2939
rect 2070 2934 2076 2935
rect 2390 2939 2396 2940
rect 2390 2935 2391 2939
rect 2395 2935 2396 2939
rect 2390 2934 2396 2935
rect 2006 2931 2012 2932
rect 2008 2903 2010 2931
rect 2146 2927 2152 2928
rect 2046 2923 2052 2924
rect 2046 2919 2047 2923
rect 2051 2919 2052 2923
rect 2146 2923 2147 2927
rect 2151 2923 2152 2927
rect 2146 2922 2152 2923
rect 2046 2918 2052 2919
rect 2070 2920 2076 2921
rect 2007 2902 2011 2903
rect 2007 2897 2011 2898
rect 2008 2877 2010 2897
rect 2048 2891 2050 2918
rect 2070 2916 2071 2920
rect 2075 2916 2076 2920
rect 2070 2915 2076 2916
rect 2072 2891 2074 2915
rect 2047 2890 2051 2891
rect 2047 2885 2051 2886
rect 2071 2890 2075 2891
rect 2071 2885 2075 2886
rect 2006 2876 2012 2877
rect 2006 2872 2007 2876
rect 2011 2872 2012 2876
rect 2006 2871 2012 2872
rect 922 2867 928 2868
rect 566 2863 572 2864
rect 110 2859 116 2860
rect 110 2855 111 2859
rect 115 2855 116 2859
rect 566 2859 567 2863
rect 571 2859 572 2863
rect 566 2858 572 2859
rect 650 2863 656 2864
rect 650 2859 651 2863
rect 655 2859 656 2863
rect 650 2858 656 2859
rect 770 2863 776 2864
rect 770 2859 771 2863
rect 775 2859 776 2863
rect 770 2858 776 2859
rect 914 2863 920 2864
rect 914 2859 915 2863
rect 919 2859 920 2863
rect 922 2863 923 2867
rect 927 2863 928 2867
rect 1922 2867 1928 2868
rect 922 2862 928 2863
rect 1226 2863 1232 2864
rect 914 2858 920 2859
rect 1226 2859 1227 2863
rect 1231 2859 1232 2863
rect 1226 2858 1232 2859
rect 1394 2863 1400 2864
rect 1394 2859 1395 2863
rect 1399 2859 1400 2863
rect 1394 2858 1400 2859
rect 1630 2863 1636 2864
rect 1630 2859 1631 2863
rect 1635 2859 1636 2863
rect 1630 2858 1636 2859
rect 1746 2863 1752 2864
rect 1746 2859 1747 2863
rect 1751 2859 1752 2863
rect 1922 2863 1923 2867
rect 1927 2863 1928 2867
rect 1922 2862 1928 2863
rect 1746 2858 1752 2859
rect 2006 2859 2012 2860
rect 110 2854 116 2855
rect 470 2856 476 2857
rect 112 2823 114 2854
rect 470 2852 471 2856
rect 475 2852 476 2856
rect 470 2851 476 2852
rect 472 2823 474 2851
rect 568 2836 570 2858
rect 574 2856 580 2857
rect 574 2852 575 2856
rect 579 2852 580 2856
rect 574 2851 580 2852
rect 566 2835 572 2836
rect 546 2831 552 2832
rect 546 2827 547 2831
rect 551 2827 552 2831
rect 566 2831 567 2835
rect 571 2831 572 2835
rect 566 2830 572 2831
rect 546 2826 552 2827
rect 111 2822 115 2823
rect 111 2817 115 2818
rect 471 2822 475 2823
rect 471 2817 475 2818
rect 479 2822 483 2823
rect 479 2817 483 2818
rect 112 2790 114 2817
rect 480 2793 482 2817
rect 478 2792 484 2793
rect 110 2789 116 2790
rect 110 2785 111 2789
rect 115 2785 116 2789
rect 478 2788 479 2792
rect 483 2788 484 2792
rect 478 2787 484 2788
rect 110 2784 116 2785
rect 548 2784 550 2826
rect 576 2823 578 2851
rect 652 2836 654 2858
rect 694 2856 700 2857
rect 694 2852 695 2856
rect 699 2852 700 2856
rect 694 2851 700 2852
rect 650 2835 656 2836
rect 650 2831 651 2835
rect 655 2831 656 2835
rect 650 2830 656 2831
rect 696 2823 698 2851
rect 772 2836 774 2858
rect 838 2856 844 2857
rect 838 2852 839 2856
rect 843 2852 844 2856
rect 838 2851 844 2852
rect 770 2835 776 2836
rect 770 2831 771 2835
rect 775 2831 776 2835
rect 770 2830 776 2831
rect 840 2823 842 2851
rect 916 2836 918 2858
rect 990 2856 996 2857
rect 990 2852 991 2856
rect 995 2852 996 2856
rect 990 2851 996 2852
rect 1150 2856 1156 2857
rect 1150 2852 1151 2856
rect 1155 2852 1156 2856
rect 1150 2851 1156 2852
rect 914 2835 920 2836
rect 914 2831 915 2835
rect 919 2831 920 2835
rect 914 2830 920 2831
rect 992 2823 994 2851
rect 1152 2823 1154 2851
rect 1228 2836 1230 2858
rect 1318 2856 1324 2857
rect 1318 2852 1319 2856
rect 1323 2852 1324 2856
rect 1318 2851 1324 2852
rect 1226 2835 1232 2836
rect 1226 2831 1227 2835
rect 1231 2831 1232 2835
rect 1226 2830 1232 2831
rect 1320 2823 1322 2851
rect 575 2822 579 2823
rect 575 2817 579 2818
rect 679 2822 683 2823
rect 679 2817 683 2818
rect 695 2822 699 2823
rect 695 2817 699 2818
rect 799 2822 803 2823
rect 799 2817 803 2818
rect 839 2822 843 2823
rect 839 2817 843 2818
rect 935 2822 939 2823
rect 935 2817 939 2818
rect 991 2822 995 2823
rect 991 2817 995 2818
rect 1079 2822 1083 2823
rect 1079 2817 1083 2818
rect 1151 2822 1155 2823
rect 1151 2817 1155 2818
rect 1239 2822 1243 2823
rect 1239 2817 1243 2818
rect 1319 2822 1323 2823
rect 1319 2817 1323 2818
rect 562 2815 568 2816
rect 562 2811 563 2815
rect 567 2811 568 2815
rect 562 2810 568 2811
rect 564 2784 566 2810
rect 576 2793 578 2817
rect 658 2815 664 2816
rect 658 2811 659 2815
rect 663 2811 664 2815
rect 658 2810 664 2811
rect 574 2792 580 2793
rect 574 2788 575 2792
rect 579 2788 580 2792
rect 574 2787 580 2788
rect 660 2784 662 2810
rect 680 2793 682 2817
rect 762 2815 768 2816
rect 762 2811 763 2815
rect 767 2811 768 2815
rect 762 2810 768 2811
rect 678 2792 684 2793
rect 678 2788 679 2792
rect 683 2788 684 2792
rect 678 2787 684 2788
rect 764 2784 766 2810
rect 800 2793 802 2817
rect 882 2815 888 2816
rect 882 2811 883 2815
rect 887 2811 888 2815
rect 882 2810 888 2811
rect 798 2792 804 2793
rect 798 2788 799 2792
rect 803 2788 804 2792
rect 798 2787 804 2788
rect 884 2784 886 2810
rect 936 2793 938 2817
rect 998 2815 1004 2816
rect 998 2811 999 2815
rect 1003 2811 1004 2815
rect 998 2810 1004 2811
rect 934 2792 940 2793
rect 934 2788 935 2792
rect 939 2788 940 2792
rect 934 2787 940 2788
rect 546 2783 552 2784
rect 546 2779 547 2783
rect 551 2779 552 2783
rect 546 2778 552 2779
rect 562 2783 568 2784
rect 562 2779 563 2783
rect 567 2779 568 2783
rect 562 2778 568 2779
rect 658 2783 664 2784
rect 658 2779 659 2783
rect 663 2779 664 2783
rect 658 2778 664 2779
rect 762 2783 768 2784
rect 762 2779 763 2783
rect 767 2779 768 2783
rect 762 2778 768 2779
rect 882 2783 888 2784
rect 882 2779 883 2783
rect 887 2779 888 2783
rect 882 2778 888 2779
rect 478 2773 484 2774
rect 110 2772 116 2773
rect 110 2768 111 2772
rect 115 2768 116 2772
rect 478 2769 479 2773
rect 483 2769 484 2773
rect 478 2768 484 2769
rect 574 2773 580 2774
rect 574 2769 575 2773
rect 579 2769 580 2773
rect 574 2768 580 2769
rect 678 2773 684 2774
rect 678 2769 679 2773
rect 683 2769 684 2773
rect 678 2768 684 2769
rect 798 2773 804 2774
rect 798 2769 799 2773
rect 803 2769 804 2773
rect 798 2768 804 2769
rect 934 2773 940 2774
rect 934 2769 935 2773
rect 939 2769 940 2773
rect 934 2768 940 2769
rect 110 2767 116 2768
rect 112 2743 114 2767
rect 480 2743 482 2768
rect 576 2743 578 2768
rect 680 2743 682 2768
rect 800 2743 802 2768
rect 936 2743 938 2768
rect 111 2742 115 2743
rect 111 2737 115 2738
rect 479 2742 483 2743
rect 479 2737 483 2738
rect 511 2742 515 2743
rect 511 2737 515 2738
rect 575 2742 579 2743
rect 575 2737 579 2738
rect 623 2742 627 2743
rect 623 2737 627 2738
rect 679 2742 683 2743
rect 679 2737 683 2738
rect 743 2742 747 2743
rect 743 2737 747 2738
rect 799 2742 803 2743
rect 799 2737 803 2738
rect 879 2742 883 2743
rect 879 2737 883 2738
rect 935 2742 939 2743
rect 935 2737 939 2738
rect 112 2717 114 2737
rect 110 2716 116 2717
rect 512 2716 514 2737
rect 624 2716 626 2737
rect 744 2716 746 2737
rect 880 2716 882 2737
rect 110 2712 111 2716
rect 115 2712 116 2716
rect 110 2711 116 2712
rect 510 2715 516 2716
rect 510 2711 511 2715
rect 515 2711 516 2715
rect 510 2710 516 2711
rect 622 2715 628 2716
rect 622 2711 623 2715
rect 627 2711 628 2715
rect 622 2710 628 2711
rect 742 2715 748 2716
rect 742 2711 743 2715
rect 747 2711 748 2715
rect 742 2710 748 2711
rect 878 2715 884 2716
rect 878 2711 879 2715
rect 883 2711 884 2715
rect 878 2710 884 2711
rect 1000 2708 1002 2810
rect 1080 2793 1082 2817
rect 1190 2815 1196 2816
rect 1190 2811 1191 2815
rect 1195 2811 1196 2815
rect 1190 2810 1196 2811
rect 1078 2792 1084 2793
rect 1078 2788 1079 2792
rect 1083 2788 1084 2792
rect 1078 2787 1084 2788
rect 1192 2784 1194 2810
rect 1240 2793 1242 2817
rect 1396 2816 1398 2858
rect 1494 2856 1500 2857
rect 1494 2852 1495 2856
rect 1499 2852 1500 2856
rect 1494 2851 1500 2852
rect 1496 2823 1498 2851
rect 1632 2836 1634 2858
rect 1670 2856 1676 2857
rect 1670 2852 1671 2856
rect 1675 2852 1676 2856
rect 1670 2851 1676 2852
rect 1630 2835 1636 2836
rect 1550 2831 1556 2832
rect 1550 2827 1551 2831
rect 1555 2827 1556 2831
rect 1630 2831 1631 2835
rect 1635 2831 1636 2835
rect 1630 2830 1636 2831
rect 1550 2826 1556 2827
rect 1415 2822 1419 2823
rect 1415 2817 1419 2818
rect 1495 2822 1499 2823
rect 1495 2817 1499 2818
rect 1326 2815 1332 2816
rect 1326 2811 1327 2815
rect 1331 2811 1332 2815
rect 1326 2810 1332 2811
rect 1394 2815 1400 2816
rect 1394 2811 1395 2815
rect 1399 2811 1400 2815
rect 1394 2810 1400 2811
rect 1238 2792 1244 2793
rect 1238 2788 1239 2792
rect 1243 2788 1244 2792
rect 1238 2787 1244 2788
rect 1328 2784 1330 2810
rect 1416 2793 1418 2817
rect 1414 2792 1420 2793
rect 1414 2788 1415 2792
rect 1419 2788 1420 2792
rect 1414 2787 1420 2788
rect 1552 2784 1554 2826
rect 1672 2823 1674 2851
rect 1748 2836 1750 2858
rect 1846 2856 1852 2857
rect 1846 2852 1847 2856
rect 1851 2852 1852 2856
rect 2006 2855 2007 2859
rect 2011 2855 2012 2859
rect 2048 2858 2050 2885
rect 2072 2861 2074 2885
rect 2148 2884 2150 2922
rect 2390 2920 2396 2921
rect 2390 2916 2391 2920
rect 2395 2916 2396 2920
rect 2390 2915 2396 2916
rect 2392 2891 2394 2915
rect 2452 2900 2454 3002
rect 2702 2997 2708 2998
rect 2702 2993 2703 2997
rect 2707 2993 2708 2997
rect 2702 2992 2708 2993
rect 2998 2997 3004 2998
rect 2998 2993 2999 2997
rect 3003 2993 3004 2997
rect 2998 2992 3004 2993
rect 3286 2997 3292 2998
rect 3286 2993 3287 2997
rect 3291 2993 3292 2997
rect 3286 2992 3292 2993
rect 3574 2997 3580 2998
rect 3574 2993 3575 2997
rect 3579 2993 3580 2997
rect 3574 2992 3580 2993
rect 3838 2997 3844 2998
rect 3838 2993 3839 2997
rect 3843 2993 3844 2997
rect 3838 2992 3844 2993
rect 2704 2967 2706 2992
rect 3000 2967 3002 2992
rect 3288 2967 3290 2992
rect 3576 2967 3578 2992
rect 3840 2967 3842 2992
rect 2703 2966 2707 2967
rect 2703 2961 2707 2962
rect 2975 2966 2979 2967
rect 2975 2961 2979 2962
rect 2999 2966 3003 2967
rect 2999 2961 3003 2962
rect 3215 2966 3219 2967
rect 3215 2961 3219 2962
rect 3287 2966 3291 2967
rect 3287 2961 3291 2962
rect 3439 2966 3443 2967
rect 3439 2961 3443 2962
rect 3575 2966 3579 2967
rect 3575 2961 3579 2962
rect 3647 2966 3651 2967
rect 3647 2961 3651 2962
rect 3839 2966 3843 2967
rect 3839 2961 3843 2962
rect 2704 2940 2706 2961
rect 2976 2940 2978 2961
rect 3216 2940 3218 2961
rect 3440 2940 3442 2961
rect 3648 2940 3650 2961
rect 3840 2940 3842 2961
rect 2702 2939 2708 2940
rect 2702 2935 2703 2939
rect 2707 2935 2708 2939
rect 2702 2934 2708 2935
rect 2974 2939 2980 2940
rect 2974 2935 2975 2939
rect 2979 2935 2980 2939
rect 2974 2934 2980 2935
rect 3214 2939 3220 2940
rect 3214 2935 3215 2939
rect 3219 2935 3220 2939
rect 3214 2934 3220 2935
rect 3438 2939 3444 2940
rect 3438 2935 3439 2939
rect 3443 2935 3444 2939
rect 3438 2934 3444 2935
rect 3646 2939 3652 2940
rect 3646 2935 3647 2939
rect 3651 2935 3652 2939
rect 3646 2934 3652 2935
rect 3838 2939 3844 2940
rect 3838 2935 3839 2939
rect 3843 2935 3844 2939
rect 3838 2934 3844 2935
rect 2778 2927 2784 2928
rect 2778 2923 2779 2927
rect 2783 2923 2784 2927
rect 2778 2922 2784 2923
rect 3050 2927 3056 2928
rect 3050 2923 3051 2927
rect 3055 2923 3056 2927
rect 3050 2922 3056 2923
rect 3290 2927 3296 2928
rect 3290 2923 3291 2927
rect 3295 2923 3296 2927
rect 3290 2922 3296 2923
rect 3514 2927 3520 2928
rect 3514 2923 3515 2927
rect 3519 2923 3520 2927
rect 3514 2922 3520 2923
rect 3722 2927 3728 2928
rect 3722 2923 3723 2927
rect 3727 2923 3728 2927
rect 3722 2922 3728 2923
rect 2702 2920 2708 2921
rect 2702 2916 2703 2920
rect 2707 2916 2708 2920
rect 2702 2915 2708 2916
rect 2446 2899 2454 2900
rect 2446 2895 2447 2899
rect 2451 2897 2454 2899
rect 2451 2895 2452 2897
rect 2446 2894 2452 2895
rect 2704 2891 2706 2915
rect 2780 2892 2782 2922
rect 2974 2920 2980 2921
rect 2974 2916 2975 2920
rect 2979 2916 2980 2920
rect 2974 2915 2980 2916
rect 2778 2891 2784 2892
rect 2976 2891 2978 2915
rect 3052 2900 3054 2922
rect 3214 2920 3220 2921
rect 3214 2916 3215 2920
rect 3219 2916 3220 2920
rect 3214 2915 3220 2916
rect 3050 2899 3056 2900
rect 3050 2895 3051 2899
rect 3055 2895 3056 2899
rect 3050 2894 3056 2895
rect 3216 2891 3218 2915
rect 3292 2900 3294 2922
rect 3438 2920 3444 2921
rect 3438 2916 3439 2920
rect 3443 2916 3444 2920
rect 3438 2915 3444 2916
rect 3290 2899 3296 2900
rect 3290 2895 3291 2899
rect 3295 2895 3296 2899
rect 3290 2894 3296 2895
rect 3440 2891 3442 2915
rect 3516 2900 3518 2922
rect 3646 2920 3652 2921
rect 3646 2916 3647 2920
rect 3651 2916 3652 2920
rect 3646 2915 3652 2916
rect 3618 2907 3624 2908
rect 3618 2903 3619 2907
rect 3623 2903 3624 2907
rect 3618 2902 3624 2903
rect 3514 2899 3520 2900
rect 3514 2895 3515 2899
rect 3519 2895 3520 2899
rect 3514 2894 3520 2895
rect 2295 2890 2299 2891
rect 2295 2885 2299 2886
rect 2391 2890 2395 2891
rect 2391 2885 2395 2886
rect 2535 2890 2539 2891
rect 2535 2885 2539 2886
rect 2703 2890 2707 2891
rect 2703 2885 2707 2886
rect 2767 2890 2771 2891
rect 2778 2887 2779 2891
rect 2783 2887 2784 2891
rect 2778 2886 2784 2887
rect 2975 2890 2979 2891
rect 2767 2885 2771 2886
rect 2975 2885 2979 2886
rect 2991 2890 2995 2891
rect 2991 2885 2995 2886
rect 3215 2890 3219 2891
rect 3215 2885 3219 2886
rect 3431 2890 3435 2891
rect 3431 2885 3435 2886
rect 3439 2890 3443 2891
rect 3439 2885 3443 2886
rect 2146 2883 2152 2884
rect 2146 2879 2147 2883
rect 2151 2879 2152 2883
rect 2146 2878 2152 2879
rect 2230 2883 2236 2884
rect 2230 2879 2231 2883
rect 2235 2879 2236 2883
rect 2230 2878 2236 2879
rect 2070 2860 2076 2861
rect 2006 2854 2012 2855
rect 2046 2857 2052 2858
rect 1846 2851 1852 2852
rect 1746 2835 1752 2836
rect 1746 2831 1747 2835
rect 1751 2831 1752 2835
rect 1746 2830 1752 2831
rect 1848 2823 1850 2851
rect 2008 2823 2010 2854
rect 2046 2853 2047 2857
rect 2051 2853 2052 2857
rect 2070 2856 2071 2860
rect 2075 2856 2076 2860
rect 2070 2855 2076 2856
rect 2046 2852 2052 2853
rect 2232 2852 2234 2878
rect 2296 2861 2298 2885
rect 2370 2883 2376 2884
rect 2370 2879 2371 2883
rect 2375 2879 2376 2883
rect 2370 2878 2376 2879
rect 2294 2860 2300 2861
rect 2294 2856 2295 2860
rect 2299 2856 2300 2860
rect 2294 2855 2300 2856
rect 2372 2852 2374 2878
rect 2536 2861 2538 2885
rect 2610 2883 2616 2884
rect 2610 2879 2611 2883
rect 2615 2879 2616 2883
rect 2610 2878 2616 2879
rect 2534 2860 2540 2861
rect 2534 2856 2535 2860
rect 2539 2856 2540 2860
rect 2534 2855 2540 2856
rect 2612 2852 2614 2878
rect 2768 2861 2770 2885
rect 2992 2861 2994 2885
rect 3066 2883 3072 2884
rect 3066 2879 3067 2883
rect 3071 2879 3072 2883
rect 3066 2878 3072 2879
rect 2766 2860 2772 2861
rect 2766 2856 2767 2860
rect 2771 2856 2772 2860
rect 2766 2855 2772 2856
rect 2990 2860 2996 2861
rect 2990 2856 2991 2860
rect 2995 2856 2996 2860
rect 2990 2855 2996 2856
rect 3068 2852 3070 2878
rect 3216 2861 3218 2885
rect 3290 2883 3296 2884
rect 3290 2879 3291 2883
rect 3295 2879 3296 2883
rect 3290 2878 3296 2879
rect 3214 2860 3220 2861
rect 3214 2856 3215 2860
rect 3219 2856 3220 2860
rect 3214 2855 3220 2856
rect 3292 2852 3294 2878
rect 3432 2861 3434 2885
rect 3506 2883 3512 2884
rect 3506 2879 3507 2883
rect 3511 2879 3512 2883
rect 3506 2878 3512 2879
rect 3438 2875 3444 2876
rect 3438 2871 3439 2875
rect 3443 2871 3444 2875
rect 3438 2870 3444 2871
rect 3430 2860 3436 2861
rect 3430 2856 3431 2860
rect 3435 2856 3436 2860
rect 3430 2855 3436 2856
rect 2230 2851 2236 2852
rect 2230 2847 2231 2851
rect 2235 2847 2236 2851
rect 2230 2846 2236 2847
rect 2370 2851 2376 2852
rect 2370 2847 2371 2851
rect 2375 2847 2376 2851
rect 2370 2846 2376 2847
rect 2610 2851 2616 2852
rect 2610 2847 2611 2851
rect 2615 2847 2616 2851
rect 2610 2846 2616 2847
rect 2718 2851 2724 2852
rect 2718 2847 2719 2851
rect 2723 2847 2724 2851
rect 2718 2846 2724 2847
rect 3066 2851 3072 2852
rect 3066 2847 3067 2851
rect 3071 2847 3072 2851
rect 3066 2846 3072 2847
rect 3290 2851 3296 2852
rect 3290 2847 3291 2851
rect 3295 2847 3296 2851
rect 3290 2846 3296 2847
rect 2070 2841 2076 2842
rect 2046 2840 2052 2841
rect 2046 2836 2047 2840
rect 2051 2836 2052 2840
rect 2070 2837 2071 2841
rect 2075 2837 2076 2841
rect 2070 2836 2076 2837
rect 2294 2841 2300 2842
rect 2294 2837 2295 2841
rect 2299 2837 2300 2841
rect 2294 2836 2300 2837
rect 2534 2841 2540 2842
rect 2534 2837 2535 2841
rect 2539 2837 2540 2841
rect 2534 2836 2540 2837
rect 2046 2835 2052 2836
rect 1599 2822 1603 2823
rect 1599 2817 1603 2818
rect 1671 2822 1675 2823
rect 1671 2817 1675 2818
rect 1783 2822 1787 2823
rect 1783 2817 1787 2818
rect 1847 2822 1851 2823
rect 1847 2817 1851 2818
rect 2007 2822 2011 2823
rect 2007 2817 2011 2818
rect 1600 2793 1602 2817
rect 1682 2815 1688 2816
rect 1682 2811 1683 2815
rect 1687 2811 1688 2815
rect 1682 2810 1688 2811
rect 1598 2792 1604 2793
rect 1598 2788 1599 2792
rect 1603 2788 1604 2792
rect 1598 2787 1604 2788
rect 1684 2784 1686 2810
rect 1784 2793 1786 2817
rect 1858 2815 1864 2816
rect 1858 2811 1859 2815
rect 1863 2811 1864 2815
rect 1858 2810 1864 2811
rect 1782 2792 1788 2793
rect 1782 2788 1783 2792
rect 1787 2788 1788 2792
rect 1782 2787 1788 2788
rect 1150 2783 1156 2784
rect 1150 2779 1151 2783
rect 1155 2779 1156 2783
rect 1150 2778 1156 2779
rect 1190 2783 1196 2784
rect 1190 2779 1191 2783
rect 1195 2779 1196 2783
rect 1190 2778 1196 2779
rect 1326 2783 1332 2784
rect 1326 2779 1327 2783
rect 1331 2779 1332 2783
rect 1326 2778 1332 2779
rect 1550 2783 1556 2784
rect 1550 2779 1551 2783
rect 1555 2779 1556 2783
rect 1550 2778 1556 2779
rect 1682 2783 1688 2784
rect 1682 2779 1683 2783
rect 1687 2779 1688 2783
rect 1682 2778 1688 2779
rect 1078 2773 1084 2774
rect 1078 2769 1079 2773
rect 1083 2769 1084 2773
rect 1078 2768 1084 2769
rect 1080 2743 1082 2768
rect 1015 2742 1019 2743
rect 1015 2737 1019 2738
rect 1079 2742 1083 2743
rect 1079 2737 1083 2738
rect 1016 2716 1018 2737
rect 1014 2715 1020 2716
rect 1014 2711 1015 2715
rect 1019 2711 1020 2715
rect 1014 2710 1020 2711
rect 998 2707 1004 2708
rect 586 2703 592 2704
rect 110 2699 116 2700
rect 110 2695 111 2699
rect 115 2695 116 2699
rect 586 2699 587 2703
rect 591 2699 592 2703
rect 586 2698 592 2699
rect 698 2703 704 2704
rect 698 2699 699 2703
rect 703 2699 704 2703
rect 698 2698 704 2699
rect 818 2703 824 2704
rect 818 2699 819 2703
rect 823 2699 824 2703
rect 818 2698 824 2699
rect 954 2703 960 2704
rect 954 2699 955 2703
rect 959 2699 960 2703
rect 998 2703 999 2707
rect 1003 2703 1004 2707
rect 998 2702 1004 2703
rect 954 2698 960 2699
rect 110 2694 116 2695
rect 510 2696 516 2697
rect 112 2663 114 2694
rect 510 2692 511 2696
rect 515 2692 516 2696
rect 510 2691 516 2692
rect 512 2663 514 2691
rect 588 2676 590 2698
rect 622 2696 628 2697
rect 622 2692 623 2696
rect 627 2692 628 2696
rect 622 2691 628 2692
rect 586 2675 592 2676
rect 586 2671 587 2675
rect 591 2671 592 2675
rect 586 2670 592 2671
rect 624 2663 626 2691
rect 700 2676 702 2698
rect 742 2696 748 2697
rect 742 2692 743 2696
rect 747 2692 748 2696
rect 742 2691 748 2692
rect 698 2675 704 2676
rect 698 2671 699 2675
rect 703 2671 704 2675
rect 698 2670 704 2671
rect 744 2663 746 2691
rect 820 2676 822 2698
rect 878 2696 884 2697
rect 878 2692 879 2696
rect 883 2692 884 2696
rect 878 2691 884 2692
rect 818 2675 824 2676
rect 818 2671 819 2675
rect 823 2671 824 2675
rect 818 2670 824 2671
rect 858 2667 864 2668
rect 858 2663 859 2667
rect 863 2663 864 2667
rect 880 2663 882 2691
rect 956 2676 958 2698
rect 1014 2696 1020 2697
rect 1014 2692 1015 2696
rect 1019 2692 1020 2696
rect 1014 2691 1020 2692
rect 954 2675 960 2676
rect 954 2671 955 2675
rect 959 2671 960 2675
rect 954 2670 960 2671
rect 1016 2663 1018 2691
rect 1152 2676 1154 2778
rect 1238 2773 1244 2774
rect 1238 2769 1239 2773
rect 1243 2769 1244 2773
rect 1238 2768 1244 2769
rect 1414 2773 1420 2774
rect 1414 2769 1415 2773
rect 1419 2769 1420 2773
rect 1414 2768 1420 2769
rect 1598 2773 1604 2774
rect 1598 2769 1599 2773
rect 1603 2769 1604 2773
rect 1598 2768 1604 2769
rect 1782 2773 1788 2774
rect 1782 2769 1783 2773
rect 1787 2769 1788 2773
rect 1782 2768 1788 2769
rect 1240 2743 1242 2768
rect 1416 2743 1418 2768
rect 1600 2743 1602 2768
rect 1784 2743 1786 2768
rect 1159 2742 1163 2743
rect 1159 2737 1163 2738
rect 1239 2742 1243 2743
rect 1239 2737 1243 2738
rect 1311 2742 1315 2743
rect 1311 2737 1315 2738
rect 1415 2742 1419 2743
rect 1415 2737 1419 2738
rect 1463 2742 1467 2743
rect 1463 2737 1467 2738
rect 1599 2742 1603 2743
rect 1599 2737 1603 2738
rect 1623 2742 1627 2743
rect 1623 2737 1627 2738
rect 1783 2742 1787 2743
rect 1783 2737 1787 2738
rect 1160 2716 1162 2737
rect 1312 2716 1314 2737
rect 1464 2716 1466 2737
rect 1624 2716 1626 2737
rect 1784 2716 1786 2737
rect 1158 2715 1164 2716
rect 1158 2711 1159 2715
rect 1163 2711 1164 2715
rect 1158 2710 1164 2711
rect 1310 2715 1316 2716
rect 1310 2711 1311 2715
rect 1315 2711 1316 2715
rect 1310 2710 1316 2711
rect 1462 2715 1468 2716
rect 1462 2711 1463 2715
rect 1467 2711 1468 2715
rect 1462 2710 1468 2711
rect 1622 2715 1628 2716
rect 1622 2711 1623 2715
rect 1627 2711 1628 2715
rect 1622 2710 1628 2711
rect 1782 2715 1788 2716
rect 1782 2711 1783 2715
rect 1787 2711 1788 2715
rect 1782 2710 1788 2711
rect 1860 2708 1862 2810
rect 2008 2790 2010 2817
rect 2048 2811 2050 2835
rect 2072 2811 2074 2836
rect 2296 2811 2298 2836
rect 2536 2811 2538 2836
rect 2047 2810 2051 2811
rect 2047 2805 2051 2806
rect 2071 2810 2075 2811
rect 2071 2805 2075 2806
rect 2199 2810 2203 2811
rect 2199 2805 2203 2806
rect 2295 2810 2299 2811
rect 2295 2805 2299 2806
rect 2367 2810 2371 2811
rect 2367 2805 2371 2806
rect 2535 2810 2539 2811
rect 2535 2805 2539 2806
rect 2551 2810 2555 2811
rect 2551 2805 2555 2806
rect 2006 2789 2012 2790
rect 2006 2785 2007 2789
rect 2011 2785 2012 2789
rect 2048 2785 2050 2805
rect 2006 2784 2012 2785
rect 2046 2784 2052 2785
rect 2072 2784 2074 2805
rect 2200 2784 2202 2805
rect 2368 2784 2370 2805
rect 2552 2784 2554 2805
rect 2046 2780 2047 2784
rect 2051 2780 2052 2784
rect 2046 2779 2052 2780
rect 2070 2783 2076 2784
rect 2070 2779 2071 2783
rect 2075 2779 2076 2783
rect 2070 2778 2076 2779
rect 2198 2783 2204 2784
rect 2198 2779 2199 2783
rect 2203 2779 2204 2783
rect 2198 2778 2204 2779
rect 2366 2783 2372 2784
rect 2366 2779 2367 2783
rect 2371 2779 2372 2783
rect 2366 2778 2372 2779
rect 2550 2783 2556 2784
rect 2550 2779 2551 2783
rect 2555 2779 2556 2783
rect 2550 2778 2556 2779
rect 2658 2775 2664 2776
rect 2006 2772 2012 2773
rect 2006 2768 2007 2772
rect 2011 2768 2012 2772
rect 2146 2771 2152 2772
rect 2006 2767 2012 2768
rect 2046 2767 2052 2768
rect 2008 2743 2010 2767
rect 2046 2763 2047 2767
rect 2051 2763 2052 2767
rect 2146 2767 2147 2771
rect 2151 2767 2152 2771
rect 2146 2766 2152 2767
rect 2274 2771 2280 2772
rect 2274 2767 2275 2771
rect 2279 2767 2280 2771
rect 2274 2766 2280 2767
rect 2442 2771 2448 2772
rect 2442 2767 2443 2771
rect 2447 2767 2448 2771
rect 2442 2766 2448 2767
rect 2626 2771 2632 2772
rect 2626 2767 2627 2771
rect 2631 2767 2632 2771
rect 2658 2771 2659 2775
rect 2663 2771 2664 2775
rect 2658 2770 2664 2771
rect 2626 2766 2632 2767
rect 2046 2762 2052 2763
rect 2070 2764 2076 2765
rect 2007 2742 2011 2743
rect 2007 2737 2011 2738
rect 2008 2717 2010 2737
rect 2048 2731 2050 2762
rect 2070 2760 2071 2764
rect 2075 2760 2076 2764
rect 2070 2759 2076 2760
rect 2072 2731 2074 2759
rect 2148 2744 2150 2766
rect 2198 2764 2204 2765
rect 2198 2760 2199 2764
rect 2203 2760 2204 2764
rect 2198 2759 2204 2760
rect 2146 2743 2152 2744
rect 2146 2739 2147 2743
rect 2151 2739 2152 2743
rect 2146 2738 2152 2739
rect 2200 2731 2202 2759
rect 2276 2744 2278 2766
rect 2366 2764 2372 2765
rect 2366 2760 2367 2764
rect 2371 2760 2372 2764
rect 2366 2759 2372 2760
rect 2274 2743 2280 2744
rect 2274 2739 2275 2743
rect 2279 2739 2280 2743
rect 2274 2738 2280 2739
rect 2368 2731 2370 2759
rect 2444 2744 2446 2766
rect 2550 2764 2556 2765
rect 2550 2760 2551 2764
rect 2555 2760 2556 2764
rect 2550 2759 2556 2760
rect 2442 2743 2448 2744
rect 2442 2739 2443 2743
rect 2447 2739 2448 2743
rect 2442 2738 2448 2739
rect 2552 2731 2554 2759
rect 2628 2744 2630 2766
rect 2626 2743 2632 2744
rect 2626 2739 2627 2743
rect 2631 2739 2632 2743
rect 2626 2738 2632 2739
rect 2660 2732 2662 2770
rect 2720 2752 2722 2846
rect 2766 2841 2772 2842
rect 2766 2837 2767 2841
rect 2771 2837 2772 2841
rect 2766 2836 2772 2837
rect 2990 2841 2996 2842
rect 2990 2837 2991 2841
rect 2995 2837 2996 2841
rect 2990 2836 2996 2837
rect 3214 2841 3220 2842
rect 3214 2837 3215 2841
rect 3219 2837 3220 2841
rect 3214 2836 3220 2837
rect 3430 2841 3436 2842
rect 3430 2837 3431 2841
rect 3435 2837 3436 2841
rect 3430 2836 3436 2837
rect 2768 2811 2770 2836
rect 2992 2811 2994 2836
rect 3216 2811 3218 2836
rect 3432 2811 3434 2836
rect 2735 2810 2739 2811
rect 2735 2805 2739 2806
rect 2767 2810 2771 2811
rect 2767 2805 2771 2806
rect 2927 2810 2931 2811
rect 2927 2805 2931 2806
rect 2991 2810 2995 2811
rect 2991 2805 2995 2806
rect 3111 2810 3115 2811
rect 3111 2805 3115 2806
rect 3215 2810 3219 2811
rect 3215 2805 3219 2806
rect 3295 2810 3299 2811
rect 3295 2805 3299 2806
rect 3431 2810 3435 2811
rect 3431 2805 3435 2806
rect 2736 2784 2738 2805
rect 2928 2784 2930 2805
rect 3112 2784 3114 2805
rect 3296 2784 3298 2805
rect 2734 2783 2740 2784
rect 2734 2779 2735 2783
rect 2739 2779 2740 2783
rect 2734 2778 2740 2779
rect 2926 2783 2932 2784
rect 2926 2779 2927 2783
rect 2931 2779 2932 2783
rect 2926 2778 2932 2779
rect 3110 2783 3116 2784
rect 3110 2779 3111 2783
rect 3115 2779 3116 2783
rect 3110 2778 3116 2779
rect 3294 2783 3300 2784
rect 3294 2779 3295 2783
rect 3299 2779 3300 2783
rect 3294 2778 3300 2779
rect 3440 2776 3442 2870
rect 3508 2852 3510 2878
rect 3620 2852 3622 2902
rect 3648 2891 3650 2915
rect 3724 2900 3726 2922
rect 3838 2920 3844 2921
rect 3838 2916 3839 2920
rect 3843 2916 3844 2920
rect 3838 2915 3844 2916
rect 3722 2899 3728 2900
rect 3722 2895 3723 2899
rect 3727 2895 3728 2899
rect 3722 2894 3728 2895
rect 3840 2891 3842 2915
rect 3647 2890 3651 2891
rect 3647 2885 3651 2886
rect 3839 2890 3843 2891
rect 3839 2885 3843 2886
rect 3648 2861 3650 2885
rect 3840 2861 3842 2885
rect 3646 2860 3652 2861
rect 3646 2856 3647 2860
rect 3651 2856 3652 2860
rect 3646 2855 3652 2856
rect 3838 2860 3844 2861
rect 3838 2856 3839 2860
rect 3843 2856 3844 2860
rect 3838 2855 3844 2856
rect 3506 2851 3512 2852
rect 3506 2847 3507 2851
rect 3511 2847 3512 2851
rect 3506 2846 3512 2847
rect 3618 2851 3624 2852
rect 3618 2847 3619 2851
rect 3623 2847 3624 2851
rect 3618 2846 3624 2847
rect 3646 2841 3652 2842
rect 3646 2837 3647 2841
rect 3651 2837 3652 2841
rect 3646 2836 3652 2837
rect 3838 2841 3844 2842
rect 3838 2837 3839 2841
rect 3843 2837 3844 2841
rect 3838 2836 3844 2837
rect 3648 2811 3650 2836
rect 3840 2811 3842 2836
rect 3479 2810 3483 2811
rect 3479 2805 3483 2806
rect 3647 2810 3651 2811
rect 3647 2805 3651 2806
rect 3671 2810 3675 2811
rect 3671 2805 3675 2806
rect 3839 2810 3843 2811
rect 3839 2805 3843 2806
rect 3480 2784 3482 2805
rect 3672 2784 3674 2805
rect 3840 2784 3842 2805
rect 3478 2783 3484 2784
rect 3478 2779 3479 2783
rect 3483 2779 3484 2783
rect 3478 2778 3484 2779
rect 3670 2783 3676 2784
rect 3670 2779 3671 2783
rect 3675 2779 3676 2783
rect 3670 2778 3676 2779
rect 3838 2783 3844 2784
rect 3838 2779 3839 2783
rect 3843 2779 3844 2783
rect 3838 2778 3844 2779
rect 3438 2775 3444 2776
rect 3002 2771 3008 2772
rect 3002 2767 3003 2771
rect 3007 2767 3008 2771
rect 3002 2766 3008 2767
rect 3186 2771 3192 2772
rect 3186 2767 3187 2771
rect 3191 2767 3192 2771
rect 3186 2766 3192 2767
rect 3370 2771 3376 2772
rect 3370 2767 3371 2771
rect 3375 2767 3376 2771
rect 3438 2771 3439 2775
rect 3443 2771 3444 2775
rect 3438 2770 3444 2771
rect 3746 2771 3752 2772
rect 3370 2766 3376 2767
rect 3746 2767 3747 2771
rect 3751 2767 3752 2771
rect 3746 2766 3752 2767
rect 2734 2764 2740 2765
rect 2734 2760 2735 2764
rect 2739 2760 2740 2764
rect 2734 2759 2740 2760
rect 2926 2764 2932 2765
rect 2926 2760 2927 2764
rect 2931 2760 2932 2764
rect 2926 2759 2932 2760
rect 2718 2751 2724 2752
rect 2718 2747 2719 2751
rect 2723 2747 2724 2751
rect 2718 2746 2724 2747
rect 2658 2731 2664 2732
rect 2736 2731 2738 2759
rect 2928 2731 2930 2759
rect 3004 2744 3006 2766
rect 3110 2764 3116 2765
rect 3110 2760 3111 2764
rect 3115 2760 3116 2764
rect 3110 2759 3116 2760
rect 3002 2743 3008 2744
rect 3002 2739 3003 2743
rect 3007 2739 3008 2743
rect 3002 2738 3008 2739
rect 3112 2731 3114 2759
rect 3188 2744 3190 2766
rect 3294 2764 3300 2765
rect 3294 2760 3295 2764
rect 3299 2760 3300 2764
rect 3294 2759 3300 2760
rect 3186 2743 3192 2744
rect 3186 2739 3187 2743
rect 3191 2739 3192 2743
rect 3186 2738 3192 2739
rect 3296 2731 3298 2759
rect 3372 2744 3374 2766
rect 3478 2764 3484 2765
rect 3478 2760 3479 2764
rect 3483 2760 3484 2764
rect 3478 2759 3484 2760
rect 3670 2764 3676 2765
rect 3670 2760 3671 2764
rect 3675 2760 3676 2764
rect 3670 2759 3676 2760
rect 3370 2743 3376 2744
rect 3370 2739 3371 2743
rect 3375 2739 3376 2743
rect 3370 2738 3376 2739
rect 3378 2735 3384 2736
rect 3378 2731 3379 2735
rect 3383 2731 3384 2735
rect 3480 2731 3482 2759
rect 3672 2731 3674 2759
rect 2047 2730 2051 2731
rect 2047 2725 2051 2726
rect 2071 2730 2075 2731
rect 2071 2725 2075 2726
rect 2191 2730 2195 2731
rect 2191 2725 2195 2726
rect 2199 2730 2203 2731
rect 2199 2725 2203 2726
rect 2319 2730 2323 2731
rect 2319 2725 2323 2726
rect 2367 2730 2371 2731
rect 2367 2725 2371 2726
rect 2447 2730 2451 2731
rect 2447 2725 2451 2726
rect 2551 2730 2555 2731
rect 2551 2725 2555 2726
rect 2583 2730 2587 2731
rect 2658 2727 2659 2731
rect 2663 2727 2664 2731
rect 2658 2726 2664 2727
rect 2727 2730 2731 2731
rect 2583 2725 2587 2726
rect 2727 2725 2731 2726
rect 2735 2730 2739 2731
rect 2735 2725 2739 2726
rect 2887 2730 2891 2731
rect 2887 2725 2891 2726
rect 2927 2730 2931 2731
rect 2927 2725 2931 2726
rect 3063 2730 3067 2731
rect 3063 2725 3067 2726
rect 3111 2730 3115 2731
rect 3111 2725 3115 2726
rect 3255 2730 3259 2731
rect 3255 2725 3259 2726
rect 3295 2730 3299 2731
rect 3378 2730 3384 2731
rect 3455 2730 3459 2731
rect 3295 2725 3299 2726
rect 2006 2716 2012 2717
rect 2006 2712 2007 2716
rect 2011 2712 2012 2716
rect 2006 2711 2012 2712
rect 1858 2707 1864 2708
rect 1234 2703 1240 2704
rect 1234 2699 1235 2703
rect 1239 2699 1240 2703
rect 1234 2698 1240 2699
rect 1386 2703 1392 2704
rect 1386 2699 1387 2703
rect 1391 2699 1392 2703
rect 1386 2698 1392 2699
rect 1538 2703 1544 2704
rect 1538 2699 1539 2703
rect 1543 2699 1544 2703
rect 1538 2698 1544 2699
rect 1698 2703 1704 2704
rect 1698 2699 1699 2703
rect 1703 2699 1704 2703
rect 1858 2703 1859 2707
rect 1863 2703 1864 2707
rect 1858 2702 1864 2703
rect 1698 2698 1704 2699
rect 2006 2699 2012 2700
rect 1158 2696 1164 2697
rect 1158 2692 1159 2696
rect 1163 2692 1164 2696
rect 1158 2691 1164 2692
rect 1150 2675 1156 2676
rect 1150 2671 1151 2675
rect 1155 2671 1156 2675
rect 1150 2670 1156 2671
rect 1160 2663 1162 2691
rect 1236 2676 1238 2698
rect 1310 2696 1316 2697
rect 1310 2692 1311 2696
rect 1315 2692 1316 2696
rect 1310 2691 1316 2692
rect 1234 2675 1240 2676
rect 1234 2671 1235 2675
rect 1239 2671 1240 2675
rect 1234 2670 1240 2671
rect 1312 2663 1314 2691
rect 111 2662 115 2663
rect 111 2657 115 2658
rect 367 2662 371 2663
rect 367 2657 371 2658
rect 487 2662 491 2663
rect 487 2657 491 2658
rect 511 2662 515 2663
rect 511 2657 515 2658
rect 615 2662 619 2663
rect 615 2657 619 2658
rect 623 2662 627 2663
rect 623 2657 627 2658
rect 743 2662 747 2663
rect 743 2657 747 2658
rect 751 2662 755 2663
rect 858 2662 864 2663
rect 879 2662 883 2663
rect 751 2657 755 2658
rect 112 2630 114 2657
rect 368 2633 370 2657
rect 442 2655 448 2656
rect 442 2651 443 2655
rect 447 2651 448 2655
rect 442 2650 448 2651
rect 366 2632 372 2633
rect 110 2629 116 2630
rect 110 2625 111 2629
rect 115 2625 116 2629
rect 366 2628 367 2632
rect 371 2628 372 2632
rect 366 2627 372 2628
rect 110 2624 116 2625
rect 444 2624 446 2650
rect 488 2633 490 2657
rect 562 2655 568 2656
rect 562 2651 563 2655
rect 567 2651 568 2655
rect 562 2650 568 2651
rect 486 2632 492 2633
rect 486 2628 487 2632
rect 491 2628 492 2632
rect 486 2627 492 2628
rect 564 2624 566 2650
rect 616 2633 618 2657
rect 690 2655 696 2656
rect 690 2651 691 2655
rect 695 2651 696 2655
rect 690 2650 696 2651
rect 614 2632 620 2633
rect 614 2628 615 2632
rect 619 2628 620 2632
rect 614 2627 620 2628
rect 692 2624 694 2650
rect 738 2647 744 2648
rect 738 2643 739 2647
rect 743 2643 744 2647
rect 738 2642 744 2643
rect 442 2623 448 2624
rect 442 2619 443 2623
rect 447 2619 448 2623
rect 442 2618 448 2619
rect 562 2623 568 2624
rect 562 2619 563 2623
rect 567 2619 568 2623
rect 562 2618 568 2619
rect 690 2623 696 2624
rect 690 2619 691 2623
rect 695 2619 696 2623
rect 690 2618 696 2619
rect 366 2613 372 2614
rect 110 2612 116 2613
rect 110 2608 111 2612
rect 115 2608 116 2612
rect 366 2609 367 2613
rect 371 2609 372 2613
rect 366 2608 372 2609
rect 486 2613 492 2614
rect 486 2609 487 2613
rect 491 2609 492 2613
rect 486 2608 492 2609
rect 614 2613 620 2614
rect 614 2609 615 2613
rect 619 2609 620 2613
rect 614 2608 620 2609
rect 110 2607 116 2608
rect 112 2587 114 2607
rect 368 2587 370 2608
rect 488 2587 490 2608
rect 616 2587 618 2608
rect 111 2586 115 2587
rect 111 2581 115 2582
rect 135 2586 139 2587
rect 135 2581 139 2582
rect 287 2586 291 2587
rect 287 2581 291 2582
rect 367 2586 371 2587
rect 367 2581 371 2582
rect 447 2586 451 2587
rect 447 2581 451 2582
rect 487 2586 491 2587
rect 487 2581 491 2582
rect 607 2586 611 2587
rect 607 2581 611 2582
rect 615 2586 619 2587
rect 615 2581 619 2582
rect 112 2561 114 2581
rect 110 2560 116 2561
rect 136 2560 138 2581
rect 288 2560 290 2581
rect 448 2560 450 2581
rect 608 2560 610 2581
rect 110 2556 111 2560
rect 115 2556 116 2560
rect 110 2555 116 2556
rect 134 2559 140 2560
rect 134 2555 135 2559
rect 139 2555 140 2559
rect 134 2554 140 2555
rect 286 2559 292 2560
rect 286 2555 287 2559
rect 291 2555 292 2559
rect 286 2554 292 2555
rect 446 2559 452 2560
rect 446 2555 447 2559
rect 451 2555 452 2559
rect 446 2554 452 2555
rect 606 2559 612 2560
rect 606 2555 607 2559
rect 611 2555 612 2559
rect 606 2554 612 2555
rect 740 2552 742 2642
rect 752 2633 754 2657
rect 826 2655 832 2656
rect 826 2651 827 2655
rect 831 2651 832 2655
rect 826 2650 832 2651
rect 750 2632 756 2633
rect 750 2628 751 2632
rect 755 2628 756 2632
rect 750 2627 756 2628
rect 828 2624 830 2650
rect 860 2624 862 2662
rect 879 2657 883 2658
rect 895 2662 899 2663
rect 895 2657 899 2658
rect 1015 2662 1019 2663
rect 1015 2657 1019 2658
rect 1031 2662 1035 2663
rect 1031 2657 1035 2658
rect 1159 2662 1163 2663
rect 1159 2657 1163 2658
rect 1167 2662 1171 2663
rect 1167 2657 1171 2658
rect 1303 2662 1307 2663
rect 1303 2657 1307 2658
rect 1311 2662 1315 2663
rect 1311 2657 1315 2658
rect 896 2633 898 2657
rect 1032 2633 1034 2657
rect 1168 2633 1170 2657
rect 1250 2655 1256 2656
rect 1250 2651 1251 2655
rect 1255 2651 1256 2655
rect 1250 2650 1256 2651
rect 894 2632 900 2633
rect 894 2628 895 2632
rect 899 2628 900 2632
rect 894 2627 900 2628
rect 1030 2632 1036 2633
rect 1030 2628 1031 2632
rect 1035 2628 1036 2632
rect 1030 2627 1036 2628
rect 1166 2632 1172 2633
rect 1166 2628 1167 2632
rect 1171 2628 1172 2632
rect 1166 2627 1172 2628
rect 1252 2624 1254 2650
rect 1304 2633 1306 2657
rect 1388 2656 1390 2698
rect 1462 2696 1468 2697
rect 1462 2692 1463 2696
rect 1467 2692 1468 2696
rect 1462 2691 1468 2692
rect 1464 2663 1466 2691
rect 1540 2676 1542 2698
rect 1622 2696 1628 2697
rect 1622 2692 1623 2696
rect 1627 2692 1628 2696
rect 1622 2691 1628 2692
rect 1538 2675 1544 2676
rect 1506 2671 1512 2672
rect 1506 2667 1507 2671
rect 1511 2667 1512 2671
rect 1538 2671 1539 2675
rect 1543 2671 1544 2675
rect 1538 2670 1544 2671
rect 1506 2666 1512 2667
rect 1431 2662 1435 2663
rect 1431 2657 1435 2658
rect 1463 2662 1467 2663
rect 1463 2657 1467 2658
rect 1386 2655 1392 2656
rect 1386 2651 1387 2655
rect 1391 2651 1392 2655
rect 1386 2650 1392 2651
rect 1432 2633 1434 2657
rect 1302 2632 1308 2633
rect 1302 2628 1303 2632
rect 1307 2628 1308 2632
rect 1302 2627 1308 2628
rect 1430 2632 1436 2633
rect 1430 2628 1431 2632
rect 1435 2628 1436 2632
rect 1430 2627 1436 2628
rect 1508 2624 1510 2666
rect 1624 2663 1626 2691
rect 1700 2676 1702 2698
rect 1782 2696 1788 2697
rect 1782 2692 1783 2696
rect 1787 2692 1788 2696
rect 2006 2695 2007 2699
rect 2011 2695 2012 2699
rect 2048 2698 2050 2725
rect 2072 2701 2074 2725
rect 2146 2723 2152 2724
rect 2146 2719 2147 2723
rect 2151 2719 2152 2723
rect 2146 2718 2152 2719
rect 2070 2700 2076 2701
rect 2006 2694 2012 2695
rect 2046 2697 2052 2698
rect 1782 2691 1788 2692
rect 1698 2675 1704 2676
rect 1698 2671 1699 2675
rect 1703 2671 1704 2675
rect 1698 2670 1704 2671
rect 1784 2663 1786 2691
rect 2008 2663 2010 2694
rect 2046 2693 2047 2697
rect 2051 2693 2052 2697
rect 2070 2696 2071 2700
rect 2075 2696 2076 2700
rect 2070 2695 2076 2696
rect 2046 2692 2052 2693
rect 2148 2692 2150 2718
rect 2192 2701 2194 2725
rect 2266 2723 2272 2724
rect 2266 2719 2267 2723
rect 2271 2719 2272 2723
rect 2266 2718 2272 2719
rect 2190 2700 2196 2701
rect 2190 2696 2191 2700
rect 2195 2696 2196 2700
rect 2190 2695 2196 2696
rect 2268 2692 2270 2718
rect 2320 2701 2322 2725
rect 2394 2723 2400 2724
rect 2394 2719 2395 2723
rect 2399 2719 2400 2723
rect 2394 2718 2400 2719
rect 2318 2700 2324 2701
rect 2318 2696 2319 2700
rect 2323 2696 2324 2700
rect 2318 2695 2324 2696
rect 2396 2692 2398 2718
rect 2448 2701 2450 2725
rect 2522 2723 2528 2724
rect 2522 2719 2523 2723
rect 2527 2719 2528 2723
rect 2522 2718 2528 2719
rect 2446 2700 2452 2701
rect 2446 2696 2447 2700
rect 2451 2696 2452 2700
rect 2446 2695 2452 2696
rect 2524 2692 2526 2718
rect 2584 2701 2586 2725
rect 2728 2701 2730 2725
rect 2782 2723 2788 2724
rect 2782 2719 2783 2723
rect 2787 2719 2788 2723
rect 2782 2718 2788 2719
rect 2802 2723 2808 2724
rect 2802 2719 2803 2723
rect 2807 2719 2808 2723
rect 2802 2718 2808 2719
rect 2582 2700 2588 2701
rect 2582 2696 2583 2700
rect 2587 2696 2588 2700
rect 2582 2695 2588 2696
rect 2726 2700 2732 2701
rect 2726 2696 2727 2700
rect 2731 2696 2732 2700
rect 2726 2695 2732 2696
rect 2146 2691 2152 2692
rect 2146 2687 2147 2691
rect 2151 2687 2152 2691
rect 2146 2686 2152 2687
rect 2266 2691 2272 2692
rect 2266 2687 2267 2691
rect 2271 2687 2272 2691
rect 2266 2686 2272 2687
rect 2394 2691 2400 2692
rect 2394 2687 2395 2691
rect 2399 2687 2400 2691
rect 2394 2686 2400 2687
rect 2522 2691 2528 2692
rect 2522 2687 2523 2691
rect 2527 2687 2528 2691
rect 2522 2686 2528 2687
rect 2538 2691 2544 2692
rect 2538 2687 2539 2691
rect 2543 2687 2544 2691
rect 2538 2686 2544 2687
rect 2070 2681 2076 2682
rect 2046 2680 2052 2681
rect 2046 2676 2047 2680
rect 2051 2676 2052 2680
rect 2070 2677 2071 2681
rect 2075 2677 2076 2681
rect 2070 2676 2076 2677
rect 2190 2681 2196 2682
rect 2190 2677 2191 2681
rect 2195 2677 2196 2681
rect 2190 2676 2196 2677
rect 2318 2681 2324 2682
rect 2318 2677 2319 2681
rect 2323 2677 2324 2681
rect 2318 2676 2324 2677
rect 2446 2681 2452 2682
rect 2446 2677 2447 2681
rect 2451 2677 2452 2681
rect 2446 2676 2452 2677
rect 2046 2675 2052 2676
rect 1567 2662 1571 2663
rect 1567 2657 1571 2658
rect 1623 2662 1627 2663
rect 1623 2657 1627 2658
rect 1703 2662 1707 2663
rect 1703 2657 1707 2658
rect 1783 2662 1787 2663
rect 1783 2657 1787 2658
rect 2007 2662 2011 2663
rect 2007 2657 2011 2658
rect 1514 2655 1520 2656
rect 1514 2651 1515 2655
rect 1519 2651 1520 2655
rect 1514 2650 1520 2651
rect 1516 2624 1518 2650
rect 1568 2633 1570 2657
rect 1650 2655 1656 2656
rect 1650 2651 1651 2655
rect 1655 2651 1656 2655
rect 1650 2650 1656 2651
rect 1566 2632 1572 2633
rect 1566 2628 1567 2632
rect 1571 2628 1572 2632
rect 1566 2627 1572 2628
rect 1652 2624 1654 2650
rect 1704 2633 1706 2657
rect 1802 2655 1808 2656
rect 1802 2651 1803 2655
rect 1807 2651 1808 2655
rect 1802 2650 1808 2651
rect 1702 2632 1708 2633
rect 1702 2628 1703 2632
rect 1707 2628 1708 2632
rect 1702 2627 1708 2628
rect 826 2623 832 2624
rect 826 2619 827 2623
rect 831 2619 832 2623
rect 826 2618 832 2619
rect 858 2623 864 2624
rect 858 2619 859 2623
rect 863 2619 864 2623
rect 858 2618 864 2619
rect 978 2623 984 2624
rect 978 2619 979 2623
rect 983 2619 984 2623
rect 978 2618 984 2619
rect 1250 2623 1256 2624
rect 1250 2619 1251 2623
rect 1255 2619 1256 2623
rect 1250 2618 1256 2619
rect 1506 2623 1512 2624
rect 1506 2619 1507 2623
rect 1511 2619 1512 2623
rect 1506 2618 1512 2619
rect 1514 2623 1520 2624
rect 1514 2619 1515 2623
rect 1519 2619 1520 2623
rect 1514 2618 1520 2619
rect 1650 2623 1656 2624
rect 1650 2619 1651 2623
rect 1655 2619 1656 2623
rect 1650 2618 1656 2619
rect 750 2613 756 2614
rect 750 2609 751 2613
rect 755 2609 756 2613
rect 750 2608 756 2609
rect 894 2613 900 2614
rect 894 2609 895 2613
rect 899 2609 900 2613
rect 894 2608 900 2609
rect 752 2587 754 2608
rect 896 2587 898 2608
rect 751 2586 755 2587
rect 751 2581 755 2582
rect 767 2586 771 2587
rect 767 2581 771 2582
rect 895 2586 899 2587
rect 895 2581 899 2582
rect 919 2586 923 2587
rect 919 2581 923 2582
rect 768 2560 770 2581
rect 920 2560 922 2581
rect 766 2559 772 2560
rect 766 2555 767 2559
rect 771 2555 772 2559
rect 766 2554 772 2555
rect 918 2559 924 2560
rect 918 2555 919 2559
rect 923 2555 924 2559
rect 918 2554 924 2555
rect 738 2551 744 2552
rect 210 2547 216 2548
rect 110 2543 116 2544
rect 110 2539 111 2543
rect 115 2539 116 2543
rect 210 2543 211 2547
rect 215 2543 216 2547
rect 210 2542 216 2543
rect 362 2547 368 2548
rect 362 2543 363 2547
rect 367 2543 368 2547
rect 362 2542 368 2543
rect 522 2547 528 2548
rect 522 2543 523 2547
rect 527 2543 528 2547
rect 522 2542 528 2543
rect 682 2547 688 2548
rect 682 2543 683 2547
rect 687 2543 688 2547
rect 738 2547 739 2551
rect 743 2547 744 2551
rect 738 2546 744 2547
rect 682 2542 688 2543
rect 110 2538 116 2539
rect 134 2540 140 2541
rect 112 2495 114 2538
rect 134 2536 135 2540
rect 139 2536 140 2540
rect 134 2535 140 2536
rect 136 2495 138 2535
rect 212 2524 214 2542
rect 286 2540 292 2541
rect 286 2536 287 2540
rect 291 2536 292 2540
rect 286 2535 292 2536
rect 210 2523 216 2524
rect 210 2519 211 2523
rect 215 2519 216 2523
rect 210 2518 216 2519
rect 288 2495 290 2535
rect 364 2520 366 2542
rect 446 2540 452 2541
rect 446 2536 447 2540
rect 451 2536 452 2540
rect 446 2535 452 2536
rect 362 2519 368 2520
rect 362 2515 363 2519
rect 367 2515 368 2519
rect 362 2514 368 2515
rect 448 2495 450 2535
rect 524 2520 526 2542
rect 606 2540 612 2541
rect 606 2536 607 2540
rect 611 2536 612 2540
rect 606 2535 612 2536
rect 522 2519 528 2520
rect 522 2515 523 2519
rect 527 2515 528 2519
rect 522 2514 528 2515
rect 506 2511 512 2512
rect 506 2507 507 2511
rect 511 2507 512 2511
rect 506 2506 512 2507
rect 111 2494 115 2495
rect 111 2489 115 2490
rect 135 2494 139 2495
rect 135 2489 139 2490
rect 231 2494 235 2495
rect 231 2489 235 2490
rect 287 2494 291 2495
rect 287 2489 291 2490
rect 327 2494 331 2495
rect 327 2489 331 2490
rect 423 2494 427 2495
rect 423 2489 427 2490
rect 447 2494 451 2495
rect 447 2489 451 2490
rect 112 2462 114 2489
rect 136 2465 138 2489
rect 202 2487 208 2488
rect 202 2483 203 2487
rect 207 2483 208 2487
rect 202 2482 208 2483
rect 210 2487 216 2488
rect 210 2483 211 2487
rect 215 2483 216 2487
rect 210 2482 216 2483
rect 134 2464 140 2465
rect 110 2461 116 2462
rect 110 2457 111 2461
rect 115 2457 116 2461
rect 134 2460 135 2464
rect 139 2460 140 2464
rect 134 2459 140 2460
rect 110 2456 116 2457
rect 134 2445 140 2446
rect 110 2444 116 2445
rect 110 2440 111 2444
rect 115 2440 116 2444
rect 134 2441 135 2445
rect 139 2441 140 2445
rect 134 2440 140 2441
rect 110 2439 116 2440
rect 112 2403 114 2439
rect 136 2403 138 2440
rect 111 2402 115 2403
rect 111 2397 115 2398
rect 135 2402 139 2403
rect 135 2397 139 2398
rect 112 2377 114 2397
rect 110 2376 116 2377
rect 136 2376 138 2397
rect 110 2372 111 2376
rect 115 2372 116 2376
rect 110 2371 116 2372
rect 134 2375 140 2376
rect 134 2371 135 2375
rect 139 2371 140 2375
rect 204 2372 206 2482
rect 212 2456 214 2482
rect 232 2465 234 2489
rect 306 2487 312 2488
rect 306 2483 307 2487
rect 311 2483 312 2487
rect 306 2482 312 2483
rect 230 2464 236 2465
rect 230 2460 231 2464
rect 235 2460 236 2464
rect 230 2459 236 2460
rect 308 2456 310 2482
rect 328 2465 330 2489
rect 402 2487 408 2488
rect 402 2483 403 2487
rect 407 2483 408 2487
rect 402 2482 408 2483
rect 326 2464 332 2465
rect 326 2460 327 2464
rect 331 2460 332 2464
rect 326 2459 332 2460
rect 404 2456 406 2482
rect 424 2465 426 2489
rect 498 2487 504 2488
rect 498 2483 499 2487
rect 503 2483 504 2487
rect 498 2482 504 2483
rect 422 2464 428 2465
rect 422 2460 423 2464
rect 427 2460 428 2464
rect 422 2459 428 2460
rect 500 2456 502 2482
rect 508 2456 510 2506
rect 608 2495 610 2535
rect 684 2520 686 2542
rect 766 2540 772 2541
rect 766 2536 767 2540
rect 771 2536 772 2540
rect 766 2535 772 2536
rect 918 2540 924 2541
rect 918 2536 919 2540
rect 923 2536 924 2540
rect 918 2535 924 2536
rect 682 2519 688 2520
rect 682 2515 683 2519
rect 687 2515 688 2519
rect 682 2514 688 2515
rect 768 2495 770 2535
rect 920 2495 922 2535
rect 980 2531 982 2618
rect 1030 2613 1036 2614
rect 1030 2609 1031 2613
rect 1035 2609 1036 2613
rect 1030 2608 1036 2609
rect 1166 2613 1172 2614
rect 1166 2609 1167 2613
rect 1171 2609 1172 2613
rect 1166 2608 1172 2609
rect 1302 2613 1308 2614
rect 1302 2609 1303 2613
rect 1307 2609 1308 2613
rect 1302 2608 1308 2609
rect 1430 2613 1436 2614
rect 1430 2609 1431 2613
rect 1435 2609 1436 2613
rect 1430 2608 1436 2609
rect 1566 2613 1572 2614
rect 1566 2609 1567 2613
rect 1571 2609 1572 2613
rect 1566 2608 1572 2609
rect 1702 2613 1708 2614
rect 1702 2609 1703 2613
rect 1707 2609 1708 2613
rect 1702 2608 1708 2609
rect 1032 2587 1034 2608
rect 1168 2587 1170 2608
rect 1304 2587 1306 2608
rect 1432 2587 1434 2608
rect 1568 2587 1570 2608
rect 1704 2587 1706 2608
rect 1031 2586 1035 2587
rect 1031 2581 1035 2582
rect 1063 2586 1067 2587
rect 1063 2581 1067 2582
rect 1167 2586 1171 2587
rect 1167 2581 1171 2582
rect 1199 2586 1203 2587
rect 1199 2581 1203 2582
rect 1303 2586 1307 2587
rect 1303 2581 1307 2582
rect 1335 2586 1339 2587
rect 1335 2581 1339 2582
rect 1431 2586 1435 2587
rect 1431 2581 1435 2582
rect 1463 2586 1467 2587
rect 1463 2581 1467 2582
rect 1567 2586 1571 2587
rect 1567 2581 1571 2582
rect 1591 2586 1595 2587
rect 1591 2581 1595 2582
rect 1703 2586 1707 2587
rect 1703 2581 1707 2582
rect 1727 2586 1731 2587
rect 1727 2581 1731 2582
rect 1064 2560 1066 2581
rect 1200 2560 1202 2581
rect 1336 2560 1338 2581
rect 1464 2560 1466 2581
rect 1592 2560 1594 2581
rect 1728 2560 1730 2581
rect 1062 2559 1068 2560
rect 1062 2555 1063 2559
rect 1067 2555 1068 2559
rect 1062 2554 1068 2555
rect 1198 2559 1204 2560
rect 1198 2555 1199 2559
rect 1203 2555 1204 2559
rect 1198 2554 1204 2555
rect 1334 2559 1340 2560
rect 1334 2555 1335 2559
rect 1339 2555 1340 2559
rect 1334 2554 1340 2555
rect 1462 2559 1468 2560
rect 1462 2555 1463 2559
rect 1467 2555 1468 2559
rect 1462 2554 1468 2555
rect 1590 2559 1596 2560
rect 1590 2555 1591 2559
rect 1595 2555 1596 2559
rect 1590 2554 1596 2555
rect 1726 2559 1732 2560
rect 1726 2555 1727 2559
rect 1731 2555 1732 2559
rect 1726 2554 1732 2555
rect 1804 2552 1806 2650
rect 2008 2630 2010 2657
rect 2048 2647 2050 2675
rect 2072 2647 2074 2676
rect 2192 2647 2194 2676
rect 2320 2647 2322 2676
rect 2448 2647 2450 2676
rect 2047 2646 2051 2647
rect 2047 2641 2051 2642
rect 2071 2646 2075 2647
rect 2071 2641 2075 2642
rect 2191 2646 2195 2647
rect 2191 2641 2195 2642
rect 2231 2646 2235 2647
rect 2231 2641 2235 2642
rect 2319 2646 2323 2647
rect 2319 2641 2323 2642
rect 2335 2646 2339 2647
rect 2335 2641 2339 2642
rect 2447 2646 2451 2647
rect 2447 2641 2451 2642
rect 2006 2629 2012 2630
rect 2006 2625 2007 2629
rect 2011 2625 2012 2629
rect 2006 2624 2012 2625
rect 2048 2621 2050 2641
rect 2046 2620 2052 2621
rect 2232 2620 2234 2641
rect 2336 2620 2338 2641
rect 2448 2620 2450 2641
rect 2046 2616 2047 2620
rect 2051 2616 2052 2620
rect 2046 2615 2052 2616
rect 2230 2619 2236 2620
rect 2230 2615 2231 2619
rect 2235 2615 2236 2619
rect 2230 2614 2236 2615
rect 2334 2619 2340 2620
rect 2334 2615 2335 2619
rect 2339 2615 2340 2619
rect 2334 2614 2340 2615
rect 2446 2619 2452 2620
rect 2446 2615 2447 2619
rect 2451 2615 2452 2619
rect 2446 2614 2452 2615
rect 2006 2612 2012 2613
rect 2006 2608 2007 2612
rect 2011 2608 2012 2612
rect 2006 2607 2012 2608
rect 2306 2607 2312 2608
rect 2008 2587 2010 2607
rect 2046 2603 2052 2604
rect 2046 2599 2047 2603
rect 2051 2599 2052 2603
rect 2306 2603 2307 2607
rect 2311 2603 2312 2607
rect 2306 2602 2312 2603
rect 2410 2607 2416 2608
rect 2410 2603 2411 2607
rect 2415 2603 2416 2607
rect 2410 2602 2416 2603
rect 2522 2607 2528 2608
rect 2522 2603 2523 2607
rect 2527 2603 2528 2607
rect 2522 2602 2528 2603
rect 2046 2598 2052 2599
rect 2230 2600 2236 2601
rect 2007 2586 2011 2587
rect 2007 2581 2011 2582
rect 2008 2561 2010 2581
rect 2048 2567 2050 2598
rect 2230 2596 2231 2600
rect 2235 2596 2236 2600
rect 2230 2595 2236 2596
rect 2232 2567 2234 2595
rect 2308 2580 2310 2602
rect 2334 2600 2340 2601
rect 2334 2596 2335 2600
rect 2339 2596 2340 2600
rect 2334 2595 2340 2596
rect 2306 2579 2312 2580
rect 2306 2575 2307 2579
rect 2311 2575 2312 2579
rect 2306 2574 2312 2575
rect 2336 2567 2338 2595
rect 2412 2580 2414 2602
rect 2446 2600 2452 2601
rect 2446 2596 2447 2600
rect 2451 2596 2452 2600
rect 2446 2595 2452 2596
rect 2410 2579 2416 2580
rect 2410 2575 2411 2579
rect 2415 2575 2416 2579
rect 2410 2574 2416 2575
rect 2448 2567 2450 2595
rect 2524 2580 2526 2602
rect 2540 2588 2542 2686
rect 2582 2681 2588 2682
rect 2582 2677 2583 2681
rect 2587 2677 2588 2681
rect 2582 2676 2588 2677
rect 2726 2681 2732 2682
rect 2726 2677 2727 2681
rect 2731 2677 2732 2681
rect 2726 2676 2732 2677
rect 2584 2647 2586 2676
rect 2728 2647 2730 2676
rect 2559 2646 2563 2647
rect 2559 2641 2563 2642
rect 2583 2646 2587 2647
rect 2583 2641 2587 2642
rect 2671 2646 2675 2647
rect 2671 2641 2675 2642
rect 2727 2646 2731 2647
rect 2727 2641 2731 2642
rect 2560 2620 2562 2641
rect 2672 2620 2674 2641
rect 2558 2619 2564 2620
rect 2558 2615 2559 2619
rect 2563 2615 2564 2619
rect 2558 2614 2564 2615
rect 2670 2619 2676 2620
rect 2670 2615 2671 2619
rect 2675 2615 2676 2619
rect 2670 2614 2676 2615
rect 2784 2612 2786 2718
rect 2804 2692 2806 2718
rect 2888 2701 2890 2725
rect 2962 2723 2968 2724
rect 2962 2719 2963 2723
rect 2967 2719 2968 2723
rect 2962 2718 2968 2719
rect 2886 2700 2892 2701
rect 2886 2696 2887 2700
rect 2891 2696 2892 2700
rect 2886 2695 2892 2696
rect 2964 2692 2966 2718
rect 3064 2701 3066 2725
rect 3138 2723 3144 2724
rect 3138 2719 3139 2723
rect 3143 2719 3144 2723
rect 3138 2718 3144 2719
rect 3062 2700 3068 2701
rect 3062 2696 3063 2700
rect 3067 2696 3068 2700
rect 3062 2695 3068 2696
rect 3140 2692 3142 2718
rect 3256 2701 3258 2725
rect 3330 2723 3336 2724
rect 3330 2719 3331 2723
rect 3335 2719 3336 2723
rect 3330 2718 3336 2719
rect 3254 2700 3260 2701
rect 3254 2696 3255 2700
rect 3259 2696 3260 2700
rect 3254 2695 3260 2696
rect 3332 2692 3334 2718
rect 3380 2692 3382 2730
rect 3455 2725 3459 2726
rect 3479 2730 3483 2731
rect 3479 2725 3483 2726
rect 3655 2730 3659 2731
rect 3655 2725 3659 2726
rect 3671 2730 3675 2731
rect 3671 2725 3675 2726
rect 3456 2701 3458 2725
rect 3656 2701 3658 2725
rect 3748 2724 3750 2766
rect 3838 2764 3844 2765
rect 3838 2760 3839 2764
rect 3843 2760 3844 2764
rect 3838 2759 3844 2760
rect 3840 2731 3842 2759
rect 3876 2744 3878 3078
rect 3916 3008 3918 3198
rect 3944 3178 3946 3205
rect 3942 3177 3948 3178
rect 3942 3173 3943 3177
rect 3947 3173 3948 3177
rect 3942 3172 3948 3173
rect 3942 3160 3948 3161
rect 3942 3156 3943 3160
rect 3947 3156 3948 3160
rect 3942 3155 3948 3156
rect 3944 3123 3946 3155
rect 3943 3122 3947 3123
rect 3943 3117 3947 3118
rect 3944 3097 3946 3117
rect 3942 3096 3948 3097
rect 3942 3092 3943 3096
rect 3947 3092 3948 3096
rect 3942 3091 3948 3092
rect 3942 3079 3948 3080
rect 3942 3075 3943 3079
rect 3947 3075 3948 3079
rect 3942 3074 3948 3075
rect 3944 3047 3946 3074
rect 3943 3046 3947 3047
rect 3943 3041 3947 3042
rect 3922 3039 3928 3040
rect 3922 3035 3923 3039
rect 3927 3035 3928 3039
rect 3922 3034 3928 3035
rect 3914 3007 3920 3008
rect 3914 3003 3915 3007
rect 3919 3003 3920 3007
rect 3914 3002 3920 3003
rect 3906 2883 3912 2884
rect 3906 2879 3907 2883
rect 3911 2879 3912 2883
rect 3906 2878 3912 2879
rect 3908 2780 3910 2878
rect 3924 2852 3926 3034
rect 3944 3014 3946 3041
rect 3942 3013 3948 3014
rect 3942 3009 3943 3013
rect 3947 3009 3948 3013
rect 3942 3008 3948 3009
rect 3942 2996 3948 2997
rect 3942 2992 3943 2996
rect 3947 2992 3948 2996
rect 3942 2991 3948 2992
rect 3944 2967 3946 2991
rect 3943 2966 3947 2967
rect 3943 2961 3947 2962
rect 3944 2941 3946 2961
rect 3942 2940 3948 2941
rect 3942 2936 3943 2940
rect 3947 2936 3948 2940
rect 3942 2935 3948 2936
rect 3942 2923 3948 2924
rect 3942 2919 3943 2923
rect 3947 2919 3948 2923
rect 3942 2918 3948 2919
rect 3944 2891 3946 2918
rect 3943 2890 3947 2891
rect 3943 2885 3947 2886
rect 3944 2858 3946 2885
rect 3942 2857 3948 2858
rect 3942 2853 3943 2857
rect 3947 2853 3948 2857
rect 3942 2852 3948 2853
rect 3922 2851 3928 2852
rect 3922 2847 3923 2851
rect 3927 2847 3928 2851
rect 3922 2846 3928 2847
rect 3942 2840 3948 2841
rect 3942 2836 3943 2840
rect 3947 2836 3948 2840
rect 3942 2835 3948 2836
rect 3944 2811 3946 2835
rect 3943 2810 3947 2811
rect 3943 2805 3947 2806
rect 3944 2785 3946 2805
rect 3942 2784 3948 2785
rect 3942 2780 3943 2784
rect 3947 2780 3948 2784
rect 3906 2779 3912 2780
rect 3942 2779 3948 2780
rect 3906 2775 3907 2779
rect 3911 2775 3912 2779
rect 3906 2774 3912 2775
rect 3942 2767 3948 2768
rect 3942 2763 3943 2767
rect 3947 2763 3948 2767
rect 3942 2762 3948 2763
rect 3874 2743 3880 2744
rect 3874 2739 3875 2743
rect 3879 2739 3880 2743
rect 3874 2738 3880 2739
rect 3906 2739 3912 2740
rect 3906 2735 3907 2739
rect 3911 2735 3912 2739
rect 3906 2734 3912 2735
rect 3839 2730 3843 2731
rect 3839 2725 3843 2726
rect 3746 2723 3752 2724
rect 3746 2719 3747 2723
rect 3751 2719 3752 2723
rect 3746 2718 3752 2719
rect 3840 2701 3842 2725
rect 3454 2700 3460 2701
rect 3454 2696 3455 2700
rect 3459 2696 3460 2700
rect 3454 2695 3460 2696
rect 3654 2700 3660 2701
rect 3654 2696 3655 2700
rect 3659 2696 3660 2700
rect 3654 2695 3660 2696
rect 3838 2700 3844 2701
rect 3838 2696 3839 2700
rect 3843 2696 3844 2700
rect 3838 2695 3844 2696
rect 3908 2692 3910 2734
rect 3944 2731 3946 2762
rect 3943 2730 3947 2731
rect 3943 2725 3947 2726
rect 3944 2698 3946 2725
rect 3942 2697 3948 2698
rect 3942 2693 3943 2697
rect 3947 2693 3948 2697
rect 3942 2692 3948 2693
rect 2802 2691 2808 2692
rect 2802 2687 2803 2691
rect 2807 2687 2808 2691
rect 2802 2686 2808 2687
rect 2962 2691 2968 2692
rect 2962 2687 2963 2691
rect 2967 2687 2968 2691
rect 2962 2686 2968 2687
rect 3138 2691 3144 2692
rect 3138 2687 3139 2691
rect 3143 2687 3144 2691
rect 3138 2686 3144 2687
rect 3330 2691 3336 2692
rect 3330 2687 3331 2691
rect 3335 2687 3336 2691
rect 3330 2686 3336 2687
rect 3378 2691 3384 2692
rect 3378 2687 3379 2691
rect 3383 2687 3384 2691
rect 3378 2686 3384 2687
rect 3906 2691 3912 2692
rect 3906 2687 3907 2691
rect 3911 2687 3912 2691
rect 3906 2686 3912 2687
rect 2886 2681 2892 2682
rect 2886 2677 2887 2681
rect 2891 2677 2892 2681
rect 2886 2676 2892 2677
rect 3062 2681 3068 2682
rect 3062 2677 3063 2681
rect 3067 2677 3068 2681
rect 3062 2676 3068 2677
rect 3254 2681 3260 2682
rect 3254 2677 3255 2681
rect 3259 2677 3260 2681
rect 3254 2676 3260 2677
rect 3454 2681 3460 2682
rect 3454 2677 3455 2681
rect 3459 2677 3460 2681
rect 3454 2676 3460 2677
rect 3654 2681 3660 2682
rect 3654 2677 3655 2681
rect 3659 2677 3660 2681
rect 3654 2676 3660 2677
rect 3838 2681 3844 2682
rect 3838 2677 3839 2681
rect 3843 2677 3844 2681
rect 3838 2676 3844 2677
rect 3942 2680 3948 2681
rect 3942 2676 3943 2680
rect 3947 2676 3948 2680
rect 2888 2647 2890 2676
rect 3064 2647 3066 2676
rect 3256 2647 3258 2676
rect 3456 2647 3458 2676
rect 3656 2647 3658 2676
rect 3840 2647 3842 2676
rect 3942 2675 3948 2676
rect 3944 2647 3946 2675
rect 2791 2646 2795 2647
rect 2791 2641 2795 2642
rect 2887 2646 2891 2647
rect 2887 2641 2891 2642
rect 2911 2646 2915 2647
rect 2911 2641 2915 2642
rect 3031 2646 3035 2647
rect 3031 2641 3035 2642
rect 3063 2646 3067 2647
rect 3063 2641 3067 2642
rect 3151 2646 3155 2647
rect 3151 2641 3155 2642
rect 3255 2646 3259 2647
rect 3255 2641 3259 2642
rect 3455 2646 3459 2647
rect 3455 2641 3459 2642
rect 3655 2646 3659 2647
rect 3655 2641 3659 2642
rect 3839 2646 3843 2647
rect 3839 2641 3843 2642
rect 3943 2646 3947 2647
rect 3943 2641 3947 2642
rect 2792 2620 2794 2641
rect 2912 2620 2914 2641
rect 3032 2620 3034 2641
rect 3152 2620 3154 2641
rect 3944 2621 3946 2641
rect 3942 2620 3948 2621
rect 2790 2619 2796 2620
rect 2790 2615 2791 2619
rect 2795 2615 2796 2619
rect 2790 2614 2796 2615
rect 2910 2619 2916 2620
rect 2910 2615 2911 2619
rect 2915 2615 2916 2619
rect 2910 2614 2916 2615
rect 3030 2619 3036 2620
rect 3030 2615 3031 2619
rect 3035 2615 3036 2619
rect 3030 2614 3036 2615
rect 3150 2619 3156 2620
rect 3150 2615 3151 2619
rect 3155 2615 3156 2619
rect 3942 2616 3943 2620
rect 3947 2616 3948 2620
rect 3942 2615 3948 2616
rect 3150 2614 3156 2615
rect 2642 2611 2648 2612
rect 2634 2607 2640 2608
rect 2634 2603 2635 2607
rect 2639 2603 2640 2607
rect 2642 2607 2643 2611
rect 2647 2607 2648 2611
rect 2642 2606 2648 2607
rect 2782 2611 2788 2612
rect 2782 2607 2783 2611
rect 2787 2607 2788 2611
rect 3114 2611 3120 2612
rect 2782 2606 2788 2607
rect 3106 2607 3112 2608
rect 2634 2602 2640 2603
rect 2558 2600 2564 2601
rect 2558 2596 2559 2600
rect 2563 2596 2564 2600
rect 2558 2595 2564 2596
rect 2538 2587 2544 2588
rect 2538 2583 2539 2587
rect 2543 2583 2544 2587
rect 2538 2582 2544 2583
rect 2522 2579 2528 2580
rect 2522 2575 2523 2579
rect 2527 2575 2528 2579
rect 2522 2574 2528 2575
rect 2560 2567 2562 2595
rect 2636 2580 2638 2602
rect 2634 2579 2640 2580
rect 2634 2575 2635 2579
rect 2639 2575 2640 2579
rect 2634 2574 2640 2575
rect 2644 2568 2646 2606
rect 3106 2603 3107 2607
rect 3111 2603 3112 2607
rect 3114 2607 3115 2611
rect 3119 2607 3120 2611
rect 3114 2606 3120 2607
rect 3106 2602 3112 2603
rect 2670 2600 2676 2601
rect 2670 2596 2671 2600
rect 2675 2596 2676 2600
rect 2670 2595 2676 2596
rect 2790 2600 2796 2601
rect 2790 2596 2791 2600
rect 2795 2596 2796 2600
rect 2790 2595 2796 2596
rect 2910 2600 2916 2601
rect 2910 2596 2911 2600
rect 2915 2596 2916 2600
rect 2910 2595 2916 2596
rect 3030 2600 3036 2601
rect 3030 2596 3031 2600
rect 3035 2596 3036 2600
rect 3030 2595 3036 2596
rect 2642 2567 2648 2568
rect 2672 2567 2674 2595
rect 2792 2567 2794 2595
rect 2912 2567 2914 2595
rect 3032 2567 3034 2595
rect 3108 2580 3110 2602
rect 3116 2588 3118 2606
rect 3942 2603 3948 2604
rect 3150 2600 3156 2601
rect 3150 2596 3151 2600
rect 3155 2596 3156 2600
rect 3942 2599 3943 2603
rect 3947 2599 3948 2603
rect 3942 2598 3948 2599
rect 3150 2595 3156 2596
rect 3114 2587 3120 2588
rect 3114 2583 3115 2587
rect 3119 2583 3120 2587
rect 3114 2582 3120 2583
rect 3106 2579 3112 2580
rect 3066 2575 3072 2576
rect 3066 2571 3067 2575
rect 3071 2571 3072 2575
rect 3106 2575 3107 2579
rect 3111 2575 3112 2579
rect 3106 2574 3112 2575
rect 3066 2570 3072 2571
rect 2047 2566 2051 2567
rect 2047 2561 2051 2562
rect 2231 2566 2235 2567
rect 2231 2561 2235 2562
rect 2335 2566 2339 2567
rect 2335 2561 2339 2562
rect 2383 2566 2387 2567
rect 2383 2561 2387 2562
rect 2447 2566 2451 2567
rect 2447 2561 2451 2562
rect 2495 2566 2499 2567
rect 2495 2561 2499 2562
rect 2559 2566 2563 2567
rect 2559 2561 2563 2562
rect 2615 2566 2619 2567
rect 2642 2563 2643 2567
rect 2647 2563 2648 2567
rect 2642 2562 2648 2563
rect 2671 2566 2675 2567
rect 2615 2561 2619 2562
rect 2671 2561 2675 2562
rect 2743 2566 2747 2567
rect 2743 2561 2747 2562
rect 2791 2566 2795 2567
rect 2791 2561 2795 2562
rect 2871 2566 2875 2567
rect 2871 2561 2875 2562
rect 2911 2566 2915 2567
rect 2911 2561 2915 2562
rect 2991 2566 2995 2567
rect 2991 2561 2995 2562
rect 3031 2566 3035 2567
rect 3031 2561 3035 2562
rect 2006 2560 2012 2561
rect 2006 2556 2007 2560
rect 2011 2556 2012 2560
rect 2006 2555 2012 2556
rect 1802 2551 1808 2552
rect 994 2547 1000 2548
rect 994 2543 995 2547
rect 999 2543 1000 2547
rect 994 2542 1000 2543
rect 1138 2547 1144 2548
rect 1138 2543 1139 2547
rect 1143 2543 1144 2547
rect 1138 2542 1144 2543
rect 1274 2547 1280 2548
rect 1274 2543 1275 2547
rect 1279 2543 1280 2547
rect 1274 2542 1280 2543
rect 1410 2547 1416 2548
rect 1410 2543 1411 2547
rect 1415 2543 1416 2547
rect 1410 2542 1416 2543
rect 1538 2547 1544 2548
rect 1538 2543 1539 2547
rect 1543 2543 1544 2547
rect 1538 2542 1544 2543
rect 1666 2547 1672 2548
rect 1666 2543 1667 2547
rect 1671 2543 1672 2547
rect 1802 2547 1803 2551
rect 1807 2547 1808 2551
rect 1802 2546 1808 2547
rect 1666 2542 1672 2543
rect 2006 2543 2012 2544
rect 976 2529 982 2531
rect 976 2520 978 2529
rect 996 2520 998 2542
rect 1062 2540 1068 2541
rect 1062 2536 1063 2540
rect 1067 2536 1068 2540
rect 1062 2535 1068 2536
rect 974 2519 980 2520
rect 974 2515 975 2519
rect 979 2515 980 2519
rect 974 2514 980 2515
rect 994 2519 1000 2520
rect 994 2515 995 2519
rect 999 2515 1000 2519
rect 994 2514 1000 2515
rect 1064 2495 1066 2535
rect 1140 2520 1142 2542
rect 1198 2540 1204 2541
rect 1198 2536 1199 2540
rect 1203 2536 1204 2540
rect 1198 2535 1204 2536
rect 1138 2519 1144 2520
rect 1138 2515 1139 2519
rect 1143 2515 1144 2519
rect 1138 2514 1144 2515
rect 1200 2495 1202 2535
rect 1276 2520 1278 2542
rect 1334 2540 1340 2541
rect 1334 2536 1335 2540
rect 1339 2536 1340 2540
rect 1334 2535 1340 2536
rect 1274 2519 1280 2520
rect 1274 2515 1275 2519
rect 1279 2515 1280 2519
rect 1274 2514 1280 2515
rect 1336 2495 1338 2535
rect 1412 2520 1414 2542
rect 1462 2540 1468 2541
rect 1462 2536 1463 2540
rect 1467 2536 1468 2540
rect 1462 2535 1468 2536
rect 1410 2519 1416 2520
rect 1410 2515 1411 2519
rect 1415 2515 1416 2519
rect 1410 2514 1416 2515
rect 1464 2495 1466 2535
rect 1540 2520 1542 2542
rect 1590 2540 1596 2541
rect 1590 2536 1591 2540
rect 1595 2536 1596 2540
rect 1590 2535 1596 2536
rect 1538 2519 1544 2520
rect 1538 2515 1539 2519
rect 1543 2515 1544 2519
rect 1538 2514 1544 2515
rect 1592 2495 1594 2535
rect 1668 2520 1670 2542
rect 1726 2540 1732 2541
rect 1726 2536 1727 2540
rect 1731 2536 1732 2540
rect 2006 2539 2007 2543
rect 2011 2539 2012 2543
rect 2006 2538 2012 2539
rect 1726 2535 1732 2536
rect 1666 2519 1672 2520
rect 1666 2515 1667 2519
rect 1671 2515 1672 2519
rect 1666 2514 1672 2515
rect 1728 2495 1730 2535
rect 2008 2495 2010 2538
rect 2048 2534 2050 2561
rect 2384 2537 2386 2561
rect 2458 2559 2464 2560
rect 2458 2555 2459 2559
rect 2463 2555 2464 2559
rect 2458 2554 2464 2555
rect 2382 2536 2388 2537
rect 2046 2533 2052 2534
rect 2046 2529 2047 2533
rect 2051 2529 2052 2533
rect 2382 2532 2383 2536
rect 2387 2532 2388 2536
rect 2382 2531 2388 2532
rect 2046 2528 2052 2529
rect 2460 2528 2462 2554
rect 2496 2537 2498 2561
rect 2570 2559 2576 2560
rect 2570 2555 2571 2559
rect 2575 2555 2576 2559
rect 2570 2554 2576 2555
rect 2494 2536 2500 2537
rect 2494 2532 2495 2536
rect 2499 2532 2500 2536
rect 2494 2531 2500 2532
rect 2572 2528 2574 2554
rect 2616 2537 2618 2561
rect 2690 2559 2696 2560
rect 2690 2555 2691 2559
rect 2695 2555 2696 2559
rect 2690 2554 2696 2555
rect 2614 2536 2620 2537
rect 2614 2532 2615 2536
rect 2619 2532 2620 2536
rect 2614 2531 2620 2532
rect 2692 2528 2694 2554
rect 2744 2537 2746 2561
rect 2818 2559 2824 2560
rect 2818 2555 2819 2559
rect 2823 2555 2824 2559
rect 2818 2554 2824 2555
rect 2742 2536 2748 2537
rect 2742 2532 2743 2536
rect 2747 2532 2748 2536
rect 2742 2531 2748 2532
rect 2820 2528 2822 2554
rect 2872 2537 2874 2561
rect 2992 2537 2994 2561
rect 2870 2536 2876 2537
rect 2870 2532 2871 2536
rect 2875 2532 2876 2536
rect 2870 2531 2876 2532
rect 2990 2536 2996 2537
rect 2990 2532 2991 2536
rect 2995 2532 2996 2536
rect 2990 2531 2996 2532
rect 3068 2528 3070 2570
rect 3152 2567 3154 2595
rect 3944 2567 3946 2598
rect 3111 2566 3115 2567
rect 3111 2561 3115 2562
rect 3151 2566 3155 2567
rect 3151 2561 3155 2562
rect 3231 2566 3235 2567
rect 3231 2561 3235 2562
rect 3359 2566 3363 2567
rect 3359 2561 3363 2562
rect 3487 2566 3491 2567
rect 3487 2561 3491 2562
rect 3943 2566 3947 2567
rect 3943 2561 3947 2562
rect 3074 2559 3080 2560
rect 3074 2555 3075 2559
rect 3079 2555 3080 2559
rect 3074 2554 3080 2555
rect 3076 2528 3078 2554
rect 3112 2537 3114 2561
rect 3194 2559 3200 2560
rect 3194 2555 3195 2559
rect 3199 2555 3200 2559
rect 3194 2554 3200 2555
rect 3110 2536 3116 2537
rect 3110 2532 3111 2536
rect 3115 2532 3116 2536
rect 3110 2531 3116 2532
rect 3196 2528 3198 2554
rect 3232 2537 3234 2561
rect 3314 2559 3320 2560
rect 3314 2555 3315 2559
rect 3319 2555 3320 2559
rect 3314 2554 3320 2555
rect 3230 2536 3236 2537
rect 3230 2532 3231 2536
rect 3235 2532 3236 2536
rect 3230 2531 3236 2532
rect 3316 2528 3318 2554
rect 3360 2537 3362 2561
rect 3442 2559 3448 2560
rect 3442 2555 3443 2559
rect 3447 2555 3448 2559
rect 3442 2554 3448 2555
rect 3434 2551 3440 2552
rect 3434 2547 3435 2551
rect 3439 2547 3440 2551
rect 3434 2546 3440 2547
rect 3358 2536 3364 2537
rect 3358 2532 3359 2536
rect 3363 2532 3364 2536
rect 3358 2531 3364 2532
rect 2458 2527 2464 2528
rect 2458 2523 2459 2527
rect 2463 2523 2464 2527
rect 2458 2522 2464 2523
rect 2570 2527 2576 2528
rect 2570 2523 2571 2527
rect 2575 2523 2576 2527
rect 2570 2522 2576 2523
rect 2690 2527 2696 2528
rect 2690 2523 2691 2527
rect 2695 2523 2696 2527
rect 2690 2522 2696 2523
rect 2818 2527 2824 2528
rect 2818 2523 2819 2527
rect 2823 2523 2824 2527
rect 2818 2522 2824 2523
rect 2826 2527 2832 2528
rect 2826 2523 2827 2527
rect 2831 2523 2832 2527
rect 2826 2522 2832 2523
rect 3066 2527 3072 2528
rect 3066 2523 3067 2527
rect 3071 2523 3072 2527
rect 3066 2522 3072 2523
rect 3074 2527 3080 2528
rect 3074 2523 3075 2527
rect 3079 2523 3080 2527
rect 3074 2522 3080 2523
rect 3194 2527 3200 2528
rect 3194 2523 3195 2527
rect 3199 2523 3200 2527
rect 3194 2522 3200 2523
rect 3314 2527 3320 2528
rect 3314 2523 3315 2527
rect 3319 2523 3320 2527
rect 3314 2522 3320 2523
rect 2382 2517 2388 2518
rect 2046 2516 2052 2517
rect 2046 2512 2047 2516
rect 2051 2512 2052 2516
rect 2382 2513 2383 2517
rect 2387 2513 2388 2517
rect 2382 2512 2388 2513
rect 2494 2517 2500 2518
rect 2494 2513 2495 2517
rect 2499 2513 2500 2517
rect 2494 2512 2500 2513
rect 2614 2517 2620 2518
rect 2614 2513 2615 2517
rect 2619 2513 2620 2517
rect 2614 2512 2620 2513
rect 2742 2517 2748 2518
rect 2742 2513 2743 2517
rect 2747 2513 2748 2517
rect 2742 2512 2748 2513
rect 2046 2511 2052 2512
rect 519 2494 523 2495
rect 519 2489 523 2490
rect 607 2494 611 2495
rect 607 2489 611 2490
rect 767 2494 771 2495
rect 767 2489 771 2490
rect 919 2494 923 2495
rect 919 2489 923 2490
rect 1063 2494 1067 2495
rect 1063 2489 1067 2490
rect 1199 2494 1203 2495
rect 1199 2489 1203 2490
rect 1335 2494 1339 2495
rect 1335 2489 1339 2490
rect 1463 2494 1467 2495
rect 1463 2489 1467 2490
rect 1591 2494 1595 2495
rect 1591 2489 1595 2490
rect 1727 2494 1731 2495
rect 1727 2489 1731 2490
rect 2007 2494 2011 2495
rect 2007 2489 2011 2490
rect 520 2465 522 2489
rect 518 2464 524 2465
rect 518 2460 519 2464
rect 523 2460 524 2464
rect 2008 2462 2010 2489
rect 2048 2487 2050 2511
rect 2384 2487 2386 2512
rect 2496 2487 2498 2512
rect 2616 2487 2618 2512
rect 2744 2487 2746 2512
rect 2047 2486 2051 2487
rect 2047 2481 2051 2482
rect 2383 2486 2387 2487
rect 2383 2481 2387 2482
rect 2495 2486 2499 2487
rect 2495 2481 2499 2482
rect 2535 2486 2539 2487
rect 2535 2481 2539 2482
rect 2615 2486 2619 2487
rect 2615 2481 2619 2482
rect 2711 2486 2715 2487
rect 2711 2481 2715 2482
rect 2743 2486 2747 2487
rect 2743 2481 2747 2482
rect 518 2459 524 2460
rect 2006 2461 2012 2462
rect 2048 2461 2050 2481
rect 2006 2457 2007 2461
rect 2011 2457 2012 2461
rect 2006 2456 2012 2457
rect 2046 2460 2052 2461
rect 2536 2460 2538 2481
rect 2712 2460 2714 2481
rect 2046 2456 2047 2460
rect 2051 2456 2052 2460
rect 210 2455 216 2456
rect 210 2451 211 2455
rect 215 2451 216 2455
rect 210 2450 216 2451
rect 306 2455 312 2456
rect 306 2451 307 2455
rect 311 2451 312 2455
rect 306 2450 312 2451
rect 402 2455 408 2456
rect 402 2451 403 2455
rect 407 2451 408 2455
rect 402 2450 408 2451
rect 498 2455 504 2456
rect 498 2451 499 2455
rect 503 2451 504 2455
rect 498 2450 504 2451
rect 506 2455 512 2456
rect 2046 2455 2052 2456
rect 2534 2459 2540 2460
rect 2534 2455 2535 2459
rect 2539 2455 2540 2459
rect 506 2451 507 2455
rect 511 2451 512 2455
rect 2534 2454 2540 2455
rect 2710 2459 2716 2460
rect 2710 2455 2711 2459
rect 2715 2455 2716 2459
rect 2710 2454 2716 2455
rect 506 2450 512 2451
rect 2610 2447 2616 2448
rect 230 2445 236 2446
rect 230 2441 231 2445
rect 235 2441 236 2445
rect 230 2440 236 2441
rect 326 2445 332 2446
rect 326 2441 327 2445
rect 331 2441 332 2445
rect 326 2440 332 2441
rect 422 2445 428 2446
rect 422 2441 423 2445
rect 427 2441 428 2445
rect 422 2440 428 2441
rect 518 2445 524 2446
rect 518 2441 519 2445
rect 523 2441 524 2445
rect 518 2440 524 2441
rect 2006 2444 2012 2445
rect 2006 2440 2007 2444
rect 2011 2440 2012 2444
rect 232 2403 234 2440
rect 328 2403 330 2440
rect 424 2403 426 2440
rect 520 2403 522 2440
rect 2006 2439 2012 2440
rect 2046 2443 2052 2444
rect 2046 2439 2047 2443
rect 2051 2439 2052 2443
rect 2610 2443 2611 2447
rect 2615 2443 2616 2447
rect 2610 2442 2616 2443
rect 2786 2447 2792 2448
rect 2786 2443 2787 2447
rect 2791 2443 2792 2447
rect 2786 2442 2792 2443
rect 2008 2403 2010 2439
rect 2046 2438 2052 2439
rect 2534 2440 2540 2441
rect 231 2402 235 2403
rect 231 2397 235 2398
rect 255 2402 259 2403
rect 255 2397 259 2398
rect 327 2402 331 2403
rect 327 2397 331 2398
rect 415 2402 419 2403
rect 415 2397 419 2398
rect 423 2402 427 2403
rect 423 2397 427 2398
rect 519 2402 523 2403
rect 519 2397 523 2398
rect 575 2402 579 2403
rect 575 2397 579 2398
rect 735 2402 739 2403
rect 735 2397 739 2398
rect 887 2402 891 2403
rect 887 2397 891 2398
rect 1039 2402 1043 2403
rect 1039 2397 1043 2398
rect 1183 2402 1187 2403
rect 1183 2397 1187 2398
rect 1327 2402 1331 2403
rect 1327 2397 1331 2398
rect 1479 2402 1483 2403
rect 1479 2397 1483 2398
rect 2007 2402 2011 2403
rect 2048 2399 2050 2438
rect 2534 2436 2535 2440
rect 2539 2436 2540 2440
rect 2534 2435 2540 2436
rect 2536 2399 2538 2435
rect 2612 2420 2614 2442
rect 2710 2440 2716 2441
rect 2710 2436 2711 2440
rect 2715 2436 2716 2440
rect 2710 2435 2716 2436
rect 2610 2419 2616 2420
rect 2610 2415 2611 2419
rect 2615 2415 2616 2419
rect 2610 2414 2616 2415
rect 2712 2399 2714 2435
rect 2788 2420 2790 2442
rect 2828 2428 2830 2522
rect 2870 2517 2876 2518
rect 2870 2513 2871 2517
rect 2875 2513 2876 2517
rect 2870 2512 2876 2513
rect 2990 2517 2996 2518
rect 2990 2513 2991 2517
rect 2995 2513 2996 2517
rect 2990 2512 2996 2513
rect 3110 2517 3116 2518
rect 3110 2513 3111 2517
rect 3115 2513 3116 2517
rect 3110 2512 3116 2513
rect 3230 2517 3236 2518
rect 3230 2513 3231 2517
rect 3235 2513 3236 2517
rect 3230 2512 3236 2513
rect 3358 2517 3364 2518
rect 3358 2513 3359 2517
rect 3363 2513 3364 2517
rect 3358 2512 3364 2513
rect 2872 2487 2874 2512
rect 2992 2487 2994 2512
rect 3112 2487 3114 2512
rect 3232 2487 3234 2512
rect 3360 2487 3362 2512
rect 2871 2486 2875 2487
rect 2871 2481 2875 2482
rect 2879 2486 2883 2487
rect 2879 2481 2883 2482
rect 2991 2486 2995 2487
rect 2991 2481 2995 2482
rect 3047 2486 3051 2487
rect 3047 2481 3051 2482
rect 3111 2486 3115 2487
rect 3111 2481 3115 2482
rect 3207 2486 3211 2487
rect 3207 2481 3211 2482
rect 3231 2486 3235 2487
rect 3231 2481 3235 2482
rect 3359 2486 3363 2487
rect 3359 2481 3363 2482
rect 2880 2460 2882 2481
rect 3048 2460 3050 2481
rect 3208 2460 3210 2481
rect 3360 2460 3362 2481
rect 2878 2459 2884 2460
rect 2878 2455 2879 2459
rect 2883 2455 2884 2459
rect 2878 2454 2884 2455
rect 3046 2459 3052 2460
rect 3046 2455 3047 2459
rect 3051 2455 3052 2459
rect 3046 2454 3052 2455
rect 3206 2459 3212 2460
rect 3206 2455 3207 2459
rect 3211 2455 3212 2459
rect 3206 2454 3212 2455
rect 3358 2459 3364 2460
rect 3358 2455 3359 2459
rect 3363 2455 3364 2459
rect 3358 2454 3364 2455
rect 3436 2452 3438 2546
rect 3444 2528 3446 2554
rect 3488 2537 3490 2561
rect 3486 2536 3492 2537
rect 3486 2532 3487 2536
rect 3491 2532 3492 2536
rect 3944 2534 3946 2561
rect 3486 2531 3492 2532
rect 3942 2533 3948 2534
rect 3942 2529 3943 2533
rect 3947 2529 3948 2533
rect 3942 2528 3948 2529
rect 3442 2527 3448 2528
rect 3442 2523 3443 2527
rect 3447 2523 3448 2527
rect 3442 2522 3448 2523
rect 3486 2517 3492 2518
rect 3486 2513 3487 2517
rect 3491 2513 3492 2517
rect 3486 2512 3492 2513
rect 3942 2516 3948 2517
rect 3942 2512 3943 2516
rect 3947 2512 3948 2516
rect 3488 2487 3490 2512
rect 3942 2511 3948 2512
rect 3944 2487 3946 2511
rect 3487 2486 3491 2487
rect 3487 2481 3491 2482
rect 3503 2486 3507 2487
rect 3503 2481 3507 2482
rect 3655 2486 3659 2487
rect 3655 2481 3659 2482
rect 3807 2486 3811 2487
rect 3807 2481 3811 2482
rect 3943 2486 3947 2487
rect 3943 2481 3947 2482
rect 3504 2460 3506 2481
rect 3656 2460 3658 2481
rect 3808 2460 3810 2481
rect 3944 2461 3946 2481
rect 3942 2460 3948 2461
rect 3502 2459 3508 2460
rect 3502 2455 3503 2459
rect 3507 2455 3508 2459
rect 3502 2454 3508 2455
rect 3654 2459 3660 2460
rect 3654 2455 3655 2459
rect 3659 2455 3660 2459
rect 3654 2454 3660 2455
rect 3806 2459 3812 2460
rect 3806 2455 3807 2459
rect 3811 2455 3812 2459
rect 3942 2456 3943 2460
rect 3947 2456 3948 2460
rect 3942 2455 3948 2456
rect 3806 2454 3812 2455
rect 3434 2451 3440 2452
rect 2954 2447 2960 2448
rect 2954 2443 2955 2447
rect 2959 2443 2960 2447
rect 2954 2442 2960 2443
rect 3122 2447 3128 2448
rect 3122 2443 3123 2447
rect 3127 2443 3128 2447
rect 3122 2442 3128 2443
rect 3282 2447 3288 2448
rect 3282 2443 3283 2447
rect 3287 2443 3288 2447
rect 3434 2447 3435 2451
rect 3439 2447 3440 2451
rect 3434 2446 3440 2447
rect 3442 2451 3448 2452
rect 3442 2447 3443 2451
rect 3447 2447 3448 2451
rect 3442 2446 3448 2447
rect 3586 2451 3592 2452
rect 3586 2447 3587 2451
rect 3591 2447 3592 2451
rect 3586 2446 3592 2447
rect 3282 2442 3288 2443
rect 2878 2440 2884 2441
rect 2878 2436 2879 2440
rect 2883 2436 2884 2440
rect 2878 2435 2884 2436
rect 2826 2427 2832 2428
rect 2826 2423 2827 2427
rect 2831 2423 2832 2427
rect 2826 2422 2832 2423
rect 2786 2419 2792 2420
rect 2786 2415 2787 2419
rect 2791 2415 2792 2419
rect 2786 2414 2792 2415
rect 2880 2399 2882 2435
rect 2956 2420 2958 2442
rect 3046 2440 3052 2441
rect 3046 2436 3047 2440
rect 3051 2436 3052 2440
rect 3046 2435 3052 2436
rect 2954 2419 2960 2420
rect 2954 2415 2955 2419
rect 2959 2415 2960 2419
rect 2954 2414 2960 2415
rect 3048 2399 3050 2435
rect 2007 2397 2011 2398
rect 2047 2398 2051 2399
rect 256 2376 258 2397
rect 416 2376 418 2397
rect 576 2376 578 2397
rect 736 2376 738 2397
rect 888 2376 890 2397
rect 1040 2376 1042 2397
rect 1184 2376 1186 2397
rect 1328 2376 1330 2397
rect 1480 2376 1482 2397
rect 2008 2377 2010 2397
rect 2047 2393 2051 2394
rect 2535 2398 2539 2399
rect 2535 2393 2539 2394
rect 2607 2398 2611 2399
rect 2607 2393 2611 2394
rect 2711 2398 2715 2399
rect 2711 2393 2715 2394
rect 2815 2398 2819 2399
rect 2815 2393 2819 2394
rect 2879 2398 2883 2399
rect 2879 2393 2883 2394
rect 3007 2398 3011 2399
rect 3007 2393 3011 2394
rect 3047 2398 3051 2399
rect 3047 2393 3051 2394
rect 2006 2376 2012 2377
rect 254 2375 260 2376
rect 134 2370 140 2371
rect 202 2371 208 2372
rect 202 2367 203 2371
rect 207 2367 208 2371
rect 254 2371 255 2375
rect 259 2371 260 2375
rect 254 2370 260 2371
rect 414 2375 420 2376
rect 414 2371 415 2375
rect 419 2371 420 2375
rect 414 2370 420 2371
rect 574 2375 580 2376
rect 574 2371 575 2375
rect 579 2371 580 2375
rect 574 2370 580 2371
rect 734 2375 740 2376
rect 734 2371 735 2375
rect 739 2371 740 2375
rect 734 2370 740 2371
rect 886 2375 892 2376
rect 886 2371 887 2375
rect 891 2371 892 2375
rect 886 2370 892 2371
rect 1038 2375 1044 2376
rect 1038 2371 1039 2375
rect 1043 2371 1044 2375
rect 1038 2370 1044 2371
rect 1182 2375 1188 2376
rect 1182 2371 1183 2375
rect 1187 2371 1188 2375
rect 1182 2370 1188 2371
rect 1326 2375 1332 2376
rect 1326 2371 1327 2375
rect 1331 2371 1332 2375
rect 1326 2370 1332 2371
rect 1478 2375 1484 2376
rect 1478 2371 1479 2375
rect 1483 2371 1484 2375
rect 2006 2372 2007 2376
rect 2011 2372 2012 2376
rect 2006 2371 2012 2372
rect 1478 2370 1484 2371
rect 202 2366 208 2367
rect 218 2367 224 2368
rect 218 2363 219 2367
rect 223 2363 224 2367
rect 218 2362 224 2363
rect 358 2367 364 2368
rect 358 2363 359 2367
rect 363 2363 364 2367
rect 358 2362 364 2363
rect 510 2367 516 2368
rect 510 2363 511 2367
rect 515 2363 516 2367
rect 510 2362 516 2363
rect 702 2367 708 2368
rect 702 2363 703 2367
rect 707 2363 708 2367
rect 970 2367 976 2368
rect 702 2362 708 2363
rect 962 2363 968 2364
rect 110 2359 116 2360
rect 110 2355 111 2359
rect 115 2355 116 2359
rect 110 2354 116 2355
rect 134 2356 140 2357
rect 112 2327 114 2354
rect 134 2352 135 2356
rect 139 2352 140 2356
rect 134 2351 140 2352
rect 136 2327 138 2351
rect 220 2336 222 2362
rect 254 2356 260 2357
rect 254 2352 255 2356
rect 259 2352 260 2356
rect 254 2351 260 2352
rect 218 2335 224 2336
rect 218 2331 219 2335
rect 223 2331 224 2335
rect 218 2330 224 2331
rect 256 2327 258 2351
rect 360 2336 362 2362
rect 414 2356 420 2357
rect 414 2352 415 2356
rect 419 2352 420 2356
rect 414 2351 420 2352
rect 358 2335 364 2336
rect 358 2331 359 2335
rect 363 2331 364 2335
rect 358 2330 364 2331
rect 416 2327 418 2351
rect 512 2336 514 2362
rect 574 2356 580 2357
rect 574 2352 575 2356
rect 579 2352 580 2356
rect 574 2351 580 2352
rect 510 2335 516 2336
rect 510 2331 511 2335
rect 515 2331 516 2335
rect 510 2330 516 2331
rect 576 2327 578 2351
rect 704 2336 706 2362
rect 962 2359 963 2363
rect 967 2359 968 2363
rect 970 2363 971 2367
rect 975 2363 976 2367
rect 970 2362 976 2363
rect 1122 2367 1128 2368
rect 1122 2363 1123 2367
rect 1127 2363 1128 2367
rect 1122 2362 1128 2363
rect 1266 2367 1272 2368
rect 1266 2363 1267 2367
rect 1271 2363 1272 2367
rect 1266 2362 1272 2363
rect 1414 2367 1420 2368
rect 1414 2363 1415 2367
rect 1419 2363 1420 2367
rect 2048 2366 2050 2393
rect 2608 2369 2610 2393
rect 2682 2391 2688 2392
rect 2682 2387 2683 2391
rect 2687 2387 2688 2391
rect 2682 2386 2688 2387
rect 2606 2368 2612 2369
rect 1414 2362 1420 2363
rect 2046 2365 2052 2366
rect 962 2358 968 2359
rect 734 2356 740 2357
rect 734 2352 735 2356
rect 739 2352 740 2356
rect 734 2351 740 2352
rect 886 2356 892 2357
rect 886 2352 887 2356
rect 891 2352 892 2356
rect 886 2351 892 2352
rect 702 2335 708 2336
rect 702 2331 703 2335
rect 707 2331 708 2335
rect 702 2330 708 2331
rect 736 2327 738 2351
rect 810 2331 816 2332
rect 810 2327 811 2331
rect 815 2327 816 2331
rect 888 2327 890 2351
rect 111 2326 115 2327
rect 111 2321 115 2322
rect 135 2326 139 2327
rect 135 2321 139 2322
rect 255 2326 259 2327
rect 255 2321 259 2322
rect 263 2326 267 2327
rect 263 2321 267 2322
rect 415 2326 419 2327
rect 415 2321 419 2322
rect 423 2326 427 2327
rect 423 2321 427 2322
rect 575 2326 579 2327
rect 575 2321 579 2322
rect 583 2326 587 2327
rect 583 2321 587 2322
rect 735 2326 739 2327
rect 735 2321 739 2322
rect 743 2326 747 2327
rect 810 2326 816 2327
rect 887 2326 891 2327
rect 743 2321 747 2322
rect 112 2294 114 2321
rect 136 2297 138 2321
rect 190 2319 196 2320
rect 190 2315 191 2319
rect 195 2315 196 2319
rect 190 2314 196 2315
rect 210 2319 216 2320
rect 210 2315 211 2319
rect 215 2315 216 2319
rect 210 2314 216 2315
rect 134 2296 140 2297
rect 110 2293 116 2294
rect 110 2289 111 2293
rect 115 2289 116 2293
rect 134 2292 135 2296
rect 139 2292 140 2296
rect 134 2291 140 2292
rect 110 2288 116 2289
rect 134 2277 140 2278
rect 110 2276 116 2277
rect 110 2272 111 2276
rect 115 2272 116 2276
rect 134 2273 135 2277
rect 139 2273 140 2277
rect 134 2272 140 2273
rect 110 2271 116 2272
rect 112 2247 114 2271
rect 136 2247 138 2272
rect 111 2246 115 2247
rect 111 2241 115 2242
rect 135 2246 139 2247
rect 135 2241 139 2242
rect 112 2221 114 2241
rect 110 2220 116 2221
rect 110 2216 111 2220
rect 115 2216 116 2220
rect 110 2215 116 2216
rect 192 2212 194 2314
rect 212 2288 214 2314
rect 264 2297 266 2321
rect 338 2319 344 2320
rect 338 2315 339 2319
rect 343 2315 344 2319
rect 338 2314 344 2315
rect 262 2296 268 2297
rect 262 2292 263 2296
rect 267 2292 268 2296
rect 262 2291 268 2292
rect 340 2288 342 2314
rect 424 2297 426 2321
rect 498 2319 504 2320
rect 498 2315 499 2319
rect 503 2315 504 2319
rect 498 2314 504 2315
rect 422 2296 428 2297
rect 422 2292 423 2296
rect 427 2292 428 2296
rect 422 2291 428 2292
rect 500 2288 502 2314
rect 584 2297 586 2321
rect 658 2319 664 2320
rect 658 2315 659 2319
rect 663 2315 664 2319
rect 658 2314 664 2315
rect 582 2296 588 2297
rect 582 2292 583 2296
rect 587 2292 588 2296
rect 582 2291 588 2292
rect 660 2288 662 2314
rect 744 2297 746 2321
rect 742 2296 748 2297
rect 742 2292 743 2296
rect 747 2292 748 2296
rect 742 2291 748 2292
rect 812 2288 814 2326
rect 887 2321 891 2322
rect 895 2326 899 2327
rect 895 2321 899 2322
rect 896 2297 898 2321
rect 964 2320 966 2358
rect 972 2336 974 2362
rect 1038 2356 1044 2357
rect 1038 2352 1039 2356
rect 1043 2352 1044 2356
rect 1038 2351 1044 2352
rect 970 2335 976 2336
rect 970 2331 971 2335
rect 975 2331 976 2335
rect 970 2330 976 2331
rect 1040 2327 1042 2351
rect 1124 2336 1126 2362
rect 1182 2356 1188 2357
rect 1182 2352 1183 2356
rect 1187 2352 1188 2356
rect 1182 2351 1188 2352
rect 1122 2335 1128 2336
rect 1122 2331 1123 2335
rect 1127 2331 1128 2335
rect 1122 2330 1128 2331
rect 1184 2327 1186 2351
rect 1268 2336 1270 2362
rect 1326 2356 1332 2357
rect 1326 2352 1327 2356
rect 1331 2352 1332 2356
rect 1326 2351 1332 2352
rect 1266 2335 1272 2336
rect 1266 2331 1267 2335
rect 1271 2331 1272 2335
rect 1266 2330 1272 2331
rect 1328 2327 1330 2351
rect 1416 2336 1418 2362
rect 2046 2361 2047 2365
rect 2051 2361 2052 2365
rect 2606 2364 2607 2368
rect 2611 2364 2612 2368
rect 2606 2363 2612 2364
rect 2046 2360 2052 2361
rect 2684 2360 2686 2386
rect 2816 2369 2818 2393
rect 2942 2383 2948 2384
rect 2942 2379 2943 2383
rect 2947 2379 2948 2383
rect 2942 2378 2948 2379
rect 2814 2368 2820 2369
rect 2814 2364 2815 2368
rect 2819 2364 2820 2368
rect 2814 2363 2820 2364
rect 2944 2360 2946 2378
rect 3008 2369 3010 2393
rect 3124 2392 3126 2442
rect 3206 2440 3212 2441
rect 3206 2436 3207 2440
rect 3211 2436 3212 2440
rect 3206 2435 3212 2436
rect 3208 2399 3210 2435
rect 3284 2420 3286 2442
rect 3358 2440 3364 2441
rect 3358 2436 3359 2440
rect 3363 2436 3364 2440
rect 3358 2435 3364 2436
rect 3282 2419 3288 2420
rect 3282 2415 3283 2419
rect 3287 2415 3288 2419
rect 3282 2414 3288 2415
rect 3360 2399 3362 2435
rect 3444 2428 3446 2446
rect 3502 2440 3508 2441
rect 3502 2436 3503 2440
rect 3507 2436 3508 2440
rect 3502 2435 3508 2436
rect 3442 2427 3448 2428
rect 3442 2423 3443 2427
rect 3447 2423 3448 2427
rect 3442 2422 3448 2423
rect 3504 2399 3506 2435
rect 3588 2420 3590 2446
rect 3942 2443 3948 2444
rect 3654 2440 3660 2441
rect 3654 2436 3655 2440
rect 3659 2436 3660 2440
rect 3654 2435 3660 2436
rect 3806 2440 3812 2441
rect 3806 2436 3807 2440
rect 3811 2436 3812 2440
rect 3942 2439 3943 2443
rect 3947 2439 3948 2443
rect 3942 2438 3948 2439
rect 3806 2435 3812 2436
rect 3586 2419 3592 2420
rect 3586 2415 3587 2419
rect 3591 2415 3592 2419
rect 3586 2414 3592 2415
rect 3656 2399 3658 2435
rect 3808 2399 3810 2435
rect 3906 2415 3912 2416
rect 3906 2411 3907 2415
rect 3911 2411 3912 2415
rect 3906 2410 3912 2411
rect 3191 2398 3195 2399
rect 3191 2393 3195 2394
rect 3207 2398 3211 2399
rect 3207 2393 3211 2394
rect 3359 2398 3363 2399
rect 3359 2393 3363 2394
rect 3503 2398 3507 2399
rect 3503 2393 3507 2394
rect 3519 2398 3523 2399
rect 3519 2393 3523 2394
rect 3655 2398 3659 2399
rect 3655 2393 3659 2394
rect 3679 2398 3683 2399
rect 3679 2393 3683 2394
rect 3807 2398 3811 2399
rect 3807 2393 3811 2394
rect 3839 2398 3843 2399
rect 3839 2393 3843 2394
rect 3122 2391 3128 2392
rect 3122 2387 3123 2391
rect 3127 2387 3128 2391
rect 3122 2386 3128 2387
rect 3192 2369 3194 2393
rect 3266 2391 3272 2392
rect 3266 2387 3267 2391
rect 3271 2387 3272 2391
rect 3266 2386 3272 2387
rect 3006 2368 3012 2369
rect 3006 2364 3007 2368
rect 3011 2364 3012 2368
rect 3006 2363 3012 2364
rect 3190 2368 3196 2369
rect 3190 2364 3191 2368
rect 3195 2364 3196 2368
rect 3190 2363 3196 2364
rect 3268 2360 3270 2386
rect 3360 2369 3362 2393
rect 3434 2391 3440 2392
rect 3434 2387 3435 2391
rect 3439 2387 3440 2391
rect 3434 2386 3440 2387
rect 3358 2368 3364 2369
rect 3358 2364 3359 2368
rect 3363 2364 3364 2368
rect 3358 2363 3364 2364
rect 3436 2360 3438 2386
rect 3520 2369 3522 2393
rect 3594 2391 3600 2392
rect 3594 2387 3595 2391
rect 3599 2387 3600 2391
rect 3594 2386 3600 2387
rect 3518 2368 3524 2369
rect 3518 2364 3519 2368
rect 3523 2364 3524 2368
rect 3518 2363 3524 2364
rect 3596 2360 3598 2386
rect 3618 2383 3624 2384
rect 3618 2379 3619 2383
rect 3623 2379 3624 2383
rect 3618 2378 3624 2379
rect 2006 2359 2012 2360
rect 1478 2356 1484 2357
rect 1478 2352 1479 2356
rect 1483 2352 1484 2356
rect 2006 2355 2007 2359
rect 2011 2355 2012 2359
rect 2006 2354 2012 2355
rect 2682 2359 2688 2360
rect 2682 2355 2683 2359
rect 2687 2355 2688 2359
rect 2682 2354 2688 2355
rect 2890 2359 2896 2360
rect 2890 2355 2891 2359
rect 2895 2355 2896 2359
rect 2890 2354 2896 2355
rect 2942 2359 2948 2360
rect 2942 2355 2943 2359
rect 2947 2355 2948 2359
rect 2942 2354 2948 2355
rect 3266 2359 3272 2360
rect 3266 2355 3267 2359
rect 3271 2355 3272 2359
rect 3266 2354 3272 2355
rect 3434 2359 3440 2360
rect 3434 2355 3435 2359
rect 3439 2355 3440 2359
rect 3434 2354 3440 2355
rect 3594 2359 3600 2360
rect 3594 2355 3595 2359
rect 3599 2355 3600 2359
rect 3594 2354 3600 2355
rect 1478 2351 1484 2352
rect 1414 2335 1420 2336
rect 1414 2331 1415 2335
rect 1419 2331 1420 2335
rect 1414 2330 1420 2331
rect 1480 2327 1482 2351
rect 1570 2331 1576 2332
rect 1570 2327 1571 2331
rect 1575 2327 1576 2331
rect 2008 2327 2010 2354
rect 2606 2349 2612 2350
rect 2046 2348 2052 2349
rect 2046 2344 2047 2348
rect 2051 2344 2052 2348
rect 2606 2345 2607 2349
rect 2611 2345 2612 2349
rect 2606 2344 2612 2345
rect 2814 2349 2820 2350
rect 2814 2345 2815 2349
rect 2819 2345 2820 2349
rect 2814 2344 2820 2345
rect 2046 2343 2052 2344
rect 1039 2326 1043 2327
rect 1039 2321 1043 2322
rect 1047 2326 1051 2327
rect 1047 2321 1051 2322
rect 1183 2326 1187 2327
rect 1183 2321 1187 2322
rect 1199 2326 1203 2327
rect 1199 2321 1203 2322
rect 1327 2326 1331 2327
rect 1327 2321 1331 2322
rect 1351 2326 1355 2327
rect 1351 2321 1355 2322
rect 1479 2326 1483 2327
rect 1479 2321 1483 2322
rect 1503 2326 1507 2327
rect 1570 2326 1576 2327
rect 2007 2326 2011 2327
rect 1503 2321 1507 2322
rect 962 2319 968 2320
rect 962 2315 963 2319
rect 967 2315 968 2319
rect 962 2314 968 2315
rect 970 2319 976 2320
rect 970 2315 971 2319
rect 975 2315 976 2319
rect 970 2314 976 2315
rect 894 2296 900 2297
rect 894 2292 895 2296
rect 899 2292 900 2296
rect 894 2291 900 2292
rect 972 2288 974 2314
rect 1048 2297 1050 2321
rect 1200 2297 1202 2321
rect 1254 2319 1260 2320
rect 1254 2315 1255 2319
rect 1259 2315 1260 2319
rect 1254 2314 1260 2315
rect 1274 2319 1280 2320
rect 1274 2315 1275 2319
rect 1279 2315 1280 2319
rect 1274 2314 1280 2315
rect 1046 2296 1052 2297
rect 1046 2292 1047 2296
rect 1051 2292 1052 2296
rect 1046 2291 1052 2292
rect 1198 2296 1204 2297
rect 1198 2292 1199 2296
rect 1203 2292 1204 2296
rect 1198 2291 1204 2292
rect 210 2287 216 2288
rect 210 2283 211 2287
rect 215 2283 216 2287
rect 210 2282 216 2283
rect 338 2287 344 2288
rect 338 2283 339 2287
rect 343 2283 344 2287
rect 338 2282 344 2283
rect 498 2287 504 2288
rect 498 2283 499 2287
rect 503 2283 504 2287
rect 498 2282 504 2283
rect 658 2287 664 2288
rect 658 2283 659 2287
rect 663 2283 664 2287
rect 658 2282 664 2283
rect 810 2287 816 2288
rect 810 2283 811 2287
rect 815 2283 816 2287
rect 810 2282 816 2283
rect 970 2287 976 2288
rect 970 2283 971 2287
rect 975 2283 976 2287
rect 970 2282 976 2283
rect 1014 2287 1020 2288
rect 1014 2283 1015 2287
rect 1019 2283 1020 2287
rect 1014 2282 1020 2283
rect 262 2277 268 2278
rect 262 2273 263 2277
rect 267 2273 268 2277
rect 262 2272 268 2273
rect 422 2277 428 2278
rect 422 2273 423 2277
rect 427 2273 428 2277
rect 422 2272 428 2273
rect 582 2277 588 2278
rect 582 2273 583 2277
rect 587 2273 588 2277
rect 582 2272 588 2273
rect 742 2277 748 2278
rect 742 2273 743 2277
rect 747 2273 748 2277
rect 742 2272 748 2273
rect 894 2277 900 2278
rect 894 2273 895 2277
rect 899 2273 900 2277
rect 894 2272 900 2273
rect 264 2247 266 2272
rect 424 2247 426 2272
rect 584 2247 586 2272
rect 744 2247 746 2272
rect 896 2247 898 2272
rect 223 2246 227 2247
rect 223 2241 227 2242
rect 263 2246 267 2247
rect 263 2241 267 2242
rect 351 2246 355 2247
rect 351 2241 355 2242
rect 423 2246 427 2247
rect 423 2241 427 2242
rect 495 2246 499 2247
rect 495 2241 499 2242
rect 583 2246 587 2247
rect 583 2241 587 2242
rect 647 2246 651 2247
rect 647 2241 651 2242
rect 743 2246 747 2247
rect 743 2241 747 2242
rect 799 2246 803 2247
rect 799 2241 803 2242
rect 895 2246 899 2247
rect 895 2241 899 2242
rect 959 2246 963 2247
rect 959 2241 963 2242
rect 224 2220 226 2241
rect 352 2220 354 2241
rect 496 2220 498 2241
rect 648 2220 650 2241
rect 800 2220 802 2241
rect 960 2220 962 2241
rect 222 2219 228 2220
rect 222 2215 223 2219
rect 227 2215 228 2219
rect 222 2214 228 2215
rect 350 2219 356 2220
rect 350 2215 351 2219
rect 355 2215 356 2219
rect 350 2214 356 2215
rect 494 2219 500 2220
rect 494 2215 495 2219
rect 499 2215 500 2219
rect 494 2214 500 2215
rect 646 2219 652 2220
rect 646 2215 647 2219
rect 651 2215 652 2219
rect 646 2214 652 2215
rect 798 2219 804 2220
rect 798 2215 799 2219
rect 803 2215 804 2219
rect 798 2214 804 2215
rect 958 2219 964 2220
rect 958 2215 959 2219
rect 963 2215 964 2219
rect 958 2214 964 2215
rect 190 2211 196 2212
rect 190 2207 191 2211
rect 195 2207 196 2211
rect 190 2206 196 2207
rect 306 2211 312 2212
rect 306 2207 307 2211
rect 311 2207 312 2211
rect 306 2206 312 2207
rect 110 2203 116 2204
rect 110 2199 111 2203
rect 115 2199 116 2203
rect 110 2198 116 2199
rect 222 2200 228 2201
rect 112 2171 114 2198
rect 222 2196 223 2200
rect 227 2196 228 2200
rect 222 2195 228 2196
rect 224 2171 226 2195
rect 308 2180 310 2206
rect 350 2200 356 2201
rect 350 2196 351 2200
rect 355 2196 356 2200
rect 350 2195 356 2196
rect 494 2200 500 2201
rect 494 2196 495 2200
rect 499 2196 500 2200
rect 494 2195 500 2196
rect 646 2200 652 2201
rect 646 2196 647 2200
rect 651 2196 652 2200
rect 646 2195 652 2196
rect 798 2200 804 2201
rect 798 2196 799 2200
rect 803 2196 804 2200
rect 798 2195 804 2196
rect 958 2200 964 2201
rect 958 2196 959 2200
rect 963 2196 964 2200
rect 958 2195 964 2196
rect 306 2179 312 2180
rect 306 2175 307 2179
rect 311 2175 312 2179
rect 306 2174 312 2175
rect 352 2171 354 2195
rect 496 2171 498 2195
rect 648 2171 650 2195
rect 800 2171 802 2195
rect 960 2171 962 2195
rect 1016 2180 1018 2282
rect 1046 2277 1052 2278
rect 1046 2273 1047 2277
rect 1051 2273 1052 2277
rect 1046 2272 1052 2273
rect 1198 2277 1204 2278
rect 1198 2273 1199 2277
rect 1203 2273 1204 2277
rect 1198 2272 1204 2273
rect 1048 2247 1050 2272
rect 1200 2247 1202 2272
rect 1047 2246 1051 2247
rect 1047 2241 1051 2242
rect 1119 2246 1123 2247
rect 1119 2241 1123 2242
rect 1199 2246 1203 2247
rect 1199 2241 1203 2242
rect 1120 2220 1122 2241
rect 1118 2219 1124 2220
rect 1118 2215 1119 2219
rect 1123 2215 1124 2219
rect 1118 2214 1124 2215
rect 1256 2212 1258 2314
rect 1276 2288 1278 2314
rect 1352 2297 1354 2321
rect 1426 2319 1432 2320
rect 1426 2315 1427 2319
rect 1431 2315 1432 2319
rect 1426 2314 1432 2315
rect 1350 2296 1356 2297
rect 1350 2292 1351 2296
rect 1355 2292 1356 2296
rect 1350 2291 1356 2292
rect 1428 2288 1430 2314
rect 1504 2297 1506 2321
rect 1502 2296 1508 2297
rect 1502 2292 1503 2296
rect 1507 2292 1508 2296
rect 1502 2291 1508 2292
rect 1572 2288 1574 2326
rect 2007 2321 2011 2322
rect 2008 2294 2010 2321
rect 2048 2307 2050 2343
rect 2608 2307 2610 2344
rect 2816 2307 2818 2344
rect 2047 2306 2051 2307
rect 2047 2301 2051 2302
rect 2071 2306 2075 2307
rect 2071 2301 2075 2302
rect 2167 2306 2171 2307
rect 2167 2301 2171 2302
rect 2271 2306 2275 2307
rect 2271 2301 2275 2302
rect 2415 2306 2419 2307
rect 2415 2301 2419 2302
rect 2575 2306 2579 2307
rect 2575 2301 2579 2302
rect 2607 2306 2611 2307
rect 2607 2301 2611 2302
rect 2743 2306 2747 2307
rect 2743 2301 2747 2302
rect 2815 2306 2819 2307
rect 2815 2301 2819 2302
rect 2006 2293 2012 2294
rect 2006 2289 2007 2293
rect 2011 2289 2012 2293
rect 2006 2288 2012 2289
rect 1274 2287 1280 2288
rect 1274 2283 1275 2287
rect 1279 2283 1280 2287
rect 1274 2282 1280 2283
rect 1426 2287 1432 2288
rect 1426 2283 1427 2287
rect 1431 2283 1432 2287
rect 1426 2282 1432 2283
rect 1570 2287 1576 2288
rect 1570 2283 1571 2287
rect 1575 2283 1576 2287
rect 1570 2282 1576 2283
rect 2048 2281 2050 2301
rect 2046 2280 2052 2281
rect 2072 2280 2074 2301
rect 2168 2280 2170 2301
rect 2272 2280 2274 2301
rect 2416 2280 2418 2301
rect 2576 2280 2578 2301
rect 2744 2280 2746 2301
rect 1350 2277 1356 2278
rect 1350 2273 1351 2277
rect 1355 2273 1356 2277
rect 1350 2272 1356 2273
rect 1502 2277 1508 2278
rect 1502 2273 1503 2277
rect 1507 2273 1508 2277
rect 1502 2272 1508 2273
rect 2006 2276 2012 2277
rect 2006 2272 2007 2276
rect 2011 2272 2012 2276
rect 2046 2276 2047 2280
rect 2051 2276 2052 2280
rect 2046 2275 2052 2276
rect 2070 2279 2076 2280
rect 2070 2275 2071 2279
rect 2075 2275 2076 2279
rect 2070 2274 2076 2275
rect 2166 2279 2172 2280
rect 2166 2275 2167 2279
rect 2171 2275 2172 2279
rect 2166 2274 2172 2275
rect 2270 2279 2276 2280
rect 2270 2275 2271 2279
rect 2275 2275 2276 2279
rect 2270 2274 2276 2275
rect 2414 2279 2420 2280
rect 2414 2275 2415 2279
rect 2419 2275 2420 2279
rect 2414 2274 2420 2275
rect 2574 2279 2580 2280
rect 2574 2275 2575 2279
rect 2579 2275 2580 2279
rect 2574 2274 2580 2275
rect 2742 2279 2748 2280
rect 2742 2275 2743 2279
rect 2747 2275 2748 2279
rect 2742 2274 2748 2275
rect 1352 2247 1354 2272
rect 1504 2247 1506 2272
rect 2006 2271 2012 2272
rect 2250 2271 2256 2272
rect 2008 2247 2010 2271
rect 2146 2267 2152 2268
rect 2046 2263 2052 2264
rect 2046 2259 2047 2263
rect 2051 2259 2052 2263
rect 2146 2263 2147 2267
rect 2151 2263 2152 2267
rect 2146 2262 2152 2263
rect 2242 2267 2248 2268
rect 2242 2263 2243 2267
rect 2247 2263 2248 2267
rect 2250 2267 2251 2271
rect 2255 2267 2256 2271
rect 2250 2266 2256 2267
rect 2358 2271 2364 2272
rect 2358 2267 2359 2271
rect 2363 2267 2364 2271
rect 2358 2266 2364 2267
rect 2534 2271 2540 2272
rect 2534 2267 2535 2271
rect 2539 2267 2540 2271
rect 2534 2266 2540 2267
rect 2658 2271 2664 2272
rect 2658 2267 2659 2271
rect 2663 2267 2664 2271
rect 2658 2266 2664 2267
rect 2870 2271 2876 2272
rect 2870 2267 2871 2271
rect 2875 2267 2876 2271
rect 2870 2266 2876 2267
rect 2242 2262 2248 2263
rect 2046 2258 2052 2259
rect 2070 2260 2076 2261
rect 1279 2246 1283 2247
rect 1279 2241 1283 2242
rect 1351 2246 1355 2247
rect 1351 2241 1355 2242
rect 1439 2246 1443 2247
rect 1439 2241 1443 2242
rect 1503 2246 1507 2247
rect 1503 2241 1507 2242
rect 1599 2246 1603 2247
rect 1599 2241 1603 2242
rect 2007 2246 2011 2247
rect 2007 2241 2011 2242
rect 1280 2220 1282 2241
rect 1440 2220 1442 2241
rect 1600 2220 1602 2241
rect 2008 2221 2010 2241
rect 2048 2231 2050 2258
rect 2070 2256 2071 2260
rect 2075 2256 2076 2260
rect 2070 2255 2076 2256
rect 2072 2231 2074 2255
rect 2148 2240 2150 2262
rect 2166 2260 2172 2261
rect 2166 2256 2167 2260
rect 2171 2256 2172 2260
rect 2166 2255 2172 2256
rect 2146 2239 2152 2240
rect 2146 2235 2147 2239
rect 2151 2235 2152 2239
rect 2146 2234 2152 2235
rect 2168 2231 2170 2255
rect 2047 2230 2051 2231
rect 2047 2225 2051 2226
rect 2071 2230 2075 2231
rect 2071 2225 2075 2226
rect 2167 2230 2171 2231
rect 2167 2225 2171 2226
rect 2175 2230 2179 2231
rect 2175 2225 2179 2226
rect 2006 2220 2012 2221
rect 1278 2219 1284 2220
rect 1278 2215 1279 2219
rect 1283 2215 1284 2219
rect 1278 2214 1284 2215
rect 1438 2219 1444 2220
rect 1438 2215 1439 2219
rect 1443 2215 1444 2219
rect 1438 2214 1444 2215
rect 1598 2219 1604 2220
rect 1598 2215 1599 2219
rect 1603 2215 1604 2219
rect 2006 2216 2007 2220
rect 2011 2216 2012 2220
rect 2006 2215 2012 2216
rect 1598 2214 1604 2215
rect 1254 2211 1260 2212
rect 1034 2207 1040 2208
rect 1034 2203 1035 2207
rect 1039 2203 1040 2207
rect 1034 2202 1040 2203
rect 1194 2207 1200 2208
rect 1194 2203 1195 2207
rect 1199 2203 1200 2207
rect 1254 2207 1255 2211
rect 1259 2207 1260 2211
rect 1254 2206 1260 2207
rect 1194 2202 1200 2203
rect 2006 2203 2012 2204
rect 1036 2180 1038 2202
rect 1118 2200 1124 2201
rect 1118 2196 1119 2200
rect 1123 2196 1124 2200
rect 1118 2195 1124 2196
rect 1014 2179 1020 2180
rect 1014 2175 1015 2179
rect 1019 2175 1020 2179
rect 1014 2174 1020 2175
rect 1034 2179 1040 2180
rect 1034 2175 1035 2179
rect 1039 2175 1040 2179
rect 1034 2174 1040 2175
rect 1120 2171 1122 2195
rect 111 2170 115 2171
rect 111 2165 115 2166
rect 223 2170 227 2171
rect 223 2165 227 2166
rect 351 2170 355 2171
rect 351 2165 355 2166
rect 471 2170 475 2171
rect 471 2165 475 2166
rect 495 2170 499 2171
rect 495 2165 499 2166
rect 567 2170 571 2171
rect 567 2165 571 2166
rect 647 2170 651 2171
rect 647 2165 651 2166
rect 679 2170 683 2171
rect 679 2165 683 2166
rect 799 2170 803 2171
rect 799 2165 803 2166
rect 807 2170 811 2171
rect 807 2165 811 2166
rect 943 2170 947 2171
rect 943 2165 947 2166
rect 959 2170 963 2171
rect 959 2165 963 2166
rect 1079 2170 1083 2171
rect 1079 2165 1083 2166
rect 1119 2170 1123 2171
rect 1119 2165 1123 2166
rect 112 2138 114 2165
rect 472 2141 474 2165
rect 546 2163 552 2164
rect 546 2159 547 2163
rect 551 2159 552 2163
rect 546 2158 552 2159
rect 470 2140 476 2141
rect 110 2137 116 2138
rect 110 2133 111 2137
rect 115 2133 116 2137
rect 470 2136 471 2140
rect 475 2136 476 2140
rect 470 2135 476 2136
rect 110 2132 116 2133
rect 548 2132 550 2158
rect 568 2141 570 2165
rect 670 2163 676 2164
rect 670 2159 671 2163
rect 675 2159 676 2163
rect 670 2158 676 2159
rect 566 2140 572 2141
rect 566 2136 567 2140
rect 571 2136 572 2140
rect 566 2135 572 2136
rect 672 2132 674 2158
rect 680 2141 682 2165
rect 808 2141 810 2165
rect 890 2163 896 2164
rect 890 2159 891 2163
rect 895 2159 896 2163
rect 890 2158 896 2159
rect 678 2140 684 2141
rect 678 2136 679 2140
rect 683 2136 684 2140
rect 678 2135 684 2136
rect 806 2140 812 2141
rect 806 2136 807 2140
rect 811 2136 812 2140
rect 806 2135 812 2136
rect 892 2132 894 2158
rect 944 2141 946 2165
rect 1080 2141 1082 2165
rect 1196 2164 1198 2202
rect 1278 2200 1284 2201
rect 1278 2196 1279 2200
rect 1283 2196 1284 2200
rect 1278 2195 1284 2196
rect 1438 2200 1444 2201
rect 1438 2196 1439 2200
rect 1443 2196 1444 2200
rect 1438 2195 1444 2196
rect 1598 2200 1604 2201
rect 1598 2196 1599 2200
rect 1603 2196 1604 2200
rect 2006 2199 2007 2203
rect 2011 2199 2012 2203
rect 2006 2198 2012 2199
rect 2048 2198 2050 2225
rect 2072 2201 2074 2225
rect 2154 2223 2160 2224
rect 2154 2219 2155 2223
rect 2159 2219 2160 2223
rect 2154 2218 2160 2219
rect 2070 2200 2076 2201
rect 1598 2195 1604 2196
rect 1280 2171 1282 2195
rect 1440 2171 1442 2195
rect 1578 2175 1584 2176
rect 1578 2171 1579 2175
rect 1583 2171 1584 2175
rect 1600 2171 1602 2195
rect 2008 2171 2010 2198
rect 2046 2197 2052 2198
rect 2046 2193 2047 2197
rect 2051 2193 2052 2197
rect 2070 2196 2071 2200
rect 2075 2196 2076 2200
rect 2070 2195 2076 2196
rect 2046 2192 2052 2193
rect 2156 2192 2158 2218
rect 2176 2201 2178 2225
rect 2244 2224 2246 2262
rect 2252 2248 2254 2266
rect 2270 2260 2276 2261
rect 2270 2256 2271 2260
rect 2275 2256 2276 2260
rect 2270 2255 2276 2256
rect 2250 2247 2256 2248
rect 2250 2243 2251 2247
rect 2255 2243 2256 2247
rect 2250 2242 2256 2243
rect 2272 2231 2274 2255
rect 2360 2240 2362 2266
rect 2414 2260 2420 2261
rect 2414 2256 2415 2260
rect 2419 2256 2420 2260
rect 2414 2255 2420 2256
rect 2358 2239 2364 2240
rect 2358 2235 2359 2239
rect 2363 2235 2364 2239
rect 2358 2234 2364 2235
rect 2416 2231 2418 2255
rect 2536 2240 2538 2266
rect 2574 2260 2580 2261
rect 2574 2256 2575 2260
rect 2579 2256 2580 2260
rect 2574 2255 2580 2256
rect 2534 2239 2540 2240
rect 2534 2235 2535 2239
rect 2539 2235 2540 2239
rect 2534 2234 2540 2235
rect 2576 2231 2578 2255
rect 2660 2240 2662 2266
rect 2742 2260 2748 2261
rect 2742 2256 2743 2260
rect 2747 2256 2748 2260
rect 2742 2255 2748 2256
rect 2658 2239 2664 2240
rect 2658 2235 2659 2239
rect 2663 2235 2664 2239
rect 2658 2234 2664 2235
rect 2698 2235 2704 2236
rect 2698 2231 2699 2235
rect 2703 2231 2704 2235
rect 2744 2231 2746 2255
rect 2271 2230 2275 2231
rect 2271 2225 2275 2226
rect 2319 2230 2323 2231
rect 2319 2225 2323 2226
rect 2415 2230 2419 2231
rect 2415 2225 2419 2226
rect 2471 2230 2475 2231
rect 2471 2225 2475 2226
rect 2575 2230 2579 2231
rect 2575 2225 2579 2226
rect 2623 2230 2627 2231
rect 2698 2230 2704 2231
rect 2743 2230 2747 2231
rect 2623 2225 2627 2226
rect 2242 2223 2248 2224
rect 2242 2219 2243 2223
rect 2247 2219 2248 2223
rect 2242 2218 2248 2219
rect 2320 2201 2322 2225
rect 2354 2223 2360 2224
rect 2354 2219 2355 2223
rect 2359 2219 2360 2223
rect 2354 2218 2360 2219
rect 2394 2223 2400 2224
rect 2394 2219 2395 2223
rect 2399 2219 2400 2223
rect 2394 2218 2400 2219
rect 2174 2200 2180 2201
rect 2174 2196 2175 2200
rect 2179 2196 2180 2200
rect 2174 2195 2180 2196
rect 2318 2200 2324 2201
rect 2318 2196 2319 2200
rect 2323 2196 2324 2200
rect 2318 2195 2324 2196
rect 2154 2191 2160 2192
rect 2154 2187 2155 2191
rect 2159 2187 2160 2191
rect 2154 2186 2160 2187
rect 2070 2181 2076 2182
rect 2046 2180 2052 2181
rect 2046 2176 2047 2180
rect 2051 2176 2052 2180
rect 2070 2177 2071 2181
rect 2075 2177 2076 2181
rect 2070 2176 2076 2177
rect 2174 2181 2180 2182
rect 2174 2177 2175 2181
rect 2179 2177 2180 2181
rect 2174 2176 2180 2177
rect 2318 2181 2324 2182
rect 2318 2177 2319 2181
rect 2323 2177 2324 2181
rect 2318 2176 2324 2177
rect 2046 2175 2052 2176
rect 1223 2170 1227 2171
rect 1223 2165 1227 2166
rect 1279 2170 1283 2171
rect 1279 2165 1283 2166
rect 1367 2170 1371 2171
rect 1367 2165 1371 2166
rect 1439 2170 1443 2171
rect 1439 2165 1443 2166
rect 1503 2170 1507 2171
rect 1578 2170 1584 2171
rect 1599 2170 1603 2171
rect 1503 2165 1507 2166
rect 1194 2163 1200 2164
rect 1194 2159 1195 2163
rect 1199 2159 1200 2163
rect 1194 2158 1200 2159
rect 1224 2141 1226 2165
rect 1368 2141 1370 2165
rect 1504 2141 1506 2165
rect 942 2140 948 2141
rect 942 2136 943 2140
rect 947 2136 948 2140
rect 942 2135 948 2136
rect 1078 2140 1084 2141
rect 1078 2136 1079 2140
rect 1083 2136 1084 2140
rect 1078 2135 1084 2136
rect 1222 2140 1228 2141
rect 1222 2136 1223 2140
rect 1227 2136 1228 2140
rect 1222 2135 1228 2136
rect 1366 2140 1372 2141
rect 1366 2136 1367 2140
rect 1371 2136 1372 2140
rect 1366 2135 1372 2136
rect 1502 2140 1508 2141
rect 1502 2136 1503 2140
rect 1507 2136 1508 2140
rect 1502 2135 1508 2136
rect 1580 2132 1582 2170
rect 1599 2165 1603 2166
rect 1639 2170 1643 2171
rect 1639 2165 1643 2166
rect 1783 2170 1787 2171
rect 1783 2165 1787 2166
rect 1903 2170 1907 2171
rect 1903 2165 1907 2166
rect 2007 2170 2011 2171
rect 2007 2165 2011 2166
rect 1586 2155 1592 2156
rect 1586 2151 1587 2155
rect 1591 2151 1592 2155
rect 1586 2150 1592 2151
rect 1588 2132 1590 2150
rect 1640 2141 1642 2165
rect 1730 2163 1736 2164
rect 1730 2159 1731 2163
rect 1735 2159 1736 2163
rect 1730 2158 1736 2159
rect 1638 2140 1644 2141
rect 1638 2136 1639 2140
rect 1643 2136 1644 2140
rect 1638 2135 1644 2136
rect 546 2131 552 2132
rect 546 2127 547 2131
rect 551 2127 552 2131
rect 546 2126 552 2127
rect 670 2131 676 2132
rect 670 2127 671 2131
rect 675 2127 676 2131
rect 670 2126 676 2127
rect 890 2131 896 2132
rect 890 2127 891 2131
rect 895 2127 896 2131
rect 890 2126 896 2127
rect 1298 2131 1304 2132
rect 1298 2127 1299 2131
rect 1303 2127 1304 2131
rect 1298 2126 1304 2127
rect 1578 2131 1584 2132
rect 1578 2127 1579 2131
rect 1583 2127 1584 2131
rect 1578 2126 1584 2127
rect 1586 2131 1592 2132
rect 1586 2127 1587 2131
rect 1591 2127 1592 2131
rect 1586 2126 1592 2127
rect 470 2121 476 2122
rect 110 2120 116 2121
rect 110 2116 111 2120
rect 115 2116 116 2120
rect 470 2117 471 2121
rect 475 2117 476 2121
rect 470 2116 476 2117
rect 566 2121 572 2122
rect 566 2117 567 2121
rect 571 2117 572 2121
rect 566 2116 572 2117
rect 678 2121 684 2122
rect 678 2117 679 2121
rect 683 2117 684 2121
rect 678 2116 684 2117
rect 806 2121 812 2122
rect 806 2117 807 2121
rect 811 2117 812 2121
rect 806 2116 812 2117
rect 942 2121 948 2122
rect 942 2117 943 2121
rect 947 2117 948 2121
rect 942 2116 948 2117
rect 1078 2121 1084 2122
rect 1078 2117 1079 2121
rect 1083 2117 1084 2121
rect 1078 2116 1084 2117
rect 1222 2121 1228 2122
rect 1222 2117 1223 2121
rect 1227 2117 1228 2121
rect 1222 2116 1228 2117
rect 110 2115 116 2116
rect 112 2095 114 2115
rect 472 2095 474 2116
rect 568 2095 570 2116
rect 680 2095 682 2116
rect 808 2095 810 2116
rect 944 2095 946 2116
rect 1080 2095 1082 2116
rect 1224 2095 1226 2116
rect 111 2094 115 2095
rect 111 2089 115 2090
rect 471 2094 475 2095
rect 471 2089 475 2090
rect 567 2094 571 2095
rect 567 2089 571 2090
rect 623 2094 627 2095
rect 623 2089 627 2090
rect 679 2094 683 2095
rect 679 2089 683 2090
rect 735 2094 739 2095
rect 735 2089 739 2090
rect 807 2094 811 2095
rect 807 2089 811 2090
rect 855 2094 859 2095
rect 855 2089 859 2090
rect 943 2094 947 2095
rect 943 2089 947 2090
rect 983 2094 987 2095
rect 983 2089 987 2090
rect 1079 2094 1083 2095
rect 1079 2089 1083 2090
rect 1119 2094 1123 2095
rect 1119 2089 1123 2090
rect 1223 2094 1227 2095
rect 1223 2089 1227 2090
rect 1255 2094 1259 2095
rect 1255 2089 1259 2090
rect 112 2069 114 2089
rect 110 2068 116 2069
rect 624 2068 626 2089
rect 736 2068 738 2089
rect 856 2068 858 2089
rect 984 2068 986 2089
rect 1120 2068 1122 2089
rect 1256 2068 1258 2089
rect 110 2064 111 2068
rect 115 2064 116 2068
rect 110 2063 116 2064
rect 622 2067 628 2068
rect 622 2063 623 2067
rect 627 2063 628 2067
rect 622 2062 628 2063
rect 734 2067 740 2068
rect 734 2063 735 2067
rect 739 2063 740 2067
rect 734 2062 740 2063
rect 854 2067 860 2068
rect 854 2063 855 2067
rect 859 2063 860 2067
rect 854 2062 860 2063
rect 982 2067 988 2068
rect 982 2063 983 2067
rect 987 2063 988 2067
rect 982 2062 988 2063
rect 1118 2067 1124 2068
rect 1118 2063 1119 2067
rect 1123 2063 1124 2067
rect 1118 2062 1124 2063
rect 1254 2067 1260 2068
rect 1254 2063 1255 2067
rect 1259 2063 1260 2067
rect 1254 2062 1260 2063
rect 698 2055 704 2056
rect 110 2051 116 2052
rect 110 2047 111 2051
rect 115 2047 116 2051
rect 698 2051 699 2055
rect 703 2051 704 2055
rect 698 2050 704 2051
rect 810 2055 816 2056
rect 810 2051 811 2055
rect 815 2051 816 2055
rect 810 2050 816 2051
rect 930 2055 936 2056
rect 930 2051 931 2055
rect 935 2051 936 2055
rect 930 2050 936 2051
rect 1058 2055 1064 2056
rect 1058 2051 1059 2055
rect 1063 2051 1064 2055
rect 1058 2050 1064 2051
rect 110 2046 116 2047
rect 622 2048 628 2049
rect 112 2015 114 2046
rect 622 2044 623 2048
rect 627 2044 628 2048
rect 622 2043 628 2044
rect 624 2015 626 2043
rect 700 2028 702 2050
rect 734 2048 740 2049
rect 734 2044 735 2048
rect 739 2044 740 2048
rect 734 2043 740 2044
rect 698 2027 704 2028
rect 698 2023 699 2027
rect 703 2023 704 2027
rect 698 2022 704 2023
rect 736 2015 738 2043
rect 812 2028 814 2050
rect 854 2048 860 2049
rect 854 2044 855 2048
rect 859 2044 860 2048
rect 854 2043 860 2044
rect 810 2027 816 2028
rect 810 2023 811 2027
rect 815 2023 816 2027
rect 810 2022 816 2023
rect 810 2019 816 2020
rect 810 2015 811 2019
rect 815 2015 816 2019
rect 856 2015 858 2043
rect 932 2028 934 2050
rect 982 2048 988 2049
rect 982 2044 983 2048
rect 987 2044 988 2048
rect 982 2043 988 2044
rect 930 2027 936 2028
rect 930 2023 931 2027
rect 935 2023 936 2027
rect 930 2022 936 2023
rect 984 2015 986 2043
rect 1060 2028 1062 2050
rect 1118 2048 1124 2049
rect 1118 2044 1119 2048
rect 1123 2044 1124 2048
rect 1118 2043 1124 2044
rect 1254 2048 1260 2049
rect 1254 2044 1255 2048
rect 1259 2044 1260 2048
rect 1254 2043 1260 2044
rect 1058 2027 1064 2028
rect 1058 2023 1059 2027
rect 1063 2023 1064 2027
rect 1058 2022 1064 2023
rect 1120 2015 1122 2043
rect 1256 2015 1258 2043
rect 1300 2028 1302 2126
rect 1366 2121 1372 2122
rect 1366 2117 1367 2121
rect 1371 2117 1372 2121
rect 1366 2116 1372 2117
rect 1502 2121 1508 2122
rect 1502 2117 1503 2121
rect 1507 2117 1508 2121
rect 1502 2116 1508 2117
rect 1638 2121 1644 2122
rect 1638 2117 1639 2121
rect 1643 2117 1644 2121
rect 1638 2116 1644 2117
rect 1368 2095 1370 2116
rect 1504 2095 1506 2116
rect 1640 2095 1642 2116
rect 1367 2094 1371 2095
rect 1367 2089 1371 2090
rect 1391 2094 1395 2095
rect 1391 2089 1395 2090
rect 1503 2094 1507 2095
rect 1503 2089 1507 2090
rect 1527 2094 1531 2095
rect 1527 2089 1531 2090
rect 1639 2094 1643 2095
rect 1639 2089 1643 2090
rect 1655 2094 1659 2095
rect 1655 2089 1659 2090
rect 1392 2068 1394 2089
rect 1528 2068 1530 2089
rect 1656 2068 1658 2089
rect 1390 2067 1396 2068
rect 1390 2063 1391 2067
rect 1395 2063 1396 2067
rect 1390 2062 1396 2063
rect 1526 2067 1532 2068
rect 1526 2063 1527 2067
rect 1531 2063 1532 2067
rect 1526 2062 1532 2063
rect 1654 2067 1660 2068
rect 1654 2063 1655 2067
rect 1659 2063 1660 2067
rect 1654 2062 1660 2063
rect 1732 2060 1734 2158
rect 1784 2141 1786 2165
rect 1866 2163 1872 2164
rect 1866 2159 1867 2163
rect 1871 2159 1872 2163
rect 1866 2158 1872 2159
rect 1782 2140 1788 2141
rect 1782 2136 1783 2140
rect 1787 2136 1788 2140
rect 1782 2135 1788 2136
rect 1868 2132 1870 2158
rect 1904 2141 1906 2165
rect 1902 2140 1908 2141
rect 1902 2136 1903 2140
rect 1907 2136 1908 2140
rect 2008 2138 2010 2165
rect 1902 2135 1908 2136
rect 2006 2137 2012 2138
rect 2006 2133 2007 2137
rect 2011 2133 2012 2137
rect 2048 2135 2050 2175
rect 2072 2135 2074 2176
rect 2176 2135 2178 2176
rect 2320 2135 2322 2176
rect 2006 2132 2012 2133
rect 2047 2134 2051 2135
rect 1850 2131 1856 2132
rect 1850 2127 1851 2131
rect 1855 2127 1856 2131
rect 1850 2126 1856 2127
rect 1866 2131 1872 2132
rect 1866 2127 1867 2131
rect 1871 2127 1872 2131
rect 2047 2129 2051 2130
rect 2071 2134 2075 2135
rect 2071 2129 2075 2130
rect 2175 2134 2179 2135
rect 2175 2129 2179 2130
rect 2279 2134 2283 2135
rect 2279 2129 2283 2130
rect 2319 2134 2323 2135
rect 2319 2129 2323 2130
rect 1866 2126 1872 2127
rect 1782 2121 1788 2122
rect 1782 2117 1783 2121
rect 1787 2117 1788 2121
rect 1782 2116 1788 2117
rect 1784 2095 1786 2116
rect 1783 2094 1787 2095
rect 1783 2089 1787 2090
rect 1791 2094 1795 2095
rect 1791 2089 1795 2090
rect 1792 2068 1794 2089
rect 1790 2067 1796 2068
rect 1790 2063 1791 2067
rect 1795 2063 1796 2067
rect 1790 2062 1796 2063
rect 1730 2059 1736 2060
rect 1330 2055 1336 2056
rect 1330 2051 1331 2055
rect 1335 2051 1336 2055
rect 1330 2050 1336 2051
rect 1602 2055 1608 2056
rect 1602 2051 1603 2055
rect 1607 2051 1608 2055
rect 1730 2055 1731 2059
rect 1735 2055 1736 2059
rect 1730 2054 1736 2055
rect 1602 2050 1608 2051
rect 1298 2027 1304 2028
rect 1298 2023 1299 2027
rect 1303 2023 1304 2027
rect 1298 2022 1304 2023
rect 111 2014 115 2015
rect 111 2009 115 2010
rect 447 2014 451 2015
rect 447 2009 451 2010
rect 575 2014 579 2015
rect 575 2009 579 2010
rect 623 2014 627 2015
rect 623 2009 627 2010
rect 727 2014 731 2015
rect 727 2009 731 2010
rect 735 2014 739 2015
rect 810 2014 816 2015
rect 855 2014 859 2015
rect 735 2009 739 2010
rect 112 1982 114 2009
rect 448 1985 450 2009
rect 514 2007 520 2008
rect 514 2003 515 2007
rect 519 2003 520 2007
rect 514 2002 520 2003
rect 522 2007 528 2008
rect 522 2003 523 2007
rect 527 2003 528 2007
rect 522 2002 528 2003
rect 446 1984 452 1985
rect 110 1981 116 1982
rect 110 1977 111 1981
rect 115 1977 116 1981
rect 446 1980 447 1984
rect 451 1980 452 1984
rect 446 1979 452 1980
rect 110 1976 116 1977
rect 446 1965 452 1966
rect 110 1964 116 1965
rect 110 1960 111 1964
rect 115 1960 116 1964
rect 446 1961 447 1965
rect 451 1961 452 1965
rect 446 1960 452 1961
rect 110 1959 116 1960
rect 112 1939 114 1959
rect 448 1939 450 1960
rect 111 1938 115 1939
rect 111 1933 115 1934
rect 447 1938 451 1939
rect 447 1933 451 1934
rect 112 1913 114 1933
rect 110 1912 116 1913
rect 110 1908 111 1912
rect 115 1908 116 1912
rect 110 1907 116 1908
rect 110 1895 116 1896
rect 110 1891 111 1895
rect 115 1891 116 1895
rect 110 1890 116 1891
rect 112 1863 114 1890
rect 111 1862 115 1863
rect 111 1857 115 1858
rect 319 1862 323 1863
rect 319 1857 323 1858
rect 447 1862 451 1863
rect 447 1857 451 1858
rect 112 1830 114 1857
rect 320 1833 322 1857
rect 330 1855 336 1856
rect 330 1851 331 1855
rect 335 1851 336 1855
rect 330 1850 336 1851
rect 394 1855 400 1856
rect 394 1851 395 1855
rect 399 1851 400 1855
rect 394 1850 400 1851
rect 318 1832 324 1833
rect 110 1829 116 1830
rect 110 1825 111 1829
rect 115 1825 116 1829
rect 318 1828 319 1832
rect 323 1828 324 1832
rect 318 1827 324 1828
rect 110 1824 116 1825
rect 318 1813 324 1814
rect 110 1812 116 1813
rect 110 1808 111 1812
rect 115 1808 116 1812
rect 318 1809 319 1813
rect 323 1809 324 1813
rect 318 1808 324 1809
rect 110 1807 116 1808
rect 112 1783 114 1807
rect 320 1783 322 1808
rect 111 1782 115 1783
rect 111 1777 115 1778
rect 255 1782 259 1783
rect 255 1777 259 1778
rect 319 1782 323 1783
rect 319 1777 323 1778
rect 112 1757 114 1777
rect 110 1756 116 1757
rect 256 1756 258 1777
rect 110 1752 111 1756
rect 115 1752 116 1756
rect 110 1751 116 1752
rect 254 1755 260 1756
rect 254 1751 255 1755
rect 259 1751 260 1755
rect 254 1750 260 1751
rect 332 1748 334 1850
rect 396 1824 398 1850
rect 448 1833 450 1857
rect 446 1832 452 1833
rect 446 1828 447 1832
rect 451 1828 452 1832
rect 446 1827 452 1828
rect 516 1824 518 2002
rect 524 1976 526 2002
rect 576 1985 578 2009
rect 650 2007 656 2008
rect 650 2003 651 2007
rect 655 2003 656 2007
rect 650 2002 656 2003
rect 574 1984 580 1985
rect 574 1980 575 1984
rect 579 1980 580 1984
rect 574 1979 580 1980
rect 652 1976 654 2002
rect 728 1985 730 2009
rect 802 2007 808 2008
rect 802 2003 803 2007
rect 807 2003 808 2007
rect 802 2002 808 2003
rect 726 1984 732 1985
rect 726 1980 727 1984
rect 731 1980 732 1984
rect 726 1979 732 1980
rect 804 1976 806 2002
rect 812 1976 814 2014
rect 855 2009 859 2010
rect 887 2014 891 2015
rect 887 2009 891 2010
rect 983 2014 987 2015
rect 983 2009 987 2010
rect 1055 2014 1059 2015
rect 1055 2009 1059 2010
rect 1119 2014 1123 2015
rect 1119 2009 1123 2010
rect 1231 2014 1235 2015
rect 1231 2009 1235 2010
rect 1255 2014 1259 2015
rect 1255 2009 1259 2010
rect 888 1985 890 2009
rect 1056 1985 1058 2009
rect 1106 2007 1112 2008
rect 1106 2003 1107 2007
rect 1111 2003 1112 2007
rect 1106 2002 1112 2003
rect 886 1984 892 1985
rect 886 1980 887 1984
rect 891 1980 892 1984
rect 886 1979 892 1980
rect 1054 1984 1060 1985
rect 1054 1980 1055 1984
rect 1059 1980 1060 1984
rect 1054 1979 1060 1980
rect 522 1975 528 1976
rect 522 1971 523 1975
rect 527 1971 528 1975
rect 522 1970 528 1971
rect 650 1975 656 1976
rect 650 1971 651 1975
rect 655 1971 656 1975
rect 650 1970 656 1971
rect 802 1975 808 1976
rect 802 1971 803 1975
rect 807 1971 808 1975
rect 802 1970 808 1971
rect 810 1975 816 1976
rect 810 1971 811 1975
rect 815 1971 816 1975
rect 810 1970 816 1971
rect 574 1965 580 1966
rect 574 1961 575 1965
rect 579 1961 580 1965
rect 574 1960 580 1961
rect 726 1965 732 1966
rect 726 1961 727 1965
rect 731 1961 732 1965
rect 726 1960 732 1961
rect 886 1965 892 1966
rect 886 1961 887 1965
rect 891 1961 892 1965
rect 886 1960 892 1961
rect 1054 1965 1060 1966
rect 1054 1961 1055 1965
rect 1059 1961 1060 1965
rect 1054 1960 1060 1961
rect 576 1939 578 1960
rect 728 1939 730 1960
rect 888 1939 890 1960
rect 1056 1939 1058 1960
rect 575 1938 579 1939
rect 575 1933 579 1934
rect 655 1938 659 1939
rect 655 1933 659 1934
rect 727 1938 731 1939
rect 727 1933 731 1934
rect 751 1938 755 1939
rect 751 1933 755 1934
rect 847 1938 851 1939
rect 847 1933 851 1934
rect 887 1938 891 1939
rect 887 1933 891 1934
rect 943 1938 947 1939
rect 943 1933 947 1934
rect 1039 1938 1043 1939
rect 1039 1933 1043 1934
rect 1055 1938 1059 1939
rect 1055 1933 1059 1934
rect 656 1912 658 1933
rect 752 1912 754 1933
rect 848 1912 850 1933
rect 944 1912 946 1933
rect 1040 1912 1042 1933
rect 654 1911 660 1912
rect 654 1907 655 1911
rect 659 1907 660 1911
rect 654 1906 660 1907
rect 750 1911 756 1912
rect 750 1907 751 1911
rect 755 1907 756 1911
rect 750 1906 756 1907
rect 846 1911 852 1912
rect 846 1907 847 1911
rect 851 1907 852 1911
rect 846 1906 852 1907
rect 942 1911 948 1912
rect 942 1907 943 1911
rect 947 1907 948 1911
rect 942 1906 948 1907
rect 1038 1911 1044 1912
rect 1038 1907 1039 1911
rect 1043 1907 1044 1911
rect 1108 1908 1110 2002
rect 1232 1985 1234 2009
rect 1332 2008 1334 2050
rect 1390 2048 1396 2049
rect 1390 2044 1391 2048
rect 1395 2044 1396 2048
rect 1390 2043 1396 2044
rect 1526 2048 1532 2049
rect 1526 2044 1527 2048
rect 1531 2044 1532 2048
rect 1526 2043 1532 2044
rect 1392 2015 1394 2043
rect 1466 2023 1472 2024
rect 1466 2019 1467 2023
rect 1471 2019 1472 2023
rect 1466 2018 1472 2019
rect 1391 2014 1395 2015
rect 1391 2009 1395 2010
rect 1399 2014 1403 2015
rect 1399 2009 1403 2010
rect 1330 2007 1336 2008
rect 1330 2003 1331 2007
rect 1335 2003 1336 2007
rect 1330 2002 1336 2003
rect 1400 1985 1402 2009
rect 1230 1984 1236 1985
rect 1230 1980 1231 1984
rect 1235 1980 1236 1984
rect 1230 1979 1236 1980
rect 1398 1984 1404 1985
rect 1398 1980 1399 1984
rect 1403 1980 1404 1984
rect 1398 1979 1404 1980
rect 1468 1976 1470 2018
rect 1528 2015 1530 2043
rect 1604 2028 1606 2050
rect 1654 2048 1660 2049
rect 1654 2044 1655 2048
rect 1659 2044 1660 2048
rect 1654 2043 1660 2044
rect 1790 2048 1796 2049
rect 1790 2044 1791 2048
rect 1795 2044 1796 2048
rect 1790 2043 1796 2044
rect 1602 2027 1608 2028
rect 1602 2023 1603 2027
rect 1607 2023 1608 2027
rect 1602 2022 1608 2023
rect 1656 2015 1658 2043
rect 1792 2015 1794 2043
rect 1852 2028 1854 2126
rect 1902 2121 1908 2122
rect 1902 2117 1903 2121
rect 1907 2117 1908 2121
rect 1902 2116 1908 2117
rect 2006 2120 2012 2121
rect 2006 2116 2007 2120
rect 2011 2116 2012 2120
rect 1904 2095 1906 2116
rect 2006 2115 2012 2116
rect 2008 2095 2010 2115
rect 2048 2109 2050 2129
rect 2046 2108 2052 2109
rect 2280 2108 2282 2129
rect 2046 2104 2047 2108
rect 2051 2104 2052 2108
rect 2046 2103 2052 2104
rect 2278 2107 2284 2108
rect 2278 2103 2279 2107
rect 2283 2103 2284 2107
rect 2278 2102 2284 2103
rect 2356 2100 2358 2218
rect 2396 2192 2398 2218
rect 2472 2201 2474 2225
rect 2546 2223 2552 2224
rect 2546 2219 2547 2223
rect 2551 2219 2552 2223
rect 2546 2218 2552 2219
rect 2470 2200 2476 2201
rect 2470 2196 2471 2200
rect 2475 2196 2476 2200
rect 2470 2195 2476 2196
rect 2548 2192 2550 2218
rect 2624 2201 2626 2225
rect 2622 2200 2628 2201
rect 2622 2196 2623 2200
rect 2627 2196 2628 2200
rect 2622 2195 2628 2196
rect 2700 2192 2702 2230
rect 2743 2225 2747 2226
rect 2783 2230 2787 2231
rect 2783 2225 2787 2226
rect 2784 2201 2786 2225
rect 2872 2224 2874 2266
rect 2892 2240 2894 2354
rect 3006 2349 3012 2350
rect 3006 2345 3007 2349
rect 3011 2345 3012 2349
rect 3006 2344 3012 2345
rect 3190 2349 3196 2350
rect 3190 2345 3191 2349
rect 3195 2345 3196 2349
rect 3190 2344 3196 2345
rect 3358 2349 3364 2350
rect 3358 2345 3359 2349
rect 3363 2345 3364 2349
rect 3358 2344 3364 2345
rect 3518 2349 3524 2350
rect 3518 2345 3519 2349
rect 3523 2345 3524 2349
rect 3518 2344 3524 2345
rect 3008 2307 3010 2344
rect 3192 2307 3194 2344
rect 3360 2307 3362 2344
rect 3520 2307 3522 2344
rect 2911 2306 2915 2307
rect 2911 2301 2915 2302
rect 3007 2306 3011 2307
rect 3007 2301 3011 2302
rect 3071 2306 3075 2307
rect 3071 2301 3075 2302
rect 3191 2306 3195 2307
rect 3191 2301 3195 2302
rect 3231 2306 3235 2307
rect 3231 2301 3235 2302
rect 3359 2306 3363 2307
rect 3359 2301 3363 2302
rect 3383 2306 3387 2307
rect 3383 2301 3387 2302
rect 3519 2306 3523 2307
rect 3519 2301 3523 2302
rect 3535 2306 3539 2307
rect 3535 2301 3539 2302
rect 2912 2280 2914 2301
rect 3072 2280 3074 2301
rect 3232 2280 3234 2301
rect 3384 2280 3386 2301
rect 3536 2280 3538 2301
rect 2910 2279 2916 2280
rect 2910 2275 2911 2279
rect 2915 2275 2916 2279
rect 2910 2274 2916 2275
rect 3070 2279 3076 2280
rect 3070 2275 3071 2279
rect 3075 2275 3076 2279
rect 3070 2274 3076 2275
rect 3230 2279 3236 2280
rect 3230 2275 3231 2279
rect 3235 2275 3236 2279
rect 3230 2274 3236 2275
rect 3382 2279 3388 2280
rect 3382 2275 3383 2279
rect 3387 2275 3388 2279
rect 3382 2274 3388 2275
rect 3534 2279 3540 2280
rect 3534 2275 3535 2279
rect 3539 2275 3540 2279
rect 3534 2274 3540 2275
rect 3620 2272 3622 2378
rect 3680 2369 3682 2393
rect 3754 2391 3760 2392
rect 3754 2387 3755 2391
rect 3759 2387 3760 2391
rect 3754 2386 3760 2387
rect 3678 2368 3684 2369
rect 3678 2364 3679 2368
rect 3683 2364 3684 2368
rect 3678 2363 3684 2364
rect 3756 2360 3758 2386
rect 3840 2369 3842 2393
rect 3838 2368 3844 2369
rect 3838 2364 3839 2368
rect 3843 2364 3844 2368
rect 3838 2363 3844 2364
rect 3908 2360 3910 2410
rect 3944 2399 3946 2438
rect 3943 2398 3947 2399
rect 3943 2393 3947 2394
rect 3944 2366 3946 2393
rect 3942 2365 3948 2366
rect 3942 2361 3943 2365
rect 3947 2361 3948 2365
rect 3942 2360 3948 2361
rect 3754 2359 3760 2360
rect 3754 2355 3755 2359
rect 3759 2355 3760 2359
rect 3754 2354 3760 2355
rect 3906 2359 3912 2360
rect 3906 2355 3907 2359
rect 3911 2355 3912 2359
rect 3906 2354 3912 2355
rect 3678 2349 3684 2350
rect 3678 2345 3679 2349
rect 3683 2345 3684 2349
rect 3678 2344 3684 2345
rect 3838 2349 3844 2350
rect 3838 2345 3839 2349
rect 3843 2345 3844 2349
rect 3838 2344 3844 2345
rect 3942 2348 3948 2349
rect 3942 2344 3943 2348
rect 3947 2344 3948 2348
rect 3680 2307 3682 2344
rect 3840 2307 3842 2344
rect 3942 2343 3948 2344
rect 3944 2307 3946 2343
rect 3679 2306 3683 2307
rect 3679 2301 3683 2302
rect 3695 2306 3699 2307
rect 3695 2301 3699 2302
rect 3839 2306 3843 2307
rect 3839 2301 3843 2302
rect 3943 2306 3947 2307
rect 3943 2301 3947 2302
rect 3696 2280 3698 2301
rect 3944 2281 3946 2301
rect 3942 2280 3948 2281
rect 3694 2279 3700 2280
rect 3694 2275 3695 2279
rect 3699 2275 3700 2279
rect 3942 2276 3943 2280
rect 3947 2276 3948 2280
rect 3942 2275 3948 2276
rect 3694 2274 3700 2275
rect 3618 2271 3624 2272
rect 3146 2267 3152 2268
rect 3146 2263 3147 2267
rect 3151 2263 3152 2267
rect 3146 2262 3152 2263
rect 3306 2267 3312 2268
rect 3306 2263 3307 2267
rect 3311 2263 3312 2267
rect 3306 2262 3312 2263
rect 3458 2267 3464 2268
rect 3458 2263 3459 2267
rect 3463 2263 3464 2267
rect 3458 2262 3464 2263
rect 3610 2267 3616 2268
rect 3610 2263 3611 2267
rect 3615 2263 3616 2267
rect 3618 2267 3619 2271
rect 3623 2267 3624 2271
rect 3618 2266 3624 2267
rect 3610 2262 3616 2263
rect 3942 2263 3948 2264
rect 2910 2260 2916 2261
rect 2910 2256 2911 2260
rect 2915 2256 2916 2260
rect 2910 2255 2916 2256
rect 3070 2260 3076 2261
rect 3070 2256 3071 2260
rect 3075 2256 3076 2260
rect 3070 2255 3076 2256
rect 2890 2239 2896 2240
rect 2890 2235 2891 2239
rect 2895 2235 2896 2239
rect 2890 2234 2896 2235
rect 2912 2231 2914 2255
rect 3072 2231 3074 2255
rect 3148 2240 3150 2262
rect 3230 2260 3236 2261
rect 3230 2256 3231 2260
rect 3235 2256 3236 2260
rect 3230 2255 3236 2256
rect 3146 2239 3152 2240
rect 3146 2235 3147 2239
rect 3151 2235 3152 2239
rect 3146 2234 3152 2235
rect 3232 2231 3234 2255
rect 3308 2240 3310 2262
rect 3382 2260 3388 2261
rect 3382 2256 3383 2260
rect 3387 2256 3388 2260
rect 3382 2255 3388 2256
rect 3306 2239 3312 2240
rect 3306 2235 3307 2239
rect 3311 2235 3312 2239
rect 3306 2234 3312 2235
rect 3384 2231 3386 2255
rect 3450 2247 3456 2248
rect 3450 2243 3451 2247
rect 3455 2243 3456 2247
rect 3450 2242 3456 2243
rect 2911 2230 2915 2231
rect 2911 2225 2915 2226
rect 2935 2230 2939 2231
rect 2935 2225 2939 2226
rect 3071 2230 3075 2231
rect 3071 2225 3075 2226
rect 3079 2230 3083 2231
rect 3079 2225 3083 2226
rect 3223 2230 3227 2231
rect 3223 2225 3227 2226
rect 3231 2230 3235 2231
rect 3231 2225 3235 2226
rect 3367 2230 3371 2231
rect 3367 2225 3371 2226
rect 3383 2230 3387 2231
rect 3383 2225 3387 2226
rect 2870 2223 2876 2224
rect 2870 2219 2871 2223
rect 2875 2219 2876 2223
rect 2870 2218 2876 2219
rect 2936 2201 2938 2225
rect 2990 2223 2996 2224
rect 2990 2219 2991 2223
rect 2995 2219 2996 2223
rect 2990 2218 2996 2219
rect 3010 2223 3016 2224
rect 3010 2219 3011 2223
rect 3015 2219 3016 2223
rect 3010 2218 3016 2219
rect 2782 2200 2788 2201
rect 2782 2196 2783 2200
rect 2787 2196 2788 2200
rect 2782 2195 2788 2196
rect 2934 2200 2940 2201
rect 2934 2196 2935 2200
rect 2939 2196 2940 2200
rect 2934 2195 2940 2196
rect 2394 2191 2400 2192
rect 2394 2187 2395 2191
rect 2399 2187 2400 2191
rect 2394 2186 2400 2187
rect 2546 2191 2552 2192
rect 2546 2187 2547 2191
rect 2551 2187 2552 2191
rect 2546 2186 2552 2187
rect 2698 2191 2704 2192
rect 2698 2187 2699 2191
rect 2703 2187 2704 2191
rect 2698 2186 2704 2187
rect 2850 2191 2856 2192
rect 2850 2187 2851 2191
rect 2855 2187 2856 2191
rect 2850 2186 2856 2187
rect 2470 2181 2476 2182
rect 2470 2177 2471 2181
rect 2475 2177 2476 2181
rect 2470 2176 2476 2177
rect 2622 2181 2628 2182
rect 2622 2177 2623 2181
rect 2627 2177 2628 2181
rect 2622 2176 2628 2177
rect 2782 2181 2788 2182
rect 2782 2177 2783 2181
rect 2787 2177 2788 2181
rect 2782 2176 2788 2177
rect 2472 2135 2474 2176
rect 2624 2135 2626 2176
rect 2784 2135 2786 2176
rect 2391 2134 2395 2135
rect 2391 2129 2395 2130
rect 2471 2134 2475 2135
rect 2471 2129 2475 2130
rect 2511 2134 2515 2135
rect 2511 2129 2515 2130
rect 2623 2134 2627 2135
rect 2623 2129 2627 2130
rect 2631 2134 2635 2135
rect 2631 2129 2635 2130
rect 2759 2134 2763 2135
rect 2759 2129 2763 2130
rect 2783 2134 2787 2135
rect 2783 2129 2787 2130
rect 2392 2108 2394 2129
rect 2512 2108 2514 2129
rect 2632 2108 2634 2129
rect 2760 2108 2762 2129
rect 2390 2107 2396 2108
rect 2390 2103 2391 2107
rect 2395 2103 2396 2107
rect 2390 2102 2396 2103
rect 2510 2107 2516 2108
rect 2510 2103 2511 2107
rect 2515 2103 2516 2107
rect 2510 2102 2516 2103
rect 2630 2107 2636 2108
rect 2630 2103 2631 2107
rect 2635 2103 2636 2107
rect 2630 2102 2636 2103
rect 2758 2107 2764 2108
rect 2758 2103 2759 2107
rect 2763 2103 2764 2107
rect 2758 2102 2764 2103
rect 2354 2099 2360 2100
rect 2354 2095 2355 2099
rect 2359 2095 2360 2099
rect 1903 2094 1907 2095
rect 1903 2089 1907 2090
rect 2007 2094 2011 2095
rect 2354 2094 2360 2095
rect 2382 2099 2388 2100
rect 2382 2095 2383 2099
rect 2387 2095 2388 2099
rect 2382 2094 2388 2095
rect 2498 2099 2504 2100
rect 2498 2095 2499 2099
rect 2503 2095 2504 2099
rect 2498 2094 2504 2095
rect 2706 2095 2712 2096
rect 2007 2089 2011 2090
rect 2046 2091 2052 2092
rect 1904 2068 1906 2089
rect 2008 2069 2010 2089
rect 2046 2087 2047 2091
rect 2051 2087 2052 2091
rect 2046 2086 2052 2087
rect 2278 2088 2284 2089
rect 2006 2068 2012 2069
rect 1902 2067 1908 2068
rect 1902 2063 1903 2067
rect 1907 2063 1908 2067
rect 2006 2064 2007 2068
rect 2011 2064 2012 2068
rect 2006 2063 2012 2064
rect 1902 2062 1908 2063
rect 1866 2055 1872 2056
rect 1866 2051 1867 2055
rect 1871 2051 1872 2055
rect 1866 2050 1872 2051
rect 1978 2055 1984 2056
rect 1978 2051 1979 2055
rect 1983 2051 1984 2055
rect 1978 2050 1984 2051
rect 2006 2051 2012 2052
rect 2048 2051 2050 2086
rect 2278 2084 2279 2088
rect 2283 2084 2284 2088
rect 2278 2083 2284 2084
rect 2280 2051 2282 2083
rect 2384 2068 2386 2094
rect 2390 2088 2396 2089
rect 2390 2084 2391 2088
rect 2395 2084 2396 2088
rect 2390 2083 2396 2084
rect 2382 2067 2388 2068
rect 2382 2063 2383 2067
rect 2387 2063 2388 2067
rect 2382 2062 2388 2063
rect 2392 2051 2394 2083
rect 2500 2068 2502 2094
rect 2706 2091 2707 2095
rect 2711 2091 2712 2095
rect 2706 2090 2712 2091
rect 2510 2088 2516 2089
rect 2510 2084 2511 2088
rect 2515 2084 2516 2088
rect 2510 2083 2516 2084
rect 2630 2088 2636 2089
rect 2630 2084 2631 2088
rect 2635 2084 2636 2088
rect 2630 2083 2636 2084
rect 2498 2067 2504 2068
rect 2498 2063 2499 2067
rect 2503 2063 2504 2067
rect 2498 2062 2504 2063
rect 2512 2051 2514 2083
rect 2518 2063 2524 2064
rect 2518 2059 2519 2063
rect 2523 2059 2524 2063
rect 2518 2058 2524 2059
rect 1868 2028 1870 2050
rect 1902 2048 1908 2049
rect 1902 2044 1903 2048
rect 1907 2044 1908 2048
rect 1902 2043 1908 2044
rect 1846 2027 1854 2028
rect 1846 2023 1847 2027
rect 1851 2025 1854 2027
rect 1866 2027 1872 2028
rect 1851 2023 1852 2025
rect 1846 2022 1852 2023
rect 1866 2023 1867 2027
rect 1871 2023 1872 2027
rect 1866 2022 1872 2023
rect 1904 2015 1906 2043
rect 1527 2014 1531 2015
rect 1527 2009 1531 2010
rect 1575 2014 1579 2015
rect 1575 2009 1579 2010
rect 1655 2014 1659 2015
rect 1655 2009 1659 2010
rect 1751 2014 1755 2015
rect 1751 2009 1755 2010
rect 1791 2014 1795 2015
rect 1791 2009 1795 2010
rect 1903 2014 1907 2015
rect 1903 2009 1907 2010
rect 1486 2007 1492 2008
rect 1486 2003 1487 2007
rect 1491 2003 1492 2007
rect 1486 2002 1492 2003
rect 1488 1976 1490 2002
rect 1576 1985 1578 2009
rect 1662 2007 1668 2008
rect 1662 2003 1663 2007
rect 1667 2003 1668 2007
rect 1662 2002 1668 2003
rect 1574 1984 1580 1985
rect 1574 1980 1575 1984
rect 1579 1980 1580 1984
rect 1574 1979 1580 1980
rect 1664 1976 1666 2002
rect 1752 1985 1754 2009
rect 1834 2007 1840 2008
rect 1834 2003 1835 2007
rect 1839 2003 1840 2007
rect 1834 2002 1840 2003
rect 1750 1984 1756 1985
rect 1750 1980 1751 1984
rect 1755 1980 1756 1984
rect 1750 1979 1756 1980
rect 1836 1976 1838 2002
rect 1904 1985 1906 2009
rect 1980 2008 1982 2050
rect 2006 2047 2007 2051
rect 2011 2047 2012 2051
rect 2006 2046 2012 2047
rect 2047 2050 2051 2051
rect 2008 2015 2010 2046
rect 2047 2045 2051 2046
rect 2279 2050 2283 2051
rect 2279 2045 2283 2046
rect 2327 2050 2331 2051
rect 2327 2045 2331 2046
rect 2391 2050 2395 2051
rect 2391 2045 2395 2046
rect 2431 2050 2435 2051
rect 2431 2045 2435 2046
rect 2511 2050 2515 2051
rect 2511 2045 2515 2046
rect 2048 2018 2050 2045
rect 2328 2021 2330 2045
rect 2402 2043 2408 2044
rect 2402 2039 2403 2043
rect 2407 2039 2408 2043
rect 2402 2038 2408 2039
rect 2326 2020 2332 2021
rect 2046 2017 2052 2018
rect 2007 2014 2011 2015
rect 2046 2013 2047 2017
rect 2051 2013 2052 2017
rect 2326 2016 2327 2020
rect 2331 2016 2332 2020
rect 2326 2015 2332 2016
rect 2046 2012 2052 2013
rect 2404 2012 2406 2038
rect 2432 2021 2434 2045
rect 2430 2020 2436 2021
rect 2430 2016 2431 2020
rect 2435 2016 2436 2020
rect 2430 2015 2436 2016
rect 2520 2012 2522 2058
rect 2632 2051 2634 2083
rect 2535 2050 2539 2051
rect 2535 2045 2539 2046
rect 2631 2050 2635 2051
rect 2631 2045 2635 2046
rect 2647 2050 2651 2051
rect 2647 2045 2651 2046
rect 2526 2035 2532 2036
rect 2526 2031 2527 2035
rect 2531 2031 2532 2035
rect 2526 2030 2532 2031
rect 2528 2012 2530 2030
rect 2536 2021 2538 2045
rect 2618 2043 2624 2044
rect 2618 2039 2619 2043
rect 2623 2039 2624 2043
rect 2618 2038 2624 2039
rect 2534 2020 2540 2021
rect 2534 2016 2535 2020
rect 2539 2016 2540 2020
rect 2534 2015 2540 2016
rect 2007 2009 2011 2010
rect 2402 2011 2408 2012
rect 1978 2007 1984 2008
rect 1978 2003 1979 2007
rect 1983 2003 1984 2007
rect 1978 2002 1984 2003
rect 1902 1984 1908 1985
rect 1902 1980 1903 1984
rect 1907 1980 1908 1984
rect 2008 1982 2010 2009
rect 2402 2007 2403 2011
rect 2407 2007 2408 2011
rect 2402 2006 2408 2007
rect 2518 2011 2524 2012
rect 2518 2007 2519 2011
rect 2523 2007 2524 2011
rect 2518 2006 2524 2007
rect 2526 2011 2532 2012
rect 2526 2007 2527 2011
rect 2531 2007 2532 2011
rect 2526 2006 2532 2007
rect 2326 2001 2332 2002
rect 2046 2000 2052 2001
rect 2046 1996 2047 2000
rect 2051 1996 2052 2000
rect 2326 1997 2327 2001
rect 2331 1997 2332 2001
rect 2326 1996 2332 1997
rect 2430 2001 2436 2002
rect 2430 1997 2431 2001
rect 2435 1997 2436 2001
rect 2430 1996 2436 1997
rect 2534 2001 2540 2002
rect 2534 1997 2535 2001
rect 2539 1997 2540 2001
rect 2534 1996 2540 1997
rect 2046 1995 2052 1996
rect 1902 1979 1908 1980
rect 2006 1981 2012 1982
rect 2006 1977 2007 1981
rect 2011 1977 2012 1981
rect 2006 1976 2012 1977
rect 1122 1975 1128 1976
rect 1122 1971 1123 1975
rect 1127 1971 1128 1975
rect 1122 1970 1128 1971
rect 1202 1975 1208 1976
rect 1202 1971 1203 1975
rect 1207 1971 1208 1975
rect 1202 1970 1208 1971
rect 1466 1975 1472 1976
rect 1466 1971 1467 1975
rect 1471 1971 1472 1975
rect 1466 1970 1472 1971
rect 1486 1975 1492 1976
rect 1486 1971 1487 1975
rect 1491 1971 1492 1975
rect 1486 1970 1492 1971
rect 1662 1975 1668 1976
rect 1662 1971 1663 1975
rect 1667 1971 1668 1975
rect 1662 1970 1668 1971
rect 1834 1975 1840 1976
rect 1834 1971 1835 1975
rect 1839 1971 1840 1975
rect 2048 1971 2050 1995
rect 2328 1971 2330 1996
rect 2432 1971 2434 1996
rect 2536 1971 2538 1996
rect 1834 1970 1840 1971
rect 2047 1970 2051 1971
rect 1038 1906 1044 1907
rect 1106 1907 1112 1908
rect 738 1903 744 1904
rect 738 1899 739 1903
rect 743 1899 744 1903
rect 738 1898 744 1899
rect 930 1903 936 1904
rect 930 1899 931 1903
rect 935 1899 936 1903
rect 1106 1903 1107 1907
rect 1111 1903 1112 1907
rect 1106 1902 1112 1903
rect 930 1898 936 1899
rect 654 1892 660 1893
rect 654 1888 655 1892
rect 659 1888 660 1892
rect 654 1887 660 1888
rect 656 1863 658 1887
rect 740 1872 742 1898
rect 750 1892 756 1893
rect 750 1888 751 1892
rect 755 1888 756 1892
rect 750 1887 756 1888
rect 846 1892 852 1893
rect 846 1888 847 1892
rect 851 1888 852 1892
rect 846 1887 852 1888
rect 738 1871 744 1872
rect 738 1867 739 1871
rect 743 1867 744 1871
rect 738 1866 744 1867
rect 752 1863 754 1887
rect 848 1863 850 1887
rect 932 1872 934 1898
rect 942 1892 948 1893
rect 942 1888 943 1892
rect 947 1888 948 1892
rect 942 1887 948 1888
rect 1038 1892 1044 1893
rect 1038 1888 1039 1892
rect 1043 1888 1044 1892
rect 1038 1887 1044 1888
rect 930 1871 936 1872
rect 930 1867 931 1871
rect 935 1867 936 1871
rect 930 1866 936 1867
rect 944 1863 946 1887
rect 1040 1863 1042 1887
rect 1124 1872 1126 1970
rect 1135 1938 1139 1939
rect 1135 1933 1139 1934
rect 1136 1912 1138 1933
rect 1134 1911 1140 1912
rect 1134 1907 1135 1911
rect 1139 1907 1140 1911
rect 1134 1906 1140 1907
rect 1134 1892 1140 1893
rect 1134 1888 1135 1892
rect 1139 1888 1140 1892
rect 1134 1887 1140 1888
rect 1122 1871 1128 1872
rect 1122 1867 1123 1871
rect 1127 1867 1128 1871
rect 1122 1866 1128 1867
rect 1136 1863 1138 1887
rect 1204 1872 1206 1970
rect 1230 1965 1236 1966
rect 1230 1961 1231 1965
rect 1235 1961 1236 1965
rect 1230 1960 1236 1961
rect 1398 1965 1404 1966
rect 1398 1961 1399 1965
rect 1403 1961 1404 1965
rect 1398 1960 1404 1961
rect 1574 1965 1580 1966
rect 1574 1961 1575 1965
rect 1579 1961 1580 1965
rect 1574 1960 1580 1961
rect 1750 1965 1756 1966
rect 1750 1961 1751 1965
rect 1755 1961 1756 1965
rect 1750 1960 1756 1961
rect 1902 1965 1908 1966
rect 2047 1965 2051 1966
rect 2255 1970 2259 1971
rect 2255 1965 2259 1966
rect 2327 1970 2331 1971
rect 2327 1965 2331 1966
rect 2351 1970 2355 1971
rect 2351 1965 2355 1966
rect 2431 1970 2435 1971
rect 2431 1965 2435 1966
rect 2447 1970 2451 1971
rect 2447 1965 2451 1966
rect 2535 1970 2539 1971
rect 2535 1965 2539 1966
rect 2543 1970 2547 1971
rect 2543 1965 2547 1966
rect 1902 1961 1903 1965
rect 1907 1961 1908 1965
rect 1902 1960 1908 1961
rect 2006 1964 2012 1965
rect 2006 1960 2007 1964
rect 2011 1960 2012 1964
rect 1232 1939 1234 1960
rect 1400 1939 1402 1960
rect 1576 1939 1578 1960
rect 1752 1939 1754 1960
rect 1904 1939 1906 1960
rect 2006 1959 2012 1960
rect 2008 1939 2010 1959
rect 2048 1945 2050 1965
rect 2046 1944 2052 1945
rect 2256 1944 2258 1965
rect 2352 1944 2354 1965
rect 2448 1944 2450 1965
rect 2544 1944 2546 1965
rect 2046 1940 2047 1944
rect 2051 1940 2052 1944
rect 2046 1939 2052 1940
rect 2254 1943 2260 1944
rect 2254 1939 2255 1943
rect 2259 1939 2260 1943
rect 1231 1938 1235 1939
rect 1231 1933 1235 1934
rect 1327 1938 1331 1939
rect 1327 1933 1331 1934
rect 1399 1938 1403 1939
rect 1399 1933 1403 1934
rect 1423 1938 1427 1939
rect 1423 1933 1427 1934
rect 1575 1938 1579 1939
rect 1575 1933 1579 1934
rect 1751 1938 1755 1939
rect 1751 1933 1755 1934
rect 1903 1938 1907 1939
rect 1903 1933 1907 1934
rect 2007 1938 2011 1939
rect 2254 1938 2260 1939
rect 2350 1943 2356 1944
rect 2350 1939 2351 1943
rect 2355 1939 2356 1943
rect 2350 1938 2356 1939
rect 2446 1943 2452 1944
rect 2446 1939 2447 1943
rect 2451 1939 2452 1943
rect 2446 1938 2452 1939
rect 2542 1943 2548 1944
rect 2542 1939 2543 1943
rect 2547 1939 2548 1943
rect 2542 1938 2548 1939
rect 2620 1936 2622 2038
rect 2648 2021 2650 2045
rect 2708 2044 2710 2090
rect 2758 2088 2764 2089
rect 2758 2084 2759 2088
rect 2763 2084 2764 2088
rect 2758 2083 2764 2084
rect 2760 2051 2762 2083
rect 2852 2068 2854 2186
rect 2934 2181 2940 2182
rect 2934 2177 2935 2181
rect 2939 2177 2940 2181
rect 2934 2176 2940 2177
rect 2936 2135 2938 2176
rect 2895 2134 2899 2135
rect 2895 2129 2899 2130
rect 2935 2134 2939 2135
rect 2935 2129 2939 2130
rect 2896 2108 2898 2129
rect 2992 2116 2994 2218
rect 3012 2192 3014 2218
rect 3080 2201 3082 2225
rect 3154 2223 3160 2224
rect 3154 2219 3155 2223
rect 3159 2219 3160 2223
rect 3154 2218 3160 2219
rect 3078 2200 3084 2201
rect 3078 2196 3079 2200
rect 3083 2196 3084 2200
rect 3078 2195 3084 2196
rect 3156 2192 3158 2218
rect 3224 2201 3226 2225
rect 3298 2223 3304 2224
rect 3298 2219 3299 2223
rect 3303 2219 3304 2223
rect 3298 2218 3304 2219
rect 3222 2200 3228 2201
rect 3222 2196 3223 2200
rect 3227 2196 3228 2200
rect 3222 2195 3228 2196
rect 3300 2192 3302 2218
rect 3368 2201 3370 2225
rect 3442 2223 3448 2224
rect 3442 2219 3443 2223
rect 3447 2219 3448 2223
rect 3442 2218 3448 2219
rect 3366 2200 3372 2201
rect 3366 2196 3367 2200
rect 3371 2196 3372 2200
rect 3366 2195 3372 2196
rect 3444 2192 3446 2218
rect 3452 2192 3454 2242
rect 3460 2240 3462 2262
rect 3534 2260 3540 2261
rect 3534 2256 3535 2260
rect 3539 2256 3540 2260
rect 3534 2255 3540 2256
rect 3458 2239 3464 2240
rect 3458 2235 3459 2239
rect 3463 2235 3464 2239
rect 3458 2234 3464 2235
rect 3536 2231 3538 2255
rect 3612 2240 3614 2262
rect 3694 2260 3700 2261
rect 3694 2256 3695 2260
rect 3699 2256 3700 2260
rect 3942 2259 3943 2263
rect 3947 2259 3948 2263
rect 3942 2258 3948 2259
rect 3694 2255 3700 2256
rect 3610 2239 3616 2240
rect 3610 2235 3611 2239
rect 3615 2235 3616 2239
rect 3610 2234 3616 2235
rect 3696 2231 3698 2255
rect 3944 2231 3946 2258
rect 3519 2230 3523 2231
rect 3519 2225 3523 2226
rect 3535 2230 3539 2231
rect 3535 2225 3539 2226
rect 3695 2230 3699 2231
rect 3695 2225 3699 2226
rect 3943 2230 3947 2231
rect 3943 2225 3947 2226
rect 3520 2201 3522 2225
rect 3518 2200 3524 2201
rect 3518 2196 3519 2200
rect 3523 2196 3524 2200
rect 3944 2198 3946 2225
rect 3518 2195 3524 2196
rect 3942 2197 3948 2198
rect 3942 2193 3943 2197
rect 3947 2193 3948 2197
rect 3942 2192 3948 2193
rect 3010 2191 3016 2192
rect 3010 2187 3011 2191
rect 3015 2187 3016 2191
rect 3010 2186 3016 2187
rect 3154 2191 3160 2192
rect 3154 2187 3155 2191
rect 3159 2187 3160 2191
rect 3154 2186 3160 2187
rect 3298 2191 3304 2192
rect 3298 2187 3299 2191
rect 3303 2187 3304 2191
rect 3298 2186 3304 2187
rect 3442 2191 3448 2192
rect 3442 2187 3443 2191
rect 3447 2187 3448 2191
rect 3442 2186 3448 2187
rect 3450 2191 3456 2192
rect 3450 2187 3451 2191
rect 3455 2187 3456 2191
rect 3450 2186 3456 2187
rect 3078 2181 3084 2182
rect 3078 2177 3079 2181
rect 3083 2177 3084 2181
rect 3078 2176 3084 2177
rect 3222 2181 3228 2182
rect 3222 2177 3223 2181
rect 3227 2177 3228 2181
rect 3222 2176 3228 2177
rect 3366 2181 3372 2182
rect 3366 2177 3367 2181
rect 3371 2177 3372 2181
rect 3366 2176 3372 2177
rect 3518 2181 3524 2182
rect 3518 2177 3519 2181
rect 3523 2177 3524 2181
rect 3518 2176 3524 2177
rect 3942 2180 3948 2181
rect 3942 2176 3943 2180
rect 3947 2176 3948 2180
rect 3080 2135 3082 2176
rect 3224 2135 3226 2176
rect 3368 2135 3370 2176
rect 3520 2135 3522 2176
rect 3942 2175 3948 2176
rect 3944 2135 3946 2175
rect 3039 2134 3043 2135
rect 3039 2129 3043 2130
rect 3079 2134 3083 2135
rect 3079 2129 3083 2130
rect 3191 2134 3195 2135
rect 3191 2129 3195 2130
rect 3223 2134 3227 2135
rect 3223 2129 3227 2130
rect 3351 2134 3355 2135
rect 3351 2129 3355 2130
rect 3367 2134 3371 2135
rect 3367 2129 3371 2130
rect 3519 2134 3523 2135
rect 3519 2129 3523 2130
rect 3687 2134 3691 2135
rect 3687 2129 3691 2130
rect 3839 2134 3843 2135
rect 3839 2129 3843 2130
rect 3943 2134 3947 2135
rect 3943 2129 3947 2130
rect 2990 2115 2996 2116
rect 2990 2111 2991 2115
rect 2995 2111 2996 2115
rect 2990 2110 2996 2111
rect 3040 2108 3042 2129
rect 3192 2108 3194 2129
rect 3352 2108 3354 2129
rect 3520 2108 3522 2129
rect 3688 2108 3690 2129
rect 3840 2108 3842 2129
rect 3944 2109 3946 2129
rect 3942 2108 3948 2109
rect 2894 2107 2900 2108
rect 2894 2103 2895 2107
rect 2899 2103 2900 2107
rect 2894 2102 2900 2103
rect 3038 2107 3044 2108
rect 3038 2103 3039 2107
rect 3043 2103 3044 2107
rect 3038 2102 3044 2103
rect 3190 2107 3196 2108
rect 3190 2103 3191 2107
rect 3195 2103 3196 2107
rect 3190 2102 3196 2103
rect 3350 2107 3356 2108
rect 3350 2103 3351 2107
rect 3355 2103 3356 2107
rect 3350 2102 3356 2103
rect 3518 2107 3524 2108
rect 3518 2103 3519 2107
rect 3523 2103 3524 2107
rect 3518 2102 3524 2103
rect 3686 2107 3692 2108
rect 3686 2103 3687 2107
rect 3691 2103 3692 2107
rect 3686 2102 3692 2103
rect 3838 2107 3844 2108
rect 3838 2103 3839 2107
rect 3843 2103 3844 2107
rect 3942 2104 3943 2108
rect 3947 2104 3948 2108
rect 3942 2103 3948 2104
rect 3838 2102 3844 2103
rect 3830 2099 3836 2100
rect 2970 2095 2976 2096
rect 2970 2091 2971 2095
rect 2975 2091 2976 2095
rect 2970 2090 2976 2091
rect 3114 2095 3120 2096
rect 3114 2091 3115 2095
rect 3119 2091 3120 2095
rect 3114 2090 3120 2091
rect 3266 2095 3272 2096
rect 3266 2091 3267 2095
rect 3271 2091 3272 2095
rect 3266 2090 3272 2091
rect 3426 2095 3432 2096
rect 3426 2091 3427 2095
rect 3431 2091 3432 2095
rect 3426 2090 3432 2091
rect 3762 2095 3768 2096
rect 3762 2091 3763 2095
rect 3767 2091 3768 2095
rect 3830 2095 3831 2099
rect 3835 2095 3836 2099
rect 3830 2094 3836 2095
rect 3762 2090 3768 2091
rect 2894 2088 2900 2089
rect 2894 2084 2895 2088
rect 2899 2084 2900 2088
rect 2894 2083 2900 2084
rect 2850 2067 2856 2068
rect 2850 2063 2851 2067
rect 2855 2063 2856 2067
rect 2850 2062 2856 2063
rect 2896 2051 2898 2083
rect 2972 2068 2974 2090
rect 3038 2088 3044 2089
rect 3038 2084 3039 2088
rect 3043 2084 3044 2088
rect 3038 2083 3044 2084
rect 2970 2067 2976 2068
rect 2970 2063 2971 2067
rect 2975 2063 2976 2067
rect 2970 2062 2976 2063
rect 3040 2051 3042 2083
rect 3116 2068 3118 2090
rect 3190 2088 3196 2089
rect 3190 2084 3191 2088
rect 3195 2084 3196 2088
rect 3190 2083 3196 2084
rect 3114 2067 3120 2068
rect 3114 2063 3115 2067
rect 3119 2063 3120 2067
rect 3114 2062 3120 2063
rect 3192 2051 3194 2083
rect 3268 2068 3270 2090
rect 3350 2088 3356 2089
rect 3350 2084 3351 2088
rect 3355 2084 3356 2088
rect 3350 2083 3356 2084
rect 3266 2067 3272 2068
rect 3266 2063 3267 2067
rect 3271 2063 3272 2067
rect 3266 2062 3272 2063
rect 3352 2051 3354 2083
rect 3428 2068 3430 2090
rect 3518 2088 3524 2089
rect 3518 2084 3519 2088
rect 3523 2084 3524 2088
rect 3518 2083 3524 2084
rect 3686 2088 3692 2089
rect 3686 2084 3687 2088
rect 3691 2084 3692 2088
rect 3686 2083 3692 2084
rect 3426 2067 3432 2068
rect 3426 2063 3427 2067
rect 3431 2063 3432 2067
rect 3426 2062 3432 2063
rect 3378 2059 3384 2060
rect 3378 2055 3379 2059
rect 3383 2055 3384 2059
rect 3378 2054 3384 2055
rect 2759 2050 2763 2051
rect 2759 2045 2763 2046
rect 2775 2050 2779 2051
rect 2775 2045 2779 2046
rect 2895 2050 2899 2051
rect 2895 2045 2899 2046
rect 2919 2050 2923 2051
rect 2919 2045 2923 2046
rect 3039 2050 3043 2051
rect 3039 2045 3043 2046
rect 3079 2050 3083 2051
rect 3079 2045 3083 2046
rect 3191 2050 3195 2051
rect 3191 2045 3195 2046
rect 3263 2050 3267 2051
rect 3263 2045 3267 2046
rect 3351 2050 3355 2051
rect 3351 2045 3355 2046
rect 2702 2043 2710 2044
rect 2702 2039 2703 2043
rect 2707 2040 2710 2043
rect 2707 2039 2708 2040
rect 2702 2038 2708 2039
rect 2776 2021 2778 2045
rect 2842 2043 2848 2044
rect 2842 2039 2843 2043
rect 2847 2039 2848 2043
rect 2842 2038 2848 2039
rect 2850 2043 2856 2044
rect 2850 2039 2851 2043
rect 2855 2039 2856 2043
rect 2850 2038 2856 2039
rect 2646 2020 2652 2021
rect 2646 2016 2647 2020
rect 2651 2016 2652 2020
rect 2646 2015 2652 2016
rect 2774 2020 2780 2021
rect 2774 2016 2775 2020
rect 2779 2016 2780 2020
rect 2774 2015 2780 2016
rect 2714 2011 2720 2012
rect 2714 2007 2715 2011
rect 2719 2007 2720 2011
rect 2714 2006 2720 2007
rect 2646 2001 2652 2002
rect 2646 1997 2647 2001
rect 2651 1997 2652 2001
rect 2646 1996 2652 1997
rect 2648 1971 2650 1996
rect 2647 1970 2651 1971
rect 2647 1965 2651 1966
rect 2648 1944 2650 1965
rect 2646 1943 2652 1944
rect 2646 1939 2647 1943
rect 2651 1939 2652 1943
rect 2646 1938 2652 1939
rect 2007 1933 2011 1934
rect 2618 1935 2624 1936
rect 1232 1912 1234 1933
rect 1328 1912 1330 1933
rect 1424 1912 1426 1933
rect 2008 1913 2010 1933
rect 2330 1931 2336 1932
rect 2046 1927 2052 1928
rect 2046 1923 2047 1927
rect 2051 1923 2052 1927
rect 2330 1927 2331 1931
rect 2335 1927 2336 1931
rect 2330 1926 2336 1927
rect 2426 1931 2432 1932
rect 2426 1927 2427 1931
rect 2431 1927 2432 1931
rect 2426 1926 2432 1927
rect 2522 1931 2528 1932
rect 2522 1927 2523 1931
rect 2527 1927 2528 1931
rect 2618 1931 2619 1935
rect 2623 1931 2624 1935
rect 2618 1930 2624 1931
rect 2638 1935 2644 1936
rect 2638 1931 2639 1935
rect 2643 1931 2644 1935
rect 2638 1930 2644 1931
rect 2522 1926 2528 1927
rect 2046 1922 2052 1923
rect 2254 1924 2260 1925
rect 2006 1912 2012 1913
rect 1230 1911 1236 1912
rect 1230 1907 1231 1911
rect 1235 1907 1236 1911
rect 1230 1906 1236 1907
rect 1326 1911 1332 1912
rect 1326 1907 1327 1911
rect 1331 1907 1332 1911
rect 1326 1906 1332 1907
rect 1422 1911 1428 1912
rect 1422 1907 1423 1911
rect 1427 1907 1428 1911
rect 2006 1908 2007 1912
rect 2011 1908 2012 1912
rect 2006 1907 2012 1908
rect 1422 1906 1428 1907
rect 1306 1899 1312 1900
rect 1306 1895 1307 1899
rect 1311 1895 1312 1899
rect 1306 1894 1312 1895
rect 1402 1899 1408 1900
rect 1402 1895 1403 1899
rect 1407 1895 1408 1899
rect 1402 1894 1408 1895
rect 1498 1899 1504 1900
rect 1498 1895 1499 1899
rect 1503 1895 1504 1899
rect 1498 1894 1504 1895
rect 2006 1895 2012 1896
rect 1230 1892 1236 1893
rect 1230 1888 1231 1892
rect 1235 1888 1236 1892
rect 1230 1887 1236 1888
rect 1202 1871 1208 1872
rect 1202 1867 1203 1871
rect 1207 1867 1208 1871
rect 1202 1866 1208 1867
rect 1232 1863 1234 1887
rect 1308 1876 1310 1894
rect 1326 1892 1332 1893
rect 1326 1888 1327 1892
rect 1331 1888 1332 1892
rect 1326 1887 1332 1888
rect 1306 1875 1312 1876
rect 1306 1871 1307 1875
rect 1311 1871 1312 1875
rect 1306 1870 1312 1871
rect 1328 1863 1330 1887
rect 1404 1872 1406 1894
rect 1422 1892 1428 1893
rect 1422 1888 1423 1892
rect 1427 1888 1428 1892
rect 1422 1887 1428 1888
rect 1402 1871 1408 1872
rect 1334 1867 1340 1868
rect 1334 1863 1335 1867
rect 1339 1863 1340 1867
rect 1402 1867 1403 1871
rect 1407 1867 1408 1871
rect 1402 1866 1408 1867
rect 1424 1863 1426 1887
rect 583 1862 587 1863
rect 583 1857 587 1858
rect 655 1862 659 1863
rect 655 1857 659 1858
rect 719 1862 723 1863
rect 719 1857 723 1858
rect 751 1862 755 1863
rect 751 1857 755 1858
rect 847 1862 851 1863
rect 847 1857 851 1858
rect 855 1862 859 1863
rect 855 1857 859 1858
rect 943 1862 947 1863
rect 943 1857 947 1858
rect 991 1862 995 1863
rect 991 1857 995 1858
rect 1039 1862 1043 1863
rect 1039 1857 1043 1858
rect 1127 1862 1131 1863
rect 1127 1857 1131 1858
rect 1135 1862 1139 1863
rect 1135 1857 1139 1858
rect 1231 1862 1235 1863
rect 1231 1857 1235 1858
rect 1263 1862 1267 1863
rect 1263 1857 1267 1858
rect 1327 1862 1331 1863
rect 1334 1862 1340 1863
rect 1399 1862 1403 1863
rect 1327 1857 1331 1858
rect 584 1833 586 1857
rect 720 1833 722 1857
rect 794 1855 800 1856
rect 794 1851 795 1855
rect 799 1851 800 1855
rect 794 1850 800 1851
rect 582 1832 588 1833
rect 582 1828 583 1832
rect 587 1828 588 1832
rect 582 1827 588 1828
rect 718 1832 724 1833
rect 718 1828 719 1832
rect 723 1828 724 1832
rect 718 1827 724 1828
rect 796 1824 798 1850
rect 856 1833 858 1857
rect 992 1833 994 1857
rect 1066 1855 1072 1856
rect 1066 1851 1067 1855
rect 1071 1851 1072 1855
rect 1066 1850 1072 1851
rect 854 1832 860 1833
rect 854 1828 855 1832
rect 859 1828 860 1832
rect 854 1827 860 1828
rect 990 1832 996 1833
rect 990 1828 991 1832
rect 995 1828 996 1832
rect 990 1827 996 1828
rect 1068 1824 1070 1850
rect 1128 1833 1130 1857
rect 1202 1855 1208 1856
rect 1202 1851 1203 1855
rect 1207 1851 1208 1855
rect 1202 1850 1208 1851
rect 1170 1847 1176 1848
rect 1170 1843 1171 1847
rect 1175 1843 1176 1847
rect 1170 1842 1176 1843
rect 1126 1832 1132 1833
rect 1126 1828 1127 1832
rect 1131 1828 1132 1832
rect 1126 1827 1132 1828
rect 394 1823 400 1824
rect 394 1819 395 1823
rect 399 1819 400 1823
rect 394 1818 400 1819
rect 514 1823 520 1824
rect 514 1819 515 1823
rect 519 1819 520 1823
rect 514 1818 520 1819
rect 794 1823 800 1824
rect 794 1819 795 1823
rect 799 1819 800 1823
rect 794 1818 800 1819
rect 922 1823 928 1824
rect 922 1819 923 1823
rect 927 1819 928 1823
rect 922 1818 928 1819
rect 1066 1823 1072 1824
rect 1066 1819 1067 1823
rect 1071 1819 1072 1823
rect 1066 1818 1072 1819
rect 446 1813 452 1814
rect 446 1809 447 1813
rect 451 1809 452 1813
rect 446 1808 452 1809
rect 582 1813 588 1814
rect 582 1809 583 1813
rect 587 1809 588 1813
rect 582 1808 588 1809
rect 718 1813 724 1814
rect 718 1809 719 1813
rect 723 1809 724 1813
rect 718 1808 724 1809
rect 854 1813 860 1814
rect 854 1809 855 1813
rect 859 1809 860 1813
rect 854 1808 860 1809
rect 448 1783 450 1808
rect 584 1783 586 1808
rect 720 1783 722 1808
rect 856 1783 858 1808
rect 391 1782 395 1783
rect 391 1777 395 1778
rect 447 1782 451 1783
rect 447 1777 451 1778
rect 535 1782 539 1783
rect 535 1777 539 1778
rect 583 1782 587 1783
rect 583 1777 587 1778
rect 695 1782 699 1783
rect 695 1777 699 1778
rect 719 1782 723 1783
rect 719 1777 723 1778
rect 855 1782 859 1783
rect 855 1777 859 1778
rect 863 1782 867 1783
rect 863 1777 867 1778
rect 392 1756 394 1777
rect 536 1756 538 1777
rect 696 1756 698 1777
rect 864 1756 866 1777
rect 390 1755 396 1756
rect 390 1751 391 1755
rect 395 1751 396 1755
rect 390 1750 396 1751
rect 534 1755 540 1756
rect 534 1751 535 1755
rect 539 1751 540 1755
rect 534 1750 540 1751
rect 694 1755 700 1756
rect 694 1751 695 1755
rect 699 1751 700 1755
rect 694 1750 700 1751
rect 862 1755 868 1756
rect 862 1751 863 1755
rect 867 1751 868 1755
rect 862 1750 868 1751
rect 330 1747 336 1748
rect 330 1743 331 1747
rect 335 1743 336 1747
rect 330 1742 336 1743
rect 342 1747 348 1748
rect 342 1743 343 1747
rect 347 1743 348 1747
rect 662 1747 668 1748
rect 342 1742 348 1743
rect 618 1743 624 1744
rect 110 1739 116 1740
rect 110 1735 111 1739
rect 115 1735 116 1739
rect 110 1734 116 1735
rect 254 1736 260 1737
rect 112 1707 114 1734
rect 254 1732 255 1736
rect 259 1732 260 1736
rect 254 1731 260 1732
rect 256 1707 258 1731
rect 344 1716 346 1742
rect 618 1739 619 1743
rect 623 1739 624 1743
rect 662 1743 663 1747
rect 667 1743 668 1747
rect 662 1742 668 1743
rect 814 1747 820 1748
rect 814 1743 815 1747
rect 819 1743 820 1747
rect 814 1742 820 1743
rect 618 1738 624 1739
rect 390 1736 396 1737
rect 390 1732 391 1736
rect 395 1732 396 1736
rect 390 1731 396 1732
rect 534 1736 540 1737
rect 534 1732 535 1736
rect 539 1732 540 1736
rect 534 1731 540 1732
rect 342 1715 348 1716
rect 342 1711 343 1715
rect 347 1711 348 1715
rect 342 1710 348 1711
rect 392 1707 394 1731
rect 498 1711 504 1712
rect 498 1707 499 1711
rect 503 1707 504 1711
rect 536 1707 538 1731
rect 111 1706 115 1707
rect 111 1701 115 1702
rect 135 1706 139 1707
rect 135 1701 139 1702
rect 255 1706 259 1707
rect 255 1701 259 1702
rect 263 1706 267 1707
rect 263 1701 267 1702
rect 391 1706 395 1707
rect 391 1701 395 1702
rect 431 1706 435 1707
rect 498 1706 504 1707
rect 535 1706 539 1707
rect 431 1701 435 1702
rect 112 1674 114 1701
rect 136 1677 138 1701
rect 202 1699 208 1700
rect 202 1695 203 1699
rect 207 1695 208 1699
rect 202 1694 208 1695
rect 210 1699 216 1700
rect 210 1695 211 1699
rect 215 1695 216 1699
rect 210 1694 216 1695
rect 134 1676 140 1677
rect 110 1673 116 1674
rect 110 1669 111 1673
rect 115 1669 116 1673
rect 134 1672 135 1676
rect 139 1672 140 1676
rect 134 1671 140 1672
rect 110 1668 116 1669
rect 134 1657 140 1658
rect 110 1656 116 1657
rect 110 1652 111 1656
rect 115 1652 116 1656
rect 134 1653 135 1657
rect 139 1653 140 1657
rect 134 1652 140 1653
rect 110 1651 116 1652
rect 112 1631 114 1651
rect 136 1631 138 1652
rect 111 1630 115 1631
rect 111 1625 115 1626
rect 135 1630 139 1631
rect 135 1625 139 1626
rect 112 1605 114 1625
rect 110 1604 116 1605
rect 136 1604 138 1625
rect 110 1600 111 1604
rect 115 1600 116 1604
rect 110 1599 116 1600
rect 134 1603 140 1604
rect 134 1599 135 1603
rect 139 1599 140 1603
rect 204 1600 206 1694
rect 212 1668 214 1694
rect 264 1677 266 1701
rect 338 1699 344 1700
rect 338 1695 339 1699
rect 343 1695 344 1699
rect 338 1694 344 1695
rect 262 1676 268 1677
rect 262 1672 263 1676
rect 267 1672 268 1676
rect 262 1671 268 1672
rect 340 1668 342 1694
rect 432 1677 434 1701
rect 430 1676 436 1677
rect 430 1672 431 1676
rect 435 1672 436 1676
rect 430 1671 436 1672
rect 500 1668 502 1706
rect 535 1701 539 1702
rect 607 1706 611 1707
rect 607 1701 611 1702
rect 608 1677 610 1701
rect 620 1700 622 1738
rect 664 1716 666 1742
rect 694 1736 700 1737
rect 694 1732 695 1736
rect 699 1732 700 1736
rect 694 1731 700 1732
rect 662 1715 668 1716
rect 662 1711 663 1715
rect 667 1711 668 1715
rect 662 1710 668 1711
rect 696 1707 698 1731
rect 816 1716 818 1742
rect 862 1736 868 1737
rect 862 1732 863 1736
rect 867 1732 868 1736
rect 862 1731 868 1732
rect 814 1715 820 1716
rect 814 1711 815 1715
rect 819 1711 820 1715
rect 814 1710 820 1711
rect 864 1707 866 1731
rect 924 1716 926 1818
rect 990 1813 996 1814
rect 990 1809 991 1813
rect 995 1809 996 1813
rect 990 1808 996 1809
rect 1126 1813 1132 1814
rect 1126 1809 1127 1813
rect 1131 1809 1132 1813
rect 1126 1808 1132 1809
rect 992 1783 994 1808
rect 1128 1783 1130 1808
rect 991 1782 995 1783
rect 991 1777 995 1778
rect 1031 1782 1035 1783
rect 1031 1777 1035 1778
rect 1127 1782 1131 1783
rect 1127 1777 1131 1778
rect 1032 1756 1034 1777
rect 1030 1755 1036 1756
rect 1030 1751 1031 1755
rect 1035 1751 1036 1755
rect 1030 1750 1036 1751
rect 1172 1748 1174 1842
rect 1204 1824 1206 1850
rect 1264 1833 1266 1857
rect 1262 1832 1268 1833
rect 1262 1828 1263 1832
rect 1267 1828 1268 1832
rect 1262 1827 1268 1828
rect 1336 1824 1338 1862
rect 1399 1857 1403 1858
rect 1423 1862 1427 1863
rect 1423 1857 1427 1858
rect 1400 1833 1402 1857
rect 1500 1856 1502 1894
rect 2006 1891 2007 1895
rect 2011 1891 2012 1895
rect 2006 1890 2012 1891
rect 2008 1863 2010 1890
rect 2048 1883 2050 1922
rect 2254 1920 2255 1924
rect 2259 1920 2260 1924
rect 2254 1919 2260 1920
rect 2256 1883 2258 1919
rect 2332 1904 2334 1926
rect 2350 1924 2356 1925
rect 2350 1920 2351 1924
rect 2355 1920 2356 1924
rect 2350 1919 2356 1920
rect 2330 1903 2336 1904
rect 2330 1899 2331 1903
rect 2335 1899 2336 1903
rect 2330 1898 2336 1899
rect 2352 1883 2354 1919
rect 2428 1904 2430 1926
rect 2446 1924 2452 1925
rect 2446 1920 2447 1924
rect 2451 1920 2452 1924
rect 2446 1919 2452 1920
rect 2426 1903 2432 1904
rect 2426 1899 2427 1903
rect 2431 1899 2432 1903
rect 2426 1898 2432 1899
rect 2448 1883 2450 1919
rect 2524 1904 2526 1926
rect 2542 1924 2548 1925
rect 2542 1920 2543 1924
rect 2547 1920 2548 1924
rect 2542 1919 2548 1920
rect 2522 1903 2528 1904
rect 2522 1899 2523 1903
rect 2527 1899 2528 1903
rect 2522 1898 2528 1899
rect 2466 1895 2472 1896
rect 2466 1891 2467 1895
rect 2471 1891 2472 1895
rect 2466 1890 2472 1891
rect 2047 1882 2051 1883
rect 2047 1877 2051 1878
rect 2183 1882 2187 1883
rect 2183 1877 2187 1878
rect 2255 1882 2259 1883
rect 2255 1877 2259 1878
rect 2279 1882 2283 1883
rect 2279 1877 2283 1878
rect 2351 1882 2355 1883
rect 2351 1877 2355 1878
rect 2383 1882 2387 1883
rect 2383 1877 2387 1878
rect 2447 1882 2451 1883
rect 2447 1877 2451 1878
rect 1535 1862 1539 1863
rect 1535 1857 1539 1858
rect 2007 1862 2011 1863
rect 2007 1857 2011 1858
rect 1482 1855 1488 1856
rect 1482 1851 1483 1855
rect 1487 1851 1488 1855
rect 1482 1850 1488 1851
rect 1498 1855 1504 1856
rect 1498 1851 1499 1855
rect 1503 1851 1504 1855
rect 1498 1850 1504 1851
rect 1398 1832 1404 1833
rect 1398 1828 1399 1832
rect 1403 1828 1404 1832
rect 1398 1827 1404 1828
rect 1484 1824 1486 1850
rect 1536 1833 1538 1857
rect 1534 1832 1540 1833
rect 1534 1828 1535 1832
rect 1539 1828 1540 1832
rect 2008 1830 2010 1857
rect 2048 1850 2050 1877
rect 2184 1853 2186 1877
rect 2202 1875 2208 1876
rect 2202 1871 2203 1875
rect 2207 1871 2208 1875
rect 2202 1870 2208 1871
rect 2182 1852 2188 1853
rect 2046 1849 2052 1850
rect 2046 1845 2047 1849
rect 2051 1845 2052 1849
rect 2182 1848 2183 1852
rect 2187 1848 2188 1852
rect 2182 1847 2188 1848
rect 2046 1844 2052 1845
rect 2182 1833 2188 1834
rect 2046 1832 2052 1833
rect 1534 1827 1540 1828
rect 2006 1829 2012 1830
rect 2006 1825 2007 1829
rect 2011 1825 2012 1829
rect 2046 1828 2047 1832
rect 2051 1828 2052 1832
rect 2182 1829 2183 1833
rect 2187 1829 2188 1833
rect 2182 1828 2188 1829
rect 2046 1827 2052 1828
rect 2006 1824 2012 1825
rect 1202 1823 1208 1824
rect 1202 1819 1203 1823
rect 1207 1819 1208 1823
rect 1202 1818 1208 1819
rect 1334 1823 1340 1824
rect 1334 1819 1335 1823
rect 1339 1819 1340 1823
rect 1334 1818 1340 1819
rect 1466 1823 1472 1824
rect 1466 1819 1467 1823
rect 1471 1819 1472 1823
rect 1466 1818 1472 1819
rect 1482 1823 1488 1824
rect 1482 1819 1483 1823
rect 1487 1819 1488 1823
rect 1482 1818 1488 1819
rect 1262 1813 1268 1814
rect 1262 1809 1263 1813
rect 1267 1809 1268 1813
rect 1262 1808 1268 1809
rect 1398 1813 1404 1814
rect 1398 1809 1399 1813
rect 1403 1809 1404 1813
rect 1398 1808 1404 1809
rect 1264 1783 1266 1808
rect 1400 1783 1402 1808
rect 1207 1782 1211 1783
rect 1207 1777 1211 1778
rect 1263 1782 1267 1783
rect 1263 1777 1267 1778
rect 1383 1782 1387 1783
rect 1383 1777 1387 1778
rect 1399 1782 1403 1783
rect 1399 1777 1403 1778
rect 1208 1756 1210 1777
rect 1384 1756 1386 1777
rect 1206 1755 1212 1756
rect 1206 1751 1207 1755
rect 1211 1751 1212 1755
rect 1206 1750 1212 1751
rect 1382 1755 1388 1756
rect 1382 1751 1383 1755
rect 1387 1751 1388 1755
rect 1382 1750 1388 1751
rect 1170 1747 1176 1748
rect 1106 1743 1112 1744
rect 1106 1739 1107 1743
rect 1111 1739 1112 1743
rect 1170 1743 1171 1747
rect 1175 1743 1176 1747
rect 1170 1742 1176 1743
rect 1106 1738 1112 1739
rect 1030 1736 1036 1737
rect 1030 1732 1031 1736
rect 1035 1732 1036 1736
rect 1030 1731 1036 1732
rect 918 1715 926 1716
rect 918 1711 919 1715
rect 923 1713 926 1715
rect 923 1711 924 1713
rect 918 1710 924 1711
rect 1032 1707 1034 1731
rect 1108 1716 1110 1738
rect 1206 1736 1212 1737
rect 1206 1732 1207 1736
rect 1211 1732 1212 1736
rect 1206 1731 1212 1732
rect 1382 1736 1388 1737
rect 1382 1732 1383 1736
rect 1387 1732 1388 1736
rect 1382 1731 1388 1732
rect 1106 1715 1112 1716
rect 1074 1711 1080 1712
rect 1074 1707 1075 1711
rect 1079 1707 1080 1711
rect 1106 1711 1107 1715
rect 1111 1711 1112 1715
rect 1106 1710 1112 1711
rect 1208 1707 1210 1731
rect 1384 1707 1386 1731
rect 1468 1716 1470 1818
rect 1534 1813 1540 1814
rect 1534 1809 1535 1813
rect 1539 1809 1540 1813
rect 1534 1808 1540 1809
rect 2006 1812 2012 1813
rect 2006 1808 2007 1812
rect 2011 1808 2012 1812
rect 1536 1783 1538 1808
rect 2006 1807 2012 1808
rect 2008 1783 2010 1807
rect 2048 1803 2050 1827
rect 2184 1803 2186 1828
rect 2047 1802 2051 1803
rect 2047 1797 2051 1798
rect 2127 1802 2131 1803
rect 2127 1797 2131 1798
rect 2183 1802 2187 1803
rect 2183 1797 2187 1798
rect 1535 1782 1539 1783
rect 1535 1777 1539 1778
rect 1559 1782 1563 1783
rect 1559 1777 1563 1778
rect 1743 1782 1747 1783
rect 1743 1777 1747 1778
rect 2007 1782 2011 1783
rect 2007 1777 2011 1778
rect 2048 1777 2050 1797
rect 1560 1756 1562 1777
rect 1744 1756 1746 1777
rect 2008 1757 2010 1777
rect 2046 1776 2052 1777
rect 2128 1776 2130 1797
rect 2046 1772 2047 1776
rect 2051 1772 2052 1776
rect 2046 1771 2052 1772
rect 2126 1775 2132 1776
rect 2126 1771 2127 1775
rect 2131 1771 2132 1775
rect 2126 1770 2132 1771
rect 2204 1768 2206 1870
rect 2280 1853 2282 1877
rect 2384 1853 2386 1877
rect 2458 1875 2464 1876
rect 2458 1871 2459 1875
rect 2463 1871 2464 1875
rect 2458 1870 2464 1871
rect 2278 1852 2284 1853
rect 2278 1848 2279 1852
rect 2283 1848 2284 1852
rect 2278 1847 2284 1848
rect 2382 1852 2388 1853
rect 2382 1848 2383 1852
rect 2387 1848 2388 1852
rect 2382 1847 2388 1848
rect 2460 1844 2462 1870
rect 2468 1844 2470 1890
rect 2544 1883 2546 1919
rect 2487 1882 2491 1883
rect 2487 1877 2491 1878
rect 2543 1882 2547 1883
rect 2543 1877 2547 1878
rect 2591 1882 2595 1883
rect 2591 1877 2595 1878
rect 2488 1853 2490 1877
rect 2592 1853 2594 1877
rect 2640 1876 2642 1930
rect 2646 1924 2652 1925
rect 2646 1920 2647 1924
rect 2651 1920 2652 1924
rect 2646 1919 2652 1920
rect 2648 1883 2650 1919
rect 2716 1904 2718 2006
rect 2774 2001 2780 2002
rect 2774 1997 2775 2001
rect 2779 1997 2780 2001
rect 2774 1996 2780 1997
rect 2776 1971 2778 1996
rect 2767 1970 2771 1971
rect 2767 1965 2771 1966
rect 2775 1970 2779 1971
rect 2775 1965 2779 1966
rect 2768 1944 2770 1965
rect 2766 1943 2772 1944
rect 2766 1939 2767 1943
rect 2771 1939 2772 1943
rect 2766 1938 2772 1939
rect 2844 1936 2846 2038
rect 2852 2012 2854 2038
rect 2920 2021 2922 2045
rect 2994 2043 3000 2044
rect 2994 2039 2995 2043
rect 2999 2039 3000 2043
rect 2994 2038 3000 2039
rect 2918 2020 2924 2021
rect 2918 2016 2919 2020
rect 2923 2016 2924 2020
rect 2918 2015 2924 2016
rect 2996 2012 2998 2038
rect 3080 2021 3082 2045
rect 3154 2043 3160 2044
rect 3154 2039 3155 2043
rect 3159 2039 3160 2043
rect 3154 2038 3160 2039
rect 3078 2020 3084 2021
rect 3078 2016 3079 2020
rect 3083 2016 3084 2020
rect 3078 2015 3084 2016
rect 3156 2012 3158 2038
rect 3264 2021 3266 2045
rect 3338 2043 3344 2044
rect 3338 2039 3339 2043
rect 3343 2039 3344 2043
rect 3338 2038 3344 2039
rect 3262 2020 3268 2021
rect 3262 2016 3263 2020
rect 3267 2016 3268 2020
rect 3262 2015 3268 2016
rect 3340 2012 3342 2038
rect 3380 2012 3382 2054
rect 3520 2051 3522 2083
rect 3688 2051 3690 2083
rect 3764 2068 3766 2090
rect 3762 2067 3768 2068
rect 3730 2063 3736 2064
rect 3730 2059 3731 2063
rect 3735 2059 3736 2063
rect 3762 2063 3763 2067
rect 3767 2063 3768 2067
rect 3762 2062 3768 2063
rect 3730 2058 3736 2059
rect 3455 2050 3459 2051
rect 3455 2045 3459 2046
rect 3519 2050 3523 2051
rect 3519 2045 3523 2046
rect 3655 2050 3659 2051
rect 3655 2045 3659 2046
rect 3687 2050 3691 2051
rect 3687 2045 3691 2046
rect 3456 2021 3458 2045
rect 3656 2021 3658 2045
rect 3454 2020 3460 2021
rect 3454 2016 3455 2020
rect 3459 2016 3460 2020
rect 3454 2015 3460 2016
rect 3654 2020 3660 2021
rect 3654 2016 3655 2020
rect 3659 2016 3660 2020
rect 3654 2015 3660 2016
rect 3732 2012 3734 2058
rect 3738 2043 3744 2044
rect 3738 2039 3739 2043
rect 3743 2039 3744 2043
rect 3738 2038 3744 2039
rect 3740 2012 3742 2038
rect 2850 2011 2856 2012
rect 2850 2007 2851 2011
rect 2855 2007 2856 2011
rect 2850 2006 2856 2007
rect 2994 2011 3000 2012
rect 2994 2007 2995 2011
rect 2999 2007 3000 2011
rect 2994 2006 3000 2007
rect 3154 2011 3160 2012
rect 3154 2007 3155 2011
rect 3159 2007 3160 2011
rect 3154 2006 3160 2007
rect 3338 2011 3344 2012
rect 3338 2007 3339 2011
rect 3343 2007 3344 2011
rect 3338 2006 3344 2007
rect 3378 2011 3384 2012
rect 3378 2007 3379 2011
rect 3383 2007 3384 2011
rect 3378 2006 3384 2007
rect 3730 2011 3736 2012
rect 3730 2007 3731 2011
rect 3735 2007 3736 2011
rect 3730 2006 3736 2007
rect 3738 2011 3744 2012
rect 3738 2007 3739 2011
rect 3743 2007 3744 2011
rect 3738 2006 3744 2007
rect 2918 2001 2924 2002
rect 2918 1997 2919 2001
rect 2923 1997 2924 2001
rect 2918 1996 2924 1997
rect 3078 2001 3084 2002
rect 3078 1997 3079 2001
rect 3083 1997 3084 2001
rect 3078 1996 3084 1997
rect 3262 2001 3268 2002
rect 3262 1997 3263 2001
rect 3267 1997 3268 2001
rect 3262 1996 3268 1997
rect 3454 2001 3460 2002
rect 3454 1997 3455 2001
rect 3459 1997 3460 2001
rect 3454 1996 3460 1997
rect 3654 2001 3660 2002
rect 3654 1997 3655 2001
rect 3659 1997 3660 2001
rect 3654 1996 3660 1997
rect 2920 1971 2922 1996
rect 3080 1971 3082 1996
rect 3264 1971 3266 1996
rect 3456 1971 3458 1996
rect 3656 1971 3658 1996
rect 2919 1970 2923 1971
rect 2919 1965 2923 1966
rect 3079 1970 3083 1971
rect 3079 1965 3083 1966
rect 3103 1970 3107 1971
rect 3103 1965 3107 1966
rect 3263 1970 3267 1971
rect 3263 1965 3267 1966
rect 3319 1970 3323 1971
rect 3319 1965 3323 1966
rect 3455 1970 3459 1971
rect 3455 1965 3459 1966
rect 3543 1970 3547 1971
rect 3543 1965 3547 1966
rect 3655 1970 3659 1971
rect 3655 1965 3659 1966
rect 3775 1970 3779 1971
rect 3775 1965 3779 1966
rect 2920 1944 2922 1965
rect 3104 1944 3106 1965
rect 3320 1944 3322 1965
rect 3544 1944 3546 1965
rect 3776 1944 3778 1965
rect 2918 1943 2924 1944
rect 2918 1939 2919 1943
rect 2923 1939 2924 1943
rect 2918 1938 2924 1939
rect 3102 1943 3108 1944
rect 3102 1939 3103 1943
rect 3107 1939 3108 1943
rect 3102 1938 3108 1939
rect 3318 1943 3324 1944
rect 3318 1939 3319 1943
rect 3323 1939 3324 1943
rect 3318 1938 3324 1939
rect 3542 1943 3548 1944
rect 3542 1939 3543 1943
rect 3547 1939 3548 1943
rect 3542 1938 3548 1939
rect 3774 1943 3780 1944
rect 3774 1939 3775 1943
rect 3779 1939 3780 1943
rect 3774 1938 3780 1939
rect 2842 1935 2848 1936
rect 2842 1931 2843 1935
rect 2847 1931 2848 1935
rect 2842 1930 2848 1931
rect 2858 1935 2864 1936
rect 2858 1931 2859 1935
rect 2863 1931 2864 1935
rect 2858 1930 2864 1931
rect 3006 1935 3012 1936
rect 3006 1931 3007 1935
rect 3011 1931 3012 1935
rect 3006 1930 3012 1931
rect 3186 1935 3192 1936
rect 3186 1931 3187 1935
rect 3191 1931 3192 1935
rect 3186 1930 3192 1931
rect 3402 1935 3408 1936
rect 3402 1931 3403 1935
rect 3407 1931 3408 1935
rect 3402 1930 3408 1931
rect 3750 1935 3756 1936
rect 3750 1931 3751 1935
rect 3755 1931 3756 1935
rect 3750 1930 3756 1931
rect 2766 1924 2772 1925
rect 2766 1920 2767 1924
rect 2771 1920 2772 1924
rect 2766 1919 2772 1920
rect 2714 1903 2720 1904
rect 2714 1899 2715 1903
rect 2719 1899 2720 1903
rect 2714 1898 2720 1899
rect 2768 1883 2770 1919
rect 2860 1904 2862 1930
rect 2918 1924 2924 1925
rect 2918 1920 2919 1924
rect 2923 1920 2924 1924
rect 2918 1919 2924 1920
rect 2858 1903 2864 1904
rect 2858 1899 2859 1903
rect 2863 1899 2864 1903
rect 2858 1898 2864 1899
rect 2920 1883 2922 1919
rect 3008 1904 3010 1930
rect 3102 1924 3108 1925
rect 3102 1920 3103 1924
rect 3107 1920 3108 1924
rect 3102 1919 3108 1920
rect 3006 1903 3012 1904
rect 3006 1899 3007 1903
rect 3011 1899 3012 1903
rect 3006 1898 3012 1899
rect 3104 1883 3106 1919
rect 3188 1904 3190 1930
rect 3318 1924 3324 1925
rect 3318 1920 3319 1924
rect 3323 1920 3324 1924
rect 3318 1919 3324 1920
rect 3186 1903 3192 1904
rect 3186 1899 3187 1903
rect 3191 1899 3192 1903
rect 3186 1898 3192 1899
rect 3320 1883 3322 1919
rect 3404 1904 3406 1930
rect 3542 1924 3548 1925
rect 3542 1920 3543 1924
rect 3547 1920 3548 1924
rect 3542 1919 3548 1920
rect 3402 1903 3408 1904
rect 3402 1899 3403 1903
rect 3407 1899 3408 1903
rect 3402 1898 3408 1899
rect 3544 1883 3546 1919
rect 2647 1882 2651 1883
rect 2647 1877 2651 1878
rect 2703 1882 2707 1883
rect 2703 1877 2707 1878
rect 2767 1882 2771 1883
rect 2767 1877 2771 1878
rect 2831 1882 2835 1883
rect 2831 1877 2835 1878
rect 2919 1882 2923 1883
rect 2919 1877 2923 1878
rect 2991 1882 2995 1883
rect 2991 1877 2995 1878
rect 3103 1882 3107 1883
rect 3103 1877 3107 1878
rect 3183 1882 3187 1883
rect 3183 1877 3187 1878
rect 3319 1882 3323 1883
rect 3319 1877 3323 1878
rect 3399 1882 3403 1883
rect 3399 1877 3403 1878
rect 3543 1882 3547 1883
rect 3543 1877 3547 1878
rect 3631 1882 3635 1883
rect 3631 1877 3635 1878
rect 2638 1875 2644 1876
rect 2638 1871 2639 1875
rect 2643 1871 2644 1875
rect 2638 1870 2644 1871
rect 2666 1875 2672 1876
rect 2666 1871 2667 1875
rect 2671 1871 2672 1875
rect 2666 1870 2672 1871
rect 2486 1852 2492 1853
rect 2486 1848 2487 1852
rect 2491 1848 2492 1852
rect 2486 1847 2492 1848
rect 2590 1852 2596 1853
rect 2590 1848 2591 1852
rect 2595 1848 2596 1852
rect 2590 1847 2596 1848
rect 2668 1844 2670 1870
rect 2704 1853 2706 1877
rect 2832 1853 2834 1877
rect 2870 1875 2876 1876
rect 2870 1871 2871 1875
rect 2875 1871 2876 1875
rect 2870 1870 2876 1871
rect 2906 1875 2912 1876
rect 2906 1871 2907 1875
rect 2911 1871 2912 1875
rect 2906 1870 2912 1871
rect 2702 1852 2708 1853
rect 2702 1848 2703 1852
rect 2707 1848 2708 1852
rect 2702 1847 2708 1848
rect 2830 1852 2836 1853
rect 2830 1848 2831 1852
rect 2835 1848 2836 1852
rect 2830 1847 2836 1848
rect 2458 1843 2464 1844
rect 2458 1839 2459 1843
rect 2463 1839 2464 1843
rect 2458 1838 2464 1839
rect 2466 1843 2472 1844
rect 2466 1839 2467 1843
rect 2471 1839 2472 1843
rect 2466 1838 2472 1839
rect 2666 1843 2672 1844
rect 2666 1839 2667 1843
rect 2671 1839 2672 1843
rect 2666 1838 2672 1839
rect 2770 1843 2776 1844
rect 2770 1839 2771 1843
rect 2775 1839 2776 1843
rect 2770 1838 2776 1839
rect 2278 1833 2284 1834
rect 2278 1829 2279 1833
rect 2283 1829 2284 1833
rect 2278 1828 2284 1829
rect 2382 1833 2388 1834
rect 2382 1829 2383 1833
rect 2387 1829 2388 1833
rect 2382 1828 2388 1829
rect 2486 1833 2492 1834
rect 2486 1829 2487 1833
rect 2491 1829 2492 1833
rect 2486 1828 2492 1829
rect 2590 1833 2596 1834
rect 2590 1829 2591 1833
rect 2595 1829 2596 1833
rect 2590 1828 2596 1829
rect 2702 1833 2708 1834
rect 2702 1829 2703 1833
rect 2707 1829 2708 1833
rect 2702 1828 2708 1829
rect 2280 1803 2282 1828
rect 2384 1803 2386 1828
rect 2488 1803 2490 1828
rect 2592 1803 2594 1828
rect 2704 1803 2706 1828
rect 2279 1802 2283 1803
rect 2279 1797 2283 1798
rect 2311 1802 2315 1803
rect 2311 1797 2315 1798
rect 2383 1802 2387 1803
rect 2383 1797 2387 1798
rect 2487 1802 2491 1803
rect 2487 1797 2491 1798
rect 2495 1802 2499 1803
rect 2495 1797 2499 1798
rect 2591 1802 2595 1803
rect 2591 1797 2595 1798
rect 2687 1802 2691 1803
rect 2687 1797 2691 1798
rect 2703 1802 2707 1803
rect 2703 1797 2707 1798
rect 2312 1776 2314 1797
rect 2496 1776 2498 1797
rect 2688 1776 2690 1797
rect 2310 1775 2316 1776
rect 2310 1771 2311 1775
rect 2315 1771 2316 1775
rect 2310 1770 2316 1771
rect 2494 1775 2500 1776
rect 2494 1771 2495 1775
rect 2499 1771 2500 1775
rect 2494 1770 2500 1771
rect 2686 1775 2692 1776
rect 2686 1771 2687 1775
rect 2691 1771 2692 1775
rect 2686 1770 2692 1771
rect 2202 1767 2208 1768
rect 2202 1763 2203 1767
rect 2207 1763 2208 1767
rect 2202 1762 2208 1763
rect 2046 1759 2052 1760
rect 2006 1756 2012 1757
rect 1558 1755 1564 1756
rect 1558 1751 1559 1755
rect 1563 1751 1564 1755
rect 1558 1750 1564 1751
rect 1742 1755 1748 1756
rect 1742 1751 1743 1755
rect 1747 1751 1748 1755
rect 2006 1752 2007 1756
rect 2011 1752 2012 1756
rect 2046 1755 2047 1759
rect 2051 1755 2052 1759
rect 2046 1754 2052 1755
rect 2126 1756 2132 1757
rect 2006 1751 2012 1752
rect 1742 1750 1748 1751
rect 1518 1743 1524 1744
rect 1518 1739 1519 1743
rect 1523 1739 1524 1743
rect 1518 1738 1524 1739
rect 1634 1743 1640 1744
rect 1634 1739 1635 1743
rect 1639 1739 1640 1743
rect 1634 1738 1640 1739
rect 1818 1743 1824 1744
rect 1818 1739 1819 1743
rect 1823 1739 1824 1743
rect 1818 1738 1824 1739
rect 2006 1739 2012 1740
rect 1520 1716 1522 1738
rect 1558 1736 1564 1737
rect 1558 1732 1559 1736
rect 1563 1732 1564 1736
rect 1558 1731 1564 1732
rect 1466 1715 1472 1716
rect 1466 1711 1467 1715
rect 1471 1711 1472 1715
rect 1466 1710 1472 1711
rect 1518 1715 1524 1716
rect 1518 1711 1519 1715
rect 1523 1711 1524 1715
rect 1518 1710 1524 1711
rect 1560 1707 1562 1731
rect 1636 1716 1638 1738
rect 1742 1736 1748 1737
rect 1742 1732 1743 1736
rect 1747 1732 1748 1736
rect 1742 1731 1748 1732
rect 1634 1715 1640 1716
rect 1634 1711 1635 1715
rect 1639 1711 1640 1715
rect 1634 1710 1640 1711
rect 1744 1707 1746 1731
rect 695 1706 699 1707
rect 695 1701 699 1702
rect 799 1706 803 1707
rect 799 1701 803 1702
rect 863 1706 867 1707
rect 863 1701 867 1702
rect 999 1706 1003 1707
rect 999 1701 1003 1702
rect 1031 1706 1035 1707
rect 1074 1706 1080 1707
rect 1199 1706 1203 1707
rect 1031 1701 1035 1702
rect 618 1699 624 1700
rect 618 1695 619 1699
rect 623 1695 624 1699
rect 618 1694 624 1695
rect 682 1699 688 1700
rect 682 1695 683 1699
rect 687 1695 688 1699
rect 682 1694 688 1695
rect 606 1676 612 1677
rect 606 1672 607 1676
rect 611 1672 612 1676
rect 606 1671 612 1672
rect 684 1668 686 1694
rect 800 1677 802 1701
rect 1000 1677 1002 1701
rect 798 1676 804 1677
rect 798 1672 799 1676
rect 803 1672 804 1676
rect 798 1671 804 1672
rect 998 1676 1004 1677
rect 998 1672 999 1676
rect 1003 1672 1004 1676
rect 998 1671 1004 1672
rect 1076 1668 1078 1706
rect 1199 1701 1203 1702
rect 1207 1706 1211 1707
rect 1207 1701 1211 1702
rect 1383 1706 1387 1707
rect 1383 1701 1387 1702
rect 1407 1706 1411 1707
rect 1407 1701 1411 1702
rect 1559 1706 1563 1707
rect 1559 1701 1563 1702
rect 1623 1706 1627 1707
rect 1623 1701 1627 1702
rect 1743 1706 1747 1707
rect 1743 1701 1747 1702
rect 1200 1677 1202 1701
rect 1254 1699 1260 1700
rect 1254 1695 1255 1699
rect 1259 1698 1260 1699
rect 1274 1699 1280 1700
rect 1259 1695 1262 1698
rect 1254 1694 1262 1695
rect 1274 1695 1275 1699
rect 1279 1695 1280 1699
rect 1274 1694 1280 1695
rect 1198 1676 1204 1677
rect 1198 1672 1199 1676
rect 1203 1672 1204 1676
rect 1198 1671 1204 1672
rect 210 1667 216 1668
rect 210 1663 211 1667
rect 215 1663 216 1667
rect 210 1662 216 1663
rect 338 1667 344 1668
rect 338 1663 339 1667
rect 343 1663 344 1667
rect 338 1662 344 1663
rect 498 1667 504 1668
rect 498 1663 499 1667
rect 503 1663 504 1667
rect 498 1662 504 1663
rect 682 1667 688 1668
rect 682 1663 683 1667
rect 687 1663 688 1667
rect 682 1662 688 1663
rect 874 1667 880 1668
rect 874 1663 875 1667
rect 879 1663 880 1667
rect 874 1662 880 1663
rect 1074 1667 1080 1668
rect 1074 1663 1075 1667
rect 1079 1663 1080 1667
rect 1074 1662 1080 1663
rect 262 1657 268 1658
rect 262 1653 263 1657
rect 267 1653 268 1657
rect 262 1652 268 1653
rect 430 1657 436 1658
rect 430 1653 431 1657
rect 435 1653 436 1657
rect 430 1652 436 1653
rect 606 1657 612 1658
rect 606 1653 607 1657
rect 611 1653 612 1657
rect 606 1652 612 1653
rect 798 1657 804 1658
rect 798 1653 799 1657
rect 803 1653 804 1657
rect 798 1652 804 1653
rect 264 1631 266 1652
rect 432 1631 434 1652
rect 608 1631 610 1652
rect 800 1631 802 1652
rect 263 1630 267 1631
rect 263 1625 267 1626
rect 287 1630 291 1631
rect 287 1625 291 1626
rect 431 1630 435 1631
rect 431 1625 435 1626
rect 471 1630 475 1631
rect 471 1625 475 1626
rect 607 1630 611 1631
rect 607 1625 611 1626
rect 655 1630 659 1631
rect 655 1625 659 1626
rect 799 1630 803 1631
rect 799 1625 803 1626
rect 839 1630 843 1631
rect 839 1625 843 1626
rect 288 1604 290 1625
rect 472 1604 474 1625
rect 656 1604 658 1625
rect 840 1604 842 1625
rect 286 1603 292 1604
rect 134 1598 140 1599
rect 202 1599 208 1600
rect 202 1595 203 1599
rect 207 1595 208 1599
rect 286 1599 287 1603
rect 291 1599 292 1603
rect 286 1598 292 1599
rect 470 1603 476 1604
rect 470 1599 471 1603
rect 475 1599 476 1603
rect 470 1598 476 1599
rect 654 1603 660 1604
rect 654 1599 655 1603
rect 659 1599 660 1603
rect 654 1598 660 1599
rect 838 1603 844 1604
rect 838 1599 839 1603
rect 843 1599 844 1603
rect 838 1598 844 1599
rect 202 1594 208 1595
rect 222 1595 228 1596
rect 222 1591 223 1595
rect 227 1591 228 1595
rect 738 1595 744 1596
rect 222 1590 228 1591
rect 546 1591 552 1592
rect 110 1587 116 1588
rect 110 1583 111 1587
rect 115 1583 116 1587
rect 110 1582 116 1583
rect 134 1584 140 1585
rect 112 1551 114 1582
rect 134 1580 135 1584
rect 139 1580 140 1584
rect 134 1579 140 1580
rect 136 1551 138 1579
rect 224 1564 226 1590
rect 546 1587 547 1591
rect 551 1587 552 1591
rect 546 1586 552 1587
rect 730 1591 736 1592
rect 730 1587 731 1591
rect 735 1587 736 1591
rect 738 1591 739 1595
rect 743 1591 744 1595
rect 738 1590 744 1591
rect 730 1586 736 1587
rect 286 1584 292 1585
rect 286 1580 287 1584
rect 291 1580 292 1584
rect 286 1579 292 1580
rect 470 1584 476 1585
rect 470 1580 471 1584
rect 475 1580 476 1584
rect 470 1579 476 1580
rect 222 1563 228 1564
rect 222 1559 223 1563
rect 227 1559 228 1563
rect 222 1558 228 1559
rect 288 1551 290 1579
rect 390 1559 396 1560
rect 390 1555 391 1559
rect 395 1555 396 1559
rect 390 1554 396 1555
rect 111 1550 115 1551
rect 111 1545 115 1546
rect 135 1550 139 1551
rect 135 1545 139 1546
rect 287 1550 291 1551
rect 287 1545 291 1546
rect 295 1550 299 1551
rect 295 1545 299 1546
rect 112 1518 114 1545
rect 136 1521 138 1545
rect 250 1543 256 1544
rect 250 1539 251 1543
rect 255 1539 256 1543
rect 250 1538 256 1539
rect 258 1543 264 1544
rect 258 1539 259 1543
rect 263 1539 264 1543
rect 258 1538 264 1539
rect 134 1520 140 1521
rect 110 1517 116 1518
rect 110 1513 111 1517
rect 115 1513 116 1517
rect 134 1516 135 1520
rect 139 1516 140 1520
rect 134 1515 140 1516
rect 110 1512 116 1513
rect 134 1501 140 1502
rect 110 1500 116 1501
rect 110 1496 111 1500
rect 115 1496 116 1500
rect 134 1497 135 1501
rect 139 1497 140 1501
rect 134 1496 140 1497
rect 110 1495 116 1496
rect 112 1475 114 1495
rect 136 1475 138 1496
rect 111 1474 115 1475
rect 111 1469 115 1470
rect 135 1474 139 1475
rect 135 1469 139 1470
rect 175 1474 179 1475
rect 175 1469 179 1470
rect 112 1449 114 1469
rect 110 1448 116 1449
rect 176 1448 178 1469
rect 110 1444 111 1448
rect 115 1444 116 1448
rect 110 1443 116 1444
rect 174 1447 180 1448
rect 174 1443 175 1447
rect 179 1443 180 1447
rect 174 1442 180 1443
rect 252 1440 254 1538
rect 260 1512 262 1538
rect 296 1521 298 1545
rect 370 1543 376 1544
rect 370 1539 371 1543
rect 375 1539 376 1543
rect 370 1538 376 1539
rect 294 1520 300 1521
rect 294 1516 295 1520
rect 299 1516 300 1520
rect 294 1515 300 1516
rect 372 1512 374 1538
rect 392 1512 394 1554
rect 472 1551 474 1579
rect 548 1564 550 1586
rect 654 1584 660 1585
rect 654 1580 655 1584
rect 659 1580 660 1584
rect 654 1579 660 1580
rect 546 1563 552 1564
rect 546 1559 547 1563
rect 551 1559 552 1563
rect 546 1558 552 1559
rect 656 1551 658 1579
rect 471 1550 475 1551
rect 471 1545 475 1546
rect 487 1550 491 1551
rect 487 1545 491 1546
rect 655 1550 659 1551
rect 655 1545 659 1546
rect 687 1550 691 1551
rect 687 1545 691 1546
rect 488 1521 490 1545
rect 688 1521 690 1545
rect 732 1544 734 1586
rect 740 1572 742 1590
rect 838 1584 844 1585
rect 838 1580 839 1584
rect 843 1580 844 1584
rect 838 1579 844 1580
rect 738 1571 744 1572
rect 738 1567 739 1571
rect 743 1567 744 1571
rect 738 1566 744 1567
rect 840 1551 842 1579
rect 876 1564 878 1662
rect 998 1657 1004 1658
rect 998 1653 999 1657
rect 1003 1653 1004 1657
rect 998 1652 1004 1653
rect 1198 1657 1204 1658
rect 1198 1653 1199 1657
rect 1203 1653 1204 1657
rect 1198 1652 1204 1653
rect 1000 1631 1002 1652
rect 1200 1631 1202 1652
rect 999 1630 1003 1631
rect 999 1625 1003 1626
rect 1015 1630 1019 1631
rect 1015 1625 1019 1626
rect 1183 1630 1187 1631
rect 1183 1625 1187 1626
rect 1199 1630 1203 1631
rect 1199 1625 1203 1626
rect 1016 1604 1018 1625
rect 1184 1604 1186 1625
rect 1014 1603 1020 1604
rect 1014 1599 1015 1603
rect 1019 1599 1020 1603
rect 1014 1598 1020 1599
rect 1182 1603 1188 1604
rect 1182 1599 1183 1603
rect 1187 1599 1188 1603
rect 1182 1598 1188 1599
rect 1260 1596 1262 1694
rect 1276 1668 1278 1694
rect 1302 1687 1308 1688
rect 1302 1683 1303 1687
rect 1307 1683 1308 1687
rect 1302 1682 1308 1683
rect 1304 1668 1306 1682
rect 1408 1677 1410 1701
rect 1624 1677 1626 1701
rect 1820 1700 1822 1738
rect 2006 1735 2007 1739
rect 2011 1735 2012 1739
rect 2006 1734 2012 1735
rect 2008 1707 2010 1734
rect 2048 1723 2050 1754
rect 2126 1752 2127 1756
rect 2131 1752 2132 1756
rect 2126 1751 2132 1752
rect 2310 1756 2316 1757
rect 2310 1752 2311 1756
rect 2315 1752 2316 1756
rect 2310 1751 2316 1752
rect 2494 1756 2500 1757
rect 2494 1752 2495 1756
rect 2499 1752 2500 1756
rect 2494 1751 2500 1752
rect 2686 1756 2692 1757
rect 2686 1752 2687 1756
rect 2691 1752 2692 1756
rect 2686 1751 2692 1752
rect 2128 1723 2130 1751
rect 2312 1723 2314 1751
rect 2496 1723 2498 1751
rect 2578 1731 2584 1732
rect 2578 1727 2579 1731
rect 2583 1727 2584 1731
rect 2578 1726 2584 1727
rect 2047 1722 2051 1723
rect 2047 1717 2051 1718
rect 2071 1722 2075 1723
rect 2071 1717 2075 1718
rect 2127 1722 2131 1723
rect 2127 1717 2131 1718
rect 2191 1722 2195 1723
rect 2191 1717 2195 1718
rect 2311 1722 2315 1723
rect 2311 1717 2315 1718
rect 2343 1722 2347 1723
rect 2343 1717 2347 1718
rect 2495 1722 2499 1723
rect 2495 1717 2499 1718
rect 2511 1722 2515 1723
rect 2511 1717 2515 1718
rect 1839 1706 1843 1707
rect 1839 1701 1843 1702
rect 2007 1706 2011 1707
rect 2007 1701 2011 1702
rect 1706 1699 1712 1700
rect 1706 1695 1707 1699
rect 1711 1695 1712 1699
rect 1706 1694 1712 1695
rect 1818 1699 1824 1700
rect 1818 1695 1819 1699
rect 1823 1695 1824 1699
rect 1818 1694 1824 1695
rect 1406 1676 1412 1677
rect 1406 1672 1407 1676
rect 1411 1672 1412 1676
rect 1406 1671 1412 1672
rect 1622 1676 1628 1677
rect 1622 1672 1623 1676
rect 1627 1672 1628 1676
rect 1622 1671 1628 1672
rect 1708 1668 1710 1694
rect 1840 1677 1842 1701
rect 1838 1676 1844 1677
rect 1838 1672 1839 1676
rect 1843 1672 1844 1676
rect 2008 1674 2010 1701
rect 2048 1690 2050 1717
rect 2072 1693 2074 1717
rect 2146 1715 2152 1716
rect 2146 1711 2147 1715
rect 2151 1711 2152 1715
rect 2146 1710 2152 1711
rect 2070 1692 2076 1693
rect 2046 1689 2052 1690
rect 2046 1685 2047 1689
rect 2051 1685 2052 1689
rect 2070 1688 2071 1692
rect 2075 1688 2076 1692
rect 2070 1687 2076 1688
rect 2046 1684 2052 1685
rect 2148 1684 2150 1710
rect 2192 1693 2194 1717
rect 2266 1715 2272 1716
rect 2266 1711 2267 1715
rect 2271 1711 2272 1715
rect 2266 1710 2272 1711
rect 2190 1692 2196 1693
rect 2190 1688 2191 1692
rect 2195 1688 2196 1692
rect 2190 1687 2196 1688
rect 2268 1684 2270 1710
rect 2298 1707 2304 1708
rect 2298 1703 2299 1707
rect 2303 1703 2304 1707
rect 2298 1702 2304 1703
rect 2146 1683 2152 1684
rect 2146 1679 2147 1683
rect 2151 1679 2152 1683
rect 2146 1678 2152 1679
rect 2266 1683 2272 1684
rect 2266 1679 2267 1683
rect 2271 1679 2272 1683
rect 2266 1678 2272 1679
rect 1838 1671 1844 1672
rect 2006 1673 2012 1674
rect 2070 1673 2076 1674
rect 2006 1669 2007 1673
rect 2011 1669 2012 1673
rect 2006 1668 2012 1669
rect 2046 1672 2052 1673
rect 2046 1668 2047 1672
rect 2051 1668 2052 1672
rect 2070 1669 2071 1673
rect 2075 1669 2076 1673
rect 2070 1668 2076 1669
rect 2190 1673 2196 1674
rect 2190 1669 2191 1673
rect 2195 1669 2196 1673
rect 2190 1668 2196 1669
rect 1274 1667 1280 1668
rect 1274 1663 1275 1667
rect 1279 1663 1280 1667
rect 1274 1662 1280 1663
rect 1302 1667 1308 1668
rect 1302 1663 1303 1667
rect 1307 1663 1308 1667
rect 1302 1662 1308 1663
rect 1558 1667 1564 1668
rect 1558 1663 1559 1667
rect 1563 1663 1564 1667
rect 1558 1662 1564 1663
rect 1706 1667 1712 1668
rect 2046 1667 2052 1668
rect 1706 1663 1707 1667
rect 1711 1663 1712 1667
rect 1706 1662 1712 1663
rect 1406 1657 1412 1658
rect 1406 1653 1407 1657
rect 1411 1653 1412 1657
rect 1406 1652 1412 1653
rect 1408 1631 1410 1652
rect 1343 1630 1347 1631
rect 1343 1625 1347 1626
rect 1407 1630 1411 1631
rect 1407 1625 1411 1626
rect 1495 1630 1499 1631
rect 1495 1625 1499 1626
rect 1344 1604 1346 1625
rect 1496 1604 1498 1625
rect 1342 1603 1348 1604
rect 1342 1599 1343 1603
rect 1347 1599 1348 1603
rect 1342 1598 1348 1599
rect 1494 1603 1500 1604
rect 1494 1599 1495 1603
rect 1499 1599 1500 1603
rect 1494 1598 1500 1599
rect 1258 1595 1264 1596
rect 1118 1591 1124 1592
rect 1118 1587 1119 1591
rect 1123 1587 1124 1591
rect 1258 1591 1259 1595
rect 1263 1591 1264 1595
rect 1258 1590 1264 1591
rect 1278 1595 1284 1596
rect 1278 1591 1279 1595
rect 1283 1591 1284 1595
rect 1278 1590 1284 1591
rect 1118 1586 1124 1587
rect 1014 1584 1020 1585
rect 1014 1580 1015 1584
rect 1019 1580 1020 1584
rect 1014 1579 1020 1580
rect 874 1563 880 1564
rect 874 1559 875 1563
rect 879 1559 880 1563
rect 874 1558 880 1559
rect 1016 1551 1018 1579
rect 1120 1560 1122 1586
rect 1182 1584 1188 1585
rect 1182 1580 1183 1584
rect 1187 1580 1188 1584
rect 1182 1579 1188 1580
rect 1118 1559 1124 1560
rect 1118 1555 1119 1559
rect 1123 1555 1124 1559
rect 1118 1554 1124 1555
rect 1184 1551 1186 1579
rect 1280 1572 1282 1590
rect 1342 1584 1348 1585
rect 1342 1580 1343 1584
rect 1347 1580 1348 1584
rect 1342 1579 1348 1580
rect 1494 1584 1500 1585
rect 1494 1580 1495 1584
rect 1499 1580 1500 1584
rect 1494 1579 1500 1580
rect 1278 1571 1284 1572
rect 1278 1567 1279 1571
rect 1283 1567 1284 1571
rect 1278 1566 1284 1567
rect 1344 1551 1346 1579
rect 1350 1559 1356 1560
rect 1350 1555 1351 1559
rect 1355 1555 1356 1559
rect 1350 1554 1356 1555
rect 839 1550 843 1551
rect 839 1545 843 1546
rect 887 1550 891 1551
rect 887 1545 891 1546
rect 1015 1550 1019 1551
rect 1015 1545 1019 1546
rect 1079 1550 1083 1551
rect 1079 1545 1083 1546
rect 1183 1550 1187 1551
rect 1183 1545 1187 1546
rect 1263 1550 1267 1551
rect 1263 1545 1267 1546
rect 1343 1550 1347 1551
rect 1343 1545 1347 1546
rect 730 1543 736 1544
rect 730 1539 731 1543
rect 735 1539 736 1543
rect 730 1538 736 1539
rect 762 1543 768 1544
rect 762 1539 763 1543
rect 767 1539 768 1543
rect 762 1538 768 1539
rect 486 1520 492 1521
rect 486 1516 487 1520
rect 491 1516 492 1520
rect 486 1515 492 1516
rect 686 1520 692 1521
rect 686 1516 687 1520
rect 691 1516 692 1520
rect 686 1515 692 1516
rect 764 1512 766 1538
rect 888 1521 890 1545
rect 1080 1521 1082 1545
rect 1154 1543 1160 1544
rect 1154 1539 1155 1543
rect 1159 1539 1160 1543
rect 1154 1538 1160 1539
rect 886 1520 892 1521
rect 886 1516 887 1520
rect 891 1516 892 1520
rect 886 1515 892 1516
rect 1078 1520 1084 1521
rect 1078 1516 1079 1520
rect 1083 1516 1084 1520
rect 1078 1515 1084 1516
rect 1156 1512 1158 1538
rect 1264 1521 1266 1545
rect 1262 1520 1268 1521
rect 1262 1516 1263 1520
rect 1267 1516 1268 1520
rect 1262 1515 1268 1516
rect 1352 1512 1354 1554
rect 1496 1551 1498 1579
rect 1560 1564 1562 1662
rect 1622 1657 1628 1658
rect 1622 1653 1623 1657
rect 1627 1653 1628 1657
rect 1622 1652 1628 1653
rect 1838 1657 1844 1658
rect 1838 1653 1839 1657
rect 1843 1653 1844 1657
rect 1838 1652 1844 1653
rect 2006 1656 2012 1657
rect 2006 1652 2007 1656
rect 2011 1652 2012 1656
rect 1624 1631 1626 1652
rect 1840 1631 1842 1652
rect 2006 1651 2012 1652
rect 2008 1631 2010 1651
rect 2048 1647 2050 1667
rect 2072 1647 2074 1668
rect 2192 1647 2194 1668
rect 2047 1646 2051 1647
rect 2047 1641 2051 1642
rect 2071 1646 2075 1647
rect 2071 1641 2075 1642
rect 2191 1646 2195 1647
rect 2191 1641 2195 1642
rect 1623 1630 1627 1631
rect 1623 1625 1627 1626
rect 1639 1630 1643 1631
rect 1639 1625 1643 1626
rect 1783 1630 1787 1631
rect 1783 1625 1787 1626
rect 1839 1630 1843 1631
rect 1839 1625 1843 1626
rect 1903 1630 1907 1631
rect 1903 1625 1907 1626
rect 2007 1630 2011 1631
rect 2007 1625 2011 1626
rect 1640 1604 1642 1625
rect 1784 1604 1786 1625
rect 1904 1604 1906 1625
rect 2008 1605 2010 1625
rect 2048 1621 2050 1641
rect 2046 1620 2052 1621
rect 2072 1620 2074 1641
rect 2046 1616 2047 1620
rect 2051 1616 2052 1620
rect 2046 1615 2052 1616
rect 2070 1619 2076 1620
rect 2070 1615 2071 1619
rect 2075 1615 2076 1619
rect 2070 1614 2076 1615
rect 2300 1612 2302 1702
rect 2344 1693 2346 1717
rect 2418 1715 2424 1716
rect 2418 1711 2419 1715
rect 2423 1711 2424 1715
rect 2418 1710 2424 1711
rect 2342 1692 2348 1693
rect 2342 1688 2343 1692
rect 2347 1688 2348 1692
rect 2342 1687 2348 1688
rect 2420 1684 2422 1710
rect 2512 1693 2514 1717
rect 2510 1692 2516 1693
rect 2510 1688 2511 1692
rect 2515 1688 2516 1692
rect 2510 1687 2516 1688
rect 2580 1684 2582 1726
rect 2688 1723 2690 1751
rect 2772 1736 2774 1838
rect 2830 1833 2836 1834
rect 2830 1829 2831 1833
rect 2835 1829 2836 1833
rect 2830 1828 2836 1829
rect 2832 1803 2834 1828
rect 2831 1802 2835 1803
rect 2831 1797 2835 1798
rect 2872 1768 2874 1870
rect 2908 1844 2910 1870
rect 2992 1853 2994 1877
rect 3066 1875 3072 1876
rect 3066 1871 3067 1875
rect 3071 1871 3072 1875
rect 3066 1870 3072 1871
rect 2990 1852 2996 1853
rect 2990 1848 2991 1852
rect 2995 1848 2996 1852
rect 2990 1847 2996 1848
rect 3068 1844 3070 1870
rect 3184 1853 3186 1877
rect 3258 1875 3264 1876
rect 3258 1871 3259 1875
rect 3263 1871 3264 1875
rect 3258 1870 3264 1871
rect 3182 1852 3188 1853
rect 3182 1848 3183 1852
rect 3187 1848 3188 1852
rect 3182 1847 3188 1848
rect 3260 1844 3262 1870
rect 3400 1853 3402 1877
rect 3474 1875 3480 1876
rect 3474 1871 3475 1875
rect 3479 1871 3480 1875
rect 3474 1870 3480 1871
rect 3398 1852 3404 1853
rect 3398 1848 3399 1852
rect 3403 1848 3404 1852
rect 3398 1847 3404 1848
rect 3476 1844 3478 1870
rect 3632 1853 3634 1877
rect 3630 1852 3636 1853
rect 3630 1848 3631 1852
rect 3635 1848 3636 1852
rect 3630 1847 3636 1848
rect 2906 1843 2912 1844
rect 2906 1839 2907 1843
rect 2911 1839 2912 1843
rect 2906 1838 2912 1839
rect 3066 1843 3072 1844
rect 3066 1839 3067 1843
rect 3071 1839 3072 1843
rect 3066 1838 3072 1839
rect 3258 1843 3264 1844
rect 3258 1839 3259 1843
rect 3263 1839 3264 1843
rect 3258 1838 3264 1839
rect 3474 1843 3480 1844
rect 3474 1839 3475 1843
rect 3479 1839 3480 1843
rect 3474 1838 3480 1839
rect 2990 1833 2996 1834
rect 2990 1829 2991 1833
rect 2995 1829 2996 1833
rect 2990 1828 2996 1829
rect 3182 1833 3188 1834
rect 3182 1829 3183 1833
rect 3187 1829 3188 1833
rect 3182 1828 3188 1829
rect 3398 1833 3404 1834
rect 3398 1829 3399 1833
rect 3403 1829 3404 1833
rect 3398 1828 3404 1829
rect 3630 1833 3636 1834
rect 3630 1829 3631 1833
rect 3635 1829 3636 1833
rect 3630 1828 3636 1829
rect 2992 1803 2994 1828
rect 3184 1803 3186 1828
rect 3400 1803 3402 1828
rect 3632 1803 3634 1828
rect 2879 1802 2883 1803
rect 2879 1797 2883 1798
rect 2991 1802 2995 1803
rect 2991 1797 2995 1798
rect 3071 1802 3075 1803
rect 3071 1797 3075 1798
rect 3183 1802 3187 1803
rect 3183 1797 3187 1798
rect 3263 1802 3267 1803
rect 3263 1797 3267 1798
rect 3399 1802 3403 1803
rect 3399 1797 3403 1798
rect 3463 1802 3467 1803
rect 3463 1797 3467 1798
rect 3631 1802 3635 1803
rect 3631 1797 3635 1798
rect 3663 1802 3667 1803
rect 3663 1797 3667 1798
rect 2880 1776 2882 1797
rect 3072 1776 3074 1797
rect 3264 1776 3266 1797
rect 3464 1776 3466 1797
rect 3664 1776 3666 1797
rect 2878 1775 2884 1776
rect 2878 1771 2879 1775
rect 2883 1771 2884 1775
rect 2878 1770 2884 1771
rect 3070 1775 3076 1776
rect 3070 1771 3071 1775
rect 3075 1771 3076 1775
rect 3070 1770 3076 1771
rect 3262 1775 3268 1776
rect 3262 1771 3263 1775
rect 3267 1771 3268 1775
rect 3262 1770 3268 1771
rect 3462 1775 3468 1776
rect 3462 1771 3463 1775
rect 3467 1771 3468 1775
rect 3462 1770 3468 1771
rect 3662 1775 3668 1776
rect 3662 1771 3663 1775
rect 3667 1771 3668 1775
rect 3662 1770 3668 1771
rect 2870 1767 2876 1768
rect 2798 1763 2804 1764
rect 2798 1759 2799 1763
rect 2803 1759 2804 1763
rect 2870 1763 2871 1767
rect 2875 1763 2876 1767
rect 2870 1762 2876 1763
rect 3158 1767 3164 1768
rect 3158 1763 3159 1767
rect 3163 1763 3164 1767
rect 3158 1762 3164 1763
rect 3346 1767 3352 1768
rect 3346 1763 3347 1767
rect 3351 1763 3352 1767
rect 3346 1762 3352 1763
rect 3738 1763 3744 1764
rect 2798 1758 2804 1759
rect 2770 1735 2776 1736
rect 2770 1731 2771 1735
rect 2775 1731 2776 1735
rect 2770 1730 2776 1731
rect 2687 1722 2691 1723
rect 2687 1717 2691 1718
rect 2688 1693 2690 1717
rect 2800 1716 2802 1758
rect 2878 1756 2884 1757
rect 2878 1752 2879 1756
rect 2883 1752 2884 1756
rect 2878 1751 2884 1752
rect 3070 1756 3076 1757
rect 3070 1752 3071 1756
rect 3075 1752 3076 1756
rect 3070 1751 3076 1752
rect 2880 1723 2882 1751
rect 3072 1723 3074 1751
rect 3160 1736 3162 1762
rect 3262 1756 3268 1757
rect 3262 1752 3263 1756
rect 3267 1752 3268 1756
rect 3262 1751 3268 1752
rect 3158 1735 3164 1736
rect 3158 1731 3159 1735
rect 3163 1731 3164 1735
rect 3158 1730 3164 1731
rect 3264 1723 3266 1751
rect 3348 1736 3350 1762
rect 3738 1759 3739 1763
rect 3743 1759 3744 1763
rect 3738 1758 3744 1759
rect 3462 1756 3468 1757
rect 3462 1752 3463 1756
rect 3467 1752 3468 1756
rect 3462 1751 3468 1752
rect 3662 1756 3668 1757
rect 3662 1752 3663 1756
rect 3667 1752 3668 1756
rect 3662 1751 3668 1752
rect 3346 1735 3352 1736
rect 3346 1731 3347 1735
rect 3351 1731 3352 1735
rect 3346 1730 3352 1731
rect 3464 1723 3466 1751
rect 3514 1731 3520 1732
rect 3514 1727 3515 1731
rect 3519 1727 3520 1731
rect 3514 1726 3520 1727
rect 2871 1722 2875 1723
rect 2871 1717 2875 1718
rect 2879 1722 2883 1723
rect 2879 1717 2883 1718
rect 3063 1722 3067 1723
rect 3063 1717 3067 1718
rect 3071 1722 3075 1723
rect 3071 1717 3075 1718
rect 3255 1722 3259 1723
rect 3255 1717 3259 1718
rect 3263 1722 3267 1723
rect 3263 1717 3267 1718
rect 3447 1722 3451 1723
rect 3447 1717 3451 1718
rect 3463 1722 3467 1723
rect 3463 1717 3467 1718
rect 2790 1715 2796 1716
rect 2790 1711 2791 1715
rect 2795 1711 2796 1715
rect 2790 1710 2796 1711
rect 2798 1715 2804 1716
rect 2798 1711 2799 1715
rect 2803 1711 2804 1715
rect 2798 1710 2804 1711
rect 2686 1692 2692 1693
rect 2686 1688 2687 1692
rect 2691 1688 2692 1692
rect 2686 1687 2692 1688
rect 2792 1684 2794 1710
rect 2872 1693 2874 1717
rect 3064 1693 3066 1717
rect 3118 1715 3124 1716
rect 3118 1711 3119 1715
rect 3123 1714 3124 1715
rect 3138 1715 3144 1716
rect 3123 1711 3126 1714
rect 3118 1710 3126 1711
rect 3138 1711 3139 1715
rect 3143 1711 3144 1715
rect 3138 1710 3144 1711
rect 2870 1692 2876 1693
rect 2870 1688 2871 1692
rect 2875 1688 2876 1692
rect 2870 1687 2876 1688
rect 3062 1692 3068 1693
rect 3062 1688 3063 1692
rect 3067 1688 3068 1692
rect 3062 1687 3068 1688
rect 2418 1683 2424 1684
rect 2418 1679 2419 1683
rect 2423 1679 2424 1683
rect 2418 1678 2424 1679
rect 2578 1683 2584 1684
rect 2578 1679 2579 1683
rect 2583 1679 2584 1683
rect 2578 1678 2584 1679
rect 2654 1683 2660 1684
rect 2654 1679 2655 1683
rect 2659 1679 2660 1683
rect 2654 1678 2660 1679
rect 2790 1683 2796 1684
rect 2790 1679 2791 1683
rect 2795 1679 2796 1683
rect 2790 1678 2796 1679
rect 2342 1673 2348 1674
rect 2342 1669 2343 1673
rect 2347 1669 2348 1673
rect 2342 1668 2348 1669
rect 2510 1673 2516 1674
rect 2510 1669 2511 1673
rect 2515 1669 2516 1673
rect 2510 1668 2516 1669
rect 2344 1647 2346 1668
rect 2512 1647 2514 1668
rect 2335 1646 2339 1647
rect 2335 1641 2339 1642
rect 2343 1646 2347 1647
rect 2343 1641 2347 1642
rect 2511 1646 2515 1647
rect 2511 1641 2515 1642
rect 2599 1646 2603 1647
rect 2599 1641 2603 1642
rect 2336 1620 2338 1641
rect 2600 1620 2602 1641
rect 2334 1619 2340 1620
rect 2334 1615 2335 1619
rect 2339 1615 2340 1619
rect 2334 1614 2340 1615
rect 2598 1619 2604 1620
rect 2598 1615 2599 1619
rect 2603 1615 2604 1619
rect 2598 1614 2604 1615
rect 2298 1611 2304 1612
rect 2146 1607 2152 1608
rect 2006 1604 2012 1605
rect 1638 1603 1644 1604
rect 1638 1599 1639 1603
rect 1643 1599 1644 1603
rect 1638 1598 1644 1599
rect 1782 1603 1788 1604
rect 1782 1599 1783 1603
rect 1787 1599 1788 1603
rect 1782 1598 1788 1599
rect 1902 1603 1908 1604
rect 1902 1599 1903 1603
rect 1907 1599 1908 1603
rect 2006 1600 2007 1604
rect 2011 1600 2012 1604
rect 2006 1599 2012 1600
rect 2046 1603 2052 1604
rect 2046 1599 2047 1603
rect 2051 1599 2052 1603
rect 2146 1603 2147 1607
rect 2151 1603 2152 1607
rect 2298 1607 2299 1611
rect 2303 1607 2304 1611
rect 2298 1606 2304 1607
rect 2146 1602 2152 1603
rect 1902 1598 1908 1599
rect 2046 1598 2052 1599
rect 2070 1600 2076 1601
rect 1570 1591 1576 1592
rect 1570 1587 1571 1591
rect 1575 1587 1576 1591
rect 1570 1586 1576 1587
rect 1714 1591 1720 1592
rect 1714 1587 1715 1591
rect 1719 1587 1720 1591
rect 1714 1586 1720 1587
rect 1858 1591 1864 1592
rect 1858 1587 1859 1591
rect 1863 1587 1864 1591
rect 1858 1586 1864 1587
rect 2006 1587 2012 1588
rect 1572 1564 1574 1586
rect 1638 1584 1644 1585
rect 1638 1580 1639 1584
rect 1643 1580 1644 1584
rect 1638 1579 1644 1580
rect 1558 1563 1564 1564
rect 1558 1559 1559 1563
rect 1563 1559 1564 1563
rect 1558 1558 1564 1559
rect 1570 1563 1576 1564
rect 1570 1559 1571 1563
rect 1575 1559 1576 1563
rect 1570 1558 1576 1559
rect 1640 1551 1642 1579
rect 1716 1564 1718 1586
rect 1782 1584 1788 1585
rect 1782 1580 1783 1584
rect 1787 1580 1788 1584
rect 1782 1579 1788 1580
rect 1714 1563 1720 1564
rect 1714 1559 1715 1563
rect 1719 1559 1720 1563
rect 1714 1558 1720 1559
rect 1784 1551 1786 1579
rect 1860 1564 1862 1586
rect 1902 1584 1908 1585
rect 1902 1580 1903 1584
rect 1907 1580 1908 1584
rect 2006 1583 2007 1587
rect 2011 1583 2012 1587
rect 2006 1582 2012 1583
rect 1902 1579 1908 1580
rect 1858 1563 1864 1564
rect 1858 1559 1859 1563
rect 1863 1559 1864 1563
rect 1858 1558 1864 1559
rect 1904 1551 1906 1579
rect 2008 1551 2010 1582
rect 2048 1567 2050 1598
rect 2070 1596 2071 1600
rect 2075 1596 2076 1600
rect 2070 1595 2076 1596
rect 2072 1567 2074 1595
rect 2148 1580 2150 1602
rect 2334 1600 2340 1601
rect 2334 1596 2335 1600
rect 2339 1596 2340 1600
rect 2334 1595 2340 1596
rect 2598 1600 2604 1601
rect 2598 1596 2599 1600
rect 2603 1596 2604 1600
rect 2598 1595 2604 1596
rect 2146 1579 2152 1580
rect 2146 1575 2147 1579
rect 2151 1575 2152 1579
rect 2146 1574 2152 1575
rect 2336 1567 2338 1595
rect 2600 1567 2602 1595
rect 2656 1580 2658 1678
rect 2686 1673 2692 1674
rect 2686 1669 2687 1673
rect 2691 1669 2692 1673
rect 2686 1668 2692 1669
rect 2870 1673 2876 1674
rect 2870 1669 2871 1673
rect 2875 1669 2876 1673
rect 2870 1668 2876 1669
rect 3062 1673 3068 1674
rect 3062 1669 3063 1673
rect 3067 1669 3068 1673
rect 3062 1668 3068 1669
rect 2688 1647 2690 1668
rect 2872 1647 2874 1668
rect 3064 1647 3066 1668
rect 2687 1646 2691 1647
rect 2687 1641 2691 1642
rect 2839 1646 2843 1647
rect 2839 1641 2843 1642
rect 2871 1646 2875 1647
rect 2871 1641 2875 1642
rect 3047 1646 3051 1647
rect 3047 1641 3051 1642
rect 3063 1646 3067 1647
rect 3063 1641 3067 1642
rect 2840 1620 2842 1641
rect 3048 1620 3050 1641
rect 2838 1619 2844 1620
rect 2838 1615 2839 1619
rect 2843 1615 2844 1619
rect 2838 1614 2844 1615
rect 3046 1619 3052 1620
rect 3046 1615 3047 1619
rect 3051 1615 3052 1619
rect 3046 1614 3052 1615
rect 3124 1612 3126 1710
rect 3140 1684 3142 1710
rect 3256 1693 3258 1717
rect 3330 1715 3336 1716
rect 3330 1711 3331 1715
rect 3335 1711 3336 1715
rect 3330 1710 3336 1711
rect 3254 1692 3260 1693
rect 3254 1688 3255 1692
rect 3259 1688 3260 1692
rect 3254 1687 3260 1688
rect 3332 1684 3334 1710
rect 3448 1693 3450 1717
rect 3446 1692 3452 1693
rect 3446 1688 3447 1692
rect 3451 1688 3452 1692
rect 3446 1687 3452 1688
rect 3516 1684 3518 1726
rect 3664 1723 3666 1751
rect 3647 1722 3651 1723
rect 3647 1717 3651 1718
rect 3663 1722 3667 1723
rect 3663 1717 3667 1718
rect 3648 1693 3650 1717
rect 3740 1716 3742 1758
rect 3752 1736 3754 1930
rect 3774 1924 3780 1925
rect 3774 1920 3775 1924
rect 3779 1920 3780 1924
rect 3774 1919 3780 1920
rect 3776 1883 3778 1919
rect 3832 1904 3834 2094
rect 3942 2091 3948 2092
rect 3838 2088 3844 2089
rect 3838 2084 3839 2088
rect 3843 2084 3844 2088
rect 3942 2087 3943 2091
rect 3947 2087 3948 2091
rect 3942 2086 3948 2087
rect 3838 2083 3844 2084
rect 3840 2051 3842 2083
rect 3944 2051 3946 2086
rect 3839 2050 3843 2051
rect 3839 2045 3843 2046
rect 3943 2050 3947 2051
rect 3943 2045 3947 2046
rect 3840 2021 3842 2045
rect 3906 2043 3912 2044
rect 3906 2039 3907 2043
rect 3911 2039 3912 2043
rect 3906 2038 3912 2039
rect 3838 2020 3844 2021
rect 3838 2016 3839 2020
rect 3843 2016 3844 2020
rect 3838 2015 3844 2016
rect 3838 2001 3844 2002
rect 3838 1997 3839 2001
rect 3843 1997 3844 2001
rect 3838 1996 3844 1997
rect 3840 1971 3842 1996
rect 3908 1993 3910 2038
rect 3944 2018 3946 2045
rect 3942 2017 3948 2018
rect 3942 2013 3943 2017
rect 3947 2013 3948 2017
rect 3942 2012 3948 2013
rect 3942 2000 3948 2001
rect 3942 1996 3943 2000
rect 3947 1996 3948 2000
rect 3942 1995 3948 1996
rect 3908 1991 3918 1993
rect 3839 1970 3843 1971
rect 3839 1965 3843 1966
rect 3830 1903 3836 1904
rect 3830 1899 3831 1903
rect 3835 1899 3836 1903
rect 3830 1898 3836 1899
rect 3775 1882 3779 1883
rect 3775 1877 3779 1878
rect 3839 1882 3843 1883
rect 3839 1877 3843 1878
rect 3840 1853 3842 1877
rect 3906 1875 3912 1876
rect 3906 1871 3907 1875
rect 3911 1871 3912 1875
rect 3906 1870 3912 1871
rect 3838 1852 3844 1853
rect 3838 1848 3839 1852
rect 3843 1848 3844 1852
rect 3838 1847 3844 1848
rect 3838 1833 3844 1834
rect 3838 1829 3839 1833
rect 3843 1829 3844 1833
rect 3838 1828 3844 1829
rect 3840 1803 3842 1828
rect 3839 1802 3843 1803
rect 3839 1797 3843 1798
rect 3840 1776 3842 1797
rect 3838 1775 3844 1776
rect 3838 1771 3839 1775
rect 3843 1771 3844 1775
rect 3908 1772 3910 1870
rect 3916 1844 3918 1991
rect 3944 1971 3946 1995
rect 3943 1970 3947 1971
rect 3943 1965 3947 1966
rect 3944 1945 3946 1965
rect 3942 1944 3948 1945
rect 3942 1940 3943 1944
rect 3947 1940 3948 1944
rect 3942 1939 3948 1940
rect 3942 1927 3948 1928
rect 3942 1923 3943 1927
rect 3947 1923 3948 1927
rect 3942 1922 3948 1923
rect 3944 1883 3946 1922
rect 3943 1882 3947 1883
rect 3943 1877 3947 1878
rect 3944 1850 3946 1877
rect 3942 1849 3948 1850
rect 3942 1845 3943 1849
rect 3947 1845 3948 1849
rect 3942 1844 3948 1845
rect 3914 1843 3920 1844
rect 3914 1839 3915 1843
rect 3919 1839 3920 1843
rect 3914 1838 3920 1839
rect 3942 1832 3948 1833
rect 3942 1828 3943 1832
rect 3947 1828 3948 1832
rect 3942 1827 3948 1828
rect 3944 1803 3946 1827
rect 3943 1802 3947 1803
rect 3943 1797 3947 1798
rect 3944 1777 3946 1797
rect 3942 1776 3948 1777
rect 3942 1772 3943 1776
rect 3947 1772 3948 1776
rect 3838 1770 3844 1771
rect 3906 1771 3912 1772
rect 3942 1771 3948 1772
rect 3906 1767 3907 1771
rect 3911 1767 3912 1771
rect 3906 1766 3912 1767
rect 3942 1759 3948 1760
rect 3838 1756 3844 1757
rect 3838 1752 3839 1756
rect 3843 1752 3844 1756
rect 3942 1755 3943 1759
rect 3947 1755 3948 1759
rect 3942 1754 3948 1755
rect 3838 1751 3844 1752
rect 3750 1735 3756 1736
rect 3750 1731 3751 1735
rect 3755 1731 3756 1735
rect 3750 1730 3756 1731
rect 3840 1723 3842 1751
rect 3906 1731 3912 1732
rect 3906 1727 3907 1731
rect 3911 1727 3912 1731
rect 3906 1726 3912 1727
rect 3839 1722 3843 1723
rect 3839 1717 3843 1718
rect 3738 1715 3744 1716
rect 3738 1711 3739 1715
rect 3743 1711 3744 1715
rect 3738 1710 3744 1711
rect 3840 1693 3842 1717
rect 3646 1692 3652 1693
rect 3646 1688 3647 1692
rect 3651 1688 3652 1692
rect 3646 1687 3652 1688
rect 3838 1692 3844 1693
rect 3838 1688 3839 1692
rect 3843 1688 3844 1692
rect 3838 1687 3844 1688
rect 3908 1684 3910 1726
rect 3944 1723 3946 1754
rect 3943 1722 3947 1723
rect 3943 1717 3947 1718
rect 3914 1715 3920 1716
rect 3914 1711 3915 1715
rect 3919 1711 3920 1715
rect 3914 1710 3920 1711
rect 3138 1683 3144 1684
rect 3138 1679 3139 1683
rect 3143 1679 3144 1683
rect 3138 1678 3144 1679
rect 3330 1683 3336 1684
rect 3330 1679 3331 1683
rect 3335 1679 3336 1683
rect 3330 1678 3336 1679
rect 3514 1683 3520 1684
rect 3514 1679 3515 1683
rect 3519 1679 3520 1683
rect 3514 1678 3520 1679
rect 3614 1683 3620 1684
rect 3614 1679 3615 1683
rect 3619 1679 3620 1683
rect 3614 1678 3620 1679
rect 3906 1683 3912 1684
rect 3906 1679 3907 1683
rect 3911 1679 3912 1683
rect 3906 1678 3912 1679
rect 3254 1673 3260 1674
rect 3254 1669 3255 1673
rect 3259 1669 3260 1673
rect 3254 1668 3260 1669
rect 3446 1673 3452 1674
rect 3446 1669 3447 1673
rect 3451 1669 3452 1673
rect 3446 1668 3452 1669
rect 3256 1647 3258 1668
rect 3448 1647 3450 1668
rect 3231 1646 3235 1647
rect 3231 1641 3235 1642
rect 3255 1646 3259 1647
rect 3255 1641 3259 1642
rect 3399 1646 3403 1647
rect 3399 1641 3403 1642
rect 3447 1646 3451 1647
rect 3447 1641 3451 1642
rect 3551 1646 3555 1647
rect 3551 1641 3555 1642
rect 3232 1620 3234 1641
rect 3400 1620 3402 1641
rect 3552 1620 3554 1641
rect 3230 1619 3236 1620
rect 3230 1615 3231 1619
rect 3235 1615 3236 1619
rect 3230 1614 3236 1615
rect 3398 1619 3404 1620
rect 3398 1615 3399 1619
rect 3403 1615 3404 1619
rect 3398 1614 3404 1615
rect 3550 1619 3556 1620
rect 3550 1615 3551 1619
rect 3555 1615 3556 1619
rect 3550 1614 3556 1615
rect 3122 1611 3128 1612
rect 2674 1607 2680 1608
rect 2674 1603 2675 1607
rect 2679 1603 2680 1607
rect 2674 1602 2680 1603
rect 2914 1607 2920 1608
rect 2914 1603 2915 1607
rect 2919 1603 2920 1607
rect 3122 1607 3123 1611
rect 3127 1607 3128 1611
rect 3122 1606 3128 1607
rect 3130 1611 3136 1612
rect 3130 1607 3131 1611
rect 3135 1607 3136 1611
rect 3130 1606 3136 1607
rect 3354 1611 3360 1612
rect 3354 1607 3355 1611
rect 3359 1607 3360 1611
rect 3354 1606 3360 1607
rect 2914 1602 2920 1603
rect 2654 1579 2660 1580
rect 2654 1575 2655 1579
rect 2659 1575 2660 1579
rect 2654 1574 2660 1575
rect 2047 1566 2051 1567
rect 2047 1561 2051 1562
rect 2071 1566 2075 1567
rect 2071 1561 2075 1562
rect 2335 1566 2339 1567
rect 2335 1561 2339 1562
rect 2583 1566 2587 1567
rect 2583 1561 2587 1562
rect 2599 1566 2603 1567
rect 2599 1561 2603 1562
rect 1447 1550 1451 1551
rect 1447 1545 1451 1546
rect 1495 1550 1499 1551
rect 1495 1545 1499 1546
rect 1623 1550 1627 1551
rect 1623 1545 1627 1546
rect 1639 1550 1643 1551
rect 1639 1545 1643 1546
rect 1783 1550 1787 1551
rect 1783 1545 1787 1546
rect 1807 1550 1811 1551
rect 1807 1545 1811 1546
rect 1903 1550 1907 1551
rect 1903 1545 1907 1546
rect 2007 1550 2011 1551
rect 2007 1545 2011 1546
rect 1398 1535 1404 1536
rect 1398 1531 1399 1535
rect 1403 1531 1404 1535
rect 1398 1530 1404 1531
rect 1400 1512 1402 1530
rect 1448 1521 1450 1545
rect 1530 1543 1536 1544
rect 1530 1539 1531 1543
rect 1535 1539 1536 1543
rect 1530 1538 1536 1539
rect 1446 1520 1452 1521
rect 1446 1516 1447 1520
rect 1451 1516 1452 1520
rect 1446 1515 1452 1516
rect 1532 1512 1534 1538
rect 1624 1521 1626 1545
rect 1706 1543 1712 1544
rect 1706 1539 1707 1543
rect 1711 1539 1712 1543
rect 1706 1538 1712 1539
rect 1622 1520 1628 1521
rect 1622 1516 1623 1520
rect 1627 1516 1628 1520
rect 1622 1515 1628 1516
rect 1708 1512 1710 1538
rect 1808 1521 1810 1545
rect 1862 1543 1868 1544
rect 1862 1539 1863 1543
rect 1867 1539 1868 1543
rect 1862 1538 1868 1539
rect 1806 1520 1812 1521
rect 1806 1516 1807 1520
rect 1811 1516 1812 1520
rect 1806 1515 1812 1516
rect 258 1511 264 1512
rect 258 1507 259 1511
rect 263 1507 264 1511
rect 258 1506 264 1507
rect 370 1511 376 1512
rect 370 1507 371 1511
rect 375 1507 376 1511
rect 370 1506 376 1507
rect 390 1511 396 1512
rect 390 1507 391 1511
rect 395 1507 396 1511
rect 390 1506 396 1507
rect 762 1511 768 1512
rect 762 1507 763 1511
rect 767 1507 768 1511
rect 762 1506 768 1507
rect 838 1511 844 1512
rect 838 1507 839 1511
rect 843 1507 844 1511
rect 838 1506 844 1507
rect 1154 1511 1160 1512
rect 1154 1507 1155 1511
rect 1159 1507 1160 1511
rect 1154 1506 1160 1507
rect 1350 1511 1356 1512
rect 1350 1507 1351 1511
rect 1355 1507 1356 1511
rect 1350 1506 1356 1507
rect 1398 1511 1404 1512
rect 1398 1507 1399 1511
rect 1403 1507 1404 1511
rect 1398 1506 1404 1507
rect 1530 1511 1536 1512
rect 1530 1507 1531 1511
rect 1535 1507 1536 1511
rect 1530 1506 1536 1507
rect 1706 1511 1712 1512
rect 1706 1507 1707 1511
rect 1711 1507 1712 1511
rect 1706 1506 1712 1507
rect 294 1501 300 1502
rect 294 1497 295 1501
rect 299 1497 300 1501
rect 294 1496 300 1497
rect 486 1501 492 1502
rect 486 1497 487 1501
rect 491 1497 492 1501
rect 486 1496 492 1497
rect 686 1501 692 1502
rect 686 1497 687 1501
rect 691 1497 692 1501
rect 686 1496 692 1497
rect 296 1475 298 1496
rect 488 1475 490 1496
rect 688 1475 690 1496
rect 295 1474 299 1475
rect 295 1469 299 1470
rect 359 1474 363 1475
rect 359 1469 363 1470
rect 487 1474 491 1475
rect 487 1469 491 1470
rect 567 1474 571 1475
rect 567 1469 571 1470
rect 687 1474 691 1475
rect 687 1469 691 1470
rect 783 1474 787 1475
rect 783 1469 787 1470
rect 360 1448 362 1469
rect 568 1448 570 1469
rect 784 1448 786 1469
rect 358 1447 364 1448
rect 358 1443 359 1447
rect 363 1443 364 1447
rect 358 1442 364 1443
rect 566 1447 572 1448
rect 566 1443 567 1447
rect 571 1443 572 1447
rect 566 1442 572 1443
rect 782 1447 788 1448
rect 782 1443 783 1447
rect 787 1443 788 1447
rect 782 1442 788 1443
rect 250 1439 256 1440
rect 250 1435 251 1439
rect 255 1435 256 1439
rect 250 1434 256 1435
rect 274 1439 280 1440
rect 274 1435 275 1439
rect 279 1435 280 1439
rect 274 1434 280 1435
rect 442 1439 448 1440
rect 442 1435 443 1439
rect 447 1435 448 1439
rect 442 1434 448 1435
rect 110 1431 116 1432
rect 110 1427 111 1431
rect 115 1427 116 1431
rect 110 1426 116 1427
rect 174 1428 180 1429
rect 112 1399 114 1426
rect 174 1424 175 1428
rect 179 1424 180 1428
rect 174 1423 180 1424
rect 176 1399 178 1423
rect 276 1408 278 1434
rect 358 1428 364 1429
rect 358 1424 359 1428
rect 363 1424 364 1428
rect 358 1423 364 1424
rect 274 1407 280 1408
rect 274 1403 275 1407
rect 279 1403 280 1407
rect 274 1402 280 1403
rect 360 1399 362 1423
rect 402 1403 408 1404
rect 402 1399 403 1403
rect 407 1399 408 1403
rect 111 1398 115 1399
rect 111 1393 115 1394
rect 175 1398 179 1399
rect 175 1393 179 1394
rect 327 1398 331 1399
rect 327 1393 331 1394
rect 359 1398 363 1399
rect 402 1398 408 1399
rect 359 1393 363 1394
rect 112 1366 114 1393
rect 328 1369 330 1393
rect 326 1368 332 1369
rect 110 1365 116 1366
rect 110 1361 111 1365
rect 115 1361 116 1365
rect 326 1364 327 1368
rect 331 1364 332 1368
rect 326 1363 332 1364
rect 110 1360 116 1361
rect 404 1360 406 1398
rect 444 1392 446 1434
rect 566 1428 572 1429
rect 566 1424 567 1428
rect 571 1424 572 1428
rect 566 1423 572 1424
rect 782 1428 788 1429
rect 782 1424 783 1428
rect 787 1424 788 1428
rect 782 1423 788 1424
rect 568 1399 570 1423
rect 784 1399 786 1423
rect 840 1408 842 1506
rect 886 1501 892 1502
rect 886 1497 887 1501
rect 891 1497 892 1501
rect 886 1496 892 1497
rect 1078 1501 1084 1502
rect 1078 1497 1079 1501
rect 1083 1497 1084 1501
rect 1078 1496 1084 1497
rect 1262 1501 1268 1502
rect 1262 1497 1263 1501
rect 1267 1497 1268 1501
rect 1262 1496 1268 1497
rect 1446 1501 1452 1502
rect 1446 1497 1447 1501
rect 1451 1497 1452 1501
rect 1446 1496 1452 1497
rect 1622 1501 1628 1502
rect 1622 1497 1623 1501
rect 1627 1497 1628 1501
rect 1622 1496 1628 1497
rect 1806 1501 1812 1502
rect 1806 1497 1807 1501
rect 1811 1497 1812 1501
rect 1806 1496 1812 1497
rect 888 1475 890 1496
rect 1080 1475 1082 1496
rect 1264 1475 1266 1496
rect 1448 1475 1450 1496
rect 1624 1475 1626 1496
rect 1808 1475 1810 1496
rect 887 1474 891 1475
rect 887 1469 891 1470
rect 1007 1474 1011 1475
rect 1007 1469 1011 1470
rect 1079 1474 1083 1475
rect 1079 1469 1083 1470
rect 1231 1474 1235 1475
rect 1231 1469 1235 1470
rect 1263 1474 1267 1475
rect 1263 1469 1267 1470
rect 1447 1474 1451 1475
rect 1447 1469 1451 1470
rect 1463 1474 1467 1475
rect 1463 1469 1467 1470
rect 1623 1474 1627 1475
rect 1623 1469 1627 1470
rect 1695 1474 1699 1475
rect 1695 1469 1699 1470
rect 1807 1474 1811 1475
rect 1807 1469 1811 1470
rect 1008 1448 1010 1469
rect 1232 1448 1234 1469
rect 1464 1448 1466 1469
rect 1696 1448 1698 1469
rect 1006 1447 1012 1448
rect 1006 1443 1007 1447
rect 1011 1443 1012 1447
rect 1006 1442 1012 1443
rect 1230 1447 1236 1448
rect 1230 1443 1231 1447
rect 1235 1443 1236 1447
rect 1230 1442 1236 1443
rect 1462 1447 1468 1448
rect 1462 1443 1463 1447
rect 1467 1443 1468 1447
rect 1462 1442 1468 1443
rect 1694 1447 1700 1448
rect 1694 1443 1695 1447
rect 1699 1443 1700 1447
rect 1694 1442 1700 1443
rect 1864 1440 1866 1538
rect 2008 1518 2010 1545
rect 2048 1534 2050 1561
rect 2584 1537 2586 1561
rect 2676 1560 2678 1602
rect 2838 1600 2844 1601
rect 2838 1596 2839 1600
rect 2843 1596 2844 1600
rect 2838 1595 2844 1596
rect 2840 1567 2842 1595
rect 2916 1580 2918 1602
rect 3046 1600 3052 1601
rect 3046 1596 3047 1600
rect 3051 1596 3052 1600
rect 3046 1595 3052 1596
rect 2914 1579 2920 1580
rect 2914 1575 2915 1579
rect 2919 1575 2920 1579
rect 2914 1574 2920 1575
rect 3048 1567 3050 1595
rect 3132 1588 3134 1606
rect 3230 1600 3236 1601
rect 3230 1596 3231 1600
rect 3235 1596 3236 1600
rect 3230 1595 3236 1596
rect 3130 1587 3136 1588
rect 3130 1583 3131 1587
rect 3135 1583 3136 1587
rect 3130 1582 3136 1583
rect 3232 1567 3234 1595
rect 3356 1580 3358 1606
rect 3398 1600 3404 1601
rect 3398 1596 3399 1600
rect 3403 1596 3404 1600
rect 3398 1595 3404 1596
rect 3550 1600 3556 1601
rect 3550 1596 3551 1600
rect 3555 1596 3556 1600
rect 3550 1595 3556 1596
rect 3354 1579 3360 1580
rect 3354 1575 3355 1579
rect 3359 1575 3360 1579
rect 3354 1574 3360 1575
rect 3400 1567 3402 1595
rect 3450 1575 3456 1576
rect 3450 1571 3451 1575
rect 3455 1571 3456 1575
rect 3450 1570 3456 1571
rect 2743 1566 2747 1567
rect 2743 1561 2747 1562
rect 2839 1566 2843 1567
rect 2839 1561 2843 1562
rect 2903 1566 2907 1567
rect 2903 1561 2907 1562
rect 3047 1566 3051 1567
rect 3047 1561 3051 1562
rect 3063 1566 3067 1567
rect 3063 1561 3067 1562
rect 3223 1566 3227 1567
rect 3223 1561 3227 1562
rect 3231 1566 3235 1567
rect 3231 1561 3235 1562
rect 3383 1566 3387 1567
rect 3383 1561 3387 1562
rect 3399 1566 3403 1567
rect 3399 1561 3403 1562
rect 2674 1559 2680 1560
rect 2674 1555 2675 1559
rect 2679 1555 2680 1559
rect 2674 1554 2680 1555
rect 2710 1559 2716 1560
rect 2710 1555 2711 1559
rect 2715 1555 2716 1559
rect 2710 1554 2716 1555
rect 2582 1536 2588 1537
rect 2046 1533 2052 1534
rect 2046 1529 2047 1533
rect 2051 1529 2052 1533
rect 2582 1532 2583 1536
rect 2587 1532 2588 1536
rect 2582 1531 2588 1532
rect 2046 1528 2052 1529
rect 2712 1528 2714 1554
rect 2744 1537 2746 1561
rect 2818 1559 2824 1560
rect 2818 1555 2819 1559
rect 2823 1555 2824 1559
rect 2818 1554 2824 1555
rect 2742 1536 2748 1537
rect 2742 1532 2743 1536
rect 2747 1532 2748 1536
rect 2742 1531 2748 1532
rect 2820 1528 2822 1554
rect 2904 1537 2906 1561
rect 2978 1559 2984 1560
rect 2978 1555 2979 1559
rect 2983 1555 2984 1559
rect 2978 1554 2984 1555
rect 2902 1536 2908 1537
rect 2902 1532 2903 1536
rect 2907 1532 2908 1536
rect 2902 1531 2908 1532
rect 2980 1528 2982 1554
rect 3064 1537 3066 1561
rect 3224 1537 3226 1561
rect 3298 1559 3304 1560
rect 3298 1555 3299 1559
rect 3303 1555 3304 1559
rect 3298 1554 3304 1555
rect 3062 1536 3068 1537
rect 3062 1532 3063 1536
rect 3067 1532 3068 1536
rect 3062 1531 3068 1532
rect 3222 1536 3228 1537
rect 3222 1532 3223 1536
rect 3227 1532 3228 1536
rect 3222 1531 3228 1532
rect 3300 1528 3302 1554
rect 3384 1537 3386 1561
rect 3382 1536 3388 1537
rect 3382 1532 3383 1536
rect 3387 1532 3388 1536
rect 3382 1531 3388 1532
rect 3452 1528 3454 1570
rect 3552 1567 3554 1595
rect 3616 1580 3618 1678
rect 3646 1673 3652 1674
rect 3646 1669 3647 1673
rect 3651 1669 3652 1673
rect 3646 1668 3652 1669
rect 3838 1673 3844 1674
rect 3838 1669 3839 1673
rect 3843 1669 3844 1673
rect 3838 1668 3844 1669
rect 3648 1647 3650 1668
rect 3840 1647 3842 1668
rect 3647 1646 3651 1647
rect 3647 1641 3651 1642
rect 3695 1646 3699 1647
rect 3695 1641 3699 1642
rect 3839 1646 3843 1647
rect 3839 1641 3843 1642
rect 3696 1620 3698 1641
rect 3840 1620 3842 1641
rect 3694 1619 3700 1620
rect 3694 1615 3695 1619
rect 3699 1615 3700 1619
rect 3694 1614 3700 1615
rect 3838 1619 3844 1620
rect 3838 1615 3839 1619
rect 3843 1615 3844 1619
rect 3838 1614 3844 1615
rect 3916 1612 3918 1710
rect 3944 1690 3946 1717
rect 3942 1689 3948 1690
rect 3942 1685 3943 1689
rect 3947 1685 3948 1689
rect 3942 1684 3948 1685
rect 3942 1672 3948 1673
rect 3942 1668 3943 1672
rect 3947 1668 3948 1672
rect 3942 1667 3948 1668
rect 3944 1647 3946 1667
rect 3943 1646 3947 1647
rect 3943 1641 3947 1642
rect 3944 1621 3946 1641
rect 3942 1620 3948 1621
rect 3942 1616 3943 1620
rect 3947 1616 3948 1620
rect 3942 1615 3948 1616
rect 3914 1611 3920 1612
rect 3626 1607 3632 1608
rect 3626 1603 3627 1607
rect 3631 1603 3632 1607
rect 3626 1602 3632 1603
rect 3770 1607 3776 1608
rect 3770 1603 3771 1607
rect 3775 1603 3776 1607
rect 3914 1607 3915 1611
rect 3919 1607 3920 1611
rect 3914 1606 3920 1607
rect 3770 1602 3776 1603
rect 3942 1603 3948 1604
rect 3628 1580 3630 1602
rect 3694 1600 3700 1601
rect 3694 1596 3695 1600
rect 3699 1596 3700 1600
rect 3694 1595 3700 1596
rect 3614 1579 3620 1580
rect 3614 1575 3615 1579
rect 3619 1575 3620 1579
rect 3614 1574 3620 1575
rect 3626 1579 3632 1580
rect 3626 1575 3627 1579
rect 3631 1575 3632 1579
rect 3626 1574 3632 1575
rect 3696 1567 3698 1595
rect 3543 1566 3547 1567
rect 3543 1561 3547 1562
rect 3551 1566 3555 1567
rect 3551 1561 3555 1562
rect 3695 1566 3699 1567
rect 3695 1561 3699 1562
rect 3703 1566 3707 1567
rect 3703 1561 3707 1562
rect 3498 1551 3504 1552
rect 3498 1547 3499 1551
rect 3503 1547 3504 1551
rect 3498 1546 3504 1547
rect 3500 1528 3502 1546
rect 3544 1537 3546 1561
rect 3638 1559 3644 1560
rect 3638 1555 3639 1559
rect 3643 1555 3644 1559
rect 3638 1554 3644 1555
rect 3542 1536 3548 1537
rect 3542 1532 3543 1536
rect 3547 1532 3548 1536
rect 3542 1531 3548 1532
rect 3640 1528 3642 1554
rect 3704 1537 3706 1561
rect 3772 1560 3774 1602
rect 3838 1600 3844 1601
rect 3838 1596 3839 1600
rect 3843 1596 3844 1600
rect 3942 1599 3943 1603
rect 3947 1599 3948 1603
rect 3942 1598 3948 1599
rect 3838 1595 3844 1596
rect 3840 1567 3842 1595
rect 3890 1575 3896 1576
rect 3890 1571 3891 1575
rect 3895 1571 3896 1575
rect 3890 1570 3896 1571
rect 3839 1566 3843 1567
rect 3839 1561 3843 1562
rect 3770 1559 3776 1560
rect 3770 1555 3771 1559
rect 3775 1555 3776 1559
rect 3770 1554 3776 1555
rect 3702 1536 3708 1537
rect 3702 1532 3703 1536
rect 3707 1532 3708 1536
rect 3702 1531 3708 1532
rect 2710 1527 2716 1528
rect 2710 1523 2711 1527
rect 2715 1523 2716 1527
rect 2710 1522 2716 1523
rect 2818 1527 2824 1528
rect 2818 1523 2819 1527
rect 2823 1523 2824 1527
rect 2818 1522 2824 1523
rect 2978 1527 2984 1528
rect 2978 1523 2979 1527
rect 2983 1523 2984 1527
rect 2978 1522 2984 1523
rect 3018 1527 3024 1528
rect 3018 1523 3019 1527
rect 3023 1523 3024 1527
rect 3018 1522 3024 1523
rect 3298 1527 3304 1528
rect 3298 1523 3299 1527
rect 3303 1523 3304 1527
rect 3298 1522 3304 1523
rect 3450 1527 3456 1528
rect 3450 1523 3451 1527
rect 3455 1523 3456 1527
rect 3450 1522 3456 1523
rect 3498 1527 3504 1528
rect 3498 1523 3499 1527
rect 3503 1523 3504 1527
rect 3498 1522 3504 1523
rect 3638 1527 3644 1528
rect 3638 1523 3639 1527
rect 3643 1523 3644 1527
rect 3638 1522 3644 1523
rect 2006 1517 2012 1518
rect 2582 1517 2588 1518
rect 2006 1513 2007 1517
rect 2011 1513 2012 1517
rect 2006 1512 2012 1513
rect 2046 1516 2052 1517
rect 2046 1512 2047 1516
rect 2051 1512 2052 1516
rect 2582 1513 2583 1517
rect 2587 1513 2588 1517
rect 2582 1512 2588 1513
rect 2742 1517 2748 1518
rect 2742 1513 2743 1517
rect 2747 1513 2748 1517
rect 2742 1512 2748 1513
rect 2902 1517 2908 1518
rect 2902 1513 2903 1517
rect 2907 1513 2908 1517
rect 2902 1512 2908 1513
rect 2046 1511 2052 1512
rect 2006 1500 2012 1501
rect 2006 1496 2007 1500
rect 2011 1496 2012 1500
rect 2006 1495 2012 1496
rect 2008 1475 2010 1495
rect 2048 1491 2050 1511
rect 2584 1491 2586 1512
rect 2744 1491 2746 1512
rect 2904 1491 2906 1512
rect 2047 1490 2051 1491
rect 2047 1485 2051 1486
rect 2415 1490 2419 1491
rect 2415 1485 2419 1486
rect 2511 1490 2515 1491
rect 2511 1485 2515 1486
rect 2583 1490 2587 1491
rect 2583 1485 2587 1486
rect 2607 1490 2611 1491
rect 2607 1485 2611 1486
rect 2703 1490 2707 1491
rect 2703 1485 2707 1486
rect 2743 1490 2747 1491
rect 2743 1485 2747 1486
rect 2799 1490 2803 1491
rect 2799 1485 2803 1486
rect 2903 1490 2907 1491
rect 2903 1485 2907 1486
rect 2919 1490 2923 1491
rect 2919 1485 2923 1486
rect 1903 1474 1907 1475
rect 1903 1469 1907 1470
rect 2007 1474 2011 1475
rect 2007 1469 2011 1470
rect 1904 1448 1906 1469
rect 2008 1449 2010 1469
rect 2048 1465 2050 1485
rect 2046 1464 2052 1465
rect 2416 1464 2418 1485
rect 2512 1464 2514 1485
rect 2608 1464 2610 1485
rect 2704 1464 2706 1485
rect 2800 1464 2802 1485
rect 2920 1464 2922 1485
rect 2046 1460 2047 1464
rect 2051 1460 2052 1464
rect 2046 1459 2052 1460
rect 2414 1463 2420 1464
rect 2414 1459 2415 1463
rect 2419 1459 2420 1463
rect 2414 1458 2420 1459
rect 2510 1463 2516 1464
rect 2510 1459 2511 1463
rect 2515 1459 2516 1463
rect 2510 1458 2516 1459
rect 2606 1463 2612 1464
rect 2606 1459 2607 1463
rect 2611 1459 2612 1463
rect 2606 1458 2612 1459
rect 2702 1463 2708 1464
rect 2702 1459 2703 1463
rect 2707 1459 2708 1463
rect 2702 1458 2708 1459
rect 2798 1463 2804 1464
rect 2798 1459 2799 1463
rect 2803 1459 2804 1463
rect 2798 1458 2804 1459
rect 2918 1463 2924 1464
rect 2918 1459 2919 1463
rect 2923 1459 2924 1463
rect 2918 1458 2924 1459
rect 2490 1451 2496 1452
rect 2006 1448 2012 1449
rect 1902 1447 1908 1448
rect 1902 1443 1903 1447
rect 1907 1443 1908 1447
rect 2006 1444 2007 1448
rect 2011 1444 2012 1448
rect 2006 1443 2012 1444
rect 2046 1447 2052 1448
rect 2046 1443 2047 1447
rect 2051 1443 2052 1447
rect 2490 1447 2491 1451
rect 2495 1447 2496 1451
rect 2490 1446 2496 1447
rect 2586 1451 2592 1452
rect 2586 1447 2587 1451
rect 2591 1447 2592 1451
rect 2586 1446 2592 1447
rect 2682 1451 2688 1452
rect 2682 1447 2683 1451
rect 2687 1447 2688 1451
rect 2682 1446 2688 1447
rect 2778 1451 2784 1452
rect 2778 1447 2779 1451
rect 2783 1447 2784 1451
rect 2778 1446 2784 1447
rect 2874 1451 2880 1452
rect 2874 1447 2875 1451
rect 2879 1447 2880 1451
rect 2874 1446 2880 1447
rect 2994 1451 3000 1452
rect 2994 1447 2995 1451
rect 2999 1447 3000 1451
rect 2994 1446 3000 1447
rect 1902 1442 1908 1443
rect 2046 1442 2052 1443
rect 2414 1444 2420 1445
rect 1862 1439 1868 1440
rect 1082 1435 1088 1436
rect 1082 1431 1083 1435
rect 1087 1431 1088 1435
rect 1082 1430 1088 1431
rect 1538 1435 1544 1436
rect 1538 1431 1539 1435
rect 1543 1431 1544 1435
rect 1538 1430 1544 1431
rect 1770 1435 1776 1436
rect 1770 1431 1771 1435
rect 1775 1431 1776 1435
rect 1862 1435 1863 1439
rect 1867 1435 1868 1439
rect 1862 1434 1868 1435
rect 1770 1430 1776 1431
rect 2006 1431 2012 1432
rect 1006 1428 1012 1429
rect 1006 1424 1007 1428
rect 1011 1424 1012 1428
rect 1006 1423 1012 1424
rect 838 1407 844 1408
rect 838 1403 839 1407
rect 843 1403 844 1407
rect 838 1402 844 1403
rect 930 1403 936 1404
rect 930 1399 931 1403
rect 935 1399 936 1403
rect 1008 1399 1010 1423
rect 1084 1408 1086 1430
rect 1230 1428 1236 1429
rect 1230 1424 1231 1428
rect 1235 1424 1236 1428
rect 1230 1423 1236 1424
rect 1462 1428 1468 1429
rect 1462 1424 1463 1428
rect 1467 1424 1468 1428
rect 1462 1423 1468 1424
rect 1082 1407 1088 1408
rect 1082 1403 1083 1407
rect 1087 1403 1088 1407
rect 1082 1402 1088 1403
rect 1232 1399 1234 1423
rect 1464 1399 1466 1423
rect 1540 1408 1542 1430
rect 1694 1428 1700 1429
rect 1694 1424 1695 1428
rect 1699 1424 1700 1428
rect 1694 1423 1700 1424
rect 1538 1407 1544 1408
rect 1538 1403 1539 1407
rect 1543 1403 1544 1407
rect 1538 1402 1544 1403
rect 1666 1399 1672 1400
rect 1696 1399 1698 1423
rect 1772 1408 1774 1430
rect 1902 1428 1908 1429
rect 1902 1424 1903 1428
rect 1907 1424 1908 1428
rect 2006 1427 2007 1431
rect 2011 1427 2012 1431
rect 2006 1426 2012 1427
rect 1902 1423 1908 1424
rect 1770 1407 1776 1408
rect 1770 1403 1771 1407
rect 1775 1403 1776 1407
rect 1770 1402 1776 1403
rect 1904 1399 1906 1423
rect 2008 1399 2010 1426
rect 463 1398 467 1399
rect 463 1393 467 1394
rect 567 1398 571 1399
rect 567 1393 571 1394
rect 599 1398 603 1399
rect 599 1393 603 1394
rect 727 1398 731 1399
rect 727 1393 731 1394
rect 783 1398 787 1399
rect 783 1393 787 1394
rect 855 1398 859 1399
rect 930 1398 936 1399
rect 983 1398 987 1399
rect 855 1393 859 1394
rect 442 1391 448 1392
rect 442 1387 443 1391
rect 447 1387 448 1391
rect 442 1386 448 1387
rect 464 1369 466 1393
rect 518 1391 524 1392
rect 518 1386 519 1391
rect 523 1386 524 1391
rect 538 1391 544 1392
rect 538 1387 539 1391
rect 543 1387 544 1391
rect 538 1386 544 1387
rect 519 1383 523 1384
rect 462 1368 468 1369
rect 462 1364 463 1368
rect 467 1364 468 1368
rect 462 1363 468 1364
rect 540 1360 542 1386
rect 600 1369 602 1393
rect 674 1391 680 1392
rect 674 1387 675 1391
rect 679 1387 680 1391
rect 674 1386 680 1387
rect 598 1368 604 1369
rect 598 1364 599 1368
rect 603 1364 604 1368
rect 598 1363 604 1364
rect 676 1360 678 1386
rect 728 1369 730 1393
rect 802 1391 808 1392
rect 802 1387 803 1391
rect 807 1387 808 1391
rect 802 1386 808 1387
rect 726 1368 732 1369
rect 726 1364 727 1368
rect 731 1364 732 1368
rect 726 1363 732 1364
rect 804 1360 806 1386
rect 856 1369 858 1393
rect 854 1368 860 1369
rect 854 1364 855 1368
rect 859 1364 860 1368
rect 854 1363 860 1364
rect 932 1360 934 1398
rect 983 1393 987 1394
rect 1007 1398 1011 1399
rect 1007 1393 1011 1394
rect 1119 1398 1123 1399
rect 1119 1393 1123 1394
rect 1231 1398 1235 1399
rect 1231 1393 1235 1394
rect 1263 1398 1267 1399
rect 1263 1393 1267 1394
rect 1423 1398 1427 1399
rect 1423 1393 1427 1394
rect 1463 1398 1467 1399
rect 1463 1393 1467 1394
rect 1583 1398 1587 1399
rect 1666 1395 1667 1399
rect 1671 1395 1672 1399
rect 1666 1394 1672 1395
rect 1695 1398 1699 1399
rect 1583 1393 1587 1394
rect 963 1388 967 1389
rect 963 1383 967 1384
rect 402 1359 408 1360
rect 402 1355 403 1359
rect 407 1355 408 1359
rect 402 1354 408 1355
rect 538 1359 544 1360
rect 538 1355 539 1359
rect 543 1355 544 1359
rect 538 1354 544 1355
rect 674 1359 680 1360
rect 674 1355 675 1359
rect 679 1355 680 1359
rect 674 1354 680 1355
rect 802 1359 808 1360
rect 802 1355 803 1359
rect 807 1355 808 1359
rect 802 1354 808 1355
rect 930 1359 936 1360
rect 930 1355 931 1359
rect 935 1355 936 1359
rect 930 1354 936 1355
rect 326 1349 332 1350
rect 110 1348 116 1349
rect 110 1344 111 1348
rect 115 1344 116 1348
rect 326 1345 327 1349
rect 331 1345 332 1349
rect 326 1344 332 1345
rect 462 1349 468 1350
rect 462 1345 463 1349
rect 467 1345 468 1349
rect 462 1344 468 1345
rect 598 1349 604 1350
rect 598 1345 599 1349
rect 603 1345 604 1349
rect 598 1344 604 1345
rect 726 1349 732 1350
rect 726 1345 727 1349
rect 731 1345 732 1349
rect 726 1344 732 1345
rect 854 1349 860 1350
rect 854 1345 855 1349
rect 859 1345 860 1349
rect 854 1344 860 1345
rect 110 1343 116 1344
rect 112 1315 114 1343
rect 328 1315 330 1344
rect 464 1315 466 1344
rect 600 1315 602 1344
rect 728 1315 730 1344
rect 856 1315 858 1344
rect 111 1314 115 1315
rect 111 1309 115 1310
rect 327 1314 331 1315
rect 327 1309 331 1310
rect 463 1314 467 1315
rect 463 1309 467 1310
rect 551 1314 555 1315
rect 551 1309 555 1310
rect 599 1314 603 1315
rect 599 1309 603 1310
rect 655 1314 659 1315
rect 655 1309 659 1310
rect 727 1314 731 1315
rect 727 1309 731 1310
rect 767 1314 771 1315
rect 767 1309 771 1310
rect 855 1314 859 1315
rect 855 1309 859 1310
rect 879 1314 883 1315
rect 879 1309 883 1310
rect 112 1289 114 1309
rect 110 1288 116 1289
rect 552 1288 554 1309
rect 656 1288 658 1309
rect 768 1288 770 1309
rect 880 1288 882 1309
rect 110 1284 111 1288
rect 115 1284 116 1288
rect 110 1283 116 1284
rect 550 1287 556 1288
rect 550 1283 551 1287
rect 555 1283 556 1287
rect 550 1282 556 1283
rect 654 1287 660 1288
rect 654 1283 655 1287
rect 659 1283 660 1287
rect 654 1282 660 1283
rect 766 1287 772 1288
rect 766 1283 767 1287
rect 771 1283 772 1287
rect 766 1282 772 1283
rect 878 1287 884 1288
rect 878 1283 879 1287
rect 883 1283 884 1287
rect 878 1282 884 1283
rect 964 1280 966 1383
rect 984 1369 986 1393
rect 1058 1391 1064 1392
rect 1058 1387 1059 1391
rect 1063 1387 1064 1391
rect 1058 1386 1064 1387
rect 982 1368 988 1369
rect 982 1364 983 1368
rect 987 1364 988 1368
rect 982 1363 988 1364
rect 1060 1360 1062 1386
rect 1120 1369 1122 1393
rect 1194 1391 1200 1392
rect 1194 1387 1195 1391
rect 1199 1387 1200 1391
rect 1194 1386 1200 1387
rect 1118 1368 1124 1369
rect 1118 1364 1119 1368
rect 1123 1364 1124 1368
rect 1118 1363 1124 1364
rect 1196 1360 1198 1386
rect 1264 1369 1266 1393
rect 1338 1391 1344 1392
rect 1338 1387 1339 1391
rect 1343 1387 1344 1391
rect 1338 1386 1344 1387
rect 1262 1368 1268 1369
rect 1262 1364 1263 1368
rect 1267 1364 1268 1368
rect 1262 1363 1268 1364
rect 1340 1360 1342 1386
rect 1402 1383 1408 1384
rect 1402 1379 1403 1383
rect 1407 1379 1408 1383
rect 1402 1378 1408 1379
rect 1058 1359 1064 1360
rect 1058 1355 1059 1359
rect 1063 1355 1064 1359
rect 1058 1354 1064 1355
rect 1194 1359 1200 1360
rect 1194 1355 1195 1359
rect 1199 1355 1200 1359
rect 1194 1354 1200 1355
rect 1338 1359 1344 1360
rect 1338 1355 1339 1359
rect 1343 1355 1344 1359
rect 1338 1354 1344 1355
rect 982 1349 988 1350
rect 982 1345 983 1349
rect 987 1345 988 1349
rect 982 1344 988 1345
rect 1118 1349 1124 1350
rect 1118 1345 1119 1349
rect 1123 1345 1124 1349
rect 1118 1344 1124 1345
rect 1262 1349 1268 1350
rect 1262 1345 1263 1349
rect 1267 1345 1268 1349
rect 1262 1344 1268 1345
rect 984 1315 986 1344
rect 1120 1315 1122 1344
rect 1178 1343 1184 1344
rect 1178 1339 1179 1343
rect 1183 1339 1184 1343
rect 1178 1338 1184 1339
rect 983 1314 987 1315
rect 983 1309 987 1310
rect 991 1314 995 1315
rect 991 1309 995 1310
rect 1103 1314 1107 1315
rect 1103 1309 1107 1310
rect 1119 1314 1123 1315
rect 1119 1309 1123 1310
rect 992 1288 994 1309
rect 1104 1288 1106 1309
rect 990 1287 996 1288
rect 990 1283 991 1287
rect 995 1283 996 1287
rect 990 1282 996 1283
rect 1102 1287 1108 1288
rect 1102 1283 1103 1287
rect 1107 1283 1108 1287
rect 1102 1282 1108 1283
rect 962 1279 968 1280
rect 626 1275 632 1276
rect 110 1271 116 1272
rect 110 1267 111 1271
rect 115 1267 116 1271
rect 626 1271 627 1275
rect 631 1271 632 1275
rect 626 1270 632 1271
rect 730 1275 736 1276
rect 730 1271 731 1275
rect 735 1271 736 1275
rect 730 1270 736 1271
rect 842 1275 848 1276
rect 842 1271 843 1275
rect 847 1271 848 1275
rect 842 1270 848 1271
rect 954 1275 960 1276
rect 954 1271 955 1275
rect 959 1271 960 1275
rect 962 1275 963 1279
rect 967 1275 968 1279
rect 962 1274 968 1275
rect 1086 1279 1092 1280
rect 1086 1275 1087 1279
rect 1091 1275 1092 1279
rect 1086 1274 1092 1275
rect 954 1270 960 1271
rect 110 1266 116 1267
rect 550 1268 556 1269
rect 112 1239 114 1266
rect 550 1264 551 1268
rect 555 1264 556 1268
rect 550 1263 556 1264
rect 552 1239 554 1263
rect 628 1248 630 1270
rect 654 1268 660 1269
rect 654 1264 655 1268
rect 659 1264 660 1268
rect 654 1263 660 1264
rect 626 1247 632 1248
rect 626 1243 627 1247
rect 631 1243 632 1247
rect 626 1242 632 1243
rect 656 1239 658 1263
rect 732 1248 734 1270
rect 766 1268 772 1269
rect 766 1264 767 1268
rect 771 1264 772 1268
rect 766 1263 772 1264
rect 730 1247 736 1248
rect 730 1243 731 1247
rect 735 1243 736 1247
rect 730 1242 736 1243
rect 768 1239 770 1263
rect 844 1248 846 1270
rect 878 1268 884 1269
rect 878 1264 879 1268
rect 883 1264 884 1268
rect 878 1263 884 1264
rect 842 1247 848 1248
rect 842 1243 843 1247
rect 847 1243 848 1247
rect 842 1242 848 1243
rect 880 1239 882 1263
rect 956 1248 958 1270
rect 990 1268 996 1269
rect 990 1264 991 1268
rect 995 1264 996 1268
rect 990 1263 996 1264
rect 954 1247 960 1248
rect 954 1243 955 1247
rect 959 1243 960 1247
rect 954 1242 960 1243
rect 938 1239 944 1240
rect 992 1239 994 1263
rect 111 1238 115 1239
rect 111 1233 115 1234
rect 391 1238 395 1239
rect 391 1233 395 1234
rect 519 1238 523 1239
rect 519 1233 523 1234
rect 551 1238 555 1239
rect 551 1233 555 1234
rect 655 1238 659 1239
rect 655 1233 659 1234
rect 663 1238 667 1239
rect 663 1233 667 1234
rect 767 1238 771 1239
rect 767 1233 771 1234
rect 807 1238 811 1239
rect 807 1233 811 1234
rect 879 1238 883 1239
rect 938 1235 939 1239
rect 943 1235 944 1239
rect 938 1234 944 1235
rect 959 1238 963 1239
rect 879 1233 883 1234
rect 112 1206 114 1233
rect 392 1209 394 1233
rect 466 1231 472 1232
rect 466 1227 467 1231
rect 471 1227 472 1231
rect 466 1226 472 1227
rect 390 1208 396 1209
rect 110 1205 116 1206
rect 110 1201 111 1205
rect 115 1201 116 1205
rect 390 1204 391 1208
rect 395 1204 396 1208
rect 390 1203 396 1204
rect 110 1200 116 1201
rect 468 1200 470 1226
rect 520 1209 522 1233
rect 594 1231 600 1232
rect 594 1227 595 1231
rect 599 1227 600 1231
rect 594 1226 600 1227
rect 518 1208 524 1209
rect 518 1204 519 1208
rect 523 1204 524 1208
rect 518 1203 524 1204
rect 596 1200 598 1226
rect 664 1209 666 1233
rect 738 1231 744 1232
rect 738 1227 739 1231
rect 743 1227 744 1231
rect 738 1226 744 1227
rect 662 1208 668 1209
rect 662 1204 663 1208
rect 667 1204 668 1208
rect 662 1203 668 1204
rect 740 1200 742 1226
rect 798 1223 804 1224
rect 798 1219 799 1223
rect 803 1219 804 1223
rect 798 1218 804 1219
rect 466 1199 472 1200
rect 466 1195 467 1199
rect 471 1195 472 1199
rect 466 1194 472 1195
rect 594 1199 600 1200
rect 594 1195 595 1199
rect 599 1195 600 1199
rect 594 1194 600 1195
rect 738 1199 744 1200
rect 738 1195 739 1199
rect 743 1195 744 1199
rect 738 1194 744 1195
rect 390 1189 396 1190
rect 110 1188 116 1189
rect 110 1184 111 1188
rect 115 1184 116 1188
rect 390 1185 391 1189
rect 395 1185 396 1189
rect 390 1184 396 1185
rect 518 1189 524 1190
rect 518 1185 519 1189
rect 523 1185 524 1189
rect 518 1184 524 1185
rect 662 1189 668 1190
rect 662 1185 663 1189
rect 667 1185 668 1189
rect 662 1184 668 1185
rect 110 1183 116 1184
rect 112 1159 114 1183
rect 392 1159 394 1184
rect 520 1159 522 1184
rect 664 1159 666 1184
rect 111 1158 115 1159
rect 111 1153 115 1154
rect 175 1158 179 1159
rect 175 1153 179 1154
rect 327 1158 331 1159
rect 327 1153 331 1154
rect 391 1158 395 1159
rect 391 1153 395 1154
rect 495 1158 499 1159
rect 495 1153 499 1154
rect 519 1158 523 1159
rect 519 1153 523 1154
rect 663 1158 667 1159
rect 663 1153 667 1154
rect 671 1158 675 1159
rect 671 1153 675 1154
rect 112 1133 114 1153
rect 110 1132 116 1133
rect 176 1132 178 1153
rect 328 1132 330 1153
rect 496 1132 498 1153
rect 672 1132 674 1153
rect 110 1128 111 1132
rect 115 1128 116 1132
rect 110 1127 116 1128
rect 174 1131 180 1132
rect 174 1127 175 1131
rect 179 1127 180 1131
rect 174 1126 180 1127
rect 326 1131 332 1132
rect 326 1127 327 1131
rect 331 1127 332 1131
rect 326 1126 332 1127
rect 494 1131 500 1132
rect 494 1127 495 1131
rect 499 1127 500 1131
rect 494 1126 500 1127
rect 670 1131 676 1132
rect 670 1127 671 1131
rect 675 1127 676 1131
rect 670 1126 676 1127
rect 800 1124 802 1218
rect 808 1209 810 1233
rect 806 1208 812 1209
rect 806 1204 807 1208
rect 811 1204 812 1208
rect 806 1203 812 1204
rect 940 1200 942 1234
rect 959 1233 963 1234
rect 991 1238 995 1239
rect 991 1233 995 1234
rect 960 1209 962 1233
rect 958 1208 964 1209
rect 958 1204 959 1208
rect 963 1204 964 1208
rect 958 1203 964 1204
rect 938 1199 944 1200
rect 938 1195 939 1199
rect 943 1195 944 1199
rect 938 1194 944 1195
rect 806 1189 812 1190
rect 806 1185 807 1189
rect 811 1185 812 1189
rect 806 1184 812 1185
rect 958 1189 964 1190
rect 958 1185 959 1189
rect 963 1185 964 1189
rect 958 1184 964 1185
rect 808 1159 810 1184
rect 960 1159 962 1184
rect 807 1158 811 1159
rect 807 1153 811 1154
rect 847 1158 851 1159
rect 847 1153 851 1154
rect 959 1158 963 1159
rect 959 1153 963 1154
rect 1031 1158 1035 1159
rect 1031 1153 1035 1154
rect 848 1132 850 1153
rect 1032 1132 1034 1153
rect 846 1131 852 1132
rect 846 1127 847 1131
rect 851 1127 852 1131
rect 846 1126 852 1127
rect 1030 1131 1036 1132
rect 1030 1127 1031 1131
rect 1035 1127 1036 1131
rect 1030 1126 1036 1127
rect 798 1123 804 1124
rect 250 1119 256 1120
rect 110 1115 116 1116
rect 110 1111 111 1115
rect 115 1111 116 1115
rect 250 1115 251 1119
rect 255 1115 256 1119
rect 250 1114 256 1115
rect 402 1119 408 1120
rect 402 1115 403 1119
rect 407 1115 408 1119
rect 402 1114 408 1115
rect 570 1119 576 1120
rect 570 1115 571 1119
rect 575 1115 576 1119
rect 570 1114 576 1115
rect 746 1119 752 1120
rect 746 1115 747 1119
rect 751 1115 752 1119
rect 798 1119 799 1123
rect 803 1119 804 1123
rect 798 1118 804 1119
rect 746 1114 752 1115
rect 110 1110 116 1111
rect 174 1112 180 1113
rect 112 1075 114 1110
rect 174 1108 175 1112
rect 179 1108 180 1112
rect 174 1107 180 1108
rect 176 1075 178 1107
rect 252 1092 254 1114
rect 326 1112 332 1113
rect 326 1108 327 1112
rect 331 1108 332 1112
rect 326 1107 332 1108
rect 250 1091 256 1092
rect 242 1087 248 1088
rect 242 1083 243 1087
rect 247 1083 248 1087
rect 250 1087 251 1091
rect 255 1087 256 1091
rect 250 1086 256 1087
rect 242 1082 248 1083
rect 111 1074 115 1075
rect 111 1069 115 1070
rect 135 1074 139 1075
rect 135 1069 139 1070
rect 175 1074 179 1075
rect 175 1069 179 1070
rect 231 1074 235 1075
rect 231 1069 235 1070
rect 112 1042 114 1069
rect 136 1045 138 1069
rect 202 1067 208 1068
rect 202 1063 203 1067
rect 207 1063 208 1067
rect 202 1062 208 1063
rect 210 1067 216 1068
rect 210 1063 211 1067
rect 215 1063 216 1067
rect 210 1062 216 1063
rect 134 1044 140 1045
rect 110 1041 116 1042
rect 110 1037 111 1041
rect 115 1037 116 1041
rect 134 1040 135 1044
rect 139 1040 140 1044
rect 134 1039 140 1040
rect 110 1036 116 1037
rect 134 1025 140 1026
rect 110 1024 116 1025
rect 110 1020 111 1024
rect 115 1020 116 1024
rect 134 1021 135 1025
rect 139 1021 140 1025
rect 134 1020 140 1021
rect 110 1019 116 1020
rect 112 999 114 1019
rect 136 999 138 1020
rect 111 998 115 999
rect 111 993 115 994
rect 135 998 139 999
rect 135 993 139 994
rect 112 973 114 993
rect 110 972 116 973
rect 136 972 138 993
rect 110 968 111 972
rect 115 968 116 972
rect 110 967 116 968
rect 134 971 140 972
rect 134 967 135 971
rect 139 967 140 971
rect 204 968 206 1062
rect 212 1036 214 1062
rect 232 1045 234 1069
rect 244 1061 246 1082
rect 328 1075 330 1107
rect 404 1092 406 1114
rect 494 1112 500 1113
rect 494 1108 495 1112
rect 499 1108 500 1112
rect 494 1107 500 1108
rect 402 1091 408 1092
rect 402 1087 403 1091
rect 407 1087 408 1091
rect 402 1086 408 1087
rect 496 1075 498 1107
rect 572 1092 574 1114
rect 670 1112 676 1113
rect 670 1108 671 1112
rect 675 1108 676 1112
rect 670 1107 676 1108
rect 570 1091 576 1092
rect 570 1087 571 1091
rect 575 1087 576 1091
rect 570 1086 576 1087
rect 672 1075 674 1107
rect 748 1092 750 1114
rect 846 1112 852 1113
rect 846 1108 847 1112
rect 851 1108 852 1112
rect 846 1107 852 1108
rect 1030 1112 1036 1113
rect 1030 1108 1031 1112
rect 1035 1108 1036 1112
rect 1030 1107 1036 1108
rect 746 1091 752 1092
rect 746 1087 747 1091
rect 751 1087 752 1091
rect 746 1086 752 1087
rect 848 1075 850 1107
rect 1032 1075 1034 1107
rect 1088 1092 1090 1274
rect 1102 1268 1108 1269
rect 1102 1264 1103 1268
rect 1107 1264 1108 1268
rect 1102 1263 1108 1264
rect 1104 1239 1106 1263
rect 1180 1248 1182 1338
rect 1264 1315 1266 1344
rect 1215 1314 1219 1315
rect 1215 1309 1219 1310
rect 1263 1314 1267 1315
rect 1263 1309 1267 1310
rect 1327 1314 1331 1315
rect 1327 1309 1331 1310
rect 1216 1288 1218 1309
rect 1328 1288 1330 1309
rect 1214 1287 1220 1288
rect 1214 1283 1215 1287
rect 1219 1283 1220 1287
rect 1214 1282 1220 1283
rect 1326 1287 1332 1288
rect 1326 1283 1327 1287
rect 1331 1283 1332 1287
rect 1326 1282 1332 1283
rect 1404 1280 1406 1378
rect 1424 1369 1426 1393
rect 1584 1369 1586 1393
rect 1422 1368 1428 1369
rect 1422 1364 1423 1368
rect 1427 1364 1428 1368
rect 1422 1363 1428 1364
rect 1582 1368 1588 1369
rect 1582 1364 1583 1368
rect 1587 1364 1588 1368
rect 1582 1363 1588 1364
rect 1668 1360 1670 1394
rect 1695 1393 1699 1394
rect 1751 1398 1755 1399
rect 1751 1393 1755 1394
rect 1903 1398 1907 1399
rect 1903 1393 1907 1394
rect 2007 1398 2011 1399
rect 2048 1395 2050 1442
rect 2414 1440 2415 1444
rect 2419 1440 2420 1444
rect 2414 1439 2420 1440
rect 2416 1395 2418 1439
rect 2492 1424 2494 1446
rect 2510 1444 2516 1445
rect 2510 1440 2511 1444
rect 2515 1440 2516 1444
rect 2510 1439 2516 1440
rect 2490 1423 2496 1424
rect 2490 1419 2491 1423
rect 2495 1419 2496 1423
rect 2490 1418 2496 1419
rect 2512 1395 2514 1439
rect 2588 1424 2590 1446
rect 2606 1444 2612 1445
rect 2606 1440 2607 1444
rect 2611 1440 2612 1444
rect 2606 1439 2612 1440
rect 2586 1423 2592 1424
rect 2586 1419 2587 1423
rect 2591 1419 2592 1423
rect 2586 1418 2592 1419
rect 2608 1395 2610 1439
rect 2626 1435 2632 1436
rect 2626 1431 2627 1435
rect 2631 1431 2632 1435
rect 2626 1430 2632 1431
rect 2007 1393 2011 1394
rect 2047 1394 2051 1395
rect 1752 1369 1754 1393
rect 1834 1391 1840 1392
rect 1834 1387 1835 1391
rect 1839 1387 1840 1391
rect 1834 1386 1840 1387
rect 1750 1368 1756 1369
rect 1750 1364 1751 1368
rect 1755 1364 1756 1368
rect 1750 1363 1756 1364
rect 1836 1360 1838 1386
rect 1904 1369 1906 1393
rect 1986 1391 1992 1392
rect 1986 1387 1987 1391
rect 1991 1387 1992 1391
rect 1986 1386 1992 1387
rect 1902 1368 1908 1369
rect 1902 1364 1903 1368
rect 1907 1364 1908 1368
rect 1902 1363 1908 1364
rect 1650 1359 1656 1360
rect 1650 1355 1651 1359
rect 1655 1355 1656 1359
rect 1650 1354 1656 1355
rect 1666 1359 1672 1360
rect 1666 1355 1667 1359
rect 1671 1355 1672 1359
rect 1666 1354 1672 1355
rect 1834 1359 1840 1360
rect 1834 1355 1835 1359
rect 1839 1355 1840 1359
rect 1988 1356 1990 1386
rect 2008 1366 2010 1393
rect 2047 1389 2051 1390
rect 2071 1394 2075 1395
rect 2071 1389 2075 1390
rect 2303 1394 2307 1395
rect 2303 1389 2307 1390
rect 2415 1394 2419 1395
rect 2415 1389 2419 1390
rect 2511 1394 2515 1395
rect 2511 1389 2515 1390
rect 2559 1394 2563 1395
rect 2559 1389 2563 1390
rect 2607 1394 2611 1395
rect 2607 1389 2611 1390
rect 2006 1365 2012 1366
rect 2006 1361 2007 1365
rect 2011 1361 2012 1365
rect 2048 1362 2050 1389
rect 2072 1365 2074 1389
rect 2154 1387 2160 1388
rect 2154 1383 2155 1387
rect 2159 1383 2160 1387
rect 2154 1382 2160 1383
rect 2070 1364 2076 1365
rect 2006 1360 2012 1361
rect 2046 1361 2052 1362
rect 2046 1357 2047 1361
rect 2051 1357 2052 1361
rect 2070 1360 2071 1364
rect 2075 1360 2076 1364
rect 2070 1359 2076 1360
rect 2046 1356 2052 1357
rect 2156 1356 2158 1382
rect 2304 1365 2306 1389
rect 2310 1387 2316 1388
rect 2310 1383 2311 1387
rect 2315 1383 2316 1387
rect 2310 1382 2316 1383
rect 2302 1364 2308 1365
rect 2302 1360 2303 1364
rect 2307 1360 2308 1364
rect 2302 1359 2308 1360
rect 1834 1354 1840 1355
rect 1986 1355 1992 1356
rect 1422 1349 1428 1350
rect 1422 1345 1423 1349
rect 1427 1345 1428 1349
rect 1422 1344 1428 1345
rect 1582 1349 1588 1350
rect 1582 1345 1583 1349
rect 1587 1345 1588 1349
rect 1582 1344 1588 1345
rect 1424 1315 1426 1344
rect 1584 1315 1586 1344
rect 1423 1314 1427 1315
rect 1423 1309 1427 1310
rect 1439 1314 1443 1315
rect 1439 1309 1443 1310
rect 1559 1314 1563 1315
rect 1559 1309 1563 1310
rect 1583 1314 1587 1315
rect 1583 1309 1587 1310
rect 1440 1288 1442 1309
rect 1560 1288 1562 1309
rect 1438 1287 1444 1288
rect 1438 1283 1439 1287
rect 1443 1283 1444 1287
rect 1438 1282 1444 1283
rect 1558 1287 1564 1288
rect 1558 1283 1559 1287
rect 1563 1283 1564 1287
rect 1558 1282 1564 1283
rect 1402 1279 1408 1280
rect 1290 1275 1296 1276
rect 1290 1271 1291 1275
rect 1295 1271 1296 1275
rect 1402 1275 1403 1279
rect 1407 1275 1408 1279
rect 1526 1279 1532 1280
rect 1402 1274 1408 1275
rect 1514 1275 1520 1276
rect 1290 1270 1296 1271
rect 1514 1271 1515 1275
rect 1519 1271 1520 1275
rect 1526 1275 1527 1279
rect 1531 1275 1532 1279
rect 1526 1274 1532 1275
rect 1514 1270 1520 1271
rect 1214 1268 1220 1269
rect 1214 1264 1215 1268
rect 1219 1264 1220 1268
rect 1214 1263 1220 1264
rect 1178 1247 1184 1248
rect 1178 1243 1179 1247
rect 1183 1243 1184 1247
rect 1178 1242 1184 1243
rect 1186 1243 1192 1244
rect 1186 1239 1187 1243
rect 1191 1239 1192 1243
rect 1216 1239 1218 1263
rect 1292 1248 1294 1270
rect 1326 1268 1332 1269
rect 1326 1264 1327 1268
rect 1331 1264 1332 1268
rect 1326 1263 1332 1264
rect 1438 1268 1444 1269
rect 1438 1264 1439 1268
rect 1443 1264 1444 1268
rect 1438 1263 1444 1264
rect 1290 1247 1296 1248
rect 1290 1243 1291 1247
rect 1295 1243 1296 1247
rect 1290 1242 1296 1243
rect 1328 1239 1330 1263
rect 1440 1239 1442 1263
rect 1103 1238 1107 1239
rect 1103 1233 1107 1234
rect 1111 1238 1115 1239
rect 1186 1238 1192 1239
rect 1215 1238 1219 1239
rect 1111 1233 1115 1234
rect 1112 1209 1114 1233
rect 1110 1208 1116 1209
rect 1110 1204 1111 1208
rect 1115 1204 1116 1208
rect 1110 1203 1116 1204
rect 1188 1200 1190 1238
rect 1215 1233 1219 1234
rect 1255 1238 1259 1239
rect 1255 1233 1259 1234
rect 1327 1238 1331 1239
rect 1327 1233 1331 1234
rect 1407 1238 1411 1239
rect 1407 1233 1411 1234
rect 1439 1238 1443 1239
rect 1439 1233 1443 1234
rect 1194 1231 1200 1232
rect 1194 1227 1195 1231
rect 1199 1227 1200 1231
rect 1194 1226 1200 1227
rect 1196 1200 1198 1226
rect 1256 1209 1258 1233
rect 1282 1231 1288 1232
rect 1282 1227 1283 1231
rect 1287 1227 1288 1231
rect 1282 1226 1288 1227
rect 1254 1208 1260 1209
rect 1254 1204 1255 1208
rect 1259 1204 1260 1208
rect 1254 1203 1260 1204
rect 1186 1199 1192 1200
rect 1186 1195 1187 1199
rect 1191 1195 1192 1199
rect 1186 1194 1192 1195
rect 1194 1199 1200 1200
rect 1194 1195 1195 1199
rect 1199 1195 1200 1199
rect 1194 1194 1200 1195
rect 1110 1189 1116 1190
rect 1110 1185 1111 1189
rect 1115 1185 1116 1189
rect 1110 1184 1116 1185
rect 1254 1189 1260 1190
rect 1254 1185 1255 1189
rect 1259 1185 1260 1189
rect 1254 1184 1260 1185
rect 1112 1159 1114 1184
rect 1256 1159 1258 1184
rect 1111 1158 1115 1159
rect 1111 1153 1115 1154
rect 1207 1158 1211 1159
rect 1207 1153 1211 1154
rect 1255 1158 1259 1159
rect 1255 1153 1259 1154
rect 1208 1132 1210 1153
rect 1206 1131 1212 1132
rect 1206 1127 1207 1131
rect 1211 1127 1212 1131
rect 1206 1126 1212 1127
rect 1284 1124 1286 1226
rect 1408 1209 1410 1233
rect 1516 1232 1518 1270
rect 1528 1248 1530 1274
rect 1558 1268 1564 1269
rect 1558 1264 1559 1268
rect 1563 1264 1564 1268
rect 1558 1263 1564 1264
rect 1526 1247 1532 1248
rect 1526 1243 1527 1247
rect 1531 1243 1532 1247
rect 1526 1242 1532 1243
rect 1560 1239 1562 1263
rect 1652 1248 1654 1354
rect 1986 1351 1987 1355
rect 1991 1351 1992 1355
rect 1986 1350 1992 1351
rect 2154 1355 2160 1356
rect 2154 1351 2155 1355
rect 2159 1351 2160 1355
rect 2154 1350 2160 1351
rect 1750 1349 1756 1350
rect 1750 1345 1751 1349
rect 1755 1345 1756 1349
rect 1750 1344 1756 1345
rect 1902 1349 1908 1350
rect 1902 1345 1903 1349
rect 1907 1345 1908 1349
rect 1902 1344 1908 1345
rect 2006 1348 2012 1349
rect 2006 1344 2007 1348
rect 2011 1344 2012 1348
rect 2070 1345 2076 1346
rect 1752 1315 1754 1344
rect 1904 1315 1906 1344
rect 2006 1343 2012 1344
rect 2046 1344 2052 1345
rect 2008 1315 2010 1343
rect 2046 1340 2047 1344
rect 2051 1340 2052 1344
rect 2070 1341 2071 1345
rect 2075 1341 2076 1345
rect 2070 1340 2076 1341
rect 2302 1345 2308 1346
rect 2302 1341 2303 1345
rect 2307 1341 2308 1345
rect 2302 1340 2308 1341
rect 2046 1339 2052 1340
rect 1751 1314 1755 1315
rect 1751 1309 1755 1310
rect 1903 1314 1907 1315
rect 1903 1309 1907 1310
rect 2007 1314 2011 1315
rect 2048 1311 2050 1339
rect 2072 1311 2074 1340
rect 2304 1311 2306 1340
rect 2007 1309 2011 1310
rect 2047 1310 2051 1311
rect 2008 1289 2010 1309
rect 2047 1305 2051 1306
rect 2071 1310 2075 1311
rect 2071 1305 2075 1306
rect 2223 1310 2227 1311
rect 2223 1305 2227 1306
rect 2303 1310 2307 1311
rect 2303 1305 2307 1306
rect 2006 1288 2012 1289
rect 2006 1284 2007 1288
rect 2011 1284 2012 1288
rect 2048 1285 2050 1305
rect 2006 1283 2012 1284
rect 2046 1284 2052 1285
rect 2072 1284 2074 1305
rect 2224 1284 2226 1305
rect 2046 1280 2047 1284
rect 2051 1280 2052 1284
rect 2046 1279 2052 1280
rect 2070 1283 2076 1284
rect 2070 1279 2071 1283
rect 2075 1279 2076 1283
rect 2070 1278 2076 1279
rect 2222 1283 2228 1284
rect 2222 1279 2223 1283
rect 2227 1279 2228 1283
rect 2222 1278 2228 1279
rect 2312 1276 2314 1382
rect 2560 1365 2562 1389
rect 2628 1388 2630 1430
rect 2684 1424 2686 1446
rect 2702 1444 2708 1445
rect 2702 1440 2703 1444
rect 2707 1440 2708 1444
rect 2702 1439 2708 1440
rect 2682 1423 2688 1424
rect 2682 1419 2683 1423
rect 2687 1419 2688 1423
rect 2682 1418 2688 1419
rect 2704 1395 2706 1439
rect 2780 1424 2782 1446
rect 2798 1444 2804 1445
rect 2798 1440 2799 1444
rect 2803 1440 2804 1444
rect 2798 1439 2804 1440
rect 2778 1423 2784 1424
rect 2778 1419 2779 1423
rect 2783 1419 2784 1423
rect 2778 1418 2784 1419
rect 2800 1395 2802 1439
rect 2876 1424 2878 1446
rect 2918 1444 2924 1445
rect 2918 1440 2919 1444
rect 2923 1440 2924 1444
rect 2918 1439 2924 1440
rect 2874 1423 2880 1424
rect 2874 1419 2875 1423
rect 2879 1419 2880 1423
rect 2874 1418 2880 1419
rect 2920 1395 2922 1439
rect 2996 1424 2998 1446
rect 2994 1423 3000 1424
rect 2994 1419 2995 1423
rect 2999 1419 3000 1423
rect 2994 1418 3000 1419
rect 3020 1416 3022 1522
rect 3062 1517 3068 1518
rect 3062 1513 3063 1517
rect 3067 1513 3068 1517
rect 3062 1512 3068 1513
rect 3222 1517 3228 1518
rect 3222 1513 3223 1517
rect 3227 1513 3228 1517
rect 3222 1512 3228 1513
rect 3382 1517 3388 1518
rect 3382 1513 3383 1517
rect 3387 1513 3388 1517
rect 3382 1512 3388 1513
rect 3542 1517 3548 1518
rect 3542 1513 3543 1517
rect 3547 1513 3548 1517
rect 3542 1512 3548 1513
rect 3702 1517 3708 1518
rect 3702 1513 3703 1517
rect 3707 1513 3708 1517
rect 3702 1512 3708 1513
rect 3064 1491 3066 1512
rect 3224 1491 3226 1512
rect 3384 1491 3386 1512
rect 3544 1491 3546 1512
rect 3704 1491 3706 1512
rect 3063 1490 3067 1491
rect 3063 1485 3067 1486
rect 3223 1490 3227 1491
rect 3223 1485 3227 1486
rect 3231 1490 3235 1491
rect 3231 1485 3235 1486
rect 3383 1490 3387 1491
rect 3383 1485 3387 1486
rect 3415 1490 3419 1491
rect 3415 1485 3419 1486
rect 3543 1490 3547 1491
rect 3543 1485 3547 1486
rect 3615 1490 3619 1491
rect 3615 1485 3619 1486
rect 3703 1490 3707 1491
rect 3703 1485 3707 1486
rect 3815 1490 3819 1491
rect 3815 1485 3819 1486
rect 3064 1464 3066 1485
rect 3232 1464 3234 1485
rect 3416 1464 3418 1485
rect 3616 1464 3618 1485
rect 3816 1464 3818 1485
rect 3062 1463 3068 1464
rect 3062 1459 3063 1463
rect 3067 1459 3068 1463
rect 3062 1458 3068 1459
rect 3230 1463 3236 1464
rect 3230 1459 3231 1463
rect 3235 1459 3236 1463
rect 3230 1458 3236 1459
rect 3414 1463 3420 1464
rect 3414 1459 3415 1463
rect 3419 1459 3420 1463
rect 3414 1458 3420 1459
rect 3614 1463 3620 1464
rect 3614 1459 3615 1463
rect 3619 1459 3620 1463
rect 3614 1458 3620 1459
rect 3814 1463 3820 1464
rect 3814 1459 3815 1463
rect 3819 1459 3820 1463
rect 3814 1458 3820 1459
rect 3892 1456 3894 1570
rect 3944 1567 3946 1598
rect 3943 1566 3947 1567
rect 3943 1561 3947 1562
rect 3944 1534 3946 1561
rect 3942 1533 3948 1534
rect 3942 1529 3943 1533
rect 3947 1529 3948 1533
rect 3942 1528 3948 1529
rect 3942 1516 3948 1517
rect 3942 1512 3943 1516
rect 3947 1512 3948 1516
rect 3942 1511 3948 1512
rect 3944 1491 3946 1511
rect 3943 1490 3947 1491
rect 3943 1485 3947 1486
rect 3944 1465 3946 1485
rect 3942 1464 3948 1465
rect 3942 1460 3943 1464
rect 3947 1460 3948 1464
rect 3942 1459 3948 1460
rect 3558 1455 3564 1456
rect 3138 1451 3144 1452
rect 3138 1447 3139 1451
rect 3143 1447 3144 1451
rect 3138 1446 3144 1447
rect 3306 1451 3312 1452
rect 3306 1447 3307 1451
rect 3311 1447 3312 1451
rect 3306 1446 3312 1447
rect 3490 1451 3496 1452
rect 3490 1447 3491 1451
rect 3495 1447 3496 1451
rect 3558 1451 3559 1455
rect 3563 1451 3564 1455
rect 3558 1450 3564 1451
rect 3890 1455 3896 1456
rect 3890 1451 3891 1455
rect 3895 1451 3896 1455
rect 3890 1450 3896 1451
rect 3490 1446 3496 1447
rect 3062 1444 3068 1445
rect 3062 1440 3063 1444
rect 3067 1440 3068 1444
rect 3062 1439 3068 1440
rect 3018 1415 3024 1416
rect 3018 1411 3019 1415
rect 3023 1411 3024 1415
rect 3018 1410 3024 1411
rect 3064 1395 3066 1439
rect 3140 1424 3142 1446
rect 3230 1444 3236 1445
rect 3230 1440 3231 1444
rect 3235 1440 3236 1444
rect 3230 1439 3236 1440
rect 3138 1423 3144 1424
rect 3138 1419 3139 1423
rect 3143 1419 3144 1423
rect 3138 1418 3144 1419
rect 3232 1395 3234 1439
rect 3308 1424 3310 1446
rect 3414 1444 3420 1445
rect 3414 1440 3415 1444
rect 3419 1440 3420 1444
rect 3414 1439 3420 1440
rect 3306 1423 3312 1424
rect 3306 1419 3307 1423
rect 3311 1419 3312 1423
rect 3306 1418 3312 1419
rect 3416 1395 3418 1439
rect 3492 1424 3494 1446
rect 3560 1436 3562 1450
rect 3942 1447 3948 1448
rect 3614 1444 3620 1445
rect 3614 1440 3615 1444
rect 3619 1440 3620 1444
rect 3614 1439 3620 1440
rect 3814 1444 3820 1445
rect 3814 1440 3815 1444
rect 3819 1440 3820 1444
rect 3942 1443 3943 1447
rect 3947 1443 3948 1447
rect 3942 1442 3948 1443
rect 3814 1439 3820 1440
rect 3558 1435 3564 1436
rect 3558 1431 3559 1435
rect 3563 1431 3564 1435
rect 3558 1430 3564 1431
rect 3490 1423 3496 1424
rect 3490 1419 3491 1423
rect 3495 1419 3496 1423
rect 3490 1418 3496 1419
rect 3616 1395 3618 1439
rect 3816 1395 3818 1439
rect 3882 1419 3888 1420
rect 3882 1415 3883 1419
rect 3887 1415 3888 1419
rect 3882 1414 3888 1415
rect 2703 1394 2707 1395
rect 2703 1389 2707 1390
rect 2799 1394 2803 1395
rect 2799 1389 2803 1390
rect 2807 1394 2811 1395
rect 2807 1389 2811 1390
rect 2919 1394 2923 1395
rect 2919 1389 2923 1390
rect 3055 1394 3059 1395
rect 3055 1389 3059 1390
rect 3063 1394 3067 1395
rect 3063 1389 3067 1390
rect 3231 1394 3235 1395
rect 3231 1389 3235 1390
rect 3303 1394 3307 1395
rect 3303 1389 3307 1390
rect 3415 1394 3419 1395
rect 3415 1389 3419 1390
rect 3559 1394 3563 1395
rect 3559 1389 3563 1390
rect 3615 1394 3619 1395
rect 3615 1389 3619 1390
rect 3815 1394 3819 1395
rect 3815 1389 3819 1390
rect 2626 1387 2632 1388
rect 2626 1383 2627 1387
rect 2631 1383 2632 1387
rect 2626 1382 2632 1383
rect 2634 1387 2640 1388
rect 2634 1383 2635 1387
rect 2639 1383 2640 1387
rect 2634 1382 2640 1383
rect 2558 1364 2564 1365
rect 2558 1360 2559 1364
rect 2563 1360 2564 1364
rect 2558 1359 2564 1360
rect 2636 1356 2638 1382
rect 2808 1365 2810 1389
rect 2882 1387 2888 1388
rect 2882 1383 2883 1387
rect 2887 1383 2888 1387
rect 2882 1382 2888 1383
rect 2806 1364 2812 1365
rect 2806 1360 2807 1364
rect 2811 1360 2812 1364
rect 2806 1359 2812 1360
rect 2884 1356 2886 1382
rect 3056 1365 3058 1389
rect 3130 1387 3136 1388
rect 3130 1383 3131 1387
rect 3135 1383 3136 1387
rect 3130 1382 3136 1383
rect 3054 1364 3060 1365
rect 3054 1360 3055 1364
rect 3059 1360 3060 1364
rect 3054 1359 3060 1360
rect 3132 1356 3134 1382
rect 3304 1365 3306 1389
rect 3378 1387 3384 1388
rect 3378 1383 3379 1387
rect 3383 1383 3384 1387
rect 3378 1382 3384 1383
rect 3302 1364 3308 1365
rect 3302 1360 3303 1364
rect 3307 1360 3308 1364
rect 3302 1359 3308 1360
rect 3380 1356 3382 1382
rect 3560 1365 3562 1389
rect 3816 1365 3818 1389
rect 3558 1364 3564 1365
rect 3558 1360 3559 1364
rect 3563 1360 3564 1364
rect 3558 1359 3564 1360
rect 3814 1364 3820 1365
rect 3814 1360 3815 1364
rect 3819 1360 3820 1364
rect 3814 1359 3820 1360
rect 3884 1356 3886 1414
rect 3944 1395 3946 1442
rect 3943 1394 3947 1395
rect 3943 1389 3947 1390
rect 3906 1387 3912 1388
rect 3906 1383 3907 1387
rect 3911 1383 3912 1387
rect 3906 1382 3912 1383
rect 2634 1355 2640 1356
rect 2634 1351 2635 1355
rect 2639 1351 2640 1355
rect 2634 1350 2640 1351
rect 2882 1355 2888 1356
rect 2882 1351 2883 1355
rect 2887 1351 2888 1355
rect 2882 1350 2888 1351
rect 3130 1355 3136 1356
rect 3130 1351 3131 1355
rect 3135 1351 3136 1355
rect 3130 1350 3136 1351
rect 3378 1355 3384 1356
rect 3378 1351 3379 1355
rect 3383 1351 3384 1355
rect 3378 1350 3384 1351
rect 3882 1355 3888 1356
rect 3882 1351 3883 1355
rect 3887 1351 3888 1355
rect 3882 1350 3888 1351
rect 2558 1345 2564 1346
rect 2558 1341 2559 1345
rect 2563 1341 2564 1345
rect 2558 1340 2564 1341
rect 2806 1345 2812 1346
rect 2806 1341 2807 1345
rect 2811 1341 2812 1345
rect 2806 1340 2812 1341
rect 3054 1345 3060 1346
rect 3054 1341 3055 1345
rect 3059 1341 3060 1345
rect 3054 1340 3060 1341
rect 3302 1345 3308 1346
rect 3302 1341 3303 1345
rect 3307 1341 3308 1345
rect 3302 1340 3308 1341
rect 3558 1345 3564 1346
rect 3558 1341 3559 1345
rect 3563 1341 3564 1345
rect 3558 1340 3564 1341
rect 3814 1345 3820 1346
rect 3814 1341 3815 1345
rect 3819 1341 3820 1345
rect 3814 1340 3820 1341
rect 2560 1311 2562 1340
rect 2808 1311 2810 1340
rect 3056 1311 3058 1340
rect 3304 1311 3306 1340
rect 3560 1311 3562 1340
rect 3816 1311 3818 1340
rect 2415 1310 2419 1311
rect 2415 1305 2419 1306
rect 2559 1310 2563 1311
rect 2559 1305 2563 1306
rect 2615 1310 2619 1311
rect 2615 1305 2619 1306
rect 2807 1310 2811 1311
rect 2807 1305 2811 1306
rect 2815 1310 2819 1311
rect 2815 1305 2819 1306
rect 2999 1310 3003 1311
rect 2999 1305 3003 1306
rect 3055 1310 3059 1311
rect 3055 1305 3059 1306
rect 3175 1310 3179 1311
rect 3175 1305 3179 1306
rect 3303 1310 3307 1311
rect 3303 1305 3307 1306
rect 3343 1310 3347 1311
rect 3343 1305 3347 1306
rect 3503 1310 3507 1311
rect 3503 1305 3507 1306
rect 3559 1310 3563 1311
rect 3559 1305 3563 1306
rect 3663 1310 3667 1311
rect 3663 1305 3667 1306
rect 3815 1310 3819 1311
rect 3815 1305 3819 1306
rect 3831 1310 3835 1311
rect 3831 1305 3835 1306
rect 2416 1284 2418 1305
rect 2616 1284 2618 1305
rect 2816 1284 2818 1305
rect 3000 1284 3002 1305
rect 3054 1299 3060 1300
rect 3054 1295 3055 1299
rect 3059 1295 3060 1299
rect 3054 1294 3060 1295
rect 2414 1283 2420 1284
rect 2414 1279 2415 1283
rect 2419 1279 2420 1283
rect 2414 1278 2420 1279
rect 2614 1283 2620 1284
rect 2614 1279 2615 1283
rect 2619 1279 2620 1283
rect 2614 1278 2620 1279
rect 2814 1283 2820 1284
rect 2814 1279 2815 1283
rect 2819 1279 2820 1283
rect 2814 1278 2820 1279
rect 2998 1283 3004 1284
rect 2998 1279 2999 1283
rect 3003 1279 3004 1283
rect 2998 1278 3004 1279
rect 2310 1275 2316 1276
rect 2006 1271 2012 1272
rect 2006 1267 2007 1271
rect 2011 1267 2012 1271
rect 2146 1271 2152 1272
rect 2006 1266 2012 1267
rect 2046 1267 2052 1268
rect 1650 1247 1656 1248
rect 1650 1243 1651 1247
rect 1655 1243 1656 1247
rect 1650 1242 1656 1243
rect 2008 1239 2010 1266
rect 2046 1263 2047 1267
rect 2051 1263 2052 1267
rect 2146 1267 2147 1271
rect 2151 1267 2152 1271
rect 2310 1271 2311 1275
rect 2315 1271 2316 1275
rect 2310 1270 2316 1271
rect 2358 1275 2364 1276
rect 2358 1271 2359 1275
rect 2363 1271 2364 1275
rect 2698 1275 2704 1276
rect 2358 1270 2364 1271
rect 2690 1271 2696 1272
rect 2146 1266 2152 1267
rect 2046 1262 2052 1263
rect 2070 1264 2076 1265
rect 1559 1238 1563 1239
rect 1559 1233 1563 1234
rect 1711 1238 1715 1239
rect 1711 1233 1715 1234
rect 2007 1238 2011 1239
rect 2007 1233 2011 1234
rect 1514 1231 1520 1232
rect 1514 1227 1515 1231
rect 1519 1227 1520 1231
rect 1514 1226 1520 1227
rect 1560 1209 1562 1233
rect 1634 1231 1640 1232
rect 1634 1227 1635 1231
rect 1639 1227 1640 1231
rect 1634 1226 1640 1227
rect 1406 1208 1412 1209
rect 1406 1204 1407 1208
rect 1411 1204 1412 1208
rect 1406 1203 1412 1204
rect 1558 1208 1564 1209
rect 1558 1204 1559 1208
rect 1563 1204 1564 1208
rect 1558 1203 1564 1204
rect 1636 1200 1638 1226
rect 1712 1209 1714 1233
rect 1710 1208 1716 1209
rect 1710 1204 1711 1208
rect 1715 1204 1716 1208
rect 2008 1206 2010 1233
rect 2048 1227 2050 1262
rect 2070 1260 2071 1264
rect 2075 1260 2076 1264
rect 2070 1259 2076 1260
rect 2072 1227 2074 1259
rect 2148 1244 2150 1266
rect 2222 1264 2228 1265
rect 2222 1260 2223 1264
rect 2227 1260 2228 1264
rect 2222 1259 2228 1260
rect 2146 1243 2152 1244
rect 2146 1239 2147 1243
rect 2151 1239 2152 1243
rect 2146 1238 2152 1239
rect 2224 1227 2226 1259
rect 2360 1252 2362 1270
rect 2690 1267 2691 1271
rect 2695 1267 2696 1271
rect 2698 1271 2699 1275
rect 2703 1271 2704 1275
rect 2698 1270 2704 1271
rect 2690 1266 2696 1267
rect 2414 1264 2420 1265
rect 2414 1260 2415 1264
rect 2419 1260 2420 1264
rect 2414 1259 2420 1260
rect 2614 1264 2620 1265
rect 2614 1260 2615 1264
rect 2619 1260 2620 1264
rect 2614 1259 2620 1260
rect 2358 1251 2364 1252
rect 2358 1247 2359 1251
rect 2363 1247 2364 1251
rect 2358 1246 2364 1247
rect 2416 1227 2418 1259
rect 2578 1239 2584 1240
rect 2578 1235 2579 1239
rect 2583 1235 2584 1239
rect 2578 1234 2584 1235
rect 2047 1226 2051 1227
rect 2047 1221 2051 1222
rect 2071 1226 2075 1227
rect 2071 1221 2075 1222
rect 2135 1226 2139 1227
rect 2135 1221 2139 1222
rect 2223 1226 2227 1227
rect 2223 1221 2227 1222
rect 2311 1226 2315 1227
rect 2311 1221 2315 1222
rect 2415 1226 2419 1227
rect 2415 1221 2419 1222
rect 2503 1226 2507 1227
rect 2503 1221 2507 1222
rect 1710 1203 1716 1204
rect 2006 1205 2012 1206
rect 2006 1201 2007 1205
rect 2011 1201 2012 1205
rect 2006 1200 2012 1201
rect 1634 1199 1640 1200
rect 1634 1195 1635 1199
rect 1639 1195 1640 1199
rect 1634 1194 1640 1195
rect 1662 1199 1668 1200
rect 1662 1195 1663 1199
rect 1667 1195 1668 1199
rect 1662 1194 1668 1195
rect 2048 1194 2050 1221
rect 2136 1197 2138 1221
rect 2210 1219 2216 1220
rect 2210 1215 2211 1219
rect 2215 1215 2216 1219
rect 2210 1214 2216 1215
rect 2134 1196 2140 1197
rect 1406 1189 1412 1190
rect 1406 1185 1407 1189
rect 1411 1185 1412 1189
rect 1406 1184 1412 1185
rect 1558 1189 1564 1190
rect 1558 1185 1559 1189
rect 1563 1185 1564 1189
rect 1558 1184 1564 1185
rect 1408 1159 1410 1184
rect 1560 1159 1562 1184
rect 1383 1158 1387 1159
rect 1383 1153 1387 1154
rect 1407 1158 1411 1159
rect 1407 1153 1411 1154
rect 1559 1158 1563 1159
rect 1559 1153 1563 1154
rect 1567 1158 1571 1159
rect 1567 1153 1571 1154
rect 1384 1132 1386 1153
rect 1568 1132 1570 1153
rect 1382 1131 1388 1132
rect 1382 1127 1383 1131
rect 1387 1127 1388 1131
rect 1382 1126 1388 1127
rect 1566 1131 1572 1132
rect 1566 1127 1567 1131
rect 1571 1127 1572 1131
rect 1566 1126 1572 1127
rect 1282 1123 1288 1124
rect 1106 1119 1112 1120
rect 1106 1115 1107 1119
rect 1111 1115 1112 1119
rect 1282 1119 1283 1123
rect 1287 1119 1288 1123
rect 1282 1118 1288 1119
rect 1326 1123 1332 1124
rect 1326 1119 1327 1123
rect 1331 1119 1332 1123
rect 1326 1118 1332 1119
rect 1106 1114 1112 1115
rect 1086 1091 1092 1092
rect 1086 1087 1087 1091
rect 1091 1087 1092 1091
rect 1086 1086 1092 1087
rect 327 1074 331 1075
rect 327 1069 331 1070
rect 375 1074 379 1075
rect 375 1069 379 1070
rect 495 1074 499 1075
rect 495 1069 499 1070
rect 543 1074 547 1075
rect 543 1069 547 1070
rect 671 1074 675 1075
rect 671 1069 675 1070
rect 727 1074 731 1075
rect 727 1069 731 1070
rect 847 1074 851 1075
rect 847 1069 851 1070
rect 911 1074 915 1075
rect 911 1069 915 1070
rect 1031 1074 1035 1075
rect 1031 1069 1035 1070
rect 1095 1074 1099 1075
rect 1095 1069 1099 1070
rect 306 1067 312 1068
rect 306 1063 307 1067
rect 311 1063 312 1067
rect 306 1062 312 1063
rect 243 1060 247 1061
rect 243 1055 247 1056
rect 230 1044 236 1045
rect 230 1040 231 1044
rect 235 1040 236 1044
rect 230 1039 236 1040
rect 308 1036 310 1062
rect 376 1045 378 1069
rect 450 1067 456 1068
rect 450 1063 451 1067
rect 455 1063 456 1067
rect 450 1062 456 1063
rect 374 1044 380 1045
rect 374 1040 375 1044
rect 379 1040 380 1044
rect 374 1039 380 1040
rect 452 1036 454 1062
rect 544 1045 546 1069
rect 618 1067 624 1068
rect 618 1063 619 1067
rect 623 1063 624 1067
rect 618 1062 624 1063
rect 542 1044 548 1045
rect 542 1040 543 1044
rect 547 1040 548 1044
rect 542 1039 548 1040
rect 620 1036 622 1062
rect 728 1045 730 1069
rect 802 1067 808 1068
rect 802 1063 803 1067
rect 807 1063 808 1067
rect 802 1062 808 1063
rect 726 1044 732 1045
rect 726 1040 727 1044
rect 731 1040 732 1044
rect 726 1039 732 1040
rect 804 1036 806 1062
rect 859 1060 863 1061
rect 859 1055 863 1056
rect 860 1036 862 1055
rect 912 1045 914 1069
rect 1096 1045 1098 1069
rect 1108 1068 1110 1114
rect 1206 1112 1212 1113
rect 1206 1108 1207 1112
rect 1211 1108 1212 1112
rect 1206 1107 1212 1108
rect 1208 1075 1210 1107
rect 1328 1092 1330 1118
rect 1382 1112 1388 1113
rect 1382 1108 1383 1112
rect 1387 1108 1388 1112
rect 1382 1107 1388 1108
rect 1566 1112 1572 1113
rect 1566 1108 1567 1112
rect 1571 1108 1572 1112
rect 1566 1107 1572 1108
rect 1326 1091 1332 1092
rect 1326 1087 1327 1091
rect 1331 1087 1332 1091
rect 1326 1086 1332 1087
rect 1384 1075 1386 1107
rect 1568 1075 1570 1107
rect 1664 1092 1666 1194
rect 2046 1193 2052 1194
rect 1710 1189 1716 1190
rect 2046 1189 2047 1193
rect 2051 1189 2052 1193
rect 2134 1192 2135 1196
rect 2139 1192 2140 1196
rect 2134 1191 2140 1192
rect 1710 1185 1711 1189
rect 1715 1185 1716 1189
rect 1710 1184 1716 1185
rect 2006 1188 2012 1189
rect 2046 1188 2052 1189
rect 2212 1188 2214 1214
rect 2312 1197 2314 1221
rect 2386 1219 2392 1220
rect 2386 1215 2387 1219
rect 2391 1215 2392 1219
rect 2386 1214 2392 1215
rect 2310 1196 2316 1197
rect 2310 1192 2311 1196
rect 2315 1192 2316 1196
rect 2310 1191 2316 1192
rect 2388 1188 2390 1214
rect 2504 1197 2506 1221
rect 2502 1196 2508 1197
rect 2502 1192 2503 1196
rect 2507 1192 2508 1196
rect 2502 1191 2508 1192
rect 2580 1188 2582 1234
rect 2616 1227 2618 1259
rect 2692 1244 2694 1266
rect 2700 1252 2702 1270
rect 2814 1264 2820 1265
rect 2814 1260 2815 1264
rect 2819 1260 2820 1264
rect 2814 1259 2820 1260
rect 2998 1264 3004 1265
rect 2998 1260 2999 1264
rect 3003 1260 3004 1264
rect 2998 1259 3004 1260
rect 2698 1251 2704 1252
rect 2698 1247 2699 1251
rect 2703 1247 2704 1251
rect 2698 1246 2704 1247
rect 2690 1243 2696 1244
rect 2690 1239 2691 1243
rect 2695 1239 2696 1243
rect 2690 1238 2696 1239
rect 2816 1227 2818 1259
rect 3000 1227 3002 1259
rect 3056 1244 3058 1294
rect 3176 1284 3178 1305
rect 3344 1284 3346 1305
rect 3504 1284 3506 1305
rect 3664 1284 3666 1305
rect 3832 1284 3834 1305
rect 3174 1283 3180 1284
rect 3174 1279 3175 1283
rect 3179 1279 3180 1283
rect 3174 1278 3180 1279
rect 3342 1283 3348 1284
rect 3342 1279 3343 1283
rect 3347 1279 3348 1283
rect 3342 1278 3348 1279
rect 3502 1283 3508 1284
rect 3502 1279 3503 1283
rect 3507 1279 3508 1283
rect 3502 1278 3508 1279
rect 3662 1283 3668 1284
rect 3662 1279 3663 1283
rect 3667 1279 3668 1283
rect 3662 1278 3668 1279
rect 3830 1283 3836 1284
rect 3830 1279 3831 1283
rect 3835 1279 3836 1283
rect 3830 1278 3836 1279
rect 3908 1276 3910 1382
rect 3944 1362 3946 1389
rect 3942 1361 3948 1362
rect 3942 1357 3943 1361
rect 3947 1357 3948 1361
rect 3942 1356 3948 1357
rect 3942 1344 3948 1345
rect 3942 1340 3943 1344
rect 3947 1340 3948 1344
rect 3942 1339 3948 1340
rect 3944 1311 3946 1339
rect 3943 1310 3947 1311
rect 3943 1305 3947 1306
rect 3944 1285 3946 1305
rect 3942 1284 3948 1285
rect 3942 1280 3943 1284
rect 3947 1280 3948 1284
rect 3942 1279 3948 1280
rect 3906 1275 3912 1276
rect 3074 1271 3080 1272
rect 3074 1267 3075 1271
rect 3079 1267 3080 1271
rect 3074 1266 3080 1267
rect 3250 1271 3256 1272
rect 3250 1267 3251 1271
rect 3255 1267 3256 1271
rect 3250 1266 3256 1267
rect 3418 1271 3424 1272
rect 3418 1267 3419 1271
rect 3423 1267 3424 1271
rect 3418 1266 3424 1267
rect 3578 1271 3584 1272
rect 3578 1267 3579 1271
rect 3583 1267 3584 1271
rect 3578 1266 3584 1267
rect 3738 1271 3744 1272
rect 3738 1267 3739 1271
rect 3743 1267 3744 1271
rect 3906 1271 3907 1275
rect 3911 1271 3912 1275
rect 3906 1270 3912 1271
rect 3738 1266 3744 1267
rect 3942 1267 3948 1268
rect 3076 1244 3078 1266
rect 3174 1264 3180 1265
rect 3174 1260 3175 1264
rect 3179 1260 3180 1264
rect 3174 1259 3180 1260
rect 3054 1243 3060 1244
rect 3054 1239 3055 1243
rect 3059 1239 3060 1243
rect 3054 1238 3060 1239
rect 3074 1243 3080 1244
rect 3074 1239 3075 1243
rect 3079 1239 3080 1243
rect 3074 1238 3080 1239
rect 3176 1227 3178 1259
rect 3252 1244 3254 1266
rect 3342 1264 3348 1265
rect 3342 1260 3343 1264
rect 3347 1260 3348 1264
rect 3342 1259 3348 1260
rect 3250 1243 3256 1244
rect 3250 1239 3251 1243
rect 3255 1239 3256 1243
rect 3250 1238 3256 1239
rect 3344 1227 3346 1259
rect 3420 1244 3422 1266
rect 3502 1264 3508 1265
rect 3502 1260 3503 1264
rect 3507 1260 3508 1264
rect 3502 1259 3508 1260
rect 3418 1243 3424 1244
rect 3418 1239 3419 1243
rect 3423 1239 3424 1243
rect 3418 1238 3424 1239
rect 3504 1227 3506 1259
rect 3580 1244 3582 1266
rect 3662 1264 3668 1265
rect 3662 1260 3663 1264
rect 3667 1260 3668 1264
rect 3662 1259 3668 1260
rect 3578 1243 3584 1244
rect 3578 1239 3579 1243
rect 3583 1239 3584 1243
rect 3578 1238 3584 1239
rect 3664 1227 3666 1259
rect 2615 1226 2619 1227
rect 2615 1221 2619 1222
rect 2695 1226 2699 1227
rect 2695 1221 2699 1222
rect 2815 1226 2819 1227
rect 2815 1221 2819 1222
rect 2887 1226 2891 1227
rect 2887 1221 2891 1222
rect 2999 1226 3003 1227
rect 2999 1221 3003 1222
rect 3071 1226 3075 1227
rect 3071 1221 3075 1222
rect 3175 1226 3179 1227
rect 3175 1221 3179 1222
rect 3239 1226 3243 1227
rect 3239 1221 3243 1222
rect 3343 1226 3347 1227
rect 3343 1221 3347 1222
rect 3399 1226 3403 1227
rect 3399 1221 3403 1222
rect 3503 1226 3507 1227
rect 3503 1221 3507 1222
rect 3551 1226 3555 1227
rect 3551 1221 3555 1222
rect 3663 1226 3667 1227
rect 3663 1221 3667 1222
rect 3703 1226 3707 1227
rect 3703 1221 3707 1222
rect 2658 1211 2664 1212
rect 2658 1207 2659 1211
rect 2663 1207 2664 1211
rect 2658 1206 2664 1207
rect 2660 1188 2662 1206
rect 2696 1197 2698 1221
rect 2888 1197 2890 1221
rect 2914 1219 2920 1220
rect 2914 1215 2915 1219
rect 2919 1215 2920 1219
rect 2914 1214 2920 1215
rect 2694 1196 2700 1197
rect 2694 1192 2695 1196
rect 2699 1192 2700 1196
rect 2694 1191 2700 1192
rect 2886 1196 2892 1197
rect 2886 1192 2887 1196
rect 2891 1192 2892 1196
rect 2886 1191 2892 1192
rect 2006 1184 2007 1188
rect 2011 1184 2012 1188
rect 1712 1159 1714 1184
rect 2006 1183 2012 1184
rect 2210 1187 2216 1188
rect 2210 1183 2211 1187
rect 2215 1183 2216 1187
rect 2008 1159 2010 1183
rect 2210 1182 2216 1183
rect 2386 1187 2392 1188
rect 2386 1183 2387 1187
rect 2391 1183 2392 1187
rect 2386 1182 2392 1183
rect 2578 1187 2584 1188
rect 2578 1183 2579 1187
rect 2583 1183 2584 1187
rect 2578 1182 2584 1183
rect 2658 1187 2664 1188
rect 2658 1183 2659 1187
rect 2663 1183 2664 1187
rect 2658 1182 2664 1183
rect 2134 1177 2140 1178
rect 2046 1176 2052 1177
rect 2046 1172 2047 1176
rect 2051 1172 2052 1176
rect 2134 1173 2135 1177
rect 2139 1173 2140 1177
rect 2134 1172 2140 1173
rect 2310 1177 2316 1178
rect 2310 1173 2311 1177
rect 2315 1173 2316 1177
rect 2310 1172 2316 1173
rect 2502 1177 2508 1178
rect 2502 1173 2503 1177
rect 2507 1173 2508 1177
rect 2502 1172 2508 1173
rect 2694 1177 2700 1178
rect 2694 1173 2695 1177
rect 2699 1173 2700 1177
rect 2694 1172 2700 1173
rect 2886 1177 2892 1178
rect 2886 1173 2887 1177
rect 2891 1173 2892 1177
rect 2886 1172 2892 1173
rect 2046 1171 2052 1172
rect 1711 1158 1715 1159
rect 1711 1153 1715 1154
rect 1751 1158 1755 1159
rect 1751 1153 1755 1154
rect 2007 1158 2011 1159
rect 2007 1153 2011 1154
rect 1752 1132 1754 1153
rect 2008 1133 2010 1153
rect 2048 1143 2050 1171
rect 2136 1143 2138 1172
rect 2312 1143 2314 1172
rect 2504 1143 2506 1172
rect 2696 1143 2698 1172
rect 2888 1143 2890 1172
rect 2047 1142 2051 1143
rect 2047 1137 2051 1138
rect 2135 1142 2139 1143
rect 2135 1137 2139 1138
rect 2295 1142 2299 1143
rect 2295 1137 2299 1138
rect 2311 1142 2315 1143
rect 2311 1137 2315 1138
rect 2423 1142 2427 1143
rect 2423 1137 2427 1138
rect 2503 1142 2507 1143
rect 2503 1137 2507 1138
rect 2559 1142 2563 1143
rect 2559 1137 2563 1138
rect 2695 1142 2699 1143
rect 2695 1137 2699 1138
rect 2839 1142 2843 1143
rect 2839 1137 2843 1138
rect 2887 1142 2891 1143
rect 2887 1137 2891 1138
rect 2006 1132 2012 1133
rect 1750 1131 1756 1132
rect 1750 1127 1751 1131
rect 1755 1127 1756 1131
rect 2006 1128 2007 1132
rect 2011 1128 2012 1132
rect 2006 1127 2012 1128
rect 1750 1126 1756 1127
rect 1838 1119 1844 1120
rect 1838 1115 1839 1119
rect 1843 1115 1844 1119
rect 2048 1117 2050 1137
rect 2046 1116 2052 1117
rect 2296 1116 2298 1137
rect 2424 1116 2426 1137
rect 2560 1116 2562 1137
rect 2696 1116 2698 1137
rect 2840 1116 2842 1137
rect 1838 1114 1844 1115
rect 2006 1115 2012 1116
rect 1750 1112 1756 1113
rect 1750 1108 1751 1112
rect 1755 1108 1756 1112
rect 1750 1107 1756 1108
rect 1662 1091 1668 1092
rect 1662 1087 1663 1091
rect 1667 1087 1668 1091
rect 1662 1086 1668 1087
rect 1752 1075 1754 1107
rect 1207 1074 1211 1075
rect 1207 1069 1211 1070
rect 1279 1074 1283 1075
rect 1279 1069 1283 1070
rect 1383 1074 1387 1075
rect 1383 1069 1387 1070
rect 1463 1074 1467 1075
rect 1463 1069 1467 1070
rect 1567 1074 1571 1075
rect 1567 1069 1571 1070
rect 1647 1074 1651 1075
rect 1647 1069 1651 1070
rect 1751 1074 1755 1075
rect 1751 1069 1755 1070
rect 1831 1074 1835 1075
rect 1831 1069 1835 1070
rect 1106 1067 1112 1068
rect 1106 1063 1107 1067
rect 1111 1063 1112 1067
rect 1106 1062 1112 1063
rect 1280 1045 1282 1069
rect 1326 1067 1332 1068
rect 1326 1063 1327 1067
rect 1331 1063 1332 1067
rect 1326 1062 1332 1063
rect 1354 1067 1360 1068
rect 1354 1063 1355 1067
rect 1359 1063 1360 1067
rect 1354 1062 1360 1063
rect 910 1044 916 1045
rect 910 1040 911 1044
rect 915 1040 916 1044
rect 910 1039 916 1040
rect 1094 1044 1100 1045
rect 1094 1040 1095 1044
rect 1099 1040 1100 1044
rect 1094 1039 1100 1040
rect 1278 1044 1284 1045
rect 1278 1040 1279 1044
rect 1283 1040 1284 1044
rect 1278 1039 1284 1040
rect 210 1035 216 1036
rect 210 1031 211 1035
rect 215 1031 216 1035
rect 210 1030 216 1031
rect 306 1035 312 1036
rect 306 1031 307 1035
rect 311 1031 312 1035
rect 306 1030 312 1031
rect 450 1035 456 1036
rect 450 1031 451 1035
rect 455 1031 456 1035
rect 450 1030 456 1031
rect 618 1035 624 1036
rect 618 1031 619 1035
rect 623 1031 624 1035
rect 618 1030 624 1031
rect 802 1035 808 1036
rect 802 1031 803 1035
rect 807 1031 808 1035
rect 802 1030 808 1031
rect 858 1035 864 1036
rect 858 1031 859 1035
rect 863 1031 864 1035
rect 858 1030 864 1031
rect 1062 1035 1068 1036
rect 1062 1031 1063 1035
rect 1067 1031 1068 1035
rect 1062 1030 1068 1031
rect 230 1025 236 1026
rect 230 1021 231 1025
rect 235 1021 236 1025
rect 230 1020 236 1021
rect 374 1025 380 1026
rect 374 1021 375 1025
rect 379 1021 380 1025
rect 374 1020 380 1021
rect 542 1025 548 1026
rect 542 1021 543 1025
rect 547 1021 548 1025
rect 542 1020 548 1021
rect 726 1025 732 1026
rect 726 1021 727 1025
rect 731 1021 732 1025
rect 726 1020 732 1021
rect 910 1025 916 1026
rect 910 1021 911 1025
rect 915 1021 916 1025
rect 910 1020 916 1021
rect 232 999 234 1020
rect 376 999 378 1020
rect 544 999 546 1020
rect 728 999 730 1020
rect 912 999 914 1020
rect 231 998 235 999
rect 231 993 235 994
rect 271 998 275 999
rect 271 993 275 994
rect 375 998 379 999
rect 375 993 379 994
rect 447 998 451 999
rect 447 993 451 994
rect 543 998 547 999
rect 543 993 547 994
rect 631 998 635 999
rect 631 993 635 994
rect 727 998 731 999
rect 727 993 731 994
rect 823 998 827 999
rect 823 993 827 994
rect 911 998 915 999
rect 911 993 915 994
rect 1007 998 1011 999
rect 1007 993 1011 994
rect 272 972 274 993
rect 448 972 450 993
rect 632 972 634 993
rect 824 972 826 993
rect 1008 972 1010 993
rect 270 971 276 972
rect 134 966 140 967
rect 202 967 208 968
rect 202 963 203 967
rect 207 963 208 967
rect 270 967 271 971
rect 275 967 276 971
rect 270 966 276 967
rect 446 971 452 972
rect 446 967 447 971
rect 451 967 452 971
rect 446 966 452 967
rect 630 971 636 972
rect 630 967 631 971
rect 635 967 636 971
rect 630 966 636 967
rect 822 971 828 972
rect 822 967 823 971
rect 827 967 828 971
rect 822 966 828 967
rect 1006 971 1012 972
rect 1006 967 1007 971
rect 1011 967 1012 971
rect 1006 966 1012 967
rect 202 962 208 963
rect 250 963 256 964
rect 250 959 251 963
rect 255 959 256 963
rect 250 958 256 959
rect 586 963 592 964
rect 586 959 587 963
rect 591 959 592 963
rect 586 958 592 959
rect 714 963 720 964
rect 714 959 715 963
rect 719 959 720 963
rect 714 958 720 959
rect 110 955 116 956
rect 110 951 111 955
rect 115 951 116 955
rect 110 950 116 951
rect 134 952 140 953
rect 112 923 114 950
rect 134 948 135 952
rect 139 948 140 952
rect 134 947 140 948
rect 136 923 138 947
rect 252 932 254 958
rect 270 952 276 953
rect 270 948 271 952
rect 275 948 276 952
rect 270 947 276 948
rect 446 952 452 953
rect 446 948 447 952
rect 451 948 452 952
rect 446 947 452 948
rect 250 931 256 932
rect 250 927 251 931
rect 255 927 256 931
rect 250 926 256 927
rect 272 923 274 947
rect 448 923 450 947
rect 588 932 590 958
rect 630 952 636 953
rect 630 948 631 952
rect 635 948 636 952
rect 630 947 636 948
rect 586 931 592 932
rect 586 927 587 931
rect 591 927 592 931
rect 586 926 592 927
rect 632 923 634 947
rect 716 932 718 958
rect 822 952 828 953
rect 822 948 823 952
rect 827 948 828 952
rect 822 947 828 948
rect 1006 952 1012 953
rect 1006 948 1007 952
rect 1011 948 1012 952
rect 1006 947 1012 948
rect 714 931 720 932
rect 714 927 715 931
rect 719 927 720 931
rect 714 926 720 927
rect 824 923 826 947
rect 922 927 928 928
rect 922 923 923 927
rect 927 923 928 927
rect 1008 923 1010 947
rect 1064 932 1066 1030
rect 1094 1025 1100 1026
rect 1094 1021 1095 1025
rect 1099 1021 1100 1025
rect 1094 1020 1100 1021
rect 1278 1025 1284 1026
rect 1278 1021 1279 1025
rect 1283 1021 1284 1025
rect 1278 1020 1284 1021
rect 1096 999 1098 1020
rect 1280 999 1282 1020
rect 1095 998 1099 999
rect 1095 993 1099 994
rect 1175 998 1179 999
rect 1175 993 1179 994
rect 1279 998 1283 999
rect 1279 993 1283 994
rect 1176 972 1178 993
rect 1174 971 1180 972
rect 1174 967 1175 971
rect 1179 967 1180 971
rect 1174 966 1180 967
rect 1328 964 1330 1062
rect 1356 1036 1358 1062
rect 1464 1045 1466 1069
rect 1648 1045 1650 1069
rect 1734 1067 1740 1068
rect 1734 1063 1735 1067
rect 1739 1063 1740 1067
rect 1734 1062 1740 1063
rect 1462 1044 1468 1045
rect 1462 1040 1463 1044
rect 1467 1040 1468 1044
rect 1462 1039 1468 1040
rect 1646 1044 1652 1045
rect 1646 1040 1647 1044
rect 1651 1040 1652 1044
rect 1646 1039 1652 1040
rect 1736 1036 1738 1062
rect 1832 1045 1834 1069
rect 1840 1068 1842 1114
rect 2006 1111 2007 1115
rect 2011 1111 2012 1115
rect 2046 1112 2047 1116
rect 2051 1112 2052 1116
rect 2046 1111 2052 1112
rect 2294 1115 2300 1116
rect 2294 1111 2295 1115
rect 2299 1111 2300 1115
rect 2006 1110 2012 1111
rect 2294 1110 2300 1111
rect 2422 1115 2428 1116
rect 2422 1111 2423 1115
rect 2427 1111 2428 1115
rect 2422 1110 2428 1111
rect 2558 1115 2564 1116
rect 2558 1111 2559 1115
rect 2563 1111 2564 1115
rect 2558 1110 2564 1111
rect 2694 1115 2700 1116
rect 2694 1111 2695 1115
rect 2699 1111 2700 1115
rect 2694 1110 2700 1111
rect 2838 1115 2844 1116
rect 2838 1111 2839 1115
rect 2843 1111 2844 1115
rect 2838 1110 2844 1111
rect 2008 1075 2010 1110
rect 2916 1108 2918 1214
rect 3072 1197 3074 1221
rect 3146 1219 3152 1220
rect 3146 1215 3147 1219
rect 3151 1215 3152 1219
rect 3146 1214 3152 1215
rect 3070 1196 3076 1197
rect 3070 1192 3071 1196
rect 3075 1192 3076 1196
rect 3070 1191 3076 1192
rect 3148 1188 3150 1214
rect 3240 1197 3242 1221
rect 3314 1219 3320 1220
rect 3314 1215 3315 1219
rect 3319 1215 3320 1219
rect 3314 1214 3320 1215
rect 3238 1196 3244 1197
rect 3238 1192 3239 1196
rect 3243 1192 3244 1196
rect 3238 1191 3244 1192
rect 3316 1188 3318 1214
rect 3400 1197 3402 1221
rect 3498 1211 3504 1212
rect 3498 1207 3499 1211
rect 3503 1207 3504 1211
rect 3498 1206 3504 1207
rect 3398 1196 3404 1197
rect 3398 1192 3399 1196
rect 3403 1192 3404 1196
rect 3398 1191 3404 1192
rect 3500 1188 3502 1206
rect 3552 1197 3554 1221
rect 3704 1197 3706 1221
rect 3740 1220 3742 1266
rect 3830 1264 3836 1265
rect 3830 1260 3831 1264
rect 3835 1260 3836 1264
rect 3942 1263 3943 1267
rect 3947 1263 3948 1267
rect 3942 1262 3948 1263
rect 3830 1259 3836 1260
rect 3832 1227 3834 1259
rect 3906 1239 3912 1240
rect 3906 1235 3907 1239
rect 3911 1235 3912 1239
rect 3906 1234 3912 1235
rect 3831 1226 3835 1227
rect 3831 1221 3835 1222
rect 3839 1226 3843 1227
rect 3839 1221 3843 1222
rect 3738 1219 3744 1220
rect 3738 1215 3739 1219
rect 3743 1215 3744 1219
rect 3738 1214 3744 1215
rect 3840 1197 3842 1221
rect 3550 1196 3556 1197
rect 3550 1192 3551 1196
rect 3555 1192 3556 1196
rect 3550 1191 3556 1192
rect 3702 1196 3708 1197
rect 3702 1192 3703 1196
rect 3707 1192 3708 1196
rect 3702 1191 3708 1192
rect 3838 1196 3844 1197
rect 3838 1192 3839 1196
rect 3843 1192 3844 1196
rect 3838 1191 3844 1192
rect 3908 1188 3910 1234
rect 3944 1227 3946 1262
rect 3943 1226 3947 1227
rect 3943 1221 3947 1222
rect 3914 1219 3920 1220
rect 3914 1215 3915 1219
rect 3919 1215 3920 1219
rect 3914 1214 3920 1215
rect 3146 1187 3152 1188
rect 3146 1183 3147 1187
rect 3151 1183 3152 1187
rect 3146 1182 3152 1183
rect 3314 1187 3320 1188
rect 3314 1183 3315 1187
rect 3319 1183 3320 1187
rect 3314 1182 3320 1183
rect 3474 1187 3480 1188
rect 3474 1183 3475 1187
rect 3479 1183 3480 1187
rect 3474 1182 3480 1183
rect 3498 1187 3504 1188
rect 3498 1183 3499 1187
rect 3503 1183 3504 1187
rect 3498 1182 3504 1183
rect 3906 1187 3912 1188
rect 3906 1183 3907 1187
rect 3911 1183 3912 1187
rect 3906 1182 3912 1183
rect 3070 1177 3076 1178
rect 3070 1173 3071 1177
rect 3075 1173 3076 1177
rect 3070 1172 3076 1173
rect 3238 1177 3244 1178
rect 3238 1173 3239 1177
rect 3243 1173 3244 1177
rect 3238 1172 3244 1173
rect 3398 1177 3404 1178
rect 3398 1173 3399 1177
rect 3403 1173 3404 1177
rect 3398 1172 3404 1173
rect 3072 1143 3074 1172
rect 3240 1143 3242 1172
rect 3400 1143 3402 1172
rect 2991 1142 2995 1143
rect 2991 1137 2995 1138
rect 3071 1142 3075 1143
rect 3071 1137 3075 1138
rect 3151 1142 3155 1143
rect 3151 1137 3155 1138
rect 3239 1142 3243 1143
rect 3239 1137 3243 1138
rect 3319 1142 3323 1143
rect 3319 1137 3323 1138
rect 3399 1142 3403 1143
rect 3399 1137 3403 1138
rect 2992 1116 2994 1137
rect 3152 1116 3154 1137
rect 3320 1116 3322 1137
rect 2990 1115 2996 1116
rect 2990 1111 2991 1115
rect 2995 1111 2996 1115
rect 2990 1110 2996 1111
rect 3150 1115 3156 1116
rect 3150 1111 3151 1115
rect 3155 1111 3156 1115
rect 3150 1110 3156 1111
rect 3318 1115 3324 1116
rect 3318 1111 3319 1115
rect 3323 1111 3324 1115
rect 3318 1110 3324 1111
rect 2914 1107 2920 1108
rect 2370 1103 2376 1104
rect 2046 1099 2052 1100
rect 2046 1095 2047 1099
rect 2051 1095 2052 1099
rect 2370 1099 2371 1103
rect 2375 1099 2376 1103
rect 2370 1098 2376 1099
rect 2498 1103 2504 1104
rect 2498 1099 2499 1103
rect 2503 1099 2504 1103
rect 2498 1098 2504 1099
rect 2634 1103 2640 1104
rect 2634 1099 2635 1103
rect 2639 1099 2640 1103
rect 2634 1098 2640 1099
rect 2770 1103 2776 1104
rect 2770 1099 2771 1103
rect 2775 1099 2776 1103
rect 2914 1103 2915 1107
rect 2919 1103 2920 1107
rect 3258 1107 3264 1108
rect 2914 1102 2920 1103
rect 3066 1103 3072 1104
rect 2770 1098 2776 1099
rect 3066 1099 3067 1103
rect 3071 1099 3072 1103
rect 3066 1098 3072 1099
rect 3226 1103 3232 1104
rect 3226 1099 3227 1103
rect 3231 1099 3232 1103
rect 3258 1103 3259 1107
rect 3263 1103 3264 1107
rect 3258 1102 3264 1103
rect 3226 1098 3232 1099
rect 2046 1094 2052 1095
rect 2294 1096 2300 1097
rect 2007 1074 2011 1075
rect 2007 1069 2011 1070
rect 1838 1067 1844 1068
rect 1838 1063 1839 1067
rect 1843 1063 1844 1067
rect 1838 1062 1844 1063
rect 1830 1044 1836 1045
rect 1830 1040 1831 1044
rect 1835 1040 1836 1044
rect 2008 1042 2010 1069
rect 2048 1063 2050 1094
rect 2294 1092 2295 1096
rect 2299 1092 2300 1096
rect 2294 1091 2300 1092
rect 2296 1063 2298 1091
rect 2372 1080 2374 1098
rect 2422 1096 2428 1097
rect 2422 1092 2423 1096
rect 2427 1092 2428 1096
rect 2422 1091 2428 1092
rect 2370 1079 2376 1080
rect 2370 1075 2371 1079
rect 2375 1075 2376 1079
rect 2370 1074 2376 1075
rect 2424 1063 2426 1091
rect 2500 1076 2502 1098
rect 2558 1096 2564 1097
rect 2558 1092 2559 1096
rect 2563 1092 2564 1096
rect 2558 1091 2564 1092
rect 2498 1075 2504 1076
rect 2498 1071 2499 1075
rect 2503 1071 2504 1075
rect 2498 1070 2504 1071
rect 2560 1063 2562 1091
rect 2636 1076 2638 1098
rect 2694 1096 2700 1097
rect 2694 1092 2695 1096
rect 2699 1092 2700 1096
rect 2694 1091 2700 1092
rect 2634 1075 2640 1076
rect 2634 1071 2635 1075
rect 2639 1071 2640 1075
rect 2634 1070 2640 1071
rect 2696 1063 2698 1091
rect 2772 1076 2774 1098
rect 2838 1096 2844 1097
rect 2838 1092 2839 1096
rect 2843 1092 2844 1096
rect 2838 1091 2844 1092
rect 2990 1096 2996 1097
rect 2990 1092 2991 1096
rect 2995 1092 2996 1096
rect 2990 1091 2996 1092
rect 2770 1075 2776 1076
rect 2770 1071 2771 1075
rect 2775 1071 2776 1075
rect 2770 1070 2776 1071
rect 2840 1063 2842 1091
rect 2992 1063 2994 1091
rect 3068 1076 3070 1098
rect 3150 1096 3156 1097
rect 3150 1092 3151 1096
rect 3155 1092 3156 1096
rect 3150 1091 3156 1092
rect 3066 1075 3072 1076
rect 3066 1071 3067 1075
rect 3071 1071 3072 1075
rect 3066 1070 3072 1071
rect 3152 1063 3154 1091
rect 2047 1062 2051 1063
rect 2047 1057 2051 1058
rect 2295 1062 2299 1063
rect 2295 1057 2299 1058
rect 2423 1062 2427 1063
rect 2423 1057 2427 1058
rect 2495 1062 2499 1063
rect 2495 1057 2499 1058
rect 2559 1062 2563 1063
rect 2559 1057 2563 1058
rect 2599 1062 2603 1063
rect 2599 1057 2603 1058
rect 2695 1062 2699 1063
rect 2695 1057 2699 1058
rect 2711 1062 2715 1063
rect 2711 1057 2715 1058
rect 2839 1062 2843 1063
rect 2839 1057 2843 1058
rect 2847 1062 2851 1063
rect 2847 1057 2851 1058
rect 2991 1062 2995 1063
rect 2991 1057 2995 1058
rect 3007 1062 3011 1063
rect 3007 1057 3011 1058
rect 3151 1062 3155 1063
rect 3151 1057 3155 1058
rect 3199 1062 3203 1063
rect 3199 1057 3203 1058
rect 1830 1039 1836 1040
rect 2006 1041 2012 1042
rect 2006 1037 2007 1041
rect 2011 1037 2012 1041
rect 2006 1036 2012 1037
rect 1354 1035 1360 1036
rect 1354 1031 1355 1035
rect 1359 1031 1360 1035
rect 1354 1030 1360 1031
rect 1554 1035 1560 1036
rect 1554 1031 1555 1035
rect 1559 1031 1560 1035
rect 1554 1030 1560 1031
rect 1734 1035 1740 1036
rect 1734 1031 1735 1035
rect 1739 1031 1740 1035
rect 1734 1030 1740 1031
rect 2048 1030 2050 1057
rect 2496 1033 2498 1057
rect 2578 1055 2584 1056
rect 2578 1051 2579 1055
rect 2583 1051 2584 1055
rect 2578 1050 2584 1051
rect 2494 1032 2500 1033
rect 1462 1025 1468 1026
rect 1462 1021 1463 1025
rect 1467 1021 1468 1025
rect 1462 1020 1468 1021
rect 1464 999 1466 1020
rect 1335 998 1339 999
rect 1335 993 1339 994
rect 1463 998 1467 999
rect 1463 993 1467 994
rect 1487 998 1491 999
rect 1487 993 1491 994
rect 1336 972 1338 993
rect 1488 972 1490 993
rect 1334 971 1340 972
rect 1334 967 1335 971
rect 1339 967 1340 971
rect 1334 966 1340 967
rect 1486 971 1492 972
rect 1486 967 1487 971
rect 1491 967 1492 971
rect 1486 966 1492 967
rect 1326 963 1332 964
rect 1082 959 1088 960
rect 1082 955 1083 959
rect 1087 955 1088 959
rect 1082 954 1088 955
rect 1250 959 1256 960
rect 1250 955 1251 959
rect 1255 955 1256 959
rect 1326 959 1327 963
rect 1331 959 1332 963
rect 1326 958 1332 959
rect 1250 954 1256 955
rect 1062 931 1068 932
rect 1062 927 1063 931
rect 1067 927 1068 931
rect 1062 926 1068 927
rect 111 922 115 923
rect 111 917 115 918
rect 135 922 139 923
rect 135 917 139 918
rect 271 922 275 923
rect 271 917 275 918
rect 447 922 451 923
rect 447 917 451 918
rect 455 922 459 923
rect 455 917 459 918
rect 631 922 635 923
rect 631 917 635 918
rect 655 922 659 923
rect 655 917 659 918
rect 823 922 827 923
rect 823 917 827 918
rect 855 922 859 923
rect 922 922 928 923
rect 1007 922 1011 923
rect 855 917 859 918
rect 112 890 114 917
rect 136 893 138 917
rect 190 915 196 916
rect 190 911 191 915
rect 195 911 196 915
rect 190 910 196 911
rect 210 915 216 916
rect 210 911 211 915
rect 215 911 216 915
rect 210 910 216 911
rect 134 892 140 893
rect 110 889 116 890
rect 110 885 111 889
rect 115 885 116 889
rect 134 888 135 892
rect 139 888 140 892
rect 134 887 140 888
rect 110 884 116 885
rect 134 873 140 874
rect 110 872 116 873
rect 110 868 111 872
rect 115 868 116 872
rect 134 869 135 873
rect 139 869 140 873
rect 134 868 140 869
rect 110 867 116 868
rect 112 847 114 867
rect 136 847 138 868
rect 111 846 115 847
rect 111 841 115 842
rect 135 846 139 847
rect 135 841 139 842
rect 112 821 114 841
rect 110 820 116 821
rect 110 816 111 820
rect 115 816 116 820
rect 110 815 116 816
rect 192 812 194 910
rect 212 884 214 910
rect 272 893 274 917
rect 346 915 352 916
rect 346 911 347 915
rect 351 911 352 915
rect 346 910 352 911
rect 270 892 276 893
rect 270 888 271 892
rect 275 888 276 892
rect 270 887 276 888
rect 348 884 350 910
rect 456 893 458 917
rect 530 915 536 916
rect 530 911 531 915
rect 535 911 536 915
rect 530 910 536 911
rect 454 892 460 893
rect 454 888 455 892
rect 459 888 460 892
rect 454 887 460 888
rect 532 884 534 910
rect 656 893 658 917
rect 730 915 736 916
rect 730 911 731 915
rect 735 911 736 915
rect 730 910 736 911
rect 654 892 660 893
rect 654 888 655 892
rect 659 888 660 892
rect 654 887 660 888
rect 732 884 734 910
rect 856 893 858 917
rect 854 892 860 893
rect 854 888 855 892
rect 859 888 860 892
rect 854 887 860 888
rect 924 884 926 922
rect 1007 917 1011 918
rect 1055 922 1059 923
rect 1055 917 1059 918
rect 1056 893 1058 917
rect 1084 916 1086 954
rect 1174 952 1180 953
rect 1174 948 1175 952
rect 1179 948 1180 952
rect 1174 947 1180 948
rect 1176 923 1178 947
rect 1252 932 1254 954
rect 1334 952 1340 953
rect 1334 948 1335 952
rect 1339 948 1340 952
rect 1334 947 1340 948
rect 1486 952 1492 953
rect 1486 948 1487 952
rect 1491 948 1492 952
rect 1486 947 1492 948
rect 1250 931 1256 932
rect 1230 927 1236 928
rect 1230 923 1231 927
rect 1235 923 1236 927
rect 1250 927 1251 931
rect 1255 927 1256 931
rect 1250 926 1256 927
rect 1336 923 1338 947
rect 1488 923 1490 947
rect 1556 932 1558 1030
rect 2046 1029 2052 1030
rect 1646 1025 1652 1026
rect 1646 1021 1647 1025
rect 1651 1021 1652 1025
rect 1646 1020 1652 1021
rect 1830 1025 1836 1026
rect 2046 1025 2047 1029
rect 2051 1025 2052 1029
rect 2494 1028 2495 1032
rect 2499 1028 2500 1032
rect 2494 1027 2500 1028
rect 1830 1021 1831 1025
rect 1835 1021 1836 1025
rect 1830 1020 1836 1021
rect 2006 1024 2012 1025
rect 2046 1024 2052 1025
rect 2580 1024 2582 1050
rect 2600 1033 2602 1057
rect 2682 1055 2688 1056
rect 2682 1051 2683 1055
rect 2687 1051 2688 1055
rect 2682 1050 2688 1051
rect 2598 1032 2604 1033
rect 2598 1028 2599 1032
rect 2603 1028 2604 1032
rect 2598 1027 2604 1028
rect 2684 1024 2686 1050
rect 2712 1033 2714 1057
rect 2848 1033 2850 1057
rect 2922 1055 2928 1056
rect 2922 1051 2923 1055
rect 2927 1051 2928 1055
rect 2922 1050 2928 1051
rect 2710 1032 2716 1033
rect 2710 1028 2711 1032
rect 2715 1028 2716 1032
rect 2710 1027 2716 1028
rect 2846 1032 2852 1033
rect 2846 1028 2847 1032
rect 2851 1028 2852 1032
rect 2846 1027 2852 1028
rect 2006 1020 2007 1024
rect 2011 1020 2012 1024
rect 1648 999 1650 1020
rect 1832 999 1834 1020
rect 2006 1019 2012 1020
rect 2578 1023 2584 1024
rect 2578 1019 2579 1023
rect 2583 1019 2584 1023
rect 2008 999 2010 1019
rect 2578 1018 2584 1019
rect 2682 1023 2688 1024
rect 2682 1019 2683 1023
rect 2687 1019 2688 1023
rect 2682 1018 2688 1019
rect 2494 1013 2500 1014
rect 2046 1012 2052 1013
rect 2046 1008 2047 1012
rect 2051 1008 2052 1012
rect 2494 1009 2495 1013
rect 2499 1009 2500 1013
rect 2494 1008 2500 1009
rect 2598 1013 2604 1014
rect 2598 1009 2599 1013
rect 2603 1009 2604 1013
rect 2598 1008 2604 1009
rect 2710 1013 2716 1014
rect 2710 1009 2711 1013
rect 2715 1009 2716 1013
rect 2710 1008 2716 1009
rect 2846 1013 2852 1014
rect 2846 1009 2847 1013
rect 2851 1009 2852 1013
rect 2846 1008 2852 1009
rect 2046 1007 2052 1008
rect 1631 998 1635 999
rect 1631 993 1635 994
rect 1647 998 1651 999
rect 1647 993 1651 994
rect 1775 998 1779 999
rect 1775 993 1779 994
rect 1831 998 1835 999
rect 1831 993 1835 994
rect 1903 998 1907 999
rect 1903 993 1907 994
rect 2007 998 2011 999
rect 2007 993 2011 994
rect 1632 972 1634 993
rect 1776 972 1778 993
rect 1904 972 1906 993
rect 2008 973 2010 993
rect 2048 987 2050 1007
rect 2496 987 2498 1008
rect 2600 987 2602 1008
rect 2712 987 2714 1008
rect 2848 987 2850 1008
rect 2047 986 2051 987
rect 2047 981 2051 982
rect 2495 986 2499 987
rect 2495 981 2499 982
rect 2599 986 2603 987
rect 2599 981 2603 982
rect 2647 986 2651 987
rect 2647 981 2651 982
rect 2711 986 2715 987
rect 2711 981 2715 982
rect 2743 986 2747 987
rect 2743 981 2747 982
rect 2847 986 2851 987
rect 2847 981 2851 982
rect 2006 972 2012 973
rect 1630 971 1636 972
rect 1630 967 1631 971
rect 1635 967 1636 971
rect 1630 966 1636 967
rect 1774 971 1780 972
rect 1774 967 1775 971
rect 1779 967 1780 971
rect 1774 966 1780 967
rect 1902 971 1908 972
rect 1902 967 1903 971
rect 1907 967 1908 971
rect 2006 968 2007 972
rect 2011 968 2012 972
rect 2006 967 2012 968
rect 1902 966 1908 967
rect 1870 963 1876 964
rect 1562 959 1568 960
rect 1562 955 1563 959
rect 1567 955 1568 959
rect 1562 954 1568 955
rect 1706 959 1712 960
rect 1706 955 1707 959
rect 1711 955 1712 959
rect 1706 954 1712 955
rect 1850 959 1856 960
rect 1850 955 1851 959
rect 1855 955 1856 959
rect 1870 959 1871 963
rect 1875 959 1876 963
rect 2048 961 2050 981
rect 1870 958 1876 959
rect 2046 960 2052 961
rect 2648 960 2650 981
rect 2744 960 2746 981
rect 2848 960 2850 981
rect 1850 954 1856 955
rect 1564 932 1566 954
rect 1630 952 1636 953
rect 1630 948 1631 952
rect 1635 948 1636 952
rect 1630 947 1636 948
rect 1554 931 1560 932
rect 1554 927 1555 931
rect 1559 927 1560 931
rect 1554 926 1560 927
rect 1562 931 1568 932
rect 1562 927 1563 931
rect 1567 927 1568 931
rect 1562 926 1568 927
rect 1632 923 1634 947
rect 1708 932 1710 954
rect 1774 952 1780 953
rect 1774 948 1775 952
rect 1779 948 1780 952
rect 1774 947 1780 948
rect 1706 931 1712 932
rect 1706 927 1707 931
rect 1711 927 1712 931
rect 1706 926 1712 927
rect 1776 923 1778 947
rect 1852 932 1854 954
rect 1850 931 1856 932
rect 1850 927 1851 931
rect 1855 927 1856 931
rect 1850 926 1856 927
rect 1872 924 1874 958
rect 2046 956 2047 960
rect 2051 956 2052 960
rect 2006 955 2012 956
rect 2046 955 2052 956
rect 2646 959 2652 960
rect 2646 955 2647 959
rect 2651 955 2652 959
rect 1902 952 1908 953
rect 1902 948 1903 952
rect 1907 948 1908 952
rect 2006 951 2007 955
rect 2011 951 2012 955
rect 2646 954 2652 955
rect 2742 959 2748 960
rect 2742 955 2743 959
rect 2747 955 2748 959
rect 2742 954 2748 955
rect 2846 959 2852 960
rect 2846 955 2847 959
rect 2851 955 2852 959
rect 2846 954 2852 955
rect 2924 952 2926 1050
rect 3008 1033 3010 1057
rect 3190 1055 3196 1056
rect 3190 1051 3191 1055
rect 3195 1051 3196 1055
rect 3190 1050 3196 1051
rect 3006 1032 3012 1033
rect 3006 1028 3007 1032
rect 3011 1028 3012 1032
rect 3192 1029 3194 1050
rect 3200 1033 3202 1057
rect 3228 1056 3230 1098
rect 3260 1084 3262 1102
rect 3318 1096 3324 1097
rect 3318 1092 3319 1096
rect 3323 1092 3324 1096
rect 3318 1091 3324 1092
rect 3258 1083 3264 1084
rect 3258 1079 3259 1083
rect 3263 1079 3264 1083
rect 3258 1078 3264 1079
rect 3320 1063 3322 1091
rect 3476 1076 3478 1182
rect 3550 1177 3556 1178
rect 3550 1173 3551 1177
rect 3555 1173 3556 1177
rect 3550 1172 3556 1173
rect 3702 1177 3708 1178
rect 3702 1173 3703 1177
rect 3707 1173 3708 1177
rect 3702 1172 3708 1173
rect 3838 1177 3844 1178
rect 3838 1173 3839 1177
rect 3843 1173 3844 1177
rect 3838 1172 3844 1173
rect 3552 1143 3554 1172
rect 3704 1143 3706 1172
rect 3840 1143 3842 1172
rect 3495 1142 3499 1143
rect 3495 1137 3499 1138
rect 3551 1142 3555 1143
rect 3551 1137 3555 1138
rect 3679 1142 3683 1143
rect 3679 1137 3683 1138
rect 3703 1142 3707 1143
rect 3703 1137 3707 1138
rect 3839 1142 3843 1143
rect 3839 1137 3843 1138
rect 3496 1116 3498 1137
rect 3680 1116 3682 1137
rect 3840 1116 3842 1137
rect 3494 1115 3500 1116
rect 3494 1111 3495 1115
rect 3499 1111 3500 1115
rect 3494 1110 3500 1111
rect 3678 1115 3684 1116
rect 3678 1111 3679 1115
rect 3683 1111 3684 1115
rect 3678 1110 3684 1111
rect 3838 1115 3844 1116
rect 3838 1111 3839 1115
rect 3843 1111 3844 1115
rect 3838 1110 3844 1111
rect 3916 1108 3918 1214
rect 3944 1194 3946 1221
rect 3942 1193 3948 1194
rect 3942 1189 3943 1193
rect 3947 1189 3948 1193
rect 3942 1188 3948 1189
rect 3942 1176 3948 1177
rect 3942 1172 3943 1176
rect 3947 1172 3948 1176
rect 3942 1171 3948 1172
rect 3944 1143 3946 1171
rect 3943 1142 3947 1143
rect 3943 1137 3947 1138
rect 3944 1117 3946 1137
rect 3942 1116 3948 1117
rect 3942 1112 3943 1116
rect 3947 1112 3948 1116
rect 3942 1111 3948 1112
rect 3578 1107 3584 1108
rect 3570 1103 3576 1104
rect 3570 1099 3571 1103
rect 3575 1099 3576 1103
rect 3578 1103 3579 1107
rect 3583 1103 3584 1107
rect 3578 1102 3584 1103
rect 3914 1107 3920 1108
rect 3914 1103 3915 1107
rect 3919 1103 3920 1107
rect 3914 1102 3920 1103
rect 3570 1098 3576 1099
rect 3494 1096 3500 1097
rect 3494 1092 3495 1096
rect 3499 1092 3500 1096
rect 3494 1091 3500 1092
rect 3474 1075 3480 1076
rect 3474 1071 3475 1075
rect 3479 1071 3480 1075
rect 3474 1070 3480 1071
rect 3496 1063 3498 1091
rect 3572 1076 3574 1098
rect 3580 1084 3582 1102
rect 3942 1099 3948 1100
rect 3678 1096 3684 1097
rect 3678 1092 3679 1096
rect 3683 1092 3684 1096
rect 3678 1091 3684 1092
rect 3838 1096 3844 1097
rect 3838 1092 3839 1096
rect 3843 1092 3844 1096
rect 3942 1095 3943 1099
rect 3947 1095 3948 1099
rect 3942 1094 3948 1095
rect 3838 1091 3844 1092
rect 3578 1083 3584 1084
rect 3578 1079 3579 1083
rect 3583 1079 3584 1083
rect 3578 1078 3584 1079
rect 3570 1075 3576 1076
rect 3570 1071 3571 1075
rect 3575 1071 3576 1075
rect 3570 1070 3576 1071
rect 3680 1063 3682 1091
rect 3840 1063 3842 1091
rect 3906 1071 3912 1072
rect 3906 1067 3907 1071
rect 3911 1067 3912 1071
rect 3906 1066 3912 1067
rect 3319 1062 3323 1063
rect 3319 1057 3323 1058
rect 3407 1062 3411 1063
rect 3407 1057 3411 1058
rect 3495 1062 3499 1063
rect 3495 1057 3499 1058
rect 3631 1062 3635 1063
rect 3631 1057 3635 1058
rect 3679 1062 3683 1063
rect 3679 1057 3683 1058
rect 3839 1062 3843 1063
rect 3839 1057 3843 1058
rect 3226 1055 3232 1056
rect 3226 1051 3227 1055
rect 3231 1051 3232 1055
rect 3226 1050 3232 1051
rect 3274 1055 3280 1056
rect 3274 1051 3275 1055
rect 3279 1051 3280 1055
rect 3274 1050 3280 1051
rect 3198 1032 3204 1033
rect 3006 1027 3012 1028
rect 3191 1028 3195 1029
rect 3198 1028 3199 1032
rect 3203 1028 3204 1032
rect 3198 1027 3204 1028
rect 3276 1024 3278 1050
rect 3408 1033 3410 1057
rect 3482 1055 3488 1056
rect 3482 1051 3483 1055
rect 3487 1051 3488 1055
rect 3482 1050 3488 1051
rect 3406 1032 3412 1033
rect 3406 1028 3407 1032
rect 3411 1028 3412 1032
rect 3406 1027 3412 1028
rect 3484 1024 3486 1050
rect 3632 1033 3634 1057
rect 3840 1033 3842 1057
rect 3630 1032 3636 1033
rect 3559 1028 3563 1029
rect 3630 1028 3631 1032
rect 3635 1028 3636 1032
rect 3630 1027 3636 1028
rect 3838 1032 3844 1033
rect 3838 1028 3839 1032
rect 3843 1028 3844 1032
rect 3838 1027 3844 1028
rect 3908 1024 3910 1066
rect 3944 1063 3946 1094
rect 3943 1062 3947 1063
rect 3943 1057 3947 1058
rect 3914 1055 3920 1056
rect 3914 1051 3915 1055
rect 3919 1051 3920 1055
rect 3914 1050 3920 1051
rect 3074 1023 3080 1024
rect 3191 1023 3195 1024
rect 3274 1023 3280 1024
rect 3074 1019 3075 1023
rect 3079 1019 3080 1023
rect 3074 1018 3080 1019
rect 3274 1019 3275 1023
rect 3279 1019 3280 1023
rect 3274 1018 3280 1019
rect 3482 1023 3488 1024
rect 3482 1019 3483 1023
rect 3487 1019 3488 1023
rect 3482 1018 3488 1019
rect 3558 1023 3564 1024
rect 3558 1019 3559 1023
rect 3563 1019 3564 1023
rect 3558 1018 3564 1019
rect 3906 1023 3912 1024
rect 3906 1019 3907 1023
rect 3911 1019 3912 1023
rect 3906 1018 3912 1019
rect 3006 1013 3012 1014
rect 3006 1009 3007 1013
rect 3011 1009 3012 1013
rect 3006 1008 3012 1009
rect 3008 987 3010 1008
rect 2967 986 2971 987
rect 2967 981 2971 982
rect 3007 986 3011 987
rect 3007 981 3011 982
rect 2968 960 2970 981
rect 2966 959 2972 960
rect 2966 955 2967 959
rect 2971 955 2972 959
rect 2966 954 2972 955
rect 2006 950 2012 951
rect 2922 951 2928 952
rect 1902 947 1908 948
rect 1870 923 1876 924
rect 1904 923 1906 947
rect 2008 923 2010 950
rect 2722 947 2728 948
rect 2046 943 2052 944
rect 2046 939 2047 943
rect 2051 939 2052 943
rect 2722 943 2723 947
rect 2727 943 2728 947
rect 2722 942 2728 943
rect 2818 947 2824 948
rect 2818 943 2819 947
rect 2823 943 2824 947
rect 2922 947 2923 951
rect 2927 947 2928 951
rect 2922 946 2928 947
rect 2818 942 2824 943
rect 2046 938 2052 939
rect 2646 940 2652 941
rect 1175 922 1179 923
rect 1230 922 1236 923
rect 1239 922 1243 923
rect 1175 917 1179 918
rect 1082 915 1088 916
rect 1082 911 1083 915
rect 1087 911 1088 915
rect 1082 910 1088 911
rect 1054 892 1060 893
rect 1054 888 1055 892
rect 1059 888 1060 892
rect 1054 887 1060 888
rect 1232 884 1234 922
rect 1239 917 1243 918
rect 1335 922 1339 923
rect 1335 917 1339 918
rect 1415 922 1419 923
rect 1415 917 1419 918
rect 1487 922 1491 923
rect 1487 917 1491 918
rect 1583 922 1587 923
rect 1583 917 1587 918
rect 1631 922 1635 923
rect 1631 917 1635 918
rect 1751 922 1755 923
rect 1751 917 1755 918
rect 1775 922 1779 923
rect 1870 919 1871 923
rect 1875 919 1876 923
rect 1870 918 1876 919
rect 1903 922 1907 923
rect 1775 917 1779 918
rect 1903 917 1907 918
rect 2007 922 2011 923
rect 2007 917 2011 918
rect 1240 893 1242 917
rect 1322 915 1328 916
rect 1322 911 1323 915
rect 1327 911 1328 915
rect 1322 910 1328 911
rect 1238 892 1244 893
rect 1238 888 1239 892
rect 1243 888 1244 892
rect 1238 887 1244 888
rect 1324 884 1326 910
rect 1416 893 1418 917
rect 1498 915 1504 916
rect 1498 911 1499 915
rect 1503 911 1504 915
rect 1498 910 1504 911
rect 1414 892 1420 893
rect 1414 888 1415 892
rect 1419 888 1420 892
rect 1414 887 1420 888
rect 1500 884 1502 910
rect 1584 893 1586 917
rect 1610 915 1616 916
rect 1610 911 1611 915
rect 1615 911 1616 915
rect 1610 910 1616 911
rect 1582 892 1588 893
rect 1582 888 1583 892
rect 1587 888 1588 892
rect 1582 887 1588 888
rect 210 883 216 884
rect 210 879 211 883
rect 215 879 216 883
rect 210 878 216 879
rect 346 883 352 884
rect 346 879 347 883
rect 351 879 352 883
rect 346 878 352 879
rect 530 883 536 884
rect 530 879 531 883
rect 535 879 536 883
rect 530 878 536 879
rect 730 883 736 884
rect 730 879 731 883
rect 735 879 736 883
rect 730 878 736 879
rect 922 883 928 884
rect 922 879 923 883
rect 927 879 928 883
rect 922 878 928 879
rect 1166 883 1172 884
rect 1166 879 1167 883
rect 1171 879 1172 883
rect 1166 878 1172 879
rect 1230 883 1236 884
rect 1230 879 1231 883
rect 1235 879 1236 883
rect 1230 878 1236 879
rect 1322 883 1328 884
rect 1322 879 1323 883
rect 1327 879 1328 883
rect 1322 878 1328 879
rect 1498 883 1504 884
rect 1498 879 1499 883
rect 1503 879 1504 883
rect 1498 878 1504 879
rect 270 873 276 874
rect 270 869 271 873
rect 275 869 276 873
rect 270 868 276 869
rect 454 873 460 874
rect 454 869 455 873
rect 459 869 460 873
rect 454 868 460 869
rect 654 873 660 874
rect 654 869 655 873
rect 659 869 660 873
rect 654 868 660 869
rect 854 873 860 874
rect 854 869 855 873
rect 859 869 860 873
rect 854 868 860 869
rect 1054 873 1060 874
rect 1054 869 1055 873
rect 1059 869 1060 873
rect 1054 868 1060 869
rect 272 847 274 868
rect 456 847 458 868
rect 656 847 658 868
rect 856 847 858 868
rect 1056 847 1058 868
rect 215 846 219 847
rect 215 841 219 842
rect 271 846 275 847
rect 271 841 275 842
rect 343 846 347 847
rect 343 841 347 842
rect 455 846 459 847
rect 455 841 459 842
rect 495 846 499 847
rect 495 841 499 842
rect 655 846 659 847
rect 655 841 659 842
rect 831 846 835 847
rect 831 841 835 842
rect 855 846 859 847
rect 855 841 859 842
rect 1007 846 1011 847
rect 1007 841 1011 842
rect 1055 846 1059 847
rect 1055 841 1059 842
rect 216 820 218 841
rect 344 820 346 841
rect 496 820 498 841
rect 656 820 658 841
rect 832 820 834 841
rect 1008 820 1010 841
rect 214 819 220 820
rect 214 815 215 819
rect 219 815 220 819
rect 214 814 220 815
rect 342 819 348 820
rect 342 815 343 819
rect 347 815 348 819
rect 342 814 348 815
rect 494 819 500 820
rect 494 815 495 819
rect 499 815 500 819
rect 494 814 500 815
rect 654 819 660 820
rect 654 815 655 819
rect 659 815 660 819
rect 654 814 660 815
rect 830 819 836 820
rect 830 815 831 819
rect 835 815 836 819
rect 830 814 836 815
rect 1006 819 1012 820
rect 1006 815 1007 819
rect 1011 815 1012 819
rect 1006 814 1012 815
rect 190 811 196 812
rect 190 807 191 811
rect 195 807 196 811
rect 190 806 196 807
rect 330 811 336 812
rect 330 807 331 811
rect 335 807 336 811
rect 330 806 336 807
rect 614 811 620 812
rect 614 807 615 811
rect 619 807 620 811
rect 1094 811 1100 812
rect 614 806 620 807
rect 1082 807 1088 808
rect 110 803 116 804
rect 110 799 111 803
rect 115 799 116 803
rect 110 798 116 799
rect 214 800 220 801
rect 112 771 114 798
rect 214 796 215 800
rect 219 796 220 800
rect 214 795 220 796
rect 216 771 218 795
rect 332 780 334 806
rect 342 800 348 801
rect 342 796 343 800
rect 347 796 348 800
rect 342 795 348 796
rect 494 800 500 801
rect 494 796 495 800
rect 499 796 500 800
rect 494 795 500 796
rect 330 779 336 780
rect 330 775 331 779
rect 335 775 336 779
rect 330 774 336 775
rect 344 771 346 795
rect 496 771 498 795
rect 616 780 618 806
rect 1082 803 1083 807
rect 1087 803 1088 807
rect 1094 807 1095 811
rect 1099 807 1100 811
rect 1094 806 1100 807
rect 1082 802 1088 803
rect 654 800 660 801
rect 654 796 655 800
rect 659 796 660 800
rect 654 795 660 796
rect 830 800 836 801
rect 830 796 831 800
rect 835 796 836 800
rect 830 795 836 796
rect 1006 800 1012 801
rect 1006 796 1007 800
rect 1011 796 1012 800
rect 1006 795 1012 796
rect 614 779 620 780
rect 614 775 615 779
rect 619 775 620 779
rect 614 774 620 775
rect 656 771 658 795
rect 832 771 834 795
rect 878 775 884 776
rect 878 771 879 775
rect 883 771 884 775
rect 1008 771 1010 795
rect 111 770 115 771
rect 111 765 115 766
rect 215 770 219 771
rect 215 765 219 766
rect 343 770 347 771
rect 343 765 347 766
rect 375 770 379 771
rect 375 765 379 766
rect 495 770 499 771
rect 495 765 499 766
rect 623 770 627 771
rect 623 765 627 766
rect 655 770 659 771
rect 655 765 659 766
rect 751 770 755 771
rect 751 765 755 766
rect 831 770 835 771
rect 878 770 884 771
rect 887 770 891 771
rect 831 765 835 766
rect 112 738 114 765
rect 376 741 378 765
rect 450 763 456 764
rect 450 759 451 763
rect 455 759 456 763
rect 450 758 456 759
rect 374 740 380 741
rect 110 737 116 738
rect 110 733 111 737
rect 115 733 116 737
rect 374 736 375 740
rect 379 736 380 740
rect 374 735 380 736
rect 110 732 116 733
rect 452 732 454 758
rect 496 741 498 765
rect 570 763 576 764
rect 570 759 571 763
rect 575 759 576 763
rect 570 758 576 759
rect 494 740 500 741
rect 494 736 495 740
rect 499 736 500 740
rect 494 735 500 736
rect 572 732 574 758
rect 624 741 626 765
rect 698 755 704 756
rect 698 751 699 755
rect 703 751 704 755
rect 698 750 704 751
rect 622 740 628 741
rect 622 736 623 740
rect 627 736 628 740
rect 622 735 628 736
rect 700 732 702 750
rect 752 741 754 765
rect 818 763 824 764
rect 818 759 819 763
rect 823 759 824 763
rect 818 758 824 759
rect 750 740 756 741
rect 750 736 751 740
rect 755 736 756 740
rect 750 735 756 736
rect 450 731 456 732
rect 450 727 451 731
rect 455 727 456 731
rect 450 726 456 727
rect 570 731 576 732
rect 570 727 571 731
rect 575 727 576 731
rect 570 726 576 727
rect 698 731 704 732
rect 698 727 699 731
rect 703 727 704 731
rect 698 726 704 727
rect 374 721 380 722
rect 110 720 116 721
rect 110 716 111 720
rect 115 716 116 720
rect 374 717 375 721
rect 379 717 380 721
rect 374 716 380 717
rect 494 721 500 722
rect 494 717 495 721
rect 499 717 500 721
rect 494 716 500 717
rect 622 721 628 722
rect 622 717 623 721
rect 627 717 628 721
rect 622 716 628 717
rect 750 721 756 722
rect 750 717 751 721
rect 755 717 756 721
rect 750 716 756 717
rect 110 715 116 716
rect 112 695 114 715
rect 376 695 378 716
rect 496 695 498 716
rect 624 695 626 716
rect 752 695 754 716
rect 111 694 115 695
rect 111 689 115 690
rect 375 694 379 695
rect 375 689 379 690
rect 495 694 499 695
rect 495 689 499 690
rect 527 694 531 695
rect 527 689 531 690
rect 623 694 627 695
rect 623 689 627 690
rect 631 694 635 695
rect 631 689 635 690
rect 743 694 747 695
rect 743 689 747 690
rect 751 694 755 695
rect 751 689 755 690
rect 112 669 114 689
rect 110 668 116 669
rect 528 668 530 689
rect 632 668 634 689
rect 744 668 746 689
rect 110 664 111 668
rect 115 664 116 668
rect 110 663 116 664
rect 526 667 532 668
rect 526 663 527 667
rect 531 663 532 667
rect 526 662 532 663
rect 630 667 636 668
rect 630 663 631 667
rect 635 663 636 667
rect 630 662 636 663
rect 742 667 748 668
rect 742 663 743 667
rect 747 663 748 667
rect 742 662 748 663
rect 820 660 822 758
rect 880 732 882 770
rect 887 765 891 766
rect 1007 770 1011 771
rect 1007 765 1011 766
rect 1023 770 1027 771
rect 1023 765 1027 766
rect 888 741 890 765
rect 1024 741 1026 765
rect 1084 764 1086 802
rect 1096 780 1098 806
rect 1168 780 1170 878
rect 1238 873 1244 874
rect 1238 869 1239 873
rect 1243 869 1244 873
rect 1238 868 1244 869
rect 1414 873 1420 874
rect 1414 869 1415 873
rect 1419 869 1420 873
rect 1414 868 1420 869
rect 1582 873 1588 874
rect 1582 869 1583 873
rect 1587 869 1588 873
rect 1582 868 1588 869
rect 1240 847 1242 868
rect 1416 847 1418 868
rect 1584 847 1586 868
rect 1183 846 1187 847
rect 1183 841 1187 842
rect 1239 846 1243 847
rect 1239 841 1243 842
rect 1359 846 1363 847
rect 1359 841 1363 842
rect 1415 846 1419 847
rect 1415 841 1419 842
rect 1535 846 1539 847
rect 1535 841 1539 842
rect 1583 846 1587 847
rect 1583 841 1587 842
rect 1184 820 1186 841
rect 1360 820 1362 841
rect 1536 820 1538 841
rect 1182 819 1188 820
rect 1182 815 1183 819
rect 1187 815 1188 819
rect 1182 814 1188 815
rect 1358 819 1364 820
rect 1358 815 1359 819
rect 1363 815 1364 819
rect 1358 814 1364 815
rect 1534 819 1540 820
rect 1534 815 1535 819
rect 1539 815 1540 819
rect 1534 814 1540 815
rect 1612 812 1614 910
rect 1752 893 1754 917
rect 1826 915 1832 916
rect 1826 911 1827 915
rect 1831 911 1832 915
rect 1826 910 1832 911
rect 1750 892 1756 893
rect 1750 888 1751 892
rect 1755 888 1756 892
rect 1750 887 1756 888
rect 1828 884 1830 910
rect 1904 893 1906 917
rect 1902 892 1908 893
rect 1902 888 1903 892
rect 1907 888 1908 892
rect 2008 890 2010 917
rect 2048 899 2050 938
rect 2646 936 2647 940
rect 2651 936 2652 940
rect 2646 935 2652 936
rect 2648 899 2650 935
rect 2724 924 2726 942
rect 2742 940 2748 941
rect 2742 936 2743 940
rect 2747 936 2748 940
rect 2742 935 2748 936
rect 2722 923 2728 924
rect 2722 919 2723 923
rect 2727 919 2728 923
rect 2722 918 2728 919
rect 2744 899 2746 935
rect 2820 920 2822 942
rect 2846 940 2852 941
rect 2846 936 2847 940
rect 2851 936 2852 940
rect 2846 935 2852 936
rect 2966 940 2972 941
rect 2966 936 2967 940
rect 2971 936 2972 940
rect 2966 935 2972 936
rect 2818 919 2824 920
rect 2750 915 2756 916
rect 2750 911 2751 915
rect 2755 911 2756 915
rect 2818 915 2819 919
rect 2823 915 2824 919
rect 2818 914 2824 915
rect 2750 910 2756 911
rect 2047 898 2051 899
rect 2047 893 2051 894
rect 2071 898 2075 899
rect 2071 893 2075 894
rect 2255 898 2259 899
rect 2255 893 2259 894
rect 2463 898 2467 899
rect 2463 893 2467 894
rect 2647 898 2651 899
rect 2647 893 2651 894
rect 2679 898 2683 899
rect 2679 893 2683 894
rect 2743 898 2747 899
rect 2743 893 2747 894
rect 1902 887 1908 888
rect 2006 889 2012 890
rect 2006 885 2007 889
rect 2011 885 2012 889
rect 2006 884 2012 885
rect 1826 883 1832 884
rect 1826 879 1827 883
rect 1831 879 1832 883
rect 1826 878 1832 879
rect 1750 873 1756 874
rect 1750 869 1751 873
rect 1755 869 1756 873
rect 1750 868 1756 869
rect 1902 873 1908 874
rect 1902 869 1903 873
rect 1907 869 1908 873
rect 1902 868 1908 869
rect 2006 872 2012 873
rect 2006 868 2007 872
rect 2011 868 2012 872
rect 1752 847 1754 868
rect 1904 847 1906 868
rect 2006 867 2012 868
rect 2008 847 2010 867
rect 2048 866 2050 893
rect 2072 869 2074 893
rect 2146 891 2152 892
rect 2146 887 2147 891
rect 2151 887 2152 891
rect 2146 886 2152 887
rect 2070 868 2076 869
rect 2046 865 2052 866
rect 2046 861 2047 865
rect 2051 861 2052 865
rect 2070 864 2071 868
rect 2075 864 2076 868
rect 2070 863 2076 864
rect 2046 860 2052 861
rect 2148 860 2150 886
rect 2256 869 2258 893
rect 2330 891 2336 892
rect 2330 887 2331 891
rect 2335 887 2336 891
rect 2330 886 2336 887
rect 2254 868 2260 869
rect 2254 864 2255 868
rect 2259 864 2260 868
rect 2254 863 2260 864
rect 2332 860 2334 886
rect 2464 869 2466 893
rect 2680 869 2682 893
rect 2462 868 2468 869
rect 2462 864 2463 868
rect 2467 864 2468 868
rect 2462 863 2468 864
rect 2678 868 2684 869
rect 2678 864 2679 868
rect 2683 864 2684 868
rect 2678 863 2684 864
rect 2752 860 2754 910
rect 2848 899 2850 935
rect 2968 899 2970 935
rect 3076 920 3078 1018
rect 3198 1013 3204 1014
rect 3198 1009 3199 1013
rect 3203 1009 3204 1013
rect 3198 1008 3204 1009
rect 3406 1013 3412 1014
rect 3406 1009 3407 1013
rect 3411 1009 3412 1013
rect 3406 1008 3412 1009
rect 3630 1013 3636 1014
rect 3630 1009 3631 1013
rect 3635 1009 3636 1013
rect 3630 1008 3636 1009
rect 3838 1013 3844 1014
rect 3838 1009 3839 1013
rect 3843 1009 3844 1013
rect 3838 1008 3844 1009
rect 3200 987 3202 1008
rect 3408 987 3410 1008
rect 3632 987 3634 1008
rect 3840 987 3842 1008
rect 3111 986 3115 987
rect 3111 981 3115 982
rect 3199 986 3203 987
rect 3199 981 3203 982
rect 3279 986 3283 987
rect 3279 981 3283 982
rect 3407 986 3411 987
rect 3407 981 3411 982
rect 3463 986 3467 987
rect 3463 981 3467 982
rect 3631 986 3635 987
rect 3631 981 3635 982
rect 3663 986 3667 987
rect 3663 981 3667 982
rect 3839 986 3843 987
rect 3839 981 3843 982
rect 3112 960 3114 981
rect 3280 960 3282 981
rect 3464 960 3466 981
rect 3664 960 3666 981
rect 3840 960 3842 981
rect 3110 959 3116 960
rect 3110 955 3111 959
rect 3115 955 3116 959
rect 3110 954 3116 955
rect 3278 959 3284 960
rect 3278 955 3279 959
rect 3283 955 3284 959
rect 3278 954 3284 955
rect 3462 959 3468 960
rect 3462 955 3463 959
rect 3467 955 3468 959
rect 3462 954 3468 955
rect 3662 959 3668 960
rect 3662 955 3663 959
rect 3667 955 3668 959
rect 3662 954 3668 955
rect 3838 959 3844 960
rect 3838 955 3839 959
rect 3843 955 3844 959
rect 3838 954 3844 955
rect 3916 952 3918 1050
rect 3944 1030 3946 1057
rect 3942 1029 3948 1030
rect 3942 1025 3943 1029
rect 3947 1025 3948 1029
rect 3942 1024 3948 1025
rect 3942 1012 3948 1013
rect 3942 1008 3943 1012
rect 3947 1008 3948 1012
rect 3942 1007 3948 1008
rect 3944 987 3946 1007
rect 3943 986 3947 987
rect 3943 981 3947 982
rect 3944 961 3946 981
rect 3942 960 3948 961
rect 3942 956 3943 960
rect 3947 956 3948 960
rect 3942 955 3948 956
rect 3622 951 3628 952
rect 3086 947 3092 948
rect 3086 943 3087 947
rect 3091 943 3092 947
rect 3086 942 3092 943
rect 3186 947 3192 948
rect 3186 943 3187 947
rect 3191 943 3192 947
rect 3186 942 3192 943
rect 3354 947 3360 948
rect 3354 943 3355 947
rect 3359 943 3360 947
rect 3354 942 3360 943
rect 3538 947 3544 948
rect 3538 943 3539 947
rect 3543 943 3544 947
rect 3622 947 3623 951
rect 3627 947 3628 951
rect 3622 946 3628 947
rect 3914 951 3920 952
rect 3914 947 3915 951
rect 3919 947 3920 951
rect 3914 946 3920 947
rect 3538 942 3544 943
rect 3088 920 3090 942
rect 3110 940 3116 941
rect 3110 936 3111 940
rect 3115 936 3116 940
rect 3110 935 3116 936
rect 3074 919 3080 920
rect 3074 915 3075 919
rect 3079 915 3080 919
rect 3074 914 3080 915
rect 3086 919 3092 920
rect 3086 915 3087 919
rect 3091 915 3092 919
rect 3086 914 3092 915
rect 3112 899 3114 935
rect 3188 920 3190 942
rect 3278 940 3284 941
rect 3278 936 3279 940
rect 3283 936 3284 940
rect 3278 935 3284 936
rect 3186 919 3192 920
rect 3186 915 3187 919
rect 3191 915 3192 919
rect 3186 914 3192 915
rect 3280 899 3282 935
rect 3356 920 3358 942
rect 3462 940 3468 941
rect 3462 936 3463 940
rect 3467 936 3468 940
rect 3462 935 3468 936
rect 3354 919 3360 920
rect 3354 915 3355 919
rect 3359 915 3360 919
rect 3354 914 3360 915
rect 3464 899 3466 935
rect 3540 920 3542 942
rect 3538 919 3544 920
rect 3538 915 3539 919
rect 3543 915 3544 919
rect 3538 914 3544 915
rect 3624 900 3626 946
rect 3942 943 3948 944
rect 3662 940 3668 941
rect 3662 936 3663 940
rect 3667 936 3668 940
rect 3662 935 3668 936
rect 3838 940 3844 941
rect 3838 936 3839 940
rect 3843 936 3844 940
rect 3942 939 3943 943
rect 3947 939 3948 943
rect 3942 938 3948 939
rect 3838 935 3844 936
rect 3622 899 3628 900
rect 3664 899 3666 935
rect 3840 899 3842 935
rect 3906 915 3912 916
rect 3906 911 3907 915
rect 3911 911 3912 915
rect 3906 910 3912 911
rect 2847 898 2851 899
rect 2847 893 2851 894
rect 2895 898 2899 899
rect 2895 893 2899 894
rect 2967 898 2971 899
rect 2967 893 2971 894
rect 3111 898 3115 899
rect 3111 893 3115 894
rect 3127 898 3131 899
rect 3127 893 3131 894
rect 3279 898 3283 899
rect 3279 893 3283 894
rect 3367 898 3371 899
rect 3367 893 3371 894
rect 3463 898 3467 899
rect 3463 893 3467 894
rect 3615 898 3619 899
rect 3622 895 3623 899
rect 3627 895 3628 899
rect 3622 894 3628 895
rect 3663 898 3667 899
rect 3615 893 3619 894
rect 3663 893 3667 894
rect 3839 898 3843 899
rect 3839 893 3843 894
rect 2896 869 2898 893
rect 2970 887 2976 888
rect 2970 883 2971 887
rect 2975 883 2976 887
rect 2970 882 2976 883
rect 2894 868 2900 869
rect 2894 864 2895 868
rect 2899 864 2900 868
rect 2894 863 2900 864
rect 2146 859 2152 860
rect 2146 855 2147 859
rect 2151 855 2152 859
rect 2146 854 2152 855
rect 2330 859 2336 860
rect 2330 855 2331 859
rect 2335 855 2336 859
rect 2330 854 2336 855
rect 2350 859 2356 860
rect 2350 855 2351 859
rect 2355 855 2356 859
rect 2350 854 2356 855
rect 2750 859 2756 860
rect 2750 855 2751 859
rect 2755 855 2756 859
rect 2750 854 2756 855
rect 2070 849 2076 850
rect 2046 848 2052 849
rect 1719 846 1723 847
rect 1719 841 1723 842
rect 1751 846 1755 847
rect 1751 841 1755 842
rect 1903 846 1907 847
rect 1903 841 1907 842
rect 2007 846 2011 847
rect 2046 844 2047 848
rect 2051 844 2052 848
rect 2070 845 2071 849
rect 2075 845 2076 849
rect 2070 844 2076 845
rect 2254 849 2260 850
rect 2254 845 2255 849
rect 2259 845 2260 849
rect 2254 844 2260 845
rect 2046 843 2052 844
rect 2007 841 2011 842
rect 1720 820 1722 841
rect 2008 821 2010 841
rect 2048 823 2050 843
rect 2072 823 2074 844
rect 2256 823 2258 844
rect 2047 822 2051 823
rect 2006 820 2012 821
rect 1718 819 1724 820
rect 1718 815 1719 819
rect 1723 815 1724 819
rect 2006 816 2007 820
rect 2011 816 2012 820
rect 2047 817 2051 818
rect 2071 822 2075 823
rect 2071 817 2075 818
rect 2215 822 2219 823
rect 2215 817 2219 818
rect 2255 822 2259 823
rect 2255 817 2259 818
rect 2327 822 2331 823
rect 2327 817 2331 818
rect 2006 815 2012 816
rect 1718 814 1724 815
rect 1610 811 1616 812
rect 1462 807 1468 808
rect 1462 803 1463 807
rect 1467 803 1468 807
rect 1610 807 1611 811
rect 1615 807 1616 811
rect 1610 806 1616 807
rect 1638 811 1644 812
rect 1638 807 1639 811
rect 1643 807 1644 811
rect 1638 806 1644 807
rect 1462 802 1468 803
rect 1182 800 1188 801
rect 1182 796 1183 800
rect 1187 796 1188 800
rect 1182 795 1188 796
rect 1358 800 1364 801
rect 1358 796 1359 800
rect 1363 796 1364 800
rect 1358 795 1364 796
rect 1094 779 1100 780
rect 1094 775 1095 779
rect 1099 775 1100 779
rect 1094 774 1100 775
rect 1166 779 1172 780
rect 1166 775 1167 779
rect 1171 775 1172 779
rect 1166 774 1172 775
rect 1184 771 1186 795
rect 1360 771 1362 795
rect 1464 776 1466 802
rect 1534 800 1540 801
rect 1534 796 1535 800
rect 1539 796 1540 800
rect 1534 795 1540 796
rect 1462 775 1468 776
rect 1462 771 1463 775
rect 1467 771 1468 775
rect 1536 771 1538 795
rect 1640 788 1642 806
rect 2006 803 2012 804
rect 1718 800 1724 801
rect 1718 796 1719 800
rect 1723 796 1724 800
rect 2006 799 2007 803
rect 2011 799 2012 803
rect 2006 798 2012 799
rect 1718 795 1724 796
rect 1638 787 1644 788
rect 1638 783 1639 787
rect 1643 783 1644 787
rect 1638 782 1644 783
rect 1674 775 1680 776
rect 1674 771 1675 775
rect 1679 771 1680 775
rect 1720 771 1722 795
rect 2008 771 2010 798
rect 2048 797 2050 817
rect 2046 796 2052 797
rect 2216 796 2218 817
rect 2328 796 2330 817
rect 2046 792 2047 796
rect 2051 792 2052 796
rect 2046 791 2052 792
rect 2214 795 2220 796
rect 2214 791 2215 795
rect 2219 791 2220 795
rect 2214 790 2220 791
rect 2326 795 2332 796
rect 2326 791 2327 795
rect 2331 791 2332 795
rect 2326 790 2332 791
rect 2290 783 2296 784
rect 2046 779 2052 780
rect 2046 775 2047 779
rect 2051 775 2052 779
rect 2290 779 2291 783
rect 2295 779 2296 783
rect 2290 778 2296 779
rect 2046 774 2052 775
rect 2214 776 2220 777
rect 1167 770 1171 771
rect 1167 765 1171 766
rect 1183 770 1187 771
rect 1183 765 1187 766
rect 1311 770 1315 771
rect 1311 765 1315 766
rect 1359 770 1363 771
rect 1359 765 1363 766
rect 1455 770 1459 771
rect 1462 770 1468 771
rect 1535 770 1539 771
rect 1455 765 1459 766
rect 1535 765 1539 766
rect 1599 770 1603 771
rect 1674 770 1680 771
rect 1719 770 1723 771
rect 1599 765 1603 766
rect 1078 763 1086 764
rect 1078 759 1079 763
rect 1083 760 1086 763
rect 1098 763 1104 764
rect 1083 759 1084 760
rect 1078 758 1084 759
rect 1098 759 1099 763
rect 1103 759 1104 763
rect 1098 758 1104 759
rect 886 740 892 741
rect 886 736 887 740
rect 891 736 892 740
rect 886 735 892 736
rect 1022 740 1028 741
rect 1022 736 1023 740
rect 1027 736 1028 740
rect 1022 735 1028 736
rect 1100 732 1102 758
rect 1168 741 1170 765
rect 1312 741 1314 765
rect 1366 763 1372 764
rect 1366 759 1367 763
rect 1371 759 1372 763
rect 1366 758 1372 759
rect 1386 763 1392 764
rect 1386 759 1387 763
rect 1391 759 1392 763
rect 1386 758 1392 759
rect 1166 740 1172 741
rect 1166 736 1167 740
rect 1171 736 1172 740
rect 1166 735 1172 736
rect 1310 740 1316 741
rect 1310 736 1311 740
rect 1315 736 1316 740
rect 1310 735 1316 736
rect 878 731 884 732
rect 878 727 879 731
rect 883 727 884 731
rect 878 726 884 727
rect 1098 731 1104 732
rect 1098 727 1099 731
rect 1103 727 1104 731
rect 1098 726 1104 727
rect 1234 731 1240 732
rect 1234 727 1235 731
rect 1239 727 1240 731
rect 1234 726 1240 727
rect 886 721 892 722
rect 886 717 887 721
rect 891 717 892 721
rect 886 716 892 717
rect 1022 721 1028 722
rect 1022 717 1023 721
rect 1027 717 1028 721
rect 1022 716 1028 717
rect 1166 721 1172 722
rect 1166 717 1167 721
rect 1171 717 1172 721
rect 1166 716 1172 717
rect 888 695 890 716
rect 1024 695 1026 716
rect 1168 695 1170 716
rect 855 694 859 695
rect 855 689 859 690
rect 887 694 891 695
rect 887 689 891 690
rect 967 694 971 695
rect 967 689 971 690
rect 1023 694 1027 695
rect 1023 689 1027 690
rect 1071 694 1075 695
rect 1071 689 1075 690
rect 1167 694 1171 695
rect 1167 689 1171 690
rect 1183 694 1187 695
rect 1183 689 1187 690
rect 856 668 858 689
rect 968 668 970 689
rect 1072 668 1074 689
rect 1184 668 1186 689
rect 854 667 860 668
rect 854 663 855 667
rect 859 663 860 667
rect 854 662 860 663
rect 966 667 972 668
rect 966 663 967 667
rect 971 663 972 667
rect 966 662 972 663
rect 1070 667 1076 668
rect 1070 663 1071 667
rect 1075 663 1076 667
rect 1070 662 1076 663
rect 1182 667 1188 668
rect 1182 663 1183 667
rect 1187 663 1188 667
rect 1182 662 1188 663
rect 818 659 824 660
rect 602 655 608 656
rect 110 651 116 652
rect 110 647 111 651
rect 115 647 116 651
rect 602 651 603 655
rect 607 651 608 655
rect 602 650 608 651
rect 706 655 712 656
rect 706 651 707 655
rect 711 651 712 655
rect 818 655 819 659
rect 823 655 824 659
rect 818 654 824 655
rect 826 659 832 660
rect 826 655 827 659
rect 831 655 832 659
rect 826 654 832 655
rect 1146 655 1152 656
rect 706 650 712 651
rect 110 646 116 647
rect 526 648 532 649
rect 112 619 114 646
rect 526 644 527 648
rect 531 644 532 648
rect 526 643 532 644
rect 528 619 530 643
rect 604 628 606 650
rect 630 648 636 649
rect 630 644 631 648
rect 635 644 636 648
rect 630 643 636 644
rect 602 627 608 628
rect 602 623 603 627
rect 607 623 608 627
rect 602 622 608 623
rect 632 619 634 643
rect 708 628 710 650
rect 742 648 748 649
rect 742 644 743 648
rect 747 644 748 648
rect 742 643 748 644
rect 706 627 712 628
rect 706 623 707 627
rect 711 623 712 627
rect 706 622 712 623
rect 744 619 746 643
rect 828 636 830 654
rect 1146 651 1147 655
rect 1151 651 1152 655
rect 1146 650 1152 651
rect 854 648 860 649
rect 854 644 855 648
rect 859 644 860 648
rect 854 643 860 644
rect 966 648 972 649
rect 966 644 967 648
rect 971 644 972 648
rect 966 643 972 644
rect 1070 648 1076 649
rect 1070 644 1071 648
rect 1075 644 1076 648
rect 1070 643 1076 644
rect 826 635 832 636
rect 826 631 827 635
rect 831 631 832 635
rect 826 630 832 631
rect 856 619 858 643
rect 968 619 970 643
rect 1072 619 1074 643
rect 111 618 115 619
rect 111 613 115 614
rect 527 618 531 619
rect 527 613 531 614
rect 631 618 635 619
rect 631 613 635 614
rect 687 618 691 619
rect 687 613 691 614
rect 743 618 747 619
rect 743 613 747 614
rect 783 618 787 619
rect 783 613 787 614
rect 855 618 859 619
rect 855 613 859 614
rect 879 618 883 619
rect 879 613 883 614
rect 967 618 971 619
rect 967 613 971 614
rect 975 618 979 619
rect 975 613 979 614
rect 1071 618 1075 619
rect 1071 613 1075 614
rect 112 586 114 613
rect 688 589 690 613
rect 762 611 768 612
rect 762 607 763 611
rect 767 607 768 611
rect 762 606 768 607
rect 686 588 692 589
rect 110 585 116 586
rect 110 581 111 585
rect 115 581 116 585
rect 686 584 687 588
rect 691 584 692 588
rect 686 583 692 584
rect 110 580 116 581
rect 764 580 766 606
rect 784 589 786 613
rect 880 589 882 613
rect 976 589 978 613
rect 1058 611 1064 612
rect 1058 607 1059 611
rect 1063 607 1064 611
rect 1058 606 1064 607
rect 1042 603 1048 604
rect 1042 599 1043 603
rect 1047 599 1048 603
rect 1042 598 1048 599
rect 782 588 788 589
rect 782 584 783 588
rect 787 584 788 588
rect 782 583 788 584
rect 878 588 884 589
rect 878 584 879 588
rect 883 584 884 588
rect 878 583 884 584
rect 974 588 980 589
rect 974 584 975 588
rect 979 584 980 588
rect 974 583 980 584
rect 1044 580 1046 598
rect 1060 580 1062 606
rect 1072 589 1074 613
rect 1148 612 1150 650
rect 1182 648 1188 649
rect 1182 644 1183 648
rect 1187 644 1188 648
rect 1182 643 1188 644
rect 1184 619 1186 643
rect 1236 628 1238 726
rect 1310 721 1316 722
rect 1310 717 1311 721
rect 1315 717 1316 721
rect 1310 716 1316 717
rect 1312 695 1314 716
rect 1295 694 1299 695
rect 1295 689 1299 690
rect 1311 694 1315 695
rect 1311 689 1315 690
rect 1296 668 1298 689
rect 1368 673 1370 758
rect 1388 732 1390 758
rect 1456 741 1458 765
rect 1600 741 1602 765
rect 1454 740 1460 741
rect 1454 736 1455 740
rect 1459 736 1460 740
rect 1454 735 1460 736
rect 1598 740 1604 741
rect 1598 736 1599 740
rect 1603 736 1604 740
rect 1598 735 1604 736
rect 1676 732 1678 770
rect 1719 765 1723 766
rect 2007 770 2011 771
rect 2007 765 2011 766
rect 2008 738 2010 765
rect 2048 743 2050 774
rect 2214 772 2215 776
rect 2219 772 2220 776
rect 2214 771 2220 772
rect 2216 743 2218 771
rect 2292 756 2294 778
rect 2326 776 2332 777
rect 2326 772 2327 776
rect 2331 772 2332 776
rect 2326 771 2332 772
rect 2290 755 2296 756
rect 2290 751 2291 755
rect 2295 751 2296 755
rect 2290 750 2296 751
rect 2328 743 2330 771
rect 2352 764 2354 854
rect 2462 849 2468 850
rect 2462 845 2463 849
rect 2467 845 2468 849
rect 2462 844 2468 845
rect 2678 849 2684 850
rect 2678 845 2679 849
rect 2683 845 2684 849
rect 2678 844 2684 845
rect 2894 849 2900 850
rect 2894 845 2895 849
rect 2899 845 2900 849
rect 2894 844 2900 845
rect 2464 823 2466 844
rect 2680 823 2682 844
rect 2896 823 2898 844
rect 2447 822 2451 823
rect 2447 817 2451 818
rect 2463 822 2467 823
rect 2463 817 2467 818
rect 2583 822 2587 823
rect 2583 817 2587 818
rect 2679 822 2683 823
rect 2679 817 2683 818
rect 2735 822 2739 823
rect 2735 817 2739 818
rect 2895 822 2899 823
rect 2895 817 2899 818
rect 2448 796 2450 817
rect 2584 796 2586 817
rect 2736 796 2738 817
rect 2896 796 2898 817
rect 2446 795 2452 796
rect 2446 791 2447 795
rect 2451 791 2452 795
rect 2446 790 2452 791
rect 2582 795 2588 796
rect 2582 791 2583 795
rect 2587 791 2588 795
rect 2582 790 2588 791
rect 2734 795 2740 796
rect 2734 791 2735 795
rect 2739 791 2740 795
rect 2734 790 2740 791
rect 2894 795 2900 796
rect 2894 791 2895 795
rect 2899 791 2900 795
rect 2894 790 2900 791
rect 2972 788 2974 882
rect 3128 869 3130 893
rect 3202 891 3208 892
rect 3202 887 3203 891
rect 3207 887 3208 891
rect 3202 886 3208 887
rect 3126 868 3132 869
rect 3126 864 3127 868
rect 3131 864 3132 868
rect 3126 863 3132 864
rect 3204 860 3206 886
rect 3368 869 3370 893
rect 3442 891 3448 892
rect 3442 887 3443 891
rect 3447 887 3448 891
rect 3442 886 3448 887
rect 3366 868 3372 869
rect 3366 864 3367 868
rect 3371 864 3372 868
rect 3366 863 3372 864
rect 3444 860 3446 886
rect 3616 869 3618 893
rect 3840 869 3842 893
rect 3614 868 3620 869
rect 3614 864 3615 868
rect 3619 864 3620 868
rect 3614 863 3620 864
rect 3838 868 3844 869
rect 3838 864 3839 868
rect 3843 864 3844 868
rect 3838 863 3844 864
rect 3908 860 3910 910
rect 3944 899 3946 938
rect 3943 898 3947 899
rect 3943 893 3947 894
rect 3914 891 3920 892
rect 3914 887 3915 891
rect 3919 887 3920 891
rect 3914 886 3920 887
rect 3202 859 3208 860
rect 3202 855 3203 859
rect 3207 855 3208 859
rect 3202 854 3208 855
rect 3442 859 3448 860
rect 3442 855 3443 859
rect 3447 855 3448 859
rect 3442 854 3448 855
rect 3690 859 3696 860
rect 3690 855 3691 859
rect 3695 855 3696 859
rect 3690 854 3696 855
rect 3906 859 3912 860
rect 3906 855 3907 859
rect 3911 855 3912 859
rect 3906 854 3912 855
rect 3126 849 3132 850
rect 3126 845 3127 849
rect 3131 845 3132 849
rect 3126 844 3132 845
rect 3366 849 3372 850
rect 3366 845 3367 849
rect 3371 845 3372 849
rect 3366 844 3372 845
rect 3614 849 3620 850
rect 3614 845 3615 849
rect 3619 845 3620 849
rect 3614 844 3620 845
rect 3128 823 3130 844
rect 3368 823 3370 844
rect 3616 823 3618 844
rect 3063 822 3067 823
rect 3063 817 3067 818
rect 3127 822 3131 823
rect 3127 817 3131 818
rect 3247 822 3251 823
rect 3247 817 3251 818
rect 3367 822 3371 823
rect 3367 817 3371 818
rect 3447 822 3451 823
rect 3447 817 3451 818
rect 3615 822 3619 823
rect 3615 817 3619 818
rect 3655 822 3659 823
rect 3655 817 3659 818
rect 3064 796 3066 817
rect 3248 796 3250 817
rect 3448 796 3450 817
rect 3656 796 3658 817
rect 3062 795 3068 796
rect 3062 791 3063 795
rect 3067 791 3068 795
rect 3062 790 3068 791
rect 3246 795 3252 796
rect 3246 791 3247 795
rect 3251 791 3252 795
rect 3246 790 3252 791
rect 3446 795 3452 796
rect 3446 791 3447 795
rect 3451 791 3452 795
rect 3446 790 3452 791
rect 3654 795 3660 796
rect 3654 791 3655 795
rect 3659 791 3660 795
rect 3654 790 3660 791
rect 2970 787 2976 788
rect 2402 783 2408 784
rect 2402 779 2403 783
rect 2407 779 2408 783
rect 2402 778 2408 779
rect 2522 783 2528 784
rect 2522 779 2523 783
rect 2527 779 2528 783
rect 2522 778 2528 779
rect 2658 783 2664 784
rect 2658 779 2659 783
rect 2663 779 2664 783
rect 2658 778 2664 779
rect 2810 783 2816 784
rect 2810 779 2811 783
rect 2815 779 2816 783
rect 2970 783 2971 787
rect 2975 783 2976 787
rect 3330 787 3336 788
rect 2970 782 2976 783
rect 3322 783 3328 784
rect 2810 778 2816 779
rect 3322 779 3323 783
rect 3327 779 3328 783
rect 3330 783 3331 787
rect 3335 783 3336 787
rect 3330 782 3336 783
rect 3530 787 3536 788
rect 3530 783 3531 787
rect 3535 783 3536 787
rect 3530 782 3536 783
rect 3322 778 3328 779
rect 2350 763 2356 764
rect 2350 759 2351 763
rect 2355 759 2356 763
rect 2350 758 2356 759
rect 2404 756 2406 778
rect 2446 776 2452 777
rect 2446 772 2447 776
rect 2451 772 2452 776
rect 2446 771 2452 772
rect 2402 755 2408 756
rect 2402 751 2403 755
rect 2407 751 2408 755
rect 2402 750 2408 751
rect 2448 743 2450 771
rect 2524 756 2526 778
rect 2582 776 2588 777
rect 2582 772 2583 776
rect 2587 772 2588 776
rect 2582 771 2588 772
rect 2522 755 2528 756
rect 2522 751 2523 755
rect 2527 751 2528 755
rect 2522 750 2528 751
rect 2584 743 2586 771
rect 2660 756 2662 778
rect 2734 776 2740 777
rect 2734 772 2735 776
rect 2739 772 2740 776
rect 2734 771 2740 772
rect 2658 755 2664 756
rect 2658 751 2659 755
rect 2663 751 2664 755
rect 2658 750 2664 751
rect 2736 743 2738 771
rect 2047 742 2051 743
rect 2006 737 2012 738
rect 2047 737 2051 738
rect 2215 742 2219 743
rect 2215 737 2219 738
rect 2327 742 2331 743
rect 2327 737 2331 738
rect 2375 742 2379 743
rect 2375 737 2379 738
rect 2447 742 2451 743
rect 2447 737 2451 738
rect 2495 742 2499 743
rect 2495 737 2499 738
rect 2583 742 2587 743
rect 2583 737 2587 738
rect 2623 742 2627 743
rect 2623 737 2627 738
rect 2735 742 2739 743
rect 2735 737 2739 738
rect 2767 742 2771 743
rect 2767 737 2771 738
rect 2006 733 2007 737
rect 2011 733 2012 737
rect 2006 732 2012 733
rect 1386 731 1392 732
rect 1386 727 1387 731
rect 1391 727 1392 731
rect 1386 726 1392 727
rect 1674 731 1680 732
rect 1674 727 1675 731
rect 1679 727 1680 731
rect 1674 726 1680 727
rect 1454 721 1460 722
rect 1454 717 1455 721
rect 1459 717 1460 721
rect 1454 716 1460 717
rect 1598 721 1604 722
rect 1598 717 1599 721
rect 1603 717 1604 721
rect 1598 716 1604 717
rect 2006 720 2012 721
rect 2006 716 2007 720
rect 2011 716 2012 720
rect 1456 695 1458 716
rect 1600 695 1602 716
rect 2006 715 2012 716
rect 2008 695 2010 715
rect 2048 710 2050 737
rect 2376 713 2378 737
rect 2466 735 2472 736
rect 2466 731 2467 735
rect 2471 731 2472 735
rect 2466 730 2472 731
rect 2374 712 2380 713
rect 2046 709 2052 710
rect 2046 705 2047 709
rect 2051 705 2052 709
rect 2374 708 2375 712
rect 2379 708 2380 712
rect 2374 707 2380 708
rect 2046 704 2052 705
rect 2468 704 2470 730
rect 2496 713 2498 737
rect 2590 727 2596 728
rect 2590 723 2591 727
rect 2595 723 2596 727
rect 2590 722 2596 723
rect 2494 712 2500 713
rect 2494 708 2495 712
rect 2499 708 2500 712
rect 2494 707 2500 708
rect 2592 704 2594 722
rect 2624 713 2626 737
rect 2768 713 2770 737
rect 2812 736 2814 778
rect 2894 776 2900 777
rect 2894 772 2895 776
rect 2899 772 2900 776
rect 2894 771 2900 772
rect 3062 776 3068 777
rect 3062 772 3063 776
rect 3067 772 3068 776
rect 3062 771 3068 772
rect 3246 776 3252 777
rect 3246 772 3247 776
rect 3251 772 3252 776
rect 3246 771 3252 772
rect 2896 743 2898 771
rect 3064 743 3066 771
rect 3130 751 3136 752
rect 3130 747 3131 751
rect 3135 747 3136 751
rect 3130 746 3136 747
rect 2895 742 2899 743
rect 2895 737 2899 738
rect 2911 742 2915 743
rect 2911 737 2915 738
rect 3063 742 3067 743
rect 3063 737 3067 738
rect 2810 735 2816 736
rect 2810 731 2811 735
rect 2815 731 2816 735
rect 2810 730 2816 731
rect 2842 735 2848 736
rect 2842 731 2843 735
rect 2847 731 2848 735
rect 2842 730 2848 731
rect 2622 712 2628 713
rect 2622 708 2623 712
rect 2627 708 2628 712
rect 2622 707 2628 708
rect 2766 712 2772 713
rect 2766 708 2767 712
rect 2771 708 2772 712
rect 2766 707 2772 708
rect 2844 704 2846 730
rect 2882 727 2888 728
rect 2882 723 2883 727
rect 2887 723 2888 727
rect 2882 722 2888 723
rect 2884 704 2886 722
rect 2912 713 2914 737
rect 3064 713 3066 737
rect 3118 735 3124 736
rect 3118 731 3119 735
rect 3123 731 3124 735
rect 3118 730 3124 731
rect 2910 712 2916 713
rect 2910 708 2911 712
rect 2915 708 2916 712
rect 2910 707 2916 708
rect 3062 712 3068 713
rect 3062 708 3063 712
rect 3067 708 3068 712
rect 3062 707 3068 708
rect 2466 703 2472 704
rect 2466 699 2467 703
rect 2471 699 2472 703
rect 2466 698 2472 699
rect 2582 703 2588 704
rect 2582 699 2583 703
rect 2587 699 2588 703
rect 2582 698 2588 699
rect 2590 703 2596 704
rect 2590 699 2591 703
rect 2595 699 2596 703
rect 2590 698 2596 699
rect 2842 703 2848 704
rect 2842 699 2843 703
rect 2847 699 2848 703
rect 2842 698 2848 699
rect 2882 703 2888 704
rect 2882 699 2883 703
rect 2887 699 2888 703
rect 2882 698 2888 699
rect 1407 694 1411 695
rect 1407 689 1411 690
rect 1455 694 1459 695
rect 1455 689 1459 690
rect 1519 694 1523 695
rect 1519 689 1523 690
rect 1599 694 1603 695
rect 1599 689 1603 690
rect 2007 694 2011 695
rect 2374 693 2380 694
rect 2007 689 2011 690
rect 2046 692 2052 693
rect 1368 671 1374 673
rect 1294 667 1300 668
rect 1294 663 1295 667
rect 1299 663 1300 667
rect 1294 662 1300 663
rect 1372 660 1374 671
rect 1408 668 1410 689
rect 1520 668 1522 689
rect 2008 669 2010 689
rect 2046 688 2047 692
rect 2051 688 2052 692
rect 2374 689 2375 693
rect 2379 689 2380 693
rect 2374 688 2380 689
rect 2494 693 2500 694
rect 2494 689 2495 693
rect 2499 689 2500 693
rect 2494 688 2500 689
rect 2046 687 2052 688
rect 2006 668 2012 669
rect 1406 667 1412 668
rect 1406 663 1407 667
rect 1411 663 1412 667
rect 1406 662 1412 663
rect 1518 667 1524 668
rect 1518 663 1519 667
rect 1523 663 1524 667
rect 2006 664 2007 668
rect 2011 664 2012 668
rect 2006 663 2012 664
rect 1518 662 1524 663
rect 1370 659 1376 660
rect 1370 655 1371 659
rect 1375 655 1376 659
rect 1370 654 1376 655
rect 1382 659 1388 660
rect 1382 655 1383 659
rect 1387 655 1388 659
rect 1382 654 1388 655
rect 1490 659 1496 660
rect 2048 659 2050 687
rect 2376 659 2378 688
rect 2496 659 2498 688
rect 1490 655 1491 659
rect 1495 655 1496 659
rect 1490 654 1496 655
rect 2047 658 2051 659
rect 1294 648 1300 649
rect 1294 644 1295 648
rect 1299 644 1300 648
rect 1294 643 1300 644
rect 1234 627 1240 628
rect 1234 623 1235 627
rect 1239 623 1240 627
rect 1234 622 1240 623
rect 1296 619 1298 643
rect 1384 628 1386 654
rect 1406 648 1412 649
rect 1406 644 1407 648
rect 1411 644 1412 648
rect 1406 643 1412 644
rect 1382 627 1388 628
rect 1382 623 1383 627
rect 1387 623 1388 627
rect 1382 622 1388 623
rect 1408 619 1410 643
rect 1492 628 1494 654
rect 2047 653 2051 654
rect 2111 658 2115 659
rect 2111 653 2115 654
rect 2247 658 2251 659
rect 2247 653 2251 654
rect 2375 658 2379 659
rect 2375 653 2379 654
rect 2399 658 2403 659
rect 2399 653 2403 654
rect 2495 658 2499 659
rect 2495 653 2499 654
rect 2575 658 2579 659
rect 2575 653 2579 654
rect 2006 651 2012 652
rect 1518 648 1524 649
rect 1518 644 1519 648
rect 1523 644 1524 648
rect 2006 647 2007 651
rect 2011 647 2012 651
rect 2006 646 2012 647
rect 1518 643 1524 644
rect 1490 627 1496 628
rect 1490 623 1491 627
rect 1495 623 1496 627
rect 1490 622 1496 623
rect 1520 619 1522 643
rect 1530 623 1536 624
rect 1530 619 1531 623
rect 1535 619 1536 623
rect 2008 619 2010 646
rect 2048 633 2050 653
rect 2046 632 2052 633
rect 2112 632 2114 653
rect 2248 632 2250 653
rect 2400 632 2402 653
rect 2576 632 2578 653
rect 2046 628 2047 632
rect 2051 628 2052 632
rect 2046 627 2052 628
rect 2110 631 2116 632
rect 2110 627 2111 631
rect 2115 627 2116 631
rect 2110 626 2116 627
rect 2246 631 2252 632
rect 2246 627 2247 631
rect 2251 627 2252 631
rect 2246 626 2252 627
rect 2398 631 2404 632
rect 2398 627 2399 631
rect 2403 627 2404 631
rect 2398 626 2404 627
rect 2574 631 2580 632
rect 2574 627 2575 631
rect 2579 627 2580 631
rect 2574 626 2580 627
rect 2194 623 2200 624
rect 2194 619 2195 623
rect 2199 619 2200 623
rect 1167 618 1171 619
rect 1167 613 1171 614
rect 1183 618 1187 619
rect 1183 613 1187 614
rect 1263 618 1267 619
rect 1263 613 1267 614
rect 1295 618 1299 619
rect 1295 613 1299 614
rect 1359 618 1363 619
rect 1359 613 1363 614
rect 1407 618 1411 619
rect 1407 613 1411 614
rect 1455 618 1459 619
rect 1455 613 1459 614
rect 1519 618 1523 619
rect 1530 618 1536 619
rect 2007 618 2011 619
rect 2194 618 2200 619
rect 1519 613 1523 614
rect 1146 611 1152 612
rect 1146 607 1147 611
rect 1151 607 1152 611
rect 1146 606 1152 607
rect 1168 589 1170 613
rect 1242 611 1248 612
rect 1242 607 1243 611
rect 1247 607 1248 611
rect 1242 606 1248 607
rect 1070 588 1076 589
rect 1070 584 1071 588
rect 1075 584 1076 588
rect 1070 583 1076 584
rect 1166 588 1172 589
rect 1166 584 1167 588
rect 1171 584 1172 588
rect 1166 583 1172 584
rect 1244 580 1246 606
rect 1264 589 1266 613
rect 1338 611 1344 612
rect 1338 607 1339 611
rect 1343 607 1344 611
rect 1338 606 1344 607
rect 1330 603 1336 604
rect 1330 599 1331 603
rect 1335 599 1336 603
rect 1330 598 1336 599
rect 1262 588 1268 589
rect 1262 584 1263 588
rect 1267 584 1268 588
rect 1262 583 1268 584
rect 762 579 768 580
rect 762 575 763 579
rect 767 575 768 579
rect 762 574 768 575
rect 1042 579 1048 580
rect 1042 575 1043 579
rect 1047 575 1048 579
rect 1042 574 1048 575
rect 1058 579 1064 580
rect 1058 575 1059 579
rect 1063 575 1064 579
rect 1058 574 1064 575
rect 1242 579 1248 580
rect 1242 575 1243 579
rect 1247 575 1248 579
rect 1242 574 1248 575
rect 686 569 692 570
rect 110 568 116 569
rect 110 564 111 568
rect 115 564 116 568
rect 686 565 687 569
rect 691 565 692 569
rect 686 564 692 565
rect 782 569 788 570
rect 782 565 783 569
rect 787 565 788 569
rect 782 564 788 565
rect 878 569 884 570
rect 878 565 879 569
rect 883 565 884 569
rect 878 564 884 565
rect 974 569 980 570
rect 974 565 975 569
rect 979 565 980 569
rect 974 564 980 565
rect 1070 569 1076 570
rect 1070 565 1071 569
rect 1075 565 1076 569
rect 1070 564 1076 565
rect 1166 569 1172 570
rect 1166 565 1167 569
rect 1171 565 1172 569
rect 1166 564 1172 565
rect 1262 569 1268 570
rect 1262 565 1263 569
rect 1267 565 1268 569
rect 1262 564 1268 565
rect 110 563 116 564
rect 112 523 114 563
rect 688 523 690 564
rect 784 523 786 564
rect 880 523 882 564
rect 976 523 978 564
rect 1072 523 1074 564
rect 1168 523 1170 564
rect 1264 523 1266 564
rect 111 522 115 523
rect 111 517 115 518
rect 383 522 387 523
rect 383 517 387 518
rect 479 522 483 523
rect 479 517 483 518
rect 575 522 579 523
rect 575 517 579 518
rect 671 522 675 523
rect 671 517 675 518
rect 687 522 691 523
rect 687 517 691 518
rect 767 522 771 523
rect 767 517 771 518
rect 783 522 787 523
rect 783 517 787 518
rect 863 522 867 523
rect 863 517 867 518
rect 879 522 883 523
rect 879 517 883 518
rect 959 522 963 523
rect 959 517 963 518
rect 975 522 979 523
rect 975 517 979 518
rect 1055 522 1059 523
rect 1055 517 1059 518
rect 1071 522 1075 523
rect 1071 517 1075 518
rect 1151 522 1155 523
rect 1151 517 1155 518
rect 1167 522 1171 523
rect 1167 517 1171 518
rect 1247 522 1251 523
rect 1247 517 1251 518
rect 1263 522 1267 523
rect 1263 517 1267 518
rect 112 497 114 517
rect 110 496 116 497
rect 384 496 386 517
rect 480 496 482 517
rect 576 496 578 517
rect 672 496 674 517
rect 768 496 770 517
rect 864 496 866 517
rect 960 496 962 517
rect 1056 496 1058 517
rect 1152 496 1154 517
rect 1248 496 1250 517
rect 110 492 111 496
rect 115 492 116 496
rect 110 491 116 492
rect 382 495 388 496
rect 382 491 383 495
rect 387 491 388 495
rect 382 490 388 491
rect 478 495 484 496
rect 478 491 479 495
rect 483 491 484 495
rect 478 490 484 491
rect 574 495 580 496
rect 574 491 575 495
rect 579 491 580 495
rect 574 490 580 491
rect 670 495 676 496
rect 670 491 671 495
rect 675 491 676 495
rect 670 490 676 491
rect 766 495 772 496
rect 766 491 767 495
rect 771 491 772 495
rect 766 490 772 491
rect 862 495 868 496
rect 862 491 863 495
rect 867 491 868 495
rect 862 490 868 491
rect 958 495 964 496
rect 958 491 959 495
rect 963 491 964 495
rect 958 490 964 491
rect 1054 495 1060 496
rect 1054 491 1055 495
rect 1059 491 1060 495
rect 1054 490 1060 491
rect 1150 495 1156 496
rect 1150 491 1151 495
rect 1155 491 1156 495
rect 1150 490 1156 491
rect 1246 495 1252 496
rect 1246 491 1247 495
rect 1251 491 1252 495
rect 1246 490 1252 491
rect 1332 488 1334 598
rect 1340 580 1342 606
rect 1360 589 1362 613
rect 1434 611 1440 612
rect 1434 607 1435 611
rect 1439 607 1440 611
rect 1434 606 1440 607
rect 1358 588 1364 589
rect 1358 584 1359 588
rect 1363 584 1364 588
rect 1358 583 1364 584
rect 1436 580 1438 606
rect 1456 589 1458 613
rect 1454 588 1460 589
rect 1454 584 1455 588
rect 1459 584 1460 588
rect 1454 583 1460 584
rect 1532 580 1534 618
rect 2007 613 2011 614
rect 2046 615 2052 616
rect 2008 586 2010 613
rect 2046 611 2047 615
rect 2051 611 2052 615
rect 2046 610 2052 611
rect 2110 612 2116 613
rect 2006 585 2012 586
rect 2006 581 2007 585
rect 2011 581 2012 585
rect 2006 580 2012 581
rect 1338 579 1344 580
rect 1338 575 1339 579
rect 1343 575 1344 579
rect 1338 574 1344 575
rect 1434 579 1440 580
rect 1434 575 1435 579
rect 1439 575 1440 579
rect 1434 574 1440 575
rect 1530 579 1536 580
rect 2048 579 2050 610
rect 2110 608 2111 612
rect 2115 608 2116 612
rect 2110 607 2116 608
rect 2112 579 2114 607
rect 2196 592 2198 618
rect 2246 612 2252 613
rect 2246 608 2247 612
rect 2251 608 2252 612
rect 2246 607 2252 608
rect 2398 612 2404 613
rect 2398 608 2399 612
rect 2403 608 2404 612
rect 2398 607 2404 608
rect 2574 612 2580 613
rect 2574 608 2575 612
rect 2579 608 2580 612
rect 2574 607 2580 608
rect 2194 591 2200 592
rect 2194 587 2195 591
rect 2199 587 2200 591
rect 2194 586 2200 587
rect 2248 579 2250 607
rect 2400 579 2402 607
rect 2576 579 2578 607
rect 2584 592 2586 698
rect 2622 693 2628 694
rect 2622 689 2623 693
rect 2627 689 2628 693
rect 2622 688 2628 689
rect 2766 693 2772 694
rect 2766 689 2767 693
rect 2771 689 2772 693
rect 2766 688 2772 689
rect 2910 693 2916 694
rect 2910 689 2911 693
rect 2915 689 2916 693
rect 2910 688 2916 689
rect 3062 693 3068 694
rect 3062 689 3063 693
rect 3067 689 3068 693
rect 3062 688 3068 689
rect 2624 659 2626 688
rect 2768 659 2770 688
rect 2912 659 2914 688
rect 3064 659 3066 688
rect 2623 658 2627 659
rect 2623 653 2627 654
rect 2759 658 2763 659
rect 2759 653 2763 654
rect 2767 658 2771 659
rect 2767 653 2771 654
rect 2911 658 2915 659
rect 2911 653 2915 654
rect 2943 658 2947 659
rect 2943 653 2947 654
rect 3063 658 3067 659
rect 3063 653 3067 654
rect 2760 632 2762 653
rect 2944 632 2946 653
rect 2758 631 2764 632
rect 2758 627 2759 631
rect 2763 627 2764 631
rect 2758 626 2764 627
rect 2942 631 2948 632
rect 2942 627 2943 631
rect 2947 627 2948 631
rect 2942 626 2948 627
rect 3120 624 3122 730
rect 3132 704 3134 746
rect 3248 743 3250 771
rect 3215 742 3219 743
rect 3215 737 3219 738
rect 3247 742 3251 743
rect 3247 737 3251 738
rect 3216 713 3218 737
rect 3324 736 3326 778
rect 3332 756 3334 782
rect 3446 776 3452 777
rect 3446 772 3447 776
rect 3451 772 3452 776
rect 3446 771 3452 772
rect 3330 755 3336 756
rect 3330 751 3331 755
rect 3335 751 3336 755
rect 3330 750 3336 751
rect 3448 743 3450 771
rect 3532 756 3534 782
rect 3654 776 3660 777
rect 3654 772 3655 776
rect 3659 772 3660 776
rect 3654 771 3660 772
rect 3530 755 3536 756
rect 3530 751 3531 755
rect 3535 751 3536 755
rect 3530 750 3536 751
rect 3656 743 3658 771
rect 3692 756 3694 854
rect 3838 849 3844 850
rect 3838 845 3839 849
rect 3843 845 3844 849
rect 3838 844 3844 845
rect 3840 823 3842 844
rect 3839 822 3843 823
rect 3839 817 3843 818
rect 3840 796 3842 817
rect 3838 795 3844 796
rect 3838 791 3839 795
rect 3843 791 3844 795
rect 3838 790 3844 791
rect 3916 788 3918 886
rect 3944 866 3946 893
rect 3942 865 3948 866
rect 3942 861 3943 865
rect 3947 861 3948 865
rect 3942 860 3948 861
rect 3942 848 3948 849
rect 3942 844 3943 848
rect 3947 844 3948 848
rect 3942 843 3948 844
rect 3944 823 3946 843
rect 3943 822 3947 823
rect 3943 817 3947 818
rect 3944 797 3946 817
rect 3942 796 3948 797
rect 3942 792 3943 796
rect 3947 792 3948 796
rect 3942 791 3948 792
rect 3914 787 3920 788
rect 3914 783 3915 787
rect 3919 783 3920 787
rect 3914 782 3920 783
rect 3942 779 3948 780
rect 3838 776 3844 777
rect 3838 772 3839 776
rect 3843 772 3844 776
rect 3942 775 3943 779
rect 3947 775 3948 779
rect 3942 774 3948 775
rect 3838 771 3844 772
rect 3690 755 3696 756
rect 3690 751 3691 755
rect 3695 751 3696 755
rect 3690 750 3696 751
rect 3840 743 3842 771
rect 3906 751 3912 752
rect 3906 747 3907 751
rect 3911 747 3912 751
rect 3906 746 3912 747
rect 3367 742 3371 743
rect 3367 737 3371 738
rect 3447 742 3451 743
rect 3447 737 3451 738
rect 3519 742 3523 743
rect 3519 737 3523 738
rect 3655 742 3659 743
rect 3655 737 3659 738
rect 3679 742 3683 743
rect 3679 737 3683 738
rect 3839 742 3843 743
rect 3839 737 3843 738
rect 3322 735 3328 736
rect 3322 731 3323 735
rect 3327 731 3328 735
rect 3322 730 3328 731
rect 3368 713 3370 737
rect 3520 713 3522 737
rect 3594 735 3600 736
rect 3594 731 3595 735
rect 3599 731 3600 735
rect 3594 730 3600 731
rect 3214 712 3220 713
rect 3214 708 3215 712
rect 3219 708 3220 712
rect 3214 707 3220 708
rect 3366 712 3372 713
rect 3366 708 3367 712
rect 3371 708 3372 712
rect 3366 707 3372 708
rect 3518 712 3524 713
rect 3518 708 3519 712
rect 3523 708 3524 712
rect 3518 707 3524 708
rect 3596 704 3598 730
rect 3680 713 3682 737
rect 3840 713 3842 737
rect 3894 735 3900 736
rect 3894 731 3895 735
rect 3899 731 3900 735
rect 3894 730 3902 731
rect 3896 729 3902 730
rect 3678 712 3684 713
rect 3678 708 3679 712
rect 3683 708 3684 712
rect 3678 707 3684 708
rect 3838 712 3844 713
rect 3838 708 3839 712
rect 3843 708 3844 712
rect 3838 707 3844 708
rect 3130 703 3136 704
rect 3130 699 3131 703
rect 3135 699 3136 703
rect 3130 698 3136 699
rect 3594 703 3600 704
rect 3594 699 3595 703
rect 3599 699 3600 703
rect 3594 698 3600 699
rect 3746 703 3752 704
rect 3746 699 3747 703
rect 3751 699 3752 703
rect 3746 698 3752 699
rect 3214 693 3220 694
rect 3214 689 3215 693
rect 3219 689 3220 693
rect 3214 688 3220 689
rect 3366 693 3372 694
rect 3366 689 3367 693
rect 3371 689 3372 693
rect 3366 688 3372 689
rect 3518 693 3524 694
rect 3518 689 3519 693
rect 3523 689 3524 693
rect 3518 688 3524 689
rect 3678 693 3684 694
rect 3678 689 3679 693
rect 3683 689 3684 693
rect 3678 688 3684 689
rect 3216 659 3218 688
rect 3368 659 3370 688
rect 3520 659 3522 688
rect 3680 659 3682 688
rect 3127 658 3131 659
rect 3127 653 3131 654
rect 3215 658 3219 659
rect 3215 653 3219 654
rect 3303 658 3307 659
rect 3303 653 3307 654
rect 3367 658 3371 659
rect 3367 653 3371 654
rect 3479 658 3483 659
rect 3479 653 3483 654
rect 3519 658 3523 659
rect 3519 653 3523 654
rect 3655 658 3659 659
rect 3655 653 3659 654
rect 3679 658 3683 659
rect 3679 653 3683 654
rect 3128 632 3130 653
rect 3304 632 3306 653
rect 3480 632 3482 653
rect 3656 632 3658 653
rect 3126 631 3132 632
rect 3126 627 3127 631
rect 3131 627 3132 631
rect 3126 626 3132 627
rect 3302 631 3308 632
rect 3302 627 3303 631
rect 3307 627 3308 631
rect 3302 626 3308 627
rect 3478 631 3484 632
rect 3478 627 3479 631
rect 3483 627 3484 631
rect 3478 626 3484 627
rect 3654 631 3660 632
rect 3654 627 3655 631
rect 3659 627 3660 631
rect 3654 626 3660 627
rect 2658 623 2664 624
rect 2650 619 2656 620
rect 2650 615 2651 619
rect 2655 615 2656 619
rect 2658 619 2659 623
rect 2663 619 2664 623
rect 3118 623 3124 624
rect 2658 618 2664 619
rect 3018 619 3024 620
rect 2650 614 2656 615
rect 2652 592 2654 614
rect 2660 600 2662 618
rect 3018 615 3019 619
rect 3023 615 3024 619
rect 3118 619 3119 623
rect 3123 619 3124 623
rect 3390 623 3396 624
rect 3118 618 3124 619
rect 3378 619 3384 620
rect 3018 614 3024 615
rect 3378 615 3379 619
rect 3383 615 3384 619
rect 3390 619 3391 623
rect 3395 619 3396 623
rect 3390 618 3396 619
rect 3598 623 3604 624
rect 3598 619 3599 623
rect 3603 619 3604 623
rect 3598 618 3604 619
rect 3378 614 3384 615
rect 2758 612 2764 613
rect 2758 608 2759 612
rect 2763 608 2764 612
rect 2758 607 2764 608
rect 2942 612 2948 613
rect 2942 608 2943 612
rect 2947 608 2948 612
rect 2942 607 2948 608
rect 2658 599 2664 600
rect 2658 595 2659 599
rect 2663 595 2664 599
rect 2658 594 2664 595
rect 2582 591 2588 592
rect 2582 587 2583 591
rect 2587 587 2588 591
rect 2582 586 2588 587
rect 2650 591 2656 592
rect 2650 587 2651 591
rect 2655 587 2656 591
rect 2650 586 2656 587
rect 2760 579 2762 607
rect 2944 579 2946 607
rect 3020 592 3022 614
rect 3126 612 3132 613
rect 3126 608 3127 612
rect 3131 608 3132 612
rect 3126 607 3132 608
rect 3302 612 3308 613
rect 3302 608 3303 612
rect 3307 608 3308 612
rect 3302 607 3308 608
rect 3018 591 3024 592
rect 2954 587 2960 588
rect 2954 583 2955 587
rect 2959 583 2960 587
rect 3018 587 3019 591
rect 3023 587 3024 591
rect 3018 586 3024 587
rect 2954 582 2960 583
rect 1530 575 1531 579
rect 1535 575 1536 579
rect 1530 574 1536 575
rect 2047 578 2051 579
rect 2047 573 2051 574
rect 2071 578 2075 579
rect 2071 573 2075 574
rect 2111 578 2115 579
rect 2111 573 2115 574
rect 2183 578 2187 579
rect 2183 573 2187 574
rect 2247 578 2251 579
rect 2247 573 2251 574
rect 2335 578 2339 579
rect 2335 573 2339 574
rect 2399 578 2403 579
rect 2399 573 2403 574
rect 2503 578 2507 579
rect 2503 573 2507 574
rect 2575 578 2579 579
rect 2575 573 2579 574
rect 2687 578 2691 579
rect 2687 573 2691 574
rect 2759 578 2763 579
rect 2759 573 2763 574
rect 2879 578 2883 579
rect 2879 573 2883 574
rect 2943 578 2947 579
rect 2943 573 2947 574
rect 1358 569 1364 570
rect 1358 565 1359 569
rect 1363 565 1364 569
rect 1358 564 1364 565
rect 1454 569 1460 570
rect 1454 565 1455 569
rect 1459 565 1460 569
rect 1454 564 1460 565
rect 2006 568 2012 569
rect 2006 564 2007 568
rect 2011 564 2012 568
rect 1360 523 1362 564
rect 1456 523 1458 564
rect 2006 563 2012 564
rect 2008 523 2010 563
rect 2048 546 2050 573
rect 2072 549 2074 573
rect 2146 571 2152 572
rect 2146 567 2147 571
rect 2151 567 2152 571
rect 2146 566 2152 567
rect 2070 548 2076 549
rect 2046 545 2052 546
rect 2046 541 2047 545
rect 2051 541 2052 545
rect 2070 544 2071 548
rect 2075 544 2076 548
rect 2070 543 2076 544
rect 2046 540 2052 541
rect 2148 540 2150 566
rect 2184 549 2186 573
rect 2258 571 2264 572
rect 2258 567 2259 571
rect 2263 567 2264 571
rect 2258 566 2264 567
rect 2182 548 2188 549
rect 2182 544 2183 548
rect 2187 544 2188 548
rect 2182 543 2188 544
rect 2260 540 2262 566
rect 2336 549 2338 573
rect 2410 571 2416 572
rect 2410 567 2411 571
rect 2415 567 2416 571
rect 2410 566 2416 567
rect 2334 548 2340 549
rect 2334 544 2335 548
rect 2339 544 2340 548
rect 2334 543 2340 544
rect 2412 540 2414 566
rect 2504 549 2506 573
rect 2688 549 2690 573
rect 2880 549 2882 573
rect 2502 548 2508 549
rect 2502 544 2503 548
rect 2507 544 2508 548
rect 2502 543 2508 544
rect 2686 548 2692 549
rect 2686 544 2687 548
rect 2691 544 2692 548
rect 2686 543 2692 544
rect 2878 548 2884 549
rect 2878 544 2879 548
rect 2883 544 2884 548
rect 2878 543 2884 544
rect 2956 540 2958 582
rect 3128 579 3130 607
rect 3304 579 3306 607
rect 3071 578 3075 579
rect 3071 573 3075 574
rect 3127 578 3131 579
rect 3127 573 3131 574
rect 3263 578 3267 579
rect 3263 573 3267 574
rect 3303 578 3307 579
rect 3303 573 3307 574
rect 2962 571 2968 572
rect 2962 567 2963 571
rect 2967 567 2968 571
rect 2962 566 2968 567
rect 2964 540 2966 566
rect 3072 549 3074 573
rect 3174 571 3180 572
rect 3174 567 3175 571
rect 3179 567 3180 571
rect 3174 566 3180 567
rect 3234 571 3240 572
rect 3234 567 3235 571
rect 3239 567 3240 571
rect 3234 566 3240 567
rect 3070 548 3076 549
rect 3070 544 3071 548
rect 3075 544 3076 548
rect 3070 543 3076 544
rect 3176 540 3178 566
rect 2146 539 2152 540
rect 2146 535 2147 539
rect 2151 535 2152 539
rect 2146 534 2152 535
rect 2258 539 2264 540
rect 2258 535 2259 539
rect 2263 535 2264 539
rect 2258 534 2264 535
rect 2410 539 2416 540
rect 2410 535 2411 539
rect 2415 535 2416 539
rect 2410 534 2416 535
rect 2658 539 2664 540
rect 2658 535 2659 539
rect 2663 535 2664 539
rect 2658 534 2664 535
rect 2954 539 2960 540
rect 2954 535 2955 539
rect 2959 535 2960 539
rect 2954 534 2960 535
rect 2962 539 2968 540
rect 2962 535 2963 539
rect 2967 535 2968 539
rect 2962 534 2968 535
rect 3174 539 3180 540
rect 3174 535 3175 539
rect 3179 535 3180 539
rect 3174 534 3180 535
rect 2070 529 2076 530
rect 2046 528 2052 529
rect 2046 524 2047 528
rect 2051 524 2052 528
rect 2070 525 2071 529
rect 2075 525 2076 529
rect 2070 524 2076 525
rect 2182 529 2188 530
rect 2182 525 2183 529
rect 2187 525 2188 529
rect 2182 524 2188 525
rect 2334 529 2340 530
rect 2334 525 2335 529
rect 2339 525 2340 529
rect 2334 524 2340 525
rect 2502 529 2508 530
rect 2502 525 2503 529
rect 2507 525 2508 529
rect 2502 524 2508 525
rect 2046 523 2052 524
rect 1343 522 1347 523
rect 1343 517 1347 518
rect 1359 522 1363 523
rect 1359 517 1363 518
rect 1439 522 1443 523
rect 1439 517 1443 518
rect 1455 522 1459 523
rect 1455 517 1459 518
rect 1535 522 1539 523
rect 1535 517 1539 518
rect 2007 522 2011 523
rect 2007 517 2011 518
rect 1344 496 1346 517
rect 1440 496 1442 517
rect 1536 496 1538 517
rect 2008 497 2010 517
rect 2048 503 2050 523
rect 2072 503 2074 524
rect 2184 503 2186 524
rect 2336 503 2338 524
rect 2504 503 2506 524
rect 2047 502 2051 503
rect 2047 497 2051 498
rect 2071 502 2075 503
rect 2071 497 2075 498
rect 2183 502 2187 503
rect 2183 497 2187 498
rect 2319 502 2323 503
rect 2319 497 2323 498
rect 2335 502 2339 503
rect 2335 497 2339 498
rect 2463 502 2467 503
rect 2463 497 2467 498
rect 2503 502 2507 503
rect 2503 497 2507 498
rect 2615 502 2619 503
rect 2615 497 2619 498
rect 2006 496 2012 497
rect 1342 495 1348 496
rect 1342 491 1343 495
rect 1347 491 1348 495
rect 1342 490 1348 491
rect 1438 495 1444 496
rect 1438 491 1439 495
rect 1443 491 1444 495
rect 1438 490 1444 491
rect 1534 495 1540 496
rect 1534 491 1535 495
rect 1539 491 1540 495
rect 2006 492 2007 496
rect 2011 492 2012 496
rect 2006 491 2012 492
rect 1534 490 1540 491
rect 1330 487 1336 488
rect 458 483 464 484
rect 110 479 116 480
rect 110 475 111 479
rect 115 475 116 479
rect 458 479 459 483
rect 463 479 464 483
rect 458 478 464 479
rect 554 483 560 484
rect 554 479 555 483
rect 559 479 560 483
rect 554 478 560 479
rect 650 483 656 484
rect 650 479 651 483
rect 655 479 656 483
rect 650 478 656 479
rect 746 483 752 484
rect 746 479 747 483
rect 751 479 752 483
rect 746 478 752 479
rect 842 483 848 484
rect 842 479 843 483
rect 847 479 848 483
rect 842 478 848 479
rect 938 483 944 484
rect 938 479 939 483
rect 943 479 944 483
rect 938 478 944 479
rect 1034 483 1040 484
rect 1034 479 1035 483
rect 1039 479 1040 483
rect 1034 478 1040 479
rect 1130 483 1136 484
rect 1130 479 1131 483
rect 1135 479 1136 483
rect 1130 478 1136 479
rect 1226 483 1232 484
rect 1226 479 1227 483
rect 1231 479 1232 483
rect 1330 483 1331 487
rect 1335 483 1336 487
rect 1330 482 1336 483
rect 1514 483 1520 484
rect 1226 478 1232 479
rect 1514 479 1515 483
rect 1519 479 1520 483
rect 1514 478 1520 479
rect 2006 479 2012 480
rect 110 474 116 475
rect 382 476 388 477
rect 112 435 114 474
rect 382 472 383 476
rect 387 472 388 476
rect 382 471 388 472
rect 384 435 386 471
rect 460 456 462 478
rect 478 476 484 477
rect 478 472 479 476
rect 483 472 484 476
rect 478 471 484 472
rect 458 455 464 456
rect 458 451 459 455
rect 463 451 464 455
rect 458 450 464 451
rect 480 435 482 471
rect 556 456 558 478
rect 574 476 580 477
rect 574 472 575 476
rect 579 472 580 476
rect 574 471 580 472
rect 554 455 560 456
rect 554 451 555 455
rect 559 451 560 455
rect 554 450 560 451
rect 576 435 578 471
rect 652 456 654 478
rect 670 476 676 477
rect 670 472 671 476
rect 675 472 676 476
rect 670 471 676 472
rect 650 455 656 456
rect 650 451 651 455
rect 655 451 656 455
rect 650 450 656 451
rect 672 435 674 471
rect 748 456 750 478
rect 766 476 772 477
rect 766 472 767 476
rect 771 472 772 476
rect 766 471 772 472
rect 746 455 752 456
rect 746 451 747 455
rect 751 451 752 455
rect 746 450 752 451
rect 768 435 770 471
rect 844 456 846 478
rect 862 476 868 477
rect 862 472 863 476
rect 867 472 868 476
rect 862 471 868 472
rect 842 455 848 456
rect 842 451 843 455
rect 847 451 848 455
rect 842 450 848 451
rect 864 435 866 471
rect 940 456 942 478
rect 958 476 964 477
rect 958 472 959 476
rect 963 472 964 476
rect 958 471 964 472
rect 938 455 944 456
rect 938 451 939 455
rect 943 451 944 455
rect 938 450 944 451
rect 960 435 962 471
rect 1036 456 1038 478
rect 1054 476 1060 477
rect 1054 472 1055 476
rect 1059 472 1060 476
rect 1054 471 1060 472
rect 1034 455 1040 456
rect 1034 451 1035 455
rect 1039 451 1040 455
rect 1034 450 1040 451
rect 966 447 972 448
rect 966 443 967 447
rect 971 443 972 447
rect 966 442 972 443
rect 111 434 115 435
rect 111 429 115 430
rect 383 434 387 435
rect 383 429 387 430
rect 479 434 483 435
rect 479 429 483 430
rect 487 434 491 435
rect 487 429 491 430
rect 575 434 579 435
rect 575 429 579 430
rect 583 434 587 435
rect 583 429 587 430
rect 671 434 675 435
rect 671 429 675 430
rect 687 434 691 435
rect 687 429 691 430
rect 767 434 771 435
rect 767 429 771 430
rect 791 434 795 435
rect 791 429 795 430
rect 863 434 867 435
rect 863 429 867 430
rect 895 434 899 435
rect 895 429 899 430
rect 959 434 963 435
rect 959 429 963 430
rect 112 402 114 429
rect 488 405 490 429
rect 562 427 568 428
rect 538 423 544 424
rect 538 418 539 423
rect 543 418 544 423
rect 562 423 563 427
rect 567 423 568 427
rect 562 422 568 423
rect 539 415 543 416
rect 486 404 492 405
rect 110 401 116 402
rect 110 397 111 401
rect 115 397 116 401
rect 486 400 487 404
rect 491 400 492 404
rect 486 399 492 400
rect 110 396 116 397
rect 564 396 566 422
rect 584 405 586 429
rect 658 427 664 428
rect 658 423 659 427
rect 663 423 664 427
rect 658 422 664 423
rect 582 404 588 405
rect 582 400 583 404
rect 587 400 588 404
rect 582 399 588 400
rect 660 396 662 422
rect 688 405 690 429
rect 792 405 794 429
rect 859 420 863 421
rect 859 415 863 416
rect 686 404 692 405
rect 686 400 687 404
rect 691 400 692 404
rect 686 399 692 400
rect 790 404 796 405
rect 790 400 791 404
rect 795 400 796 404
rect 790 399 796 400
rect 562 395 568 396
rect 562 391 563 395
rect 567 391 568 395
rect 562 390 568 391
rect 658 395 664 396
rect 658 391 659 395
rect 663 391 664 395
rect 658 390 664 391
rect 486 385 492 386
rect 110 384 116 385
rect 110 380 111 384
rect 115 380 116 384
rect 486 381 487 385
rect 491 381 492 385
rect 486 380 492 381
rect 582 385 588 386
rect 582 381 583 385
rect 587 381 588 385
rect 582 380 588 381
rect 686 385 692 386
rect 686 381 687 385
rect 691 381 692 385
rect 686 380 692 381
rect 790 385 796 386
rect 790 381 791 385
rect 795 381 796 385
rect 790 380 796 381
rect 110 379 116 380
rect 112 355 114 379
rect 488 355 490 380
rect 584 355 586 380
rect 688 355 690 380
rect 792 355 794 380
rect 111 354 115 355
rect 111 349 115 350
rect 327 354 331 355
rect 327 349 331 350
rect 463 354 467 355
rect 463 349 467 350
rect 487 354 491 355
rect 487 349 491 350
rect 583 354 587 355
rect 583 349 587 350
rect 615 354 619 355
rect 615 349 619 350
rect 687 354 691 355
rect 687 349 691 350
rect 767 354 771 355
rect 767 349 771 350
rect 791 354 795 355
rect 791 349 795 350
rect 112 329 114 349
rect 110 328 116 329
rect 328 328 330 349
rect 464 328 466 349
rect 616 328 618 349
rect 768 328 770 349
rect 110 324 111 328
rect 115 324 116 328
rect 110 323 116 324
rect 326 327 332 328
rect 326 323 327 327
rect 331 323 332 327
rect 326 322 332 323
rect 462 327 468 328
rect 462 323 463 327
rect 467 323 468 327
rect 462 322 468 323
rect 614 327 620 328
rect 614 323 615 327
rect 619 323 620 327
rect 614 322 620 323
rect 766 327 772 328
rect 766 323 767 327
rect 771 323 772 327
rect 766 322 772 323
rect 860 320 862 415
rect 896 405 898 429
rect 894 404 900 405
rect 894 400 895 404
rect 899 400 900 404
rect 894 399 900 400
rect 968 396 970 442
rect 1056 435 1058 471
rect 1132 456 1134 478
rect 1150 476 1156 477
rect 1150 472 1151 476
rect 1155 472 1156 476
rect 1150 471 1156 472
rect 1130 455 1136 456
rect 1130 451 1131 455
rect 1135 451 1136 455
rect 1130 450 1136 451
rect 1152 435 1154 471
rect 1228 456 1230 478
rect 1246 476 1252 477
rect 1246 472 1247 476
rect 1251 472 1252 476
rect 1246 471 1252 472
rect 1342 476 1348 477
rect 1342 472 1343 476
rect 1347 472 1348 476
rect 1342 471 1348 472
rect 1438 476 1444 477
rect 1438 472 1439 476
rect 1443 472 1444 476
rect 1438 471 1444 472
rect 1226 455 1232 456
rect 1226 451 1227 455
rect 1231 451 1232 455
rect 1226 450 1232 451
rect 1248 435 1250 471
rect 1344 435 1346 471
rect 1440 435 1442 471
rect 1516 456 1518 478
rect 1534 476 1540 477
rect 1534 472 1535 476
rect 1539 472 1540 476
rect 2006 475 2007 479
rect 2011 475 2012 479
rect 2048 477 2050 497
rect 2006 474 2012 475
rect 2046 476 2052 477
rect 2184 476 2186 497
rect 2320 476 2322 497
rect 2464 476 2466 497
rect 2616 476 2618 497
rect 1534 471 1540 472
rect 1514 455 1520 456
rect 1494 451 1500 452
rect 1494 447 1495 451
rect 1499 447 1500 451
rect 1514 451 1515 455
rect 1519 451 1520 455
rect 1514 450 1520 451
rect 1494 446 1500 447
rect 999 434 1003 435
rect 999 429 1003 430
rect 1055 434 1059 435
rect 1055 429 1059 430
rect 1103 434 1107 435
rect 1103 429 1107 430
rect 1151 434 1155 435
rect 1151 429 1155 430
rect 1207 434 1211 435
rect 1207 429 1211 430
rect 1247 434 1251 435
rect 1247 429 1251 430
rect 1319 434 1323 435
rect 1319 429 1323 430
rect 1343 434 1347 435
rect 1343 429 1347 430
rect 1431 434 1435 435
rect 1431 429 1435 430
rect 1439 434 1443 435
rect 1439 429 1443 430
rect 1000 405 1002 429
rect 1104 405 1106 429
rect 1186 427 1192 428
rect 1186 423 1187 427
rect 1191 423 1192 427
rect 1186 422 1192 423
rect 998 404 1004 405
rect 998 400 999 404
rect 1003 400 1004 404
rect 998 399 1004 400
rect 1102 404 1108 405
rect 1102 400 1103 404
rect 1107 400 1108 404
rect 1102 399 1108 400
rect 1188 396 1190 422
rect 1208 405 1210 429
rect 1320 405 1322 429
rect 1418 427 1424 428
rect 1418 423 1419 427
rect 1423 423 1424 427
rect 1418 422 1424 423
rect 1394 419 1400 420
rect 1394 415 1395 419
rect 1399 415 1400 419
rect 1394 414 1400 415
rect 1206 404 1212 405
rect 1206 400 1207 404
rect 1211 400 1212 404
rect 1206 399 1212 400
rect 1318 404 1324 405
rect 1318 400 1319 404
rect 1323 400 1324 404
rect 1318 399 1324 400
rect 1396 396 1398 414
rect 966 395 972 396
rect 966 391 967 395
rect 971 391 972 395
rect 966 390 972 391
rect 1074 395 1080 396
rect 1074 391 1075 395
rect 1079 391 1080 395
rect 1074 390 1080 391
rect 1186 395 1192 396
rect 1186 391 1187 395
rect 1191 391 1192 395
rect 1186 390 1192 391
rect 1394 395 1400 396
rect 1394 391 1395 395
rect 1399 391 1400 395
rect 1394 390 1400 391
rect 894 385 900 386
rect 894 381 895 385
rect 899 381 900 385
rect 894 380 900 381
rect 998 385 1004 386
rect 998 381 999 385
rect 1003 381 1004 385
rect 998 380 1004 381
rect 896 355 898 380
rect 1000 355 1002 380
rect 895 354 899 355
rect 895 349 899 350
rect 919 354 923 355
rect 919 349 923 350
rect 999 354 1003 355
rect 999 349 1003 350
rect 1063 354 1067 355
rect 1063 349 1067 350
rect 920 328 922 349
rect 1064 328 1066 349
rect 918 327 924 328
rect 918 323 919 327
rect 923 323 924 327
rect 918 322 924 323
rect 1062 327 1068 328
rect 1062 323 1063 327
rect 1067 323 1068 327
rect 1062 322 1068 323
rect 858 319 864 320
rect 402 315 408 316
rect 110 311 116 312
rect 110 307 111 311
rect 115 307 116 311
rect 402 311 403 315
rect 407 311 408 315
rect 402 310 408 311
rect 538 315 544 316
rect 538 311 539 315
rect 543 311 544 315
rect 538 310 544 311
rect 690 315 696 316
rect 690 311 691 315
rect 695 311 696 315
rect 690 310 696 311
rect 842 315 848 316
rect 842 311 843 315
rect 847 311 848 315
rect 858 315 859 319
rect 863 315 864 319
rect 858 314 864 315
rect 842 310 848 311
rect 110 306 116 307
rect 326 308 332 309
rect 112 271 114 306
rect 326 304 327 308
rect 331 304 332 308
rect 326 303 332 304
rect 328 271 330 303
rect 404 288 406 310
rect 462 308 468 309
rect 462 304 463 308
rect 467 304 468 308
rect 462 303 468 304
rect 402 287 408 288
rect 402 283 403 287
rect 407 283 408 287
rect 402 282 408 283
rect 464 271 466 303
rect 540 288 542 310
rect 614 308 620 309
rect 614 304 615 308
rect 619 304 620 308
rect 614 303 620 304
rect 538 287 544 288
rect 538 283 539 287
rect 543 283 544 287
rect 538 282 544 283
rect 616 271 618 303
rect 692 288 694 310
rect 766 308 772 309
rect 766 304 767 308
rect 771 304 772 308
rect 766 303 772 304
rect 690 287 696 288
rect 690 283 691 287
rect 695 283 696 287
rect 690 282 696 283
rect 768 271 770 303
rect 844 288 846 310
rect 918 308 924 309
rect 918 304 919 308
rect 923 304 924 308
rect 918 303 924 304
rect 1062 308 1068 309
rect 1062 304 1063 308
rect 1067 304 1068 308
rect 1062 303 1068 304
rect 842 287 848 288
rect 842 283 843 287
rect 847 283 848 287
rect 842 282 848 283
rect 920 271 922 303
rect 1064 271 1066 303
rect 1076 288 1078 390
rect 1102 385 1108 386
rect 1102 381 1103 385
rect 1107 381 1108 385
rect 1102 380 1108 381
rect 1206 385 1212 386
rect 1206 381 1207 385
rect 1211 381 1212 385
rect 1206 380 1212 381
rect 1318 385 1324 386
rect 1318 381 1319 385
rect 1323 381 1324 385
rect 1318 380 1324 381
rect 1104 355 1106 380
rect 1208 355 1210 380
rect 1320 355 1322 380
rect 1103 354 1107 355
rect 1103 349 1107 350
rect 1207 354 1211 355
rect 1207 349 1211 350
rect 1319 354 1323 355
rect 1319 349 1323 350
rect 1351 354 1355 355
rect 1351 349 1355 350
rect 1208 328 1210 349
rect 1352 328 1354 349
rect 1206 327 1212 328
rect 1206 323 1207 327
rect 1211 323 1212 327
rect 1206 322 1212 323
rect 1350 327 1356 328
rect 1350 323 1351 327
rect 1355 323 1356 327
rect 1420 324 1422 422
rect 1432 405 1434 429
rect 1430 404 1436 405
rect 1430 400 1431 404
rect 1435 400 1436 404
rect 1430 399 1436 400
rect 1496 396 1498 446
rect 1536 435 1538 471
rect 2008 435 2010 474
rect 2046 472 2047 476
rect 2051 472 2052 476
rect 2046 471 2052 472
rect 2182 475 2188 476
rect 2182 471 2183 475
rect 2187 471 2188 475
rect 2182 470 2188 471
rect 2318 475 2324 476
rect 2318 471 2319 475
rect 2323 471 2324 475
rect 2318 470 2324 471
rect 2462 475 2468 476
rect 2462 471 2463 475
rect 2467 471 2468 475
rect 2462 470 2468 471
rect 2614 475 2620 476
rect 2614 471 2615 475
rect 2619 471 2620 475
rect 2614 470 2620 471
rect 2258 463 2264 464
rect 2046 459 2052 460
rect 2046 455 2047 459
rect 2051 455 2052 459
rect 2258 459 2259 463
rect 2263 459 2264 463
rect 2258 458 2264 459
rect 2394 463 2400 464
rect 2394 459 2395 463
rect 2399 459 2400 463
rect 2394 458 2400 459
rect 2538 463 2544 464
rect 2538 459 2539 463
rect 2543 459 2544 463
rect 2538 458 2544 459
rect 2046 454 2052 455
rect 2182 456 2188 457
rect 1535 434 1539 435
rect 1535 429 1539 430
rect 2007 434 2011 435
rect 2007 429 2011 430
rect 2008 402 2010 429
rect 2048 427 2050 454
rect 2182 452 2183 456
rect 2187 452 2188 456
rect 2182 451 2188 452
rect 2184 427 2186 451
rect 2260 436 2262 458
rect 2318 456 2324 457
rect 2318 452 2319 456
rect 2323 452 2324 456
rect 2318 451 2324 452
rect 2258 435 2264 436
rect 2258 431 2259 435
rect 2263 431 2264 435
rect 2258 430 2264 431
rect 2320 427 2322 451
rect 2396 436 2398 458
rect 2462 456 2468 457
rect 2462 452 2463 456
rect 2467 452 2468 456
rect 2462 451 2468 452
rect 2394 435 2400 436
rect 2394 431 2395 435
rect 2399 431 2400 435
rect 2394 430 2400 431
rect 2464 427 2466 451
rect 2540 436 2542 458
rect 2614 456 2620 457
rect 2614 452 2615 456
rect 2619 452 2620 456
rect 2614 451 2620 452
rect 2538 435 2544 436
rect 2538 431 2539 435
rect 2543 431 2544 435
rect 2538 430 2544 431
rect 2616 427 2618 451
rect 2660 444 2662 534
rect 2686 529 2692 530
rect 2686 525 2687 529
rect 2691 525 2692 529
rect 2686 524 2692 525
rect 2878 529 2884 530
rect 2878 525 2879 529
rect 2883 525 2884 529
rect 2878 524 2884 525
rect 3070 529 3076 530
rect 3070 525 3071 529
rect 3075 525 3076 529
rect 3070 524 3076 525
rect 2688 503 2690 524
rect 2880 503 2882 524
rect 3072 503 3074 524
rect 2687 502 2691 503
rect 2687 497 2691 498
rect 2775 502 2779 503
rect 2775 497 2779 498
rect 2879 502 2883 503
rect 2879 497 2883 498
rect 2959 502 2963 503
rect 2959 497 2963 498
rect 3071 502 3075 503
rect 3071 497 3075 498
rect 3159 502 3163 503
rect 3159 497 3163 498
rect 2776 476 2778 497
rect 2960 476 2962 497
rect 3160 476 3162 497
rect 2774 475 2780 476
rect 2774 471 2775 475
rect 2779 471 2780 475
rect 2774 470 2780 471
rect 2958 475 2964 476
rect 2958 471 2959 475
rect 2963 471 2964 475
rect 2958 470 2964 471
rect 3158 475 3164 476
rect 3158 471 3159 475
rect 3163 471 3164 475
rect 3158 470 3164 471
rect 3236 468 3238 566
rect 3264 549 3266 573
rect 3380 572 3382 614
rect 3392 592 3394 618
rect 3478 612 3484 613
rect 3478 608 3479 612
rect 3483 608 3484 612
rect 3478 607 3484 608
rect 3390 591 3396 592
rect 3390 587 3391 591
rect 3395 587 3396 591
rect 3390 586 3396 587
rect 3480 579 3482 607
rect 3600 592 3602 618
rect 3654 612 3660 613
rect 3654 608 3655 612
rect 3659 608 3660 612
rect 3654 607 3660 608
rect 3598 591 3604 592
rect 3598 587 3599 591
rect 3603 587 3604 591
rect 3598 586 3604 587
rect 3656 579 3658 607
rect 3748 592 3750 698
rect 3838 693 3844 694
rect 3838 689 3839 693
rect 3843 689 3844 693
rect 3838 688 3844 689
rect 3840 659 3842 688
rect 3831 658 3835 659
rect 3831 653 3835 654
rect 3839 658 3843 659
rect 3839 653 3843 654
rect 3832 632 3834 653
rect 3830 631 3836 632
rect 3830 627 3831 631
rect 3835 627 3836 631
rect 3900 628 3902 729
rect 3908 704 3910 746
rect 3944 743 3946 774
rect 3943 742 3947 743
rect 3943 737 3947 738
rect 3944 710 3946 737
rect 3942 709 3948 710
rect 3942 705 3943 709
rect 3947 705 3948 709
rect 3942 704 3948 705
rect 3906 703 3912 704
rect 3906 699 3907 703
rect 3911 699 3912 703
rect 3906 698 3912 699
rect 3942 692 3948 693
rect 3942 688 3943 692
rect 3947 688 3948 692
rect 3942 687 3948 688
rect 3944 659 3946 687
rect 3943 658 3947 659
rect 3943 653 3947 654
rect 3944 633 3946 653
rect 3942 632 3948 633
rect 3942 628 3943 632
rect 3947 628 3948 632
rect 3830 626 3836 627
rect 3898 627 3904 628
rect 3942 627 3948 628
rect 3898 623 3899 627
rect 3903 623 3904 627
rect 3898 622 3904 623
rect 3942 615 3948 616
rect 3830 612 3836 613
rect 3830 608 3831 612
rect 3835 608 3836 612
rect 3942 611 3943 615
rect 3947 611 3948 615
rect 3942 610 3948 611
rect 3830 607 3836 608
rect 3746 591 3752 592
rect 3746 587 3747 591
rect 3751 587 3752 591
rect 3746 586 3752 587
rect 3832 579 3834 607
rect 3906 587 3912 588
rect 3906 583 3907 587
rect 3911 583 3912 587
rect 3906 582 3912 583
rect 3455 578 3459 579
rect 3455 573 3459 574
rect 3479 578 3483 579
rect 3479 573 3483 574
rect 3647 578 3651 579
rect 3647 573 3651 574
rect 3655 578 3659 579
rect 3655 573 3659 574
rect 3831 578 3835 579
rect 3831 573 3835 574
rect 3839 578 3843 579
rect 3839 573 3843 574
rect 3378 571 3384 572
rect 3378 567 3379 571
rect 3383 567 3384 571
rect 3378 566 3384 567
rect 3456 549 3458 573
rect 3530 571 3536 572
rect 3530 567 3531 571
rect 3535 567 3536 571
rect 3530 566 3536 567
rect 3262 548 3268 549
rect 3262 544 3263 548
rect 3267 544 3268 548
rect 3262 543 3268 544
rect 3454 548 3460 549
rect 3454 544 3455 548
rect 3459 544 3460 548
rect 3454 543 3460 544
rect 3532 540 3534 566
rect 3648 549 3650 573
rect 3722 571 3728 572
rect 3722 567 3723 571
rect 3727 567 3728 571
rect 3722 566 3728 567
rect 3646 548 3652 549
rect 3646 544 3647 548
rect 3651 544 3652 548
rect 3646 543 3652 544
rect 3724 540 3726 566
rect 3840 549 3842 573
rect 3838 548 3844 549
rect 3838 544 3839 548
rect 3843 544 3844 548
rect 3838 543 3844 544
rect 3908 540 3910 582
rect 3944 579 3946 610
rect 3943 578 3947 579
rect 3943 573 3947 574
rect 3944 546 3946 573
rect 3942 545 3948 546
rect 3942 541 3943 545
rect 3947 541 3948 545
rect 3942 540 3948 541
rect 3530 539 3536 540
rect 3530 535 3531 539
rect 3535 535 3536 539
rect 3530 534 3536 535
rect 3722 539 3728 540
rect 3722 535 3723 539
rect 3727 535 3728 539
rect 3722 534 3728 535
rect 3906 539 3912 540
rect 3906 535 3907 539
rect 3911 535 3912 539
rect 3906 534 3912 535
rect 3262 529 3268 530
rect 3262 525 3263 529
rect 3267 525 3268 529
rect 3262 524 3268 525
rect 3454 529 3460 530
rect 3454 525 3455 529
rect 3459 525 3460 529
rect 3454 524 3460 525
rect 3646 529 3652 530
rect 3646 525 3647 529
rect 3651 525 3652 529
rect 3646 524 3652 525
rect 3838 529 3844 530
rect 3838 525 3839 529
rect 3843 525 3844 529
rect 3838 524 3844 525
rect 3942 528 3948 529
rect 3942 524 3943 528
rect 3947 524 3948 528
rect 3264 503 3266 524
rect 3456 503 3458 524
rect 3648 503 3650 524
rect 3840 503 3842 524
rect 3942 523 3948 524
rect 3944 503 3946 523
rect 3263 502 3267 503
rect 3263 497 3267 498
rect 3367 502 3371 503
rect 3367 497 3371 498
rect 3455 502 3459 503
rect 3455 497 3459 498
rect 3583 502 3587 503
rect 3583 497 3587 498
rect 3647 502 3651 503
rect 3647 497 3651 498
rect 3807 502 3811 503
rect 3807 497 3811 498
rect 3839 502 3843 503
rect 3839 497 3843 498
rect 3943 502 3947 503
rect 3943 497 3947 498
rect 3368 476 3370 497
rect 3584 476 3586 497
rect 3808 476 3810 497
rect 3944 477 3946 497
rect 3942 476 3948 477
rect 3366 475 3372 476
rect 3366 471 3367 475
rect 3371 471 3372 475
rect 3366 470 3372 471
rect 3582 475 3588 476
rect 3582 471 3583 475
rect 3587 471 3588 475
rect 3582 470 3588 471
rect 3806 475 3812 476
rect 3806 471 3807 475
rect 3811 471 3812 475
rect 3942 472 3943 476
rect 3947 472 3948 476
rect 3942 471 3948 472
rect 3806 470 3812 471
rect 2698 467 2704 468
rect 2690 463 2696 464
rect 2690 459 2691 463
rect 2695 459 2696 463
rect 2698 463 2699 467
rect 2703 463 2704 467
rect 3234 467 3240 468
rect 2698 462 2704 463
rect 3034 463 3040 464
rect 2690 458 2696 459
rect 2658 443 2664 444
rect 2658 439 2659 443
rect 2663 439 2664 443
rect 2658 438 2664 439
rect 2692 436 2694 458
rect 2690 435 2696 436
rect 2690 431 2691 435
rect 2695 431 2696 435
rect 2690 430 2696 431
rect 2700 428 2702 462
rect 3034 459 3035 463
rect 3039 459 3040 463
rect 3234 463 3235 467
rect 3239 463 3240 467
rect 3234 462 3240 463
rect 3242 467 3248 468
rect 3242 463 3243 467
rect 3247 463 3248 467
rect 3242 462 3248 463
rect 3766 467 3772 468
rect 3766 463 3767 467
rect 3771 463 3772 467
rect 3766 462 3772 463
rect 3034 458 3040 459
rect 2774 456 2780 457
rect 2774 452 2775 456
rect 2779 452 2780 456
rect 2774 451 2780 452
rect 2958 456 2964 457
rect 2958 452 2959 456
rect 2963 452 2964 456
rect 2958 451 2964 452
rect 2698 427 2704 428
rect 2776 427 2778 451
rect 2960 427 2962 451
rect 3036 436 3038 458
rect 3158 456 3164 457
rect 3158 452 3159 456
rect 3163 452 3164 456
rect 3158 451 3164 452
rect 3034 435 3040 436
rect 3034 431 3035 435
rect 3039 431 3040 435
rect 3034 430 3040 431
rect 3160 427 3162 451
rect 3244 444 3246 462
rect 3366 456 3372 457
rect 3366 452 3367 456
rect 3371 452 3372 456
rect 3366 451 3372 452
rect 3582 456 3588 457
rect 3582 452 3583 456
rect 3587 452 3588 456
rect 3582 451 3588 452
rect 3242 443 3248 444
rect 3242 439 3243 443
rect 3247 439 3248 443
rect 3242 438 3248 439
rect 3368 427 3370 451
rect 3490 431 3496 432
rect 3490 427 3491 431
rect 3495 427 3496 431
rect 3584 427 3586 451
rect 2047 426 2051 427
rect 2047 421 2051 422
rect 2183 426 2187 427
rect 2183 421 2187 422
rect 2319 426 2323 427
rect 2319 421 2323 422
rect 2343 426 2347 427
rect 2343 421 2347 422
rect 2463 426 2467 427
rect 2463 421 2467 422
rect 2487 426 2491 427
rect 2487 421 2491 422
rect 2615 426 2619 427
rect 2615 421 2619 422
rect 2639 426 2643 427
rect 2698 423 2699 427
rect 2703 423 2704 427
rect 2698 422 2704 423
rect 2775 426 2779 427
rect 2639 421 2643 422
rect 2775 421 2779 422
rect 2799 426 2803 427
rect 2799 421 2803 422
rect 2959 426 2963 427
rect 2959 421 2963 422
rect 3111 426 3115 427
rect 3111 421 3115 422
rect 3159 426 3163 427
rect 3159 421 3163 422
rect 3263 426 3267 427
rect 3263 421 3267 422
rect 3367 426 3371 427
rect 3367 421 3371 422
rect 3415 426 3419 427
rect 3490 426 3496 427
rect 3559 426 3563 427
rect 3415 421 3419 422
rect 2006 401 2012 402
rect 2006 397 2007 401
rect 2011 397 2012 401
rect 2006 396 2012 397
rect 1496 395 1504 396
rect 1496 392 1499 395
rect 1498 391 1499 392
rect 1503 391 1504 395
rect 2048 394 2050 421
rect 2344 397 2346 421
rect 2418 419 2424 420
rect 2418 415 2419 419
rect 2423 415 2424 419
rect 2418 414 2424 415
rect 2342 396 2348 397
rect 1498 390 1504 391
rect 2046 393 2052 394
rect 2046 389 2047 393
rect 2051 389 2052 393
rect 2342 392 2343 396
rect 2347 392 2348 396
rect 2342 391 2348 392
rect 2046 388 2052 389
rect 2420 388 2422 414
rect 2488 397 2490 421
rect 2562 419 2568 420
rect 2562 415 2563 419
rect 2567 415 2568 419
rect 2562 414 2568 415
rect 2486 396 2492 397
rect 2486 392 2487 396
rect 2491 392 2492 396
rect 2486 391 2492 392
rect 2564 388 2566 414
rect 2640 397 2642 421
rect 2714 419 2720 420
rect 2714 415 2715 419
rect 2719 415 2720 419
rect 2714 414 2720 415
rect 2638 396 2644 397
rect 2638 392 2639 396
rect 2643 392 2644 396
rect 2638 391 2644 392
rect 2716 388 2718 414
rect 2800 397 2802 421
rect 2874 419 2880 420
rect 2874 415 2875 419
rect 2879 415 2880 419
rect 2874 414 2880 415
rect 2798 396 2804 397
rect 2798 392 2799 396
rect 2803 392 2804 396
rect 2798 391 2804 392
rect 2876 388 2878 414
rect 2960 397 2962 421
rect 3112 397 3114 421
rect 3186 419 3192 420
rect 3186 415 3187 419
rect 3191 415 3192 419
rect 3186 414 3192 415
rect 2958 396 2964 397
rect 2958 392 2959 396
rect 2963 392 2964 396
rect 2958 391 2964 392
rect 3110 396 3116 397
rect 3110 392 3111 396
rect 3115 392 3116 396
rect 3110 391 3116 392
rect 3188 388 3190 414
rect 3264 397 3266 421
rect 3338 419 3344 420
rect 3338 415 3339 419
rect 3343 415 3344 419
rect 3338 414 3344 415
rect 3262 396 3268 397
rect 3262 392 3263 396
rect 3267 392 3268 396
rect 3262 391 3268 392
rect 3340 388 3342 414
rect 3416 397 3418 421
rect 3414 396 3420 397
rect 3414 392 3415 396
rect 3419 392 3420 396
rect 3414 391 3420 392
rect 3492 388 3494 426
rect 3559 421 3563 422
rect 3583 426 3587 427
rect 3583 421 3587 422
rect 3711 426 3715 427
rect 3711 421 3715 422
rect 3498 411 3504 412
rect 3498 407 3499 411
rect 3503 407 3504 411
rect 3498 406 3504 407
rect 3500 388 3502 406
rect 3560 397 3562 421
rect 3646 419 3652 420
rect 3646 415 3647 419
rect 3651 415 3652 419
rect 3646 414 3652 415
rect 3558 396 3564 397
rect 3558 392 3559 396
rect 3563 392 3564 396
rect 3558 391 3564 392
rect 3648 388 3650 414
rect 3712 397 3714 421
rect 3710 396 3716 397
rect 3710 392 3711 396
rect 3715 392 3716 396
rect 3710 391 3716 392
rect 2418 387 2424 388
rect 1430 385 1436 386
rect 1430 381 1431 385
rect 1435 381 1436 385
rect 1430 380 1436 381
rect 2006 384 2012 385
rect 2006 380 2007 384
rect 2011 380 2012 384
rect 2418 383 2419 387
rect 2423 383 2424 387
rect 2418 382 2424 383
rect 2562 387 2568 388
rect 2562 383 2563 387
rect 2567 383 2568 387
rect 2562 382 2568 383
rect 2714 387 2720 388
rect 2714 383 2715 387
rect 2719 383 2720 387
rect 2714 382 2720 383
rect 2874 387 2880 388
rect 2874 383 2875 387
rect 2879 383 2880 387
rect 2874 382 2880 383
rect 2898 387 2904 388
rect 2898 383 2899 387
rect 2903 383 2904 387
rect 2898 382 2904 383
rect 3186 387 3192 388
rect 3186 383 3187 387
rect 3191 383 3192 387
rect 3186 382 3192 383
rect 3338 387 3344 388
rect 3338 383 3339 387
rect 3343 383 3344 387
rect 3338 382 3344 383
rect 3490 387 3496 388
rect 3490 383 3491 387
rect 3495 383 3496 387
rect 3490 382 3496 383
rect 3498 387 3504 388
rect 3498 383 3499 387
rect 3503 383 3504 387
rect 3498 382 3504 383
rect 3646 387 3652 388
rect 3646 383 3647 387
rect 3651 383 3652 387
rect 3646 382 3652 383
rect 1432 355 1434 380
rect 2006 379 2012 380
rect 2008 355 2010 379
rect 2342 377 2348 378
rect 2046 376 2052 377
rect 2046 372 2047 376
rect 2051 372 2052 376
rect 2342 373 2343 377
rect 2347 373 2348 377
rect 2342 372 2348 373
rect 2486 377 2492 378
rect 2486 373 2487 377
rect 2491 373 2492 377
rect 2486 372 2492 373
rect 2638 377 2644 378
rect 2638 373 2639 377
rect 2643 373 2644 377
rect 2638 372 2644 373
rect 2798 377 2804 378
rect 2798 373 2799 377
rect 2803 373 2804 377
rect 2798 372 2804 373
rect 2046 371 2052 372
rect 1431 354 1435 355
rect 1431 349 1435 350
rect 1495 354 1499 355
rect 1495 349 1499 350
rect 1639 354 1643 355
rect 1639 349 1643 350
rect 2007 354 2011 355
rect 2007 349 2011 350
rect 1496 328 1498 349
rect 1640 328 1642 349
rect 2008 329 2010 349
rect 2048 347 2050 371
rect 2344 347 2346 372
rect 2488 347 2490 372
rect 2640 347 2642 372
rect 2800 347 2802 372
rect 2047 346 2051 347
rect 2047 341 2051 342
rect 2343 346 2347 347
rect 2343 341 2347 342
rect 2487 346 2491 347
rect 2487 341 2491 342
rect 2495 346 2499 347
rect 2495 341 2499 342
rect 2639 346 2643 347
rect 2639 341 2643 342
rect 2799 346 2803 347
rect 2799 341 2803 342
rect 2006 328 2012 329
rect 1494 327 1500 328
rect 1350 322 1356 323
rect 1418 323 1424 324
rect 1418 319 1419 323
rect 1423 319 1424 323
rect 1494 323 1495 327
rect 1499 323 1500 327
rect 1494 322 1500 323
rect 1638 327 1644 328
rect 1638 323 1639 327
rect 1643 323 1644 327
rect 2006 324 2007 328
rect 2011 324 2012 328
rect 2006 323 2012 324
rect 1638 322 1644 323
rect 2048 321 2050 341
rect 2046 320 2052 321
rect 2496 320 2498 341
rect 2640 320 2642 341
rect 2800 320 2802 341
rect 1418 318 1424 319
rect 1434 319 1440 320
rect 1138 315 1144 316
rect 1138 311 1139 315
rect 1143 311 1144 315
rect 1138 310 1144 311
rect 1282 315 1288 316
rect 1282 311 1283 315
rect 1287 311 1288 315
rect 1434 315 1435 319
rect 1439 315 1440 319
rect 1434 314 1440 315
rect 1578 319 1584 320
rect 1578 315 1579 319
rect 1583 315 1584 319
rect 2046 316 2047 320
rect 2051 316 2052 320
rect 2046 315 2052 316
rect 2494 319 2500 320
rect 2494 315 2495 319
rect 2499 315 2500 319
rect 1578 314 1584 315
rect 2494 314 2500 315
rect 2638 319 2644 320
rect 2638 315 2639 319
rect 2643 315 2644 319
rect 2638 314 2644 315
rect 2798 319 2804 320
rect 2798 315 2799 319
rect 2803 315 2804 319
rect 2798 314 2804 315
rect 1282 310 1288 311
rect 1140 288 1142 310
rect 1206 308 1212 309
rect 1206 304 1207 308
rect 1211 304 1212 308
rect 1206 303 1212 304
rect 1074 287 1080 288
rect 1074 283 1075 287
rect 1079 283 1080 287
rect 1074 282 1080 283
rect 1138 287 1144 288
rect 1138 283 1139 287
rect 1143 283 1144 287
rect 1138 282 1144 283
rect 1208 271 1210 303
rect 111 270 115 271
rect 111 265 115 266
rect 167 270 171 271
rect 167 265 171 266
rect 327 270 331 271
rect 327 265 331 266
rect 463 270 467 271
rect 463 265 467 266
rect 503 270 507 271
rect 503 265 507 266
rect 615 270 619 271
rect 615 265 619 266
rect 687 270 691 271
rect 687 265 691 266
rect 767 270 771 271
rect 767 265 771 266
rect 871 270 875 271
rect 871 265 875 266
rect 919 270 923 271
rect 919 265 923 266
rect 1047 270 1051 271
rect 1047 265 1051 266
rect 1063 270 1067 271
rect 1063 265 1067 266
rect 1207 270 1211 271
rect 1207 265 1211 266
rect 1215 270 1219 271
rect 1215 265 1219 266
rect 112 238 114 265
rect 168 241 170 265
rect 242 263 248 264
rect 242 259 243 263
rect 247 259 248 263
rect 242 258 248 259
rect 166 240 172 241
rect 110 237 116 238
rect 110 233 111 237
rect 115 233 116 237
rect 166 236 167 240
rect 171 236 172 240
rect 166 235 172 236
rect 110 232 116 233
rect 244 232 246 258
rect 328 241 330 265
rect 402 263 408 264
rect 402 259 403 263
rect 407 259 408 263
rect 402 258 408 259
rect 326 240 332 241
rect 326 236 327 240
rect 331 236 332 240
rect 326 235 332 236
rect 404 232 406 258
rect 504 241 506 265
rect 578 263 584 264
rect 578 259 579 263
rect 583 259 584 263
rect 578 258 584 259
rect 502 240 508 241
rect 502 236 503 240
rect 507 236 508 240
rect 502 235 508 236
rect 580 232 582 258
rect 688 241 690 265
rect 858 251 864 252
rect 858 247 859 251
rect 863 247 864 251
rect 858 246 864 247
rect 686 240 692 241
rect 686 236 687 240
rect 691 236 692 240
rect 686 235 692 236
rect 242 231 248 232
rect 242 227 243 231
rect 247 227 248 231
rect 242 226 248 227
rect 402 231 408 232
rect 402 227 403 231
rect 407 227 408 231
rect 402 226 408 227
rect 578 231 584 232
rect 578 227 579 231
rect 583 227 584 231
rect 578 226 584 227
rect 166 221 172 222
rect 110 220 116 221
rect 110 216 111 220
rect 115 216 116 220
rect 166 217 167 221
rect 171 217 172 221
rect 166 216 172 217
rect 326 221 332 222
rect 326 217 327 221
rect 331 217 332 221
rect 326 216 332 217
rect 502 221 508 222
rect 502 217 503 221
rect 507 217 508 221
rect 502 216 508 217
rect 686 221 692 222
rect 686 217 687 221
rect 691 217 692 221
rect 686 216 692 217
rect 110 215 116 216
rect 112 167 114 215
rect 168 167 170 216
rect 328 167 330 216
rect 504 167 506 216
rect 688 167 690 216
rect 111 166 115 167
rect 111 161 115 162
rect 135 166 139 167
rect 135 161 139 162
rect 167 166 171 167
rect 167 161 171 162
rect 231 166 235 167
rect 231 161 235 162
rect 327 166 331 167
rect 327 161 331 162
rect 423 166 427 167
rect 423 161 427 162
rect 503 166 507 167
rect 503 161 507 162
rect 527 166 531 167
rect 527 161 531 162
rect 647 166 651 167
rect 647 161 651 162
rect 687 166 691 167
rect 687 161 691 162
rect 775 166 779 167
rect 775 161 779 162
rect 112 141 114 161
rect 110 140 116 141
rect 136 140 138 161
rect 232 140 234 161
rect 328 140 330 161
rect 424 140 426 161
rect 528 140 530 161
rect 648 140 650 161
rect 776 140 778 161
rect 110 136 111 140
rect 115 136 116 140
rect 110 135 116 136
rect 134 139 140 140
rect 134 135 135 139
rect 139 135 140 139
rect 134 134 140 135
rect 230 139 236 140
rect 230 135 231 139
rect 235 135 236 139
rect 230 134 236 135
rect 326 139 332 140
rect 326 135 327 139
rect 331 135 332 139
rect 326 134 332 135
rect 422 139 428 140
rect 422 135 423 139
rect 427 135 428 139
rect 422 134 428 135
rect 526 139 532 140
rect 526 135 527 139
rect 531 135 532 139
rect 526 134 532 135
rect 646 139 652 140
rect 646 135 647 139
rect 651 135 652 139
rect 646 134 652 135
rect 774 139 780 140
rect 774 135 775 139
rect 779 135 780 139
rect 774 134 780 135
rect 860 132 862 246
rect 872 241 874 265
rect 1048 241 1050 265
rect 1216 241 1218 265
rect 1284 264 1286 310
rect 1350 308 1356 309
rect 1350 304 1351 308
rect 1355 304 1356 308
rect 1350 303 1356 304
rect 1352 271 1354 303
rect 1436 288 1438 314
rect 1494 308 1500 309
rect 1494 304 1495 308
rect 1499 304 1500 308
rect 1494 303 1500 304
rect 1434 287 1440 288
rect 1434 283 1435 287
rect 1439 283 1440 287
rect 1434 282 1440 283
rect 1496 271 1498 303
rect 1580 288 1582 314
rect 2006 311 2012 312
rect 1638 308 1644 309
rect 1638 304 1639 308
rect 1643 304 1644 308
rect 2006 307 2007 311
rect 2011 307 2012 311
rect 2006 306 2012 307
rect 2570 307 2576 308
rect 1638 303 1644 304
rect 1578 287 1584 288
rect 1578 283 1579 287
rect 1583 283 1584 287
rect 1578 282 1584 283
rect 1586 283 1592 284
rect 1586 279 1587 283
rect 1591 279 1592 283
rect 1586 278 1592 279
rect 1351 270 1355 271
rect 1351 265 1355 266
rect 1367 270 1371 271
rect 1367 265 1371 266
rect 1495 270 1499 271
rect 1495 265 1499 266
rect 1511 270 1515 271
rect 1511 265 1515 266
rect 1282 263 1288 264
rect 1282 259 1283 263
rect 1287 259 1288 263
rect 1282 258 1288 259
rect 1290 263 1296 264
rect 1290 259 1291 263
rect 1295 259 1296 263
rect 1290 258 1296 259
rect 870 240 876 241
rect 870 236 871 240
rect 875 236 876 240
rect 870 235 876 236
rect 1046 240 1052 241
rect 1046 236 1047 240
rect 1051 236 1052 240
rect 1046 235 1052 236
rect 1214 240 1220 241
rect 1214 236 1215 240
rect 1219 236 1220 240
rect 1214 235 1220 236
rect 1292 232 1294 258
rect 1338 255 1344 256
rect 1338 251 1339 255
rect 1343 251 1344 255
rect 1338 250 1344 251
rect 1340 232 1342 250
rect 1368 241 1370 265
rect 1512 241 1514 265
rect 1366 240 1372 241
rect 1366 236 1367 240
rect 1371 236 1372 240
rect 1366 235 1372 236
rect 1510 240 1516 241
rect 1510 236 1511 240
rect 1515 236 1516 240
rect 1510 235 1516 236
rect 1588 232 1590 278
rect 1640 271 1642 303
rect 2008 271 2010 306
rect 2046 303 2052 304
rect 2046 299 2047 303
rect 2051 299 2052 303
rect 2570 303 2571 307
rect 2575 303 2576 307
rect 2570 302 2576 303
rect 2714 307 2720 308
rect 2714 303 2715 307
rect 2719 303 2720 307
rect 2714 302 2720 303
rect 2874 307 2880 308
rect 2874 303 2875 307
rect 2879 303 2880 307
rect 2874 302 2880 303
rect 2046 298 2052 299
rect 2494 300 2500 301
rect 2048 271 2050 298
rect 2494 296 2495 300
rect 2499 296 2500 300
rect 2494 295 2500 296
rect 2496 271 2498 295
rect 2551 284 2555 285
rect 2572 280 2574 302
rect 2638 300 2644 301
rect 2638 296 2639 300
rect 2643 296 2644 300
rect 2638 295 2644 296
rect 2550 279 2556 280
rect 2550 275 2551 279
rect 2555 275 2556 279
rect 2550 274 2556 275
rect 2570 279 2576 280
rect 2570 275 2571 279
rect 2575 275 2576 279
rect 2570 274 2576 275
rect 2640 271 2642 295
rect 2716 280 2718 302
rect 2798 300 2804 301
rect 2798 296 2799 300
rect 2803 296 2804 300
rect 2798 295 2804 296
rect 2714 279 2720 280
rect 2714 275 2715 279
rect 2719 275 2720 279
rect 2714 274 2720 275
rect 2800 271 2802 295
rect 2876 280 2878 302
rect 2900 285 2902 382
rect 2958 377 2964 378
rect 2958 373 2959 377
rect 2963 373 2964 377
rect 2958 372 2964 373
rect 3110 377 3116 378
rect 3110 373 3111 377
rect 3115 373 3116 377
rect 3110 372 3116 373
rect 3262 377 3268 378
rect 3262 373 3263 377
rect 3267 373 3268 377
rect 3262 372 3268 373
rect 3414 377 3420 378
rect 3414 373 3415 377
rect 3419 373 3420 377
rect 3414 372 3420 373
rect 3558 377 3564 378
rect 3558 373 3559 377
rect 3563 373 3564 377
rect 3558 372 3564 373
rect 3710 377 3716 378
rect 3710 373 3711 377
rect 3715 373 3716 377
rect 3710 372 3716 373
rect 2960 347 2962 372
rect 3112 347 3114 372
rect 3264 347 3266 372
rect 3416 347 3418 372
rect 3560 347 3562 372
rect 3712 347 3714 372
rect 2959 346 2963 347
rect 2959 341 2963 342
rect 3111 346 3115 347
rect 3111 341 3115 342
rect 3119 346 3123 347
rect 3119 341 3123 342
rect 3263 346 3267 347
rect 3263 341 3267 342
rect 3271 346 3275 347
rect 3271 341 3275 342
rect 3415 346 3419 347
rect 3415 341 3419 342
rect 3423 346 3427 347
rect 3423 341 3427 342
rect 3559 346 3563 347
rect 3559 341 3563 342
rect 3567 346 3571 347
rect 3567 341 3571 342
rect 3711 346 3715 347
rect 3711 341 3715 342
rect 2960 320 2962 341
rect 3120 320 3122 341
rect 3272 320 3274 341
rect 3424 320 3426 341
rect 3568 320 3570 341
rect 3712 320 3714 341
rect 2958 319 2964 320
rect 2958 315 2959 319
rect 2963 315 2964 319
rect 2958 314 2964 315
rect 3118 319 3124 320
rect 3118 315 3119 319
rect 3123 315 3124 319
rect 3118 314 3124 315
rect 3270 319 3276 320
rect 3270 315 3271 319
rect 3275 315 3276 319
rect 3270 314 3276 315
rect 3422 319 3428 320
rect 3422 315 3423 319
rect 3427 315 3428 319
rect 3422 314 3428 315
rect 3566 319 3572 320
rect 3566 315 3567 319
rect 3571 315 3572 319
rect 3566 314 3572 315
rect 3710 319 3716 320
rect 3710 315 3711 319
rect 3715 315 3716 319
rect 3710 314 3716 315
rect 3042 311 3048 312
rect 3034 307 3040 308
rect 3034 303 3035 307
rect 3039 303 3040 307
rect 3042 307 3043 311
rect 3047 307 3048 311
rect 3042 306 3048 307
rect 3346 307 3352 308
rect 3034 302 3040 303
rect 2958 300 2964 301
rect 2958 296 2959 300
rect 2963 296 2964 300
rect 2958 295 2964 296
rect 2899 284 2903 285
rect 2874 279 2880 280
rect 2899 279 2903 280
rect 2874 275 2875 279
rect 2879 275 2880 279
rect 2874 274 2880 275
rect 2960 271 2962 295
rect 3036 280 3038 302
rect 3034 279 3040 280
rect 3034 275 3035 279
rect 3039 275 3040 279
rect 3034 274 3040 275
rect 1639 270 1643 271
rect 1639 265 1643 266
rect 1647 270 1651 271
rect 1647 265 1651 266
rect 1783 270 1787 271
rect 1783 265 1787 266
rect 1903 270 1907 271
rect 1903 265 1907 266
rect 2007 270 2011 271
rect 2007 265 2011 266
rect 2047 270 2051 271
rect 2047 265 2051 266
rect 2071 270 2075 271
rect 2071 265 2075 266
rect 2271 270 2275 271
rect 2271 265 2275 266
rect 2495 270 2499 271
rect 2495 265 2499 266
rect 2639 270 2643 271
rect 2639 265 2643 266
rect 2703 270 2707 271
rect 2703 265 2707 266
rect 2799 270 2803 271
rect 2799 265 2803 266
rect 2903 270 2907 271
rect 2903 265 2907 266
rect 2959 270 2963 271
rect 2959 265 2963 266
rect 1594 263 1600 264
rect 1594 259 1595 263
rect 1599 259 1600 263
rect 1594 258 1600 259
rect 1596 232 1598 258
rect 1648 241 1650 265
rect 1730 263 1736 264
rect 1730 259 1731 263
rect 1735 259 1736 263
rect 1730 258 1736 259
rect 1646 240 1652 241
rect 1646 236 1647 240
rect 1651 236 1652 240
rect 1646 235 1652 236
rect 1732 232 1734 258
rect 1784 241 1786 265
rect 1866 263 1872 264
rect 1866 259 1867 263
rect 1871 259 1872 263
rect 1866 258 1872 259
rect 1782 240 1788 241
rect 1782 236 1783 240
rect 1787 236 1788 240
rect 1782 235 1788 236
rect 1868 232 1870 258
rect 1904 241 1906 265
rect 1986 263 1992 264
rect 1986 259 1987 263
rect 1991 259 1992 263
rect 1986 258 1992 259
rect 1902 240 1908 241
rect 1902 236 1903 240
rect 1907 236 1908 240
rect 1902 235 1908 236
rect 1988 232 1990 258
rect 2008 238 2010 265
rect 2048 238 2050 265
rect 2072 241 2074 265
rect 2154 263 2160 264
rect 2154 259 2155 263
rect 2159 259 2160 263
rect 2154 258 2160 259
rect 2070 240 2076 241
rect 2006 237 2012 238
rect 2006 233 2007 237
rect 2011 233 2012 237
rect 2006 232 2012 233
rect 2046 237 2052 238
rect 2046 233 2047 237
rect 2051 233 2052 237
rect 2070 236 2071 240
rect 2075 236 2076 240
rect 2070 235 2076 236
rect 2046 232 2052 233
rect 2156 232 2158 258
rect 2272 241 2274 265
rect 2496 241 2498 265
rect 2538 263 2544 264
rect 2538 259 2539 263
rect 2543 259 2544 263
rect 2538 258 2544 259
rect 2578 263 2584 264
rect 2578 259 2579 263
rect 2583 259 2584 263
rect 2578 258 2584 259
rect 2270 240 2276 241
rect 2270 236 2271 240
rect 2275 236 2276 240
rect 2270 235 2276 236
rect 2494 240 2500 241
rect 2494 236 2495 240
rect 2499 236 2500 240
rect 2494 235 2500 236
rect 1114 231 1120 232
rect 1114 227 1115 231
rect 1119 227 1120 231
rect 1114 226 1120 227
rect 1290 231 1296 232
rect 1290 227 1291 231
rect 1295 227 1296 231
rect 1290 226 1296 227
rect 1338 231 1344 232
rect 1338 227 1339 231
rect 1343 227 1344 231
rect 1338 226 1344 227
rect 1586 231 1592 232
rect 1586 227 1587 231
rect 1591 227 1592 231
rect 1586 226 1592 227
rect 1594 231 1600 232
rect 1594 227 1595 231
rect 1599 227 1600 231
rect 1594 226 1600 227
rect 1730 231 1736 232
rect 1730 227 1731 231
rect 1735 227 1736 231
rect 1730 226 1736 227
rect 1866 231 1872 232
rect 1866 227 1867 231
rect 1871 227 1872 231
rect 1866 226 1872 227
rect 1986 231 1992 232
rect 1986 227 1987 231
rect 1991 227 1992 231
rect 1986 226 1992 227
rect 2154 231 2160 232
rect 2154 227 2155 231
rect 2159 227 2160 231
rect 2154 226 2160 227
rect 870 221 876 222
rect 870 217 871 221
rect 875 217 876 221
rect 870 216 876 217
rect 1046 221 1052 222
rect 1046 217 1047 221
rect 1051 217 1052 221
rect 1046 216 1052 217
rect 872 167 874 216
rect 1048 167 1050 216
rect 871 166 875 167
rect 871 161 875 162
rect 903 166 907 167
rect 903 161 907 162
rect 1031 166 1035 167
rect 1031 161 1035 162
rect 1047 166 1051 167
rect 1047 161 1051 162
rect 904 140 906 161
rect 1032 140 1034 161
rect 902 139 908 140
rect 902 135 903 139
rect 907 135 908 139
rect 902 134 908 135
rect 1030 139 1036 140
rect 1030 135 1031 139
rect 1035 135 1036 139
rect 1030 134 1036 135
rect 858 131 864 132
rect 210 127 216 128
rect 110 123 116 124
rect 110 119 111 123
rect 115 119 116 123
rect 210 123 211 127
rect 215 123 216 127
rect 210 122 216 123
rect 306 127 312 128
rect 306 123 307 127
rect 311 123 312 127
rect 306 122 312 123
rect 402 127 408 128
rect 402 123 403 127
rect 407 123 408 127
rect 402 122 408 123
rect 498 127 504 128
rect 498 123 499 127
rect 503 123 504 127
rect 498 122 504 123
rect 602 127 608 128
rect 602 123 603 127
rect 607 123 608 127
rect 602 122 608 123
rect 722 127 728 128
rect 722 123 723 127
rect 727 123 728 127
rect 722 122 728 123
rect 850 127 856 128
rect 850 123 851 127
rect 855 123 856 127
rect 858 127 859 131
rect 863 127 864 131
rect 858 126 864 127
rect 850 122 856 123
rect 110 118 116 119
rect 134 120 140 121
rect 112 91 114 118
rect 134 116 135 120
rect 139 116 140 120
rect 134 115 140 116
rect 136 91 138 115
rect 212 100 214 122
rect 230 120 236 121
rect 230 116 231 120
rect 235 116 236 120
rect 230 115 236 116
rect 210 99 216 100
rect 210 95 211 99
rect 215 95 216 99
rect 210 94 216 95
rect 232 91 234 115
rect 308 100 310 122
rect 326 120 332 121
rect 326 116 327 120
rect 331 116 332 120
rect 326 115 332 116
rect 306 99 312 100
rect 306 95 307 99
rect 311 95 312 99
rect 306 94 312 95
rect 328 91 330 115
rect 404 100 406 122
rect 422 120 428 121
rect 422 116 423 120
rect 427 116 428 120
rect 422 115 428 116
rect 402 99 408 100
rect 402 95 403 99
rect 407 95 408 99
rect 402 94 408 95
rect 424 91 426 115
rect 500 100 502 122
rect 526 120 532 121
rect 526 116 527 120
rect 531 116 532 120
rect 526 115 532 116
rect 498 99 504 100
rect 498 95 499 99
rect 503 95 504 99
rect 498 94 504 95
rect 528 91 530 115
rect 604 100 606 122
rect 646 120 652 121
rect 646 116 647 120
rect 651 116 652 120
rect 646 115 652 116
rect 602 99 608 100
rect 602 95 603 99
rect 607 95 608 99
rect 602 94 608 95
rect 648 91 650 115
rect 724 100 726 122
rect 774 120 780 121
rect 774 116 775 120
rect 779 116 780 120
rect 774 115 780 116
rect 722 99 728 100
rect 722 95 723 99
rect 727 95 728 99
rect 722 94 728 95
rect 776 91 778 115
rect 852 100 854 122
rect 902 120 908 121
rect 902 116 903 120
rect 907 116 908 120
rect 902 115 908 116
rect 1030 120 1036 121
rect 1030 116 1031 120
rect 1035 116 1036 120
rect 1030 115 1036 116
rect 850 99 856 100
rect 850 95 851 99
rect 855 95 856 99
rect 850 94 856 95
rect 904 91 906 115
rect 1032 91 1034 115
rect 1116 100 1118 226
rect 1214 221 1220 222
rect 1214 217 1215 221
rect 1219 217 1220 221
rect 1214 216 1220 217
rect 1366 221 1372 222
rect 1366 217 1367 221
rect 1371 217 1372 221
rect 1366 216 1372 217
rect 1510 221 1516 222
rect 1510 217 1511 221
rect 1515 217 1516 221
rect 1510 216 1516 217
rect 1646 221 1652 222
rect 1646 217 1647 221
rect 1651 217 1652 221
rect 1646 216 1652 217
rect 1782 221 1788 222
rect 1782 217 1783 221
rect 1787 217 1788 221
rect 1782 216 1788 217
rect 1902 221 1908 222
rect 2070 221 2076 222
rect 1902 217 1903 221
rect 1907 217 1908 221
rect 1902 216 1908 217
rect 2006 220 2012 221
rect 2006 216 2007 220
rect 2011 216 2012 220
rect 1216 167 1218 216
rect 1368 167 1370 216
rect 1512 167 1514 216
rect 1648 167 1650 216
rect 1784 167 1786 216
rect 1904 167 1906 216
rect 2006 215 2012 216
rect 2046 220 2052 221
rect 2046 216 2047 220
rect 2051 216 2052 220
rect 2070 217 2071 221
rect 2075 217 2076 221
rect 2070 216 2076 217
rect 2270 221 2276 222
rect 2270 217 2271 221
rect 2275 217 2276 221
rect 2270 216 2276 217
rect 2494 221 2500 222
rect 2494 217 2495 221
rect 2499 217 2500 221
rect 2494 216 2500 217
rect 2046 215 2052 216
rect 2008 167 2010 215
rect 2048 171 2050 215
rect 2072 171 2074 216
rect 2272 171 2274 216
rect 2496 171 2498 216
rect 2047 170 2051 171
rect 1151 166 1155 167
rect 1151 161 1155 162
rect 1215 166 1219 167
rect 1215 161 1219 162
rect 1271 166 1275 167
rect 1271 161 1275 162
rect 1367 166 1371 167
rect 1367 161 1371 162
rect 1383 166 1387 167
rect 1383 161 1387 162
rect 1487 166 1491 167
rect 1487 161 1491 162
rect 1511 166 1515 167
rect 1511 161 1515 162
rect 1591 166 1595 167
rect 1591 161 1595 162
rect 1647 166 1651 167
rect 1647 161 1651 162
rect 1703 166 1707 167
rect 1703 161 1707 162
rect 1783 166 1787 167
rect 1783 161 1787 162
rect 1807 166 1811 167
rect 1807 161 1811 162
rect 1903 166 1907 167
rect 1903 161 1907 162
rect 2007 166 2011 167
rect 2047 165 2051 166
rect 2071 170 2075 171
rect 2071 165 2075 166
rect 2167 170 2171 171
rect 2167 165 2171 166
rect 2263 170 2267 171
rect 2263 165 2267 166
rect 2271 170 2275 171
rect 2271 165 2275 166
rect 2359 170 2363 171
rect 2359 165 2363 166
rect 2455 170 2459 171
rect 2455 165 2459 166
rect 2495 170 2499 171
rect 2495 165 2499 166
rect 2007 161 2011 162
rect 1152 140 1154 161
rect 1272 140 1274 161
rect 1384 140 1386 161
rect 1488 140 1490 161
rect 1592 140 1594 161
rect 1704 140 1706 161
rect 1808 140 1810 161
rect 1904 140 1906 161
rect 2008 141 2010 161
rect 2048 145 2050 165
rect 2046 144 2052 145
rect 2072 144 2074 165
rect 2168 144 2170 165
rect 2264 144 2266 165
rect 2360 144 2362 165
rect 2456 144 2458 165
rect 2006 140 2012 141
rect 1150 139 1156 140
rect 1150 135 1151 139
rect 1155 135 1156 139
rect 1150 134 1156 135
rect 1270 139 1276 140
rect 1270 135 1271 139
rect 1275 135 1276 139
rect 1270 134 1276 135
rect 1382 139 1388 140
rect 1382 135 1383 139
rect 1387 135 1388 139
rect 1382 134 1388 135
rect 1486 139 1492 140
rect 1486 135 1487 139
rect 1491 135 1492 139
rect 1486 134 1492 135
rect 1590 139 1596 140
rect 1590 135 1591 139
rect 1595 135 1596 139
rect 1590 134 1596 135
rect 1702 139 1708 140
rect 1702 135 1703 139
rect 1707 135 1708 139
rect 1702 134 1708 135
rect 1806 139 1812 140
rect 1806 135 1807 139
rect 1811 135 1812 139
rect 1806 134 1812 135
rect 1902 139 1908 140
rect 1902 135 1903 139
rect 1907 135 1908 139
rect 2006 136 2007 140
rect 2011 136 2012 140
rect 2046 140 2047 144
rect 2051 140 2052 144
rect 2046 139 2052 140
rect 2070 143 2076 144
rect 2070 139 2071 143
rect 2075 139 2076 143
rect 2070 138 2076 139
rect 2166 143 2172 144
rect 2166 139 2167 143
rect 2171 139 2172 143
rect 2166 138 2172 139
rect 2262 143 2268 144
rect 2262 139 2263 143
rect 2267 139 2268 143
rect 2262 138 2268 139
rect 2358 143 2364 144
rect 2358 139 2359 143
rect 2363 139 2364 143
rect 2358 138 2364 139
rect 2454 143 2460 144
rect 2454 139 2455 143
rect 2459 139 2460 143
rect 2454 138 2460 139
rect 2540 136 2542 258
rect 2580 232 2582 258
rect 2704 241 2706 265
rect 2904 241 2906 265
rect 3044 264 3046 306
rect 3346 303 3347 307
rect 3351 303 3352 307
rect 3346 302 3352 303
rect 3498 307 3504 308
rect 3498 303 3499 307
rect 3503 303 3504 307
rect 3498 302 3504 303
rect 3642 307 3648 308
rect 3642 303 3643 307
rect 3647 303 3648 307
rect 3642 302 3648 303
rect 3118 300 3124 301
rect 3118 296 3119 300
rect 3123 296 3124 300
rect 3118 295 3124 296
rect 3270 300 3276 301
rect 3270 296 3271 300
rect 3275 296 3276 300
rect 3270 295 3276 296
rect 3120 271 3122 295
rect 3272 271 3274 295
rect 3348 280 3350 302
rect 3422 300 3428 301
rect 3422 296 3423 300
rect 3427 296 3428 300
rect 3422 295 3428 296
rect 3346 279 3352 280
rect 3346 275 3347 279
rect 3351 275 3352 279
rect 3346 274 3352 275
rect 3424 271 3426 295
rect 3500 280 3502 302
rect 3566 300 3572 301
rect 3566 296 3567 300
rect 3571 296 3572 300
rect 3566 295 3572 296
rect 3498 279 3504 280
rect 3498 275 3499 279
rect 3503 275 3504 279
rect 3498 274 3504 275
rect 3568 271 3570 295
rect 3618 271 3624 272
rect 3095 270 3099 271
rect 3095 265 3099 266
rect 3119 270 3123 271
rect 3119 265 3123 266
rect 3271 270 3275 271
rect 3271 265 3275 266
rect 3287 270 3291 271
rect 3287 265 3291 266
rect 3423 270 3427 271
rect 3423 265 3427 266
rect 3479 270 3483 271
rect 3479 265 3483 266
rect 3567 270 3571 271
rect 3618 267 3619 271
rect 3623 267 3624 271
rect 3618 266 3624 267
rect 3567 265 3571 266
rect 3042 263 3048 264
rect 3042 259 3043 263
rect 3047 259 3048 263
rect 3042 258 3048 259
rect 3096 241 3098 265
rect 3170 263 3176 264
rect 3170 259 3171 263
rect 3175 259 3176 263
rect 3170 258 3176 259
rect 2702 240 2708 241
rect 2702 236 2703 240
rect 2707 236 2708 240
rect 2702 235 2708 236
rect 2902 240 2908 241
rect 2902 236 2903 240
rect 2907 236 2908 240
rect 2902 235 2908 236
rect 3094 240 3100 241
rect 3094 236 3095 240
rect 3099 236 3100 240
rect 3094 235 3100 236
rect 3172 232 3174 258
rect 3288 241 3290 265
rect 3362 263 3368 264
rect 3362 259 3363 263
rect 3367 259 3368 263
rect 3362 258 3368 259
rect 3286 240 3292 241
rect 3286 236 3287 240
rect 3291 236 3292 240
rect 3286 235 3292 236
rect 3364 232 3366 258
rect 3480 241 3482 265
rect 3554 263 3560 264
rect 3554 259 3555 263
rect 3559 259 3560 263
rect 3554 258 3560 259
rect 3498 255 3504 256
rect 3498 251 3499 255
rect 3503 251 3504 255
rect 3498 250 3504 251
rect 3478 240 3484 241
rect 3478 236 3479 240
rect 3483 236 3484 240
rect 3478 235 3484 236
rect 2578 231 2584 232
rect 2578 227 2579 231
rect 2583 227 2584 231
rect 2578 226 2584 227
rect 3170 231 3176 232
rect 3170 227 3171 231
rect 3175 227 3176 231
rect 3170 226 3176 227
rect 3362 231 3368 232
rect 3362 227 3363 231
rect 3367 227 3368 231
rect 3362 226 3368 227
rect 2614 223 2620 224
rect 2614 219 2615 223
rect 2619 219 2620 223
rect 2614 218 2620 219
rect 2702 221 2708 222
rect 2551 170 2555 171
rect 2551 165 2555 166
rect 2552 144 2554 165
rect 2550 143 2556 144
rect 2550 139 2551 143
rect 2555 139 2556 143
rect 2550 138 2556 139
rect 2006 135 2012 136
rect 2538 135 2544 136
rect 1902 134 1908 135
rect 2146 131 2152 132
rect 1122 127 1128 128
rect 1122 123 1123 127
rect 1127 123 1128 127
rect 1122 122 1128 123
rect 1226 127 1232 128
rect 1226 123 1227 127
rect 1231 123 1232 127
rect 1226 122 1232 123
rect 1346 127 1352 128
rect 1346 123 1347 127
rect 1351 123 1352 127
rect 1346 122 1352 123
rect 1458 127 1464 128
rect 1458 123 1459 127
rect 1463 123 1464 127
rect 1458 122 1464 123
rect 1562 127 1568 128
rect 1562 123 1563 127
rect 1567 123 1568 127
rect 1562 122 1568 123
rect 1666 127 1672 128
rect 1666 123 1667 127
rect 1671 123 1672 127
rect 1666 122 1672 123
rect 1778 127 1784 128
rect 1778 123 1779 127
rect 1783 123 1784 127
rect 1778 122 1784 123
rect 1882 127 1888 128
rect 1882 123 1883 127
rect 1887 123 1888 127
rect 1882 122 1888 123
rect 1978 127 1984 128
rect 1978 123 1979 127
rect 1983 123 1984 127
rect 2046 127 2052 128
rect 1978 122 1984 123
rect 2006 123 2012 124
rect 1124 100 1126 122
rect 1150 120 1156 121
rect 1150 116 1151 120
rect 1155 116 1156 120
rect 1150 115 1156 116
rect 1114 99 1120 100
rect 1114 95 1115 99
rect 1119 95 1120 99
rect 1114 94 1120 95
rect 1122 99 1128 100
rect 1122 95 1123 99
rect 1127 95 1128 99
rect 1122 94 1128 95
rect 1152 91 1154 115
rect 1228 100 1230 122
rect 1270 120 1276 121
rect 1270 116 1271 120
rect 1275 116 1276 120
rect 1270 115 1276 116
rect 1226 99 1232 100
rect 1226 95 1227 99
rect 1231 95 1232 99
rect 1226 94 1232 95
rect 1272 91 1274 115
rect 1348 100 1350 122
rect 1382 120 1388 121
rect 1382 116 1383 120
rect 1387 116 1388 120
rect 1382 115 1388 116
rect 1346 99 1352 100
rect 1346 95 1347 99
rect 1351 95 1352 99
rect 1346 94 1352 95
rect 1384 91 1386 115
rect 1460 100 1462 122
rect 1486 120 1492 121
rect 1486 116 1487 120
rect 1491 116 1492 120
rect 1486 115 1492 116
rect 1458 99 1464 100
rect 1458 95 1459 99
rect 1463 95 1464 99
rect 1458 94 1464 95
rect 1488 91 1490 115
rect 1564 100 1566 122
rect 1590 120 1596 121
rect 1590 116 1591 120
rect 1595 116 1596 120
rect 1590 115 1596 116
rect 1562 99 1568 100
rect 1562 95 1563 99
rect 1567 95 1568 99
rect 1562 94 1568 95
rect 1592 91 1594 115
rect 1668 100 1670 122
rect 1702 120 1708 121
rect 1702 116 1703 120
rect 1707 116 1708 120
rect 1702 115 1708 116
rect 1666 99 1672 100
rect 1666 95 1667 99
rect 1671 95 1672 99
rect 1666 94 1672 95
rect 1704 91 1706 115
rect 1780 100 1782 122
rect 1806 120 1812 121
rect 1806 116 1807 120
rect 1811 116 1812 120
rect 1806 115 1812 116
rect 1778 99 1784 100
rect 1778 95 1779 99
rect 1783 95 1784 99
rect 1778 94 1784 95
rect 1808 91 1810 115
rect 1884 100 1886 122
rect 1902 120 1908 121
rect 1902 116 1903 120
rect 1907 116 1908 120
rect 1902 115 1908 116
rect 1882 99 1888 100
rect 1882 95 1883 99
rect 1887 95 1888 99
rect 1882 94 1888 95
rect 1904 91 1906 115
rect 1980 104 1982 122
rect 2006 119 2007 123
rect 2011 119 2012 123
rect 2046 123 2047 127
rect 2051 123 2052 127
rect 2146 127 2147 131
rect 2151 127 2152 131
rect 2146 126 2152 127
rect 2242 131 2248 132
rect 2242 127 2243 131
rect 2247 127 2248 131
rect 2242 126 2248 127
rect 2338 131 2344 132
rect 2338 127 2339 131
rect 2343 127 2344 131
rect 2338 126 2344 127
rect 2434 131 2440 132
rect 2434 127 2435 131
rect 2439 127 2440 131
rect 2434 126 2440 127
rect 2530 131 2536 132
rect 2530 127 2531 131
rect 2535 127 2536 131
rect 2538 131 2539 135
rect 2543 131 2544 135
rect 2538 130 2544 131
rect 2530 126 2536 127
rect 2046 122 2052 123
rect 2070 124 2076 125
rect 2006 118 2012 119
rect 1978 103 1984 104
rect 1978 99 1979 103
rect 1983 99 1984 103
rect 1978 98 1984 99
rect 2008 91 2010 118
rect 2048 95 2050 122
rect 2070 120 2071 124
rect 2075 120 2076 124
rect 2070 119 2076 120
rect 2072 95 2074 119
rect 2148 104 2150 126
rect 2166 124 2172 125
rect 2166 120 2167 124
rect 2171 120 2172 124
rect 2166 119 2172 120
rect 2146 103 2152 104
rect 2146 99 2147 103
rect 2151 99 2152 103
rect 2146 98 2152 99
rect 2168 95 2170 119
rect 2244 104 2246 126
rect 2262 124 2268 125
rect 2262 120 2263 124
rect 2267 120 2268 124
rect 2262 119 2268 120
rect 2242 103 2248 104
rect 2242 99 2243 103
rect 2247 99 2248 103
rect 2242 98 2248 99
rect 2264 95 2266 119
rect 2340 104 2342 126
rect 2358 124 2364 125
rect 2358 120 2359 124
rect 2363 120 2364 124
rect 2358 119 2364 120
rect 2338 103 2344 104
rect 2338 99 2339 103
rect 2343 99 2344 103
rect 2338 98 2344 99
rect 2360 95 2362 119
rect 2436 104 2438 126
rect 2454 124 2460 125
rect 2454 120 2455 124
rect 2459 120 2460 124
rect 2454 119 2460 120
rect 2434 103 2440 104
rect 2434 99 2435 103
rect 2439 99 2440 103
rect 2434 98 2440 99
rect 2456 95 2458 119
rect 2532 104 2534 126
rect 2550 124 2556 125
rect 2550 120 2551 124
rect 2555 120 2556 124
rect 2550 119 2556 120
rect 2530 103 2536 104
rect 2530 99 2531 103
rect 2535 99 2536 103
rect 2530 98 2536 99
rect 2552 95 2554 119
rect 2616 104 2618 218
rect 2702 217 2703 221
rect 2707 217 2708 221
rect 2702 216 2708 217
rect 2902 221 2908 222
rect 2902 217 2903 221
rect 2907 217 2908 221
rect 2902 216 2908 217
rect 3094 221 3100 222
rect 3094 217 3095 221
rect 3099 217 3100 221
rect 3094 216 3100 217
rect 3286 221 3292 222
rect 3286 217 3287 221
rect 3291 217 3292 221
rect 3286 216 3292 217
rect 3478 221 3484 222
rect 3478 217 3479 221
rect 3483 217 3484 221
rect 3478 216 3484 217
rect 2704 171 2706 216
rect 2904 171 2906 216
rect 3096 171 3098 216
rect 3288 171 3290 216
rect 3480 171 3482 216
rect 2655 170 2659 171
rect 2655 165 2659 166
rect 2703 170 2707 171
rect 2703 165 2707 166
rect 2759 170 2763 171
rect 2759 165 2763 166
rect 2863 170 2867 171
rect 2863 165 2867 166
rect 2903 170 2907 171
rect 2903 165 2907 166
rect 2975 170 2979 171
rect 2975 165 2979 166
rect 3095 170 3099 171
rect 3095 165 3099 166
rect 3103 170 3107 171
rect 3103 165 3107 166
rect 3239 170 3243 171
rect 3239 165 3243 166
rect 3287 170 3291 171
rect 3287 165 3291 166
rect 3383 170 3387 171
rect 3383 165 3387 166
rect 3479 170 3483 171
rect 3479 165 3483 166
rect 2656 144 2658 165
rect 2760 144 2762 165
rect 2864 144 2866 165
rect 2976 144 2978 165
rect 3104 144 3106 165
rect 3240 144 3242 165
rect 3384 144 3386 165
rect 2654 143 2660 144
rect 2654 139 2655 143
rect 2659 139 2660 143
rect 2654 138 2660 139
rect 2758 143 2764 144
rect 2758 139 2759 143
rect 2763 139 2764 143
rect 2758 138 2764 139
rect 2862 143 2868 144
rect 2862 139 2863 143
rect 2867 139 2868 143
rect 2862 138 2868 139
rect 2974 143 2980 144
rect 2974 139 2975 143
rect 2979 139 2980 143
rect 2974 138 2980 139
rect 3102 143 3108 144
rect 3102 139 3103 143
rect 3107 139 3108 143
rect 3102 138 3108 139
rect 3238 143 3244 144
rect 3238 139 3239 143
rect 3243 139 3244 143
rect 3238 138 3244 139
rect 3382 143 3388 144
rect 3382 139 3383 143
rect 3387 139 3388 143
rect 3382 138 3388 139
rect 3500 136 3502 250
rect 3556 232 3558 258
rect 3620 232 3622 266
rect 3554 231 3560 232
rect 3554 227 3555 231
rect 3559 227 3560 231
rect 3554 226 3560 227
rect 3618 231 3624 232
rect 3618 227 3619 231
rect 3623 227 3624 231
rect 3618 226 3624 227
rect 3535 170 3539 171
rect 3535 165 3539 166
rect 3536 144 3538 165
rect 3534 143 3540 144
rect 3534 139 3535 143
rect 3539 139 3540 143
rect 3534 138 3540 139
rect 3498 135 3504 136
rect 2730 131 2736 132
rect 2730 127 2731 131
rect 2735 127 2736 131
rect 2730 126 2736 127
rect 2834 131 2840 132
rect 2834 127 2835 131
rect 2839 127 2840 131
rect 2834 126 2840 127
rect 2938 131 2944 132
rect 2938 127 2939 131
rect 2943 127 2944 131
rect 2938 126 2944 127
rect 3050 131 3056 132
rect 3050 127 3051 131
rect 3055 127 3056 131
rect 3050 126 3056 127
rect 3178 131 3184 132
rect 3178 127 3179 131
rect 3183 127 3184 131
rect 3178 126 3184 127
rect 3314 131 3320 132
rect 3314 127 3315 131
rect 3319 127 3320 131
rect 3314 126 3320 127
rect 3458 131 3464 132
rect 3458 127 3459 131
rect 3463 127 3464 131
rect 3498 131 3499 135
rect 3503 131 3504 135
rect 3498 130 3504 131
rect 3458 126 3464 127
rect 2654 124 2660 125
rect 2654 120 2655 124
rect 2659 120 2660 124
rect 2654 119 2660 120
rect 2614 103 2620 104
rect 2614 99 2615 103
rect 2619 99 2620 103
rect 2614 98 2620 99
rect 2656 95 2658 119
rect 2732 104 2734 126
rect 2758 124 2764 125
rect 2758 120 2759 124
rect 2763 120 2764 124
rect 2758 119 2764 120
rect 2730 103 2736 104
rect 2730 99 2731 103
rect 2735 99 2736 103
rect 2730 98 2736 99
rect 2760 95 2762 119
rect 2836 104 2838 126
rect 2862 124 2868 125
rect 2862 120 2863 124
rect 2867 120 2868 124
rect 2862 119 2868 120
rect 2834 103 2840 104
rect 2834 99 2835 103
rect 2839 99 2840 103
rect 2834 98 2840 99
rect 2864 95 2866 119
rect 2940 104 2942 126
rect 2974 124 2980 125
rect 2974 120 2975 124
rect 2979 120 2980 124
rect 2974 119 2980 120
rect 2938 103 2944 104
rect 2938 99 2939 103
rect 2943 99 2944 103
rect 2938 98 2944 99
rect 2976 95 2978 119
rect 3052 104 3054 126
rect 3102 124 3108 125
rect 3102 120 3103 124
rect 3107 120 3108 124
rect 3102 119 3108 120
rect 3050 103 3056 104
rect 3050 99 3051 103
rect 3055 99 3056 103
rect 3050 98 3056 99
rect 3104 95 3106 119
rect 3180 104 3182 126
rect 3238 124 3244 125
rect 3238 120 3239 124
rect 3243 120 3244 124
rect 3238 119 3244 120
rect 3178 103 3184 104
rect 3178 99 3179 103
rect 3183 99 3184 103
rect 3178 98 3184 99
rect 3240 95 3242 119
rect 3316 104 3318 126
rect 3382 124 3388 125
rect 3382 120 3383 124
rect 3387 120 3388 124
rect 3382 119 3388 120
rect 3314 103 3320 104
rect 3314 99 3315 103
rect 3319 99 3320 103
rect 3314 98 3320 99
rect 3384 95 3386 119
rect 3460 104 3462 126
rect 3534 124 3540 125
rect 3534 120 3535 124
rect 3539 120 3540 124
rect 3534 119 3540 120
rect 3458 103 3464 104
rect 3458 99 3459 103
rect 3463 99 3464 103
rect 3458 98 3464 99
rect 3536 95 3538 119
rect 3644 104 3646 302
rect 3710 300 3716 301
rect 3710 296 3711 300
rect 3715 296 3716 300
rect 3710 295 3716 296
rect 3712 271 3714 295
rect 3768 280 3770 462
rect 3942 459 3948 460
rect 3806 456 3812 457
rect 3806 452 3807 456
rect 3811 452 3812 456
rect 3942 455 3943 459
rect 3947 455 3948 459
rect 3942 454 3948 455
rect 3806 451 3812 452
rect 3808 427 3810 451
rect 3906 431 3912 432
rect 3906 427 3907 431
rect 3911 427 3912 431
rect 3944 427 3946 454
rect 3807 426 3811 427
rect 3807 421 3811 422
rect 3839 426 3843 427
rect 3906 426 3912 427
rect 3943 426 3947 427
rect 3839 421 3843 422
rect 3786 419 3792 420
rect 3786 415 3787 419
rect 3791 415 3792 419
rect 3786 414 3792 415
rect 3788 312 3790 414
rect 3840 397 3842 421
rect 3838 396 3844 397
rect 3838 392 3839 396
rect 3843 392 3844 396
rect 3838 391 3844 392
rect 3908 388 3910 426
rect 3943 421 3947 422
rect 3914 419 3920 420
rect 3914 415 3915 419
rect 3919 415 3920 419
rect 3914 414 3920 415
rect 3906 387 3912 388
rect 3906 383 3907 387
rect 3911 383 3912 387
rect 3906 382 3912 383
rect 3838 377 3844 378
rect 3838 373 3839 377
rect 3843 373 3844 377
rect 3838 372 3844 373
rect 3840 347 3842 372
rect 3839 346 3843 347
rect 3839 341 3843 342
rect 3840 320 3842 341
rect 3838 319 3844 320
rect 3838 315 3839 319
rect 3843 315 3844 319
rect 3838 314 3844 315
rect 3916 312 3918 414
rect 3944 394 3946 421
rect 3942 393 3948 394
rect 3942 389 3943 393
rect 3947 389 3948 393
rect 3942 388 3948 389
rect 3942 376 3948 377
rect 3942 372 3943 376
rect 3947 372 3948 376
rect 3942 371 3948 372
rect 3944 347 3946 371
rect 3943 346 3947 347
rect 3943 341 3947 342
rect 3944 321 3946 341
rect 3942 320 3948 321
rect 3942 316 3943 320
rect 3947 316 3948 320
rect 3942 315 3948 316
rect 3786 311 3792 312
rect 3786 307 3787 311
rect 3791 307 3792 311
rect 3786 306 3792 307
rect 3914 311 3920 312
rect 3914 307 3915 311
rect 3919 307 3920 311
rect 3914 306 3920 307
rect 3942 303 3948 304
rect 3838 300 3844 301
rect 3838 296 3839 300
rect 3843 296 3844 300
rect 3942 299 3943 303
rect 3947 299 3948 303
rect 3942 298 3948 299
rect 3838 295 3844 296
rect 3766 279 3772 280
rect 3766 275 3767 279
rect 3771 275 3772 279
rect 3766 274 3772 275
rect 3840 271 3842 295
rect 3906 275 3912 276
rect 3906 271 3907 275
rect 3911 271 3912 275
rect 3944 271 3946 298
rect 3671 270 3675 271
rect 3671 265 3675 266
rect 3711 270 3715 271
rect 3711 265 3715 266
rect 3839 270 3843 271
rect 3906 270 3912 271
rect 3943 270 3947 271
rect 3839 265 3843 266
rect 3672 241 3674 265
rect 3840 241 3842 265
rect 3670 240 3676 241
rect 3670 236 3671 240
rect 3675 236 3676 240
rect 3670 235 3676 236
rect 3838 240 3844 241
rect 3838 236 3839 240
rect 3843 236 3844 240
rect 3838 235 3844 236
rect 3908 232 3910 270
rect 3943 265 3947 266
rect 3914 263 3920 264
rect 3914 259 3915 263
rect 3919 259 3920 263
rect 3914 258 3920 259
rect 3906 231 3912 232
rect 3906 227 3907 231
rect 3911 227 3912 231
rect 3906 226 3912 227
rect 3670 221 3676 222
rect 3670 217 3671 221
rect 3675 217 3676 221
rect 3670 216 3676 217
rect 3838 221 3844 222
rect 3838 217 3839 221
rect 3843 217 3844 221
rect 3838 216 3844 217
rect 3672 171 3674 216
rect 3840 171 3842 216
rect 3671 170 3675 171
rect 3671 165 3675 166
rect 3695 170 3699 171
rect 3695 165 3699 166
rect 3839 170 3843 171
rect 3839 165 3843 166
rect 3696 144 3698 165
rect 3840 144 3842 165
rect 3694 143 3700 144
rect 3694 139 3695 143
rect 3699 139 3700 143
rect 3694 138 3700 139
rect 3838 143 3844 144
rect 3838 139 3839 143
rect 3843 139 3844 143
rect 3838 138 3844 139
rect 3916 136 3918 258
rect 3944 238 3946 265
rect 3942 237 3948 238
rect 3942 233 3943 237
rect 3947 233 3948 237
rect 3942 232 3948 233
rect 3942 220 3948 221
rect 3942 216 3943 220
rect 3947 216 3948 220
rect 3942 215 3948 216
rect 3944 171 3946 215
rect 3943 170 3947 171
rect 3943 165 3947 166
rect 3944 145 3946 165
rect 3942 144 3948 145
rect 3942 140 3943 144
rect 3947 140 3948 144
rect 3942 139 3948 140
rect 3914 135 3920 136
rect 3770 131 3776 132
rect 3770 127 3771 131
rect 3775 127 3776 131
rect 3914 131 3915 135
rect 3919 131 3920 135
rect 3914 130 3920 131
rect 3770 126 3776 127
rect 3942 127 3948 128
rect 3694 124 3700 125
rect 3694 120 3695 124
rect 3699 120 3700 124
rect 3694 119 3700 120
rect 3642 103 3648 104
rect 3642 99 3643 103
rect 3647 99 3648 103
rect 3642 98 3648 99
rect 3696 95 3698 119
rect 3772 104 3774 126
rect 3838 124 3844 125
rect 3838 120 3839 124
rect 3843 120 3844 124
rect 3942 123 3943 127
rect 3947 123 3948 127
rect 3942 122 3948 123
rect 3838 119 3844 120
rect 3770 103 3776 104
rect 3770 99 3771 103
rect 3775 99 3776 103
rect 3770 98 3776 99
rect 3840 95 3842 119
rect 3944 95 3946 122
rect 2047 94 2051 95
rect 111 90 115 91
rect 111 85 115 86
rect 135 90 139 91
rect 135 85 139 86
rect 231 90 235 91
rect 231 85 235 86
rect 327 90 331 91
rect 327 85 331 86
rect 423 90 427 91
rect 423 85 427 86
rect 527 90 531 91
rect 527 85 531 86
rect 647 90 651 91
rect 647 85 651 86
rect 775 90 779 91
rect 775 85 779 86
rect 903 90 907 91
rect 903 85 907 86
rect 1031 90 1035 91
rect 1031 85 1035 86
rect 1151 90 1155 91
rect 1151 85 1155 86
rect 1271 90 1275 91
rect 1271 85 1275 86
rect 1383 90 1387 91
rect 1383 85 1387 86
rect 1487 90 1491 91
rect 1487 85 1491 86
rect 1591 90 1595 91
rect 1591 85 1595 86
rect 1703 90 1707 91
rect 1703 85 1707 86
rect 1807 90 1811 91
rect 1807 85 1811 86
rect 1903 90 1907 91
rect 1903 85 1907 86
rect 2007 90 2011 91
rect 2047 89 2051 90
rect 2071 94 2075 95
rect 2071 89 2075 90
rect 2167 94 2171 95
rect 2167 89 2171 90
rect 2263 94 2267 95
rect 2263 89 2267 90
rect 2359 94 2363 95
rect 2359 89 2363 90
rect 2455 94 2459 95
rect 2455 89 2459 90
rect 2551 94 2555 95
rect 2551 89 2555 90
rect 2655 94 2659 95
rect 2655 89 2659 90
rect 2759 94 2763 95
rect 2759 89 2763 90
rect 2863 94 2867 95
rect 2863 89 2867 90
rect 2975 94 2979 95
rect 2975 89 2979 90
rect 3103 94 3107 95
rect 3103 89 3107 90
rect 3239 94 3243 95
rect 3239 89 3243 90
rect 3383 94 3387 95
rect 3383 89 3387 90
rect 3535 94 3539 95
rect 3535 89 3539 90
rect 3695 94 3699 95
rect 3695 89 3699 90
rect 3839 94 3843 95
rect 3839 89 3843 90
rect 3943 94 3947 95
rect 3943 89 3947 90
rect 2007 85 2011 86
<< m4c >>
rect 111 4026 115 4030
rect 1519 4026 1523 4030
rect 1615 4026 1619 4030
rect 1711 4026 1715 4030
rect 1807 4026 1811 4030
rect 1903 4026 1907 4030
rect 2007 4026 2011 4030
rect 2047 4014 2051 4018
rect 2071 4014 2075 4018
rect 2167 4014 2171 4018
rect 2263 4014 2267 4018
rect 3943 4014 3947 4018
rect 111 3950 115 3954
rect 199 3950 203 3954
rect 295 3950 299 3954
rect 391 3950 395 3954
rect 495 3950 499 3954
rect 615 3950 619 3954
rect 743 3950 747 3954
rect 871 3950 875 3954
rect 999 3950 1003 3954
rect 1127 3950 1131 3954
rect 1255 3950 1259 3954
rect 1383 3950 1387 3954
rect 1511 3950 1515 3954
rect 1519 3950 1523 3954
rect 1615 3950 1619 3954
rect 1647 3950 1651 3954
rect 1711 3950 1715 3954
rect 1807 3950 1811 3954
rect 1903 3950 1907 3954
rect 2007 3950 2011 3954
rect 111 3874 115 3878
rect 199 3874 203 3878
rect 295 3874 299 3878
rect 335 3874 339 3878
rect 391 3874 395 3878
rect 455 3874 459 3878
rect 495 3874 499 3878
rect 583 3874 587 3878
rect 615 3874 619 3878
rect 719 3874 723 3878
rect 743 3874 747 3878
rect 847 3874 851 3878
rect 871 3874 875 3878
rect 975 3874 979 3878
rect 999 3874 1003 3878
rect 1103 3874 1107 3878
rect 1127 3874 1131 3878
rect 2047 3938 2051 3942
rect 2071 3938 2075 3942
rect 2159 3938 2163 3942
rect 2167 3938 2171 3942
rect 2263 3938 2267 3942
rect 2287 3938 2291 3942
rect 2415 3938 2419 3942
rect 2551 3938 2555 3942
rect 2687 3938 2691 3942
rect 2823 3938 2827 3942
rect 2951 3938 2955 3942
rect 3071 3938 3075 3942
rect 3191 3938 3195 3942
rect 3303 3938 3307 3942
rect 3407 3938 3411 3942
rect 3519 3938 3523 3942
rect 3631 3938 3635 3942
rect 3743 3938 3747 3942
rect 3943 3938 3947 3942
rect 1231 3874 1235 3878
rect 1255 3874 1259 3878
rect 1359 3874 1363 3878
rect 1383 3874 1387 3878
rect 1487 3874 1491 3878
rect 1511 3874 1515 3878
rect 1647 3874 1651 3878
rect 2007 3874 2011 3878
rect 2047 3854 2051 3858
rect 2159 3854 2163 3858
rect 2207 3854 2211 3858
rect 2287 3854 2291 3858
rect 2343 3854 2347 3858
rect 2415 3854 2419 3858
rect 2487 3854 2491 3858
rect 2551 3854 2555 3858
rect 2647 3854 2651 3858
rect 2687 3854 2691 3858
rect 111 3794 115 3798
rect 335 3794 339 3798
rect 455 3794 459 3798
rect 503 3794 507 3798
rect 583 3794 587 3798
rect 615 3794 619 3798
rect 719 3794 723 3798
rect 735 3794 739 3798
rect 847 3794 851 3798
rect 863 3794 867 3798
rect 975 3794 979 3798
rect 999 3794 1003 3798
rect 111 3710 115 3714
rect 495 3710 499 3714
rect 503 3710 507 3714
rect 591 3710 595 3714
rect 615 3710 619 3714
rect 687 3710 691 3714
rect 735 3710 739 3714
rect 791 3710 795 3714
rect 863 3710 867 3714
rect 1103 3794 1107 3798
rect 1143 3794 1147 3798
rect 1231 3794 1235 3798
rect 1287 3794 1291 3798
rect 1359 3794 1363 3798
rect 1431 3794 1435 3798
rect 1487 3794 1491 3798
rect 2823 3854 2827 3858
rect 2951 3854 2955 3858
rect 3015 3854 3019 3858
rect 3071 3854 3075 3858
rect 3191 3854 3195 3858
rect 3223 3854 3227 3858
rect 3303 3854 3307 3858
rect 3407 3854 3411 3858
rect 3439 3854 3443 3858
rect 3519 3854 3523 3858
rect 3631 3854 3635 3858
rect 3655 3854 3659 3858
rect 1583 3794 1587 3798
rect 2007 3794 2011 3798
rect 911 3710 915 3714
rect 999 3710 1003 3714
rect 1039 3710 1043 3714
rect 1143 3710 1147 3714
rect 1183 3710 1187 3714
rect 111 3626 115 3630
rect 335 3626 339 3630
rect 463 3626 467 3630
rect 495 3626 499 3630
rect 591 3626 595 3630
rect 607 3626 611 3630
rect 687 3626 691 3630
rect 759 3626 763 3630
rect 791 3626 795 3630
rect 111 3538 115 3542
rect 159 3538 163 3542
rect 303 3538 307 3542
rect 335 3538 339 3542
rect 463 3538 467 3542
rect 607 3538 611 3542
rect 639 3538 643 3542
rect 911 3626 915 3630
rect 927 3626 931 3630
rect 1039 3626 1043 3630
rect 1095 3626 1099 3630
rect 1287 3710 1291 3714
rect 1335 3710 1339 3714
rect 1431 3710 1435 3714
rect 1495 3710 1499 3714
rect 2047 3778 2051 3782
rect 2191 3778 2195 3782
rect 2207 3778 2211 3782
rect 1583 3710 1587 3714
rect 1655 3710 1659 3714
rect 2007 3710 2011 3714
rect 2343 3778 2347 3782
rect 2375 3778 2379 3782
rect 2487 3778 2491 3782
rect 2559 3778 2563 3782
rect 2647 3778 2651 3782
rect 2743 3778 2747 3782
rect 2823 3778 2827 3782
rect 2935 3778 2939 3782
rect 3015 3778 3019 3782
rect 3127 3778 3131 3782
rect 3223 3778 3227 3782
rect 3319 3778 3323 3782
rect 3743 3854 3747 3858
rect 3943 3854 3947 3858
rect 3439 3778 3443 3782
rect 3511 3778 3515 3782
rect 3655 3778 3659 3782
rect 3711 3778 3715 3782
rect 2047 3698 2051 3702
rect 2127 3698 2131 3702
rect 2191 3698 2195 3702
rect 2351 3698 2355 3702
rect 2375 3698 2379 3702
rect 2559 3698 2563 3702
rect 2583 3698 2587 3702
rect 2743 3698 2747 3702
rect 2815 3698 2819 3702
rect 1183 3626 1187 3630
rect 1263 3626 1267 3630
rect 1335 3626 1339 3630
rect 1439 3626 1443 3630
rect 1495 3626 1499 3630
rect 1615 3626 1619 3630
rect 1655 3626 1659 3630
rect 2935 3698 2939 3702
rect 3047 3698 3051 3702
rect 3127 3698 3131 3702
rect 3279 3698 3283 3702
rect 3319 3698 3323 3702
rect 3511 3698 3515 3702
rect 1791 3626 1795 3630
rect 2007 3626 2011 3630
rect 759 3538 763 3542
rect 815 3538 819 3542
rect 927 3538 931 3542
rect 999 3538 1003 3542
rect 1095 3538 1099 3542
rect 1175 3538 1179 3542
rect 1263 3538 1267 3542
rect 111 3454 115 3458
rect 135 3454 139 3458
rect 159 3454 163 3458
rect 303 3454 307 3458
rect 319 3454 323 3458
rect 463 3454 467 3458
rect 535 3454 539 3458
rect 639 3454 643 3458
rect 255 3424 259 3428
rect 751 3454 755 3458
rect 815 3454 819 3458
rect 959 3454 963 3458
rect 999 3454 1003 3458
rect 1351 3538 1355 3542
rect 1439 3538 1443 3542
rect 1527 3538 1531 3542
rect 1615 3538 1619 3542
rect 1703 3538 1707 3542
rect 1791 3538 1795 3542
rect 2047 3614 2051 3618
rect 2127 3614 2131 3618
rect 2191 3614 2195 3618
rect 2327 3614 2331 3618
rect 2351 3614 2355 3618
rect 2455 3614 2459 3618
rect 2583 3614 2587 3618
rect 2719 3614 2723 3618
rect 2815 3614 2819 3618
rect 2855 3614 2859 3618
rect 2999 3614 3003 3618
rect 3047 3614 3051 3618
rect 3143 3614 3147 3618
rect 3279 3614 3283 3618
rect 3295 3614 3299 3618
rect 3943 3778 3947 3782
rect 3711 3698 3715 3702
rect 3751 3698 3755 3702
rect 3943 3698 3947 3702
rect 3455 3614 3459 3618
rect 3511 3614 3515 3618
rect 3623 3614 3627 3618
rect 3751 3614 3755 3618
rect 1879 3538 1883 3542
rect 2007 3538 2011 3542
rect 2047 3538 2051 3542
rect 2103 3538 2107 3542
rect 2191 3538 2195 3542
rect 2271 3538 2275 3542
rect 2327 3538 2331 3542
rect 2447 3538 2451 3542
rect 2455 3538 2459 3542
rect 2583 3538 2587 3542
rect 2631 3538 2635 3542
rect 2719 3538 2723 3542
rect 2815 3538 2819 3542
rect 2855 3538 2859 3542
rect 2999 3538 3003 3542
rect 3143 3538 3147 3542
rect 3175 3538 3179 3542
rect 3295 3538 3299 3542
rect 3351 3538 3355 3542
rect 3455 3538 3459 3542
rect 3519 3538 3523 3542
rect 1159 3454 1163 3458
rect 1175 3454 1179 3458
rect 1351 3454 1355 3458
rect 1527 3454 1531 3458
rect 1535 3454 1539 3458
rect 799 3424 803 3428
rect 111 3378 115 3382
rect 135 3378 139 3382
rect 231 3378 235 3382
rect 319 3378 323 3382
rect 375 3378 379 3382
rect 535 3378 539 3382
rect 703 3378 707 3382
rect 751 3378 755 3382
rect 1703 3454 1707 3458
rect 1719 3454 1723 3458
rect 1879 3454 1883 3458
rect 1903 3454 1907 3458
rect 2007 3454 2011 3458
rect 2047 3458 2051 3462
rect 2103 3458 2107 3462
rect 2127 3458 2131 3462
rect 871 3378 875 3382
rect 959 3378 963 3382
rect 1047 3378 1051 3382
rect 1159 3378 1163 3382
rect 1215 3378 1219 3382
rect 1351 3378 1355 3382
rect 1383 3378 1387 3382
rect 111 3302 115 3306
rect 135 3302 139 3306
rect 231 3302 235 3306
rect 279 3302 283 3306
rect 375 3302 379 3306
rect 463 3302 467 3306
rect 535 3302 539 3306
rect 663 3302 667 3306
rect 703 3302 707 3306
rect 871 3302 875 3306
rect 1047 3302 1051 3306
rect 1079 3302 1083 3306
rect 111 3226 115 3230
rect 135 3226 139 3230
rect 279 3226 283 3230
rect 287 3226 291 3230
rect 447 3226 451 3230
rect 463 3226 467 3230
rect 1535 3378 1539 3382
rect 1543 3378 1547 3382
rect 1703 3378 1707 3382
rect 1719 3378 1723 3382
rect 1871 3378 1875 3382
rect 1903 3378 1907 3382
rect 2007 3378 2011 3382
rect 2271 3458 2275 3462
rect 2311 3458 2315 3462
rect 2447 3458 2451 3462
rect 2495 3458 2499 3462
rect 2631 3458 2635 3462
rect 2679 3458 2683 3462
rect 2815 3458 2819 3462
rect 2863 3458 2867 3462
rect 2999 3458 3003 3462
rect 3047 3458 3051 3462
rect 3175 3458 3179 3462
rect 3223 3458 3227 3462
rect 2047 3366 2051 3370
rect 2071 3366 2075 3370
rect 2127 3366 2131 3370
rect 2215 3366 2219 3370
rect 2311 3366 2315 3370
rect 2359 3366 2363 3370
rect 2495 3366 2499 3370
rect 2511 3366 2515 3370
rect 2655 3366 2659 3370
rect 2679 3366 2683 3370
rect 2799 3366 2803 3370
rect 2863 3366 2867 3370
rect 2935 3366 2939 3370
rect 1215 3302 1219 3306
rect 1295 3302 1299 3306
rect 1383 3302 1387 3306
rect 1519 3302 1523 3306
rect 1543 3302 1547 3306
rect 1703 3302 1707 3306
rect 1743 3302 1747 3306
rect 1871 3302 1875 3306
rect 2007 3302 2011 3306
rect 615 3226 619 3230
rect 663 3226 667 3230
rect 791 3226 795 3230
rect 871 3226 875 3230
rect 967 3226 971 3230
rect 1079 3226 1083 3230
rect 1143 3226 1147 3230
rect 1295 3226 1299 3230
rect 1327 3226 1331 3230
rect 111 3146 115 3150
rect 135 3146 139 3150
rect 287 3146 291 3150
rect 311 3146 315 3150
rect 439 3146 443 3150
rect 447 3146 451 3150
rect 583 3146 587 3150
rect 615 3146 619 3150
rect 743 3146 747 3150
rect 791 3146 795 3150
rect 903 3146 907 3150
rect 967 3146 971 3150
rect 111 3062 115 3066
rect 311 3062 315 3066
rect 1511 3226 1515 3230
rect 1519 3226 1523 3230
rect 1695 3226 1699 3230
rect 1743 3226 1747 3230
rect 2047 3282 2051 3286
rect 2071 3282 2075 3286
rect 2111 3282 2115 3286
rect 2007 3226 2011 3230
rect 2215 3282 2219 3286
rect 2247 3282 2251 3286
rect 2359 3282 2363 3286
rect 2399 3282 2403 3286
rect 2511 3282 2515 3286
rect 2575 3282 2579 3286
rect 2655 3282 2659 3286
rect 2783 3282 2787 3286
rect 2799 3282 2803 3286
rect 3351 3458 3355 3462
rect 3623 3538 3627 3542
rect 3687 3538 3691 3542
rect 3407 3458 3411 3462
rect 3519 3458 3523 3462
rect 3591 3458 3595 3462
rect 3687 3458 3691 3462
rect 3775 3458 3779 3462
rect 3047 3366 3051 3370
rect 3079 3366 3083 3370
rect 3223 3366 3227 3370
rect 3375 3366 3379 3370
rect 3407 3366 3411 3370
rect 3535 3366 3539 3370
rect 3591 3366 3595 3370
rect 3299 3304 3303 3308
rect 2935 3282 2939 3286
rect 3015 3282 3019 3286
rect 3079 3282 3083 3286
rect 3223 3282 3227 3286
rect 3263 3282 3267 3286
rect 3375 3282 3379 3286
rect 3943 3614 3947 3618
rect 3839 3538 3843 3542
rect 3943 3538 3947 3542
rect 3839 3458 3843 3462
rect 3695 3366 3699 3370
rect 3775 3366 3779 3370
rect 3839 3366 3843 3370
rect 3507 3304 3511 3308
rect 2047 3206 2051 3210
rect 2071 3206 2075 3210
rect 2111 3206 2115 3210
rect 2167 3206 2171 3210
rect 1063 3146 1067 3150
rect 1143 3146 1147 3150
rect 1223 3146 1227 3150
rect 1327 3146 1331 3150
rect 1391 3146 1395 3150
rect 2247 3206 2251 3210
rect 2263 3206 2267 3210
rect 2359 3206 2363 3210
rect 2399 3206 2403 3210
rect 2455 3206 2459 3210
rect 2551 3206 2555 3210
rect 2575 3206 2579 3210
rect 2647 3206 2651 3210
rect 2743 3206 2747 3210
rect 2783 3206 2787 3210
rect 2839 3206 2843 3210
rect 2935 3206 2939 3210
rect 3015 3206 3019 3210
rect 3031 3206 3035 3210
rect 3127 3206 3131 3210
rect 3223 3206 3227 3210
rect 3263 3206 3267 3210
rect 3319 3206 3323 3210
rect 3527 3282 3531 3286
rect 3535 3282 3539 3286
rect 3695 3282 3699 3286
rect 3791 3282 3795 3286
rect 3839 3282 3843 3286
rect 3439 3206 3443 3210
rect 3527 3206 3531 3210
rect 3575 3206 3579 3210
rect 3719 3206 3723 3210
rect 3791 3206 3795 3210
rect 3839 3206 3843 3210
rect 1511 3146 1515 3150
rect 1559 3146 1563 3150
rect 1695 3146 1699 3150
rect 1727 3146 1731 3150
rect 2007 3146 2011 3150
rect 439 3062 443 3066
rect 503 3062 507 3066
rect 583 3062 587 3066
rect 599 3062 603 3066
rect 703 3062 707 3066
rect 743 3062 747 3066
rect 815 3062 819 3066
rect 903 3062 907 3066
rect 935 3062 939 3066
rect 1063 3062 1067 3066
rect 1071 3062 1075 3066
rect 1223 3062 1227 3066
rect 111 2982 115 2986
rect 503 2982 507 2986
rect 551 2982 555 2986
rect 599 2982 603 2986
rect 647 2982 651 2986
rect 703 2982 707 2986
rect 759 2982 763 2986
rect 815 2982 819 2986
rect 887 2982 891 2986
rect 935 2982 939 2986
rect 111 2898 115 2902
rect 471 2898 475 2902
rect 551 2898 555 2902
rect 575 2898 579 2902
rect 647 2898 651 2902
rect 695 2898 699 2902
rect 759 2898 763 2902
rect 839 2898 843 2902
rect 887 2898 891 2902
rect 1023 2982 1027 2986
rect 1071 2982 1075 2986
rect 1383 3062 1387 3066
rect 1391 3062 1395 3066
rect 1551 3062 1555 3066
rect 1559 3062 1563 3066
rect 1719 3062 1723 3066
rect 1727 3062 1731 3066
rect 2047 3118 2051 3122
rect 2071 3118 2075 3122
rect 2167 3118 2171 3122
rect 2263 3118 2267 3122
rect 2007 3062 2011 3066
rect 2047 3042 2051 3046
rect 2071 3042 2075 3046
rect 1175 2982 1179 2986
rect 1223 2982 1227 2986
rect 1327 2982 1331 2986
rect 1383 2982 1387 2986
rect 1487 2982 1491 2986
rect 1551 2982 1555 2986
rect 2335 3118 2339 3122
rect 2359 3118 2363 3122
rect 2455 3118 2459 3122
rect 2551 3118 2555 3122
rect 2623 3118 2627 3122
rect 2647 3118 2651 3122
rect 2743 3118 2747 3122
rect 2839 3118 2843 3122
rect 2911 3118 2915 3122
rect 2935 3118 2939 3122
rect 3031 3118 3035 3122
rect 3127 3118 3131 3122
rect 3207 3118 3211 3122
rect 3223 3118 3227 3122
rect 3319 3118 3323 3122
rect 3439 3118 3443 3122
rect 3503 3118 3507 3122
rect 3575 3118 3579 3122
rect 3719 3118 3723 3122
rect 3799 3118 3803 3122
rect 3839 3118 3843 3122
rect 3943 3458 3947 3462
rect 3943 3366 3947 3370
rect 3943 3282 3947 3286
rect 3943 3206 3947 3210
rect 2335 3042 2339 3046
rect 2383 3042 2387 3046
rect 2623 3042 2627 3046
rect 2703 3042 2707 3046
rect 2911 3042 2915 3046
rect 2999 3042 3003 3046
rect 3207 3042 3211 3046
rect 3287 3042 3291 3046
rect 3503 3042 3507 3046
rect 3575 3042 3579 3046
rect 3799 3042 3803 3046
rect 3839 3042 3843 3046
rect 1655 2982 1659 2986
rect 1719 2982 1723 2986
rect 1823 2982 1827 2986
rect 2007 2982 2011 2986
rect 991 2898 995 2902
rect 1023 2898 1027 2902
rect 1151 2898 1155 2902
rect 1175 2898 1179 2902
rect 1319 2898 1323 2902
rect 1327 2898 1331 2902
rect 1487 2898 1491 2902
rect 1495 2898 1499 2902
rect 1655 2898 1659 2902
rect 1671 2898 1675 2902
rect 1823 2898 1827 2902
rect 1847 2898 1851 2902
rect 2047 2962 2051 2966
rect 2071 2962 2075 2966
rect 2383 2962 2387 2966
rect 2391 2962 2395 2966
rect 2007 2898 2011 2902
rect 2047 2886 2051 2890
rect 2071 2886 2075 2890
rect 111 2818 115 2822
rect 471 2818 475 2822
rect 479 2818 483 2822
rect 575 2818 579 2822
rect 679 2818 683 2822
rect 695 2818 699 2822
rect 799 2818 803 2822
rect 839 2818 843 2822
rect 935 2818 939 2822
rect 991 2818 995 2822
rect 1079 2818 1083 2822
rect 1151 2818 1155 2822
rect 1239 2818 1243 2822
rect 1319 2818 1323 2822
rect 111 2738 115 2742
rect 479 2738 483 2742
rect 511 2738 515 2742
rect 575 2738 579 2742
rect 623 2738 627 2742
rect 679 2738 683 2742
rect 743 2738 747 2742
rect 799 2738 803 2742
rect 879 2738 883 2742
rect 935 2738 939 2742
rect 1415 2818 1419 2822
rect 1495 2818 1499 2822
rect 2703 2962 2707 2966
rect 2975 2962 2979 2966
rect 2999 2962 3003 2966
rect 3215 2962 3219 2966
rect 3287 2962 3291 2966
rect 3439 2962 3443 2966
rect 3575 2962 3579 2966
rect 3647 2962 3651 2966
rect 3839 2962 3843 2966
rect 2295 2886 2299 2890
rect 2391 2886 2395 2890
rect 2535 2886 2539 2890
rect 2703 2886 2707 2890
rect 2767 2886 2771 2890
rect 2975 2886 2979 2890
rect 2991 2886 2995 2890
rect 3215 2886 3219 2890
rect 3431 2886 3435 2890
rect 3439 2886 3443 2890
rect 1599 2818 1603 2822
rect 1671 2818 1675 2822
rect 1783 2818 1787 2822
rect 1847 2818 1851 2822
rect 2007 2818 2011 2822
rect 1015 2738 1019 2742
rect 1079 2738 1083 2742
rect 1159 2738 1163 2742
rect 1239 2738 1243 2742
rect 1311 2738 1315 2742
rect 1415 2738 1419 2742
rect 1463 2738 1467 2742
rect 1599 2738 1603 2742
rect 1623 2738 1627 2742
rect 1783 2738 1787 2742
rect 2047 2806 2051 2810
rect 2071 2806 2075 2810
rect 2199 2806 2203 2810
rect 2295 2806 2299 2810
rect 2367 2806 2371 2810
rect 2535 2806 2539 2810
rect 2551 2806 2555 2810
rect 2007 2738 2011 2742
rect 2735 2806 2739 2810
rect 2767 2806 2771 2810
rect 2927 2806 2931 2810
rect 2991 2806 2995 2810
rect 3111 2806 3115 2810
rect 3215 2806 3219 2810
rect 3295 2806 3299 2810
rect 3431 2806 3435 2810
rect 3647 2886 3651 2890
rect 3839 2886 3843 2890
rect 3479 2806 3483 2810
rect 3647 2806 3651 2810
rect 3671 2806 3675 2810
rect 3839 2806 3843 2810
rect 2047 2726 2051 2730
rect 2071 2726 2075 2730
rect 2191 2726 2195 2730
rect 2199 2726 2203 2730
rect 2319 2726 2323 2730
rect 2367 2726 2371 2730
rect 2447 2726 2451 2730
rect 2551 2726 2555 2730
rect 2583 2726 2587 2730
rect 2727 2726 2731 2730
rect 2735 2726 2739 2730
rect 2887 2726 2891 2730
rect 2927 2726 2931 2730
rect 3063 2726 3067 2730
rect 3111 2726 3115 2730
rect 3255 2726 3259 2730
rect 3295 2726 3299 2730
rect 111 2658 115 2662
rect 367 2658 371 2662
rect 487 2658 491 2662
rect 511 2658 515 2662
rect 615 2658 619 2662
rect 623 2658 627 2662
rect 743 2658 747 2662
rect 751 2658 755 2662
rect 111 2582 115 2586
rect 135 2582 139 2586
rect 287 2582 291 2586
rect 367 2582 371 2586
rect 447 2582 451 2586
rect 487 2582 491 2586
rect 607 2582 611 2586
rect 615 2582 619 2586
rect 879 2658 883 2662
rect 895 2658 899 2662
rect 1015 2658 1019 2662
rect 1031 2658 1035 2662
rect 1159 2658 1163 2662
rect 1167 2658 1171 2662
rect 1303 2658 1307 2662
rect 1311 2658 1315 2662
rect 1431 2658 1435 2662
rect 1463 2658 1467 2662
rect 1567 2658 1571 2662
rect 1623 2658 1627 2662
rect 1703 2658 1707 2662
rect 1783 2658 1787 2662
rect 2007 2658 2011 2662
rect 751 2582 755 2586
rect 767 2582 771 2586
rect 895 2582 899 2586
rect 919 2582 923 2586
rect 111 2490 115 2494
rect 135 2490 139 2494
rect 231 2490 235 2494
rect 287 2490 291 2494
rect 327 2490 331 2494
rect 423 2490 427 2494
rect 447 2490 451 2494
rect 111 2398 115 2402
rect 135 2398 139 2402
rect 1031 2582 1035 2586
rect 1063 2582 1067 2586
rect 1167 2582 1171 2586
rect 1199 2582 1203 2586
rect 1303 2582 1307 2586
rect 1335 2582 1339 2586
rect 1431 2582 1435 2586
rect 1463 2582 1467 2586
rect 1567 2582 1571 2586
rect 1591 2582 1595 2586
rect 1703 2582 1707 2586
rect 1727 2582 1731 2586
rect 2047 2642 2051 2646
rect 2071 2642 2075 2646
rect 2191 2642 2195 2646
rect 2231 2642 2235 2646
rect 2319 2642 2323 2646
rect 2335 2642 2339 2646
rect 2447 2642 2451 2646
rect 2007 2582 2011 2586
rect 2559 2642 2563 2646
rect 2583 2642 2587 2646
rect 2671 2642 2675 2646
rect 2727 2642 2731 2646
rect 3455 2726 3459 2730
rect 3479 2726 3483 2730
rect 3655 2726 3659 2730
rect 3671 2726 3675 2730
rect 3943 3118 3947 3122
rect 3943 3042 3947 3046
rect 3943 2962 3947 2966
rect 3943 2886 3947 2890
rect 3943 2806 3947 2810
rect 3839 2726 3843 2730
rect 3943 2726 3947 2730
rect 2791 2642 2795 2646
rect 2887 2642 2891 2646
rect 2911 2642 2915 2646
rect 3031 2642 3035 2646
rect 3063 2642 3067 2646
rect 3151 2642 3155 2646
rect 3255 2642 3259 2646
rect 3455 2642 3459 2646
rect 3655 2642 3659 2646
rect 3839 2642 3843 2646
rect 3943 2642 3947 2646
rect 2047 2562 2051 2566
rect 2231 2562 2235 2566
rect 2335 2562 2339 2566
rect 2383 2562 2387 2566
rect 2447 2562 2451 2566
rect 2495 2562 2499 2566
rect 2559 2562 2563 2566
rect 2615 2562 2619 2566
rect 2671 2562 2675 2566
rect 2743 2562 2747 2566
rect 2791 2562 2795 2566
rect 2871 2562 2875 2566
rect 2911 2562 2915 2566
rect 2991 2562 2995 2566
rect 3031 2562 3035 2566
rect 3111 2562 3115 2566
rect 3151 2562 3155 2566
rect 3231 2562 3235 2566
rect 3359 2562 3363 2566
rect 3487 2562 3491 2566
rect 3943 2562 3947 2566
rect 519 2490 523 2494
rect 607 2490 611 2494
rect 767 2490 771 2494
rect 919 2490 923 2494
rect 1063 2490 1067 2494
rect 1199 2490 1203 2494
rect 1335 2490 1339 2494
rect 1463 2490 1467 2494
rect 1591 2490 1595 2494
rect 1727 2490 1731 2494
rect 2007 2490 2011 2494
rect 2047 2482 2051 2486
rect 2383 2482 2387 2486
rect 2495 2482 2499 2486
rect 2535 2482 2539 2486
rect 2615 2482 2619 2486
rect 2711 2482 2715 2486
rect 2743 2482 2747 2486
rect 231 2398 235 2402
rect 255 2398 259 2402
rect 327 2398 331 2402
rect 415 2398 419 2402
rect 423 2398 427 2402
rect 519 2398 523 2402
rect 575 2398 579 2402
rect 735 2398 739 2402
rect 887 2398 891 2402
rect 1039 2398 1043 2402
rect 1183 2398 1187 2402
rect 1327 2398 1331 2402
rect 1479 2398 1483 2402
rect 2007 2398 2011 2402
rect 2871 2482 2875 2486
rect 2879 2482 2883 2486
rect 2991 2482 2995 2486
rect 3047 2482 3051 2486
rect 3111 2482 3115 2486
rect 3207 2482 3211 2486
rect 3231 2482 3235 2486
rect 3359 2482 3363 2486
rect 3487 2482 3491 2486
rect 3503 2482 3507 2486
rect 3655 2482 3659 2486
rect 3807 2482 3811 2486
rect 3943 2482 3947 2486
rect 2047 2394 2051 2398
rect 2535 2394 2539 2398
rect 2607 2394 2611 2398
rect 2711 2394 2715 2398
rect 2815 2394 2819 2398
rect 2879 2394 2883 2398
rect 3007 2394 3011 2398
rect 3047 2394 3051 2398
rect 111 2322 115 2326
rect 135 2322 139 2326
rect 255 2322 259 2326
rect 263 2322 267 2326
rect 415 2322 419 2326
rect 423 2322 427 2326
rect 575 2322 579 2326
rect 583 2322 587 2326
rect 735 2322 739 2326
rect 743 2322 747 2326
rect 111 2242 115 2246
rect 135 2242 139 2246
rect 887 2322 891 2326
rect 895 2322 899 2326
rect 3191 2394 3195 2398
rect 3207 2394 3211 2398
rect 3359 2394 3363 2398
rect 3503 2394 3507 2398
rect 3519 2394 3523 2398
rect 3655 2394 3659 2398
rect 3679 2394 3683 2398
rect 3807 2394 3811 2398
rect 3839 2394 3843 2398
rect 1039 2322 1043 2326
rect 1047 2322 1051 2326
rect 1183 2322 1187 2326
rect 1199 2322 1203 2326
rect 1327 2322 1331 2326
rect 1351 2322 1355 2326
rect 1479 2322 1483 2326
rect 1503 2322 1507 2326
rect 223 2242 227 2246
rect 263 2242 267 2246
rect 351 2242 355 2246
rect 423 2242 427 2246
rect 495 2242 499 2246
rect 583 2242 587 2246
rect 647 2242 651 2246
rect 743 2242 747 2246
rect 799 2242 803 2246
rect 895 2242 899 2246
rect 959 2242 963 2246
rect 1047 2242 1051 2246
rect 1119 2242 1123 2246
rect 1199 2242 1203 2246
rect 2007 2322 2011 2326
rect 2047 2302 2051 2306
rect 2071 2302 2075 2306
rect 2167 2302 2171 2306
rect 2271 2302 2275 2306
rect 2415 2302 2419 2306
rect 2575 2302 2579 2306
rect 2607 2302 2611 2306
rect 2743 2302 2747 2306
rect 2815 2302 2819 2306
rect 1279 2242 1283 2246
rect 1351 2242 1355 2246
rect 1439 2242 1443 2246
rect 1503 2242 1507 2246
rect 1599 2242 1603 2246
rect 2007 2242 2011 2246
rect 2047 2226 2051 2230
rect 2071 2226 2075 2230
rect 2167 2226 2171 2230
rect 2175 2226 2179 2230
rect 111 2166 115 2170
rect 223 2166 227 2170
rect 351 2166 355 2170
rect 471 2166 475 2170
rect 495 2166 499 2170
rect 567 2166 571 2170
rect 647 2166 651 2170
rect 679 2166 683 2170
rect 799 2166 803 2170
rect 807 2166 811 2170
rect 943 2166 947 2170
rect 959 2166 963 2170
rect 1079 2166 1083 2170
rect 1119 2166 1123 2170
rect 2271 2226 2275 2230
rect 2319 2226 2323 2230
rect 2415 2226 2419 2230
rect 2471 2226 2475 2230
rect 2575 2226 2579 2230
rect 2623 2226 2627 2230
rect 1223 2166 1227 2170
rect 1279 2166 1283 2170
rect 1367 2166 1371 2170
rect 1439 2166 1443 2170
rect 1503 2166 1507 2170
rect 1599 2166 1603 2170
rect 1639 2166 1643 2170
rect 1783 2166 1787 2170
rect 1903 2166 1907 2170
rect 2007 2166 2011 2170
rect 111 2090 115 2094
rect 471 2090 475 2094
rect 567 2090 571 2094
rect 623 2090 627 2094
rect 679 2090 683 2094
rect 735 2090 739 2094
rect 807 2090 811 2094
rect 855 2090 859 2094
rect 943 2090 947 2094
rect 983 2090 987 2094
rect 1079 2090 1083 2094
rect 1119 2090 1123 2094
rect 1223 2090 1227 2094
rect 1255 2090 1259 2094
rect 1367 2090 1371 2094
rect 1391 2090 1395 2094
rect 1503 2090 1507 2094
rect 1527 2090 1531 2094
rect 1639 2090 1643 2094
rect 1655 2090 1659 2094
rect 2047 2130 2051 2134
rect 2071 2130 2075 2134
rect 2175 2130 2179 2134
rect 2279 2130 2283 2134
rect 2319 2130 2323 2134
rect 1783 2090 1787 2094
rect 1791 2090 1795 2094
rect 111 2010 115 2014
rect 447 2010 451 2014
rect 575 2010 579 2014
rect 623 2010 627 2014
rect 727 2010 731 2014
rect 735 2010 739 2014
rect 111 1934 115 1938
rect 447 1934 451 1938
rect 111 1858 115 1862
rect 319 1858 323 1862
rect 447 1858 451 1862
rect 111 1778 115 1782
rect 255 1778 259 1782
rect 319 1778 323 1782
rect 855 2010 859 2014
rect 887 2010 891 2014
rect 983 2010 987 2014
rect 1055 2010 1059 2014
rect 1119 2010 1123 2014
rect 1231 2010 1235 2014
rect 1255 2010 1259 2014
rect 575 1934 579 1938
rect 655 1934 659 1938
rect 727 1934 731 1938
rect 751 1934 755 1938
rect 847 1934 851 1938
rect 887 1934 891 1938
rect 943 1934 947 1938
rect 1039 1934 1043 1938
rect 1055 1934 1059 1938
rect 1391 2010 1395 2014
rect 1399 2010 1403 2014
rect 2743 2226 2747 2230
rect 2783 2226 2787 2230
rect 2911 2302 2915 2306
rect 3007 2302 3011 2306
rect 3071 2302 3075 2306
rect 3191 2302 3195 2306
rect 3231 2302 3235 2306
rect 3359 2302 3363 2306
rect 3383 2302 3387 2306
rect 3519 2302 3523 2306
rect 3535 2302 3539 2306
rect 3943 2394 3947 2398
rect 3679 2302 3683 2306
rect 3695 2302 3699 2306
rect 3839 2302 3843 2306
rect 3943 2302 3947 2306
rect 2911 2226 2915 2230
rect 2935 2226 2939 2230
rect 3071 2226 3075 2230
rect 3079 2226 3083 2230
rect 3223 2226 3227 2230
rect 3231 2226 3235 2230
rect 3367 2226 3371 2230
rect 3383 2226 3387 2230
rect 2391 2130 2395 2134
rect 2471 2130 2475 2134
rect 2511 2130 2515 2134
rect 2623 2130 2627 2134
rect 2631 2130 2635 2134
rect 2759 2130 2763 2134
rect 2783 2130 2787 2134
rect 1903 2090 1907 2094
rect 2007 2090 2011 2094
rect 1527 2010 1531 2014
rect 1575 2010 1579 2014
rect 1655 2010 1659 2014
rect 1751 2010 1755 2014
rect 1791 2010 1795 2014
rect 1903 2010 1907 2014
rect 2047 2046 2051 2050
rect 2279 2046 2283 2050
rect 2327 2046 2331 2050
rect 2391 2046 2395 2050
rect 2431 2046 2435 2050
rect 2511 2046 2515 2050
rect 2007 2010 2011 2014
rect 2535 2046 2539 2050
rect 2631 2046 2635 2050
rect 2647 2046 2651 2050
rect 1135 1934 1139 1938
rect 2047 1966 2051 1970
rect 2255 1966 2259 1970
rect 2327 1966 2331 1970
rect 2351 1966 2355 1970
rect 2431 1966 2435 1970
rect 2447 1966 2451 1970
rect 2535 1966 2539 1970
rect 2543 1966 2547 1970
rect 1231 1934 1235 1938
rect 1327 1934 1331 1938
rect 1399 1934 1403 1938
rect 1423 1934 1427 1938
rect 1575 1934 1579 1938
rect 1751 1934 1755 1938
rect 1903 1934 1907 1938
rect 2007 1934 2011 1938
rect 2895 2130 2899 2134
rect 2935 2130 2939 2134
rect 3519 2226 3523 2230
rect 3535 2226 3539 2230
rect 3695 2226 3699 2230
rect 3943 2226 3947 2230
rect 3039 2130 3043 2134
rect 3079 2130 3083 2134
rect 3191 2130 3195 2134
rect 3223 2130 3227 2134
rect 3351 2130 3355 2134
rect 3367 2130 3371 2134
rect 3519 2130 3523 2134
rect 3687 2130 3691 2134
rect 3839 2130 3843 2134
rect 3943 2130 3947 2134
rect 2759 2046 2763 2050
rect 2775 2046 2779 2050
rect 2895 2046 2899 2050
rect 2919 2046 2923 2050
rect 3039 2046 3043 2050
rect 3079 2046 3083 2050
rect 3191 2046 3195 2050
rect 3263 2046 3267 2050
rect 3351 2046 3355 2050
rect 2647 1966 2651 1970
rect 583 1858 587 1862
rect 655 1858 659 1862
rect 719 1858 723 1862
rect 751 1858 755 1862
rect 847 1858 851 1862
rect 855 1858 859 1862
rect 943 1858 947 1862
rect 991 1858 995 1862
rect 1039 1858 1043 1862
rect 1127 1858 1131 1862
rect 1135 1858 1139 1862
rect 1231 1858 1235 1862
rect 1263 1858 1267 1862
rect 1327 1858 1331 1862
rect 391 1778 395 1782
rect 447 1778 451 1782
rect 535 1778 539 1782
rect 583 1778 587 1782
rect 695 1778 699 1782
rect 719 1778 723 1782
rect 855 1778 859 1782
rect 863 1778 867 1782
rect 111 1702 115 1706
rect 135 1702 139 1706
rect 255 1702 259 1706
rect 263 1702 267 1706
rect 391 1702 395 1706
rect 431 1702 435 1706
rect 111 1626 115 1630
rect 135 1626 139 1630
rect 535 1702 539 1706
rect 607 1702 611 1706
rect 991 1778 995 1782
rect 1031 1778 1035 1782
rect 1127 1778 1131 1782
rect 1399 1858 1403 1862
rect 1423 1858 1427 1862
rect 2047 1878 2051 1882
rect 2183 1878 2187 1882
rect 2255 1878 2259 1882
rect 2279 1878 2283 1882
rect 2351 1878 2355 1882
rect 2383 1878 2387 1882
rect 2447 1878 2451 1882
rect 1535 1858 1539 1862
rect 2007 1858 2011 1862
rect 1207 1778 1211 1782
rect 1263 1778 1267 1782
rect 1383 1778 1387 1782
rect 1399 1778 1403 1782
rect 2047 1798 2051 1802
rect 2127 1798 2131 1802
rect 2183 1798 2187 1802
rect 1535 1778 1539 1782
rect 1559 1778 1563 1782
rect 1743 1778 1747 1782
rect 2007 1778 2011 1782
rect 2487 1878 2491 1882
rect 2543 1878 2547 1882
rect 2591 1878 2595 1882
rect 2767 1966 2771 1970
rect 2775 1966 2779 1970
rect 3455 2046 3459 2050
rect 3519 2046 3523 2050
rect 3655 2046 3659 2050
rect 3687 2046 3691 2050
rect 2919 1966 2923 1970
rect 3079 1966 3083 1970
rect 3103 1966 3107 1970
rect 3263 1966 3267 1970
rect 3319 1966 3323 1970
rect 3455 1966 3459 1970
rect 3543 1966 3547 1970
rect 3655 1966 3659 1970
rect 3775 1966 3779 1970
rect 2647 1878 2651 1882
rect 2703 1878 2707 1882
rect 2767 1878 2771 1882
rect 2831 1878 2835 1882
rect 2919 1878 2923 1882
rect 2991 1878 2995 1882
rect 3103 1878 3107 1882
rect 3183 1878 3187 1882
rect 3319 1878 3323 1882
rect 3399 1878 3403 1882
rect 3543 1878 3547 1882
rect 3631 1878 3635 1882
rect 2279 1798 2283 1802
rect 2311 1798 2315 1802
rect 2383 1798 2387 1802
rect 2487 1798 2491 1802
rect 2495 1798 2499 1802
rect 2591 1798 2595 1802
rect 2687 1798 2691 1802
rect 2703 1798 2707 1802
rect 695 1702 699 1706
rect 799 1702 803 1706
rect 863 1702 867 1706
rect 999 1702 1003 1706
rect 1031 1702 1035 1706
rect 1199 1702 1203 1706
rect 1207 1702 1211 1706
rect 1383 1702 1387 1706
rect 1407 1702 1411 1706
rect 1559 1702 1563 1706
rect 1623 1702 1627 1706
rect 1743 1702 1747 1706
rect 263 1626 267 1630
rect 287 1626 291 1630
rect 431 1626 435 1630
rect 471 1626 475 1630
rect 607 1626 611 1630
rect 655 1626 659 1630
rect 799 1626 803 1630
rect 839 1626 843 1630
rect 111 1546 115 1550
rect 135 1546 139 1550
rect 287 1546 291 1550
rect 295 1546 299 1550
rect 111 1470 115 1474
rect 135 1470 139 1474
rect 175 1470 179 1474
rect 471 1546 475 1550
rect 487 1546 491 1550
rect 655 1546 659 1550
rect 687 1546 691 1550
rect 999 1626 1003 1630
rect 1015 1626 1019 1630
rect 1183 1626 1187 1630
rect 1199 1626 1203 1630
rect 2047 1718 2051 1722
rect 2071 1718 2075 1722
rect 2127 1718 2131 1722
rect 2191 1718 2195 1722
rect 2311 1718 2315 1722
rect 2343 1718 2347 1722
rect 2495 1718 2499 1722
rect 2511 1718 2515 1722
rect 1839 1702 1843 1706
rect 2007 1702 2011 1706
rect 1343 1626 1347 1630
rect 1407 1626 1411 1630
rect 1495 1626 1499 1630
rect 839 1546 843 1550
rect 887 1546 891 1550
rect 1015 1546 1019 1550
rect 1079 1546 1083 1550
rect 1183 1546 1187 1550
rect 1263 1546 1267 1550
rect 1343 1546 1347 1550
rect 2047 1642 2051 1646
rect 2071 1642 2075 1646
rect 2191 1642 2195 1646
rect 1623 1626 1627 1630
rect 1639 1626 1643 1630
rect 1783 1626 1787 1630
rect 1839 1626 1843 1630
rect 1903 1626 1907 1630
rect 2007 1626 2011 1630
rect 2831 1798 2835 1802
rect 2879 1798 2883 1802
rect 2991 1798 2995 1802
rect 3071 1798 3075 1802
rect 3183 1798 3187 1802
rect 3263 1798 3267 1802
rect 3399 1798 3403 1802
rect 3463 1798 3467 1802
rect 3631 1798 3635 1802
rect 3663 1798 3667 1802
rect 2687 1718 2691 1722
rect 2871 1718 2875 1722
rect 2879 1718 2883 1722
rect 3063 1718 3067 1722
rect 3071 1718 3075 1722
rect 3255 1718 3259 1722
rect 3263 1718 3267 1722
rect 3447 1718 3451 1722
rect 3463 1718 3467 1722
rect 2335 1642 2339 1646
rect 2343 1642 2347 1646
rect 2511 1642 2515 1646
rect 2599 1642 2603 1646
rect 2687 1642 2691 1646
rect 2839 1642 2843 1646
rect 2871 1642 2875 1646
rect 3047 1642 3051 1646
rect 3063 1642 3067 1646
rect 3647 1718 3651 1722
rect 3663 1718 3667 1722
rect 3839 2046 3843 2050
rect 3943 2046 3947 2050
rect 3839 1966 3843 1970
rect 3775 1878 3779 1882
rect 3839 1878 3843 1882
rect 3839 1798 3843 1802
rect 3943 1966 3947 1970
rect 3943 1878 3947 1882
rect 3943 1798 3947 1802
rect 3839 1718 3843 1722
rect 3943 1718 3947 1722
rect 3231 1642 3235 1646
rect 3255 1642 3259 1646
rect 3399 1642 3403 1646
rect 3447 1642 3451 1646
rect 3551 1642 3555 1646
rect 2047 1562 2051 1566
rect 2071 1562 2075 1566
rect 2335 1562 2339 1566
rect 2583 1562 2587 1566
rect 2599 1562 2603 1566
rect 1447 1546 1451 1550
rect 1495 1546 1499 1550
rect 1623 1546 1627 1550
rect 1639 1546 1643 1550
rect 1783 1546 1787 1550
rect 1807 1546 1811 1550
rect 1903 1546 1907 1550
rect 2007 1546 2011 1550
rect 295 1470 299 1474
rect 359 1470 363 1474
rect 487 1470 491 1474
rect 567 1470 571 1474
rect 687 1470 691 1474
rect 783 1470 787 1474
rect 111 1394 115 1398
rect 175 1394 179 1398
rect 327 1394 331 1398
rect 359 1394 363 1398
rect 887 1470 891 1474
rect 1007 1470 1011 1474
rect 1079 1470 1083 1474
rect 1231 1470 1235 1474
rect 1263 1470 1267 1474
rect 1447 1470 1451 1474
rect 1463 1470 1467 1474
rect 1623 1470 1627 1474
rect 1695 1470 1699 1474
rect 1807 1470 1811 1474
rect 2743 1562 2747 1566
rect 2839 1562 2843 1566
rect 2903 1562 2907 1566
rect 3047 1562 3051 1566
rect 3063 1562 3067 1566
rect 3223 1562 3227 1566
rect 3231 1562 3235 1566
rect 3383 1562 3387 1566
rect 3399 1562 3403 1566
rect 3647 1642 3651 1646
rect 3695 1642 3699 1646
rect 3839 1642 3843 1646
rect 3943 1642 3947 1646
rect 3543 1562 3547 1566
rect 3551 1562 3555 1566
rect 3695 1562 3699 1566
rect 3703 1562 3707 1566
rect 3839 1562 3843 1566
rect 2047 1486 2051 1490
rect 2415 1486 2419 1490
rect 2511 1486 2515 1490
rect 2583 1486 2587 1490
rect 2607 1486 2611 1490
rect 2703 1486 2707 1490
rect 2743 1486 2747 1490
rect 2799 1486 2803 1490
rect 2903 1486 2907 1490
rect 2919 1486 2923 1490
rect 1903 1470 1907 1474
rect 2007 1470 2011 1474
rect 463 1394 467 1398
rect 567 1394 571 1398
rect 599 1394 603 1398
rect 727 1394 731 1398
rect 783 1394 787 1398
rect 855 1394 859 1398
rect 519 1387 523 1388
rect 519 1384 523 1387
rect 983 1394 987 1398
rect 1007 1394 1011 1398
rect 1119 1394 1123 1398
rect 1231 1394 1235 1398
rect 1263 1394 1267 1398
rect 1423 1394 1427 1398
rect 1463 1394 1467 1398
rect 1583 1394 1587 1398
rect 1695 1394 1699 1398
rect 963 1384 967 1388
rect 111 1310 115 1314
rect 327 1310 331 1314
rect 463 1310 467 1314
rect 551 1310 555 1314
rect 599 1310 603 1314
rect 655 1310 659 1314
rect 727 1310 731 1314
rect 767 1310 771 1314
rect 855 1310 859 1314
rect 879 1310 883 1314
rect 983 1310 987 1314
rect 991 1310 995 1314
rect 1103 1310 1107 1314
rect 1119 1310 1123 1314
rect 111 1234 115 1238
rect 391 1234 395 1238
rect 519 1234 523 1238
rect 551 1234 555 1238
rect 655 1234 659 1238
rect 663 1234 667 1238
rect 767 1234 771 1238
rect 807 1234 811 1238
rect 879 1234 883 1238
rect 959 1234 963 1238
rect 111 1154 115 1158
rect 175 1154 179 1158
rect 327 1154 331 1158
rect 391 1154 395 1158
rect 495 1154 499 1158
rect 519 1154 523 1158
rect 663 1154 667 1158
rect 671 1154 675 1158
rect 991 1234 995 1238
rect 807 1154 811 1158
rect 847 1154 851 1158
rect 959 1154 963 1158
rect 1031 1154 1035 1158
rect 111 1070 115 1074
rect 135 1070 139 1074
rect 175 1070 179 1074
rect 231 1070 235 1074
rect 111 994 115 998
rect 135 994 139 998
rect 1215 1310 1219 1314
rect 1263 1310 1267 1314
rect 1327 1310 1331 1314
rect 1751 1394 1755 1398
rect 1903 1394 1907 1398
rect 2007 1394 2011 1398
rect 2047 1390 2051 1394
rect 2071 1390 2075 1394
rect 2303 1390 2307 1394
rect 2415 1390 2419 1394
rect 2511 1390 2515 1394
rect 2559 1390 2563 1394
rect 2607 1390 2611 1394
rect 1423 1310 1427 1314
rect 1439 1310 1443 1314
rect 1559 1310 1563 1314
rect 1583 1310 1587 1314
rect 1103 1234 1107 1238
rect 1111 1234 1115 1238
rect 1215 1234 1219 1238
rect 1255 1234 1259 1238
rect 1327 1234 1331 1238
rect 1407 1234 1411 1238
rect 1439 1234 1443 1238
rect 1111 1154 1115 1158
rect 1207 1154 1211 1158
rect 1255 1154 1259 1158
rect 1751 1310 1755 1314
rect 1903 1310 1907 1314
rect 2007 1310 2011 1314
rect 2047 1306 2051 1310
rect 2071 1306 2075 1310
rect 2223 1306 2227 1310
rect 2303 1306 2307 1310
rect 3063 1486 3067 1490
rect 3223 1486 3227 1490
rect 3231 1486 3235 1490
rect 3383 1486 3387 1490
rect 3415 1486 3419 1490
rect 3543 1486 3547 1490
rect 3615 1486 3619 1490
rect 3703 1486 3707 1490
rect 3815 1486 3819 1490
rect 3943 1562 3947 1566
rect 3943 1486 3947 1490
rect 2703 1390 2707 1394
rect 2799 1390 2803 1394
rect 2807 1390 2811 1394
rect 2919 1390 2923 1394
rect 3055 1390 3059 1394
rect 3063 1390 3067 1394
rect 3231 1390 3235 1394
rect 3303 1390 3307 1394
rect 3415 1390 3419 1394
rect 3559 1390 3563 1394
rect 3615 1390 3619 1394
rect 3815 1390 3819 1394
rect 3943 1390 3947 1394
rect 2415 1306 2419 1310
rect 2559 1306 2563 1310
rect 2615 1306 2619 1310
rect 2807 1306 2811 1310
rect 2815 1306 2819 1310
rect 2999 1306 3003 1310
rect 3055 1306 3059 1310
rect 3175 1306 3179 1310
rect 3303 1306 3307 1310
rect 3343 1306 3347 1310
rect 3503 1306 3507 1310
rect 3559 1306 3563 1310
rect 3663 1306 3667 1310
rect 3815 1306 3819 1310
rect 3831 1306 3835 1310
rect 1559 1234 1563 1238
rect 1711 1234 1715 1238
rect 2007 1234 2011 1238
rect 2047 1222 2051 1226
rect 2071 1222 2075 1226
rect 2135 1222 2139 1226
rect 2223 1222 2227 1226
rect 2311 1222 2315 1226
rect 2415 1222 2419 1226
rect 2503 1222 2507 1226
rect 1383 1154 1387 1158
rect 1407 1154 1411 1158
rect 1559 1154 1563 1158
rect 1567 1154 1571 1158
rect 327 1070 331 1074
rect 375 1070 379 1074
rect 495 1070 499 1074
rect 543 1070 547 1074
rect 671 1070 675 1074
rect 727 1070 731 1074
rect 847 1070 851 1074
rect 911 1070 915 1074
rect 1031 1070 1035 1074
rect 1095 1070 1099 1074
rect 243 1056 247 1060
rect 859 1056 863 1060
rect 3943 1306 3947 1310
rect 2615 1222 2619 1226
rect 2695 1222 2699 1226
rect 2815 1222 2819 1226
rect 2887 1222 2891 1226
rect 2999 1222 3003 1226
rect 3071 1222 3075 1226
rect 3175 1222 3179 1226
rect 3239 1222 3243 1226
rect 3343 1222 3347 1226
rect 3399 1222 3403 1226
rect 3503 1222 3507 1226
rect 3551 1222 3555 1226
rect 3663 1222 3667 1226
rect 3703 1222 3707 1226
rect 1711 1154 1715 1158
rect 1751 1154 1755 1158
rect 2007 1154 2011 1158
rect 2047 1138 2051 1142
rect 2135 1138 2139 1142
rect 2295 1138 2299 1142
rect 2311 1138 2315 1142
rect 2423 1138 2427 1142
rect 2503 1138 2507 1142
rect 2559 1138 2563 1142
rect 2695 1138 2699 1142
rect 2839 1138 2843 1142
rect 2887 1138 2891 1142
rect 1207 1070 1211 1074
rect 1279 1070 1283 1074
rect 1383 1070 1387 1074
rect 1463 1070 1467 1074
rect 1567 1070 1571 1074
rect 1647 1070 1651 1074
rect 1751 1070 1755 1074
rect 1831 1070 1835 1074
rect 231 994 235 998
rect 271 994 275 998
rect 375 994 379 998
rect 447 994 451 998
rect 543 994 547 998
rect 631 994 635 998
rect 727 994 731 998
rect 823 994 827 998
rect 911 994 915 998
rect 1007 994 1011 998
rect 1095 994 1099 998
rect 1175 994 1179 998
rect 1279 994 1283 998
rect 3831 1222 3835 1226
rect 3839 1222 3843 1226
rect 3943 1222 3947 1226
rect 2991 1138 2995 1142
rect 3071 1138 3075 1142
rect 3151 1138 3155 1142
rect 3239 1138 3243 1142
rect 3319 1138 3323 1142
rect 3399 1138 3403 1142
rect 2007 1070 2011 1074
rect 2047 1058 2051 1062
rect 2295 1058 2299 1062
rect 2423 1058 2427 1062
rect 2495 1058 2499 1062
rect 2559 1058 2563 1062
rect 2599 1058 2603 1062
rect 2695 1058 2699 1062
rect 2711 1058 2715 1062
rect 2839 1058 2843 1062
rect 2847 1058 2851 1062
rect 2991 1058 2995 1062
rect 3007 1058 3011 1062
rect 3151 1058 3155 1062
rect 3199 1058 3203 1062
rect 1335 994 1339 998
rect 1463 994 1467 998
rect 1487 994 1491 998
rect 111 918 115 922
rect 135 918 139 922
rect 271 918 275 922
rect 447 918 451 922
rect 455 918 459 922
rect 631 918 635 922
rect 655 918 659 922
rect 823 918 827 922
rect 855 918 859 922
rect 111 842 115 846
rect 135 842 139 846
rect 1007 918 1011 922
rect 1055 918 1059 922
rect 1631 994 1635 998
rect 1647 994 1651 998
rect 1775 994 1779 998
rect 1831 994 1835 998
rect 1903 994 1907 998
rect 2007 994 2011 998
rect 2047 982 2051 986
rect 2495 982 2499 986
rect 2599 982 2603 986
rect 2647 982 2651 986
rect 2711 982 2715 986
rect 2743 982 2747 986
rect 2847 982 2851 986
rect 3495 1138 3499 1142
rect 3551 1138 3555 1142
rect 3679 1138 3683 1142
rect 3703 1138 3707 1142
rect 3839 1138 3843 1142
rect 3943 1138 3947 1142
rect 3319 1058 3323 1062
rect 3407 1058 3411 1062
rect 3495 1058 3499 1062
rect 3631 1058 3635 1062
rect 3679 1058 3683 1062
rect 3839 1058 3843 1062
rect 3191 1024 3195 1028
rect 3559 1024 3563 1028
rect 3943 1058 3947 1062
rect 2967 982 2971 986
rect 3007 982 3011 986
rect 1175 918 1179 922
rect 1239 918 1243 922
rect 1335 918 1339 922
rect 1415 918 1419 922
rect 1487 918 1491 922
rect 1583 918 1587 922
rect 1631 918 1635 922
rect 1751 918 1755 922
rect 1775 918 1779 922
rect 1903 918 1907 922
rect 2007 918 2011 922
rect 215 842 219 846
rect 271 842 275 846
rect 343 842 347 846
rect 455 842 459 846
rect 495 842 499 846
rect 655 842 659 846
rect 831 842 835 846
rect 855 842 859 846
rect 1007 842 1011 846
rect 1055 842 1059 846
rect 111 766 115 770
rect 215 766 219 770
rect 343 766 347 770
rect 375 766 379 770
rect 495 766 499 770
rect 623 766 627 770
rect 655 766 659 770
rect 751 766 755 770
rect 831 766 835 770
rect 111 690 115 694
rect 375 690 379 694
rect 495 690 499 694
rect 527 690 531 694
rect 623 690 627 694
rect 631 690 635 694
rect 743 690 747 694
rect 751 690 755 694
rect 887 766 891 770
rect 1007 766 1011 770
rect 1023 766 1027 770
rect 1183 842 1187 846
rect 1239 842 1243 846
rect 1359 842 1363 846
rect 1415 842 1419 846
rect 1535 842 1539 846
rect 1583 842 1587 846
rect 2047 894 2051 898
rect 2071 894 2075 898
rect 2255 894 2259 898
rect 2463 894 2467 898
rect 2647 894 2651 898
rect 2679 894 2683 898
rect 2743 894 2747 898
rect 3111 982 3115 986
rect 3199 982 3203 986
rect 3279 982 3283 986
rect 3407 982 3411 986
rect 3463 982 3467 986
rect 3631 982 3635 986
rect 3663 982 3667 986
rect 3839 982 3843 986
rect 3943 982 3947 986
rect 2847 894 2851 898
rect 2895 894 2899 898
rect 2967 894 2971 898
rect 3111 894 3115 898
rect 3127 894 3131 898
rect 3279 894 3283 898
rect 3367 894 3371 898
rect 3463 894 3467 898
rect 3615 894 3619 898
rect 3663 894 3667 898
rect 3839 894 3843 898
rect 1719 842 1723 846
rect 1751 842 1755 846
rect 1903 842 1907 846
rect 2007 842 2011 846
rect 2047 818 2051 822
rect 2071 818 2075 822
rect 2215 818 2219 822
rect 2255 818 2259 822
rect 2327 818 2331 822
rect 1167 766 1171 770
rect 1183 766 1187 770
rect 1311 766 1315 770
rect 1359 766 1363 770
rect 1455 766 1459 770
rect 1535 766 1539 770
rect 1599 766 1603 770
rect 855 690 859 694
rect 887 690 891 694
rect 967 690 971 694
rect 1023 690 1027 694
rect 1071 690 1075 694
rect 1167 690 1171 694
rect 1183 690 1187 694
rect 111 614 115 618
rect 527 614 531 618
rect 631 614 635 618
rect 687 614 691 618
rect 743 614 747 618
rect 783 614 787 618
rect 855 614 859 618
rect 879 614 883 618
rect 967 614 971 618
rect 975 614 979 618
rect 1071 614 1075 618
rect 1295 690 1299 694
rect 1311 690 1315 694
rect 1719 766 1723 770
rect 2007 766 2011 770
rect 2447 818 2451 822
rect 2463 818 2467 822
rect 2583 818 2587 822
rect 2679 818 2683 822
rect 2735 818 2739 822
rect 2895 818 2899 822
rect 3943 894 3947 898
rect 3063 818 3067 822
rect 3127 818 3131 822
rect 3247 818 3251 822
rect 3367 818 3371 822
rect 3447 818 3451 822
rect 3615 818 3619 822
rect 3655 818 3659 822
rect 2047 738 2051 742
rect 2215 738 2219 742
rect 2327 738 2331 742
rect 2375 738 2379 742
rect 2447 738 2451 742
rect 2495 738 2499 742
rect 2583 738 2587 742
rect 2623 738 2627 742
rect 2735 738 2739 742
rect 2767 738 2771 742
rect 2895 738 2899 742
rect 2911 738 2915 742
rect 3063 738 3067 742
rect 1407 690 1411 694
rect 1455 690 1459 694
rect 1519 690 1523 694
rect 1599 690 1603 694
rect 2007 690 2011 694
rect 2047 654 2051 658
rect 2111 654 2115 658
rect 2247 654 2251 658
rect 2375 654 2379 658
rect 2399 654 2403 658
rect 2495 654 2499 658
rect 2575 654 2579 658
rect 1167 614 1171 618
rect 1183 614 1187 618
rect 1263 614 1267 618
rect 1295 614 1299 618
rect 1359 614 1363 618
rect 1407 614 1411 618
rect 1455 614 1459 618
rect 1519 614 1523 618
rect 111 518 115 522
rect 383 518 387 522
rect 479 518 483 522
rect 575 518 579 522
rect 671 518 675 522
rect 687 518 691 522
rect 767 518 771 522
rect 783 518 787 522
rect 863 518 867 522
rect 879 518 883 522
rect 959 518 963 522
rect 975 518 979 522
rect 1055 518 1059 522
rect 1071 518 1075 522
rect 1151 518 1155 522
rect 1167 518 1171 522
rect 1247 518 1251 522
rect 1263 518 1267 522
rect 2007 614 2011 618
rect 2623 654 2627 658
rect 2759 654 2763 658
rect 2767 654 2771 658
rect 2911 654 2915 658
rect 2943 654 2947 658
rect 3063 654 3067 658
rect 3215 738 3219 742
rect 3247 738 3251 742
rect 3839 818 3843 822
rect 3943 818 3947 822
rect 3367 738 3371 742
rect 3447 738 3451 742
rect 3519 738 3523 742
rect 3655 738 3659 742
rect 3679 738 3683 742
rect 3839 738 3843 742
rect 3127 654 3131 658
rect 3215 654 3219 658
rect 3303 654 3307 658
rect 3367 654 3371 658
rect 3479 654 3483 658
rect 3519 654 3523 658
rect 3655 654 3659 658
rect 3679 654 3683 658
rect 2047 574 2051 578
rect 2071 574 2075 578
rect 2111 574 2115 578
rect 2183 574 2187 578
rect 2247 574 2251 578
rect 2335 574 2339 578
rect 2399 574 2403 578
rect 2503 574 2507 578
rect 2575 574 2579 578
rect 2687 574 2691 578
rect 2759 574 2763 578
rect 2879 574 2883 578
rect 2943 574 2947 578
rect 3071 574 3075 578
rect 3127 574 3131 578
rect 3263 574 3267 578
rect 3303 574 3307 578
rect 1343 518 1347 522
rect 1359 518 1363 522
rect 1439 518 1443 522
rect 1455 518 1459 522
rect 1535 518 1539 522
rect 2007 518 2011 522
rect 2047 498 2051 502
rect 2071 498 2075 502
rect 2183 498 2187 502
rect 2319 498 2323 502
rect 2335 498 2339 502
rect 2463 498 2467 502
rect 2503 498 2507 502
rect 2615 498 2619 502
rect 111 430 115 434
rect 383 430 387 434
rect 479 430 483 434
rect 487 430 491 434
rect 575 430 579 434
rect 583 430 587 434
rect 671 430 675 434
rect 687 430 691 434
rect 767 430 771 434
rect 791 430 795 434
rect 863 430 867 434
rect 895 430 899 434
rect 959 430 963 434
rect 539 419 543 420
rect 539 416 543 419
rect 859 416 863 420
rect 111 350 115 354
rect 327 350 331 354
rect 463 350 467 354
rect 487 350 491 354
rect 583 350 587 354
rect 615 350 619 354
rect 687 350 691 354
rect 767 350 771 354
rect 791 350 795 354
rect 999 430 1003 434
rect 1055 430 1059 434
rect 1103 430 1107 434
rect 1151 430 1155 434
rect 1207 430 1211 434
rect 1247 430 1251 434
rect 1319 430 1323 434
rect 1343 430 1347 434
rect 1431 430 1435 434
rect 1439 430 1443 434
rect 895 350 899 354
rect 919 350 923 354
rect 999 350 1003 354
rect 1063 350 1067 354
rect 1103 350 1107 354
rect 1207 350 1211 354
rect 1319 350 1323 354
rect 1351 350 1355 354
rect 1535 430 1539 434
rect 2007 430 2011 434
rect 2687 498 2691 502
rect 2775 498 2779 502
rect 2879 498 2883 502
rect 2959 498 2963 502
rect 3071 498 3075 502
rect 3159 498 3163 502
rect 3831 654 3835 658
rect 3839 654 3843 658
rect 3943 738 3947 742
rect 3943 654 3947 658
rect 3455 574 3459 578
rect 3479 574 3483 578
rect 3647 574 3651 578
rect 3655 574 3659 578
rect 3831 574 3835 578
rect 3839 574 3843 578
rect 3943 574 3947 578
rect 3263 498 3267 502
rect 3367 498 3371 502
rect 3455 498 3459 502
rect 3583 498 3587 502
rect 3647 498 3651 502
rect 3807 498 3811 502
rect 3839 498 3843 502
rect 3943 498 3947 502
rect 2047 422 2051 426
rect 2183 422 2187 426
rect 2319 422 2323 426
rect 2343 422 2347 426
rect 2463 422 2467 426
rect 2487 422 2491 426
rect 2615 422 2619 426
rect 2639 422 2643 426
rect 2775 422 2779 426
rect 2799 422 2803 426
rect 2959 422 2963 426
rect 3111 422 3115 426
rect 3159 422 3163 426
rect 3263 422 3267 426
rect 3367 422 3371 426
rect 3415 422 3419 426
rect 3559 422 3563 426
rect 3583 422 3587 426
rect 3711 422 3715 426
rect 1431 350 1435 354
rect 1495 350 1499 354
rect 1639 350 1643 354
rect 2007 350 2011 354
rect 2047 342 2051 346
rect 2343 342 2347 346
rect 2487 342 2491 346
rect 2495 342 2499 346
rect 2639 342 2643 346
rect 2799 342 2803 346
rect 111 266 115 270
rect 167 266 171 270
rect 327 266 331 270
rect 463 266 467 270
rect 503 266 507 270
rect 615 266 619 270
rect 687 266 691 270
rect 767 266 771 270
rect 871 266 875 270
rect 919 266 923 270
rect 1047 266 1051 270
rect 1063 266 1067 270
rect 1207 266 1211 270
rect 1215 266 1219 270
rect 111 162 115 166
rect 135 162 139 166
rect 167 162 171 166
rect 231 162 235 166
rect 327 162 331 166
rect 423 162 427 166
rect 503 162 507 166
rect 527 162 531 166
rect 647 162 651 166
rect 687 162 691 166
rect 775 162 779 166
rect 1351 266 1355 270
rect 1367 266 1371 270
rect 1495 266 1499 270
rect 1511 266 1515 270
rect 2551 280 2555 284
rect 2959 342 2963 346
rect 3111 342 3115 346
rect 3119 342 3123 346
rect 3263 342 3267 346
rect 3271 342 3275 346
rect 3415 342 3419 346
rect 3423 342 3427 346
rect 3559 342 3563 346
rect 3567 342 3571 346
rect 3711 342 3715 346
rect 2899 280 2903 284
rect 1639 266 1643 270
rect 1647 266 1651 270
rect 1783 266 1787 270
rect 1903 266 1907 270
rect 2007 266 2011 270
rect 2047 266 2051 270
rect 2071 266 2075 270
rect 2271 266 2275 270
rect 2495 266 2499 270
rect 2639 266 2643 270
rect 2703 266 2707 270
rect 2799 266 2803 270
rect 2903 266 2907 270
rect 2959 266 2963 270
rect 871 162 875 166
rect 903 162 907 166
rect 1031 162 1035 166
rect 1047 162 1051 166
rect 1151 162 1155 166
rect 1215 162 1219 166
rect 1271 162 1275 166
rect 1367 162 1371 166
rect 1383 162 1387 166
rect 1487 162 1491 166
rect 1511 162 1515 166
rect 1591 162 1595 166
rect 1647 162 1651 166
rect 1703 162 1707 166
rect 1783 162 1787 166
rect 1807 162 1811 166
rect 1903 162 1907 166
rect 2007 162 2011 166
rect 2047 166 2051 170
rect 2071 166 2075 170
rect 2167 166 2171 170
rect 2263 166 2267 170
rect 2271 166 2275 170
rect 2359 166 2363 170
rect 2455 166 2459 170
rect 2495 166 2499 170
rect 3095 266 3099 270
rect 3119 266 3123 270
rect 3271 266 3275 270
rect 3287 266 3291 270
rect 3423 266 3427 270
rect 3479 266 3483 270
rect 3567 266 3571 270
rect 2551 166 2555 170
rect 2655 166 2659 170
rect 2703 166 2707 170
rect 2759 166 2763 170
rect 2863 166 2867 170
rect 2903 166 2907 170
rect 2975 166 2979 170
rect 3095 166 3099 170
rect 3103 166 3107 170
rect 3239 166 3243 170
rect 3287 166 3291 170
rect 3383 166 3387 170
rect 3479 166 3483 170
rect 3535 166 3539 170
rect 3807 422 3811 426
rect 3839 422 3843 426
rect 3943 422 3947 426
rect 3839 342 3843 346
rect 3943 342 3947 346
rect 3671 266 3675 270
rect 3711 266 3715 270
rect 3839 266 3843 270
rect 3943 266 3947 270
rect 3671 166 3675 170
rect 3695 166 3699 170
rect 3839 166 3843 170
rect 3943 166 3947 170
rect 111 86 115 90
rect 135 86 139 90
rect 231 86 235 90
rect 327 86 331 90
rect 423 86 427 90
rect 527 86 531 90
rect 647 86 651 90
rect 775 86 779 90
rect 903 86 907 90
rect 1031 86 1035 90
rect 1151 86 1155 90
rect 1271 86 1275 90
rect 1383 86 1387 90
rect 1487 86 1491 90
rect 1591 86 1595 90
rect 1703 86 1707 90
rect 1807 86 1811 90
rect 1903 86 1907 90
rect 2007 86 2011 90
rect 2047 90 2051 94
rect 2071 90 2075 94
rect 2167 90 2171 94
rect 2263 90 2267 94
rect 2359 90 2363 94
rect 2455 90 2459 94
rect 2551 90 2555 94
rect 2655 90 2659 94
rect 2759 90 2763 94
rect 2863 90 2867 94
rect 2975 90 2979 94
rect 3103 90 3107 94
rect 3239 90 3243 94
rect 3383 90 3387 94
rect 3535 90 3539 94
rect 3695 90 3699 94
rect 3839 90 3843 94
rect 3943 90 3947 94
<< m4 >>
rect 96 4025 97 4031
rect 103 4030 2031 4031
rect 103 4026 111 4030
rect 115 4026 1519 4030
rect 1523 4026 1615 4030
rect 1619 4026 1711 4030
rect 1715 4026 1807 4030
rect 1811 4026 1903 4030
rect 1907 4026 2007 4030
rect 2011 4026 2031 4030
rect 103 4025 2031 4026
rect 2037 4025 2038 4031
rect 2018 4013 2019 4019
rect 2025 4018 3967 4019
rect 2025 4014 2047 4018
rect 2051 4014 2071 4018
rect 2075 4014 2167 4018
rect 2171 4014 2263 4018
rect 2267 4014 3943 4018
rect 3947 4014 3967 4018
rect 2025 4013 3967 4014
rect 3973 4013 3974 4019
rect 84 3949 85 3955
rect 91 3954 2019 3955
rect 91 3950 111 3954
rect 115 3950 199 3954
rect 203 3950 295 3954
rect 299 3950 391 3954
rect 395 3950 495 3954
rect 499 3950 615 3954
rect 619 3950 743 3954
rect 747 3950 871 3954
rect 875 3950 999 3954
rect 1003 3950 1127 3954
rect 1131 3950 1255 3954
rect 1259 3950 1383 3954
rect 1387 3950 1511 3954
rect 1515 3950 1519 3954
rect 1523 3950 1615 3954
rect 1619 3950 1647 3954
rect 1651 3950 1711 3954
rect 1715 3950 1807 3954
rect 1811 3950 1903 3954
rect 1907 3950 2007 3954
rect 2011 3950 2019 3954
rect 91 3949 2019 3950
rect 2025 3949 2026 3955
rect 2030 3937 2031 3943
rect 2037 3942 3979 3943
rect 2037 3938 2047 3942
rect 2051 3938 2071 3942
rect 2075 3938 2159 3942
rect 2163 3938 2167 3942
rect 2171 3938 2263 3942
rect 2267 3938 2287 3942
rect 2291 3938 2415 3942
rect 2419 3938 2551 3942
rect 2555 3938 2687 3942
rect 2691 3938 2823 3942
rect 2827 3938 2951 3942
rect 2955 3938 3071 3942
rect 3075 3938 3191 3942
rect 3195 3938 3303 3942
rect 3307 3938 3407 3942
rect 3411 3938 3519 3942
rect 3523 3938 3631 3942
rect 3635 3938 3743 3942
rect 3747 3938 3943 3942
rect 3947 3938 3979 3942
rect 2037 3937 3979 3938
rect 3985 3937 3986 3943
rect 96 3873 97 3879
rect 103 3878 2031 3879
rect 103 3874 111 3878
rect 115 3874 199 3878
rect 203 3874 295 3878
rect 299 3874 335 3878
rect 339 3874 391 3878
rect 395 3874 455 3878
rect 459 3874 495 3878
rect 499 3874 583 3878
rect 587 3874 615 3878
rect 619 3874 719 3878
rect 723 3874 743 3878
rect 747 3874 847 3878
rect 851 3874 871 3878
rect 875 3874 975 3878
rect 979 3874 999 3878
rect 1003 3874 1103 3878
rect 1107 3874 1127 3878
rect 1131 3874 1231 3878
rect 1235 3874 1255 3878
rect 1259 3874 1359 3878
rect 1363 3874 1383 3878
rect 1387 3874 1487 3878
rect 1491 3874 1511 3878
rect 1515 3874 1647 3878
rect 1651 3874 2007 3878
rect 2011 3874 2031 3878
rect 103 3873 2031 3874
rect 2037 3873 2038 3879
rect 2018 3853 2019 3859
rect 2025 3858 3967 3859
rect 2025 3854 2047 3858
rect 2051 3854 2159 3858
rect 2163 3854 2207 3858
rect 2211 3854 2287 3858
rect 2291 3854 2343 3858
rect 2347 3854 2415 3858
rect 2419 3854 2487 3858
rect 2491 3854 2551 3858
rect 2555 3854 2647 3858
rect 2651 3854 2687 3858
rect 2691 3854 2823 3858
rect 2827 3854 2951 3858
rect 2955 3854 3015 3858
rect 3019 3854 3071 3858
rect 3075 3854 3191 3858
rect 3195 3854 3223 3858
rect 3227 3854 3303 3858
rect 3307 3854 3407 3858
rect 3411 3854 3439 3858
rect 3443 3854 3519 3858
rect 3523 3854 3631 3858
rect 3635 3854 3655 3858
rect 3659 3854 3743 3858
rect 3747 3854 3943 3858
rect 3947 3854 3967 3858
rect 2025 3853 3967 3854
rect 3973 3853 3974 3859
rect 84 3793 85 3799
rect 91 3798 2019 3799
rect 91 3794 111 3798
rect 115 3794 335 3798
rect 339 3794 455 3798
rect 459 3794 503 3798
rect 507 3794 583 3798
rect 587 3794 615 3798
rect 619 3794 719 3798
rect 723 3794 735 3798
rect 739 3794 847 3798
rect 851 3794 863 3798
rect 867 3794 975 3798
rect 979 3794 999 3798
rect 1003 3794 1103 3798
rect 1107 3794 1143 3798
rect 1147 3794 1231 3798
rect 1235 3794 1287 3798
rect 1291 3794 1359 3798
rect 1363 3794 1431 3798
rect 1435 3794 1487 3798
rect 1491 3794 1583 3798
rect 1587 3794 2007 3798
rect 2011 3794 2019 3798
rect 91 3793 2019 3794
rect 2025 3793 2026 3799
rect 2030 3777 2031 3783
rect 2037 3782 3979 3783
rect 2037 3778 2047 3782
rect 2051 3778 2191 3782
rect 2195 3778 2207 3782
rect 2211 3778 2343 3782
rect 2347 3778 2375 3782
rect 2379 3778 2487 3782
rect 2491 3778 2559 3782
rect 2563 3778 2647 3782
rect 2651 3778 2743 3782
rect 2747 3778 2823 3782
rect 2827 3778 2935 3782
rect 2939 3778 3015 3782
rect 3019 3778 3127 3782
rect 3131 3778 3223 3782
rect 3227 3778 3319 3782
rect 3323 3778 3439 3782
rect 3443 3778 3511 3782
rect 3515 3778 3655 3782
rect 3659 3778 3711 3782
rect 3715 3778 3943 3782
rect 3947 3778 3979 3782
rect 2037 3777 3979 3778
rect 3985 3777 3986 3783
rect 96 3709 97 3715
rect 103 3714 2031 3715
rect 103 3710 111 3714
rect 115 3710 495 3714
rect 499 3710 503 3714
rect 507 3710 591 3714
rect 595 3710 615 3714
rect 619 3710 687 3714
rect 691 3710 735 3714
rect 739 3710 791 3714
rect 795 3710 863 3714
rect 867 3710 911 3714
rect 915 3710 999 3714
rect 1003 3710 1039 3714
rect 1043 3710 1143 3714
rect 1147 3710 1183 3714
rect 1187 3710 1287 3714
rect 1291 3710 1335 3714
rect 1339 3710 1431 3714
rect 1435 3710 1495 3714
rect 1499 3710 1583 3714
rect 1587 3710 1655 3714
rect 1659 3710 2007 3714
rect 2011 3710 2031 3714
rect 103 3709 2031 3710
rect 2037 3709 2038 3715
rect 2018 3697 2019 3703
rect 2025 3702 3967 3703
rect 2025 3698 2047 3702
rect 2051 3698 2127 3702
rect 2131 3698 2191 3702
rect 2195 3698 2351 3702
rect 2355 3698 2375 3702
rect 2379 3698 2559 3702
rect 2563 3698 2583 3702
rect 2587 3698 2743 3702
rect 2747 3698 2815 3702
rect 2819 3698 2935 3702
rect 2939 3698 3047 3702
rect 3051 3698 3127 3702
rect 3131 3698 3279 3702
rect 3283 3698 3319 3702
rect 3323 3698 3511 3702
rect 3515 3698 3711 3702
rect 3715 3698 3751 3702
rect 3755 3698 3943 3702
rect 3947 3698 3967 3702
rect 2025 3697 3967 3698
rect 3973 3697 3974 3703
rect 84 3625 85 3631
rect 91 3630 2019 3631
rect 91 3626 111 3630
rect 115 3626 335 3630
rect 339 3626 463 3630
rect 467 3626 495 3630
rect 499 3626 591 3630
rect 595 3626 607 3630
rect 611 3626 687 3630
rect 691 3626 759 3630
rect 763 3626 791 3630
rect 795 3626 911 3630
rect 915 3626 927 3630
rect 931 3626 1039 3630
rect 1043 3626 1095 3630
rect 1099 3626 1183 3630
rect 1187 3626 1263 3630
rect 1267 3626 1335 3630
rect 1339 3626 1439 3630
rect 1443 3626 1495 3630
rect 1499 3626 1615 3630
rect 1619 3626 1655 3630
rect 1659 3626 1791 3630
rect 1795 3626 2007 3630
rect 2011 3626 2019 3630
rect 91 3625 2019 3626
rect 2025 3625 2026 3631
rect 2030 3613 2031 3619
rect 2037 3618 3979 3619
rect 2037 3614 2047 3618
rect 2051 3614 2127 3618
rect 2131 3614 2191 3618
rect 2195 3614 2327 3618
rect 2331 3614 2351 3618
rect 2355 3614 2455 3618
rect 2459 3614 2583 3618
rect 2587 3614 2719 3618
rect 2723 3614 2815 3618
rect 2819 3614 2855 3618
rect 2859 3614 2999 3618
rect 3003 3614 3047 3618
rect 3051 3614 3143 3618
rect 3147 3614 3279 3618
rect 3283 3614 3295 3618
rect 3299 3614 3455 3618
rect 3459 3614 3511 3618
rect 3515 3614 3623 3618
rect 3627 3614 3751 3618
rect 3755 3614 3943 3618
rect 3947 3614 3979 3618
rect 2037 3613 3979 3614
rect 3985 3613 3986 3619
rect 2018 3547 2019 3553
rect 2025 3547 2050 3553
rect 2044 3543 2050 3547
rect 96 3537 97 3543
rect 103 3542 2031 3543
rect 103 3538 111 3542
rect 115 3538 159 3542
rect 163 3538 303 3542
rect 307 3538 335 3542
rect 339 3538 463 3542
rect 467 3538 607 3542
rect 611 3538 639 3542
rect 643 3538 759 3542
rect 763 3538 815 3542
rect 819 3538 927 3542
rect 931 3538 999 3542
rect 1003 3538 1095 3542
rect 1099 3538 1175 3542
rect 1179 3538 1263 3542
rect 1267 3538 1351 3542
rect 1355 3538 1439 3542
rect 1443 3538 1527 3542
rect 1531 3538 1615 3542
rect 1619 3538 1703 3542
rect 1707 3538 1791 3542
rect 1795 3538 1879 3542
rect 1883 3538 2007 3542
rect 2011 3538 2031 3542
rect 103 3537 2031 3538
rect 2037 3537 2038 3543
rect 2044 3542 3967 3543
rect 2044 3538 2047 3542
rect 2051 3538 2103 3542
rect 2107 3538 2191 3542
rect 2195 3538 2271 3542
rect 2275 3538 2327 3542
rect 2331 3538 2447 3542
rect 2451 3538 2455 3542
rect 2459 3538 2583 3542
rect 2587 3538 2631 3542
rect 2635 3538 2719 3542
rect 2723 3538 2815 3542
rect 2819 3538 2855 3542
rect 2859 3538 2999 3542
rect 3003 3538 3143 3542
rect 3147 3538 3175 3542
rect 3179 3538 3295 3542
rect 3299 3538 3351 3542
rect 3355 3538 3455 3542
rect 3459 3538 3519 3542
rect 3523 3538 3623 3542
rect 3627 3538 3687 3542
rect 3691 3538 3839 3542
rect 3843 3538 3943 3542
rect 3947 3538 3967 3542
rect 2044 3537 3967 3538
rect 3973 3537 3974 3543
rect 84 3453 85 3459
rect 91 3458 2019 3459
rect 91 3454 111 3458
rect 115 3454 135 3458
rect 139 3454 159 3458
rect 163 3454 303 3458
rect 307 3454 319 3458
rect 323 3454 463 3458
rect 467 3454 535 3458
rect 539 3454 639 3458
rect 643 3454 751 3458
rect 755 3454 815 3458
rect 819 3454 959 3458
rect 963 3454 999 3458
rect 1003 3454 1159 3458
rect 1163 3454 1175 3458
rect 1179 3454 1351 3458
rect 1355 3454 1527 3458
rect 1531 3454 1535 3458
rect 1539 3454 1703 3458
rect 1707 3454 1719 3458
rect 1723 3454 1879 3458
rect 1883 3454 1903 3458
rect 1907 3454 2007 3458
rect 2011 3454 2019 3458
rect 91 3453 2019 3454
rect 2025 3453 2026 3459
rect 2030 3457 2031 3463
rect 2037 3462 3979 3463
rect 2037 3458 2047 3462
rect 2051 3458 2103 3462
rect 2107 3458 2127 3462
rect 2131 3458 2271 3462
rect 2275 3458 2311 3462
rect 2315 3458 2447 3462
rect 2451 3458 2495 3462
rect 2499 3458 2631 3462
rect 2635 3458 2679 3462
rect 2683 3458 2815 3462
rect 2819 3458 2863 3462
rect 2867 3458 2999 3462
rect 3003 3458 3047 3462
rect 3051 3458 3175 3462
rect 3179 3458 3223 3462
rect 3227 3458 3351 3462
rect 3355 3458 3407 3462
rect 3411 3458 3519 3462
rect 3523 3458 3591 3462
rect 3595 3458 3687 3462
rect 3691 3458 3775 3462
rect 3779 3458 3839 3462
rect 3843 3458 3943 3462
rect 3947 3458 3979 3462
rect 2037 3457 3979 3458
rect 3985 3457 3986 3463
rect 254 3428 260 3429
rect 798 3428 804 3429
rect 254 3424 255 3428
rect 259 3424 799 3428
rect 803 3424 804 3428
rect 254 3423 260 3424
rect 798 3423 804 3424
rect 96 3377 97 3383
rect 103 3382 2031 3383
rect 103 3378 111 3382
rect 115 3378 135 3382
rect 139 3378 231 3382
rect 235 3378 319 3382
rect 323 3378 375 3382
rect 379 3378 535 3382
rect 539 3378 703 3382
rect 707 3378 751 3382
rect 755 3378 871 3382
rect 875 3378 959 3382
rect 963 3378 1047 3382
rect 1051 3378 1159 3382
rect 1163 3378 1215 3382
rect 1219 3378 1351 3382
rect 1355 3378 1383 3382
rect 1387 3378 1535 3382
rect 1539 3378 1543 3382
rect 1547 3378 1703 3382
rect 1707 3378 1719 3382
rect 1723 3378 1871 3382
rect 1875 3378 1903 3382
rect 1907 3378 2007 3382
rect 2011 3378 2031 3382
rect 103 3377 2031 3378
rect 2037 3377 2038 3383
rect 2018 3365 2019 3371
rect 2025 3370 3967 3371
rect 2025 3366 2047 3370
rect 2051 3366 2071 3370
rect 2075 3366 2127 3370
rect 2131 3366 2215 3370
rect 2219 3366 2311 3370
rect 2315 3366 2359 3370
rect 2363 3366 2495 3370
rect 2499 3366 2511 3370
rect 2515 3366 2655 3370
rect 2659 3366 2679 3370
rect 2683 3366 2799 3370
rect 2803 3366 2863 3370
rect 2867 3366 2935 3370
rect 2939 3366 3047 3370
rect 3051 3366 3079 3370
rect 3083 3366 3223 3370
rect 3227 3366 3375 3370
rect 3379 3366 3407 3370
rect 3411 3366 3535 3370
rect 3539 3366 3591 3370
rect 3595 3366 3695 3370
rect 3699 3366 3775 3370
rect 3779 3366 3839 3370
rect 3843 3366 3943 3370
rect 3947 3366 3967 3370
rect 2025 3365 3967 3366
rect 3973 3365 3974 3371
rect 3298 3308 3304 3309
rect 3506 3308 3512 3309
rect 84 3301 85 3307
rect 91 3306 2019 3307
rect 91 3302 111 3306
rect 115 3302 135 3306
rect 139 3302 231 3306
rect 235 3302 279 3306
rect 283 3302 375 3306
rect 379 3302 463 3306
rect 467 3302 535 3306
rect 539 3302 663 3306
rect 667 3302 703 3306
rect 707 3302 871 3306
rect 875 3302 1047 3306
rect 1051 3302 1079 3306
rect 1083 3302 1215 3306
rect 1219 3302 1295 3306
rect 1299 3302 1383 3306
rect 1387 3302 1519 3306
rect 1523 3302 1543 3306
rect 1547 3302 1703 3306
rect 1707 3302 1743 3306
rect 1747 3302 1871 3306
rect 1875 3302 2007 3306
rect 2011 3302 2019 3306
rect 91 3301 2019 3302
rect 2025 3301 2026 3307
rect 3298 3304 3299 3308
rect 3303 3304 3507 3308
rect 3511 3304 3512 3308
rect 3298 3303 3304 3304
rect 3506 3303 3512 3304
rect 2030 3281 2031 3287
rect 2037 3286 3979 3287
rect 2037 3282 2047 3286
rect 2051 3282 2071 3286
rect 2075 3282 2111 3286
rect 2115 3282 2215 3286
rect 2219 3282 2247 3286
rect 2251 3282 2359 3286
rect 2363 3282 2399 3286
rect 2403 3282 2511 3286
rect 2515 3282 2575 3286
rect 2579 3282 2655 3286
rect 2659 3282 2783 3286
rect 2787 3282 2799 3286
rect 2803 3282 2935 3286
rect 2939 3282 3015 3286
rect 3019 3282 3079 3286
rect 3083 3282 3223 3286
rect 3227 3282 3263 3286
rect 3267 3282 3375 3286
rect 3379 3282 3527 3286
rect 3531 3282 3535 3286
rect 3539 3282 3695 3286
rect 3699 3282 3791 3286
rect 3795 3282 3839 3286
rect 3843 3282 3943 3286
rect 3947 3282 3979 3286
rect 2037 3281 3979 3282
rect 3985 3281 3986 3287
rect 96 3225 97 3231
rect 103 3230 2031 3231
rect 103 3226 111 3230
rect 115 3226 135 3230
rect 139 3226 279 3230
rect 283 3226 287 3230
rect 291 3226 447 3230
rect 451 3226 463 3230
rect 467 3226 615 3230
rect 619 3226 663 3230
rect 667 3226 791 3230
rect 795 3226 871 3230
rect 875 3226 967 3230
rect 971 3226 1079 3230
rect 1083 3226 1143 3230
rect 1147 3226 1295 3230
rect 1299 3226 1327 3230
rect 1331 3226 1511 3230
rect 1515 3226 1519 3230
rect 1523 3226 1695 3230
rect 1699 3226 1743 3230
rect 1747 3226 2007 3230
rect 2011 3226 2031 3230
rect 103 3225 2031 3226
rect 2037 3225 2038 3231
rect 2018 3205 2019 3211
rect 2025 3210 3967 3211
rect 2025 3206 2047 3210
rect 2051 3206 2071 3210
rect 2075 3206 2111 3210
rect 2115 3206 2167 3210
rect 2171 3206 2247 3210
rect 2251 3206 2263 3210
rect 2267 3206 2359 3210
rect 2363 3206 2399 3210
rect 2403 3206 2455 3210
rect 2459 3206 2551 3210
rect 2555 3206 2575 3210
rect 2579 3206 2647 3210
rect 2651 3206 2743 3210
rect 2747 3206 2783 3210
rect 2787 3206 2839 3210
rect 2843 3206 2935 3210
rect 2939 3206 3015 3210
rect 3019 3206 3031 3210
rect 3035 3206 3127 3210
rect 3131 3206 3223 3210
rect 3227 3206 3263 3210
rect 3267 3206 3319 3210
rect 3323 3206 3439 3210
rect 3443 3206 3527 3210
rect 3531 3206 3575 3210
rect 3579 3206 3719 3210
rect 3723 3206 3791 3210
rect 3795 3206 3839 3210
rect 3843 3206 3943 3210
rect 3947 3206 3967 3210
rect 2025 3205 3967 3206
rect 3973 3205 3974 3211
rect 84 3145 85 3151
rect 91 3150 2019 3151
rect 91 3146 111 3150
rect 115 3146 135 3150
rect 139 3146 287 3150
rect 291 3146 311 3150
rect 315 3146 439 3150
rect 443 3146 447 3150
rect 451 3146 583 3150
rect 587 3146 615 3150
rect 619 3146 743 3150
rect 747 3146 791 3150
rect 795 3146 903 3150
rect 907 3146 967 3150
rect 971 3146 1063 3150
rect 1067 3146 1143 3150
rect 1147 3146 1223 3150
rect 1227 3146 1327 3150
rect 1331 3146 1391 3150
rect 1395 3146 1511 3150
rect 1515 3146 1559 3150
rect 1563 3146 1695 3150
rect 1699 3146 1727 3150
rect 1731 3146 2007 3150
rect 2011 3146 2019 3150
rect 91 3145 2019 3146
rect 2025 3145 2026 3151
rect 2030 3117 2031 3123
rect 2037 3122 3979 3123
rect 2037 3118 2047 3122
rect 2051 3118 2071 3122
rect 2075 3118 2167 3122
rect 2171 3118 2263 3122
rect 2267 3118 2335 3122
rect 2339 3118 2359 3122
rect 2363 3118 2455 3122
rect 2459 3118 2551 3122
rect 2555 3118 2623 3122
rect 2627 3118 2647 3122
rect 2651 3118 2743 3122
rect 2747 3118 2839 3122
rect 2843 3118 2911 3122
rect 2915 3118 2935 3122
rect 2939 3118 3031 3122
rect 3035 3118 3127 3122
rect 3131 3118 3207 3122
rect 3211 3118 3223 3122
rect 3227 3118 3319 3122
rect 3323 3118 3439 3122
rect 3443 3118 3503 3122
rect 3507 3118 3575 3122
rect 3579 3118 3719 3122
rect 3723 3118 3799 3122
rect 3803 3118 3839 3122
rect 3843 3118 3943 3122
rect 3947 3118 3979 3122
rect 2037 3117 3979 3118
rect 3985 3117 3986 3123
rect 96 3061 97 3067
rect 103 3066 2031 3067
rect 103 3062 111 3066
rect 115 3062 311 3066
rect 315 3062 439 3066
rect 443 3062 503 3066
rect 507 3062 583 3066
rect 587 3062 599 3066
rect 603 3062 703 3066
rect 707 3062 743 3066
rect 747 3062 815 3066
rect 819 3062 903 3066
rect 907 3062 935 3066
rect 939 3062 1063 3066
rect 1067 3062 1071 3066
rect 1075 3062 1223 3066
rect 1227 3062 1383 3066
rect 1387 3062 1391 3066
rect 1395 3062 1551 3066
rect 1555 3062 1559 3066
rect 1563 3062 1719 3066
rect 1723 3062 1727 3066
rect 1731 3062 2007 3066
rect 2011 3062 2031 3066
rect 103 3061 2031 3062
rect 2037 3061 2038 3067
rect 2018 3041 2019 3047
rect 2025 3046 3967 3047
rect 2025 3042 2047 3046
rect 2051 3042 2071 3046
rect 2075 3042 2335 3046
rect 2339 3042 2383 3046
rect 2387 3042 2623 3046
rect 2627 3042 2703 3046
rect 2707 3042 2911 3046
rect 2915 3042 2999 3046
rect 3003 3042 3207 3046
rect 3211 3042 3287 3046
rect 3291 3042 3503 3046
rect 3507 3042 3575 3046
rect 3579 3042 3799 3046
rect 3803 3042 3839 3046
rect 3843 3042 3943 3046
rect 3947 3042 3967 3046
rect 2025 3041 3967 3042
rect 3973 3041 3974 3047
rect 84 2981 85 2987
rect 91 2986 2019 2987
rect 91 2982 111 2986
rect 115 2982 503 2986
rect 507 2982 551 2986
rect 555 2982 599 2986
rect 603 2982 647 2986
rect 651 2982 703 2986
rect 707 2982 759 2986
rect 763 2982 815 2986
rect 819 2982 887 2986
rect 891 2982 935 2986
rect 939 2982 1023 2986
rect 1027 2982 1071 2986
rect 1075 2982 1175 2986
rect 1179 2982 1223 2986
rect 1227 2982 1327 2986
rect 1331 2982 1383 2986
rect 1387 2982 1487 2986
rect 1491 2982 1551 2986
rect 1555 2982 1655 2986
rect 1659 2982 1719 2986
rect 1723 2982 1823 2986
rect 1827 2982 2007 2986
rect 2011 2982 2019 2986
rect 91 2981 2019 2982
rect 2025 2981 2026 2987
rect 2030 2961 2031 2967
rect 2037 2966 3979 2967
rect 2037 2962 2047 2966
rect 2051 2962 2071 2966
rect 2075 2962 2383 2966
rect 2387 2962 2391 2966
rect 2395 2962 2703 2966
rect 2707 2962 2975 2966
rect 2979 2962 2999 2966
rect 3003 2962 3215 2966
rect 3219 2962 3287 2966
rect 3291 2962 3439 2966
rect 3443 2962 3575 2966
rect 3579 2962 3647 2966
rect 3651 2962 3839 2966
rect 3843 2962 3943 2966
rect 3947 2962 3979 2966
rect 2037 2961 3979 2962
rect 3985 2961 3986 2967
rect 96 2897 97 2903
rect 103 2902 2031 2903
rect 103 2898 111 2902
rect 115 2898 471 2902
rect 475 2898 551 2902
rect 555 2898 575 2902
rect 579 2898 647 2902
rect 651 2898 695 2902
rect 699 2898 759 2902
rect 763 2898 839 2902
rect 843 2898 887 2902
rect 891 2898 991 2902
rect 995 2898 1023 2902
rect 1027 2898 1151 2902
rect 1155 2898 1175 2902
rect 1179 2898 1319 2902
rect 1323 2898 1327 2902
rect 1331 2898 1487 2902
rect 1491 2898 1495 2902
rect 1499 2898 1655 2902
rect 1659 2898 1671 2902
rect 1675 2898 1823 2902
rect 1827 2898 1847 2902
rect 1851 2898 2007 2902
rect 2011 2898 2031 2902
rect 103 2897 2031 2898
rect 2037 2897 2038 2903
rect 2018 2885 2019 2891
rect 2025 2890 3967 2891
rect 2025 2886 2047 2890
rect 2051 2886 2071 2890
rect 2075 2886 2295 2890
rect 2299 2886 2391 2890
rect 2395 2886 2535 2890
rect 2539 2886 2703 2890
rect 2707 2886 2767 2890
rect 2771 2886 2975 2890
rect 2979 2886 2991 2890
rect 2995 2886 3215 2890
rect 3219 2886 3431 2890
rect 3435 2886 3439 2890
rect 3443 2886 3647 2890
rect 3651 2886 3839 2890
rect 3843 2886 3943 2890
rect 3947 2886 3967 2890
rect 2025 2885 3967 2886
rect 3973 2885 3974 2891
rect 84 2817 85 2823
rect 91 2822 2019 2823
rect 91 2818 111 2822
rect 115 2818 471 2822
rect 475 2818 479 2822
rect 483 2818 575 2822
rect 579 2818 679 2822
rect 683 2818 695 2822
rect 699 2818 799 2822
rect 803 2818 839 2822
rect 843 2818 935 2822
rect 939 2818 991 2822
rect 995 2818 1079 2822
rect 1083 2818 1151 2822
rect 1155 2818 1239 2822
rect 1243 2818 1319 2822
rect 1323 2818 1415 2822
rect 1419 2818 1495 2822
rect 1499 2818 1599 2822
rect 1603 2818 1671 2822
rect 1675 2818 1783 2822
rect 1787 2818 1847 2822
rect 1851 2818 2007 2822
rect 2011 2818 2019 2822
rect 91 2817 2019 2818
rect 2025 2817 2026 2823
rect 2030 2805 2031 2811
rect 2037 2810 3979 2811
rect 2037 2806 2047 2810
rect 2051 2806 2071 2810
rect 2075 2806 2199 2810
rect 2203 2806 2295 2810
rect 2299 2806 2367 2810
rect 2371 2806 2535 2810
rect 2539 2806 2551 2810
rect 2555 2806 2735 2810
rect 2739 2806 2767 2810
rect 2771 2806 2927 2810
rect 2931 2806 2991 2810
rect 2995 2806 3111 2810
rect 3115 2806 3215 2810
rect 3219 2806 3295 2810
rect 3299 2806 3431 2810
rect 3435 2806 3479 2810
rect 3483 2806 3647 2810
rect 3651 2806 3671 2810
rect 3675 2806 3839 2810
rect 3843 2806 3943 2810
rect 3947 2806 3979 2810
rect 2037 2805 3979 2806
rect 3985 2805 3986 2811
rect 96 2737 97 2743
rect 103 2742 2031 2743
rect 103 2738 111 2742
rect 115 2738 479 2742
rect 483 2738 511 2742
rect 515 2738 575 2742
rect 579 2738 623 2742
rect 627 2738 679 2742
rect 683 2738 743 2742
rect 747 2738 799 2742
rect 803 2738 879 2742
rect 883 2738 935 2742
rect 939 2738 1015 2742
rect 1019 2738 1079 2742
rect 1083 2738 1159 2742
rect 1163 2738 1239 2742
rect 1243 2738 1311 2742
rect 1315 2738 1415 2742
rect 1419 2738 1463 2742
rect 1467 2738 1599 2742
rect 1603 2738 1623 2742
rect 1627 2738 1783 2742
rect 1787 2738 2007 2742
rect 2011 2738 2031 2742
rect 103 2737 2031 2738
rect 2037 2737 2038 2743
rect 2018 2725 2019 2731
rect 2025 2730 3967 2731
rect 2025 2726 2047 2730
rect 2051 2726 2071 2730
rect 2075 2726 2191 2730
rect 2195 2726 2199 2730
rect 2203 2726 2319 2730
rect 2323 2726 2367 2730
rect 2371 2726 2447 2730
rect 2451 2726 2551 2730
rect 2555 2726 2583 2730
rect 2587 2726 2727 2730
rect 2731 2726 2735 2730
rect 2739 2726 2887 2730
rect 2891 2726 2927 2730
rect 2931 2726 3063 2730
rect 3067 2726 3111 2730
rect 3115 2726 3255 2730
rect 3259 2726 3295 2730
rect 3299 2726 3455 2730
rect 3459 2726 3479 2730
rect 3483 2726 3655 2730
rect 3659 2726 3671 2730
rect 3675 2726 3839 2730
rect 3843 2726 3943 2730
rect 3947 2726 3967 2730
rect 2025 2725 3967 2726
rect 3973 2725 3974 2731
rect 84 2657 85 2663
rect 91 2662 2019 2663
rect 91 2658 111 2662
rect 115 2658 367 2662
rect 371 2658 487 2662
rect 491 2658 511 2662
rect 515 2658 615 2662
rect 619 2658 623 2662
rect 627 2658 743 2662
rect 747 2658 751 2662
rect 755 2658 879 2662
rect 883 2658 895 2662
rect 899 2658 1015 2662
rect 1019 2658 1031 2662
rect 1035 2658 1159 2662
rect 1163 2658 1167 2662
rect 1171 2658 1303 2662
rect 1307 2658 1311 2662
rect 1315 2658 1431 2662
rect 1435 2658 1463 2662
rect 1467 2658 1567 2662
rect 1571 2658 1623 2662
rect 1627 2658 1703 2662
rect 1707 2658 1783 2662
rect 1787 2658 2007 2662
rect 2011 2658 2019 2662
rect 91 2657 2019 2658
rect 2025 2657 2026 2663
rect 2030 2641 2031 2647
rect 2037 2646 3979 2647
rect 2037 2642 2047 2646
rect 2051 2642 2071 2646
rect 2075 2642 2191 2646
rect 2195 2642 2231 2646
rect 2235 2642 2319 2646
rect 2323 2642 2335 2646
rect 2339 2642 2447 2646
rect 2451 2642 2559 2646
rect 2563 2642 2583 2646
rect 2587 2642 2671 2646
rect 2675 2642 2727 2646
rect 2731 2642 2791 2646
rect 2795 2642 2887 2646
rect 2891 2642 2911 2646
rect 2915 2642 3031 2646
rect 3035 2642 3063 2646
rect 3067 2642 3151 2646
rect 3155 2642 3255 2646
rect 3259 2642 3455 2646
rect 3459 2642 3655 2646
rect 3659 2642 3839 2646
rect 3843 2642 3943 2646
rect 3947 2642 3979 2646
rect 2037 2641 3979 2642
rect 3985 2641 3986 2647
rect 96 2581 97 2587
rect 103 2586 2031 2587
rect 103 2582 111 2586
rect 115 2582 135 2586
rect 139 2582 287 2586
rect 291 2582 367 2586
rect 371 2582 447 2586
rect 451 2582 487 2586
rect 491 2582 607 2586
rect 611 2582 615 2586
rect 619 2582 751 2586
rect 755 2582 767 2586
rect 771 2582 895 2586
rect 899 2582 919 2586
rect 923 2582 1031 2586
rect 1035 2582 1063 2586
rect 1067 2582 1167 2586
rect 1171 2582 1199 2586
rect 1203 2582 1303 2586
rect 1307 2582 1335 2586
rect 1339 2582 1431 2586
rect 1435 2582 1463 2586
rect 1467 2582 1567 2586
rect 1571 2582 1591 2586
rect 1595 2582 1703 2586
rect 1707 2582 1727 2586
rect 1731 2582 2007 2586
rect 2011 2582 2031 2586
rect 103 2581 2031 2582
rect 2037 2581 2038 2587
rect 2018 2561 2019 2567
rect 2025 2566 3967 2567
rect 2025 2562 2047 2566
rect 2051 2562 2231 2566
rect 2235 2562 2335 2566
rect 2339 2562 2383 2566
rect 2387 2562 2447 2566
rect 2451 2562 2495 2566
rect 2499 2562 2559 2566
rect 2563 2562 2615 2566
rect 2619 2562 2671 2566
rect 2675 2562 2743 2566
rect 2747 2562 2791 2566
rect 2795 2562 2871 2566
rect 2875 2562 2911 2566
rect 2915 2562 2991 2566
rect 2995 2562 3031 2566
rect 3035 2562 3111 2566
rect 3115 2562 3151 2566
rect 3155 2562 3231 2566
rect 3235 2562 3359 2566
rect 3363 2562 3487 2566
rect 3491 2562 3943 2566
rect 3947 2562 3967 2566
rect 2025 2561 3967 2562
rect 3973 2561 3974 2567
rect 84 2489 85 2495
rect 91 2494 2019 2495
rect 91 2490 111 2494
rect 115 2490 135 2494
rect 139 2490 231 2494
rect 235 2490 287 2494
rect 291 2490 327 2494
rect 331 2490 423 2494
rect 427 2490 447 2494
rect 451 2490 519 2494
rect 523 2490 607 2494
rect 611 2490 767 2494
rect 771 2490 919 2494
rect 923 2490 1063 2494
rect 1067 2490 1199 2494
rect 1203 2490 1335 2494
rect 1339 2490 1463 2494
rect 1467 2490 1591 2494
rect 1595 2490 1727 2494
rect 1731 2490 2007 2494
rect 2011 2490 2019 2494
rect 91 2489 2019 2490
rect 2025 2489 2026 2495
rect 2030 2481 2031 2487
rect 2037 2486 3979 2487
rect 2037 2482 2047 2486
rect 2051 2482 2383 2486
rect 2387 2482 2495 2486
rect 2499 2482 2535 2486
rect 2539 2482 2615 2486
rect 2619 2482 2711 2486
rect 2715 2482 2743 2486
rect 2747 2482 2871 2486
rect 2875 2482 2879 2486
rect 2883 2482 2991 2486
rect 2995 2482 3047 2486
rect 3051 2482 3111 2486
rect 3115 2482 3207 2486
rect 3211 2482 3231 2486
rect 3235 2482 3359 2486
rect 3363 2482 3487 2486
rect 3491 2482 3503 2486
rect 3507 2482 3655 2486
rect 3659 2482 3807 2486
rect 3811 2482 3943 2486
rect 3947 2482 3979 2486
rect 2037 2481 3979 2482
rect 3985 2481 3986 2487
rect 2018 2407 2019 2413
rect 2025 2407 2050 2413
rect 96 2397 97 2403
rect 103 2402 2031 2403
rect 103 2398 111 2402
rect 115 2398 135 2402
rect 139 2398 231 2402
rect 235 2398 255 2402
rect 259 2398 327 2402
rect 331 2398 415 2402
rect 419 2398 423 2402
rect 427 2398 519 2402
rect 523 2398 575 2402
rect 579 2398 735 2402
rect 739 2398 887 2402
rect 891 2398 1039 2402
rect 1043 2398 1183 2402
rect 1187 2398 1327 2402
rect 1331 2398 1479 2402
rect 1483 2398 2007 2402
rect 2011 2398 2031 2402
rect 103 2397 2031 2398
rect 2037 2397 2038 2403
rect 2044 2399 2050 2407
rect 2044 2398 3967 2399
rect 2044 2394 2047 2398
rect 2051 2394 2535 2398
rect 2539 2394 2607 2398
rect 2611 2394 2711 2398
rect 2715 2394 2815 2398
rect 2819 2394 2879 2398
rect 2883 2394 3007 2398
rect 3011 2394 3047 2398
rect 3051 2394 3191 2398
rect 3195 2394 3207 2398
rect 3211 2394 3359 2398
rect 3363 2394 3503 2398
rect 3507 2394 3519 2398
rect 3523 2394 3655 2398
rect 3659 2394 3679 2398
rect 3683 2394 3807 2398
rect 3811 2394 3839 2398
rect 3843 2394 3943 2398
rect 3947 2394 3967 2398
rect 2044 2393 3967 2394
rect 3973 2393 3974 2399
rect 84 2321 85 2327
rect 91 2326 2019 2327
rect 91 2322 111 2326
rect 115 2322 135 2326
rect 139 2322 255 2326
rect 259 2322 263 2326
rect 267 2322 415 2326
rect 419 2322 423 2326
rect 427 2322 575 2326
rect 579 2322 583 2326
rect 587 2322 735 2326
rect 739 2322 743 2326
rect 747 2322 887 2326
rect 891 2322 895 2326
rect 899 2322 1039 2326
rect 1043 2322 1047 2326
rect 1051 2322 1183 2326
rect 1187 2322 1199 2326
rect 1203 2322 1327 2326
rect 1331 2322 1351 2326
rect 1355 2322 1479 2326
rect 1483 2322 1503 2326
rect 1507 2322 2007 2326
rect 2011 2322 2019 2326
rect 91 2321 2019 2322
rect 2025 2321 2026 2327
rect 2030 2301 2031 2307
rect 2037 2306 3979 2307
rect 2037 2302 2047 2306
rect 2051 2302 2071 2306
rect 2075 2302 2167 2306
rect 2171 2302 2271 2306
rect 2275 2302 2415 2306
rect 2419 2302 2575 2306
rect 2579 2302 2607 2306
rect 2611 2302 2743 2306
rect 2747 2302 2815 2306
rect 2819 2302 2911 2306
rect 2915 2302 3007 2306
rect 3011 2302 3071 2306
rect 3075 2302 3191 2306
rect 3195 2302 3231 2306
rect 3235 2302 3359 2306
rect 3363 2302 3383 2306
rect 3387 2302 3519 2306
rect 3523 2302 3535 2306
rect 3539 2302 3679 2306
rect 3683 2302 3695 2306
rect 3699 2302 3839 2306
rect 3843 2302 3943 2306
rect 3947 2302 3979 2306
rect 2037 2301 3979 2302
rect 3985 2301 3986 2307
rect 96 2241 97 2247
rect 103 2246 2031 2247
rect 103 2242 111 2246
rect 115 2242 135 2246
rect 139 2242 223 2246
rect 227 2242 263 2246
rect 267 2242 351 2246
rect 355 2242 423 2246
rect 427 2242 495 2246
rect 499 2242 583 2246
rect 587 2242 647 2246
rect 651 2242 743 2246
rect 747 2242 799 2246
rect 803 2242 895 2246
rect 899 2242 959 2246
rect 963 2242 1047 2246
rect 1051 2242 1119 2246
rect 1123 2242 1199 2246
rect 1203 2242 1279 2246
rect 1283 2242 1351 2246
rect 1355 2242 1439 2246
rect 1443 2242 1503 2246
rect 1507 2242 1599 2246
rect 1603 2242 2007 2246
rect 2011 2242 2031 2246
rect 103 2241 2031 2242
rect 2037 2241 2038 2247
rect 2018 2225 2019 2231
rect 2025 2230 3967 2231
rect 2025 2226 2047 2230
rect 2051 2226 2071 2230
rect 2075 2226 2167 2230
rect 2171 2226 2175 2230
rect 2179 2226 2271 2230
rect 2275 2226 2319 2230
rect 2323 2226 2415 2230
rect 2419 2226 2471 2230
rect 2475 2226 2575 2230
rect 2579 2226 2623 2230
rect 2627 2226 2743 2230
rect 2747 2226 2783 2230
rect 2787 2226 2911 2230
rect 2915 2226 2935 2230
rect 2939 2226 3071 2230
rect 3075 2226 3079 2230
rect 3083 2226 3223 2230
rect 3227 2226 3231 2230
rect 3235 2226 3367 2230
rect 3371 2226 3383 2230
rect 3387 2226 3519 2230
rect 3523 2226 3535 2230
rect 3539 2226 3695 2230
rect 3699 2226 3943 2230
rect 3947 2226 3967 2230
rect 2025 2225 3967 2226
rect 3973 2225 3974 2231
rect 84 2165 85 2171
rect 91 2170 2019 2171
rect 91 2166 111 2170
rect 115 2166 223 2170
rect 227 2166 351 2170
rect 355 2166 471 2170
rect 475 2166 495 2170
rect 499 2166 567 2170
rect 571 2166 647 2170
rect 651 2166 679 2170
rect 683 2166 799 2170
rect 803 2166 807 2170
rect 811 2166 943 2170
rect 947 2166 959 2170
rect 963 2166 1079 2170
rect 1083 2166 1119 2170
rect 1123 2166 1223 2170
rect 1227 2166 1279 2170
rect 1283 2166 1367 2170
rect 1371 2166 1439 2170
rect 1443 2166 1503 2170
rect 1507 2166 1599 2170
rect 1603 2166 1639 2170
rect 1643 2166 1783 2170
rect 1787 2166 1903 2170
rect 1907 2166 2007 2170
rect 2011 2166 2019 2170
rect 91 2165 2019 2166
rect 2025 2165 2026 2171
rect 2030 2129 2031 2135
rect 2037 2134 3979 2135
rect 2037 2130 2047 2134
rect 2051 2130 2071 2134
rect 2075 2130 2175 2134
rect 2179 2130 2279 2134
rect 2283 2130 2319 2134
rect 2323 2130 2391 2134
rect 2395 2130 2471 2134
rect 2475 2130 2511 2134
rect 2515 2130 2623 2134
rect 2627 2130 2631 2134
rect 2635 2130 2759 2134
rect 2763 2130 2783 2134
rect 2787 2130 2895 2134
rect 2899 2130 2935 2134
rect 2939 2130 3039 2134
rect 3043 2130 3079 2134
rect 3083 2130 3191 2134
rect 3195 2130 3223 2134
rect 3227 2130 3351 2134
rect 3355 2130 3367 2134
rect 3371 2130 3519 2134
rect 3523 2130 3687 2134
rect 3691 2130 3839 2134
rect 3843 2130 3943 2134
rect 3947 2130 3979 2134
rect 2037 2129 3979 2130
rect 3985 2129 3986 2135
rect 96 2089 97 2095
rect 103 2094 2031 2095
rect 103 2090 111 2094
rect 115 2090 471 2094
rect 475 2090 567 2094
rect 571 2090 623 2094
rect 627 2090 679 2094
rect 683 2090 735 2094
rect 739 2090 807 2094
rect 811 2090 855 2094
rect 859 2090 943 2094
rect 947 2090 983 2094
rect 987 2090 1079 2094
rect 1083 2090 1119 2094
rect 1123 2090 1223 2094
rect 1227 2090 1255 2094
rect 1259 2090 1367 2094
rect 1371 2090 1391 2094
rect 1395 2090 1503 2094
rect 1507 2090 1527 2094
rect 1531 2090 1639 2094
rect 1643 2090 1655 2094
rect 1659 2090 1783 2094
rect 1787 2090 1791 2094
rect 1795 2090 1903 2094
rect 1907 2090 2007 2094
rect 2011 2090 2031 2094
rect 103 2089 2031 2090
rect 2037 2089 2038 2095
rect 2018 2045 2019 2051
rect 2025 2050 3967 2051
rect 2025 2046 2047 2050
rect 2051 2046 2279 2050
rect 2283 2046 2327 2050
rect 2331 2046 2391 2050
rect 2395 2046 2431 2050
rect 2435 2046 2511 2050
rect 2515 2046 2535 2050
rect 2539 2046 2631 2050
rect 2635 2046 2647 2050
rect 2651 2046 2759 2050
rect 2763 2046 2775 2050
rect 2779 2046 2895 2050
rect 2899 2046 2919 2050
rect 2923 2046 3039 2050
rect 3043 2046 3079 2050
rect 3083 2046 3191 2050
rect 3195 2046 3263 2050
rect 3267 2046 3351 2050
rect 3355 2046 3455 2050
rect 3459 2046 3519 2050
rect 3523 2046 3655 2050
rect 3659 2046 3687 2050
rect 3691 2046 3839 2050
rect 3843 2046 3943 2050
rect 3947 2046 3967 2050
rect 2025 2045 3967 2046
rect 3973 2045 3974 2051
rect 84 2009 85 2015
rect 91 2014 2019 2015
rect 91 2010 111 2014
rect 115 2010 447 2014
rect 451 2010 575 2014
rect 579 2010 623 2014
rect 627 2010 727 2014
rect 731 2010 735 2014
rect 739 2010 855 2014
rect 859 2010 887 2014
rect 891 2010 983 2014
rect 987 2010 1055 2014
rect 1059 2010 1119 2014
rect 1123 2010 1231 2014
rect 1235 2010 1255 2014
rect 1259 2010 1391 2014
rect 1395 2010 1399 2014
rect 1403 2010 1527 2014
rect 1531 2010 1575 2014
rect 1579 2010 1655 2014
rect 1659 2010 1751 2014
rect 1755 2010 1791 2014
rect 1795 2010 1903 2014
rect 1907 2010 2007 2014
rect 2011 2010 2019 2014
rect 91 2009 2019 2010
rect 2025 2009 2026 2015
rect 2030 1965 2031 1971
rect 2037 1970 3979 1971
rect 2037 1966 2047 1970
rect 2051 1966 2255 1970
rect 2259 1966 2327 1970
rect 2331 1966 2351 1970
rect 2355 1966 2431 1970
rect 2435 1966 2447 1970
rect 2451 1966 2535 1970
rect 2539 1966 2543 1970
rect 2547 1966 2647 1970
rect 2651 1966 2767 1970
rect 2771 1966 2775 1970
rect 2779 1966 2919 1970
rect 2923 1966 3079 1970
rect 3083 1966 3103 1970
rect 3107 1966 3263 1970
rect 3267 1966 3319 1970
rect 3323 1966 3455 1970
rect 3459 1966 3543 1970
rect 3547 1966 3655 1970
rect 3659 1966 3775 1970
rect 3779 1966 3839 1970
rect 3843 1966 3943 1970
rect 3947 1966 3979 1970
rect 2037 1965 3979 1966
rect 3985 1965 3986 1971
rect 96 1933 97 1939
rect 103 1938 2031 1939
rect 103 1934 111 1938
rect 115 1934 447 1938
rect 451 1934 575 1938
rect 579 1934 655 1938
rect 659 1934 727 1938
rect 731 1934 751 1938
rect 755 1934 847 1938
rect 851 1934 887 1938
rect 891 1934 943 1938
rect 947 1934 1039 1938
rect 1043 1934 1055 1938
rect 1059 1934 1135 1938
rect 1139 1934 1231 1938
rect 1235 1934 1327 1938
rect 1331 1934 1399 1938
rect 1403 1934 1423 1938
rect 1427 1934 1575 1938
rect 1579 1934 1751 1938
rect 1755 1934 1903 1938
rect 1907 1934 2007 1938
rect 2011 1934 2031 1938
rect 103 1933 2031 1934
rect 2037 1933 2038 1939
rect 2018 1877 2019 1883
rect 2025 1882 3967 1883
rect 2025 1878 2047 1882
rect 2051 1878 2183 1882
rect 2187 1878 2255 1882
rect 2259 1878 2279 1882
rect 2283 1878 2351 1882
rect 2355 1878 2383 1882
rect 2387 1878 2447 1882
rect 2451 1878 2487 1882
rect 2491 1878 2543 1882
rect 2547 1878 2591 1882
rect 2595 1878 2647 1882
rect 2651 1878 2703 1882
rect 2707 1878 2767 1882
rect 2771 1878 2831 1882
rect 2835 1878 2919 1882
rect 2923 1878 2991 1882
rect 2995 1878 3103 1882
rect 3107 1878 3183 1882
rect 3187 1878 3319 1882
rect 3323 1878 3399 1882
rect 3403 1878 3543 1882
rect 3547 1878 3631 1882
rect 3635 1878 3775 1882
rect 3779 1878 3839 1882
rect 3843 1878 3943 1882
rect 3947 1878 3967 1882
rect 2025 1877 3967 1878
rect 3973 1877 3974 1883
rect 84 1857 85 1863
rect 91 1862 2019 1863
rect 91 1858 111 1862
rect 115 1858 319 1862
rect 323 1858 447 1862
rect 451 1858 583 1862
rect 587 1858 655 1862
rect 659 1858 719 1862
rect 723 1858 751 1862
rect 755 1858 847 1862
rect 851 1858 855 1862
rect 859 1858 943 1862
rect 947 1858 991 1862
rect 995 1858 1039 1862
rect 1043 1858 1127 1862
rect 1131 1858 1135 1862
rect 1139 1858 1231 1862
rect 1235 1858 1263 1862
rect 1267 1858 1327 1862
rect 1331 1858 1399 1862
rect 1403 1858 1423 1862
rect 1427 1858 1535 1862
rect 1539 1858 2007 1862
rect 2011 1858 2019 1862
rect 91 1857 2019 1858
rect 2025 1857 2026 1863
rect 2030 1797 2031 1803
rect 2037 1802 3979 1803
rect 2037 1798 2047 1802
rect 2051 1798 2127 1802
rect 2131 1798 2183 1802
rect 2187 1798 2279 1802
rect 2283 1798 2311 1802
rect 2315 1798 2383 1802
rect 2387 1798 2487 1802
rect 2491 1798 2495 1802
rect 2499 1798 2591 1802
rect 2595 1798 2687 1802
rect 2691 1798 2703 1802
rect 2707 1798 2831 1802
rect 2835 1798 2879 1802
rect 2883 1798 2991 1802
rect 2995 1798 3071 1802
rect 3075 1798 3183 1802
rect 3187 1798 3263 1802
rect 3267 1798 3399 1802
rect 3403 1798 3463 1802
rect 3467 1798 3631 1802
rect 3635 1798 3663 1802
rect 3667 1798 3839 1802
rect 3843 1798 3943 1802
rect 3947 1798 3979 1802
rect 2037 1797 3979 1798
rect 3985 1797 3986 1803
rect 96 1777 97 1783
rect 103 1782 2031 1783
rect 103 1778 111 1782
rect 115 1778 255 1782
rect 259 1778 319 1782
rect 323 1778 391 1782
rect 395 1778 447 1782
rect 451 1778 535 1782
rect 539 1778 583 1782
rect 587 1778 695 1782
rect 699 1778 719 1782
rect 723 1778 855 1782
rect 859 1778 863 1782
rect 867 1778 991 1782
rect 995 1778 1031 1782
rect 1035 1778 1127 1782
rect 1131 1778 1207 1782
rect 1211 1778 1263 1782
rect 1267 1778 1383 1782
rect 1387 1778 1399 1782
rect 1403 1778 1535 1782
rect 1539 1778 1559 1782
rect 1563 1778 1743 1782
rect 1747 1778 2007 1782
rect 2011 1778 2031 1782
rect 103 1777 2031 1778
rect 2037 1777 2038 1783
rect 2018 1717 2019 1723
rect 2025 1722 3967 1723
rect 2025 1718 2047 1722
rect 2051 1718 2071 1722
rect 2075 1718 2127 1722
rect 2131 1718 2191 1722
rect 2195 1718 2311 1722
rect 2315 1718 2343 1722
rect 2347 1718 2495 1722
rect 2499 1718 2511 1722
rect 2515 1718 2687 1722
rect 2691 1718 2871 1722
rect 2875 1718 2879 1722
rect 2883 1718 3063 1722
rect 3067 1718 3071 1722
rect 3075 1718 3255 1722
rect 3259 1718 3263 1722
rect 3267 1718 3447 1722
rect 3451 1718 3463 1722
rect 3467 1718 3647 1722
rect 3651 1718 3663 1722
rect 3667 1718 3839 1722
rect 3843 1718 3943 1722
rect 3947 1718 3967 1722
rect 2025 1717 3967 1718
rect 3973 1717 3974 1723
rect 84 1701 85 1707
rect 91 1706 2019 1707
rect 91 1702 111 1706
rect 115 1702 135 1706
rect 139 1702 255 1706
rect 259 1702 263 1706
rect 267 1702 391 1706
rect 395 1702 431 1706
rect 435 1702 535 1706
rect 539 1702 607 1706
rect 611 1702 695 1706
rect 699 1702 799 1706
rect 803 1702 863 1706
rect 867 1702 999 1706
rect 1003 1702 1031 1706
rect 1035 1702 1199 1706
rect 1203 1702 1207 1706
rect 1211 1702 1383 1706
rect 1387 1702 1407 1706
rect 1411 1702 1559 1706
rect 1563 1702 1623 1706
rect 1627 1702 1743 1706
rect 1747 1702 1839 1706
rect 1843 1702 2007 1706
rect 2011 1702 2019 1706
rect 91 1701 2019 1702
rect 2025 1701 2026 1707
rect 2030 1641 2031 1647
rect 2037 1646 3979 1647
rect 2037 1642 2047 1646
rect 2051 1642 2071 1646
rect 2075 1642 2191 1646
rect 2195 1642 2335 1646
rect 2339 1642 2343 1646
rect 2347 1642 2511 1646
rect 2515 1642 2599 1646
rect 2603 1642 2687 1646
rect 2691 1642 2839 1646
rect 2843 1642 2871 1646
rect 2875 1642 3047 1646
rect 3051 1642 3063 1646
rect 3067 1642 3231 1646
rect 3235 1642 3255 1646
rect 3259 1642 3399 1646
rect 3403 1642 3447 1646
rect 3451 1642 3551 1646
rect 3555 1642 3647 1646
rect 3651 1642 3695 1646
rect 3699 1642 3839 1646
rect 3843 1642 3943 1646
rect 3947 1642 3979 1646
rect 2037 1641 3979 1642
rect 3985 1641 3986 1647
rect 96 1625 97 1631
rect 103 1630 2031 1631
rect 103 1626 111 1630
rect 115 1626 135 1630
rect 139 1626 263 1630
rect 267 1626 287 1630
rect 291 1626 431 1630
rect 435 1626 471 1630
rect 475 1626 607 1630
rect 611 1626 655 1630
rect 659 1626 799 1630
rect 803 1626 839 1630
rect 843 1626 999 1630
rect 1003 1626 1015 1630
rect 1019 1626 1183 1630
rect 1187 1626 1199 1630
rect 1203 1626 1343 1630
rect 1347 1626 1407 1630
rect 1411 1626 1495 1630
rect 1499 1626 1623 1630
rect 1627 1626 1639 1630
rect 1643 1626 1783 1630
rect 1787 1626 1839 1630
rect 1843 1626 1903 1630
rect 1907 1626 2007 1630
rect 2011 1626 2031 1630
rect 103 1625 2031 1626
rect 2037 1625 2038 1631
rect 2018 1561 2019 1567
rect 2025 1566 3967 1567
rect 2025 1562 2047 1566
rect 2051 1562 2071 1566
rect 2075 1562 2335 1566
rect 2339 1562 2583 1566
rect 2587 1562 2599 1566
rect 2603 1562 2743 1566
rect 2747 1562 2839 1566
rect 2843 1562 2903 1566
rect 2907 1562 3047 1566
rect 3051 1562 3063 1566
rect 3067 1562 3223 1566
rect 3227 1562 3231 1566
rect 3235 1562 3383 1566
rect 3387 1562 3399 1566
rect 3403 1562 3543 1566
rect 3547 1562 3551 1566
rect 3555 1562 3695 1566
rect 3699 1562 3703 1566
rect 3707 1562 3839 1566
rect 3843 1562 3943 1566
rect 3947 1562 3967 1566
rect 2025 1561 3967 1562
rect 3973 1561 3974 1567
rect 84 1545 85 1551
rect 91 1550 2019 1551
rect 91 1546 111 1550
rect 115 1546 135 1550
rect 139 1546 287 1550
rect 291 1546 295 1550
rect 299 1546 471 1550
rect 475 1546 487 1550
rect 491 1546 655 1550
rect 659 1546 687 1550
rect 691 1546 839 1550
rect 843 1546 887 1550
rect 891 1546 1015 1550
rect 1019 1546 1079 1550
rect 1083 1546 1183 1550
rect 1187 1546 1263 1550
rect 1267 1546 1343 1550
rect 1347 1546 1447 1550
rect 1451 1546 1495 1550
rect 1499 1546 1623 1550
rect 1627 1546 1639 1550
rect 1643 1546 1783 1550
rect 1787 1546 1807 1550
rect 1811 1546 1903 1550
rect 1907 1546 2007 1550
rect 2011 1546 2019 1550
rect 91 1545 2019 1546
rect 2025 1545 2026 1551
rect 2030 1485 2031 1491
rect 2037 1490 3979 1491
rect 2037 1486 2047 1490
rect 2051 1486 2415 1490
rect 2419 1486 2511 1490
rect 2515 1486 2583 1490
rect 2587 1486 2607 1490
rect 2611 1486 2703 1490
rect 2707 1486 2743 1490
rect 2747 1486 2799 1490
rect 2803 1486 2903 1490
rect 2907 1486 2919 1490
rect 2923 1486 3063 1490
rect 3067 1486 3223 1490
rect 3227 1486 3231 1490
rect 3235 1486 3383 1490
rect 3387 1486 3415 1490
rect 3419 1486 3543 1490
rect 3547 1486 3615 1490
rect 3619 1486 3703 1490
rect 3707 1486 3815 1490
rect 3819 1486 3943 1490
rect 3947 1486 3979 1490
rect 2037 1485 3979 1486
rect 3985 1485 3986 1491
rect 96 1469 97 1475
rect 103 1474 2031 1475
rect 103 1470 111 1474
rect 115 1470 135 1474
rect 139 1470 175 1474
rect 179 1470 295 1474
rect 299 1470 359 1474
rect 363 1470 487 1474
rect 491 1470 567 1474
rect 571 1470 687 1474
rect 691 1470 783 1474
rect 787 1470 887 1474
rect 891 1470 1007 1474
rect 1011 1470 1079 1474
rect 1083 1470 1231 1474
rect 1235 1470 1263 1474
rect 1267 1470 1447 1474
rect 1451 1470 1463 1474
rect 1467 1470 1623 1474
rect 1627 1470 1695 1474
rect 1699 1470 1807 1474
rect 1811 1470 1903 1474
rect 1907 1470 2007 1474
rect 2011 1470 2031 1474
rect 103 1469 2031 1470
rect 2037 1469 2038 1475
rect 84 1393 85 1399
rect 91 1398 2019 1399
rect 91 1394 111 1398
rect 115 1394 175 1398
rect 179 1394 327 1398
rect 331 1394 359 1398
rect 363 1394 463 1398
rect 467 1394 567 1398
rect 571 1394 599 1398
rect 603 1394 727 1398
rect 731 1394 783 1398
rect 787 1394 855 1398
rect 859 1394 983 1398
rect 987 1394 1007 1398
rect 1011 1394 1119 1398
rect 1123 1394 1231 1398
rect 1235 1394 1263 1398
rect 1267 1394 1423 1398
rect 1427 1394 1463 1398
rect 1467 1394 1583 1398
rect 1587 1394 1695 1398
rect 1699 1394 1751 1398
rect 1755 1394 1903 1398
rect 1907 1394 2007 1398
rect 2011 1394 2019 1398
rect 91 1393 2019 1394
rect 2025 1395 2026 1399
rect 2025 1394 3974 1395
rect 2025 1393 2047 1394
rect 2018 1390 2047 1393
rect 2051 1390 2071 1394
rect 2075 1390 2303 1394
rect 2307 1390 2415 1394
rect 2419 1390 2511 1394
rect 2515 1390 2559 1394
rect 2563 1390 2607 1394
rect 2611 1390 2703 1394
rect 2707 1390 2799 1394
rect 2803 1390 2807 1394
rect 2811 1390 2919 1394
rect 2923 1390 3055 1394
rect 3059 1390 3063 1394
rect 3067 1390 3231 1394
rect 3235 1390 3303 1394
rect 3307 1390 3415 1394
rect 3419 1390 3559 1394
rect 3563 1390 3615 1394
rect 3619 1390 3815 1394
rect 3819 1390 3943 1394
rect 3947 1390 3974 1394
rect 2018 1389 3974 1390
rect 518 1388 524 1389
rect 962 1388 968 1389
rect 518 1384 519 1388
rect 523 1384 963 1388
rect 967 1384 968 1388
rect 518 1383 524 1384
rect 962 1383 968 1384
rect 96 1309 97 1315
rect 103 1314 2031 1315
rect 103 1310 111 1314
rect 115 1310 327 1314
rect 331 1310 463 1314
rect 467 1310 551 1314
rect 555 1310 599 1314
rect 603 1310 655 1314
rect 659 1310 727 1314
rect 731 1310 767 1314
rect 771 1310 855 1314
rect 859 1310 879 1314
rect 883 1310 983 1314
rect 987 1310 991 1314
rect 995 1310 1103 1314
rect 1107 1310 1119 1314
rect 1123 1310 1215 1314
rect 1219 1310 1263 1314
rect 1267 1310 1327 1314
rect 1331 1310 1423 1314
rect 1427 1310 1439 1314
rect 1443 1310 1559 1314
rect 1563 1310 1583 1314
rect 1587 1310 1751 1314
rect 1755 1310 1903 1314
rect 1907 1310 2007 1314
rect 2011 1310 2031 1314
rect 103 1309 2031 1310
rect 2037 1311 2038 1315
rect 2037 1310 3986 1311
rect 2037 1309 2047 1310
rect 2030 1306 2047 1309
rect 2051 1306 2071 1310
rect 2075 1306 2223 1310
rect 2227 1306 2303 1310
rect 2307 1306 2415 1310
rect 2419 1306 2559 1310
rect 2563 1306 2615 1310
rect 2619 1306 2807 1310
rect 2811 1306 2815 1310
rect 2819 1306 2999 1310
rect 3003 1306 3055 1310
rect 3059 1306 3175 1310
rect 3179 1306 3303 1310
rect 3307 1306 3343 1310
rect 3347 1306 3503 1310
rect 3507 1306 3559 1310
rect 3563 1306 3663 1310
rect 3667 1306 3815 1310
rect 3819 1306 3831 1310
rect 3835 1306 3943 1310
rect 3947 1306 3986 1310
rect 2030 1305 3986 1306
rect 84 1233 85 1239
rect 91 1238 2019 1239
rect 91 1234 111 1238
rect 115 1234 391 1238
rect 395 1234 519 1238
rect 523 1234 551 1238
rect 555 1234 655 1238
rect 659 1234 663 1238
rect 667 1234 767 1238
rect 771 1234 807 1238
rect 811 1234 879 1238
rect 883 1234 959 1238
rect 963 1234 991 1238
rect 995 1234 1103 1238
rect 1107 1234 1111 1238
rect 1115 1234 1215 1238
rect 1219 1234 1255 1238
rect 1259 1234 1327 1238
rect 1331 1234 1407 1238
rect 1411 1234 1439 1238
rect 1443 1234 1559 1238
rect 1563 1234 1711 1238
rect 1715 1234 2007 1238
rect 2011 1234 2019 1238
rect 91 1233 2019 1234
rect 2025 1233 2026 1239
rect 2018 1221 2019 1227
rect 2025 1226 3967 1227
rect 2025 1222 2047 1226
rect 2051 1222 2071 1226
rect 2075 1222 2135 1226
rect 2139 1222 2223 1226
rect 2227 1222 2311 1226
rect 2315 1222 2415 1226
rect 2419 1222 2503 1226
rect 2507 1222 2615 1226
rect 2619 1222 2695 1226
rect 2699 1222 2815 1226
rect 2819 1222 2887 1226
rect 2891 1222 2999 1226
rect 3003 1222 3071 1226
rect 3075 1222 3175 1226
rect 3179 1222 3239 1226
rect 3243 1222 3343 1226
rect 3347 1222 3399 1226
rect 3403 1222 3503 1226
rect 3507 1222 3551 1226
rect 3555 1222 3663 1226
rect 3667 1222 3703 1226
rect 3707 1222 3831 1226
rect 3835 1222 3839 1226
rect 3843 1222 3943 1226
rect 3947 1222 3967 1226
rect 2025 1221 3967 1222
rect 3973 1221 3974 1227
rect 96 1153 97 1159
rect 103 1158 2031 1159
rect 103 1154 111 1158
rect 115 1154 175 1158
rect 179 1154 327 1158
rect 331 1154 391 1158
rect 395 1154 495 1158
rect 499 1154 519 1158
rect 523 1154 663 1158
rect 667 1154 671 1158
rect 675 1154 807 1158
rect 811 1154 847 1158
rect 851 1154 959 1158
rect 963 1154 1031 1158
rect 1035 1154 1111 1158
rect 1115 1154 1207 1158
rect 1211 1154 1255 1158
rect 1259 1154 1383 1158
rect 1387 1154 1407 1158
rect 1411 1154 1559 1158
rect 1563 1154 1567 1158
rect 1571 1154 1711 1158
rect 1715 1154 1751 1158
rect 1755 1154 2007 1158
rect 2011 1154 2031 1158
rect 103 1153 2031 1154
rect 2037 1153 2038 1159
rect 2030 1137 2031 1143
rect 2037 1142 3979 1143
rect 2037 1138 2047 1142
rect 2051 1138 2135 1142
rect 2139 1138 2295 1142
rect 2299 1138 2311 1142
rect 2315 1138 2423 1142
rect 2427 1138 2503 1142
rect 2507 1138 2559 1142
rect 2563 1138 2695 1142
rect 2699 1138 2839 1142
rect 2843 1138 2887 1142
rect 2891 1138 2991 1142
rect 2995 1138 3071 1142
rect 3075 1138 3151 1142
rect 3155 1138 3239 1142
rect 3243 1138 3319 1142
rect 3323 1138 3399 1142
rect 3403 1138 3495 1142
rect 3499 1138 3551 1142
rect 3555 1138 3679 1142
rect 3683 1138 3703 1142
rect 3707 1138 3839 1142
rect 3843 1138 3943 1142
rect 3947 1138 3979 1142
rect 2037 1137 3979 1138
rect 3985 1137 3986 1143
rect 84 1069 85 1075
rect 91 1074 2019 1075
rect 91 1070 111 1074
rect 115 1070 135 1074
rect 139 1070 175 1074
rect 179 1070 231 1074
rect 235 1070 327 1074
rect 331 1070 375 1074
rect 379 1070 495 1074
rect 499 1070 543 1074
rect 547 1070 671 1074
rect 675 1070 727 1074
rect 731 1070 847 1074
rect 851 1070 911 1074
rect 915 1070 1031 1074
rect 1035 1070 1095 1074
rect 1099 1070 1207 1074
rect 1211 1070 1279 1074
rect 1283 1070 1383 1074
rect 1387 1070 1463 1074
rect 1467 1070 1567 1074
rect 1571 1070 1647 1074
rect 1651 1070 1751 1074
rect 1755 1070 1831 1074
rect 1835 1070 2007 1074
rect 2011 1070 2019 1074
rect 91 1069 2019 1070
rect 2025 1069 2026 1075
rect 242 1060 248 1061
rect 858 1060 864 1061
rect 242 1056 243 1060
rect 247 1056 859 1060
rect 863 1056 864 1060
rect 2018 1057 2019 1063
rect 2025 1062 3967 1063
rect 2025 1058 2047 1062
rect 2051 1058 2295 1062
rect 2299 1058 2423 1062
rect 2427 1058 2495 1062
rect 2499 1058 2559 1062
rect 2563 1058 2599 1062
rect 2603 1058 2695 1062
rect 2699 1058 2711 1062
rect 2715 1058 2839 1062
rect 2843 1058 2847 1062
rect 2851 1058 2991 1062
rect 2995 1058 3007 1062
rect 3011 1058 3151 1062
rect 3155 1058 3199 1062
rect 3203 1058 3319 1062
rect 3323 1058 3407 1062
rect 3411 1058 3495 1062
rect 3499 1058 3631 1062
rect 3635 1058 3679 1062
rect 3683 1058 3839 1062
rect 3843 1058 3943 1062
rect 3947 1058 3967 1062
rect 2025 1057 3967 1058
rect 3973 1057 3974 1063
rect 242 1055 248 1056
rect 858 1055 864 1056
rect 3190 1028 3196 1029
rect 3558 1028 3564 1029
rect 3190 1024 3191 1028
rect 3195 1024 3559 1028
rect 3563 1024 3564 1028
rect 3190 1023 3196 1024
rect 3558 1023 3564 1024
rect 96 993 97 999
rect 103 998 2031 999
rect 103 994 111 998
rect 115 994 135 998
rect 139 994 231 998
rect 235 994 271 998
rect 275 994 375 998
rect 379 994 447 998
rect 451 994 543 998
rect 547 994 631 998
rect 635 994 727 998
rect 731 994 823 998
rect 827 994 911 998
rect 915 994 1007 998
rect 1011 994 1095 998
rect 1099 994 1175 998
rect 1179 994 1279 998
rect 1283 994 1335 998
rect 1339 994 1463 998
rect 1467 994 1487 998
rect 1491 994 1631 998
rect 1635 994 1647 998
rect 1651 994 1775 998
rect 1779 994 1831 998
rect 1835 994 1903 998
rect 1907 994 2007 998
rect 2011 994 2031 998
rect 103 993 2031 994
rect 2037 993 2038 999
rect 2030 981 2031 987
rect 2037 986 3979 987
rect 2037 982 2047 986
rect 2051 982 2495 986
rect 2499 982 2599 986
rect 2603 982 2647 986
rect 2651 982 2711 986
rect 2715 982 2743 986
rect 2747 982 2847 986
rect 2851 982 2967 986
rect 2971 982 3007 986
rect 3011 982 3111 986
rect 3115 982 3199 986
rect 3203 982 3279 986
rect 3283 982 3407 986
rect 3411 982 3463 986
rect 3467 982 3631 986
rect 3635 982 3663 986
rect 3667 982 3839 986
rect 3843 982 3943 986
rect 3947 982 3979 986
rect 2037 981 3979 982
rect 3985 981 3986 987
rect 84 917 85 923
rect 91 922 2019 923
rect 91 918 111 922
rect 115 918 135 922
rect 139 918 271 922
rect 275 918 447 922
rect 451 918 455 922
rect 459 918 631 922
rect 635 918 655 922
rect 659 918 823 922
rect 827 918 855 922
rect 859 918 1007 922
rect 1011 918 1055 922
rect 1059 918 1175 922
rect 1179 918 1239 922
rect 1243 918 1335 922
rect 1339 918 1415 922
rect 1419 918 1487 922
rect 1491 918 1583 922
rect 1587 918 1631 922
rect 1635 918 1751 922
rect 1755 918 1775 922
rect 1779 918 1903 922
rect 1907 918 2007 922
rect 2011 918 2019 922
rect 91 917 2019 918
rect 2025 917 2026 923
rect 2018 893 2019 899
rect 2025 898 3967 899
rect 2025 894 2047 898
rect 2051 894 2071 898
rect 2075 894 2255 898
rect 2259 894 2463 898
rect 2467 894 2647 898
rect 2651 894 2679 898
rect 2683 894 2743 898
rect 2747 894 2847 898
rect 2851 894 2895 898
rect 2899 894 2967 898
rect 2971 894 3111 898
rect 3115 894 3127 898
rect 3131 894 3279 898
rect 3283 894 3367 898
rect 3371 894 3463 898
rect 3467 894 3615 898
rect 3619 894 3663 898
rect 3667 894 3839 898
rect 3843 894 3943 898
rect 3947 894 3967 898
rect 2025 893 3967 894
rect 3973 893 3974 899
rect 96 841 97 847
rect 103 846 2031 847
rect 103 842 111 846
rect 115 842 135 846
rect 139 842 215 846
rect 219 842 271 846
rect 275 842 343 846
rect 347 842 455 846
rect 459 842 495 846
rect 499 842 655 846
rect 659 842 831 846
rect 835 842 855 846
rect 859 842 1007 846
rect 1011 842 1055 846
rect 1059 842 1183 846
rect 1187 842 1239 846
rect 1243 842 1359 846
rect 1363 842 1415 846
rect 1419 842 1535 846
rect 1539 842 1583 846
rect 1587 842 1719 846
rect 1723 842 1751 846
rect 1755 842 1903 846
rect 1907 842 2007 846
rect 2011 842 2031 846
rect 103 841 2031 842
rect 2037 841 2038 847
rect 2030 817 2031 823
rect 2037 822 3979 823
rect 2037 818 2047 822
rect 2051 818 2071 822
rect 2075 818 2215 822
rect 2219 818 2255 822
rect 2259 818 2327 822
rect 2331 818 2447 822
rect 2451 818 2463 822
rect 2467 818 2583 822
rect 2587 818 2679 822
rect 2683 818 2735 822
rect 2739 818 2895 822
rect 2899 818 3063 822
rect 3067 818 3127 822
rect 3131 818 3247 822
rect 3251 818 3367 822
rect 3371 818 3447 822
rect 3451 818 3615 822
rect 3619 818 3655 822
rect 3659 818 3839 822
rect 3843 818 3943 822
rect 3947 818 3979 822
rect 2037 817 3979 818
rect 3985 817 3986 823
rect 84 765 85 771
rect 91 770 2019 771
rect 91 766 111 770
rect 115 766 215 770
rect 219 766 343 770
rect 347 766 375 770
rect 379 766 495 770
rect 499 766 623 770
rect 627 766 655 770
rect 659 766 751 770
rect 755 766 831 770
rect 835 766 887 770
rect 891 766 1007 770
rect 1011 766 1023 770
rect 1027 766 1167 770
rect 1171 766 1183 770
rect 1187 766 1311 770
rect 1315 766 1359 770
rect 1363 766 1455 770
rect 1459 766 1535 770
rect 1539 766 1599 770
rect 1603 766 1719 770
rect 1723 766 2007 770
rect 2011 766 2019 770
rect 91 765 2019 766
rect 2025 765 2026 771
rect 2018 737 2019 743
rect 2025 742 3967 743
rect 2025 738 2047 742
rect 2051 738 2215 742
rect 2219 738 2327 742
rect 2331 738 2375 742
rect 2379 738 2447 742
rect 2451 738 2495 742
rect 2499 738 2583 742
rect 2587 738 2623 742
rect 2627 738 2735 742
rect 2739 738 2767 742
rect 2771 738 2895 742
rect 2899 738 2911 742
rect 2915 738 3063 742
rect 3067 738 3215 742
rect 3219 738 3247 742
rect 3251 738 3367 742
rect 3371 738 3447 742
rect 3451 738 3519 742
rect 3523 738 3655 742
rect 3659 738 3679 742
rect 3683 738 3839 742
rect 3843 738 3943 742
rect 3947 738 3967 742
rect 2025 737 3967 738
rect 3973 737 3974 743
rect 96 689 97 695
rect 103 694 2031 695
rect 103 690 111 694
rect 115 690 375 694
rect 379 690 495 694
rect 499 690 527 694
rect 531 690 623 694
rect 627 690 631 694
rect 635 690 743 694
rect 747 690 751 694
rect 755 690 855 694
rect 859 690 887 694
rect 891 690 967 694
rect 971 690 1023 694
rect 1027 690 1071 694
rect 1075 690 1167 694
rect 1171 690 1183 694
rect 1187 690 1295 694
rect 1299 690 1311 694
rect 1315 690 1407 694
rect 1411 690 1455 694
rect 1459 690 1519 694
rect 1523 690 1599 694
rect 1603 690 2007 694
rect 2011 690 2031 694
rect 103 689 2031 690
rect 2037 689 2038 695
rect 2030 653 2031 659
rect 2037 658 3979 659
rect 2037 654 2047 658
rect 2051 654 2111 658
rect 2115 654 2247 658
rect 2251 654 2375 658
rect 2379 654 2399 658
rect 2403 654 2495 658
rect 2499 654 2575 658
rect 2579 654 2623 658
rect 2627 654 2759 658
rect 2763 654 2767 658
rect 2771 654 2911 658
rect 2915 654 2943 658
rect 2947 654 3063 658
rect 3067 654 3127 658
rect 3131 654 3215 658
rect 3219 654 3303 658
rect 3307 654 3367 658
rect 3371 654 3479 658
rect 3483 654 3519 658
rect 3523 654 3655 658
rect 3659 654 3679 658
rect 3683 654 3831 658
rect 3835 654 3839 658
rect 3843 654 3943 658
rect 3947 654 3979 658
rect 2037 653 3979 654
rect 3985 653 3986 659
rect 84 613 85 619
rect 91 618 2019 619
rect 91 614 111 618
rect 115 614 527 618
rect 531 614 631 618
rect 635 614 687 618
rect 691 614 743 618
rect 747 614 783 618
rect 787 614 855 618
rect 859 614 879 618
rect 883 614 967 618
rect 971 614 975 618
rect 979 614 1071 618
rect 1075 614 1167 618
rect 1171 614 1183 618
rect 1187 614 1263 618
rect 1267 614 1295 618
rect 1299 614 1359 618
rect 1363 614 1407 618
rect 1411 614 1455 618
rect 1459 614 1519 618
rect 1523 614 2007 618
rect 2011 614 2019 618
rect 91 613 2019 614
rect 2025 613 2026 619
rect 2018 573 2019 579
rect 2025 578 3967 579
rect 2025 574 2047 578
rect 2051 574 2071 578
rect 2075 574 2111 578
rect 2115 574 2183 578
rect 2187 574 2247 578
rect 2251 574 2335 578
rect 2339 574 2399 578
rect 2403 574 2503 578
rect 2507 574 2575 578
rect 2579 574 2687 578
rect 2691 574 2759 578
rect 2763 574 2879 578
rect 2883 574 2943 578
rect 2947 574 3071 578
rect 3075 574 3127 578
rect 3131 574 3263 578
rect 3267 574 3303 578
rect 3307 574 3455 578
rect 3459 574 3479 578
rect 3483 574 3647 578
rect 3651 574 3655 578
rect 3659 574 3831 578
rect 3835 574 3839 578
rect 3843 574 3943 578
rect 3947 574 3967 578
rect 2025 573 3967 574
rect 3973 573 3974 579
rect 96 517 97 523
rect 103 522 2031 523
rect 103 518 111 522
rect 115 518 383 522
rect 387 518 479 522
rect 483 518 575 522
rect 579 518 671 522
rect 675 518 687 522
rect 691 518 767 522
rect 771 518 783 522
rect 787 518 863 522
rect 867 518 879 522
rect 883 518 959 522
rect 963 518 975 522
rect 979 518 1055 522
rect 1059 518 1071 522
rect 1075 518 1151 522
rect 1155 518 1167 522
rect 1171 518 1247 522
rect 1251 518 1263 522
rect 1267 518 1343 522
rect 1347 518 1359 522
rect 1363 518 1439 522
rect 1443 518 1455 522
rect 1459 518 1535 522
rect 1539 518 2007 522
rect 2011 518 2031 522
rect 103 517 2031 518
rect 2037 517 2038 523
rect 2030 497 2031 503
rect 2037 502 3979 503
rect 2037 498 2047 502
rect 2051 498 2071 502
rect 2075 498 2183 502
rect 2187 498 2319 502
rect 2323 498 2335 502
rect 2339 498 2463 502
rect 2467 498 2503 502
rect 2507 498 2615 502
rect 2619 498 2687 502
rect 2691 498 2775 502
rect 2779 498 2879 502
rect 2883 498 2959 502
rect 2963 498 3071 502
rect 3075 498 3159 502
rect 3163 498 3263 502
rect 3267 498 3367 502
rect 3371 498 3455 502
rect 3459 498 3583 502
rect 3587 498 3647 502
rect 3651 498 3807 502
rect 3811 498 3839 502
rect 3843 498 3943 502
rect 3947 498 3979 502
rect 2037 497 3979 498
rect 3985 497 3986 503
rect 84 429 85 435
rect 91 434 2019 435
rect 91 430 111 434
rect 115 430 383 434
rect 387 430 479 434
rect 483 430 487 434
rect 491 430 575 434
rect 579 430 583 434
rect 587 430 671 434
rect 675 430 687 434
rect 691 430 767 434
rect 771 430 791 434
rect 795 430 863 434
rect 867 430 895 434
rect 899 430 959 434
rect 963 430 999 434
rect 1003 430 1055 434
rect 1059 430 1103 434
rect 1107 430 1151 434
rect 1155 430 1207 434
rect 1211 430 1247 434
rect 1251 430 1319 434
rect 1323 430 1343 434
rect 1347 430 1431 434
rect 1435 430 1439 434
rect 1443 430 1535 434
rect 1539 430 2007 434
rect 2011 430 2019 434
rect 91 429 2019 430
rect 2025 429 2026 435
rect 2018 427 2026 429
rect 2018 421 2019 427
rect 2025 426 3967 427
rect 2025 422 2047 426
rect 2051 422 2183 426
rect 2187 422 2319 426
rect 2323 422 2343 426
rect 2347 422 2463 426
rect 2467 422 2487 426
rect 2491 422 2615 426
rect 2619 422 2639 426
rect 2643 422 2775 426
rect 2779 422 2799 426
rect 2803 422 2959 426
rect 2963 422 3111 426
rect 3115 422 3159 426
rect 3163 422 3263 426
rect 3267 422 3367 426
rect 3371 422 3415 426
rect 3419 422 3559 426
rect 3563 422 3583 426
rect 3587 422 3711 426
rect 3715 422 3807 426
rect 3811 422 3839 426
rect 3843 422 3943 426
rect 3947 422 3967 426
rect 2025 421 3967 422
rect 3973 421 3974 427
rect 538 420 544 421
rect 858 420 864 421
rect 538 416 539 420
rect 543 416 859 420
rect 863 416 864 420
rect 538 415 544 416
rect 858 415 864 416
rect 96 349 97 355
rect 103 354 2031 355
rect 103 350 111 354
rect 115 350 327 354
rect 331 350 463 354
rect 467 350 487 354
rect 491 350 583 354
rect 587 350 615 354
rect 619 350 687 354
rect 691 350 767 354
rect 771 350 791 354
rect 795 350 895 354
rect 899 350 919 354
rect 923 350 999 354
rect 1003 350 1063 354
rect 1067 350 1103 354
rect 1107 350 1207 354
rect 1211 350 1319 354
rect 1323 350 1351 354
rect 1355 350 1431 354
rect 1435 350 1495 354
rect 1499 350 1639 354
rect 1643 350 2007 354
rect 2011 350 2031 354
rect 103 349 2031 350
rect 2037 349 2038 355
rect 2030 347 2038 349
rect 2030 341 2031 347
rect 2037 346 3979 347
rect 2037 342 2047 346
rect 2051 342 2343 346
rect 2347 342 2487 346
rect 2491 342 2495 346
rect 2499 342 2639 346
rect 2643 342 2799 346
rect 2803 342 2959 346
rect 2963 342 3111 346
rect 3115 342 3119 346
rect 3123 342 3263 346
rect 3267 342 3271 346
rect 3275 342 3415 346
rect 3419 342 3423 346
rect 3427 342 3559 346
rect 3563 342 3567 346
rect 3571 342 3711 346
rect 3715 342 3839 346
rect 3843 342 3943 346
rect 3947 342 3979 346
rect 2037 341 3979 342
rect 3985 341 3986 347
rect 2550 284 2556 285
rect 2898 284 2904 285
rect 2550 280 2551 284
rect 2555 280 2899 284
rect 2903 280 2904 284
rect 2550 279 2556 280
rect 2898 279 2904 280
rect 84 265 85 271
rect 91 270 2019 271
rect 91 266 111 270
rect 115 266 167 270
rect 171 266 327 270
rect 331 266 463 270
rect 467 266 503 270
rect 507 266 615 270
rect 619 266 687 270
rect 691 266 767 270
rect 771 266 871 270
rect 875 266 919 270
rect 923 266 1047 270
rect 1051 266 1063 270
rect 1067 266 1207 270
rect 1211 266 1215 270
rect 1219 266 1351 270
rect 1355 266 1367 270
rect 1371 266 1495 270
rect 1499 266 1511 270
rect 1515 266 1639 270
rect 1643 266 1647 270
rect 1651 266 1783 270
rect 1787 266 1903 270
rect 1907 266 2007 270
rect 2011 266 2019 270
rect 91 265 2019 266
rect 2025 270 3974 271
rect 2025 266 2047 270
rect 2051 266 2071 270
rect 2075 266 2271 270
rect 2275 266 2495 270
rect 2499 266 2639 270
rect 2643 266 2703 270
rect 2707 266 2799 270
rect 2803 266 2903 270
rect 2907 266 2959 270
rect 2963 266 3095 270
rect 3099 266 3119 270
rect 3123 266 3271 270
rect 3275 266 3287 270
rect 3291 266 3423 270
rect 3427 266 3479 270
rect 3483 266 3567 270
rect 3571 266 3671 270
rect 3675 266 3711 270
rect 3715 266 3839 270
rect 3843 266 3943 270
rect 3947 266 3974 270
rect 2025 265 3974 266
rect 2030 170 3986 171
rect 2030 167 2047 170
rect 96 161 97 167
rect 103 166 2031 167
rect 103 162 111 166
rect 115 162 135 166
rect 139 162 167 166
rect 171 162 231 166
rect 235 162 327 166
rect 331 162 423 166
rect 427 162 503 166
rect 507 162 527 166
rect 531 162 647 166
rect 651 162 687 166
rect 691 162 775 166
rect 779 162 871 166
rect 875 162 903 166
rect 907 162 1031 166
rect 1035 162 1047 166
rect 1051 162 1151 166
rect 1155 162 1215 166
rect 1219 162 1271 166
rect 1275 162 1367 166
rect 1371 162 1383 166
rect 1387 162 1487 166
rect 1491 162 1511 166
rect 1515 162 1591 166
rect 1595 162 1647 166
rect 1651 162 1703 166
rect 1707 162 1783 166
rect 1787 162 1807 166
rect 1811 162 1903 166
rect 1907 162 2007 166
rect 2011 162 2031 166
rect 103 161 2031 162
rect 2037 166 2047 167
rect 2051 166 2071 170
rect 2075 166 2167 170
rect 2171 166 2263 170
rect 2267 166 2271 170
rect 2275 166 2359 170
rect 2363 166 2455 170
rect 2459 166 2495 170
rect 2499 166 2551 170
rect 2555 166 2655 170
rect 2659 166 2703 170
rect 2707 166 2759 170
rect 2763 166 2863 170
rect 2867 166 2903 170
rect 2907 166 2975 170
rect 2979 166 3095 170
rect 3099 166 3103 170
rect 3107 166 3239 170
rect 3243 166 3287 170
rect 3291 166 3383 170
rect 3387 166 3479 170
rect 3483 166 3535 170
rect 3539 166 3671 170
rect 3675 166 3695 170
rect 3699 166 3839 170
rect 3843 166 3943 170
rect 3947 166 3986 170
rect 2037 165 3986 166
rect 2037 161 2038 165
rect 2018 94 3974 95
rect 2018 91 2047 94
rect 84 85 85 91
rect 91 90 2019 91
rect 91 86 111 90
rect 115 86 135 90
rect 139 86 231 90
rect 235 86 327 90
rect 331 86 423 90
rect 427 86 527 90
rect 531 86 647 90
rect 651 86 775 90
rect 779 86 903 90
rect 907 86 1031 90
rect 1035 86 1151 90
rect 1155 86 1271 90
rect 1275 86 1383 90
rect 1387 86 1487 90
rect 1491 86 1591 90
rect 1595 86 1703 90
rect 1707 86 1807 90
rect 1811 86 1903 90
rect 1907 86 2007 90
rect 2011 86 2019 90
rect 91 85 2019 86
rect 2025 90 2047 91
rect 2051 90 2071 94
rect 2075 90 2167 94
rect 2171 90 2263 94
rect 2267 90 2359 94
rect 2363 90 2455 94
rect 2459 90 2551 94
rect 2555 90 2655 94
rect 2659 90 2759 94
rect 2763 90 2863 94
rect 2867 90 2975 94
rect 2979 90 3103 94
rect 3107 90 3239 94
rect 3243 90 3383 94
rect 3387 90 3535 94
rect 3539 90 3695 94
rect 3699 90 3839 94
rect 3843 90 3943 94
rect 3947 90 3974 94
rect 2025 89 3974 90
rect 2025 85 2026 89
<< m5c >>
rect 97 4025 103 4031
rect 2031 4025 2037 4031
rect 2019 4013 2025 4019
rect 3967 4013 3973 4019
rect 85 3949 91 3955
rect 2019 3949 2025 3955
rect 2031 3937 2037 3943
rect 3979 3937 3985 3943
rect 97 3873 103 3879
rect 2031 3873 2037 3879
rect 2019 3853 2025 3859
rect 3967 3853 3973 3859
rect 85 3793 91 3799
rect 2019 3793 2025 3799
rect 2031 3777 2037 3783
rect 3979 3777 3985 3783
rect 97 3709 103 3715
rect 2031 3709 2037 3715
rect 2019 3697 2025 3703
rect 3967 3697 3973 3703
rect 85 3625 91 3631
rect 2019 3625 2025 3631
rect 2031 3613 2037 3619
rect 3979 3613 3985 3619
rect 2019 3547 2025 3553
rect 97 3537 103 3543
rect 2031 3537 2037 3543
rect 3967 3537 3973 3543
rect 85 3453 91 3459
rect 2019 3453 2025 3459
rect 2031 3457 2037 3463
rect 3979 3457 3985 3463
rect 97 3377 103 3383
rect 2031 3377 2037 3383
rect 2019 3365 2025 3371
rect 3967 3365 3973 3371
rect 85 3301 91 3307
rect 2019 3301 2025 3307
rect 2031 3281 2037 3287
rect 3979 3281 3985 3287
rect 97 3225 103 3231
rect 2031 3225 2037 3231
rect 2019 3205 2025 3211
rect 3967 3205 3973 3211
rect 85 3145 91 3151
rect 2019 3145 2025 3151
rect 2031 3117 2037 3123
rect 3979 3117 3985 3123
rect 97 3061 103 3067
rect 2031 3061 2037 3067
rect 2019 3041 2025 3047
rect 3967 3041 3973 3047
rect 85 2981 91 2987
rect 2019 2981 2025 2987
rect 2031 2961 2037 2967
rect 3979 2961 3985 2967
rect 97 2897 103 2903
rect 2031 2897 2037 2903
rect 2019 2885 2025 2891
rect 3967 2885 3973 2891
rect 85 2817 91 2823
rect 2019 2817 2025 2823
rect 2031 2805 2037 2811
rect 3979 2805 3985 2811
rect 97 2737 103 2743
rect 2031 2737 2037 2743
rect 2019 2725 2025 2731
rect 3967 2725 3973 2731
rect 85 2657 91 2663
rect 2019 2657 2025 2663
rect 2031 2641 2037 2647
rect 3979 2641 3985 2647
rect 97 2581 103 2587
rect 2031 2581 2037 2587
rect 2019 2561 2025 2567
rect 3967 2561 3973 2567
rect 85 2489 91 2495
rect 2019 2489 2025 2495
rect 2031 2481 2037 2487
rect 3979 2481 3985 2487
rect 2019 2407 2025 2413
rect 97 2397 103 2403
rect 2031 2397 2037 2403
rect 3967 2393 3973 2399
rect 85 2321 91 2327
rect 2019 2321 2025 2327
rect 2031 2301 2037 2307
rect 3979 2301 3985 2307
rect 97 2241 103 2247
rect 2031 2241 2037 2247
rect 2019 2225 2025 2231
rect 3967 2225 3973 2231
rect 85 2165 91 2171
rect 2019 2165 2025 2171
rect 2031 2129 2037 2135
rect 3979 2129 3985 2135
rect 97 2089 103 2095
rect 2031 2089 2037 2095
rect 2019 2045 2025 2051
rect 3967 2045 3973 2051
rect 85 2009 91 2015
rect 2019 2009 2025 2015
rect 2031 1965 2037 1971
rect 3979 1965 3985 1971
rect 97 1933 103 1939
rect 2031 1933 2037 1939
rect 2019 1877 2025 1883
rect 3967 1877 3973 1883
rect 85 1857 91 1863
rect 2019 1857 2025 1863
rect 2031 1797 2037 1803
rect 3979 1797 3985 1803
rect 97 1777 103 1783
rect 2031 1777 2037 1783
rect 2019 1717 2025 1723
rect 3967 1717 3973 1723
rect 85 1701 91 1707
rect 2019 1701 2025 1707
rect 2031 1641 2037 1647
rect 3979 1641 3985 1647
rect 97 1625 103 1631
rect 2031 1625 2037 1631
rect 2019 1561 2025 1567
rect 3967 1561 3973 1567
rect 85 1545 91 1551
rect 2019 1545 2025 1551
rect 2031 1485 2037 1491
rect 3979 1485 3985 1491
rect 97 1469 103 1475
rect 2031 1469 2037 1475
rect 85 1393 91 1399
rect 2019 1393 2025 1399
rect 97 1309 103 1315
rect 2031 1309 2037 1315
rect 85 1233 91 1239
rect 2019 1233 2025 1239
rect 2019 1221 2025 1227
rect 3967 1221 3973 1227
rect 97 1153 103 1159
rect 2031 1153 2037 1159
rect 2031 1137 2037 1143
rect 3979 1137 3985 1143
rect 85 1069 91 1075
rect 2019 1069 2025 1075
rect 2019 1057 2025 1063
rect 3967 1057 3973 1063
rect 97 993 103 999
rect 2031 993 2037 999
rect 2031 981 2037 987
rect 3979 981 3985 987
rect 85 917 91 923
rect 2019 917 2025 923
rect 2019 893 2025 899
rect 3967 893 3973 899
rect 97 841 103 847
rect 2031 841 2037 847
rect 2031 817 2037 823
rect 3979 817 3985 823
rect 85 765 91 771
rect 2019 765 2025 771
rect 2019 737 2025 743
rect 3967 737 3973 743
rect 97 689 103 695
rect 2031 689 2037 695
rect 2031 653 2037 659
rect 3979 653 3985 659
rect 85 613 91 619
rect 2019 613 2025 619
rect 2019 573 2025 579
rect 3967 573 3973 579
rect 97 517 103 523
rect 2031 517 2037 523
rect 2031 497 2037 503
rect 3979 497 3985 503
rect 85 429 91 435
rect 2019 429 2025 435
rect 2019 421 2025 427
rect 3967 421 3973 427
rect 97 349 103 355
rect 2031 349 2037 355
rect 2031 341 2037 347
rect 3979 341 3985 347
rect 85 265 91 271
rect 2019 265 2025 271
rect 97 161 103 167
rect 2031 161 2037 167
rect 85 85 91 91
rect 2019 85 2025 91
<< m5 >>
rect 84 3955 92 4032
rect 84 3949 85 3955
rect 91 3949 92 3955
rect 84 3799 92 3949
rect 84 3793 85 3799
rect 91 3793 92 3799
rect 84 3631 92 3793
rect 84 3625 85 3631
rect 91 3625 92 3631
rect 84 3459 92 3625
rect 84 3453 85 3459
rect 91 3453 92 3459
rect 84 3307 92 3453
rect 84 3301 85 3307
rect 91 3301 92 3307
rect 84 3151 92 3301
rect 84 3145 85 3151
rect 91 3145 92 3151
rect 84 2987 92 3145
rect 84 2981 85 2987
rect 91 2981 92 2987
rect 84 2823 92 2981
rect 84 2817 85 2823
rect 91 2817 92 2823
rect 84 2663 92 2817
rect 84 2657 85 2663
rect 91 2657 92 2663
rect 84 2495 92 2657
rect 84 2489 85 2495
rect 91 2489 92 2495
rect 84 2327 92 2489
rect 84 2321 85 2327
rect 91 2321 92 2327
rect 84 2171 92 2321
rect 84 2165 85 2171
rect 91 2165 92 2171
rect 84 2015 92 2165
rect 84 2009 85 2015
rect 91 2009 92 2015
rect 84 1863 92 2009
rect 84 1857 85 1863
rect 91 1857 92 1863
rect 84 1707 92 1857
rect 84 1701 85 1707
rect 91 1701 92 1707
rect 84 1551 92 1701
rect 84 1545 85 1551
rect 91 1545 92 1551
rect 84 1399 92 1545
rect 84 1393 85 1399
rect 91 1393 92 1399
rect 84 1239 92 1393
rect 84 1233 85 1239
rect 91 1233 92 1239
rect 84 1075 92 1233
rect 84 1069 85 1075
rect 91 1069 92 1075
rect 84 923 92 1069
rect 84 917 85 923
rect 91 917 92 923
rect 84 771 92 917
rect 84 765 85 771
rect 91 765 92 771
rect 84 619 92 765
rect 84 613 85 619
rect 91 613 92 619
rect 84 435 92 613
rect 84 429 85 435
rect 91 429 92 435
rect 84 271 92 429
rect 84 265 85 271
rect 91 265 92 271
rect 84 91 92 265
rect 84 85 85 91
rect 91 85 92 91
rect 84 72 92 85
rect 96 4031 104 4032
rect 96 4025 97 4031
rect 103 4025 104 4031
rect 96 3879 104 4025
rect 96 3873 97 3879
rect 103 3873 104 3879
rect 96 3715 104 3873
rect 96 3709 97 3715
rect 103 3709 104 3715
rect 96 3543 104 3709
rect 96 3537 97 3543
rect 103 3537 104 3543
rect 96 3383 104 3537
rect 96 3377 97 3383
rect 103 3377 104 3383
rect 96 3231 104 3377
rect 96 3225 97 3231
rect 103 3225 104 3231
rect 96 3067 104 3225
rect 96 3061 97 3067
rect 103 3061 104 3067
rect 96 2903 104 3061
rect 96 2897 97 2903
rect 103 2897 104 2903
rect 96 2743 104 2897
rect 96 2737 97 2743
rect 103 2737 104 2743
rect 96 2587 104 2737
rect 96 2581 97 2587
rect 103 2581 104 2587
rect 96 2403 104 2581
rect 96 2397 97 2403
rect 103 2397 104 2403
rect 96 2247 104 2397
rect 96 2241 97 2247
rect 103 2241 104 2247
rect 96 2095 104 2241
rect 96 2089 97 2095
rect 103 2089 104 2095
rect 96 1939 104 2089
rect 96 1933 97 1939
rect 103 1933 104 1939
rect 96 1783 104 1933
rect 96 1777 97 1783
rect 103 1777 104 1783
rect 96 1631 104 1777
rect 96 1625 97 1631
rect 103 1625 104 1631
rect 96 1475 104 1625
rect 96 1469 97 1475
rect 103 1469 104 1475
rect 96 1315 104 1469
rect 96 1309 97 1315
rect 103 1309 104 1315
rect 96 1159 104 1309
rect 96 1153 97 1159
rect 103 1153 104 1159
rect 96 999 104 1153
rect 96 993 97 999
rect 103 993 104 999
rect 96 847 104 993
rect 96 841 97 847
rect 103 841 104 847
rect 96 695 104 841
rect 96 689 97 695
rect 103 689 104 695
rect 96 523 104 689
rect 96 517 97 523
rect 103 517 104 523
rect 96 355 104 517
rect 96 349 97 355
rect 103 349 104 355
rect 96 167 104 349
rect 96 161 97 167
rect 103 161 104 167
rect 96 72 104 161
rect 2018 4019 2026 4032
rect 2018 4013 2019 4019
rect 2025 4013 2026 4019
rect 2018 3955 2026 4013
rect 2018 3949 2019 3955
rect 2025 3949 2026 3955
rect 2018 3859 2026 3949
rect 2018 3853 2019 3859
rect 2025 3853 2026 3859
rect 2018 3799 2026 3853
rect 2018 3793 2019 3799
rect 2025 3793 2026 3799
rect 2018 3703 2026 3793
rect 2018 3697 2019 3703
rect 2025 3697 2026 3703
rect 2018 3631 2026 3697
rect 2018 3625 2019 3631
rect 2025 3625 2026 3631
rect 2018 3553 2026 3625
rect 2018 3547 2019 3553
rect 2025 3547 2026 3553
rect 2018 3459 2026 3547
rect 2018 3453 2019 3459
rect 2025 3453 2026 3459
rect 2018 3371 2026 3453
rect 2018 3365 2019 3371
rect 2025 3365 2026 3371
rect 2018 3307 2026 3365
rect 2018 3301 2019 3307
rect 2025 3301 2026 3307
rect 2018 3211 2026 3301
rect 2018 3205 2019 3211
rect 2025 3205 2026 3211
rect 2018 3151 2026 3205
rect 2018 3145 2019 3151
rect 2025 3145 2026 3151
rect 2018 3047 2026 3145
rect 2018 3041 2019 3047
rect 2025 3041 2026 3047
rect 2018 2987 2026 3041
rect 2018 2981 2019 2987
rect 2025 2981 2026 2987
rect 2018 2891 2026 2981
rect 2018 2885 2019 2891
rect 2025 2885 2026 2891
rect 2018 2823 2026 2885
rect 2018 2817 2019 2823
rect 2025 2817 2026 2823
rect 2018 2731 2026 2817
rect 2018 2725 2019 2731
rect 2025 2725 2026 2731
rect 2018 2663 2026 2725
rect 2018 2657 2019 2663
rect 2025 2657 2026 2663
rect 2018 2567 2026 2657
rect 2018 2561 2019 2567
rect 2025 2561 2026 2567
rect 2018 2495 2026 2561
rect 2018 2489 2019 2495
rect 2025 2489 2026 2495
rect 2018 2413 2026 2489
rect 2018 2407 2019 2413
rect 2025 2407 2026 2413
rect 2018 2327 2026 2407
rect 2018 2321 2019 2327
rect 2025 2321 2026 2327
rect 2018 2231 2026 2321
rect 2018 2225 2019 2231
rect 2025 2225 2026 2231
rect 2018 2171 2026 2225
rect 2018 2165 2019 2171
rect 2025 2165 2026 2171
rect 2018 2051 2026 2165
rect 2018 2045 2019 2051
rect 2025 2045 2026 2051
rect 2018 2015 2026 2045
rect 2018 2009 2019 2015
rect 2025 2009 2026 2015
rect 2018 1883 2026 2009
rect 2018 1877 2019 1883
rect 2025 1877 2026 1883
rect 2018 1863 2026 1877
rect 2018 1857 2019 1863
rect 2025 1857 2026 1863
rect 2018 1723 2026 1857
rect 2018 1717 2019 1723
rect 2025 1717 2026 1723
rect 2018 1707 2026 1717
rect 2018 1701 2019 1707
rect 2025 1701 2026 1707
rect 2018 1567 2026 1701
rect 2018 1561 2019 1567
rect 2025 1561 2026 1567
rect 2018 1551 2026 1561
rect 2018 1545 2019 1551
rect 2025 1545 2026 1551
rect 2018 1399 2026 1545
rect 2018 1393 2019 1399
rect 2025 1393 2026 1399
rect 2018 1239 2026 1393
rect 2018 1233 2019 1239
rect 2025 1233 2026 1239
rect 2018 1227 2026 1233
rect 2018 1221 2019 1227
rect 2025 1221 2026 1227
rect 2018 1075 2026 1221
rect 2018 1069 2019 1075
rect 2025 1069 2026 1075
rect 2018 1063 2026 1069
rect 2018 1057 2019 1063
rect 2025 1057 2026 1063
rect 2018 923 2026 1057
rect 2018 917 2019 923
rect 2025 917 2026 923
rect 2018 899 2026 917
rect 2018 893 2019 899
rect 2025 893 2026 899
rect 2018 771 2026 893
rect 2018 765 2019 771
rect 2025 765 2026 771
rect 2018 743 2026 765
rect 2018 737 2019 743
rect 2025 737 2026 743
rect 2018 619 2026 737
rect 2018 613 2019 619
rect 2025 613 2026 619
rect 2018 579 2026 613
rect 2018 573 2019 579
rect 2025 573 2026 579
rect 2018 435 2026 573
rect 2018 429 2019 435
rect 2025 429 2026 435
rect 2018 427 2026 429
rect 2018 421 2019 427
rect 2025 421 2026 427
rect 2018 271 2026 421
rect 2018 265 2019 271
rect 2025 265 2026 271
rect 2018 91 2026 265
rect 2018 85 2019 91
rect 2025 85 2026 91
rect 2018 72 2026 85
rect 2030 4031 2038 4032
rect 2030 4025 2031 4031
rect 2037 4025 2038 4031
rect 2030 3943 2038 4025
rect 2030 3937 2031 3943
rect 2037 3937 2038 3943
rect 2030 3879 2038 3937
rect 2030 3873 2031 3879
rect 2037 3873 2038 3879
rect 2030 3783 2038 3873
rect 2030 3777 2031 3783
rect 2037 3777 2038 3783
rect 2030 3715 2038 3777
rect 2030 3709 2031 3715
rect 2037 3709 2038 3715
rect 2030 3619 2038 3709
rect 2030 3613 2031 3619
rect 2037 3613 2038 3619
rect 2030 3543 2038 3613
rect 2030 3537 2031 3543
rect 2037 3537 2038 3543
rect 2030 3463 2038 3537
rect 2030 3457 2031 3463
rect 2037 3457 2038 3463
rect 2030 3383 2038 3457
rect 2030 3377 2031 3383
rect 2037 3377 2038 3383
rect 2030 3287 2038 3377
rect 2030 3281 2031 3287
rect 2037 3281 2038 3287
rect 2030 3231 2038 3281
rect 2030 3225 2031 3231
rect 2037 3225 2038 3231
rect 2030 3123 2038 3225
rect 2030 3117 2031 3123
rect 2037 3117 2038 3123
rect 2030 3067 2038 3117
rect 2030 3061 2031 3067
rect 2037 3061 2038 3067
rect 2030 2967 2038 3061
rect 2030 2961 2031 2967
rect 2037 2961 2038 2967
rect 2030 2903 2038 2961
rect 2030 2897 2031 2903
rect 2037 2897 2038 2903
rect 2030 2811 2038 2897
rect 2030 2805 2031 2811
rect 2037 2805 2038 2811
rect 2030 2743 2038 2805
rect 2030 2737 2031 2743
rect 2037 2737 2038 2743
rect 2030 2647 2038 2737
rect 2030 2641 2031 2647
rect 2037 2641 2038 2647
rect 2030 2587 2038 2641
rect 2030 2581 2031 2587
rect 2037 2581 2038 2587
rect 2030 2487 2038 2581
rect 2030 2481 2031 2487
rect 2037 2481 2038 2487
rect 2030 2403 2038 2481
rect 2030 2397 2031 2403
rect 2037 2397 2038 2403
rect 2030 2307 2038 2397
rect 2030 2301 2031 2307
rect 2037 2301 2038 2307
rect 2030 2247 2038 2301
rect 2030 2241 2031 2247
rect 2037 2241 2038 2247
rect 2030 2135 2038 2241
rect 2030 2129 2031 2135
rect 2037 2129 2038 2135
rect 2030 2095 2038 2129
rect 2030 2089 2031 2095
rect 2037 2089 2038 2095
rect 2030 1971 2038 2089
rect 2030 1965 2031 1971
rect 2037 1965 2038 1971
rect 2030 1939 2038 1965
rect 2030 1933 2031 1939
rect 2037 1933 2038 1939
rect 2030 1803 2038 1933
rect 2030 1797 2031 1803
rect 2037 1797 2038 1803
rect 2030 1783 2038 1797
rect 2030 1777 2031 1783
rect 2037 1777 2038 1783
rect 2030 1647 2038 1777
rect 2030 1641 2031 1647
rect 2037 1641 2038 1647
rect 2030 1631 2038 1641
rect 2030 1625 2031 1631
rect 2037 1625 2038 1631
rect 2030 1491 2038 1625
rect 2030 1485 2031 1491
rect 2037 1485 2038 1491
rect 2030 1475 2038 1485
rect 2030 1469 2031 1475
rect 2037 1469 2038 1475
rect 2030 1315 2038 1469
rect 2030 1309 2031 1315
rect 2037 1309 2038 1315
rect 2030 1159 2038 1309
rect 2030 1153 2031 1159
rect 2037 1153 2038 1159
rect 2030 1143 2038 1153
rect 2030 1137 2031 1143
rect 2037 1137 2038 1143
rect 2030 999 2038 1137
rect 2030 993 2031 999
rect 2037 993 2038 999
rect 2030 987 2038 993
rect 2030 981 2031 987
rect 2037 981 2038 987
rect 2030 847 2038 981
rect 2030 841 2031 847
rect 2037 841 2038 847
rect 2030 823 2038 841
rect 2030 817 2031 823
rect 2037 817 2038 823
rect 2030 695 2038 817
rect 2030 689 2031 695
rect 2037 689 2038 695
rect 2030 659 2038 689
rect 2030 653 2031 659
rect 2037 653 2038 659
rect 2030 523 2038 653
rect 2030 517 2031 523
rect 2037 517 2038 523
rect 2030 503 2038 517
rect 2030 497 2031 503
rect 2037 497 2038 503
rect 2030 355 2038 497
rect 2030 349 2031 355
rect 2037 349 2038 355
rect 2030 347 2038 349
rect 2030 341 2031 347
rect 2037 341 2038 347
rect 2030 167 2038 341
rect 2030 161 2031 167
rect 2037 161 2038 167
rect 2030 72 2038 161
rect 3966 4019 3974 4032
rect 3966 4013 3967 4019
rect 3973 4013 3974 4019
rect 3966 3859 3974 4013
rect 3966 3853 3967 3859
rect 3973 3853 3974 3859
rect 3966 3703 3974 3853
rect 3966 3697 3967 3703
rect 3973 3697 3974 3703
rect 3966 3543 3974 3697
rect 3966 3537 3967 3543
rect 3973 3537 3974 3543
rect 3966 3371 3974 3537
rect 3966 3365 3967 3371
rect 3973 3365 3974 3371
rect 3966 3211 3974 3365
rect 3966 3205 3967 3211
rect 3973 3205 3974 3211
rect 3966 3047 3974 3205
rect 3966 3041 3967 3047
rect 3973 3041 3974 3047
rect 3966 2891 3974 3041
rect 3966 2885 3967 2891
rect 3973 2885 3974 2891
rect 3966 2731 3974 2885
rect 3966 2725 3967 2731
rect 3973 2725 3974 2731
rect 3966 2567 3974 2725
rect 3966 2561 3967 2567
rect 3973 2561 3974 2567
rect 3966 2399 3974 2561
rect 3966 2393 3967 2399
rect 3973 2393 3974 2399
rect 3966 2231 3974 2393
rect 3966 2225 3967 2231
rect 3973 2225 3974 2231
rect 3966 2051 3974 2225
rect 3966 2045 3967 2051
rect 3973 2045 3974 2051
rect 3966 1883 3974 2045
rect 3966 1877 3967 1883
rect 3973 1877 3974 1883
rect 3966 1723 3974 1877
rect 3966 1717 3967 1723
rect 3973 1717 3974 1723
rect 3966 1567 3974 1717
rect 3966 1561 3967 1567
rect 3973 1561 3974 1567
rect 3966 1227 3974 1561
rect 3966 1221 3967 1227
rect 3973 1221 3974 1227
rect 3966 1063 3974 1221
rect 3966 1057 3967 1063
rect 3973 1057 3974 1063
rect 3966 899 3974 1057
rect 3966 893 3967 899
rect 3973 893 3974 899
rect 3966 743 3974 893
rect 3966 737 3967 743
rect 3973 737 3974 743
rect 3966 579 3974 737
rect 3966 573 3967 579
rect 3973 573 3974 579
rect 3966 427 3974 573
rect 3966 421 3967 427
rect 3973 421 3974 427
rect 3966 72 3974 421
rect 3978 3943 3986 4032
rect 3978 3937 3979 3943
rect 3985 3937 3986 3943
rect 3978 3783 3986 3937
rect 3978 3777 3979 3783
rect 3985 3777 3986 3783
rect 3978 3619 3986 3777
rect 3978 3613 3979 3619
rect 3985 3613 3986 3619
rect 3978 3463 3986 3613
rect 3978 3457 3979 3463
rect 3985 3457 3986 3463
rect 3978 3287 3986 3457
rect 3978 3281 3979 3287
rect 3985 3281 3986 3287
rect 3978 3123 3986 3281
rect 3978 3117 3979 3123
rect 3985 3117 3986 3123
rect 3978 2967 3986 3117
rect 3978 2961 3979 2967
rect 3985 2961 3986 2967
rect 3978 2811 3986 2961
rect 3978 2805 3979 2811
rect 3985 2805 3986 2811
rect 3978 2647 3986 2805
rect 3978 2641 3979 2647
rect 3985 2641 3986 2647
rect 3978 2487 3986 2641
rect 3978 2481 3979 2487
rect 3985 2481 3986 2487
rect 3978 2307 3986 2481
rect 3978 2301 3979 2307
rect 3985 2301 3986 2307
rect 3978 2135 3986 2301
rect 3978 2129 3979 2135
rect 3985 2129 3986 2135
rect 3978 1971 3986 2129
rect 3978 1965 3979 1971
rect 3985 1965 3986 1971
rect 3978 1803 3986 1965
rect 3978 1797 3979 1803
rect 3985 1797 3986 1803
rect 3978 1647 3986 1797
rect 3978 1641 3979 1647
rect 3985 1641 3986 1647
rect 3978 1491 3986 1641
rect 3978 1485 3979 1491
rect 3985 1485 3986 1491
rect 3978 1143 3986 1485
rect 3978 1137 3979 1143
rect 3985 1137 3986 1143
rect 3978 987 3986 1137
rect 3978 981 3979 987
rect 3985 981 3986 987
rect 3978 823 3986 981
rect 3978 817 3979 823
rect 3985 817 3986 823
rect 3978 659 3986 817
rect 3978 653 3979 659
rect 3985 653 3986 659
rect 3978 503 3986 653
rect 3978 497 3979 503
rect 3985 497 3986 503
rect 3978 347 3986 497
rect 3978 341 3979 347
rect 3985 341 3986 347
rect 3978 72 3986 341
use circuitwell  npwells
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use circuitppnp  ppnps
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use welltap_svt  __well_tap__193
timestamp 1731220359
transform 1 0 3936 0 -1 3988
box 7 3 12 24
use welltap_svt  __well_tap__192
timestamp 1731220359
transform 1 0 2040 0 -1 3988
box 7 3 12 24
use welltap_svt  __well_tap__191
timestamp 1731220359
transform 1 0 3936 0 1 3892
box 7 3 12 24
use welltap_svt  __well_tap__190
timestamp 1731220359
transform 1 0 2040 0 1 3892
box 7 3 12 24
use welltap_svt  __well_tap__189
timestamp 1731220359
transform 1 0 3936 0 -1 3828
box 7 3 12 24
use welltap_svt  __well_tap__188
timestamp 1731220359
transform 1 0 2040 0 -1 3828
box 7 3 12 24
use welltap_svt  __well_tap__187
timestamp 1731220359
transform 1 0 3936 0 1 3732
box 7 3 12 24
use welltap_svt  __well_tap__186
timestamp 1731220359
transform 1 0 2040 0 1 3732
box 7 3 12 24
use welltap_svt  __well_tap__185
timestamp 1731220359
transform 1 0 3936 0 -1 3672
box 7 3 12 24
use welltap_svt  __well_tap__184
timestamp 1731220359
transform 1 0 2040 0 -1 3672
box 7 3 12 24
use welltap_svt  __well_tap__183
timestamp 1731220359
transform 1 0 3936 0 1 3568
box 7 3 12 24
use welltap_svt  __well_tap__182
timestamp 1731220359
transform 1 0 2040 0 1 3568
box 7 3 12 24
use welltap_svt  __well_tap__181
timestamp 1731220359
transform 1 0 3936 0 -1 3512
box 7 3 12 24
use welltap_svt  __well_tap__180
timestamp 1731220359
transform 1 0 2040 0 -1 3512
box 7 3 12 24
use welltap_svt  __well_tap__179
timestamp 1731220359
transform 1 0 3936 0 1 3412
box 7 3 12 24
use welltap_svt  __well_tap__178
timestamp 1731220359
transform 1 0 2040 0 1 3412
box 7 3 12 24
use welltap_svt  __well_tap__177
timestamp 1731220359
transform 1 0 3936 0 -1 3340
box 7 3 12 24
use welltap_svt  __well_tap__176
timestamp 1731220359
transform 1 0 2040 0 -1 3340
box 7 3 12 24
use welltap_svt  __well_tap__175
timestamp 1731220359
transform 1 0 3936 0 1 3236
box 7 3 12 24
use welltap_svt  __well_tap__174
timestamp 1731220359
transform 1 0 2040 0 1 3236
box 7 3 12 24
use welltap_svt  __well_tap__173
timestamp 1731220359
transform 1 0 3936 0 -1 3180
box 7 3 12 24
use welltap_svt  __well_tap__172
timestamp 1731220359
transform 1 0 2040 0 -1 3180
box 7 3 12 24
use welltap_svt  __well_tap__171
timestamp 1731220359
transform 1 0 3936 0 1 3072
box 7 3 12 24
use welltap_svt  __well_tap__170
timestamp 1731220359
transform 1 0 2040 0 1 3072
box 7 3 12 24
use welltap_svt  __well_tap__169
timestamp 1731220359
transform 1 0 3936 0 -1 3016
box 7 3 12 24
use welltap_svt  __well_tap__168
timestamp 1731220359
transform 1 0 2040 0 -1 3016
box 7 3 12 24
use welltap_svt  __well_tap__167
timestamp 1731220359
transform 1 0 3936 0 1 2916
box 7 3 12 24
use welltap_svt  __well_tap__166
timestamp 1731220359
transform 1 0 2040 0 1 2916
box 7 3 12 24
use welltap_svt  __well_tap__165
timestamp 1731220359
transform 1 0 3936 0 -1 2860
box 7 3 12 24
use welltap_svt  __well_tap__164
timestamp 1731220359
transform 1 0 2040 0 -1 2860
box 7 3 12 24
use welltap_svt  __well_tap__163
timestamp 1731220359
transform 1 0 3936 0 1 2760
box 7 3 12 24
use welltap_svt  __well_tap__162
timestamp 1731220359
transform 1 0 2040 0 1 2760
box 7 3 12 24
use welltap_svt  __well_tap__161
timestamp 1731220359
transform 1 0 3936 0 -1 2700
box 7 3 12 24
use welltap_svt  __well_tap__160
timestamp 1731220359
transform 1 0 2040 0 -1 2700
box 7 3 12 24
use welltap_svt  __well_tap__159
timestamp 1731220359
transform 1 0 3936 0 1 2596
box 7 3 12 24
use welltap_svt  __well_tap__158
timestamp 1731220359
transform 1 0 2040 0 1 2596
box 7 3 12 24
use welltap_svt  __well_tap__157
timestamp 1731220359
transform 1 0 3936 0 -1 2536
box 7 3 12 24
use welltap_svt  __well_tap__156
timestamp 1731220359
transform 1 0 2040 0 -1 2536
box 7 3 12 24
use welltap_svt  __well_tap__155
timestamp 1731220359
transform 1 0 3936 0 1 2436
box 7 3 12 24
use welltap_svt  __well_tap__154
timestamp 1731220359
transform 1 0 2040 0 1 2436
box 7 3 12 24
use welltap_svt  __well_tap__153
timestamp 1731220359
transform 1 0 3936 0 -1 2368
box 7 3 12 24
use welltap_svt  __well_tap__152
timestamp 1731220359
transform 1 0 2040 0 -1 2368
box 7 3 12 24
use welltap_svt  __well_tap__151
timestamp 1731220359
transform 1 0 3936 0 1 2256
box 7 3 12 24
use welltap_svt  __well_tap__150
timestamp 1731220359
transform 1 0 2040 0 1 2256
box 7 3 12 24
use welltap_svt  __well_tap__149
timestamp 1731220359
transform 1 0 3936 0 -1 2200
box 7 3 12 24
use welltap_svt  __well_tap__148
timestamp 1731220359
transform 1 0 2040 0 -1 2200
box 7 3 12 24
use welltap_svt  __well_tap__147
timestamp 1731220359
transform 1 0 3936 0 1 2084
box 7 3 12 24
use welltap_svt  __well_tap__146
timestamp 1731220359
transform 1 0 2040 0 1 2084
box 7 3 12 24
use welltap_svt  __well_tap__145
timestamp 1731220359
transform 1 0 3936 0 -1 2020
box 7 3 12 24
use welltap_svt  __well_tap__144
timestamp 1731220359
transform 1 0 2040 0 -1 2020
box 7 3 12 24
use welltap_svt  __well_tap__143
timestamp 1731220359
transform 1 0 3936 0 1 1920
box 7 3 12 24
use welltap_svt  __well_tap__142
timestamp 1731220359
transform 1 0 2040 0 1 1920
box 7 3 12 24
use welltap_svt  __well_tap__141
timestamp 1731220359
transform 1 0 3936 0 -1 1852
box 7 3 12 24
use welltap_svt  __well_tap__140
timestamp 1731220359
transform 1 0 2040 0 -1 1852
box 7 3 12 24
use welltap_svt  __well_tap__139
timestamp 1731220359
transform 1 0 3936 0 1 1752
box 7 3 12 24
use welltap_svt  __well_tap__138
timestamp 1731220359
transform 1 0 2040 0 1 1752
box 7 3 12 24
use welltap_svt  __well_tap__137
timestamp 1731220359
transform 1 0 3936 0 -1 1692
box 7 3 12 24
use welltap_svt  __well_tap__136
timestamp 1731220359
transform 1 0 2040 0 -1 1692
box 7 3 12 24
use welltap_svt  __well_tap__135
timestamp 1731220359
transform 1 0 3936 0 1 1596
box 7 3 12 24
use welltap_svt  __well_tap__134
timestamp 1731220359
transform 1 0 2040 0 1 1596
box 7 3 12 24
use welltap_svt  __well_tap__133
timestamp 1731220359
transform 1 0 3936 0 -1 1536
box 7 3 12 24
use welltap_svt  __well_tap__132
timestamp 1731220359
transform 1 0 2040 0 -1 1536
box 7 3 12 24
use welltap_svt  __well_tap__131
timestamp 1731220359
transform 1 0 3936 0 1 1440
box 7 3 12 24
use welltap_svt  __well_tap__130
timestamp 1731220359
transform 1 0 2040 0 1 1440
box 7 3 12 24
use welltap_svt  __well_tap__129
timestamp 1731220359
transform 1 0 3936 0 -1 1364
box 7 3 12 24
use welltap_svt  __well_tap__128
timestamp 1731220359
transform 1 0 2040 0 -1 1364
box 7 3 12 24
use welltap_svt  __well_tap__127
timestamp 1731220359
transform 1 0 3936 0 1 1260
box 7 3 12 24
use welltap_svt  __well_tap__126
timestamp 1731220359
transform 1 0 2040 0 1 1260
box 7 3 12 24
use welltap_svt  __well_tap__125
timestamp 1731220359
transform 1 0 3936 0 -1 1196
box 7 3 12 24
use welltap_svt  __well_tap__124
timestamp 1731220359
transform 1 0 2040 0 -1 1196
box 7 3 12 24
use welltap_svt  __well_tap__123
timestamp 1731220359
transform 1 0 3936 0 1 1092
box 7 3 12 24
use welltap_svt  __well_tap__122
timestamp 1731220359
transform 1 0 2040 0 1 1092
box 7 3 12 24
use welltap_svt  __well_tap__121
timestamp 1731220359
transform 1 0 3936 0 -1 1032
box 7 3 12 24
use welltap_svt  __well_tap__120
timestamp 1731220359
transform 1 0 2040 0 -1 1032
box 7 3 12 24
use welltap_svt  __well_tap__119
timestamp 1731220359
transform 1 0 3936 0 1 936
box 7 3 12 24
use welltap_svt  __well_tap__118
timestamp 1731220359
transform 1 0 2040 0 1 936
box 7 3 12 24
use welltap_svt  __well_tap__117
timestamp 1731220359
transform 1 0 3936 0 -1 868
box 7 3 12 24
use welltap_svt  __well_tap__116
timestamp 1731220359
transform 1 0 2040 0 -1 868
box 7 3 12 24
use welltap_svt  __well_tap__115
timestamp 1731220359
transform 1 0 3936 0 1 772
box 7 3 12 24
use welltap_svt  __well_tap__114
timestamp 1731220359
transform 1 0 2040 0 1 772
box 7 3 12 24
use welltap_svt  __well_tap__113
timestamp 1731220359
transform 1 0 3936 0 -1 712
box 7 3 12 24
use welltap_svt  __well_tap__112
timestamp 1731220359
transform 1 0 2040 0 -1 712
box 7 3 12 24
use welltap_svt  __well_tap__111
timestamp 1731220359
transform 1 0 3936 0 1 608
box 7 3 12 24
use welltap_svt  __well_tap__110
timestamp 1731220359
transform 1 0 2040 0 1 608
box 7 3 12 24
use welltap_svt  __well_tap__109
timestamp 1731220359
transform 1 0 3936 0 -1 548
box 7 3 12 24
use welltap_svt  __well_tap__108
timestamp 1731220359
transform 1 0 2040 0 -1 548
box 7 3 12 24
use welltap_svt  __well_tap__107
timestamp 1731220359
transform 1 0 3936 0 1 452
box 7 3 12 24
use welltap_svt  __well_tap__106
timestamp 1731220359
transform 1 0 2040 0 1 452
box 7 3 12 24
use welltap_svt  __well_tap__105
timestamp 1731220359
transform 1 0 3936 0 -1 396
box 7 3 12 24
use welltap_svt  __well_tap__104
timestamp 1731220359
transform 1 0 2040 0 -1 396
box 7 3 12 24
use welltap_svt  __well_tap__103
timestamp 1731220359
transform 1 0 3936 0 1 296
box 7 3 12 24
use welltap_svt  __well_tap__102
timestamp 1731220359
transform 1 0 2040 0 1 296
box 7 3 12 24
use welltap_svt  __well_tap__101
timestamp 1731220359
transform 1 0 3936 0 -1 240
box 7 3 12 24
use welltap_svt  __well_tap__100
timestamp 1731220359
transform 1 0 2040 0 -1 240
box 7 3 12 24
use welltap_svt  __well_tap__99
timestamp 1731220359
transform 1 0 3936 0 1 120
box 7 3 12 24
use welltap_svt  __well_tap__98
timestamp 1731220359
transform 1 0 2040 0 1 120
box 7 3 12 24
use welltap_svt  __well_tap__97
timestamp 1731220359
transform 1 0 2000 0 1 3980
box 7 3 12 24
use welltap_svt  __well_tap__96
timestamp 1731220359
transform 1 0 104 0 1 3980
box 7 3 12 24
use welltap_svt  __well_tap__95
timestamp 1731220359
transform 1 0 2000 0 -1 3924
box 7 3 12 24
use welltap_svt  __well_tap__94
timestamp 1731220359
transform 1 0 104 0 -1 3924
box 7 3 12 24
use welltap_svt  __well_tap__93
timestamp 1731220359
transform 1 0 2000 0 1 3828
box 7 3 12 24
use welltap_svt  __well_tap__92
timestamp 1731220359
transform 1 0 104 0 1 3828
box 7 3 12 24
use welltap_svt  __well_tap__91
timestamp 1731220359
transform 1 0 2000 0 -1 3768
box 7 3 12 24
use welltap_svt  __well_tap__90
timestamp 1731220359
transform 1 0 104 0 -1 3768
box 7 3 12 24
use welltap_svt  __well_tap__89
timestamp 1731220359
transform 1 0 2000 0 1 3664
box 7 3 12 24
use welltap_svt  __well_tap__88
timestamp 1731220359
transform 1 0 104 0 1 3664
box 7 3 12 24
use welltap_svt  __well_tap__87
timestamp 1731220359
transform 1 0 2000 0 -1 3600
box 7 3 12 24
use welltap_svt  __well_tap__86
timestamp 1731220359
transform 1 0 104 0 -1 3600
box 7 3 12 24
use welltap_svt  __well_tap__85
timestamp 1731220359
transform 1 0 2000 0 1 3492
box 7 3 12 24
use welltap_svt  __well_tap__84
timestamp 1731220359
transform 1 0 104 0 1 3492
box 7 3 12 24
use welltap_svt  __well_tap__83
timestamp 1731220359
transform 1 0 2000 0 -1 3428
box 7 3 12 24
use welltap_svt  __well_tap__82
timestamp 1731220359
transform 1 0 104 0 -1 3428
box 7 3 12 24
use welltap_svt  __well_tap__81
timestamp 1731220359
transform 1 0 2000 0 1 3332
box 7 3 12 24
use welltap_svt  __well_tap__80
timestamp 1731220359
transform 1 0 104 0 1 3332
box 7 3 12 24
use welltap_svt  __well_tap__79
timestamp 1731220359
transform 1 0 2000 0 -1 3276
box 7 3 12 24
use welltap_svt  __well_tap__78
timestamp 1731220359
transform 1 0 104 0 -1 3276
box 7 3 12 24
use welltap_svt  __well_tap__77
timestamp 1731220359
transform 1 0 2000 0 1 3180
box 7 3 12 24
use welltap_svt  __well_tap__76
timestamp 1731220359
transform 1 0 104 0 1 3180
box 7 3 12 24
use welltap_svt  __well_tap__75
timestamp 1731220359
transform 1 0 2000 0 -1 3120
box 7 3 12 24
use welltap_svt  __well_tap__74
timestamp 1731220359
transform 1 0 104 0 -1 3120
box 7 3 12 24
use welltap_svt  __well_tap__73
timestamp 1731220359
transform 1 0 2000 0 1 3016
box 7 3 12 24
use welltap_svt  __well_tap__72
timestamp 1731220359
transform 1 0 104 0 1 3016
box 7 3 12 24
use welltap_svt  __well_tap__71
timestamp 1731220359
transform 1 0 2000 0 -1 2956
box 7 3 12 24
use welltap_svt  __well_tap__70
timestamp 1731220359
transform 1 0 104 0 -1 2956
box 7 3 12 24
use welltap_svt  __well_tap__69
timestamp 1731220359
transform 1 0 2000 0 1 2852
box 7 3 12 24
use welltap_svt  __well_tap__68
timestamp 1731220359
transform 1 0 104 0 1 2852
box 7 3 12 24
use welltap_svt  __well_tap__67
timestamp 1731220359
transform 1 0 2000 0 -1 2792
box 7 3 12 24
use welltap_svt  __well_tap__66
timestamp 1731220359
transform 1 0 104 0 -1 2792
box 7 3 12 24
use welltap_svt  __well_tap__65
timestamp 1731220359
transform 1 0 2000 0 1 2692
box 7 3 12 24
use welltap_svt  __well_tap__64
timestamp 1731220359
transform 1 0 104 0 1 2692
box 7 3 12 24
use welltap_svt  __well_tap__63
timestamp 1731220359
transform 1 0 2000 0 -1 2632
box 7 3 12 24
use welltap_svt  __well_tap__62
timestamp 1731220359
transform 1 0 104 0 -1 2632
box 7 3 12 24
use welltap_svt  __well_tap__61
timestamp 1731220359
transform 1 0 2000 0 1 2536
box 7 3 12 24
use welltap_svt  __well_tap__60
timestamp 1731220359
transform 1 0 104 0 1 2536
box 7 3 12 24
use welltap_svt  __well_tap__59
timestamp 1731220359
transform 1 0 2000 0 -1 2464
box 7 3 12 24
use welltap_svt  __well_tap__58
timestamp 1731220359
transform 1 0 104 0 -1 2464
box 7 3 12 24
use welltap_svt  __well_tap__57
timestamp 1731220359
transform 1 0 2000 0 1 2352
box 7 3 12 24
use welltap_svt  __well_tap__56
timestamp 1731220359
transform 1 0 104 0 1 2352
box 7 3 12 24
use welltap_svt  __well_tap__55
timestamp 1731220359
transform 1 0 2000 0 -1 2296
box 7 3 12 24
use welltap_svt  __well_tap__54
timestamp 1731220359
transform 1 0 104 0 -1 2296
box 7 3 12 24
use welltap_svt  __well_tap__53
timestamp 1731220359
transform 1 0 2000 0 1 2196
box 7 3 12 24
use welltap_svt  __well_tap__52
timestamp 1731220359
transform 1 0 104 0 1 2196
box 7 3 12 24
use welltap_svt  __well_tap__51
timestamp 1731220359
transform 1 0 2000 0 -1 2140
box 7 3 12 24
use welltap_svt  __well_tap__50
timestamp 1731220359
transform 1 0 104 0 -1 2140
box 7 3 12 24
use welltap_svt  __well_tap__49
timestamp 1731220359
transform 1 0 2000 0 1 2044
box 7 3 12 24
use welltap_svt  __well_tap__48
timestamp 1731220359
transform 1 0 104 0 1 2044
box 7 3 12 24
use welltap_svt  __well_tap__47
timestamp 1731220359
transform 1 0 2000 0 -1 1984
box 7 3 12 24
use welltap_svt  __well_tap__46
timestamp 1731220359
transform 1 0 104 0 -1 1984
box 7 3 12 24
use welltap_svt  __well_tap__45
timestamp 1731220359
transform 1 0 2000 0 1 1888
box 7 3 12 24
use welltap_svt  __well_tap__44
timestamp 1731220359
transform 1 0 104 0 1 1888
box 7 3 12 24
use welltap_svt  __well_tap__43
timestamp 1731220359
transform 1 0 2000 0 -1 1832
box 7 3 12 24
use welltap_svt  __well_tap__42
timestamp 1731220359
transform 1 0 104 0 -1 1832
box 7 3 12 24
use welltap_svt  __well_tap__41
timestamp 1731220359
transform 1 0 2000 0 1 1732
box 7 3 12 24
use welltap_svt  __well_tap__40
timestamp 1731220359
transform 1 0 104 0 1 1732
box 7 3 12 24
use welltap_svt  __well_tap__39
timestamp 1731220359
transform 1 0 2000 0 -1 1676
box 7 3 12 24
use welltap_svt  __well_tap__38
timestamp 1731220359
transform 1 0 104 0 -1 1676
box 7 3 12 24
use welltap_svt  __well_tap__37
timestamp 1731220359
transform 1 0 2000 0 1 1580
box 7 3 12 24
use welltap_svt  __well_tap__36
timestamp 1731220359
transform 1 0 104 0 1 1580
box 7 3 12 24
use welltap_svt  __well_tap__35
timestamp 1731220359
transform 1 0 2000 0 -1 1520
box 7 3 12 24
use welltap_svt  __well_tap__34
timestamp 1731220359
transform 1 0 104 0 -1 1520
box 7 3 12 24
use welltap_svt  __well_tap__33
timestamp 1731220359
transform 1 0 2000 0 1 1424
box 7 3 12 24
use welltap_svt  __well_tap__32
timestamp 1731220359
transform 1 0 104 0 1 1424
box 7 3 12 24
use welltap_svt  __well_tap__31
timestamp 1731220359
transform 1 0 2000 0 -1 1368
box 7 3 12 24
use welltap_svt  __well_tap__30
timestamp 1731220359
transform 1 0 104 0 -1 1368
box 7 3 12 24
use welltap_svt  __well_tap__29
timestamp 1731220359
transform 1 0 2000 0 1 1264
box 7 3 12 24
use welltap_svt  __well_tap__28
timestamp 1731220359
transform 1 0 104 0 1 1264
box 7 3 12 24
use welltap_svt  __well_tap__27
timestamp 1731220359
transform 1 0 2000 0 -1 1208
box 7 3 12 24
use welltap_svt  __well_tap__26
timestamp 1731220359
transform 1 0 104 0 -1 1208
box 7 3 12 24
use welltap_svt  __well_tap__25
timestamp 1731220359
transform 1 0 2000 0 1 1108
box 7 3 12 24
use welltap_svt  __well_tap__24
timestamp 1731220359
transform 1 0 104 0 1 1108
box 7 3 12 24
use welltap_svt  __well_tap__23
timestamp 1731220359
transform 1 0 2000 0 -1 1044
box 7 3 12 24
use welltap_svt  __well_tap__22
timestamp 1731220359
transform 1 0 104 0 -1 1044
box 7 3 12 24
use welltap_svt  __well_tap__21
timestamp 1731220359
transform 1 0 2000 0 1 948
box 7 3 12 24
use welltap_svt  __well_tap__20
timestamp 1731220359
transform 1 0 104 0 1 948
box 7 3 12 24
use welltap_svt  __well_tap__19
timestamp 1731220359
transform 1 0 2000 0 -1 892
box 7 3 12 24
use welltap_svt  __well_tap__18
timestamp 1731220359
transform 1 0 104 0 -1 892
box 7 3 12 24
use welltap_svt  __well_tap__17
timestamp 1731220359
transform 1 0 2000 0 1 796
box 7 3 12 24
use welltap_svt  __well_tap__16
timestamp 1731220359
transform 1 0 104 0 1 796
box 7 3 12 24
use welltap_svt  __well_tap__15
timestamp 1731220359
transform 1 0 2000 0 -1 740
box 7 3 12 24
use welltap_svt  __well_tap__14
timestamp 1731220359
transform 1 0 104 0 -1 740
box 7 3 12 24
use welltap_svt  __well_tap__13
timestamp 1731220359
transform 1 0 2000 0 1 644
box 7 3 12 24
use welltap_svt  __well_tap__12
timestamp 1731220359
transform 1 0 104 0 1 644
box 7 3 12 24
use welltap_svt  __well_tap__11
timestamp 1731220359
transform 1 0 2000 0 -1 588
box 7 3 12 24
use welltap_svt  __well_tap__10
timestamp 1731220359
transform 1 0 104 0 -1 588
box 7 3 12 24
use welltap_svt  __well_tap__9
timestamp 1731220359
transform 1 0 2000 0 1 472
box 7 3 12 24
use welltap_svt  __well_tap__8
timestamp 1731220359
transform 1 0 104 0 1 472
box 7 3 12 24
use welltap_svt  __well_tap__7
timestamp 1731220359
transform 1 0 2000 0 -1 404
box 7 3 12 24
use welltap_svt  __well_tap__6
timestamp 1731220359
transform 1 0 104 0 -1 404
box 7 3 12 24
use welltap_svt  __well_tap__5
timestamp 1731220359
transform 1 0 2000 0 1 304
box 7 3 12 24
use welltap_svt  __well_tap__4
timestamp 1731220359
transform 1 0 104 0 1 304
box 7 3 12 24
use welltap_svt  __well_tap__3
timestamp 1731220359
transform 1 0 2000 0 -1 240
box 7 3 12 24
use welltap_svt  __well_tap__2
timestamp 1731220359
transform 1 0 104 0 -1 240
box 7 3 12 24
use welltap_svt  __well_tap__1
timestamp 1731220359
transform 1 0 2000 0 1 116
box 7 3 12 24
use welltap_svt  __well_tap__0
timestamp 1731220359
transform 1 0 104 0 1 116
box 7 3 12 24
use _0_0cell_0_0gcelem3x0  tst_5999_6
timestamp 1731220359
transform 1 0 3680 0 -1 3540
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5998_6
timestamp 1731220359
transform 1 0 3832 0 -1 3540
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5997_6
timestamp 1731220359
transform 1 0 3832 0 -1 3368
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5996_6
timestamp 1731220359
transform 1 0 3832 0 -1 3208
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5995_6
timestamp 1731220359
transform 1 0 3832 0 -1 3044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5994_6
timestamp 1731220359
transform 1 0 3832 0 -1 2888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5993_6
timestamp 1731220359
transform 1 0 3832 0 1 2732
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5992_6
timestamp 1731220359
transform 1 0 3832 0 -1 2728
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5991_6
timestamp 1731220359
transform 1 0 3648 0 -1 2728
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5990_6
timestamp 1731220359
transform 1 0 3664 0 1 2732
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5989_6
timestamp 1731220359
transform 1 0 3792 0 1 3044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5988_6
timestamp 1731220359
transform 1 0 3784 0 1 3208
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5987_6
timestamp 1731220359
transform 1 0 3768 0 1 3384
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5986_6
timestamp 1731220359
transform 1 0 3744 0 -1 3700
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5985_6
timestamp 1731220359
transform 1 0 3704 0 1 3704
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5984_6
timestamp 1731220359
transform 1 0 3648 0 -1 3856
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5983_6
timestamp 1731220359
transform 1 0 3736 0 1 3864
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5982_6
timestamp 1731220359
transform 1 0 3624 0 1 3864
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5981_6
timestamp 1731220359
transform 1 0 3512 0 1 3864
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5980_6
timestamp 1731220359
transform 1 0 3400 0 1 3864
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5979_6
timestamp 1731220359
transform 1 0 3296 0 1 3864
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5978_6
timestamp 1731220359
transform 1 0 3184 0 1 3864
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5977_6
timestamp 1731220359
transform 1 0 3064 0 1 3864
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5976_6
timestamp 1731220359
transform 1 0 2944 0 1 3864
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5975_6
timestamp 1731220359
transform 1 0 2816 0 1 3864
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5974_6
timestamp 1731220359
transform 1 0 3008 0 -1 3856
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5973_6
timestamp 1731220359
transform 1 0 3216 0 -1 3856
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5972_6
timestamp 1731220359
transform 1 0 3432 0 -1 3856
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5971_6
timestamp 1731220359
transform 1 0 3312 0 1 3704
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5970_6
timestamp 1731220359
transform 1 0 3120 0 1 3704
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5969_6
timestamp 1731220359
transform 1 0 2928 0 1 3704
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5968_6
timestamp 1731220359
transform 1 0 3504 0 1 3704
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5967_6
timestamp 1731220359
transform 1 0 3504 0 -1 3700
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5966_6
timestamp 1731220359
transform 1 0 3272 0 -1 3700
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5965_6
timestamp 1731220359
transform 1 0 3040 0 -1 3700
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5964_6
timestamp 1731220359
transform 1 0 3448 0 1 3540
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5963_6
timestamp 1731220359
transform 1 0 3616 0 1 3540
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5962_6
timestamp 1731220359
transform 1 0 3512 0 -1 3540
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5961_6
timestamp 1731220359
transform 1 0 3344 0 -1 3540
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5960_6
timestamp 1731220359
transform 1 0 3400 0 1 3384
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5959_6
timestamp 1731220359
transform 1 0 3584 0 1 3384
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5958_6
timestamp 1731220359
transform 1 0 3688 0 -1 3368
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5957_6
timestamp 1731220359
transform 1 0 3528 0 -1 3368
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5956_6
timestamp 1731220359
transform 1 0 3368 0 -1 3368
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5955_6
timestamp 1731220359
transform 1 0 3520 0 1 3208
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5954_6
timestamp 1731220359
transform 1 0 3216 0 -1 3368
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5953_6
timestamp 1731220359
transform 1 0 3072 0 -1 3368
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5952_6
timestamp 1731220359
transform 1 0 2928 0 -1 3368
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5951_6
timestamp 1731220359
transform 1 0 2856 0 1 3384
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5950_6
timestamp 1731220359
transform 1 0 3040 0 1 3384
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5949_6
timestamp 1731220359
transform 1 0 3216 0 1 3384
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5948_6
timestamp 1731220359
transform 1 0 3168 0 -1 3540
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5947_6
timestamp 1731220359
transform 1 0 2992 0 -1 3540
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5946_6
timestamp 1731220359
transform 1 0 3288 0 1 3540
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5945_6
timestamp 1731220359
transform 1 0 3136 0 1 3540
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5944_6
timestamp 1731220359
transform 1 0 2992 0 1 3540
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5943_6
timestamp 1731220359
transform 1 0 2848 0 1 3540
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5942_6
timestamp 1731220359
transform 1 0 2712 0 1 3540
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5941_6
timestamp 1731220359
transform 1 0 2576 0 1 3540
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5940_6
timestamp 1731220359
transform 1 0 2448 0 1 3540
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5939_6
timestamp 1731220359
transform 1 0 2320 0 1 3540
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5938_6
timestamp 1731220359
transform 1 0 2440 0 -1 3540
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5937_6
timestamp 1731220359
transform 1 0 2624 0 -1 3540
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5936_6
timestamp 1731220359
transform 1 0 2808 0 -1 3540
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5935_6
timestamp 1731220359
transform 1 0 2672 0 1 3384
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5934_6
timestamp 1731220359
transform 1 0 2488 0 1 3384
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5933_6
timestamp 1731220359
transform 1 0 2304 0 1 3384
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5932_6
timestamp 1731220359
transform 1 0 2352 0 -1 3368
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5931_6
timestamp 1731220359
transform 1 0 2504 0 -1 3368
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5930_6
timestamp 1731220359
transform 1 0 2648 0 -1 3368
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5929_6
timestamp 1731220359
transform 1 0 2792 0 -1 3368
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5928_6
timestamp 1731220359
transform 1 0 3008 0 1 3208
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5927_6
timestamp 1731220359
transform 1 0 2776 0 1 3208
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5926_6
timestamp 1731220359
transform 1 0 2568 0 1 3208
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5925_6
timestamp 1731220359
transform 1 0 2392 0 1 3208
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5924_6
timestamp 1731220359
transform 1 0 2240 0 1 3208
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5923_6
timestamp 1731220359
transform 1 0 2256 0 -1 3208
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5922_6
timestamp 1731220359
transform 1 0 2352 0 -1 3208
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5921_6
timestamp 1731220359
transform 1 0 2448 0 -1 3208
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5920_6
timestamp 1731220359
transform 1 0 2544 0 -1 3208
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5919_6
timestamp 1731220359
transform 1 0 2640 0 -1 3208
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5918_6
timestamp 1731220359
transform 1 0 2736 0 -1 3208
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5917_6
timestamp 1731220359
transform 1 0 2832 0 -1 3208
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5916_6
timestamp 1731220359
transform 1 0 2928 0 -1 3208
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5915_6
timestamp 1731220359
transform 1 0 3024 0 -1 3208
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5914_6
timestamp 1731220359
transform 1 0 3120 0 -1 3208
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5913_6
timestamp 1731220359
transform 1 0 3216 0 -1 3208
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5912_6
timestamp 1731220359
transform 1 0 3256 0 1 3208
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5911_6
timestamp 1731220359
transform 1 0 3312 0 -1 3208
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5910_6
timestamp 1731220359
transform 1 0 3432 0 -1 3208
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5909_6
timestamp 1731220359
transform 1 0 3712 0 -1 3208
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5908_6
timestamp 1731220359
transform 1 0 3568 0 -1 3208
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5907_6
timestamp 1731220359
transform 1 0 3496 0 1 3044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5906_6
timestamp 1731220359
transform 1 0 3200 0 1 3044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5905_6
timestamp 1731220359
transform 1 0 2904 0 1 3044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5904_6
timestamp 1731220359
transform 1 0 2616 0 1 3044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5903_6
timestamp 1731220359
transform 1 0 2696 0 -1 3044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5902_6
timestamp 1731220359
transform 1 0 2992 0 -1 3044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5901_6
timestamp 1731220359
transform 1 0 3280 0 -1 3044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5900_6
timestamp 1731220359
transform 1 0 3568 0 -1 3044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5899_6
timestamp 1731220359
transform 1 0 3832 0 1 2888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5898_6
timestamp 1731220359
transform 1 0 3640 0 1 2888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5897_6
timestamp 1731220359
transform 1 0 3432 0 1 2888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5896_6
timestamp 1731220359
transform 1 0 3208 0 1 2888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5895_6
timestamp 1731220359
transform 1 0 2968 0 1 2888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5894_6
timestamp 1731220359
transform 1 0 2696 0 1 2888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5893_6
timestamp 1731220359
transform 1 0 3640 0 -1 2888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5892_6
timestamp 1731220359
transform 1 0 3424 0 -1 2888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5891_6
timestamp 1731220359
transform 1 0 3208 0 -1 2888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5890_6
timestamp 1731220359
transform 1 0 2984 0 -1 2888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5889_6
timestamp 1731220359
transform 1 0 3472 0 1 2732
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5888_6
timestamp 1731220359
transform 1 0 3288 0 1 2732
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5887_6
timestamp 1731220359
transform 1 0 3104 0 1 2732
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5886_6
timestamp 1731220359
transform 1 0 2920 0 1 2732
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5885_6
timestamp 1731220359
transform 1 0 3448 0 -1 2728
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5884_6
timestamp 1731220359
transform 1 0 3248 0 -1 2728
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5883_6
timestamp 1731220359
transform 1 0 3056 0 -1 2728
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5882_6
timestamp 1731220359
transform 1 0 2880 0 -1 2728
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5881_6
timestamp 1731220359
transform 1 0 2720 0 -1 2728
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5880_6
timestamp 1731220359
transform 1 0 2784 0 1 2568
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5879_6
timestamp 1731220359
transform 1 0 2904 0 1 2568
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5878_6
timestamp 1731220359
transform 1 0 3144 0 1 2568
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5877_6
timestamp 1731220359
transform 1 0 3024 0 1 2568
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5876_6
timestamp 1731220359
transform 1 0 2984 0 -1 2564
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5875_6
timestamp 1731220359
transform 1 0 3104 0 -1 2564
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5874_6
timestamp 1731220359
transform 1 0 3224 0 -1 2564
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5873_6
timestamp 1731220359
transform 1 0 3352 0 -1 2564
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5872_6
timestamp 1731220359
transform 1 0 3480 0 -1 2564
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5871_6
timestamp 1731220359
transform 1 0 3352 0 1 2408
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5870_6
timestamp 1731220359
transform 1 0 3200 0 1 2408
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5869_6
timestamp 1731220359
transform 1 0 3496 0 1 2408
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5868_6
timestamp 1731220359
transform 1 0 3648 0 1 2408
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5867_6
timestamp 1731220359
transform 1 0 3800 0 1 2408
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5866_6
timestamp 1731220359
transform 1 0 3832 0 -1 2396
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5865_6
timestamp 1731220359
transform 1 0 3672 0 -1 2396
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5864_6
timestamp 1731220359
transform 1 0 3512 0 -1 2396
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5863_6
timestamp 1731220359
transform 1 0 3352 0 -1 2396
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5862_6
timestamp 1731220359
transform 1 0 3184 0 -1 2396
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5861_6
timestamp 1731220359
transform 1 0 3688 0 1 2228
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5860_6
timestamp 1731220359
transform 1 0 3528 0 1 2228
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5859_6
timestamp 1731220359
transform 1 0 3376 0 1 2228
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5858_6
timestamp 1731220359
transform 1 0 3224 0 1 2228
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5857_6
timestamp 1731220359
transform 1 0 3064 0 1 2228
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5856_6
timestamp 1731220359
transform 1 0 3512 0 -1 2228
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5855_6
timestamp 1731220359
transform 1 0 3360 0 -1 2228
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5854_6
timestamp 1731220359
transform 1 0 3216 0 -1 2228
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5853_6
timestamp 1731220359
transform 1 0 3072 0 -1 2228
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5852_6
timestamp 1731220359
transform 1 0 2928 0 -1 2228
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5851_6
timestamp 1731220359
transform 1 0 3512 0 1 2056
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5850_6
timestamp 1731220359
transform 1 0 3344 0 1 2056
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5849_6
timestamp 1731220359
transform 1 0 3184 0 1 2056
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5848_6
timestamp 1731220359
transform 1 0 3032 0 1 2056
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5847_6
timestamp 1731220359
transform 1 0 2888 0 1 2056
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5846_6
timestamp 1731220359
transform 1 0 3448 0 -1 2048
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5845_6
timestamp 1731220359
transform 1 0 3256 0 -1 2048
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5844_6
timestamp 1731220359
transform 1 0 3072 0 -1 2048
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5843_6
timestamp 1731220359
transform 1 0 2912 0 -1 2048
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5842_6
timestamp 1731220359
transform 1 0 2768 0 -1 2048
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5841_6
timestamp 1731220359
transform 1 0 2760 0 1 1892
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5840_6
timestamp 1731220359
transform 1 0 2912 0 1 1892
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5839_6
timestamp 1731220359
transform 1 0 3096 0 1 1892
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5838_6
timestamp 1731220359
transform 1 0 3312 0 1 1892
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5837_6
timestamp 1731220359
transform 1 0 3536 0 1 1892
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5836_6
timestamp 1731220359
transform 1 0 3624 0 -1 1880
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5835_6
timestamp 1731220359
transform 1 0 3392 0 -1 1880
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5834_6
timestamp 1731220359
transform 1 0 3176 0 -1 1880
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5833_6
timestamp 1731220359
transform 1 0 2984 0 -1 1880
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5832_6
timestamp 1731220359
transform 1 0 2824 0 -1 1880
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5831_6
timestamp 1731220359
transform 1 0 2872 0 1 1724
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5830_6
timestamp 1731220359
transform 1 0 3064 0 1 1724
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5829_6
timestamp 1731220359
transform 1 0 3256 0 1 1724
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5828_6
timestamp 1731220359
transform 1 0 3456 0 1 1724
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5827_6
timestamp 1731220359
transform 1 0 3440 0 -1 1720
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5826_6
timestamp 1731220359
transform 1 0 3248 0 -1 1720
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5825_6
timestamp 1731220359
transform 1 0 3056 0 -1 1720
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5824_6
timestamp 1731220359
transform 1 0 3040 0 1 1568
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5823_6
timestamp 1731220359
transform 1 0 2832 0 1 1568
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5822_6
timestamp 1731220359
transform 1 0 3224 0 1 1568
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5821_6
timestamp 1731220359
transform 1 0 3392 0 1 1568
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5820_6
timestamp 1731220359
transform 1 0 3376 0 -1 1564
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5819_6
timestamp 1731220359
transform 1 0 3216 0 -1 1564
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5818_6
timestamp 1731220359
transform 1 0 3536 0 -1 1564
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5817_6
timestamp 1731220359
transform 1 0 3696 0 -1 1564
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5816_6
timestamp 1731220359
transform 1 0 3688 0 1 1568
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5815_6
timestamp 1731220359
transform 1 0 3544 0 1 1568
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5814_6
timestamp 1731220359
transform 1 0 3640 0 -1 1720
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5813_6
timestamp 1731220359
transform 1 0 3656 0 1 1724
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5812_6
timestamp 1731220359
transform 1 0 3768 0 1 1892
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5811_6
timestamp 1731220359
transform 1 0 3832 0 1 2056
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5810_6
timestamp 1731220359
transform 1 0 3680 0 1 2056
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5809_6
timestamp 1731220359
transform 1 0 3648 0 -1 2048
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5808_6
timestamp 1731220359
transform 1 0 3832 0 -1 2048
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5807_6
timestamp 1731220359
transform 1 0 3832 0 -1 1880
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5806_6
timestamp 1731220359
transform 1 0 3832 0 1 1724
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5805_6
timestamp 1731220359
transform 1 0 3832 0 -1 1720
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5804_6
timestamp 1731220359
transform 1 0 3832 0 1 1568
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5803_6
timestamp 1731220359
transform 1 0 3808 0 1 1412
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5802_6
timestamp 1731220359
transform 1 0 3808 0 -1 1392
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5801_6
timestamp 1731220359
transform 1 0 3824 0 1 1232
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5800_6
timestamp 1731220359
transform 1 0 3832 0 -1 1224
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5799_6
timestamp 1731220359
transform 1 0 3832 0 1 1064
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5798_6
timestamp 1731220359
transform 1 0 3832 0 -1 1060
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5797_6
timestamp 1731220359
transform 1 0 3832 0 1 908
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5796_6
timestamp 1731220359
transform 1 0 3832 0 -1 896
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5795_6
timestamp 1731220359
transform 1 0 3832 0 1 744
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5794_6
timestamp 1731220359
transform 1 0 3832 0 -1 740
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5793_6
timestamp 1731220359
transform 1 0 3824 0 1 580
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5792_6
timestamp 1731220359
transform 1 0 3832 0 -1 576
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5791_6
timestamp 1731220359
transform 1 0 3640 0 -1 576
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5790_6
timestamp 1731220359
transform 1 0 3448 0 -1 576
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5789_6
timestamp 1731220359
transform 1 0 3296 0 1 580
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5788_6
timestamp 1731220359
transform 1 0 3472 0 1 580
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5787_6
timestamp 1731220359
transform 1 0 3648 0 1 580
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5786_6
timestamp 1731220359
transform 1 0 3672 0 -1 740
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5785_6
timestamp 1731220359
transform 1 0 3512 0 -1 740
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5784_6
timestamp 1731220359
transform 1 0 3360 0 -1 740
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5783_6
timestamp 1731220359
transform 1 0 3208 0 -1 740
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5782_6
timestamp 1731220359
transform 1 0 3240 0 1 744
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5781_6
timestamp 1731220359
transform 1 0 3440 0 1 744
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5780_6
timestamp 1731220359
transform 1 0 3648 0 1 744
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5779_6
timestamp 1731220359
transform 1 0 3608 0 -1 896
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5778_6
timestamp 1731220359
transform 1 0 3360 0 -1 896
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5777_6
timestamp 1731220359
transform 1 0 3120 0 -1 896
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5776_6
timestamp 1731220359
transform 1 0 3656 0 1 908
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5775_6
timestamp 1731220359
transform 1 0 3456 0 1 908
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5774_6
timestamp 1731220359
transform 1 0 3272 0 1 908
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5773_6
timestamp 1731220359
transform 1 0 3104 0 1 908
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5772_6
timestamp 1731220359
transform 1 0 2960 0 1 908
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5771_6
timestamp 1731220359
transform 1 0 3000 0 -1 1060
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5770_6
timestamp 1731220359
transform 1 0 3624 0 -1 1060
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5769_6
timestamp 1731220359
transform 1 0 3400 0 -1 1060
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5768_6
timestamp 1731220359
transform 1 0 3192 0 -1 1060
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5767_6
timestamp 1731220359
transform 1 0 3144 0 1 1064
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5766_6
timestamp 1731220359
transform 1 0 2984 0 1 1064
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5765_6
timestamp 1731220359
transform 1 0 3312 0 1 1064
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5764_6
timestamp 1731220359
transform 1 0 3672 0 1 1064
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5763_6
timestamp 1731220359
transform 1 0 3488 0 1 1064
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5762_6
timestamp 1731220359
transform 1 0 3392 0 -1 1224
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5761_6
timestamp 1731220359
transform 1 0 3232 0 -1 1224
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5760_6
timestamp 1731220359
transform 1 0 3064 0 -1 1224
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5759_6
timestamp 1731220359
transform 1 0 3544 0 -1 1224
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5758_6
timestamp 1731220359
transform 1 0 3696 0 -1 1224
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5757_6
timestamp 1731220359
transform 1 0 3656 0 1 1232
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5756_6
timestamp 1731220359
transform 1 0 3496 0 1 1232
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5755_6
timestamp 1731220359
transform 1 0 3336 0 1 1232
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5754_6
timestamp 1731220359
transform 1 0 3168 0 1 1232
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5753_6
timestamp 1731220359
transform 1 0 2992 0 1 1232
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5752_6
timestamp 1731220359
transform 1 0 3552 0 -1 1392
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5751_6
timestamp 1731220359
transform 1 0 3296 0 -1 1392
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5750_6
timestamp 1731220359
transform 1 0 3048 0 -1 1392
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5749_6
timestamp 1731220359
transform 1 0 2800 0 -1 1392
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5748_6
timestamp 1731220359
transform 1 0 2552 0 -1 1392
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5747_6
timestamp 1731220359
transform 1 0 3608 0 1 1412
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5746_6
timestamp 1731220359
transform 1 0 3408 0 1 1412
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5745_6
timestamp 1731220359
transform 1 0 3224 0 1 1412
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5744_6
timestamp 1731220359
transform 1 0 3056 0 1 1412
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5743_6
timestamp 1731220359
transform 1 0 2912 0 1 1412
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5742_6
timestamp 1731220359
transform 1 0 2792 0 1 1412
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5741_6
timestamp 1731220359
transform 1 0 2696 0 1 1412
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5740_6
timestamp 1731220359
transform 1 0 2600 0 1 1412
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5739_6
timestamp 1731220359
transform 1 0 2504 0 1 1412
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5738_6
timestamp 1731220359
transform 1 0 2408 0 1 1412
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5737_6
timestamp 1731220359
transform 1 0 3056 0 -1 1564
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5736_6
timestamp 1731220359
transform 1 0 2896 0 -1 1564
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5735_6
timestamp 1731220359
transform 1 0 2736 0 -1 1564
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5734_6
timestamp 1731220359
transform 1 0 2576 0 -1 1564
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5733_6
timestamp 1731220359
transform 1 0 2592 0 1 1568
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5732_6
timestamp 1731220359
transform 1 0 2680 0 -1 1720
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5731_6
timestamp 1731220359
transform 1 0 2864 0 -1 1720
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5730_6
timestamp 1731220359
transform 1 0 2680 0 1 1724
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5729_6
timestamp 1731220359
transform 1 0 2696 0 -1 1880
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5728_6
timestamp 1731220359
transform 1 0 2584 0 -1 1880
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5727_6
timestamp 1731220359
transform 1 0 2640 0 1 1892
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5726_6
timestamp 1731220359
transform 1 0 2640 0 -1 2048
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5725_6
timestamp 1731220359
transform 1 0 2624 0 1 2056
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5724_6
timestamp 1731220359
transform 1 0 2752 0 1 2056
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5723_6
timestamp 1731220359
transform 1 0 2776 0 -1 2228
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5722_6
timestamp 1731220359
transform 1 0 2904 0 1 2228
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5721_6
timestamp 1731220359
transform 1 0 2808 0 -1 2396
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5720_6
timestamp 1731220359
transform 1 0 2600 0 -1 2396
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5719_6
timestamp 1731220359
transform 1 0 3000 0 -1 2396
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5718_6
timestamp 1731220359
transform 1 0 3040 0 1 2408
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5717_6
timestamp 1731220359
transform 1 0 2872 0 1 2408
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5716_6
timestamp 1731220359
transform 1 0 2704 0 1 2408
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5715_6
timestamp 1731220359
transform 1 0 2528 0 1 2408
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5714_6
timestamp 1731220359
transform 1 0 2864 0 -1 2564
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5713_6
timestamp 1731220359
transform 1 0 2736 0 -1 2564
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5712_6
timestamp 1731220359
transform 1 0 2608 0 -1 2564
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5711_6
timestamp 1731220359
transform 1 0 2488 0 -1 2564
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5710_6
timestamp 1731220359
transform 1 0 2376 0 -1 2564
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5709_6
timestamp 1731220359
transform 1 0 2664 0 1 2568
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5708_6
timestamp 1731220359
transform 1 0 2552 0 1 2568
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5707_6
timestamp 1731220359
transform 1 0 2440 0 1 2568
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5706_6
timestamp 1731220359
transform 1 0 2328 0 1 2568
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5705_6
timestamp 1731220359
transform 1 0 2224 0 1 2568
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5704_6
timestamp 1731220359
transform 1 0 2576 0 -1 2728
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5703_6
timestamp 1731220359
transform 1 0 2440 0 -1 2728
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5702_6
timestamp 1731220359
transform 1 0 2312 0 -1 2728
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5701_6
timestamp 1731220359
transform 1 0 2184 0 -1 2728
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5700_6
timestamp 1731220359
transform 1 0 2064 0 -1 2728
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5699_6
timestamp 1731220359
transform 1 0 2728 0 1 2732
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5698_6
timestamp 1731220359
transform 1 0 2544 0 1 2732
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5697_6
timestamp 1731220359
transform 1 0 2360 0 1 2732
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5696_6
timestamp 1731220359
transform 1 0 2192 0 1 2732
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5695_6
timestamp 1731220359
transform 1 0 2064 0 1 2732
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5694_6
timestamp 1731220359
transform 1 0 2760 0 -1 2888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5693_6
timestamp 1731220359
transform 1 0 2528 0 -1 2888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5692_6
timestamp 1731220359
transform 1 0 2288 0 -1 2888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5691_6
timestamp 1731220359
transform 1 0 2064 0 -1 2888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5690_6
timestamp 1731220359
transform 1 0 2064 0 1 2888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5689_6
timestamp 1731220359
transform 1 0 2384 0 1 2888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5688_6
timestamp 1731220359
transform 1 0 2376 0 -1 3044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5687_6
timestamp 1731220359
transform 1 0 2064 0 -1 3044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5686_6
timestamp 1731220359
transform 1 0 2064 0 1 3044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5685_6
timestamp 1731220359
transform 1 0 2328 0 1 3044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5684_6
timestamp 1731220359
transform 1 0 2160 0 -1 3208
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5683_6
timestamp 1731220359
transform 1 0 2064 0 -1 3208
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5682_6
timestamp 1731220359
transform 1 0 2104 0 1 3208
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5681_6
timestamp 1731220359
transform 1 0 2064 0 -1 3368
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5680_6
timestamp 1731220359
transform 1 0 2208 0 -1 3368
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5679_6
timestamp 1731220359
transform 1 0 2120 0 1 3384
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5678_6
timestamp 1731220359
transform 1 0 2096 0 -1 3540
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5677_6
timestamp 1731220359
transform 1 0 2264 0 -1 3540
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5676_6
timestamp 1731220359
transform 1 0 2184 0 1 3540
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5675_6
timestamp 1731220359
transform 1 0 2120 0 -1 3700
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5674_6
timestamp 1731220359
transform 1 0 2344 0 -1 3700
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5673_6
timestamp 1731220359
transform 1 0 2576 0 -1 3700
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5672_6
timestamp 1731220359
transform 1 0 2808 0 -1 3700
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5671_6
timestamp 1731220359
transform 1 0 2736 0 1 3704
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5670_6
timestamp 1731220359
transform 1 0 2552 0 1 3704
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5669_6
timestamp 1731220359
transform 1 0 2368 0 1 3704
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5668_6
timestamp 1731220359
transform 1 0 2184 0 1 3704
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5667_6
timestamp 1731220359
transform 1 0 2200 0 -1 3856
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5666_6
timestamp 1731220359
transform 1 0 2336 0 -1 3856
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5665_6
timestamp 1731220359
transform 1 0 2480 0 -1 3856
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5664_6
timestamp 1731220359
transform 1 0 2640 0 -1 3856
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5663_6
timestamp 1731220359
transform 1 0 2816 0 -1 3856
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5662_6
timestamp 1731220359
transform 1 0 2680 0 1 3864
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5661_6
timestamp 1731220359
transform 1 0 2544 0 1 3864
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5660_6
timestamp 1731220359
transform 1 0 2408 0 1 3864
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5659_6
timestamp 1731220359
transform 1 0 2280 0 1 3864
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5658_6
timestamp 1731220359
transform 1 0 2152 0 1 3864
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5657_6
timestamp 1731220359
transform 1 0 2256 0 -1 4016
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5656_6
timestamp 1731220359
transform 1 0 2160 0 -1 4016
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5655_6
timestamp 1731220359
transform 1 0 2064 0 -1 4016
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5654_6
timestamp 1731220359
transform 1 0 1896 0 1 3952
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5653_6
timestamp 1731220359
transform 1 0 1800 0 1 3952
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5652_6
timestamp 1731220359
transform 1 0 1704 0 1 3952
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5651_6
timestamp 1731220359
transform 1 0 1608 0 1 3952
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5650_6
timestamp 1731220359
transform 1 0 1512 0 1 3952
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5649_6
timestamp 1731220359
transform 1 0 1640 0 -1 3952
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5648_6
timestamp 1731220359
transform 1 0 1504 0 -1 3952
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5647_6
timestamp 1731220359
transform 1 0 1376 0 -1 3952
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5646_6
timestamp 1731220359
transform 1 0 1248 0 -1 3952
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5645_6
timestamp 1731220359
transform 1 0 1120 0 -1 3952
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5644_6
timestamp 1731220359
transform 1 0 1096 0 1 3800
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5643_6
timestamp 1731220359
transform 1 0 1224 0 1 3800
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5642_6
timestamp 1731220359
transform 1 0 1352 0 1 3800
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5641_6
timestamp 1731220359
transform 1 0 1480 0 1 3800
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5640_6
timestamp 1731220359
transform 1 0 1424 0 -1 3796
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5639_6
timestamp 1731220359
transform 1 0 1280 0 -1 3796
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5638_6
timestamp 1731220359
transform 1 0 1576 0 -1 3796
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5637_6
timestamp 1731220359
transform 1 0 1488 0 1 3636
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5636_6
timestamp 1731220359
transform 1 0 1648 0 1 3636
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5635_6
timestamp 1731220359
transform 1 0 1608 0 -1 3628
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5634_6
timestamp 1731220359
transform 1 0 1432 0 -1 3628
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5633_6
timestamp 1731220359
transform 1 0 1784 0 -1 3628
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5632_6
timestamp 1731220359
transform 1 0 1872 0 1 3464
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5631_6
timestamp 1731220359
transform 1 0 1696 0 1 3464
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5630_6
timestamp 1731220359
transform 1 0 1520 0 1 3464
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5629_6
timestamp 1731220359
transform 1 0 1528 0 -1 3456
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5628_6
timestamp 1731220359
transform 1 0 1712 0 -1 3456
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5627_6
timestamp 1731220359
transform 1 0 1896 0 -1 3456
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5626_6
timestamp 1731220359
transform 1 0 1864 0 1 3304
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5625_6
timestamp 1731220359
transform 1 0 1696 0 1 3304
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5624_6
timestamp 1731220359
transform 1 0 1536 0 1 3304
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5623_6
timestamp 1731220359
transform 1 0 1512 0 -1 3304
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5622_6
timestamp 1731220359
transform 1 0 1736 0 -1 3304
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5621_6
timestamp 1731220359
transform 1 0 1688 0 1 3152
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5620_6
timestamp 1731220359
transform 1 0 1504 0 1 3152
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5619_6
timestamp 1731220359
transform 1 0 1384 0 -1 3148
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5618_6
timestamp 1731220359
transform 1 0 1552 0 -1 3148
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5617_6
timestamp 1731220359
transform 1 0 1720 0 -1 3148
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5616_6
timestamp 1731220359
transform 1 0 1712 0 1 2988
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5615_6
timestamp 1731220359
transform 1 0 1544 0 1 2988
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5614_6
timestamp 1731220359
transform 1 0 1480 0 -1 2984
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5613_6
timestamp 1731220359
transform 1 0 1648 0 -1 2984
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5612_6
timestamp 1731220359
transform 1 0 1816 0 -1 2984
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5611_6
timestamp 1731220359
transform 1 0 1840 0 1 2824
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5610_6
timestamp 1731220359
transform 1 0 1664 0 1 2824
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5609_6
timestamp 1731220359
transform 1 0 1488 0 1 2824
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5608_6
timestamp 1731220359
transform 1 0 1592 0 -1 2820
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5607_6
timestamp 1731220359
transform 1 0 1776 0 -1 2820
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5606_6
timestamp 1731220359
transform 1 0 1776 0 1 2664
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5605_6
timestamp 1731220359
transform 1 0 1616 0 1 2664
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5604_6
timestamp 1731220359
transform 1 0 1456 0 1 2664
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5603_6
timestamp 1731220359
transform 1 0 1424 0 -1 2660
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5602_6
timestamp 1731220359
transform 1 0 1560 0 -1 2660
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5601_6
timestamp 1731220359
transform 1 0 1696 0 -1 2660
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5600_6
timestamp 1731220359
transform 1 0 1720 0 1 2508
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5599_6
timestamp 1731220359
transform 1 0 1584 0 1 2508
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5598_6
timestamp 1731220359
transform 1 0 1456 0 1 2508
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5597_6
timestamp 1731220359
transform 1 0 1328 0 1 2508
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5596_6
timestamp 1731220359
transform 1 0 1192 0 1 2508
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5595_6
timestamp 1731220359
transform 1 0 1056 0 1 2508
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5594_6
timestamp 1731220359
transform 1 0 912 0 1 2508
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5593_6
timestamp 1731220359
transform 1 0 1024 0 -1 2660
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5592_6
timestamp 1731220359
transform 1 0 1160 0 -1 2660
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5591_6
timestamp 1731220359
transform 1 0 1296 0 -1 2660
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5590_6
timestamp 1731220359
transform 1 0 1304 0 1 2664
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5589_6
timestamp 1731220359
transform 1 0 1152 0 1 2664
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5588_6
timestamp 1731220359
transform 1 0 1072 0 -1 2820
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5587_6
timestamp 1731220359
transform 1 0 1232 0 -1 2820
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5586_6
timestamp 1731220359
transform 1 0 1408 0 -1 2820
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5585_6
timestamp 1731220359
transform 1 0 1312 0 1 2824
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5584_6
timestamp 1731220359
transform 1 0 1144 0 1 2824
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5583_6
timestamp 1731220359
transform 1 0 1320 0 -1 2984
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5582_6
timestamp 1731220359
transform 1 0 1168 0 -1 2984
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5581_6
timestamp 1731220359
transform 1 0 1064 0 1 2988
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5580_6
timestamp 1731220359
transform 1 0 1216 0 1 2988
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5579_6
timestamp 1731220359
transform 1 0 1376 0 1 2988
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5578_6
timestamp 1731220359
transform 1 0 1216 0 -1 3148
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5577_6
timestamp 1731220359
transform 1 0 1056 0 -1 3148
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5576_6
timestamp 1731220359
transform 1 0 960 0 1 3152
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5575_6
timestamp 1731220359
transform 1 0 1136 0 1 3152
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5574_6
timestamp 1731220359
transform 1 0 1320 0 1 3152
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5573_6
timestamp 1731220359
transform 1 0 1288 0 -1 3304
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5572_6
timestamp 1731220359
transform 1 0 1072 0 -1 3304
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5571_6
timestamp 1731220359
transform 1 0 1040 0 1 3304
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5570_6
timestamp 1731220359
transform 1 0 1208 0 1 3304
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5569_6
timestamp 1731220359
transform 1 0 1376 0 1 3304
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5568_6
timestamp 1731220359
transform 1 0 1344 0 -1 3456
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5567_6
timestamp 1731220359
transform 1 0 1152 0 -1 3456
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5566_6
timestamp 1731220359
transform 1 0 952 0 -1 3456
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5565_6
timestamp 1731220359
transform 1 0 992 0 1 3464
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5564_6
timestamp 1731220359
transform 1 0 1168 0 1 3464
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5563_6
timestamp 1731220359
transform 1 0 1344 0 1 3464
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5562_6
timestamp 1731220359
transform 1 0 1256 0 -1 3628
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5561_6
timestamp 1731220359
transform 1 0 1088 0 -1 3628
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5560_6
timestamp 1731220359
transform 1 0 1032 0 1 3636
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5559_6
timestamp 1731220359
transform 1 0 1328 0 1 3636
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5558_6
timestamp 1731220359
transform 1 0 1176 0 1 3636
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5557_6
timestamp 1731220359
transform 1 0 1136 0 -1 3796
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5556_6
timestamp 1731220359
transform 1 0 992 0 -1 3796
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5555_6
timestamp 1731220359
transform 1 0 968 0 1 3800
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5554_6
timestamp 1731220359
transform 1 0 840 0 1 3800
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5553_6
timestamp 1731220359
transform 1 0 712 0 1 3800
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5552_6
timestamp 1731220359
transform 1 0 992 0 -1 3952
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5551_6
timestamp 1731220359
transform 1 0 864 0 -1 3952
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5550_6
timestamp 1731220359
transform 1 0 736 0 -1 3952
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5549_6
timestamp 1731220359
transform 1 0 608 0 -1 3952
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5548_6
timestamp 1731220359
transform 1 0 488 0 -1 3952
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5547_6
timestamp 1731220359
transform 1 0 384 0 -1 3952
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5546_6
timestamp 1731220359
transform 1 0 288 0 -1 3952
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5545_6
timestamp 1731220359
transform 1 0 192 0 -1 3952
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5544_6
timestamp 1731220359
transform 1 0 328 0 1 3800
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5543_6
timestamp 1731220359
transform 1 0 448 0 1 3800
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5542_6
timestamp 1731220359
transform 1 0 576 0 1 3800
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5541_6
timestamp 1731220359
transform 1 0 496 0 -1 3796
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5540_6
timestamp 1731220359
transform 1 0 608 0 -1 3796
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5539_6
timestamp 1731220359
transform 1 0 728 0 -1 3796
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5538_6
timestamp 1731220359
transform 1 0 856 0 -1 3796
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5537_6
timestamp 1731220359
transform 1 0 904 0 1 3636
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5536_6
timestamp 1731220359
transform 1 0 784 0 1 3636
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5535_6
timestamp 1731220359
transform 1 0 680 0 1 3636
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5534_6
timestamp 1731220359
transform 1 0 584 0 1 3636
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5533_6
timestamp 1731220359
transform 1 0 488 0 1 3636
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5532_6
timestamp 1731220359
transform 1 0 920 0 -1 3628
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5531_6
timestamp 1731220359
transform 1 0 752 0 -1 3628
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5530_6
timestamp 1731220359
transform 1 0 600 0 -1 3628
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5529_6
timestamp 1731220359
transform 1 0 456 0 -1 3628
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5528_6
timestamp 1731220359
transform 1 0 328 0 -1 3628
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5527_6
timestamp 1731220359
transform 1 0 808 0 1 3464
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5526_6
timestamp 1731220359
transform 1 0 632 0 1 3464
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5525_6
timestamp 1731220359
transform 1 0 456 0 1 3464
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5524_6
timestamp 1731220359
transform 1 0 296 0 1 3464
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5523_6
timestamp 1731220359
transform 1 0 152 0 1 3464
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5522_6
timestamp 1731220359
transform 1 0 744 0 -1 3456
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5521_6
timestamp 1731220359
transform 1 0 528 0 -1 3456
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5520_6
timestamp 1731220359
transform 1 0 312 0 -1 3456
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5519_6
timestamp 1731220359
transform 1 0 128 0 -1 3456
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5518_6
timestamp 1731220359
transform 1 0 864 0 1 3304
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5517_6
timestamp 1731220359
transform 1 0 696 0 1 3304
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5516_6
timestamp 1731220359
transform 1 0 528 0 1 3304
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5515_6
timestamp 1731220359
transform 1 0 368 0 1 3304
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5514_6
timestamp 1731220359
transform 1 0 224 0 1 3304
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5513_6
timestamp 1731220359
transform 1 0 128 0 1 3304
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5512_6
timestamp 1731220359
transform 1 0 128 0 -1 3304
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5511_6
timestamp 1731220359
transform 1 0 272 0 -1 3304
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5510_6
timestamp 1731220359
transform 1 0 864 0 -1 3304
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5509_6
timestamp 1731220359
transform 1 0 656 0 -1 3304
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5508_6
timestamp 1731220359
transform 1 0 456 0 -1 3304
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5507_6
timestamp 1731220359
transform 1 0 440 0 1 3152
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5506_6
timestamp 1731220359
transform 1 0 280 0 1 3152
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5505_6
timestamp 1731220359
transform 1 0 128 0 1 3152
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5504_6
timestamp 1731220359
transform 1 0 608 0 1 3152
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5503_6
timestamp 1731220359
transform 1 0 784 0 1 3152
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5502_6
timestamp 1731220359
transform 1 0 896 0 -1 3148
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5501_6
timestamp 1731220359
transform 1 0 736 0 -1 3148
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5500_6
timestamp 1731220359
transform 1 0 576 0 -1 3148
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5499_6
timestamp 1731220359
transform 1 0 432 0 -1 3148
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5498_6
timestamp 1731220359
transform 1 0 304 0 -1 3148
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5497_6
timestamp 1731220359
transform 1 0 496 0 1 2988
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5496_6
timestamp 1731220359
transform 1 0 592 0 1 2988
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5495_6
timestamp 1731220359
transform 1 0 696 0 1 2988
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5494_6
timestamp 1731220359
transform 1 0 808 0 1 2988
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5493_6
timestamp 1731220359
transform 1 0 928 0 1 2988
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5492_6
timestamp 1731220359
transform 1 0 1016 0 -1 2984
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5491_6
timestamp 1731220359
transform 1 0 880 0 -1 2984
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5490_6
timestamp 1731220359
transform 1 0 752 0 -1 2984
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5489_6
timestamp 1731220359
transform 1 0 640 0 -1 2984
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5488_6
timestamp 1731220359
transform 1 0 544 0 -1 2984
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5487_6
timestamp 1731220359
transform 1 0 984 0 1 2824
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5486_6
timestamp 1731220359
transform 1 0 832 0 1 2824
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5485_6
timestamp 1731220359
transform 1 0 688 0 1 2824
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5484_6
timestamp 1731220359
transform 1 0 568 0 1 2824
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5483_6
timestamp 1731220359
transform 1 0 464 0 1 2824
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5482_6
timestamp 1731220359
transform 1 0 472 0 -1 2820
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5481_6
timestamp 1731220359
transform 1 0 568 0 -1 2820
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5480_6
timestamp 1731220359
transform 1 0 672 0 -1 2820
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5479_6
timestamp 1731220359
transform 1 0 792 0 -1 2820
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5478_6
timestamp 1731220359
transform 1 0 928 0 -1 2820
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5477_6
timestamp 1731220359
transform 1 0 1008 0 1 2664
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5476_6
timestamp 1731220359
transform 1 0 872 0 1 2664
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5475_6
timestamp 1731220359
transform 1 0 736 0 1 2664
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5474_6
timestamp 1731220359
transform 1 0 616 0 1 2664
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5473_6
timestamp 1731220359
transform 1 0 504 0 1 2664
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5472_6
timestamp 1731220359
transform 1 0 888 0 -1 2660
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5471_6
timestamp 1731220359
transform 1 0 744 0 -1 2660
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5470_6
timestamp 1731220359
transform 1 0 608 0 -1 2660
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5469_6
timestamp 1731220359
transform 1 0 480 0 -1 2660
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5468_6
timestamp 1731220359
transform 1 0 360 0 -1 2660
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5467_6
timestamp 1731220359
transform 1 0 760 0 1 2508
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5466_6
timestamp 1731220359
transform 1 0 600 0 1 2508
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5465_6
timestamp 1731220359
transform 1 0 440 0 1 2508
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5464_6
timestamp 1731220359
transform 1 0 280 0 1 2508
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5463_6
timestamp 1731220359
transform 1 0 128 0 1 2508
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5462_6
timestamp 1731220359
transform 1 0 512 0 -1 2492
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5461_6
timestamp 1731220359
transform 1 0 416 0 -1 2492
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5460_6
timestamp 1731220359
transform 1 0 320 0 -1 2492
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5459_6
timestamp 1731220359
transform 1 0 224 0 -1 2492
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5458_6
timestamp 1731220359
transform 1 0 128 0 -1 2492
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5457_6
timestamp 1731220359
transform 1 0 128 0 1 2324
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5456_6
timestamp 1731220359
transform 1 0 248 0 1 2324
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5455_6
timestamp 1731220359
transform 1 0 408 0 1 2324
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5454_6
timestamp 1731220359
transform 1 0 568 0 1 2324
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5453_6
timestamp 1731220359
transform 1 0 728 0 1 2324
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5452_6
timestamp 1731220359
transform 1 0 736 0 -1 2324
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5451_6
timestamp 1731220359
transform 1 0 576 0 -1 2324
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5450_6
timestamp 1731220359
transform 1 0 416 0 -1 2324
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5449_6
timestamp 1731220359
transform 1 0 256 0 -1 2324
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5448_6
timestamp 1731220359
transform 1 0 128 0 -1 2324
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5447_6
timestamp 1731220359
transform 1 0 216 0 1 2168
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5446_6
timestamp 1731220359
transform 1 0 344 0 1 2168
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5445_6
timestamp 1731220359
transform 1 0 488 0 1 2168
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5444_6
timestamp 1731220359
transform 1 0 640 0 1 2168
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5443_6
timestamp 1731220359
transform 1 0 792 0 1 2168
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5442_6
timestamp 1731220359
transform 1 0 672 0 -1 2168
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5441_6
timestamp 1731220359
transform 1 0 560 0 -1 2168
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5440_6
timestamp 1731220359
transform 1 0 464 0 -1 2168
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5439_6
timestamp 1731220359
transform 1 0 800 0 -1 2168
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5438_6
timestamp 1731220359
transform 1 0 936 0 -1 2168
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5437_6
timestamp 1731220359
transform 1 0 1112 0 1 2016
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5436_6
timestamp 1731220359
transform 1 0 976 0 1 2016
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5435_6
timestamp 1731220359
transform 1 0 848 0 1 2016
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5434_6
timestamp 1731220359
transform 1 0 728 0 1 2016
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5433_6
timestamp 1731220359
transform 1 0 616 0 1 2016
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5432_6
timestamp 1731220359
transform 1 0 880 0 -1 2012
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5431_6
timestamp 1731220359
transform 1 0 720 0 -1 2012
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5430_6
timestamp 1731220359
transform 1 0 568 0 -1 2012
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5429_6
timestamp 1731220359
transform 1 0 440 0 -1 2012
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5428_6
timestamp 1731220359
transform 1 0 440 0 -1 1860
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5427_6
timestamp 1731220359
transform 1 0 312 0 -1 1860
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5426_6
timestamp 1731220359
transform 1 0 248 0 1 1704
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5425_6
timestamp 1731220359
transform 1 0 384 0 1 1704
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5424_6
timestamp 1731220359
transform 1 0 424 0 -1 1704
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5423_6
timestamp 1731220359
transform 1 0 256 0 -1 1704
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5422_6
timestamp 1731220359
transform 1 0 128 0 -1 1704
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5421_6
timestamp 1731220359
transform 1 0 128 0 1 1552
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5420_6
timestamp 1731220359
transform 1 0 280 0 1 1552
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5419_6
timestamp 1731220359
transform 1 0 480 0 -1 1548
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5418_6
timestamp 1731220359
transform 1 0 288 0 -1 1548
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5417_6
timestamp 1731220359
transform 1 0 128 0 -1 1548
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5416_6
timestamp 1731220359
transform 1 0 168 0 1 1396
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5415_6
timestamp 1731220359
transform 1 0 352 0 1 1396
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5414_6
timestamp 1731220359
transform 1 0 320 0 -1 1396
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5413_6
timestamp 1731220359
transform 1 0 560 0 1 1396
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5412_6
timestamp 1731220359
transform 1 0 776 0 1 1396
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5411_6
timestamp 1731220359
transform 1 0 880 0 -1 1548
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5410_6
timestamp 1731220359
transform 1 0 680 0 -1 1548
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5409_6
timestamp 1731220359
transform 1 0 648 0 1 1552
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5408_6
timestamp 1731220359
transform 1 0 464 0 1 1552
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5407_6
timestamp 1731220359
transform 1 0 832 0 1 1552
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5406_6
timestamp 1731220359
transform 1 0 792 0 -1 1704
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5405_6
timestamp 1731220359
transform 1 0 600 0 -1 1704
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5404_6
timestamp 1731220359
transform 1 0 528 0 1 1704
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5403_6
timestamp 1731220359
transform 1 0 688 0 1 1704
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5402_6
timestamp 1731220359
transform 1 0 856 0 1 1704
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5401_6
timestamp 1731220359
transform 1 0 848 0 -1 1860
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5400_6
timestamp 1731220359
transform 1 0 712 0 -1 1860
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5399_6
timestamp 1731220359
transform 1 0 576 0 -1 1860
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5398_6
timestamp 1731220359
transform 1 0 648 0 1 1860
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5397_6
timestamp 1731220359
transform 1 0 744 0 1 1860
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5396_6
timestamp 1731220359
transform 1 0 840 0 1 1860
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5395_6
timestamp 1731220359
transform 1 0 936 0 1 1860
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5394_6
timestamp 1731220359
transform 1 0 1032 0 1 1860
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5393_6
timestamp 1731220359
transform 1 0 1048 0 -1 2012
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5392_6
timestamp 1731220359
transform 1 0 1128 0 1 1860
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5391_6
timestamp 1731220359
transform 1 0 1224 0 -1 2012
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5390_6
timestamp 1731220359
transform 1 0 1248 0 1 2016
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5389_6
timestamp 1731220359
transform 1 0 1216 0 -1 2168
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5388_6
timestamp 1731220359
transform 1 0 1072 0 -1 2168
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5387_6
timestamp 1731220359
transform 1 0 1112 0 1 2168
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5386_6
timestamp 1731220359
transform 1 0 952 0 1 2168
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5385_6
timestamp 1731220359
transform 1 0 1040 0 -1 2324
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5384_6
timestamp 1731220359
transform 1 0 888 0 -1 2324
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5383_6
timestamp 1731220359
transform 1 0 880 0 1 2324
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5382_6
timestamp 1731220359
transform 1 0 1032 0 1 2324
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5381_6
timestamp 1731220359
transform 1 0 1176 0 1 2324
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5380_6
timestamp 1731220359
transform 1 0 1320 0 1 2324
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5379_6
timestamp 1731220359
transform 1 0 1472 0 1 2324
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5378_6
timestamp 1731220359
transform 1 0 1496 0 -1 2324
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5377_6
timestamp 1731220359
transform 1 0 1344 0 -1 2324
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5376_6
timestamp 1731220359
transform 1 0 1192 0 -1 2324
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5375_6
timestamp 1731220359
transform 1 0 1272 0 1 2168
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5374_6
timestamp 1731220359
transform 1 0 1432 0 1 2168
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5373_6
timestamp 1731220359
transform 1 0 1592 0 1 2168
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5372_6
timestamp 1731220359
transform 1 0 1496 0 -1 2168
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5371_6
timestamp 1731220359
transform 1 0 1360 0 -1 2168
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5370_6
timestamp 1731220359
transform 1 0 1632 0 -1 2168
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5369_6
timestamp 1731220359
transform 1 0 1648 0 1 2016
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5368_6
timestamp 1731220359
transform 1 0 1520 0 1 2016
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5367_6
timestamp 1731220359
transform 1 0 1384 0 1 2016
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5366_6
timestamp 1731220359
transform 1 0 1392 0 -1 2012
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5365_6
timestamp 1731220359
transform 1 0 1568 0 -1 2012
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5364_6
timestamp 1731220359
transform 1 0 1744 0 -1 2012
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5363_6
timestamp 1731220359
transform 1 0 1896 0 -1 2012
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5362_6
timestamp 1731220359
transform 1 0 1896 0 1 2016
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5361_6
timestamp 1731220359
transform 1 0 1784 0 1 2016
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5360_6
timestamp 1731220359
transform 1 0 1776 0 -1 2168
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5359_6
timestamp 1731220359
transform 1 0 1896 0 -1 2168
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5358_6
timestamp 1731220359
transform 1 0 2064 0 -1 2228
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5357_6
timestamp 1731220359
transform 1 0 2168 0 -1 2228
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5356_6
timestamp 1731220359
transform 1 0 2160 0 1 2228
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5355_6
timestamp 1731220359
transform 1 0 2064 0 1 2228
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5354_6
timestamp 1731220359
transform 1 0 2264 0 1 2228
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5353_6
timestamp 1731220359
transform 1 0 2408 0 1 2228
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5352_6
timestamp 1731220359
transform 1 0 2568 0 1 2228
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5351_6
timestamp 1731220359
transform 1 0 2736 0 1 2228
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5350_6
timestamp 1731220359
transform 1 0 2616 0 -1 2228
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5349_6
timestamp 1731220359
transform 1 0 2464 0 -1 2228
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5348_6
timestamp 1731220359
transform 1 0 2312 0 -1 2228
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5347_6
timestamp 1731220359
transform 1 0 2272 0 1 2056
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5346_6
timestamp 1731220359
transform 1 0 2384 0 1 2056
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5345_6
timestamp 1731220359
transform 1 0 2504 0 1 2056
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5344_6
timestamp 1731220359
transform 1 0 2424 0 -1 2048
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5343_6
timestamp 1731220359
transform 1 0 2320 0 -1 2048
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5342_6
timestamp 1731220359
transform 1 0 2528 0 -1 2048
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5341_6
timestamp 1731220359
transform 1 0 2536 0 1 1892
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5340_6
timestamp 1731220359
transform 1 0 2440 0 1 1892
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5339_6
timestamp 1731220359
transform 1 0 2344 0 1 1892
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5338_6
timestamp 1731220359
transform 1 0 2248 0 1 1892
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5337_6
timestamp 1731220359
transform 1 0 2480 0 -1 1880
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5336_6
timestamp 1731220359
transform 1 0 2376 0 -1 1880
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5335_6
timestamp 1731220359
transform 1 0 2272 0 -1 1880
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5334_6
timestamp 1731220359
transform 1 0 2176 0 -1 1880
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5333_6
timestamp 1731220359
transform 1 0 2120 0 1 1724
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5332_6
timestamp 1731220359
transform 1 0 2304 0 1 1724
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5331_6
timestamp 1731220359
transform 1 0 2488 0 1 1724
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5330_6
timestamp 1731220359
transform 1 0 2504 0 -1 1720
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5329_6
timestamp 1731220359
transform 1 0 2336 0 -1 1720
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5328_6
timestamp 1731220359
transform 1 0 2184 0 -1 1720
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5327_6
timestamp 1731220359
transform 1 0 2064 0 -1 1720
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5326_6
timestamp 1731220359
transform 1 0 2328 0 1 1568
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5325_6
timestamp 1731220359
transform 1 0 2064 0 1 1568
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5324_6
timestamp 1731220359
transform 1 0 1896 0 1 1552
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5323_6
timestamp 1731220359
transform 1 0 1776 0 1 1552
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5322_6
timestamp 1731220359
transform 1 0 1632 0 1 1552
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5321_6
timestamp 1731220359
transform 1 0 1488 0 1 1552
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5320_6
timestamp 1731220359
transform 1 0 1616 0 -1 1704
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5319_6
timestamp 1731220359
transform 1 0 1832 0 -1 1704
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5318_6
timestamp 1731220359
transform 1 0 1736 0 1 1704
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5317_6
timestamp 1731220359
transform 1 0 1552 0 1 1704
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5316_6
timestamp 1731220359
transform 1 0 1376 0 1 1704
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5315_6
timestamp 1731220359
transform 1 0 1392 0 -1 1860
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5314_6
timestamp 1731220359
transform 1 0 1528 0 -1 1860
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5313_6
timestamp 1731220359
transform 1 0 1416 0 1 1860
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5312_6
timestamp 1731220359
transform 1 0 1320 0 1 1860
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5311_6
timestamp 1731220359
transform 1 0 1224 0 1 1860
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5310_6
timestamp 1731220359
transform 1 0 1256 0 -1 1860
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5309_6
timestamp 1731220359
transform 1 0 1120 0 -1 1860
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5308_6
timestamp 1731220359
transform 1 0 984 0 -1 1860
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5307_6
timestamp 1731220359
transform 1 0 1200 0 1 1704
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5306_6
timestamp 1731220359
transform 1 0 1024 0 1 1704
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5305_6
timestamp 1731220359
transform 1 0 992 0 -1 1704
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5304_6
timestamp 1731220359
transform 1 0 1400 0 -1 1704
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5303_6
timestamp 1731220359
transform 1 0 1192 0 -1 1704
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5302_6
timestamp 1731220359
transform 1 0 1176 0 1 1552
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5301_6
timestamp 1731220359
transform 1 0 1008 0 1 1552
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5300_6
timestamp 1731220359
transform 1 0 1336 0 1 1552
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5299_6
timestamp 1731220359
transform 1 0 1256 0 -1 1548
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5298_6
timestamp 1731220359
transform 1 0 1072 0 -1 1548
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5297_6
timestamp 1731220359
transform 1 0 1440 0 -1 1548
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5296_6
timestamp 1731220359
transform 1 0 1616 0 -1 1548
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5295_6
timestamp 1731220359
transform 1 0 1800 0 -1 1548
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5294_6
timestamp 1731220359
transform 1 0 1896 0 1 1396
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5293_6
timestamp 1731220359
transform 1 0 1688 0 1 1396
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5292_6
timestamp 1731220359
transform 1 0 1456 0 1 1396
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5291_6
timestamp 1731220359
transform 1 0 1744 0 -1 1396
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5290_6
timestamp 1731220359
transform 1 0 1896 0 -1 1396
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5289_6
timestamp 1731220359
transform 1 0 2064 0 -1 1392
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5288_6
timestamp 1731220359
transform 1 0 2296 0 -1 1392
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5287_6
timestamp 1731220359
transform 1 0 2216 0 1 1232
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5286_6
timestamp 1731220359
transform 1 0 2064 0 1 1232
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5285_6
timestamp 1731220359
transform 1 0 2408 0 1 1232
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5284_6
timestamp 1731220359
transform 1 0 2808 0 1 1232
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5283_6
timestamp 1731220359
transform 1 0 2608 0 1 1232
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5282_6
timestamp 1731220359
transform 1 0 2496 0 -1 1224
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5281_6
timestamp 1731220359
transform 1 0 2304 0 -1 1224
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5280_6
timestamp 1731220359
transform 1 0 2128 0 -1 1224
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5279_6
timestamp 1731220359
transform 1 0 2688 0 -1 1224
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5278_6
timestamp 1731220359
transform 1 0 2880 0 -1 1224
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5277_6
timestamp 1731220359
transform 1 0 2832 0 1 1064
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5276_6
timestamp 1731220359
transform 1 0 2688 0 1 1064
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5275_6
timestamp 1731220359
transform 1 0 2552 0 1 1064
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5274_6
timestamp 1731220359
transform 1 0 2416 0 1 1064
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5273_6
timestamp 1731220359
transform 1 0 2288 0 1 1064
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5272_6
timestamp 1731220359
transform 1 0 2488 0 -1 1060
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5271_6
timestamp 1731220359
transform 1 0 2592 0 -1 1060
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5270_6
timestamp 1731220359
transform 1 0 2704 0 -1 1060
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5269_6
timestamp 1731220359
transform 1 0 2840 0 -1 1060
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5268_6
timestamp 1731220359
transform 1 0 2840 0 1 908
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5267_6
timestamp 1731220359
transform 1 0 2736 0 1 908
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5266_6
timestamp 1731220359
transform 1 0 2640 0 1 908
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5265_6
timestamp 1731220359
transform 1 0 2672 0 -1 896
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5264_6
timestamp 1731220359
transform 1 0 2888 0 -1 896
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5263_6
timestamp 1731220359
transform 1 0 2888 0 1 744
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5262_6
timestamp 1731220359
transform 1 0 3056 0 1 744
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5261_6
timestamp 1731220359
transform 1 0 3056 0 -1 740
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5260_6
timestamp 1731220359
transform 1 0 3120 0 1 580
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5259_6
timestamp 1731220359
transform 1 0 2936 0 1 580
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5258_6
timestamp 1731220359
transform 1 0 2872 0 -1 576
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5257_6
timestamp 1731220359
transform 1 0 3064 0 -1 576
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5256_6
timestamp 1731220359
transform 1 0 3256 0 -1 576
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5255_6
timestamp 1731220359
transform 1 0 3152 0 1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5254_6
timestamp 1731220359
transform 1 0 2952 0 1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5253_6
timestamp 1731220359
transform 1 0 3360 0 1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5252_6
timestamp 1731220359
transform 1 0 3576 0 1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5251_6
timestamp 1731220359
transform 1 0 3408 0 -1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5250_6
timestamp 1731220359
transform 1 0 3256 0 -1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5249_6
timestamp 1731220359
transform 1 0 3104 0 -1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5248_6
timestamp 1731220359
transform 1 0 3552 0 -1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5247_6
timestamp 1731220359
transform 1 0 3704 0 -1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5246_6
timestamp 1731220359
transform 1 0 3704 0 1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5245_6
timestamp 1731220359
transform 1 0 3800 0 1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5244_6
timestamp 1731220359
transform 1 0 3832 0 -1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5243_6
timestamp 1731220359
transform 1 0 3832 0 1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5242_6
timestamp 1731220359
transform 1 0 3832 0 -1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5241_6
timestamp 1731220359
transform 1 0 3832 0 1 92
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5240_6
timestamp 1731220359
transform 1 0 3688 0 1 92
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5239_6
timestamp 1731220359
transform 1 0 3560 0 1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5238_6
timestamp 1731220359
transform 1 0 3416 0 1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5237_6
timestamp 1731220359
transform 1 0 3264 0 1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5236_6
timestamp 1731220359
transform 1 0 3664 0 -1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5235_6
timestamp 1731220359
transform 1 0 3472 0 -1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5234_6
timestamp 1731220359
transform 1 0 3280 0 -1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5233_6
timestamp 1731220359
transform 1 0 3088 0 -1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5232_6
timestamp 1731220359
transform 1 0 3528 0 1 92
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5231_6
timestamp 1731220359
transform 1 0 3376 0 1 92
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5230_6
timestamp 1731220359
transform 1 0 3232 0 1 92
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5229_6
timestamp 1731220359
transform 1 0 3096 0 1 92
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5228_6
timestamp 1731220359
transform 1 0 2968 0 1 92
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5227_6
timestamp 1731220359
transform 1 0 2856 0 1 92
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5226_6
timestamp 1731220359
transform 1 0 2752 0 1 92
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5225_6
timestamp 1731220359
transform 1 0 2648 0 1 92
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5224_6
timestamp 1731220359
transform 1 0 2488 0 -1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5223_6
timestamp 1731220359
transform 1 0 2696 0 -1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5222_6
timestamp 1731220359
transform 1 0 2896 0 -1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5221_6
timestamp 1731220359
transform 1 0 3112 0 1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5220_6
timestamp 1731220359
transform 1 0 2952 0 1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5219_6
timestamp 1731220359
transform 1 0 2792 0 1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5218_6
timestamp 1731220359
transform 1 0 2632 0 1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5217_6
timestamp 1731220359
transform 1 0 2488 0 1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5216_6
timestamp 1731220359
transform 1 0 2952 0 -1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5215_6
timestamp 1731220359
transform 1 0 2792 0 -1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5214_6
timestamp 1731220359
transform 1 0 2632 0 -1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5213_6
timestamp 1731220359
transform 1 0 2480 0 -1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5212_6
timestamp 1731220359
transform 1 0 2336 0 -1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5211_6
timestamp 1731220359
transform 1 0 2768 0 1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5210_6
timestamp 1731220359
transform 1 0 2608 0 1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5209_6
timestamp 1731220359
transform 1 0 2456 0 1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5208_6
timestamp 1731220359
transform 1 0 2312 0 1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5207_6
timestamp 1731220359
transform 1 0 2176 0 1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5206_6
timestamp 1731220359
transform 1 0 2680 0 -1 576
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5205_6
timestamp 1731220359
transform 1 0 2496 0 -1 576
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5204_6
timestamp 1731220359
transform 1 0 2328 0 -1 576
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5203_6
timestamp 1731220359
transform 1 0 2176 0 -1 576
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5202_6
timestamp 1731220359
transform 1 0 2064 0 -1 576
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5201_6
timestamp 1731220359
transform 1 0 2104 0 1 580
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5200_6
timestamp 1731220359
transform 1 0 2240 0 1 580
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5199_6
timestamp 1731220359
transform 1 0 2392 0 1 580
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5198_6
timestamp 1731220359
transform 1 0 2752 0 1 580
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5197_6
timestamp 1731220359
transform 1 0 2568 0 1 580
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5196_6
timestamp 1731220359
transform 1 0 2488 0 -1 740
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5195_6
timestamp 1731220359
transform 1 0 2368 0 -1 740
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5194_6
timestamp 1731220359
transform 1 0 2616 0 -1 740
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5193_6
timestamp 1731220359
transform 1 0 2904 0 -1 740
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5192_6
timestamp 1731220359
transform 1 0 2760 0 -1 740
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5191_6
timestamp 1731220359
transform 1 0 2728 0 1 744
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5190_6
timestamp 1731220359
transform 1 0 2576 0 1 744
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5189_6
timestamp 1731220359
transform 1 0 2440 0 1 744
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5188_6
timestamp 1731220359
transform 1 0 2320 0 1 744
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5187_6
timestamp 1731220359
transform 1 0 2208 0 1 744
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5186_6
timestamp 1731220359
transform 1 0 2456 0 -1 896
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5185_6
timestamp 1731220359
transform 1 0 2248 0 -1 896
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5184_6
timestamp 1731220359
transform 1 0 2064 0 -1 896
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5183_6
timestamp 1731220359
transform 1 0 1896 0 -1 920
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5182_6
timestamp 1731220359
transform 1 0 1744 0 -1 920
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5181_6
timestamp 1731220359
transform 1 0 1896 0 1 920
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5180_6
timestamp 1731220359
transform 1 0 1768 0 1 920
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5179_6
timestamp 1731220359
transform 1 0 1624 0 1 920
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5178_6
timestamp 1731220359
transform 1 0 1480 0 1 920
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5177_6
timestamp 1731220359
transform 1 0 1640 0 -1 1072
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5176_6
timestamp 1731220359
transform 1 0 1824 0 -1 1072
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5175_6
timestamp 1731220359
transform 1 0 1744 0 1 1080
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5174_6
timestamp 1731220359
transform 1 0 1560 0 1 1080
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5173_6
timestamp 1731220359
transform 1 0 1704 0 -1 1236
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5172_6
timestamp 1731220359
transform 1 0 1552 0 -1 1236
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5171_6
timestamp 1731220359
transform 1 0 1400 0 -1 1236
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5170_6
timestamp 1731220359
transform 1 0 1432 0 1 1236
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5169_6
timestamp 1731220359
transform 1 0 1552 0 1 1236
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5168_6
timestamp 1731220359
transform 1 0 1576 0 -1 1396
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5167_6
timestamp 1731220359
transform 1 0 1320 0 1 1236
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5166_6
timestamp 1731220359
transform 1 0 1208 0 1 1236
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5165_6
timestamp 1731220359
transform 1 0 1104 0 -1 1236
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5164_6
timestamp 1731220359
transform 1 0 1248 0 -1 1236
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5163_6
timestamp 1731220359
transform 1 0 1200 0 1 1080
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5162_6
timestamp 1731220359
transform 1 0 1376 0 1 1080
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5161_6
timestamp 1731220359
transform 1 0 1456 0 -1 1072
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5160_6
timestamp 1731220359
transform 1 0 1272 0 -1 1072
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5159_6
timestamp 1731220359
transform 1 0 1328 0 1 920
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5158_6
timestamp 1731220359
transform 1 0 1168 0 1 920
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5157_6
timestamp 1731220359
transform 1 0 1232 0 -1 920
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5156_6
timestamp 1731220359
transform 1 0 1408 0 -1 920
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5155_6
timestamp 1731220359
transform 1 0 1576 0 -1 920
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5154_6
timestamp 1731220359
transform 1 0 1528 0 1 768
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5153_6
timestamp 1731220359
transform 1 0 1352 0 1 768
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5152_6
timestamp 1731220359
transform 1 0 1712 0 1 768
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5151_6
timestamp 1731220359
transform 1 0 1592 0 -1 768
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5150_6
timestamp 1731220359
transform 1 0 1448 0 -1 768
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5149_6
timestamp 1731220359
transform 1 0 1304 0 -1 768
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5148_6
timestamp 1731220359
transform 1 0 1288 0 1 616
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5147_6
timestamp 1731220359
transform 1 0 1400 0 1 616
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5146_6
timestamp 1731220359
transform 1 0 1512 0 1 616
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5145_6
timestamp 1731220359
transform 1 0 1448 0 -1 616
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5144_6
timestamp 1731220359
transform 1 0 1352 0 -1 616
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5143_6
timestamp 1731220359
transform 1 0 1256 0 -1 616
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5142_6
timestamp 1731220359
transform 1 0 1160 0 -1 616
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5141_6
timestamp 1731220359
transform 1 0 1064 0 1 616
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5140_6
timestamp 1731220359
transform 1 0 1176 0 1 616
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5139_6
timestamp 1731220359
transform 1 0 1160 0 -1 768
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5138_6
timestamp 1731220359
transform 1 0 1016 0 -1 768
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5137_6
timestamp 1731220359
transform 1 0 1000 0 1 768
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5136_6
timestamp 1731220359
transform 1 0 1176 0 1 768
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5135_6
timestamp 1731220359
transform 1 0 1048 0 -1 920
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5134_6
timestamp 1731220359
transform 1 0 1000 0 1 920
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5133_6
timestamp 1731220359
transform 1 0 1088 0 -1 1072
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5132_6
timestamp 1731220359
transform 1 0 1024 0 1 1080
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5131_6
timestamp 1731220359
transform 1 0 1096 0 1 1236
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5130_6
timestamp 1731220359
transform 1 0 1416 0 -1 1396
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5129_6
timestamp 1731220359
transform 1 0 1256 0 -1 1396
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5128_6
timestamp 1731220359
transform 1 0 1112 0 -1 1396
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5127_6
timestamp 1731220359
transform 1 0 976 0 -1 1396
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5126_6
timestamp 1731220359
transform 1 0 1224 0 1 1396
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5125_6
timestamp 1731220359
transform 1 0 1000 0 1 1396
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5124_6
timestamp 1731220359
transform 1 0 848 0 -1 1396
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5123_6
timestamp 1731220359
transform 1 0 720 0 -1 1396
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5122_6
timestamp 1731220359
transform 1 0 592 0 -1 1396
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5121_6
timestamp 1731220359
transform 1 0 456 0 -1 1396
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5120_6
timestamp 1731220359
transform 1 0 984 0 1 1236
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5119_6
timestamp 1731220359
transform 1 0 872 0 1 1236
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5118_6
timestamp 1731220359
transform 1 0 760 0 1 1236
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5117_6
timestamp 1731220359
transform 1 0 648 0 1 1236
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5116_6
timestamp 1731220359
transform 1 0 544 0 1 1236
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5115_6
timestamp 1731220359
transform 1 0 952 0 -1 1236
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5114_6
timestamp 1731220359
transform 1 0 800 0 -1 1236
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5113_6
timestamp 1731220359
transform 1 0 656 0 -1 1236
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5112_6
timestamp 1731220359
transform 1 0 512 0 -1 1236
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5111_6
timestamp 1731220359
transform 1 0 384 0 -1 1236
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5110_6
timestamp 1731220359
transform 1 0 840 0 1 1080
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5109_6
timestamp 1731220359
transform 1 0 664 0 1 1080
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5108_6
timestamp 1731220359
transform 1 0 488 0 1 1080
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5107_6
timestamp 1731220359
transform 1 0 320 0 1 1080
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5106_6
timestamp 1731220359
transform 1 0 168 0 1 1080
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5105_6
timestamp 1731220359
transform 1 0 904 0 -1 1072
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5104_6
timestamp 1731220359
transform 1 0 720 0 -1 1072
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5103_6
timestamp 1731220359
transform 1 0 536 0 -1 1072
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5102_6
timestamp 1731220359
transform 1 0 368 0 -1 1072
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5101_6
timestamp 1731220359
transform 1 0 224 0 -1 1072
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5100_6
timestamp 1731220359
transform 1 0 128 0 -1 1072
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_599_6
timestamp 1731220359
transform 1 0 128 0 1 920
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_598_6
timestamp 1731220359
transform 1 0 264 0 1 920
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_597_6
timestamp 1731220359
transform 1 0 440 0 1 920
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_596_6
timestamp 1731220359
transform 1 0 624 0 1 920
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_595_6
timestamp 1731220359
transform 1 0 816 0 1 920
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_594_6
timestamp 1731220359
transform 1 0 848 0 -1 920
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_593_6
timestamp 1731220359
transform 1 0 648 0 -1 920
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_592_6
timestamp 1731220359
transform 1 0 448 0 -1 920
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_591_6
timestamp 1731220359
transform 1 0 264 0 -1 920
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_590_6
timestamp 1731220359
transform 1 0 128 0 -1 920
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_589_6
timestamp 1731220359
transform 1 0 208 0 1 768
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_588_6
timestamp 1731220359
transform 1 0 336 0 1 768
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_587_6
timestamp 1731220359
transform 1 0 488 0 1 768
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_586_6
timestamp 1731220359
transform 1 0 648 0 1 768
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_585_6
timestamp 1731220359
transform 1 0 824 0 1 768
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_584_6
timestamp 1731220359
transform 1 0 880 0 -1 768
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_583_6
timestamp 1731220359
transform 1 0 616 0 -1 768
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_582_6
timestamp 1731220359
transform 1 0 488 0 -1 768
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_581_6
timestamp 1731220359
transform 1 0 368 0 -1 768
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_580_6
timestamp 1731220359
transform 1 0 744 0 -1 768
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_579_6
timestamp 1731220359
transform 1 0 736 0 1 616
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_578_6
timestamp 1731220359
transform 1 0 624 0 1 616
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_577_6
timestamp 1731220359
transform 1 0 520 0 1 616
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_576_6
timestamp 1731220359
transform 1 0 848 0 1 616
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_575_6
timestamp 1731220359
transform 1 0 960 0 1 616
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_574_6
timestamp 1731220359
transform 1 0 872 0 -1 616
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_573_6
timestamp 1731220359
transform 1 0 776 0 -1 616
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_572_6
timestamp 1731220359
transform 1 0 680 0 -1 616
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_571_6
timestamp 1731220359
transform 1 0 968 0 -1 616
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_570_6
timestamp 1731220359
transform 1 0 1064 0 -1 616
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_569_6
timestamp 1731220359
transform 1 0 1336 0 1 444
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_568_6
timestamp 1731220359
transform 1 0 1528 0 1 444
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_567_6
timestamp 1731220359
transform 1 0 1432 0 1 444
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_566_6
timestamp 1731220359
transform 1 0 1424 0 -1 432
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_565_6
timestamp 1731220359
transform 1 0 1312 0 -1 432
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_564_6
timestamp 1731220359
transform 1 0 1344 0 1 276
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_563_6
timestamp 1731220359
transform 1 0 1488 0 1 276
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_562_6
timestamp 1731220359
transform 1 0 1632 0 1 276
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_561_6
timestamp 1731220359
transform 1 0 1504 0 -1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_560_6
timestamp 1731220359
transform 1 0 1640 0 -1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_559_6
timestamp 1731220359
transform 1 0 1776 0 -1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_558_6
timestamp 1731220359
transform 1 0 1896 0 -1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_557_6
timestamp 1731220359
transform 1 0 2064 0 -1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_556_6
timestamp 1731220359
transform 1 0 2264 0 -1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_555_6
timestamp 1731220359
transform 1 0 2544 0 1 92
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_554_6
timestamp 1731220359
transform 1 0 2448 0 1 92
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_553_6
timestamp 1731220359
transform 1 0 2352 0 1 92
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_552_6
timestamp 1731220359
transform 1 0 2256 0 1 92
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_551_6
timestamp 1731220359
transform 1 0 2160 0 1 92
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_550_6
timestamp 1731220359
transform 1 0 2064 0 1 92
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_549_6
timestamp 1731220359
transform 1 0 1896 0 1 88
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_548_6
timestamp 1731220359
transform 1 0 1800 0 1 88
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_547_6
timestamp 1731220359
transform 1 0 1696 0 1 88
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_546_6
timestamp 1731220359
transform 1 0 1584 0 1 88
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_545_6
timestamp 1731220359
transform 1 0 1480 0 1 88
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_544_6
timestamp 1731220359
transform 1 0 1376 0 1 88
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_543_6
timestamp 1731220359
transform 1 0 1264 0 1 88
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_542_6
timestamp 1731220359
transform 1 0 1144 0 1 88
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_541_6
timestamp 1731220359
transform 1 0 1024 0 1 88
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_540_6
timestamp 1731220359
transform 1 0 1040 0 -1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_539_6
timestamp 1731220359
transform 1 0 1360 0 -1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_538_6
timestamp 1731220359
transform 1 0 1208 0 -1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_537_6
timestamp 1731220359
transform 1 0 1200 0 1 276
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_536_6
timestamp 1731220359
transform 1 0 1056 0 1 276
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_535_6
timestamp 1731220359
transform 1 0 992 0 -1 432
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_534_6
timestamp 1731220359
transform 1 0 1096 0 -1 432
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_533_6
timestamp 1731220359
transform 1 0 1200 0 -1 432
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_532_6
timestamp 1731220359
transform 1 0 1240 0 1 444
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_531_6
timestamp 1731220359
transform 1 0 1144 0 1 444
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_530_6
timestamp 1731220359
transform 1 0 1048 0 1 444
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_529_6
timestamp 1731220359
transform 1 0 952 0 1 444
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_528_6
timestamp 1731220359
transform 1 0 856 0 1 444
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_527_6
timestamp 1731220359
transform 1 0 760 0 1 444
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_526_6
timestamp 1731220359
transform 1 0 664 0 1 444
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_525_6
timestamp 1731220359
transform 1 0 568 0 1 444
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_524_6
timestamp 1731220359
transform 1 0 472 0 1 444
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_523_6
timestamp 1731220359
transform 1 0 376 0 1 444
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_522_6
timestamp 1731220359
transform 1 0 888 0 -1 432
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_521_6
timestamp 1731220359
transform 1 0 784 0 -1 432
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_520_6
timestamp 1731220359
transform 1 0 680 0 -1 432
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_519_6
timestamp 1731220359
transform 1 0 576 0 -1 432
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_518_6
timestamp 1731220359
transform 1 0 480 0 -1 432
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_517_6
timestamp 1731220359
transform 1 0 912 0 1 276
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_516_6
timestamp 1731220359
transform 1 0 760 0 1 276
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_515_6
timestamp 1731220359
transform 1 0 608 0 1 276
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_514_6
timestamp 1731220359
transform 1 0 456 0 1 276
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_513_6
timestamp 1731220359
transform 1 0 320 0 1 276
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_512_6
timestamp 1731220359
transform 1 0 864 0 -1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_511_6
timestamp 1731220359
transform 1 0 680 0 -1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_510_6
timestamp 1731220359
transform 1 0 496 0 -1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_59_6
timestamp 1731220359
transform 1 0 320 0 -1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_58_6
timestamp 1731220359
transform 1 0 160 0 -1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_57_6
timestamp 1731220359
transform 1 0 896 0 1 88
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_56_6
timestamp 1731220359
transform 1 0 768 0 1 88
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_55_6
timestamp 1731220359
transform 1 0 640 0 1 88
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_54_6
timestamp 1731220359
transform 1 0 520 0 1 88
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_53_6
timestamp 1731220359
transform 1 0 416 0 1 88
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_52_6
timestamp 1731220359
transform 1 0 320 0 1 88
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_51_6
timestamp 1731220359
transform 1 0 224 0 1 88
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_50_6
timestamp 1731220359
transform 1 0 128 0 1 88
box 8 5 92 72
<< end >>
