magic
tech sky130l
timestamp 1731220306
<< checkpaint >>
rect -19 66 50 67
rect -19 64 59 66
rect -19 59 60 64
rect -24 -20 60 59
rect -24 -26 52 -20
rect -19 -28 47 -26
<< ndiffusion >>
rect 8 11 13 12
rect 8 8 9 11
rect 12 8 13 11
rect 8 6 13 8
rect 15 11 20 12
rect 15 8 16 11
rect 19 8 20 11
rect 15 6 20 8
<< ndc >>
rect 9 8 12 11
rect 16 8 19 11
<< ntransistor >>
rect 13 6 15 12
<< pdiffusion >>
rect 8 23 13 27
rect 8 20 9 23
rect 12 20 13 23
rect 8 19 13 20
rect 15 23 20 27
rect 15 20 16 23
rect 19 20 20 23
rect 15 19 20 20
<< pdc >>
rect 9 20 12 23
rect 16 20 19 23
<< ptransistor >>
rect 13 19 15 27
<< polysilicon >>
rect 13 34 18 35
rect 13 31 14 34
rect 17 31 18 34
rect 13 30 18 31
rect 13 27 15 30
rect 13 12 15 19
rect 13 4 15 6
<< pc >>
rect 14 31 17 34
<< m1 >>
rect 13 31 14 34
rect 17 32 27 34
rect 17 31 28 32
rect 24 28 28 31
rect 8 23 12 24
rect 16 23 19 24
rect 8 20 9 23
rect 12 20 13 23
rect 16 16 19 20
rect 16 13 28 16
rect 8 11 12 12
rect 16 11 19 13
rect 24 12 28 13
rect 8 8 9 11
rect 12 8 13 11
rect 16 7 19 8
<< m2c >>
rect 9 20 12 23
rect 9 8 12 11
<< m2 >>
rect 8 23 13 24
rect 8 20 9 23
rect 12 20 13 23
rect 8 19 13 20
rect 8 11 13 12
rect 8 8 9 11
rect 12 8 13 11
rect 8 7 13 8
<< labels >>
rlabel space 0 0 32 40 6 prboundary
rlabel ndiffusion 20 9 20 9 3 Y
rlabel pdiffusion 20 21 20 21 3 Y
rlabel ndiffusion 16 7 16 7 3 Y
rlabel ndiffusion 16 9 16 9 3 Y
rlabel ndiffusion 16 12 16 12 3 Y
rlabel pdiffusion 16 20 16 20 3 Y
rlabel pdiffusion 16 21 16 21 3 Y
rlabel pdiffusion 16 24 16 24 3 Y
rlabel polysilicon 14 5 14 5 3 A
rlabel ntransistor 14 7 14 7 3 A
rlabel polysilicon 14 13 14 13 3 A
rlabel ptransistor 14 20 14 20 3 A
rlabel polysilicon 14 28 14 28 3 A
rlabel polysilicon 14 31 14 31 3 A
rlabel polysilicon 14 35 14 35 3 A
rlabel ndiffusion 9 7 9 7 3 GND
rlabel m1 25 13 25 13 3 Y
port 1 e
rlabel m1 25 29 25 29 3 A
port 2 e
rlabel ndc 17 9 17 9 3 Y
port 1 e
rlabel m1 17 12 17 12 3 Y
port 1 e
rlabel m1 17 14 17 14 3 Y
port 1 e
rlabel m1 17 17 17 17 3 Y
port 1 e
rlabel pdc 17 21 17 21 3 Y
port 1 e
rlabel m1 17 24 17 24 3 Y
port 1 e
rlabel m1 18 32 18 32 3 A
port 2 e
rlabel m1 18 33 18 33 3 A
port 2 e
rlabel pc 15 32 15 32 3 A
port 2 e
rlabel m1 17 8 17 8 3 Y
port 1 e
rlabel m1 14 32 14 32 3 A
port 2 e
rlabel m2 13 9 13 9 3 GND
rlabel m2 13 21 13 21 3 Vdd
rlabel m2c 10 9 10 9 3 GND
rlabel m2c 10 21 10 21 3 Vdd
rlabel m2 9 8 9 8 3 GND
rlabel m2 9 9 9 9 3 GND
rlabel m2 9 12 9 12 3 GND
rlabel m2 9 20 9 20 3 Vdd
rlabel m2 9 21 9 21 3 Vdd
rlabel m2 9 24 9 24 3 Vdd
<< end >>
