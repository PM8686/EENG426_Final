magic
tech sky130l
timestamp 1731220528
<< m2 >>
rect 110 1704 116 1705
rect 110 1700 111 1704
rect 115 1700 116 1704
rect 1662 1704 1668 1705
rect 110 1699 116 1700
rect 254 1702 260 1703
rect 254 1698 255 1702
rect 259 1698 260 1702
rect 254 1697 260 1698
rect 286 1702 292 1703
rect 286 1698 287 1702
rect 291 1698 292 1702
rect 286 1697 292 1698
rect 318 1702 324 1703
rect 318 1698 319 1702
rect 323 1698 324 1702
rect 318 1697 324 1698
rect 358 1702 364 1703
rect 358 1698 359 1702
rect 363 1698 364 1702
rect 358 1697 364 1698
rect 406 1702 412 1703
rect 406 1698 407 1702
rect 411 1698 412 1702
rect 406 1697 412 1698
rect 454 1702 460 1703
rect 454 1698 455 1702
rect 459 1698 460 1702
rect 454 1697 460 1698
rect 502 1702 508 1703
rect 502 1698 503 1702
rect 507 1698 508 1702
rect 502 1697 508 1698
rect 550 1702 556 1703
rect 550 1698 551 1702
rect 555 1698 556 1702
rect 550 1697 556 1698
rect 606 1702 612 1703
rect 606 1698 607 1702
rect 611 1698 612 1702
rect 606 1697 612 1698
rect 662 1702 668 1703
rect 662 1698 663 1702
rect 667 1698 668 1702
rect 662 1697 668 1698
rect 726 1702 732 1703
rect 726 1698 727 1702
rect 731 1698 732 1702
rect 726 1697 732 1698
rect 782 1702 788 1703
rect 782 1698 783 1702
rect 787 1698 788 1702
rect 782 1697 788 1698
rect 838 1702 844 1703
rect 838 1698 839 1702
rect 843 1698 844 1702
rect 838 1697 844 1698
rect 894 1702 900 1703
rect 894 1698 895 1702
rect 899 1698 900 1702
rect 894 1697 900 1698
rect 950 1702 956 1703
rect 950 1698 951 1702
rect 955 1698 956 1702
rect 950 1697 956 1698
rect 1006 1702 1012 1703
rect 1006 1698 1007 1702
rect 1011 1698 1012 1702
rect 1006 1697 1012 1698
rect 1062 1702 1068 1703
rect 1062 1698 1063 1702
rect 1067 1698 1068 1702
rect 1062 1697 1068 1698
rect 1118 1702 1124 1703
rect 1118 1698 1119 1702
rect 1123 1698 1124 1702
rect 1118 1697 1124 1698
rect 1174 1702 1180 1703
rect 1174 1698 1175 1702
rect 1179 1698 1180 1702
rect 1174 1697 1180 1698
rect 1230 1702 1236 1703
rect 1230 1698 1231 1702
rect 1235 1698 1236 1702
rect 1230 1697 1236 1698
rect 1286 1702 1292 1703
rect 1286 1698 1287 1702
rect 1291 1698 1292 1702
rect 1286 1697 1292 1698
rect 1334 1702 1340 1703
rect 1334 1698 1335 1702
rect 1339 1698 1340 1702
rect 1334 1697 1340 1698
rect 1374 1702 1380 1703
rect 1374 1698 1375 1702
rect 1379 1698 1380 1702
rect 1374 1697 1380 1698
rect 1422 1702 1428 1703
rect 1422 1698 1423 1702
rect 1427 1698 1428 1702
rect 1422 1697 1428 1698
rect 1470 1702 1476 1703
rect 1470 1698 1471 1702
rect 1475 1698 1476 1702
rect 1470 1697 1476 1698
rect 1518 1702 1524 1703
rect 1518 1698 1519 1702
rect 1523 1698 1524 1702
rect 1662 1700 1663 1704
rect 1667 1700 1668 1704
rect 1662 1699 1668 1700
rect 1518 1697 1524 1698
rect 110 1687 116 1688
rect 110 1683 111 1687
rect 115 1683 116 1687
rect 1662 1687 1668 1688
rect 110 1682 116 1683
rect 254 1685 260 1686
rect 254 1681 255 1685
rect 259 1681 260 1685
rect 254 1680 260 1681
rect 286 1685 292 1686
rect 286 1681 287 1685
rect 291 1681 292 1685
rect 286 1680 292 1681
rect 318 1685 324 1686
rect 318 1681 319 1685
rect 323 1681 324 1685
rect 318 1680 324 1681
rect 358 1685 364 1686
rect 358 1681 359 1685
rect 363 1681 364 1685
rect 358 1680 364 1681
rect 406 1685 412 1686
rect 406 1681 407 1685
rect 411 1681 412 1685
rect 406 1680 412 1681
rect 454 1685 460 1686
rect 454 1681 455 1685
rect 459 1681 460 1685
rect 454 1680 460 1681
rect 502 1685 508 1686
rect 502 1681 503 1685
rect 507 1681 508 1685
rect 502 1680 508 1681
rect 550 1685 556 1686
rect 550 1681 551 1685
rect 555 1681 556 1685
rect 550 1680 556 1681
rect 606 1685 612 1686
rect 606 1681 607 1685
rect 611 1681 612 1685
rect 606 1680 612 1681
rect 662 1685 668 1686
rect 662 1681 663 1685
rect 667 1681 668 1685
rect 662 1680 668 1681
rect 726 1685 732 1686
rect 726 1681 727 1685
rect 731 1681 732 1685
rect 726 1680 732 1681
rect 782 1685 788 1686
rect 782 1681 783 1685
rect 787 1681 788 1685
rect 782 1680 788 1681
rect 838 1685 844 1686
rect 838 1681 839 1685
rect 843 1681 844 1685
rect 838 1680 844 1681
rect 894 1685 900 1686
rect 894 1681 895 1685
rect 899 1681 900 1685
rect 894 1680 900 1681
rect 950 1685 956 1686
rect 950 1681 951 1685
rect 955 1681 956 1685
rect 950 1680 956 1681
rect 1006 1685 1012 1686
rect 1006 1681 1007 1685
rect 1011 1681 1012 1685
rect 1006 1680 1012 1681
rect 1062 1685 1068 1686
rect 1062 1681 1063 1685
rect 1067 1681 1068 1685
rect 1062 1680 1068 1681
rect 1118 1685 1124 1686
rect 1118 1681 1119 1685
rect 1123 1681 1124 1685
rect 1118 1680 1124 1681
rect 1174 1685 1180 1686
rect 1174 1681 1175 1685
rect 1179 1681 1180 1685
rect 1174 1680 1180 1681
rect 1230 1685 1236 1686
rect 1230 1681 1231 1685
rect 1235 1681 1236 1685
rect 1230 1680 1236 1681
rect 1286 1685 1292 1686
rect 1286 1681 1287 1685
rect 1291 1681 1292 1685
rect 1286 1680 1292 1681
rect 1334 1685 1340 1686
rect 1334 1681 1335 1685
rect 1339 1681 1340 1685
rect 1334 1680 1340 1681
rect 1374 1685 1380 1686
rect 1374 1681 1375 1685
rect 1379 1681 1380 1685
rect 1374 1680 1380 1681
rect 1422 1685 1428 1686
rect 1422 1681 1423 1685
rect 1427 1681 1428 1685
rect 1422 1680 1428 1681
rect 1470 1685 1476 1686
rect 1470 1681 1471 1685
rect 1475 1681 1476 1685
rect 1470 1680 1476 1681
rect 1518 1685 1524 1686
rect 1518 1681 1519 1685
rect 1523 1681 1524 1685
rect 1662 1683 1663 1687
rect 1667 1683 1668 1687
rect 1662 1682 1668 1683
rect 1518 1680 1524 1681
rect 134 1671 140 1672
rect 110 1669 116 1670
rect 110 1665 111 1669
rect 115 1665 116 1669
rect 134 1667 135 1671
rect 139 1667 140 1671
rect 134 1666 140 1667
rect 166 1671 172 1672
rect 166 1667 167 1671
rect 171 1667 172 1671
rect 166 1666 172 1667
rect 214 1671 220 1672
rect 214 1667 215 1671
rect 219 1667 220 1671
rect 214 1666 220 1667
rect 278 1671 284 1672
rect 278 1667 279 1671
rect 283 1667 284 1671
rect 278 1666 284 1667
rect 342 1671 348 1672
rect 342 1667 343 1671
rect 347 1667 348 1671
rect 342 1666 348 1667
rect 414 1671 420 1672
rect 414 1667 415 1671
rect 419 1667 420 1671
rect 414 1666 420 1667
rect 486 1671 492 1672
rect 486 1667 487 1671
rect 491 1667 492 1671
rect 486 1666 492 1667
rect 558 1671 564 1672
rect 558 1667 559 1671
rect 563 1667 564 1671
rect 558 1666 564 1667
rect 630 1671 636 1672
rect 630 1667 631 1671
rect 635 1667 636 1671
rect 630 1666 636 1667
rect 710 1671 716 1672
rect 710 1667 711 1671
rect 715 1667 716 1671
rect 710 1666 716 1667
rect 790 1671 796 1672
rect 790 1667 791 1671
rect 795 1667 796 1671
rect 790 1666 796 1667
rect 870 1671 876 1672
rect 870 1667 871 1671
rect 875 1667 876 1671
rect 870 1666 876 1667
rect 950 1671 956 1672
rect 950 1667 951 1671
rect 955 1667 956 1671
rect 950 1666 956 1667
rect 1030 1671 1036 1672
rect 1030 1667 1031 1671
rect 1035 1667 1036 1671
rect 1030 1666 1036 1667
rect 1102 1671 1108 1672
rect 1102 1667 1103 1671
rect 1107 1667 1108 1671
rect 1102 1666 1108 1667
rect 1174 1671 1180 1672
rect 1174 1667 1175 1671
rect 1179 1667 1180 1671
rect 1174 1666 1180 1667
rect 1246 1671 1252 1672
rect 1246 1667 1247 1671
rect 1251 1667 1252 1671
rect 1246 1666 1252 1667
rect 1318 1671 1324 1672
rect 1318 1667 1319 1671
rect 1323 1667 1324 1671
rect 1318 1666 1324 1667
rect 1390 1671 1396 1672
rect 1390 1667 1391 1671
rect 1395 1667 1396 1671
rect 1390 1666 1396 1667
rect 1454 1671 1460 1672
rect 1454 1667 1455 1671
rect 1459 1667 1460 1671
rect 1454 1666 1460 1667
rect 1518 1671 1524 1672
rect 1518 1667 1519 1671
rect 1523 1667 1524 1671
rect 1518 1666 1524 1667
rect 1582 1671 1588 1672
rect 1582 1667 1583 1671
rect 1587 1667 1588 1671
rect 1582 1666 1588 1667
rect 1622 1671 1628 1672
rect 1622 1667 1623 1671
rect 1627 1667 1628 1671
rect 1622 1666 1628 1667
rect 1662 1669 1668 1670
rect 110 1664 116 1665
rect 1662 1665 1663 1669
rect 1667 1665 1668 1669
rect 1662 1664 1668 1665
rect 134 1654 140 1655
rect 110 1652 116 1653
rect 110 1648 111 1652
rect 115 1648 116 1652
rect 134 1650 135 1654
rect 139 1650 140 1654
rect 134 1649 140 1650
rect 166 1654 172 1655
rect 166 1650 167 1654
rect 171 1650 172 1654
rect 166 1649 172 1650
rect 214 1654 220 1655
rect 214 1650 215 1654
rect 219 1650 220 1654
rect 214 1649 220 1650
rect 278 1654 284 1655
rect 278 1650 279 1654
rect 283 1650 284 1654
rect 278 1649 284 1650
rect 342 1654 348 1655
rect 342 1650 343 1654
rect 347 1650 348 1654
rect 342 1649 348 1650
rect 414 1654 420 1655
rect 414 1650 415 1654
rect 419 1650 420 1654
rect 414 1649 420 1650
rect 486 1654 492 1655
rect 486 1650 487 1654
rect 491 1650 492 1654
rect 486 1649 492 1650
rect 558 1654 564 1655
rect 558 1650 559 1654
rect 563 1650 564 1654
rect 558 1649 564 1650
rect 630 1654 636 1655
rect 630 1650 631 1654
rect 635 1650 636 1654
rect 630 1649 636 1650
rect 710 1654 716 1655
rect 710 1650 711 1654
rect 715 1650 716 1654
rect 710 1649 716 1650
rect 790 1654 796 1655
rect 790 1650 791 1654
rect 795 1650 796 1654
rect 790 1649 796 1650
rect 870 1654 876 1655
rect 870 1650 871 1654
rect 875 1650 876 1654
rect 870 1649 876 1650
rect 950 1654 956 1655
rect 950 1650 951 1654
rect 955 1650 956 1654
rect 950 1649 956 1650
rect 1030 1654 1036 1655
rect 1030 1650 1031 1654
rect 1035 1650 1036 1654
rect 1030 1649 1036 1650
rect 1102 1654 1108 1655
rect 1102 1650 1103 1654
rect 1107 1650 1108 1654
rect 1102 1649 1108 1650
rect 1174 1654 1180 1655
rect 1174 1650 1175 1654
rect 1179 1650 1180 1654
rect 1174 1649 1180 1650
rect 1246 1654 1252 1655
rect 1246 1650 1247 1654
rect 1251 1650 1252 1654
rect 1246 1649 1252 1650
rect 1318 1654 1324 1655
rect 1318 1650 1319 1654
rect 1323 1650 1324 1654
rect 1318 1649 1324 1650
rect 1390 1654 1396 1655
rect 1390 1650 1391 1654
rect 1395 1650 1396 1654
rect 1390 1649 1396 1650
rect 1454 1654 1460 1655
rect 1454 1650 1455 1654
rect 1459 1650 1460 1654
rect 1454 1649 1460 1650
rect 1518 1654 1524 1655
rect 1518 1650 1519 1654
rect 1523 1650 1524 1654
rect 1518 1649 1524 1650
rect 1582 1654 1588 1655
rect 1582 1650 1583 1654
rect 1587 1650 1588 1654
rect 1582 1649 1588 1650
rect 1622 1654 1628 1655
rect 1622 1650 1623 1654
rect 1627 1650 1628 1654
rect 1622 1649 1628 1650
rect 1662 1652 1668 1653
rect 110 1647 116 1648
rect 1662 1648 1663 1652
rect 1667 1648 1668 1652
rect 1662 1647 1668 1648
rect 110 1624 116 1625
rect 110 1620 111 1624
rect 115 1620 116 1624
rect 1662 1624 1668 1625
rect 110 1619 116 1620
rect 134 1622 140 1623
rect 134 1618 135 1622
rect 139 1618 140 1622
rect 134 1617 140 1618
rect 182 1622 188 1623
rect 182 1618 183 1622
rect 187 1618 188 1622
rect 182 1617 188 1618
rect 246 1622 252 1623
rect 246 1618 247 1622
rect 251 1618 252 1622
rect 246 1617 252 1618
rect 302 1622 308 1623
rect 302 1618 303 1622
rect 307 1618 308 1622
rect 302 1617 308 1618
rect 358 1622 364 1623
rect 358 1618 359 1622
rect 363 1618 364 1622
rect 358 1617 364 1618
rect 414 1622 420 1623
rect 414 1618 415 1622
rect 419 1618 420 1622
rect 414 1617 420 1618
rect 470 1622 476 1623
rect 470 1618 471 1622
rect 475 1618 476 1622
rect 470 1617 476 1618
rect 534 1622 540 1623
rect 534 1618 535 1622
rect 539 1618 540 1622
rect 534 1617 540 1618
rect 598 1622 604 1623
rect 598 1618 599 1622
rect 603 1618 604 1622
rect 598 1617 604 1618
rect 662 1622 668 1623
rect 662 1618 663 1622
rect 667 1618 668 1622
rect 662 1617 668 1618
rect 726 1622 732 1623
rect 726 1618 727 1622
rect 731 1618 732 1622
rect 726 1617 732 1618
rect 798 1622 804 1623
rect 798 1618 799 1622
rect 803 1618 804 1622
rect 798 1617 804 1618
rect 870 1622 876 1623
rect 870 1618 871 1622
rect 875 1618 876 1622
rect 870 1617 876 1618
rect 942 1622 948 1623
rect 942 1618 943 1622
rect 947 1618 948 1622
rect 942 1617 948 1618
rect 1022 1622 1028 1623
rect 1022 1618 1023 1622
rect 1027 1618 1028 1622
rect 1022 1617 1028 1618
rect 1102 1622 1108 1623
rect 1102 1618 1103 1622
rect 1107 1618 1108 1622
rect 1102 1617 1108 1618
rect 1174 1622 1180 1623
rect 1174 1618 1175 1622
rect 1179 1618 1180 1622
rect 1174 1617 1180 1618
rect 1246 1622 1252 1623
rect 1246 1618 1247 1622
rect 1251 1618 1252 1622
rect 1246 1617 1252 1618
rect 1318 1622 1324 1623
rect 1318 1618 1319 1622
rect 1323 1618 1324 1622
rect 1318 1617 1324 1618
rect 1398 1622 1404 1623
rect 1398 1618 1399 1622
rect 1403 1618 1404 1622
rect 1398 1617 1404 1618
rect 1478 1622 1484 1623
rect 1478 1618 1479 1622
rect 1483 1618 1484 1622
rect 1478 1617 1484 1618
rect 1558 1622 1564 1623
rect 1558 1618 1559 1622
rect 1563 1618 1564 1622
rect 1558 1617 1564 1618
rect 1622 1622 1628 1623
rect 1622 1618 1623 1622
rect 1627 1618 1628 1622
rect 1662 1620 1663 1624
rect 1667 1620 1668 1624
rect 1662 1619 1668 1620
rect 1622 1617 1628 1618
rect 110 1607 116 1608
rect 110 1603 111 1607
rect 115 1603 116 1607
rect 1662 1607 1668 1608
rect 110 1602 116 1603
rect 134 1605 140 1606
rect 134 1601 135 1605
rect 139 1601 140 1605
rect 134 1600 140 1601
rect 182 1605 188 1606
rect 182 1601 183 1605
rect 187 1601 188 1605
rect 182 1600 188 1601
rect 246 1605 252 1606
rect 246 1601 247 1605
rect 251 1601 252 1605
rect 246 1600 252 1601
rect 302 1605 308 1606
rect 302 1601 303 1605
rect 307 1601 308 1605
rect 302 1600 308 1601
rect 358 1605 364 1606
rect 358 1601 359 1605
rect 363 1601 364 1605
rect 358 1600 364 1601
rect 414 1605 420 1606
rect 414 1601 415 1605
rect 419 1601 420 1605
rect 414 1600 420 1601
rect 470 1605 476 1606
rect 470 1601 471 1605
rect 475 1601 476 1605
rect 470 1600 476 1601
rect 534 1605 540 1606
rect 534 1601 535 1605
rect 539 1601 540 1605
rect 534 1600 540 1601
rect 598 1605 604 1606
rect 598 1601 599 1605
rect 603 1601 604 1605
rect 598 1600 604 1601
rect 662 1605 668 1606
rect 662 1601 663 1605
rect 667 1601 668 1605
rect 662 1600 668 1601
rect 726 1605 732 1606
rect 726 1601 727 1605
rect 731 1601 732 1605
rect 726 1600 732 1601
rect 798 1605 804 1606
rect 798 1601 799 1605
rect 803 1601 804 1605
rect 798 1600 804 1601
rect 870 1605 876 1606
rect 870 1601 871 1605
rect 875 1601 876 1605
rect 870 1600 876 1601
rect 942 1605 948 1606
rect 942 1601 943 1605
rect 947 1601 948 1605
rect 942 1600 948 1601
rect 1022 1605 1028 1606
rect 1022 1601 1023 1605
rect 1027 1601 1028 1605
rect 1022 1600 1028 1601
rect 1102 1605 1108 1606
rect 1102 1601 1103 1605
rect 1107 1601 1108 1605
rect 1102 1600 1108 1601
rect 1174 1605 1180 1606
rect 1174 1601 1175 1605
rect 1179 1601 1180 1605
rect 1174 1600 1180 1601
rect 1246 1605 1252 1606
rect 1246 1601 1247 1605
rect 1251 1601 1252 1605
rect 1246 1600 1252 1601
rect 1318 1605 1324 1606
rect 1318 1601 1319 1605
rect 1323 1601 1324 1605
rect 1318 1600 1324 1601
rect 1398 1605 1404 1606
rect 1398 1601 1399 1605
rect 1403 1601 1404 1605
rect 1398 1600 1404 1601
rect 1478 1605 1484 1606
rect 1478 1601 1479 1605
rect 1483 1601 1484 1605
rect 1478 1600 1484 1601
rect 1558 1605 1564 1606
rect 1558 1601 1559 1605
rect 1563 1601 1564 1605
rect 1558 1600 1564 1601
rect 1622 1605 1628 1606
rect 1622 1601 1623 1605
rect 1627 1601 1628 1605
rect 1662 1603 1663 1607
rect 1667 1603 1668 1607
rect 1662 1602 1668 1603
rect 1622 1600 1628 1601
rect 134 1591 140 1592
rect 110 1589 116 1590
rect 110 1585 111 1589
rect 115 1585 116 1589
rect 134 1587 135 1591
rect 139 1587 140 1591
rect 134 1586 140 1587
rect 166 1591 172 1592
rect 166 1587 167 1591
rect 171 1587 172 1591
rect 166 1586 172 1587
rect 222 1591 228 1592
rect 222 1587 223 1591
rect 227 1587 228 1591
rect 222 1586 228 1587
rect 278 1591 284 1592
rect 278 1587 279 1591
rect 283 1587 284 1591
rect 278 1586 284 1587
rect 334 1591 340 1592
rect 334 1587 335 1591
rect 339 1587 340 1591
rect 334 1586 340 1587
rect 382 1591 388 1592
rect 382 1587 383 1591
rect 387 1587 388 1591
rect 382 1586 388 1587
rect 430 1591 436 1592
rect 430 1587 431 1591
rect 435 1587 436 1591
rect 430 1586 436 1587
rect 478 1591 484 1592
rect 478 1587 479 1591
rect 483 1587 484 1591
rect 478 1586 484 1587
rect 534 1591 540 1592
rect 534 1587 535 1591
rect 539 1587 540 1591
rect 534 1586 540 1587
rect 598 1591 604 1592
rect 598 1587 599 1591
rect 603 1587 604 1591
rect 598 1586 604 1587
rect 662 1591 668 1592
rect 662 1587 663 1591
rect 667 1587 668 1591
rect 662 1586 668 1587
rect 726 1591 732 1592
rect 726 1587 727 1591
rect 731 1587 732 1591
rect 726 1586 732 1587
rect 798 1591 804 1592
rect 798 1587 799 1591
rect 803 1587 804 1591
rect 798 1586 804 1587
rect 870 1591 876 1592
rect 870 1587 871 1591
rect 875 1587 876 1591
rect 870 1586 876 1587
rect 950 1591 956 1592
rect 950 1587 951 1591
rect 955 1587 956 1591
rect 950 1586 956 1587
rect 1038 1591 1044 1592
rect 1038 1587 1039 1591
rect 1043 1587 1044 1591
rect 1038 1586 1044 1587
rect 1118 1591 1124 1592
rect 1118 1587 1119 1591
rect 1123 1587 1124 1591
rect 1118 1586 1124 1587
rect 1198 1591 1204 1592
rect 1198 1587 1199 1591
rect 1203 1587 1204 1591
rect 1198 1586 1204 1587
rect 1278 1591 1284 1592
rect 1278 1587 1279 1591
rect 1283 1587 1284 1591
rect 1278 1586 1284 1587
rect 1350 1591 1356 1592
rect 1350 1587 1351 1591
rect 1355 1587 1356 1591
rect 1350 1586 1356 1587
rect 1414 1591 1420 1592
rect 1414 1587 1415 1591
rect 1419 1587 1420 1591
rect 1414 1586 1420 1587
rect 1470 1591 1476 1592
rect 1470 1587 1471 1591
rect 1475 1587 1476 1591
rect 1470 1586 1476 1587
rect 1526 1591 1532 1592
rect 1526 1587 1527 1591
rect 1531 1587 1532 1591
rect 1526 1586 1532 1587
rect 1582 1591 1588 1592
rect 1582 1587 1583 1591
rect 1587 1587 1588 1591
rect 1582 1586 1588 1587
rect 1622 1591 1628 1592
rect 1622 1587 1623 1591
rect 1627 1587 1628 1591
rect 1622 1586 1628 1587
rect 1662 1589 1668 1590
rect 110 1584 116 1585
rect 1662 1585 1663 1589
rect 1667 1585 1668 1589
rect 1662 1584 1668 1585
rect 134 1574 140 1575
rect 110 1572 116 1573
rect 110 1568 111 1572
rect 115 1568 116 1572
rect 134 1570 135 1574
rect 139 1570 140 1574
rect 134 1569 140 1570
rect 166 1574 172 1575
rect 166 1570 167 1574
rect 171 1570 172 1574
rect 166 1569 172 1570
rect 222 1574 228 1575
rect 222 1570 223 1574
rect 227 1570 228 1574
rect 222 1569 228 1570
rect 278 1574 284 1575
rect 278 1570 279 1574
rect 283 1570 284 1574
rect 278 1569 284 1570
rect 334 1574 340 1575
rect 334 1570 335 1574
rect 339 1570 340 1574
rect 334 1569 340 1570
rect 382 1574 388 1575
rect 382 1570 383 1574
rect 387 1570 388 1574
rect 382 1569 388 1570
rect 430 1574 436 1575
rect 430 1570 431 1574
rect 435 1570 436 1574
rect 430 1569 436 1570
rect 478 1574 484 1575
rect 478 1570 479 1574
rect 483 1570 484 1574
rect 478 1569 484 1570
rect 534 1574 540 1575
rect 534 1570 535 1574
rect 539 1570 540 1574
rect 534 1569 540 1570
rect 598 1574 604 1575
rect 598 1570 599 1574
rect 603 1570 604 1574
rect 598 1569 604 1570
rect 662 1574 668 1575
rect 662 1570 663 1574
rect 667 1570 668 1574
rect 662 1569 668 1570
rect 726 1574 732 1575
rect 726 1570 727 1574
rect 731 1570 732 1574
rect 726 1569 732 1570
rect 798 1574 804 1575
rect 798 1570 799 1574
rect 803 1570 804 1574
rect 798 1569 804 1570
rect 870 1574 876 1575
rect 870 1570 871 1574
rect 875 1570 876 1574
rect 870 1569 876 1570
rect 950 1574 956 1575
rect 950 1570 951 1574
rect 955 1570 956 1574
rect 950 1569 956 1570
rect 1038 1574 1044 1575
rect 1038 1570 1039 1574
rect 1043 1570 1044 1574
rect 1038 1569 1044 1570
rect 1118 1574 1124 1575
rect 1118 1570 1119 1574
rect 1123 1570 1124 1574
rect 1118 1569 1124 1570
rect 1198 1574 1204 1575
rect 1198 1570 1199 1574
rect 1203 1570 1204 1574
rect 1198 1569 1204 1570
rect 1278 1574 1284 1575
rect 1278 1570 1279 1574
rect 1283 1570 1284 1574
rect 1278 1569 1284 1570
rect 1350 1574 1356 1575
rect 1350 1570 1351 1574
rect 1355 1570 1356 1574
rect 1350 1569 1356 1570
rect 1414 1574 1420 1575
rect 1414 1570 1415 1574
rect 1419 1570 1420 1574
rect 1414 1569 1420 1570
rect 1470 1574 1476 1575
rect 1470 1570 1471 1574
rect 1475 1570 1476 1574
rect 1470 1569 1476 1570
rect 1526 1574 1532 1575
rect 1526 1570 1527 1574
rect 1531 1570 1532 1574
rect 1526 1569 1532 1570
rect 1582 1574 1588 1575
rect 1582 1570 1583 1574
rect 1587 1570 1588 1574
rect 1582 1569 1588 1570
rect 1622 1574 1628 1575
rect 1622 1570 1623 1574
rect 1627 1570 1628 1574
rect 1622 1569 1628 1570
rect 1662 1572 1668 1573
rect 110 1567 116 1568
rect 1662 1568 1663 1572
rect 1667 1568 1668 1572
rect 1662 1567 1668 1568
rect 110 1544 116 1545
rect 110 1540 111 1544
rect 115 1540 116 1544
rect 1662 1544 1668 1545
rect 110 1539 116 1540
rect 134 1542 140 1543
rect 134 1538 135 1542
rect 139 1538 140 1542
rect 134 1537 140 1538
rect 166 1542 172 1543
rect 166 1538 167 1542
rect 171 1538 172 1542
rect 166 1537 172 1538
rect 214 1542 220 1543
rect 214 1538 215 1542
rect 219 1538 220 1542
rect 214 1537 220 1538
rect 262 1542 268 1543
rect 262 1538 263 1542
rect 267 1538 268 1542
rect 262 1537 268 1538
rect 310 1542 316 1543
rect 310 1538 311 1542
rect 315 1538 316 1542
rect 310 1537 316 1538
rect 358 1542 364 1543
rect 358 1538 359 1542
rect 363 1538 364 1542
rect 358 1537 364 1538
rect 406 1542 412 1543
rect 406 1538 407 1542
rect 411 1538 412 1542
rect 406 1537 412 1538
rect 454 1542 460 1543
rect 454 1538 455 1542
rect 459 1538 460 1542
rect 454 1537 460 1538
rect 510 1542 516 1543
rect 510 1538 511 1542
rect 515 1538 516 1542
rect 510 1537 516 1538
rect 566 1542 572 1543
rect 566 1538 567 1542
rect 571 1538 572 1542
rect 566 1537 572 1538
rect 630 1542 636 1543
rect 630 1538 631 1542
rect 635 1538 636 1542
rect 630 1537 636 1538
rect 694 1542 700 1543
rect 694 1538 695 1542
rect 699 1538 700 1542
rect 694 1537 700 1538
rect 758 1542 764 1543
rect 758 1538 759 1542
rect 763 1538 764 1542
rect 758 1537 764 1538
rect 830 1542 836 1543
rect 830 1538 831 1542
rect 835 1538 836 1542
rect 830 1537 836 1538
rect 918 1542 924 1543
rect 918 1538 919 1542
rect 923 1538 924 1542
rect 918 1537 924 1538
rect 1006 1542 1012 1543
rect 1006 1538 1007 1542
rect 1011 1538 1012 1542
rect 1006 1537 1012 1538
rect 1094 1542 1100 1543
rect 1094 1538 1095 1542
rect 1099 1538 1100 1542
rect 1094 1537 1100 1538
rect 1182 1542 1188 1543
rect 1182 1538 1183 1542
rect 1187 1538 1188 1542
rect 1182 1537 1188 1538
rect 1262 1542 1268 1543
rect 1262 1538 1263 1542
rect 1267 1538 1268 1542
rect 1262 1537 1268 1538
rect 1334 1542 1340 1543
rect 1334 1538 1335 1542
rect 1339 1538 1340 1542
rect 1334 1537 1340 1538
rect 1406 1542 1412 1543
rect 1406 1538 1407 1542
rect 1411 1538 1412 1542
rect 1406 1537 1412 1538
rect 1470 1542 1476 1543
rect 1470 1538 1471 1542
rect 1475 1538 1476 1542
rect 1470 1537 1476 1538
rect 1526 1542 1532 1543
rect 1526 1538 1527 1542
rect 1531 1538 1532 1542
rect 1526 1537 1532 1538
rect 1582 1542 1588 1543
rect 1582 1538 1583 1542
rect 1587 1538 1588 1542
rect 1582 1537 1588 1538
rect 1622 1542 1628 1543
rect 1622 1538 1623 1542
rect 1627 1538 1628 1542
rect 1662 1540 1663 1544
rect 1667 1540 1668 1544
rect 1662 1539 1668 1540
rect 1622 1537 1628 1538
rect 110 1527 116 1528
rect 110 1523 111 1527
rect 115 1523 116 1527
rect 1662 1527 1668 1528
rect 110 1522 116 1523
rect 134 1525 140 1526
rect 134 1521 135 1525
rect 139 1521 140 1525
rect 134 1520 140 1521
rect 166 1525 172 1526
rect 166 1521 167 1525
rect 171 1521 172 1525
rect 166 1520 172 1521
rect 214 1525 220 1526
rect 214 1521 215 1525
rect 219 1521 220 1525
rect 214 1520 220 1521
rect 262 1525 268 1526
rect 262 1521 263 1525
rect 267 1521 268 1525
rect 262 1520 268 1521
rect 310 1525 316 1526
rect 310 1521 311 1525
rect 315 1521 316 1525
rect 310 1520 316 1521
rect 358 1525 364 1526
rect 358 1521 359 1525
rect 363 1521 364 1525
rect 358 1520 364 1521
rect 406 1525 412 1526
rect 406 1521 407 1525
rect 411 1521 412 1525
rect 406 1520 412 1521
rect 454 1525 460 1526
rect 454 1521 455 1525
rect 459 1521 460 1525
rect 454 1520 460 1521
rect 510 1525 516 1526
rect 510 1521 511 1525
rect 515 1521 516 1525
rect 510 1520 516 1521
rect 566 1525 572 1526
rect 566 1521 567 1525
rect 571 1521 572 1525
rect 566 1520 572 1521
rect 630 1525 636 1526
rect 630 1521 631 1525
rect 635 1521 636 1525
rect 630 1520 636 1521
rect 694 1525 700 1526
rect 694 1521 695 1525
rect 699 1521 700 1525
rect 694 1520 700 1521
rect 758 1525 764 1526
rect 758 1521 759 1525
rect 763 1521 764 1525
rect 758 1520 764 1521
rect 830 1525 836 1526
rect 830 1521 831 1525
rect 835 1521 836 1525
rect 830 1520 836 1521
rect 918 1525 924 1526
rect 918 1521 919 1525
rect 923 1521 924 1525
rect 918 1520 924 1521
rect 1006 1525 1012 1526
rect 1006 1521 1007 1525
rect 1011 1521 1012 1525
rect 1006 1520 1012 1521
rect 1094 1525 1100 1526
rect 1094 1521 1095 1525
rect 1099 1521 1100 1525
rect 1094 1520 1100 1521
rect 1182 1525 1188 1526
rect 1182 1521 1183 1525
rect 1187 1521 1188 1525
rect 1182 1520 1188 1521
rect 1262 1525 1268 1526
rect 1262 1521 1263 1525
rect 1267 1521 1268 1525
rect 1262 1520 1268 1521
rect 1334 1525 1340 1526
rect 1334 1521 1335 1525
rect 1339 1521 1340 1525
rect 1334 1520 1340 1521
rect 1406 1525 1412 1526
rect 1406 1521 1407 1525
rect 1411 1521 1412 1525
rect 1406 1520 1412 1521
rect 1470 1525 1476 1526
rect 1470 1521 1471 1525
rect 1475 1521 1476 1525
rect 1470 1520 1476 1521
rect 1526 1525 1532 1526
rect 1526 1521 1527 1525
rect 1531 1521 1532 1525
rect 1526 1520 1532 1521
rect 1582 1525 1588 1526
rect 1582 1521 1583 1525
rect 1587 1521 1588 1525
rect 1582 1520 1588 1521
rect 1622 1525 1628 1526
rect 1622 1521 1623 1525
rect 1627 1521 1628 1525
rect 1662 1523 1663 1527
rect 1667 1523 1668 1527
rect 1662 1522 1668 1523
rect 1622 1520 1628 1521
rect 134 1507 140 1508
rect 110 1505 116 1506
rect 110 1501 111 1505
rect 115 1501 116 1505
rect 134 1503 135 1507
rect 139 1503 140 1507
rect 134 1502 140 1503
rect 166 1507 172 1508
rect 166 1503 167 1507
rect 171 1503 172 1507
rect 166 1502 172 1503
rect 222 1507 228 1508
rect 222 1503 223 1507
rect 227 1503 228 1507
rect 222 1502 228 1503
rect 294 1507 300 1508
rect 294 1503 295 1507
rect 299 1503 300 1507
rect 294 1502 300 1503
rect 374 1507 380 1508
rect 374 1503 375 1507
rect 379 1503 380 1507
rect 374 1502 380 1503
rect 454 1507 460 1508
rect 454 1503 455 1507
rect 459 1503 460 1507
rect 454 1502 460 1503
rect 526 1507 532 1508
rect 526 1503 527 1507
rect 531 1503 532 1507
rect 526 1502 532 1503
rect 598 1507 604 1508
rect 598 1503 599 1507
rect 603 1503 604 1507
rect 598 1502 604 1503
rect 670 1507 676 1508
rect 670 1503 671 1507
rect 675 1503 676 1507
rect 670 1502 676 1503
rect 742 1507 748 1508
rect 742 1503 743 1507
rect 747 1503 748 1507
rect 742 1502 748 1503
rect 814 1507 820 1508
rect 814 1503 815 1507
rect 819 1503 820 1507
rect 814 1502 820 1503
rect 878 1507 884 1508
rect 878 1503 879 1507
rect 883 1503 884 1507
rect 878 1502 884 1503
rect 942 1507 948 1508
rect 942 1503 943 1507
rect 947 1503 948 1507
rect 942 1502 948 1503
rect 1006 1507 1012 1508
rect 1006 1503 1007 1507
rect 1011 1503 1012 1507
rect 1006 1502 1012 1503
rect 1062 1507 1068 1508
rect 1062 1503 1063 1507
rect 1067 1503 1068 1507
rect 1062 1502 1068 1503
rect 1110 1507 1116 1508
rect 1110 1503 1111 1507
rect 1115 1503 1116 1507
rect 1110 1502 1116 1503
rect 1150 1507 1156 1508
rect 1150 1503 1151 1507
rect 1155 1503 1156 1507
rect 1150 1502 1156 1503
rect 1182 1507 1188 1508
rect 1182 1503 1183 1507
rect 1187 1503 1188 1507
rect 1182 1502 1188 1503
rect 1214 1507 1220 1508
rect 1214 1503 1215 1507
rect 1219 1503 1220 1507
rect 1214 1502 1220 1503
rect 1254 1507 1260 1508
rect 1254 1503 1255 1507
rect 1259 1503 1260 1507
rect 1254 1502 1260 1503
rect 1294 1507 1300 1508
rect 1294 1503 1295 1507
rect 1299 1503 1300 1507
rect 1294 1502 1300 1503
rect 1350 1507 1356 1508
rect 1350 1503 1351 1507
rect 1355 1503 1356 1507
rect 1350 1502 1356 1503
rect 1414 1507 1420 1508
rect 1414 1503 1415 1507
rect 1419 1503 1420 1507
rect 1414 1502 1420 1503
rect 1486 1507 1492 1508
rect 1486 1503 1487 1507
rect 1491 1503 1492 1507
rect 1486 1502 1492 1503
rect 1566 1507 1572 1508
rect 1566 1503 1567 1507
rect 1571 1503 1572 1507
rect 1566 1502 1572 1503
rect 1622 1507 1628 1508
rect 1622 1503 1623 1507
rect 1627 1503 1628 1507
rect 1622 1502 1628 1503
rect 1662 1505 1668 1506
rect 110 1500 116 1501
rect 1662 1501 1663 1505
rect 1667 1501 1668 1505
rect 1662 1500 1668 1501
rect 134 1490 140 1491
rect 110 1488 116 1489
rect 110 1484 111 1488
rect 115 1484 116 1488
rect 134 1486 135 1490
rect 139 1486 140 1490
rect 134 1485 140 1486
rect 166 1490 172 1491
rect 166 1486 167 1490
rect 171 1486 172 1490
rect 166 1485 172 1486
rect 222 1490 228 1491
rect 222 1486 223 1490
rect 227 1486 228 1490
rect 222 1485 228 1486
rect 294 1490 300 1491
rect 294 1486 295 1490
rect 299 1486 300 1490
rect 294 1485 300 1486
rect 374 1490 380 1491
rect 374 1486 375 1490
rect 379 1486 380 1490
rect 374 1485 380 1486
rect 454 1490 460 1491
rect 454 1486 455 1490
rect 459 1486 460 1490
rect 454 1485 460 1486
rect 526 1490 532 1491
rect 526 1486 527 1490
rect 531 1486 532 1490
rect 526 1485 532 1486
rect 598 1490 604 1491
rect 598 1486 599 1490
rect 603 1486 604 1490
rect 598 1485 604 1486
rect 670 1490 676 1491
rect 670 1486 671 1490
rect 675 1486 676 1490
rect 670 1485 676 1486
rect 742 1490 748 1491
rect 742 1486 743 1490
rect 747 1486 748 1490
rect 742 1485 748 1486
rect 814 1490 820 1491
rect 814 1486 815 1490
rect 819 1486 820 1490
rect 814 1485 820 1486
rect 878 1490 884 1491
rect 878 1486 879 1490
rect 883 1486 884 1490
rect 878 1485 884 1486
rect 942 1490 948 1491
rect 942 1486 943 1490
rect 947 1486 948 1490
rect 942 1485 948 1486
rect 1006 1490 1012 1491
rect 1006 1486 1007 1490
rect 1011 1486 1012 1490
rect 1006 1485 1012 1486
rect 1062 1490 1068 1491
rect 1062 1486 1063 1490
rect 1067 1486 1068 1490
rect 1062 1485 1068 1486
rect 1110 1490 1116 1491
rect 1110 1486 1111 1490
rect 1115 1486 1116 1490
rect 1110 1485 1116 1486
rect 1150 1490 1156 1491
rect 1150 1486 1151 1490
rect 1155 1486 1156 1490
rect 1150 1485 1156 1486
rect 1182 1490 1188 1491
rect 1182 1486 1183 1490
rect 1187 1486 1188 1490
rect 1182 1485 1188 1486
rect 1214 1490 1220 1491
rect 1214 1486 1215 1490
rect 1219 1486 1220 1490
rect 1214 1485 1220 1486
rect 1254 1490 1260 1491
rect 1254 1486 1255 1490
rect 1259 1486 1260 1490
rect 1254 1485 1260 1486
rect 1294 1490 1300 1491
rect 1294 1486 1295 1490
rect 1299 1486 1300 1490
rect 1294 1485 1300 1486
rect 1350 1490 1356 1491
rect 1350 1486 1351 1490
rect 1355 1486 1356 1490
rect 1350 1485 1356 1486
rect 1414 1490 1420 1491
rect 1414 1486 1415 1490
rect 1419 1486 1420 1490
rect 1414 1485 1420 1486
rect 1486 1490 1492 1491
rect 1486 1486 1487 1490
rect 1491 1486 1492 1490
rect 1486 1485 1492 1486
rect 1566 1490 1572 1491
rect 1566 1486 1567 1490
rect 1571 1486 1572 1490
rect 1566 1485 1572 1486
rect 1622 1490 1628 1491
rect 1622 1486 1623 1490
rect 1627 1486 1628 1490
rect 1622 1485 1628 1486
rect 1662 1488 1668 1489
rect 110 1483 116 1484
rect 1662 1484 1663 1488
rect 1667 1484 1668 1488
rect 1662 1483 1668 1484
rect 110 1460 116 1461
rect 110 1456 111 1460
rect 115 1456 116 1460
rect 1662 1460 1668 1461
rect 110 1455 116 1456
rect 134 1458 140 1459
rect 134 1454 135 1458
rect 139 1454 140 1458
rect 134 1453 140 1454
rect 166 1458 172 1459
rect 166 1454 167 1458
rect 171 1454 172 1458
rect 166 1453 172 1454
rect 222 1458 228 1459
rect 222 1454 223 1458
rect 227 1454 228 1458
rect 222 1453 228 1454
rect 294 1458 300 1459
rect 294 1454 295 1458
rect 299 1454 300 1458
rect 294 1453 300 1454
rect 374 1458 380 1459
rect 374 1454 375 1458
rect 379 1454 380 1458
rect 374 1453 380 1454
rect 454 1458 460 1459
rect 454 1454 455 1458
rect 459 1454 460 1458
rect 454 1453 460 1454
rect 526 1458 532 1459
rect 526 1454 527 1458
rect 531 1454 532 1458
rect 526 1453 532 1454
rect 598 1458 604 1459
rect 598 1454 599 1458
rect 603 1454 604 1458
rect 598 1453 604 1454
rect 662 1458 668 1459
rect 662 1454 663 1458
rect 667 1454 668 1458
rect 662 1453 668 1454
rect 718 1458 724 1459
rect 718 1454 719 1458
rect 723 1454 724 1458
rect 718 1453 724 1454
rect 782 1458 788 1459
rect 782 1454 783 1458
rect 787 1454 788 1458
rect 782 1453 788 1454
rect 846 1458 852 1459
rect 846 1454 847 1458
rect 851 1454 852 1458
rect 846 1453 852 1454
rect 902 1458 908 1459
rect 902 1454 903 1458
rect 907 1454 908 1458
rect 902 1453 908 1454
rect 958 1458 964 1459
rect 958 1454 959 1458
rect 963 1454 964 1458
rect 958 1453 964 1454
rect 1014 1458 1020 1459
rect 1014 1454 1015 1458
rect 1019 1454 1020 1458
rect 1014 1453 1020 1454
rect 1070 1458 1076 1459
rect 1070 1454 1071 1458
rect 1075 1454 1076 1458
rect 1070 1453 1076 1454
rect 1118 1458 1124 1459
rect 1118 1454 1119 1458
rect 1123 1454 1124 1458
rect 1118 1453 1124 1454
rect 1158 1458 1164 1459
rect 1158 1454 1159 1458
rect 1163 1454 1164 1458
rect 1158 1453 1164 1454
rect 1206 1458 1212 1459
rect 1206 1454 1207 1458
rect 1211 1454 1212 1458
rect 1206 1453 1212 1454
rect 1262 1458 1268 1459
rect 1262 1454 1263 1458
rect 1267 1454 1268 1458
rect 1262 1453 1268 1454
rect 1326 1458 1332 1459
rect 1326 1454 1327 1458
rect 1331 1454 1332 1458
rect 1326 1453 1332 1454
rect 1398 1458 1404 1459
rect 1398 1454 1399 1458
rect 1403 1454 1404 1458
rect 1398 1453 1404 1454
rect 1478 1458 1484 1459
rect 1478 1454 1479 1458
rect 1483 1454 1484 1458
rect 1478 1453 1484 1454
rect 1558 1458 1564 1459
rect 1558 1454 1559 1458
rect 1563 1454 1564 1458
rect 1558 1453 1564 1454
rect 1622 1458 1628 1459
rect 1622 1454 1623 1458
rect 1627 1454 1628 1458
rect 1662 1456 1663 1460
rect 1667 1456 1668 1460
rect 1662 1455 1668 1456
rect 1622 1453 1628 1454
rect 110 1443 116 1444
rect 110 1439 111 1443
rect 115 1439 116 1443
rect 1662 1443 1668 1444
rect 110 1438 116 1439
rect 134 1441 140 1442
rect 134 1437 135 1441
rect 139 1437 140 1441
rect 134 1436 140 1437
rect 166 1441 172 1442
rect 166 1437 167 1441
rect 171 1437 172 1441
rect 166 1436 172 1437
rect 222 1441 228 1442
rect 222 1437 223 1441
rect 227 1437 228 1441
rect 222 1436 228 1437
rect 294 1441 300 1442
rect 294 1437 295 1441
rect 299 1437 300 1441
rect 294 1436 300 1437
rect 374 1441 380 1442
rect 374 1437 375 1441
rect 379 1437 380 1441
rect 374 1436 380 1437
rect 454 1441 460 1442
rect 454 1437 455 1441
rect 459 1437 460 1441
rect 454 1436 460 1437
rect 526 1441 532 1442
rect 526 1437 527 1441
rect 531 1437 532 1441
rect 526 1436 532 1437
rect 598 1441 604 1442
rect 598 1437 599 1441
rect 603 1437 604 1441
rect 598 1436 604 1437
rect 662 1441 668 1442
rect 662 1437 663 1441
rect 667 1437 668 1441
rect 662 1436 668 1437
rect 718 1441 724 1442
rect 718 1437 719 1441
rect 723 1437 724 1441
rect 718 1436 724 1437
rect 782 1441 788 1442
rect 782 1437 783 1441
rect 787 1437 788 1441
rect 782 1436 788 1437
rect 846 1441 852 1442
rect 846 1437 847 1441
rect 851 1437 852 1441
rect 846 1436 852 1437
rect 902 1441 908 1442
rect 902 1437 903 1441
rect 907 1437 908 1441
rect 902 1436 908 1437
rect 958 1441 964 1442
rect 958 1437 959 1441
rect 963 1437 964 1441
rect 958 1436 964 1437
rect 1014 1441 1020 1442
rect 1014 1437 1015 1441
rect 1019 1437 1020 1441
rect 1014 1436 1020 1437
rect 1070 1441 1076 1442
rect 1070 1437 1071 1441
rect 1075 1437 1076 1441
rect 1070 1436 1076 1437
rect 1118 1441 1124 1442
rect 1118 1437 1119 1441
rect 1123 1437 1124 1441
rect 1118 1436 1124 1437
rect 1158 1441 1164 1442
rect 1158 1437 1159 1441
rect 1163 1437 1164 1441
rect 1158 1436 1164 1437
rect 1206 1441 1212 1442
rect 1206 1437 1207 1441
rect 1211 1437 1212 1441
rect 1206 1436 1212 1437
rect 1262 1441 1268 1442
rect 1262 1437 1263 1441
rect 1267 1437 1268 1441
rect 1262 1436 1268 1437
rect 1326 1441 1332 1442
rect 1326 1437 1327 1441
rect 1331 1437 1332 1441
rect 1326 1436 1332 1437
rect 1398 1441 1404 1442
rect 1398 1437 1399 1441
rect 1403 1437 1404 1441
rect 1398 1436 1404 1437
rect 1478 1441 1484 1442
rect 1478 1437 1479 1441
rect 1483 1437 1484 1441
rect 1478 1436 1484 1437
rect 1558 1441 1564 1442
rect 1558 1437 1559 1441
rect 1563 1437 1564 1441
rect 1558 1436 1564 1437
rect 1622 1441 1628 1442
rect 1622 1437 1623 1441
rect 1627 1437 1628 1441
rect 1662 1439 1663 1443
rect 1667 1439 1668 1443
rect 1662 1438 1668 1439
rect 1622 1436 1628 1437
rect 134 1423 140 1424
rect 110 1421 116 1422
rect 110 1417 111 1421
rect 115 1417 116 1421
rect 134 1419 135 1423
rect 139 1419 140 1423
rect 134 1418 140 1419
rect 166 1423 172 1424
rect 166 1419 167 1423
rect 171 1419 172 1423
rect 166 1418 172 1419
rect 214 1423 220 1424
rect 214 1419 215 1423
rect 219 1419 220 1423
rect 214 1418 220 1419
rect 286 1423 292 1424
rect 286 1419 287 1423
rect 291 1419 292 1423
rect 286 1418 292 1419
rect 358 1423 364 1424
rect 358 1419 359 1423
rect 363 1419 364 1423
rect 358 1418 364 1419
rect 438 1423 444 1424
rect 438 1419 439 1423
rect 443 1419 444 1423
rect 438 1418 444 1419
rect 518 1423 524 1424
rect 518 1419 519 1423
rect 523 1419 524 1423
rect 518 1418 524 1419
rect 598 1423 604 1424
rect 598 1419 599 1423
rect 603 1419 604 1423
rect 598 1418 604 1419
rect 678 1423 684 1424
rect 678 1419 679 1423
rect 683 1419 684 1423
rect 678 1418 684 1419
rect 758 1423 764 1424
rect 758 1419 759 1423
rect 763 1419 764 1423
rect 758 1418 764 1419
rect 830 1423 836 1424
rect 830 1419 831 1423
rect 835 1419 836 1423
rect 830 1418 836 1419
rect 902 1423 908 1424
rect 902 1419 903 1423
rect 907 1419 908 1423
rect 902 1418 908 1419
rect 966 1423 972 1424
rect 966 1419 967 1423
rect 971 1419 972 1423
rect 966 1418 972 1419
rect 1030 1423 1036 1424
rect 1030 1419 1031 1423
rect 1035 1419 1036 1423
rect 1030 1418 1036 1419
rect 1102 1423 1108 1424
rect 1102 1419 1103 1423
rect 1107 1419 1108 1423
rect 1102 1418 1108 1419
rect 1166 1423 1172 1424
rect 1166 1419 1167 1423
rect 1171 1419 1172 1423
rect 1166 1418 1172 1419
rect 1230 1423 1236 1424
rect 1230 1419 1231 1423
rect 1235 1419 1236 1423
rect 1230 1418 1236 1419
rect 1294 1423 1300 1424
rect 1294 1419 1295 1423
rect 1299 1419 1300 1423
rect 1294 1418 1300 1419
rect 1358 1423 1364 1424
rect 1358 1419 1359 1423
rect 1363 1419 1364 1423
rect 1358 1418 1364 1419
rect 1414 1423 1420 1424
rect 1414 1419 1415 1423
rect 1419 1419 1420 1423
rect 1414 1418 1420 1419
rect 1462 1423 1468 1424
rect 1462 1419 1463 1423
rect 1467 1419 1468 1423
rect 1462 1418 1468 1419
rect 1502 1423 1508 1424
rect 1502 1419 1503 1423
rect 1507 1419 1508 1423
rect 1502 1418 1508 1419
rect 1550 1423 1556 1424
rect 1550 1419 1551 1423
rect 1555 1419 1556 1423
rect 1550 1418 1556 1419
rect 1590 1423 1596 1424
rect 1590 1419 1591 1423
rect 1595 1419 1596 1423
rect 1590 1418 1596 1419
rect 1622 1423 1628 1424
rect 1622 1419 1623 1423
rect 1627 1419 1628 1423
rect 1622 1418 1628 1419
rect 1662 1421 1668 1422
rect 110 1416 116 1417
rect 1662 1417 1663 1421
rect 1667 1417 1668 1421
rect 1662 1416 1668 1417
rect 134 1406 140 1407
rect 110 1404 116 1405
rect 110 1400 111 1404
rect 115 1400 116 1404
rect 134 1402 135 1406
rect 139 1402 140 1406
rect 134 1401 140 1402
rect 166 1406 172 1407
rect 166 1402 167 1406
rect 171 1402 172 1406
rect 166 1401 172 1402
rect 214 1406 220 1407
rect 214 1402 215 1406
rect 219 1402 220 1406
rect 214 1401 220 1402
rect 286 1406 292 1407
rect 286 1402 287 1406
rect 291 1402 292 1406
rect 286 1401 292 1402
rect 358 1406 364 1407
rect 358 1402 359 1406
rect 363 1402 364 1406
rect 358 1401 364 1402
rect 438 1406 444 1407
rect 438 1402 439 1406
rect 443 1402 444 1406
rect 438 1401 444 1402
rect 518 1406 524 1407
rect 518 1402 519 1406
rect 523 1402 524 1406
rect 518 1401 524 1402
rect 598 1406 604 1407
rect 598 1402 599 1406
rect 603 1402 604 1406
rect 598 1401 604 1402
rect 678 1406 684 1407
rect 678 1402 679 1406
rect 683 1402 684 1406
rect 678 1401 684 1402
rect 758 1406 764 1407
rect 758 1402 759 1406
rect 763 1402 764 1406
rect 758 1401 764 1402
rect 830 1406 836 1407
rect 830 1402 831 1406
rect 835 1402 836 1406
rect 830 1401 836 1402
rect 902 1406 908 1407
rect 902 1402 903 1406
rect 907 1402 908 1406
rect 902 1401 908 1402
rect 966 1406 972 1407
rect 966 1402 967 1406
rect 971 1402 972 1406
rect 966 1401 972 1402
rect 1030 1406 1036 1407
rect 1030 1402 1031 1406
rect 1035 1402 1036 1406
rect 1030 1401 1036 1402
rect 1102 1406 1108 1407
rect 1102 1402 1103 1406
rect 1107 1402 1108 1406
rect 1102 1401 1108 1402
rect 1166 1406 1172 1407
rect 1166 1402 1167 1406
rect 1171 1402 1172 1406
rect 1166 1401 1172 1402
rect 1230 1406 1236 1407
rect 1230 1402 1231 1406
rect 1235 1402 1236 1406
rect 1230 1401 1236 1402
rect 1294 1406 1300 1407
rect 1294 1402 1295 1406
rect 1299 1402 1300 1406
rect 1294 1401 1300 1402
rect 1358 1406 1364 1407
rect 1358 1402 1359 1406
rect 1363 1402 1364 1406
rect 1358 1401 1364 1402
rect 1414 1406 1420 1407
rect 1414 1402 1415 1406
rect 1419 1402 1420 1406
rect 1414 1401 1420 1402
rect 1462 1406 1468 1407
rect 1462 1402 1463 1406
rect 1467 1402 1468 1406
rect 1462 1401 1468 1402
rect 1502 1406 1508 1407
rect 1502 1402 1503 1406
rect 1507 1402 1508 1406
rect 1502 1401 1508 1402
rect 1550 1406 1556 1407
rect 1550 1402 1551 1406
rect 1555 1402 1556 1406
rect 1550 1401 1556 1402
rect 1590 1406 1596 1407
rect 1590 1402 1591 1406
rect 1595 1402 1596 1406
rect 1590 1401 1596 1402
rect 1622 1406 1628 1407
rect 1622 1402 1623 1406
rect 1627 1402 1628 1406
rect 1622 1401 1628 1402
rect 1662 1404 1668 1405
rect 110 1399 116 1400
rect 1662 1400 1663 1404
rect 1667 1400 1668 1404
rect 1662 1399 1668 1400
rect 110 1376 116 1377
rect 110 1372 111 1376
rect 115 1372 116 1376
rect 1662 1376 1668 1377
rect 110 1371 116 1372
rect 134 1374 140 1375
rect 134 1370 135 1374
rect 139 1370 140 1374
rect 134 1369 140 1370
rect 166 1374 172 1375
rect 166 1370 167 1374
rect 171 1370 172 1374
rect 166 1369 172 1370
rect 222 1374 228 1375
rect 222 1370 223 1374
rect 227 1370 228 1374
rect 222 1369 228 1370
rect 286 1374 292 1375
rect 286 1370 287 1374
rect 291 1370 292 1374
rect 286 1369 292 1370
rect 358 1374 364 1375
rect 358 1370 359 1374
rect 363 1370 364 1374
rect 358 1369 364 1370
rect 430 1374 436 1375
rect 430 1370 431 1374
rect 435 1370 436 1374
rect 430 1369 436 1370
rect 502 1374 508 1375
rect 502 1370 503 1374
rect 507 1370 508 1374
rect 502 1369 508 1370
rect 582 1374 588 1375
rect 582 1370 583 1374
rect 587 1370 588 1374
rect 582 1369 588 1370
rect 662 1374 668 1375
rect 662 1370 663 1374
rect 667 1370 668 1374
rect 662 1369 668 1370
rect 742 1374 748 1375
rect 742 1370 743 1374
rect 747 1370 748 1374
rect 742 1369 748 1370
rect 814 1374 820 1375
rect 814 1370 815 1374
rect 819 1370 820 1374
rect 814 1369 820 1370
rect 886 1374 892 1375
rect 886 1370 887 1374
rect 891 1370 892 1374
rect 886 1369 892 1370
rect 958 1374 964 1375
rect 958 1370 959 1374
rect 963 1370 964 1374
rect 958 1369 964 1370
rect 1030 1374 1036 1375
rect 1030 1370 1031 1374
rect 1035 1370 1036 1374
rect 1030 1369 1036 1370
rect 1102 1374 1108 1375
rect 1102 1370 1103 1374
rect 1107 1370 1108 1374
rect 1102 1369 1108 1370
rect 1174 1374 1180 1375
rect 1174 1370 1175 1374
rect 1179 1370 1180 1374
rect 1174 1369 1180 1370
rect 1238 1374 1244 1375
rect 1238 1370 1239 1374
rect 1243 1370 1244 1374
rect 1238 1369 1244 1370
rect 1302 1374 1308 1375
rect 1302 1370 1303 1374
rect 1307 1370 1308 1374
rect 1302 1369 1308 1370
rect 1366 1374 1372 1375
rect 1366 1370 1367 1374
rect 1371 1370 1372 1374
rect 1366 1369 1372 1370
rect 1430 1374 1436 1375
rect 1430 1370 1431 1374
rect 1435 1370 1436 1374
rect 1430 1369 1436 1370
rect 1494 1374 1500 1375
rect 1494 1370 1495 1374
rect 1499 1370 1500 1374
rect 1494 1369 1500 1370
rect 1566 1374 1572 1375
rect 1566 1370 1567 1374
rect 1571 1370 1572 1374
rect 1566 1369 1572 1370
rect 1622 1374 1628 1375
rect 1622 1370 1623 1374
rect 1627 1370 1628 1374
rect 1662 1372 1663 1376
rect 1667 1372 1668 1376
rect 1662 1371 1668 1372
rect 1622 1369 1628 1370
rect 110 1359 116 1360
rect 110 1355 111 1359
rect 115 1355 116 1359
rect 1662 1359 1668 1360
rect 110 1354 116 1355
rect 134 1357 140 1358
rect 134 1353 135 1357
rect 139 1353 140 1357
rect 134 1352 140 1353
rect 166 1357 172 1358
rect 166 1353 167 1357
rect 171 1353 172 1357
rect 166 1352 172 1353
rect 222 1357 228 1358
rect 222 1353 223 1357
rect 227 1353 228 1357
rect 222 1352 228 1353
rect 286 1357 292 1358
rect 286 1353 287 1357
rect 291 1353 292 1357
rect 286 1352 292 1353
rect 358 1357 364 1358
rect 358 1353 359 1357
rect 363 1353 364 1357
rect 358 1352 364 1353
rect 430 1357 436 1358
rect 430 1353 431 1357
rect 435 1353 436 1357
rect 430 1352 436 1353
rect 502 1357 508 1358
rect 502 1353 503 1357
rect 507 1353 508 1357
rect 502 1352 508 1353
rect 582 1357 588 1358
rect 582 1353 583 1357
rect 587 1353 588 1357
rect 582 1352 588 1353
rect 662 1357 668 1358
rect 662 1353 663 1357
rect 667 1353 668 1357
rect 662 1352 668 1353
rect 742 1357 748 1358
rect 742 1353 743 1357
rect 747 1353 748 1357
rect 742 1352 748 1353
rect 814 1357 820 1358
rect 814 1353 815 1357
rect 819 1353 820 1357
rect 814 1352 820 1353
rect 886 1357 892 1358
rect 886 1353 887 1357
rect 891 1353 892 1357
rect 886 1352 892 1353
rect 958 1357 964 1358
rect 958 1353 959 1357
rect 963 1353 964 1357
rect 958 1352 964 1353
rect 1030 1357 1036 1358
rect 1030 1353 1031 1357
rect 1035 1353 1036 1357
rect 1030 1352 1036 1353
rect 1102 1357 1108 1358
rect 1102 1353 1103 1357
rect 1107 1353 1108 1357
rect 1102 1352 1108 1353
rect 1174 1357 1180 1358
rect 1174 1353 1175 1357
rect 1179 1353 1180 1357
rect 1174 1352 1180 1353
rect 1238 1357 1244 1358
rect 1238 1353 1239 1357
rect 1243 1353 1244 1357
rect 1238 1352 1244 1353
rect 1302 1357 1308 1358
rect 1302 1353 1303 1357
rect 1307 1353 1308 1357
rect 1302 1352 1308 1353
rect 1366 1357 1372 1358
rect 1366 1353 1367 1357
rect 1371 1353 1372 1357
rect 1366 1352 1372 1353
rect 1430 1357 1436 1358
rect 1430 1353 1431 1357
rect 1435 1353 1436 1357
rect 1430 1352 1436 1353
rect 1494 1357 1500 1358
rect 1494 1353 1495 1357
rect 1499 1353 1500 1357
rect 1494 1352 1500 1353
rect 1566 1357 1572 1358
rect 1566 1353 1567 1357
rect 1571 1353 1572 1357
rect 1566 1352 1572 1353
rect 1622 1357 1628 1358
rect 1622 1353 1623 1357
rect 1627 1353 1628 1357
rect 1662 1355 1663 1359
rect 1667 1355 1668 1359
rect 1662 1354 1668 1355
rect 1622 1352 1628 1353
rect 134 1343 140 1344
rect 110 1341 116 1342
rect 110 1337 111 1341
rect 115 1337 116 1341
rect 134 1339 135 1343
rect 139 1339 140 1343
rect 134 1338 140 1339
rect 182 1343 188 1344
rect 182 1339 183 1343
rect 187 1339 188 1343
rect 182 1338 188 1339
rect 238 1343 244 1344
rect 238 1339 239 1343
rect 243 1339 244 1343
rect 238 1338 244 1339
rect 294 1343 300 1344
rect 294 1339 295 1343
rect 299 1339 300 1343
rect 294 1338 300 1339
rect 350 1343 356 1344
rect 350 1339 351 1343
rect 355 1339 356 1343
rect 350 1338 356 1339
rect 398 1343 404 1344
rect 398 1339 399 1343
rect 403 1339 404 1343
rect 398 1338 404 1339
rect 454 1343 460 1344
rect 454 1339 455 1343
rect 459 1339 460 1343
rect 454 1338 460 1339
rect 510 1343 516 1344
rect 510 1339 511 1343
rect 515 1339 516 1343
rect 510 1338 516 1339
rect 566 1343 572 1344
rect 566 1339 567 1343
rect 571 1339 572 1343
rect 566 1338 572 1339
rect 630 1343 636 1344
rect 630 1339 631 1343
rect 635 1339 636 1343
rect 630 1338 636 1339
rect 694 1343 700 1344
rect 694 1339 695 1343
rect 699 1339 700 1343
rect 694 1338 700 1339
rect 758 1343 764 1344
rect 758 1339 759 1343
rect 763 1339 764 1343
rect 758 1338 764 1339
rect 822 1343 828 1344
rect 822 1339 823 1343
rect 827 1339 828 1343
rect 822 1338 828 1339
rect 886 1343 892 1344
rect 886 1339 887 1343
rect 891 1339 892 1343
rect 886 1338 892 1339
rect 958 1343 964 1344
rect 958 1339 959 1343
rect 963 1339 964 1343
rect 958 1338 964 1339
rect 1022 1343 1028 1344
rect 1022 1339 1023 1343
rect 1027 1339 1028 1343
rect 1022 1338 1028 1339
rect 1086 1343 1092 1344
rect 1086 1339 1087 1343
rect 1091 1339 1092 1343
rect 1086 1338 1092 1339
rect 1150 1343 1156 1344
rect 1150 1339 1151 1343
rect 1155 1339 1156 1343
rect 1150 1338 1156 1339
rect 1214 1343 1220 1344
rect 1214 1339 1215 1343
rect 1219 1339 1220 1343
rect 1214 1338 1220 1339
rect 1278 1343 1284 1344
rect 1278 1339 1279 1343
rect 1283 1339 1284 1343
rect 1278 1338 1284 1339
rect 1342 1343 1348 1344
rect 1342 1339 1343 1343
rect 1347 1339 1348 1343
rect 1342 1338 1348 1339
rect 1406 1343 1412 1344
rect 1406 1339 1407 1343
rect 1411 1339 1412 1343
rect 1406 1338 1412 1339
rect 1478 1343 1484 1344
rect 1478 1339 1479 1343
rect 1483 1339 1484 1343
rect 1478 1338 1484 1339
rect 1558 1343 1564 1344
rect 1558 1339 1559 1343
rect 1563 1339 1564 1343
rect 1558 1338 1564 1339
rect 1622 1343 1628 1344
rect 1622 1339 1623 1343
rect 1627 1339 1628 1343
rect 1622 1338 1628 1339
rect 1662 1341 1668 1342
rect 110 1336 116 1337
rect 1662 1337 1663 1341
rect 1667 1337 1668 1341
rect 1662 1336 1668 1337
rect 134 1326 140 1327
rect 110 1324 116 1325
rect 110 1320 111 1324
rect 115 1320 116 1324
rect 134 1322 135 1326
rect 139 1322 140 1326
rect 134 1321 140 1322
rect 182 1326 188 1327
rect 182 1322 183 1326
rect 187 1322 188 1326
rect 182 1321 188 1322
rect 238 1326 244 1327
rect 238 1322 239 1326
rect 243 1322 244 1326
rect 238 1321 244 1322
rect 294 1326 300 1327
rect 294 1322 295 1326
rect 299 1322 300 1326
rect 294 1321 300 1322
rect 350 1326 356 1327
rect 350 1322 351 1326
rect 355 1322 356 1326
rect 350 1321 356 1322
rect 398 1326 404 1327
rect 398 1322 399 1326
rect 403 1322 404 1326
rect 398 1321 404 1322
rect 454 1326 460 1327
rect 454 1322 455 1326
rect 459 1322 460 1326
rect 454 1321 460 1322
rect 510 1326 516 1327
rect 510 1322 511 1326
rect 515 1322 516 1326
rect 510 1321 516 1322
rect 566 1326 572 1327
rect 566 1322 567 1326
rect 571 1322 572 1326
rect 566 1321 572 1322
rect 630 1326 636 1327
rect 630 1322 631 1326
rect 635 1322 636 1326
rect 630 1321 636 1322
rect 694 1326 700 1327
rect 694 1322 695 1326
rect 699 1322 700 1326
rect 694 1321 700 1322
rect 758 1326 764 1327
rect 758 1322 759 1326
rect 763 1322 764 1326
rect 758 1321 764 1322
rect 822 1326 828 1327
rect 822 1322 823 1326
rect 827 1322 828 1326
rect 822 1321 828 1322
rect 886 1326 892 1327
rect 886 1322 887 1326
rect 891 1322 892 1326
rect 886 1321 892 1322
rect 958 1326 964 1327
rect 958 1322 959 1326
rect 963 1322 964 1326
rect 958 1321 964 1322
rect 1022 1326 1028 1327
rect 1022 1322 1023 1326
rect 1027 1322 1028 1326
rect 1022 1321 1028 1322
rect 1086 1326 1092 1327
rect 1086 1322 1087 1326
rect 1091 1322 1092 1326
rect 1086 1321 1092 1322
rect 1150 1326 1156 1327
rect 1150 1322 1151 1326
rect 1155 1322 1156 1326
rect 1150 1321 1156 1322
rect 1214 1326 1220 1327
rect 1214 1322 1215 1326
rect 1219 1322 1220 1326
rect 1214 1321 1220 1322
rect 1278 1326 1284 1327
rect 1278 1322 1279 1326
rect 1283 1322 1284 1326
rect 1278 1321 1284 1322
rect 1342 1326 1348 1327
rect 1342 1322 1343 1326
rect 1347 1322 1348 1326
rect 1342 1321 1348 1322
rect 1406 1326 1412 1327
rect 1406 1322 1407 1326
rect 1411 1322 1412 1326
rect 1406 1321 1412 1322
rect 1478 1326 1484 1327
rect 1478 1322 1479 1326
rect 1483 1322 1484 1326
rect 1478 1321 1484 1322
rect 1558 1326 1564 1327
rect 1558 1322 1559 1326
rect 1563 1322 1564 1326
rect 1558 1321 1564 1322
rect 1622 1326 1628 1327
rect 1622 1322 1623 1326
rect 1627 1322 1628 1326
rect 1622 1321 1628 1322
rect 1662 1324 1668 1325
rect 110 1319 116 1320
rect 1662 1320 1663 1324
rect 1667 1320 1668 1324
rect 1662 1319 1668 1320
rect 110 1292 116 1293
rect 110 1288 111 1292
rect 115 1288 116 1292
rect 1662 1292 1668 1293
rect 110 1287 116 1288
rect 134 1290 140 1291
rect 134 1286 135 1290
rect 139 1286 140 1290
rect 134 1285 140 1286
rect 182 1290 188 1291
rect 182 1286 183 1290
rect 187 1286 188 1290
rect 182 1285 188 1286
rect 230 1290 236 1291
rect 230 1286 231 1290
rect 235 1286 236 1290
rect 230 1285 236 1286
rect 278 1290 284 1291
rect 278 1286 279 1290
rect 283 1286 284 1290
rect 278 1285 284 1286
rect 326 1290 332 1291
rect 326 1286 327 1290
rect 331 1286 332 1290
rect 326 1285 332 1286
rect 374 1290 380 1291
rect 374 1286 375 1290
rect 379 1286 380 1290
rect 374 1285 380 1286
rect 430 1290 436 1291
rect 430 1286 431 1290
rect 435 1286 436 1290
rect 430 1285 436 1286
rect 486 1290 492 1291
rect 486 1286 487 1290
rect 491 1286 492 1290
rect 486 1285 492 1286
rect 542 1290 548 1291
rect 542 1286 543 1290
rect 547 1286 548 1290
rect 542 1285 548 1286
rect 606 1290 612 1291
rect 606 1286 607 1290
rect 611 1286 612 1290
rect 606 1285 612 1286
rect 662 1290 668 1291
rect 662 1286 663 1290
rect 667 1286 668 1290
rect 662 1285 668 1286
rect 718 1290 724 1291
rect 718 1286 719 1290
rect 723 1286 724 1290
rect 718 1285 724 1286
rect 774 1290 780 1291
rect 774 1286 775 1290
rect 779 1286 780 1290
rect 774 1285 780 1286
rect 830 1290 836 1291
rect 830 1286 831 1290
rect 835 1286 836 1290
rect 830 1285 836 1286
rect 894 1290 900 1291
rect 894 1286 895 1290
rect 899 1286 900 1290
rect 894 1285 900 1286
rect 958 1290 964 1291
rect 958 1286 959 1290
rect 963 1286 964 1290
rect 958 1285 964 1286
rect 1022 1290 1028 1291
rect 1022 1286 1023 1290
rect 1027 1286 1028 1290
rect 1022 1285 1028 1286
rect 1078 1290 1084 1291
rect 1078 1286 1079 1290
rect 1083 1286 1084 1290
rect 1078 1285 1084 1286
rect 1142 1290 1148 1291
rect 1142 1286 1143 1290
rect 1147 1286 1148 1290
rect 1142 1285 1148 1286
rect 1206 1290 1212 1291
rect 1206 1286 1207 1290
rect 1211 1286 1212 1290
rect 1206 1285 1212 1286
rect 1278 1290 1284 1291
rect 1278 1286 1279 1290
rect 1283 1286 1284 1290
rect 1278 1285 1284 1286
rect 1358 1290 1364 1291
rect 1358 1286 1359 1290
rect 1363 1286 1364 1290
rect 1358 1285 1364 1286
rect 1446 1290 1452 1291
rect 1446 1286 1447 1290
rect 1451 1286 1452 1290
rect 1446 1285 1452 1286
rect 1542 1290 1548 1291
rect 1542 1286 1543 1290
rect 1547 1286 1548 1290
rect 1542 1285 1548 1286
rect 1622 1290 1628 1291
rect 1622 1286 1623 1290
rect 1627 1286 1628 1290
rect 1662 1288 1663 1292
rect 1667 1288 1668 1292
rect 1662 1287 1668 1288
rect 1622 1285 1628 1286
rect 110 1275 116 1276
rect 110 1271 111 1275
rect 115 1271 116 1275
rect 1662 1275 1668 1276
rect 110 1270 116 1271
rect 134 1273 140 1274
rect 134 1269 135 1273
rect 139 1269 140 1273
rect 134 1268 140 1269
rect 182 1273 188 1274
rect 182 1269 183 1273
rect 187 1269 188 1273
rect 182 1268 188 1269
rect 230 1273 236 1274
rect 230 1269 231 1273
rect 235 1269 236 1273
rect 230 1268 236 1269
rect 278 1273 284 1274
rect 278 1269 279 1273
rect 283 1269 284 1273
rect 278 1268 284 1269
rect 326 1273 332 1274
rect 326 1269 327 1273
rect 331 1269 332 1273
rect 326 1268 332 1269
rect 374 1273 380 1274
rect 374 1269 375 1273
rect 379 1269 380 1273
rect 374 1268 380 1269
rect 430 1273 436 1274
rect 430 1269 431 1273
rect 435 1269 436 1273
rect 430 1268 436 1269
rect 486 1273 492 1274
rect 486 1269 487 1273
rect 491 1269 492 1273
rect 486 1268 492 1269
rect 542 1273 548 1274
rect 542 1269 543 1273
rect 547 1269 548 1273
rect 542 1268 548 1269
rect 606 1273 612 1274
rect 606 1269 607 1273
rect 611 1269 612 1273
rect 606 1268 612 1269
rect 662 1273 668 1274
rect 662 1269 663 1273
rect 667 1269 668 1273
rect 662 1268 668 1269
rect 718 1273 724 1274
rect 718 1269 719 1273
rect 723 1269 724 1273
rect 718 1268 724 1269
rect 774 1273 780 1274
rect 774 1269 775 1273
rect 779 1269 780 1273
rect 774 1268 780 1269
rect 830 1273 836 1274
rect 830 1269 831 1273
rect 835 1269 836 1273
rect 830 1268 836 1269
rect 894 1273 900 1274
rect 894 1269 895 1273
rect 899 1269 900 1273
rect 894 1268 900 1269
rect 958 1273 964 1274
rect 958 1269 959 1273
rect 963 1269 964 1273
rect 958 1268 964 1269
rect 1022 1273 1028 1274
rect 1022 1269 1023 1273
rect 1027 1269 1028 1273
rect 1022 1268 1028 1269
rect 1078 1273 1084 1274
rect 1078 1269 1079 1273
rect 1083 1269 1084 1273
rect 1078 1268 1084 1269
rect 1142 1273 1148 1274
rect 1142 1269 1143 1273
rect 1147 1269 1148 1273
rect 1142 1268 1148 1269
rect 1206 1273 1212 1274
rect 1206 1269 1207 1273
rect 1211 1269 1212 1273
rect 1206 1268 1212 1269
rect 1278 1273 1284 1274
rect 1278 1269 1279 1273
rect 1283 1269 1284 1273
rect 1278 1268 1284 1269
rect 1358 1273 1364 1274
rect 1358 1269 1359 1273
rect 1363 1269 1364 1273
rect 1358 1268 1364 1269
rect 1446 1273 1452 1274
rect 1446 1269 1447 1273
rect 1451 1269 1452 1273
rect 1446 1268 1452 1269
rect 1542 1273 1548 1274
rect 1542 1269 1543 1273
rect 1547 1269 1548 1273
rect 1542 1268 1548 1269
rect 1622 1273 1628 1274
rect 1622 1269 1623 1273
rect 1627 1269 1628 1273
rect 1662 1271 1663 1275
rect 1667 1271 1668 1275
rect 1662 1270 1668 1271
rect 1622 1268 1628 1269
rect 134 1259 140 1260
rect 110 1257 116 1258
rect 110 1253 111 1257
rect 115 1253 116 1257
rect 134 1255 135 1259
rect 139 1255 140 1259
rect 134 1254 140 1255
rect 166 1259 172 1260
rect 166 1255 167 1259
rect 171 1255 172 1259
rect 166 1254 172 1255
rect 222 1259 228 1260
rect 222 1255 223 1259
rect 227 1255 228 1259
rect 222 1254 228 1255
rect 278 1259 284 1260
rect 278 1255 279 1259
rect 283 1255 284 1259
rect 278 1254 284 1255
rect 326 1259 332 1260
rect 326 1255 327 1259
rect 331 1255 332 1259
rect 326 1254 332 1255
rect 382 1259 388 1260
rect 382 1255 383 1259
rect 387 1255 388 1259
rect 382 1254 388 1255
rect 438 1259 444 1260
rect 438 1255 439 1259
rect 443 1255 444 1259
rect 438 1254 444 1255
rect 494 1259 500 1260
rect 494 1255 495 1259
rect 499 1255 500 1259
rect 494 1254 500 1255
rect 550 1259 556 1260
rect 550 1255 551 1259
rect 555 1255 556 1259
rect 550 1254 556 1255
rect 606 1259 612 1260
rect 606 1255 607 1259
rect 611 1255 612 1259
rect 606 1254 612 1255
rect 662 1259 668 1260
rect 662 1255 663 1259
rect 667 1255 668 1259
rect 662 1254 668 1255
rect 718 1259 724 1260
rect 718 1255 719 1259
rect 723 1255 724 1259
rect 718 1254 724 1255
rect 766 1259 772 1260
rect 766 1255 767 1259
rect 771 1255 772 1259
rect 766 1254 772 1255
rect 814 1259 820 1260
rect 814 1255 815 1259
rect 819 1255 820 1259
rect 814 1254 820 1255
rect 870 1259 876 1260
rect 870 1255 871 1259
rect 875 1255 876 1259
rect 870 1254 876 1255
rect 926 1259 932 1260
rect 926 1255 927 1259
rect 931 1255 932 1259
rect 926 1254 932 1255
rect 982 1259 988 1260
rect 982 1255 983 1259
rect 987 1255 988 1259
rect 982 1254 988 1255
rect 1038 1259 1044 1260
rect 1038 1255 1039 1259
rect 1043 1255 1044 1259
rect 1038 1254 1044 1255
rect 1094 1259 1100 1260
rect 1094 1255 1095 1259
rect 1099 1255 1100 1259
rect 1094 1254 1100 1255
rect 1158 1259 1164 1260
rect 1158 1255 1159 1259
rect 1163 1255 1164 1259
rect 1158 1254 1164 1255
rect 1230 1259 1236 1260
rect 1230 1255 1231 1259
rect 1235 1255 1236 1259
rect 1230 1254 1236 1255
rect 1318 1259 1324 1260
rect 1318 1255 1319 1259
rect 1323 1255 1324 1259
rect 1318 1254 1324 1255
rect 1422 1259 1428 1260
rect 1422 1255 1423 1259
rect 1427 1255 1428 1259
rect 1422 1254 1428 1255
rect 1534 1259 1540 1260
rect 1534 1255 1535 1259
rect 1539 1255 1540 1259
rect 1534 1254 1540 1255
rect 1622 1259 1628 1260
rect 1622 1255 1623 1259
rect 1627 1255 1628 1259
rect 1622 1254 1628 1255
rect 1662 1257 1668 1258
rect 110 1252 116 1253
rect 1662 1253 1663 1257
rect 1667 1253 1668 1257
rect 1662 1252 1668 1253
rect 134 1242 140 1243
rect 110 1240 116 1241
rect 110 1236 111 1240
rect 115 1236 116 1240
rect 134 1238 135 1242
rect 139 1238 140 1242
rect 134 1237 140 1238
rect 166 1242 172 1243
rect 166 1238 167 1242
rect 171 1238 172 1242
rect 166 1237 172 1238
rect 222 1242 228 1243
rect 222 1238 223 1242
rect 227 1238 228 1242
rect 222 1237 228 1238
rect 278 1242 284 1243
rect 278 1238 279 1242
rect 283 1238 284 1242
rect 278 1237 284 1238
rect 326 1242 332 1243
rect 326 1238 327 1242
rect 331 1238 332 1242
rect 326 1237 332 1238
rect 382 1242 388 1243
rect 382 1238 383 1242
rect 387 1238 388 1242
rect 382 1237 388 1238
rect 438 1242 444 1243
rect 438 1238 439 1242
rect 443 1238 444 1242
rect 438 1237 444 1238
rect 494 1242 500 1243
rect 494 1238 495 1242
rect 499 1238 500 1242
rect 494 1237 500 1238
rect 550 1242 556 1243
rect 550 1238 551 1242
rect 555 1238 556 1242
rect 550 1237 556 1238
rect 606 1242 612 1243
rect 606 1238 607 1242
rect 611 1238 612 1242
rect 606 1237 612 1238
rect 662 1242 668 1243
rect 662 1238 663 1242
rect 667 1238 668 1242
rect 662 1237 668 1238
rect 718 1242 724 1243
rect 718 1238 719 1242
rect 723 1238 724 1242
rect 718 1237 724 1238
rect 766 1242 772 1243
rect 766 1238 767 1242
rect 771 1238 772 1242
rect 766 1237 772 1238
rect 814 1242 820 1243
rect 814 1238 815 1242
rect 819 1238 820 1242
rect 814 1237 820 1238
rect 870 1242 876 1243
rect 870 1238 871 1242
rect 875 1238 876 1242
rect 870 1237 876 1238
rect 926 1242 932 1243
rect 926 1238 927 1242
rect 931 1238 932 1242
rect 926 1237 932 1238
rect 982 1242 988 1243
rect 982 1238 983 1242
rect 987 1238 988 1242
rect 982 1237 988 1238
rect 1038 1242 1044 1243
rect 1038 1238 1039 1242
rect 1043 1238 1044 1242
rect 1038 1237 1044 1238
rect 1094 1242 1100 1243
rect 1094 1238 1095 1242
rect 1099 1238 1100 1242
rect 1094 1237 1100 1238
rect 1158 1242 1164 1243
rect 1158 1238 1159 1242
rect 1163 1238 1164 1242
rect 1158 1237 1164 1238
rect 1230 1242 1236 1243
rect 1230 1238 1231 1242
rect 1235 1238 1236 1242
rect 1230 1237 1236 1238
rect 1318 1242 1324 1243
rect 1318 1238 1319 1242
rect 1323 1238 1324 1242
rect 1318 1237 1324 1238
rect 1422 1242 1428 1243
rect 1422 1238 1423 1242
rect 1427 1238 1428 1242
rect 1422 1237 1428 1238
rect 1534 1242 1540 1243
rect 1534 1238 1535 1242
rect 1539 1238 1540 1242
rect 1534 1237 1540 1238
rect 1622 1242 1628 1243
rect 1622 1238 1623 1242
rect 1627 1238 1628 1242
rect 1622 1237 1628 1238
rect 1662 1240 1668 1241
rect 110 1235 116 1236
rect 1662 1236 1663 1240
rect 1667 1236 1668 1240
rect 1662 1235 1668 1236
rect 110 1208 116 1209
rect 110 1204 111 1208
rect 115 1204 116 1208
rect 1662 1208 1668 1209
rect 110 1203 116 1204
rect 134 1206 140 1207
rect 134 1202 135 1206
rect 139 1202 140 1206
rect 134 1201 140 1202
rect 166 1206 172 1207
rect 166 1202 167 1206
rect 171 1202 172 1206
rect 166 1201 172 1202
rect 222 1206 228 1207
rect 222 1202 223 1206
rect 227 1202 228 1206
rect 222 1201 228 1202
rect 278 1206 284 1207
rect 278 1202 279 1206
rect 283 1202 284 1206
rect 278 1201 284 1202
rect 334 1206 340 1207
rect 334 1202 335 1206
rect 339 1202 340 1206
rect 334 1201 340 1202
rect 382 1206 388 1207
rect 382 1202 383 1206
rect 387 1202 388 1206
rect 382 1201 388 1202
rect 430 1206 436 1207
rect 430 1202 431 1206
rect 435 1202 436 1206
rect 430 1201 436 1202
rect 486 1206 492 1207
rect 486 1202 487 1206
rect 491 1202 492 1206
rect 486 1201 492 1202
rect 542 1206 548 1207
rect 542 1202 543 1206
rect 547 1202 548 1206
rect 542 1201 548 1202
rect 598 1206 604 1207
rect 598 1202 599 1206
rect 603 1202 604 1206
rect 598 1201 604 1202
rect 654 1206 660 1207
rect 654 1202 655 1206
rect 659 1202 660 1206
rect 654 1201 660 1202
rect 710 1206 716 1207
rect 710 1202 711 1206
rect 715 1202 716 1206
rect 710 1201 716 1202
rect 766 1206 772 1207
rect 766 1202 767 1206
rect 771 1202 772 1206
rect 766 1201 772 1202
rect 822 1206 828 1207
rect 822 1202 823 1206
rect 827 1202 828 1206
rect 822 1201 828 1202
rect 886 1206 892 1207
rect 886 1202 887 1206
rect 891 1202 892 1206
rect 886 1201 892 1202
rect 950 1206 956 1207
rect 950 1202 951 1206
rect 955 1202 956 1206
rect 950 1201 956 1202
rect 1014 1206 1020 1207
rect 1014 1202 1015 1206
rect 1019 1202 1020 1206
rect 1014 1201 1020 1202
rect 1078 1206 1084 1207
rect 1078 1202 1079 1206
rect 1083 1202 1084 1206
rect 1078 1201 1084 1202
rect 1142 1206 1148 1207
rect 1142 1202 1143 1206
rect 1147 1202 1148 1206
rect 1142 1201 1148 1202
rect 1206 1206 1212 1207
rect 1206 1202 1207 1206
rect 1211 1202 1212 1206
rect 1206 1201 1212 1202
rect 1278 1206 1284 1207
rect 1278 1202 1279 1206
rect 1283 1202 1284 1206
rect 1278 1201 1284 1202
rect 1358 1206 1364 1207
rect 1358 1202 1359 1206
rect 1363 1202 1364 1206
rect 1358 1201 1364 1202
rect 1446 1206 1452 1207
rect 1446 1202 1447 1206
rect 1451 1202 1452 1206
rect 1446 1201 1452 1202
rect 1542 1206 1548 1207
rect 1542 1202 1543 1206
rect 1547 1202 1548 1206
rect 1542 1201 1548 1202
rect 1622 1206 1628 1207
rect 1622 1202 1623 1206
rect 1627 1202 1628 1206
rect 1662 1204 1663 1208
rect 1667 1204 1668 1208
rect 1662 1203 1668 1204
rect 1622 1201 1628 1202
rect 110 1191 116 1192
rect 110 1187 111 1191
rect 115 1187 116 1191
rect 1662 1191 1668 1192
rect 110 1186 116 1187
rect 134 1189 140 1190
rect 134 1185 135 1189
rect 139 1185 140 1189
rect 134 1184 140 1185
rect 166 1189 172 1190
rect 166 1185 167 1189
rect 171 1185 172 1189
rect 166 1184 172 1185
rect 222 1189 228 1190
rect 222 1185 223 1189
rect 227 1185 228 1189
rect 222 1184 228 1185
rect 278 1189 284 1190
rect 278 1185 279 1189
rect 283 1185 284 1189
rect 278 1184 284 1185
rect 334 1189 340 1190
rect 334 1185 335 1189
rect 339 1185 340 1189
rect 334 1184 340 1185
rect 382 1189 388 1190
rect 382 1185 383 1189
rect 387 1185 388 1189
rect 382 1184 388 1185
rect 430 1189 436 1190
rect 430 1185 431 1189
rect 435 1185 436 1189
rect 430 1184 436 1185
rect 486 1189 492 1190
rect 486 1185 487 1189
rect 491 1185 492 1189
rect 486 1184 492 1185
rect 542 1189 548 1190
rect 542 1185 543 1189
rect 547 1185 548 1189
rect 542 1184 548 1185
rect 598 1189 604 1190
rect 598 1185 599 1189
rect 603 1185 604 1189
rect 598 1184 604 1185
rect 654 1189 660 1190
rect 654 1185 655 1189
rect 659 1185 660 1189
rect 654 1184 660 1185
rect 710 1189 716 1190
rect 710 1185 711 1189
rect 715 1185 716 1189
rect 710 1184 716 1185
rect 766 1189 772 1190
rect 766 1185 767 1189
rect 771 1185 772 1189
rect 766 1184 772 1185
rect 822 1189 828 1190
rect 822 1185 823 1189
rect 827 1185 828 1189
rect 822 1184 828 1185
rect 886 1189 892 1190
rect 886 1185 887 1189
rect 891 1185 892 1189
rect 886 1184 892 1185
rect 950 1189 956 1190
rect 950 1185 951 1189
rect 955 1185 956 1189
rect 950 1184 956 1185
rect 1014 1189 1020 1190
rect 1014 1185 1015 1189
rect 1019 1185 1020 1189
rect 1014 1184 1020 1185
rect 1078 1189 1084 1190
rect 1078 1185 1079 1189
rect 1083 1185 1084 1189
rect 1078 1184 1084 1185
rect 1142 1189 1148 1190
rect 1142 1185 1143 1189
rect 1147 1185 1148 1189
rect 1142 1184 1148 1185
rect 1206 1189 1212 1190
rect 1206 1185 1207 1189
rect 1211 1185 1212 1189
rect 1206 1184 1212 1185
rect 1278 1189 1284 1190
rect 1278 1185 1279 1189
rect 1283 1185 1284 1189
rect 1278 1184 1284 1185
rect 1358 1189 1364 1190
rect 1358 1185 1359 1189
rect 1363 1185 1364 1189
rect 1358 1184 1364 1185
rect 1446 1189 1452 1190
rect 1446 1185 1447 1189
rect 1451 1185 1452 1189
rect 1446 1184 1452 1185
rect 1542 1189 1548 1190
rect 1542 1185 1543 1189
rect 1547 1185 1548 1189
rect 1542 1184 1548 1185
rect 1622 1189 1628 1190
rect 1622 1185 1623 1189
rect 1627 1185 1628 1189
rect 1662 1187 1663 1191
rect 1667 1187 1668 1191
rect 1662 1186 1668 1187
rect 1622 1184 1628 1185
rect 134 1171 140 1172
rect 110 1169 116 1170
rect 110 1165 111 1169
rect 115 1165 116 1169
rect 134 1167 135 1171
rect 139 1167 140 1171
rect 134 1166 140 1167
rect 166 1171 172 1172
rect 166 1167 167 1171
rect 171 1167 172 1171
rect 166 1166 172 1167
rect 222 1171 228 1172
rect 222 1167 223 1171
rect 227 1167 228 1171
rect 222 1166 228 1167
rect 286 1171 292 1172
rect 286 1167 287 1171
rect 291 1167 292 1171
rect 286 1166 292 1167
rect 350 1171 356 1172
rect 350 1167 351 1171
rect 355 1167 356 1171
rect 350 1166 356 1167
rect 414 1171 420 1172
rect 414 1167 415 1171
rect 419 1167 420 1171
rect 414 1166 420 1167
rect 470 1171 476 1172
rect 470 1167 471 1171
rect 475 1167 476 1171
rect 470 1166 476 1167
rect 534 1171 540 1172
rect 534 1167 535 1171
rect 539 1167 540 1171
rect 534 1166 540 1167
rect 598 1171 604 1172
rect 598 1167 599 1171
rect 603 1167 604 1171
rect 598 1166 604 1167
rect 662 1171 668 1172
rect 662 1167 663 1171
rect 667 1167 668 1171
rect 662 1166 668 1167
rect 726 1171 732 1172
rect 726 1167 727 1171
rect 731 1167 732 1171
rect 726 1166 732 1167
rect 782 1171 788 1172
rect 782 1167 783 1171
rect 787 1167 788 1171
rect 782 1166 788 1167
rect 838 1171 844 1172
rect 838 1167 839 1171
rect 843 1167 844 1171
rect 838 1166 844 1167
rect 902 1171 908 1172
rect 902 1167 903 1171
rect 907 1167 908 1171
rect 902 1166 908 1167
rect 966 1171 972 1172
rect 966 1167 967 1171
rect 971 1167 972 1171
rect 966 1166 972 1167
rect 1030 1171 1036 1172
rect 1030 1167 1031 1171
rect 1035 1167 1036 1171
rect 1030 1166 1036 1167
rect 1094 1171 1100 1172
rect 1094 1167 1095 1171
rect 1099 1167 1100 1171
rect 1094 1166 1100 1167
rect 1158 1171 1164 1172
rect 1158 1167 1159 1171
rect 1163 1167 1164 1171
rect 1158 1166 1164 1167
rect 1214 1171 1220 1172
rect 1214 1167 1215 1171
rect 1219 1167 1220 1171
rect 1214 1166 1220 1167
rect 1278 1171 1284 1172
rect 1278 1167 1279 1171
rect 1283 1167 1284 1171
rect 1278 1166 1284 1167
rect 1342 1171 1348 1172
rect 1342 1167 1343 1171
rect 1347 1167 1348 1171
rect 1342 1166 1348 1167
rect 1406 1171 1412 1172
rect 1406 1167 1407 1171
rect 1411 1167 1412 1171
rect 1406 1166 1412 1167
rect 1478 1171 1484 1172
rect 1478 1167 1479 1171
rect 1483 1167 1484 1171
rect 1478 1166 1484 1167
rect 1558 1171 1564 1172
rect 1558 1167 1559 1171
rect 1563 1167 1564 1171
rect 1558 1166 1564 1167
rect 1622 1171 1628 1172
rect 1622 1167 1623 1171
rect 1627 1167 1628 1171
rect 1622 1166 1628 1167
rect 1662 1169 1668 1170
rect 110 1164 116 1165
rect 1662 1165 1663 1169
rect 1667 1165 1668 1169
rect 1662 1164 1668 1165
rect 134 1154 140 1155
rect 110 1152 116 1153
rect 110 1148 111 1152
rect 115 1148 116 1152
rect 134 1150 135 1154
rect 139 1150 140 1154
rect 134 1149 140 1150
rect 166 1154 172 1155
rect 166 1150 167 1154
rect 171 1150 172 1154
rect 166 1149 172 1150
rect 222 1154 228 1155
rect 222 1150 223 1154
rect 227 1150 228 1154
rect 222 1149 228 1150
rect 286 1154 292 1155
rect 286 1150 287 1154
rect 291 1150 292 1154
rect 286 1149 292 1150
rect 350 1154 356 1155
rect 350 1150 351 1154
rect 355 1150 356 1154
rect 350 1149 356 1150
rect 414 1154 420 1155
rect 414 1150 415 1154
rect 419 1150 420 1154
rect 414 1149 420 1150
rect 470 1154 476 1155
rect 470 1150 471 1154
rect 475 1150 476 1154
rect 470 1149 476 1150
rect 534 1154 540 1155
rect 534 1150 535 1154
rect 539 1150 540 1154
rect 534 1149 540 1150
rect 598 1154 604 1155
rect 598 1150 599 1154
rect 603 1150 604 1154
rect 598 1149 604 1150
rect 662 1154 668 1155
rect 662 1150 663 1154
rect 667 1150 668 1154
rect 662 1149 668 1150
rect 726 1154 732 1155
rect 726 1150 727 1154
rect 731 1150 732 1154
rect 726 1149 732 1150
rect 782 1154 788 1155
rect 782 1150 783 1154
rect 787 1150 788 1154
rect 782 1149 788 1150
rect 838 1154 844 1155
rect 838 1150 839 1154
rect 843 1150 844 1154
rect 838 1149 844 1150
rect 902 1154 908 1155
rect 902 1150 903 1154
rect 907 1150 908 1154
rect 902 1149 908 1150
rect 966 1154 972 1155
rect 966 1150 967 1154
rect 971 1150 972 1154
rect 966 1149 972 1150
rect 1030 1154 1036 1155
rect 1030 1150 1031 1154
rect 1035 1150 1036 1154
rect 1030 1149 1036 1150
rect 1094 1154 1100 1155
rect 1094 1150 1095 1154
rect 1099 1150 1100 1154
rect 1094 1149 1100 1150
rect 1158 1154 1164 1155
rect 1158 1150 1159 1154
rect 1163 1150 1164 1154
rect 1158 1149 1164 1150
rect 1214 1154 1220 1155
rect 1214 1150 1215 1154
rect 1219 1150 1220 1154
rect 1214 1149 1220 1150
rect 1278 1154 1284 1155
rect 1278 1150 1279 1154
rect 1283 1150 1284 1154
rect 1278 1149 1284 1150
rect 1342 1154 1348 1155
rect 1342 1150 1343 1154
rect 1347 1150 1348 1154
rect 1342 1149 1348 1150
rect 1406 1154 1412 1155
rect 1406 1150 1407 1154
rect 1411 1150 1412 1154
rect 1406 1149 1412 1150
rect 1478 1154 1484 1155
rect 1478 1150 1479 1154
rect 1483 1150 1484 1154
rect 1478 1149 1484 1150
rect 1558 1154 1564 1155
rect 1558 1150 1559 1154
rect 1563 1150 1564 1154
rect 1558 1149 1564 1150
rect 1622 1154 1628 1155
rect 1622 1150 1623 1154
rect 1627 1150 1628 1154
rect 1622 1149 1628 1150
rect 1662 1152 1668 1153
rect 110 1147 116 1148
rect 1662 1148 1663 1152
rect 1667 1148 1668 1152
rect 1662 1147 1668 1148
rect 110 1120 116 1121
rect 110 1116 111 1120
rect 115 1116 116 1120
rect 1662 1120 1668 1121
rect 110 1115 116 1116
rect 142 1118 148 1119
rect 142 1114 143 1118
rect 147 1114 148 1118
rect 142 1113 148 1114
rect 174 1118 180 1119
rect 174 1114 175 1118
rect 179 1114 180 1118
rect 174 1113 180 1114
rect 214 1118 220 1119
rect 214 1114 215 1118
rect 219 1114 220 1118
rect 214 1113 220 1114
rect 270 1118 276 1119
rect 270 1114 271 1118
rect 275 1114 276 1118
rect 270 1113 276 1114
rect 334 1118 340 1119
rect 334 1114 335 1118
rect 339 1114 340 1118
rect 334 1113 340 1114
rect 398 1118 404 1119
rect 398 1114 399 1118
rect 403 1114 404 1118
rect 398 1113 404 1114
rect 462 1118 468 1119
rect 462 1114 463 1118
rect 467 1114 468 1118
rect 462 1113 468 1114
rect 526 1118 532 1119
rect 526 1114 527 1118
rect 531 1114 532 1118
rect 526 1113 532 1114
rect 598 1118 604 1119
rect 598 1114 599 1118
rect 603 1114 604 1118
rect 598 1113 604 1114
rect 662 1118 668 1119
rect 662 1114 663 1118
rect 667 1114 668 1118
rect 662 1113 668 1114
rect 726 1118 732 1119
rect 726 1114 727 1118
rect 731 1114 732 1118
rect 726 1113 732 1114
rect 790 1118 796 1119
rect 790 1114 791 1118
rect 795 1114 796 1118
rect 790 1113 796 1114
rect 854 1118 860 1119
rect 854 1114 855 1118
rect 859 1114 860 1118
rect 854 1113 860 1114
rect 910 1118 916 1119
rect 910 1114 911 1118
rect 915 1114 916 1118
rect 910 1113 916 1114
rect 966 1118 972 1119
rect 966 1114 967 1118
rect 971 1114 972 1118
rect 966 1113 972 1114
rect 1022 1118 1028 1119
rect 1022 1114 1023 1118
rect 1027 1114 1028 1118
rect 1022 1113 1028 1114
rect 1086 1118 1092 1119
rect 1086 1114 1087 1118
rect 1091 1114 1092 1118
rect 1086 1113 1092 1114
rect 1150 1118 1156 1119
rect 1150 1114 1151 1118
rect 1155 1114 1156 1118
rect 1150 1113 1156 1114
rect 1214 1118 1220 1119
rect 1214 1114 1215 1118
rect 1219 1114 1220 1118
rect 1214 1113 1220 1114
rect 1278 1118 1284 1119
rect 1278 1114 1279 1118
rect 1283 1114 1284 1118
rect 1278 1113 1284 1114
rect 1334 1118 1340 1119
rect 1334 1114 1335 1118
rect 1339 1114 1340 1118
rect 1334 1113 1340 1114
rect 1390 1118 1396 1119
rect 1390 1114 1391 1118
rect 1395 1114 1396 1118
rect 1390 1113 1396 1114
rect 1446 1118 1452 1119
rect 1446 1114 1447 1118
rect 1451 1114 1452 1118
rect 1446 1113 1452 1114
rect 1494 1118 1500 1119
rect 1494 1114 1495 1118
rect 1499 1114 1500 1118
rect 1494 1113 1500 1114
rect 1542 1118 1548 1119
rect 1542 1114 1543 1118
rect 1547 1114 1548 1118
rect 1542 1113 1548 1114
rect 1590 1118 1596 1119
rect 1590 1114 1591 1118
rect 1595 1114 1596 1118
rect 1590 1113 1596 1114
rect 1622 1118 1628 1119
rect 1622 1114 1623 1118
rect 1627 1114 1628 1118
rect 1662 1116 1663 1120
rect 1667 1116 1668 1120
rect 1662 1115 1668 1116
rect 1622 1113 1628 1114
rect 110 1103 116 1104
rect 110 1099 111 1103
rect 115 1099 116 1103
rect 1662 1103 1668 1104
rect 110 1098 116 1099
rect 142 1101 148 1102
rect 142 1097 143 1101
rect 147 1097 148 1101
rect 142 1096 148 1097
rect 174 1101 180 1102
rect 174 1097 175 1101
rect 179 1097 180 1101
rect 174 1096 180 1097
rect 214 1101 220 1102
rect 214 1097 215 1101
rect 219 1097 220 1101
rect 214 1096 220 1097
rect 270 1101 276 1102
rect 270 1097 271 1101
rect 275 1097 276 1101
rect 270 1096 276 1097
rect 334 1101 340 1102
rect 334 1097 335 1101
rect 339 1097 340 1101
rect 334 1096 340 1097
rect 398 1101 404 1102
rect 398 1097 399 1101
rect 403 1097 404 1101
rect 398 1096 404 1097
rect 462 1101 468 1102
rect 462 1097 463 1101
rect 467 1097 468 1101
rect 462 1096 468 1097
rect 526 1101 532 1102
rect 526 1097 527 1101
rect 531 1097 532 1101
rect 526 1096 532 1097
rect 598 1101 604 1102
rect 598 1097 599 1101
rect 603 1097 604 1101
rect 598 1096 604 1097
rect 662 1101 668 1102
rect 662 1097 663 1101
rect 667 1097 668 1101
rect 662 1096 668 1097
rect 726 1101 732 1102
rect 726 1097 727 1101
rect 731 1097 732 1101
rect 726 1096 732 1097
rect 790 1101 796 1102
rect 790 1097 791 1101
rect 795 1097 796 1101
rect 790 1096 796 1097
rect 854 1101 860 1102
rect 854 1097 855 1101
rect 859 1097 860 1101
rect 854 1096 860 1097
rect 910 1101 916 1102
rect 910 1097 911 1101
rect 915 1097 916 1101
rect 910 1096 916 1097
rect 966 1101 972 1102
rect 966 1097 967 1101
rect 971 1097 972 1101
rect 966 1096 972 1097
rect 1022 1101 1028 1102
rect 1022 1097 1023 1101
rect 1027 1097 1028 1101
rect 1022 1096 1028 1097
rect 1086 1101 1092 1102
rect 1086 1097 1087 1101
rect 1091 1097 1092 1101
rect 1086 1096 1092 1097
rect 1150 1101 1156 1102
rect 1150 1097 1151 1101
rect 1155 1097 1156 1101
rect 1150 1096 1156 1097
rect 1214 1101 1220 1102
rect 1214 1097 1215 1101
rect 1219 1097 1220 1101
rect 1214 1096 1220 1097
rect 1278 1101 1284 1102
rect 1278 1097 1279 1101
rect 1283 1097 1284 1101
rect 1278 1096 1284 1097
rect 1334 1101 1340 1102
rect 1334 1097 1335 1101
rect 1339 1097 1340 1101
rect 1334 1096 1340 1097
rect 1390 1101 1396 1102
rect 1390 1097 1391 1101
rect 1395 1097 1396 1101
rect 1390 1096 1396 1097
rect 1446 1101 1452 1102
rect 1446 1097 1447 1101
rect 1451 1097 1452 1101
rect 1446 1096 1452 1097
rect 1494 1101 1500 1102
rect 1494 1097 1495 1101
rect 1499 1097 1500 1101
rect 1494 1096 1500 1097
rect 1542 1101 1548 1102
rect 1542 1097 1543 1101
rect 1547 1097 1548 1101
rect 1542 1096 1548 1097
rect 1590 1101 1596 1102
rect 1590 1097 1591 1101
rect 1595 1097 1596 1101
rect 1590 1096 1596 1097
rect 1622 1101 1628 1102
rect 1622 1097 1623 1101
rect 1627 1097 1628 1101
rect 1662 1099 1663 1103
rect 1667 1099 1668 1103
rect 1662 1098 1668 1099
rect 1622 1096 1628 1097
rect 214 1083 220 1084
rect 110 1081 116 1082
rect 110 1077 111 1081
rect 115 1077 116 1081
rect 214 1079 215 1083
rect 219 1079 220 1083
rect 214 1078 220 1079
rect 246 1083 252 1084
rect 246 1079 247 1083
rect 251 1079 252 1083
rect 246 1078 252 1079
rect 278 1083 284 1084
rect 278 1079 279 1083
rect 283 1079 284 1083
rect 278 1078 284 1079
rect 310 1083 316 1084
rect 310 1079 311 1083
rect 315 1079 316 1083
rect 310 1078 316 1079
rect 350 1083 356 1084
rect 350 1079 351 1083
rect 355 1079 356 1083
rect 350 1078 356 1079
rect 390 1083 396 1084
rect 390 1079 391 1083
rect 395 1079 396 1083
rect 390 1078 396 1079
rect 438 1083 444 1084
rect 438 1079 439 1083
rect 443 1079 444 1083
rect 438 1078 444 1079
rect 502 1083 508 1084
rect 502 1079 503 1083
rect 507 1079 508 1083
rect 502 1078 508 1079
rect 574 1083 580 1084
rect 574 1079 575 1083
rect 579 1079 580 1083
rect 574 1078 580 1079
rect 654 1083 660 1084
rect 654 1079 655 1083
rect 659 1079 660 1083
rect 654 1078 660 1079
rect 734 1083 740 1084
rect 734 1079 735 1083
rect 739 1079 740 1083
rect 734 1078 740 1079
rect 814 1083 820 1084
rect 814 1079 815 1083
rect 819 1079 820 1083
rect 814 1078 820 1079
rect 894 1083 900 1084
rect 894 1079 895 1083
rect 899 1079 900 1083
rect 894 1078 900 1079
rect 966 1083 972 1084
rect 966 1079 967 1083
rect 971 1079 972 1083
rect 966 1078 972 1079
rect 1038 1083 1044 1084
rect 1038 1079 1039 1083
rect 1043 1079 1044 1083
rect 1038 1078 1044 1079
rect 1110 1083 1116 1084
rect 1110 1079 1111 1083
rect 1115 1079 1116 1083
rect 1110 1078 1116 1079
rect 1174 1083 1180 1084
rect 1174 1079 1175 1083
rect 1179 1079 1180 1083
rect 1174 1078 1180 1079
rect 1238 1083 1244 1084
rect 1238 1079 1239 1083
rect 1243 1079 1244 1083
rect 1238 1078 1244 1079
rect 1302 1083 1308 1084
rect 1302 1079 1303 1083
rect 1307 1079 1308 1083
rect 1302 1078 1308 1079
rect 1358 1083 1364 1084
rect 1358 1079 1359 1083
rect 1363 1079 1364 1083
rect 1358 1078 1364 1079
rect 1414 1083 1420 1084
rect 1414 1079 1415 1083
rect 1419 1079 1420 1083
rect 1414 1078 1420 1079
rect 1462 1083 1468 1084
rect 1462 1079 1463 1083
rect 1467 1079 1468 1083
rect 1462 1078 1468 1079
rect 1502 1083 1508 1084
rect 1502 1079 1503 1083
rect 1507 1079 1508 1083
rect 1502 1078 1508 1079
rect 1550 1083 1556 1084
rect 1550 1079 1551 1083
rect 1555 1079 1556 1083
rect 1550 1078 1556 1079
rect 1590 1083 1596 1084
rect 1590 1079 1591 1083
rect 1595 1079 1596 1083
rect 1590 1078 1596 1079
rect 1622 1083 1628 1084
rect 1622 1079 1623 1083
rect 1627 1079 1628 1083
rect 1622 1078 1628 1079
rect 1662 1081 1668 1082
rect 110 1076 116 1077
rect 1662 1077 1663 1081
rect 1667 1077 1668 1081
rect 1662 1076 1668 1077
rect 214 1066 220 1067
rect 110 1064 116 1065
rect 110 1060 111 1064
rect 115 1060 116 1064
rect 214 1062 215 1066
rect 219 1062 220 1066
rect 214 1061 220 1062
rect 246 1066 252 1067
rect 246 1062 247 1066
rect 251 1062 252 1066
rect 246 1061 252 1062
rect 278 1066 284 1067
rect 278 1062 279 1066
rect 283 1062 284 1066
rect 278 1061 284 1062
rect 310 1066 316 1067
rect 310 1062 311 1066
rect 315 1062 316 1066
rect 310 1061 316 1062
rect 350 1066 356 1067
rect 350 1062 351 1066
rect 355 1062 356 1066
rect 350 1061 356 1062
rect 390 1066 396 1067
rect 390 1062 391 1066
rect 395 1062 396 1066
rect 390 1061 396 1062
rect 438 1066 444 1067
rect 438 1062 439 1066
rect 443 1062 444 1066
rect 438 1061 444 1062
rect 502 1066 508 1067
rect 502 1062 503 1066
rect 507 1062 508 1066
rect 502 1061 508 1062
rect 574 1066 580 1067
rect 574 1062 575 1066
rect 579 1062 580 1066
rect 574 1061 580 1062
rect 654 1066 660 1067
rect 654 1062 655 1066
rect 659 1062 660 1066
rect 654 1061 660 1062
rect 734 1066 740 1067
rect 734 1062 735 1066
rect 739 1062 740 1066
rect 734 1061 740 1062
rect 814 1066 820 1067
rect 814 1062 815 1066
rect 819 1062 820 1066
rect 814 1061 820 1062
rect 894 1066 900 1067
rect 894 1062 895 1066
rect 899 1062 900 1066
rect 894 1061 900 1062
rect 966 1066 972 1067
rect 966 1062 967 1066
rect 971 1062 972 1066
rect 966 1061 972 1062
rect 1038 1066 1044 1067
rect 1038 1062 1039 1066
rect 1043 1062 1044 1066
rect 1038 1061 1044 1062
rect 1110 1066 1116 1067
rect 1110 1062 1111 1066
rect 1115 1062 1116 1066
rect 1110 1061 1116 1062
rect 1174 1066 1180 1067
rect 1174 1062 1175 1066
rect 1179 1062 1180 1066
rect 1174 1061 1180 1062
rect 1238 1066 1244 1067
rect 1238 1062 1239 1066
rect 1243 1062 1244 1066
rect 1238 1061 1244 1062
rect 1302 1066 1308 1067
rect 1302 1062 1303 1066
rect 1307 1062 1308 1066
rect 1302 1061 1308 1062
rect 1358 1066 1364 1067
rect 1358 1062 1359 1066
rect 1363 1062 1364 1066
rect 1358 1061 1364 1062
rect 1414 1066 1420 1067
rect 1414 1062 1415 1066
rect 1419 1062 1420 1066
rect 1414 1061 1420 1062
rect 1462 1066 1468 1067
rect 1462 1062 1463 1066
rect 1467 1062 1468 1066
rect 1462 1061 1468 1062
rect 1502 1066 1508 1067
rect 1502 1062 1503 1066
rect 1507 1062 1508 1066
rect 1502 1061 1508 1062
rect 1550 1066 1556 1067
rect 1550 1062 1551 1066
rect 1555 1062 1556 1066
rect 1550 1061 1556 1062
rect 1590 1066 1596 1067
rect 1590 1062 1591 1066
rect 1595 1062 1596 1066
rect 1590 1061 1596 1062
rect 1622 1066 1628 1067
rect 1622 1062 1623 1066
rect 1627 1062 1628 1066
rect 1622 1061 1628 1062
rect 1662 1064 1668 1065
rect 110 1059 116 1060
rect 1662 1060 1663 1064
rect 1667 1060 1668 1064
rect 1662 1059 1668 1060
rect 110 1032 116 1033
rect 110 1028 111 1032
rect 115 1028 116 1032
rect 1662 1032 1668 1033
rect 110 1027 116 1028
rect 294 1030 300 1031
rect 294 1026 295 1030
rect 299 1026 300 1030
rect 294 1025 300 1026
rect 326 1030 332 1031
rect 326 1026 327 1030
rect 331 1026 332 1030
rect 326 1025 332 1026
rect 358 1030 364 1031
rect 358 1026 359 1030
rect 363 1026 364 1030
rect 358 1025 364 1026
rect 390 1030 396 1031
rect 390 1026 391 1030
rect 395 1026 396 1030
rect 390 1025 396 1026
rect 422 1030 428 1031
rect 422 1026 423 1030
rect 427 1026 428 1030
rect 422 1025 428 1026
rect 454 1030 460 1031
rect 454 1026 455 1030
rect 459 1026 460 1030
rect 454 1025 460 1026
rect 502 1030 508 1031
rect 502 1026 503 1030
rect 507 1026 508 1030
rect 502 1025 508 1026
rect 558 1030 564 1031
rect 558 1026 559 1030
rect 563 1026 564 1030
rect 558 1025 564 1026
rect 630 1030 636 1031
rect 630 1026 631 1030
rect 635 1026 636 1030
rect 630 1025 636 1026
rect 710 1030 716 1031
rect 710 1026 711 1030
rect 715 1026 716 1030
rect 710 1025 716 1026
rect 798 1030 804 1031
rect 798 1026 799 1030
rect 803 1026 804 1030
rect 798 1025 804 1026
rect 878 1030 884 1031
rect 878 1026 879 1030
rect 883 1026 884 1030
rect 878 1025 884 1026
rect 958 1030 964 1031
rect 958 1026 959 1030
rect 963 1026 964 1030
rect 958 1025 964 1026
rect 1030 1030 1036 1031
rect 1030 1026 1031 1030
rect 1035 1026 1036 1030
rect 1030 1025 1036 1026
rect 1094 1030 1100 1031
rect 1094 1026 1095 1030
rect 1099 1026 1100 1030
rect 1094 1025 1100 1026
rect 1158 1030 1164 1031
rect 1158 1026 1159 1030
rect 1163 1026 1164 1030
rect 1158 1025 1164 1026
rect 1222 1030 1228 1031
rect 1222 1026 1223 1030
rect 1227 1026 1228 1030
rect 1222 1025 1228 1026
rect 1278 1030 1284 1031
rect 1278 1026 1279 1030
rect 1283 1026 1284 1030
rect 1278 1025 1284 1026
rect 1334 1030 1340 1031
rect 1334 1026 1335 1030
rect 1339 1026 1340 1030
rect 1334 1025 1340 1026
rect 1382 1030 1388 1031
rect 1382 1026 1383 1030
rect 1387 1026 1388 1030
rect 1382 1025 1388 1026
rect 1430 1030 1436 1031
rect 1430 1026 1431 1030
rect 1435 1026 1436 1030
rect 1430 1025 1436 1026
rect 1478 1030 1484 1031
rect 1478 1026 1479 1030
rect 1483 1026 1484 1030
rect 1478 1025 1484 1026
rect 1534 1030 1540 1031
rect 1534 1026 1535 1030
rect 1539 1026 1540 1030
rect 1534 1025 1540 1026
rect 1590 1030 1596 1031
rect 1590 1026 1591 1030
rect 1595 1026 1596 1030
rect 1590 1025 1596 1026
rect 1622 1030 1628 1031
rect 1622 1026 1623 1030
rect 1627 1026 1628 1030
rect 1662 1028 1663 1032
rect 1667 1028 1668 1032
rect 1662 1027 1668 1028
rect 1622 1025 1628 1026
rect 110 1015 116 1016
rect 110 1011 111 1015
rect 115 1011 116 1015
rect 1662 1015 1668 1016
rect 110 1010 116 1011
rect 294 1013 300 1014
rect 294 1009 295 1013
rect 299 1009 300 1013
rect 294 1008 300 1009
rect 326 1013 332 1014
rect 326 1009 327 1013
rect 331 1009 332 1013
rect 326 1008 332 1009
rect 358 1013 364 1014
rect 358 1009 359 1013
rect 363 1009 364 1013
rect 358 1008 364 1009
rect 390 1013 396 1014
rect 390 1009 391 1013
rect 395 1009 396 1013
rect 390 1008 396 1009
rect 422 1013 428 1014
rect 422 1009 423 1013
rect 427 1009 428 1013
rect 422 1008 428 1009
rect 454 1013 460 1014
rect 454 1009 455 1013
rect 459 1009 460 1013
rect 454 1008 460 1009
rect 502 1013 508 1014
rect 502 1009 503 1013
rect 507 1009 508 1013
rect 502 1008 508 1009
rect 558 1013 564 1014
rect 558 1009 559 1013
rect 563 1009 564 1013
rect 558 1008 564 1009
rect 630 1013 636 1014
rect 630 1009 631 1013
rect 635 1009 636 1013
rect 630 1008 636 1009
rect 710 1013 716 1014
rect 710 1009 711 1013
rect 715 1009 716 1013
rect 710 1008 716 1009
rect 798 1013 804 1014
rect 798 1009 799 1013
rect 803 1009 804 1013
rect 798 1008 804 1009
rect 878 1013 884 1014
rect 878 1009 879 1013
rect 883 1009 884 1013
rect 878 1008 884 1009
rect 958 1013 964 1014
rect 958 1009 959 1013
rect 963 1009 964 1013
rect 958 1008 964 1009
rect 1030 1013 1036 1014
rect 1030 1009 1031 1013
rect 1035 1009 1036 1013
rect 1030 1008 1036 1009
rect 1094 1013 1100 1014
rect 1094 1009 1095 1013
rect 1099 1009 1100 1013
rect 1094 1008 1100 1009
rect 1158 1013 1164 1014
rect 1158 1009 1159 1013
rect 1163 1009 1164 1013
rect 1158 1008 1164 1009
rect 1222 1013 1228 1014
rect 1222 1009 1223 1013
rect 1227 1009 1228 1013
rect 1222 1008 1228 1009
rect 1278 1013 1284 1014
rect 1278 1009 1279 1013
rect 1283 1009 1284 1013
rect 1278 1008 1284 1009
rect 1334 1013 1340 1014
rect 1334 1009 1335 1013
rect 1339 1009 1340 1013
rect 1334 1008 1340 1009
rect 1382 1013 1388 1014
rect 1382 1009 1383 1013
rect 1387 1009 1388 1013
rect 1382 1008 1388 1009
rect 1430 1013 1436 1014
rect 1430 1009 1431 1013
rect 1435 1009 1436 1013
rect 1430 1008 1436 1009
rect 1478 1013 1484 1014
rect 1478 1009 1479 1013
rect 1483 1009 1484 1013
rect 1478 1008 1484 1009
rect 1534 1013 1540 1014
rect 1534 1009 1535 1013
rect 1539 1009 1540 1013
rect 1534 1008 1540 1009
rect 1590 1013 1596 1014
rect 1590 1009 1591 1013
rect 1595 1009 1596 1013
rect 1590 1008 1596 1009
rect 1622 1013 1628 1014
rect 1622 1009 1623 1013
rect 1627 1009 1628 1013
rect 1662 1011 1663 1015
rect 1667 1011 1668 1015
rect 1662 1010 1668 1011
rect 1622 1008 1628 1009
rect 246 999 252 1000
rect 110 997 116 998
rect 110 993 111 997
rect 115 993 116 997
rect 246 995 247 999
rect 251 995 252 999
rect 246 994 252 995
rect 278 999 284 1000
rect 278 995 279 999
rect 283 995 284 999
rect 278 994 284 995
rect 310 999 316 1000
rect 310 995 311 999
rect 315 995 316 999
rect 310 994 316 995
rect 342 999 348 1000
rect 342 995 343 999
rect 347 995 348 999
rect 342 994 348 995
rect 382 999 388 1000
rect 382 995 383 999
rect 387 995 388 999
rect 382 994 388 995
rect 422 999 428 1000
rect 422 995 423 999
rect 427 995 428 999
rect 422 994 428 995
rect 478 999 484 1000
rect 478 995 479 999
rect 483 995 484 999
rect 478 994 484 995
rect 542 999 548 1000
rect 542 995 543 999
rect 547 995 548 999
rect 542 994 548 995
rect 614 999 620 1000
rect 614 995 615 999
rect 619 995 620 999
rect 614 994 620 995
rect 686 999 692 1000
rect 686 995 687 999
rect 691 995 692 999
rect 686 994 692 995
rect 758 999 764 1000
rect 758 995 759 999
rect 763 995 764 999
rect 758 994 764 995
rect 830 999 836 1000
rect 830 995 831 999
rect 835 995 836 999
rect 830 994 836 995
rect 902 999 908 1000
rect 902 995 903 999
rect 907 995 908 999
rect 902 994 908 995
rect 966 999 972 1000
rect 966 995 967 999
rect 971 995 972 999
rect 966 994 972 995
rect 1030 999 1036 1000
rect 1030 995 1031 999
rect 1035 995 1036 999
rect 1030 994 1036 995
rect 1094 999 1100 1000
rect 1094 995 1095 999
rect 1099 995 1100 999
rect 1094 994 1100 995
rect 1158 999 1164 1000
rect 1158 995 1159 999
rect 1163 995 1164 999
rect 1158 994 1164 995
rect 1222 999 1228 1000
rect 1222 995 1223 999
rect 1227 995 1228 999
rect 1222 994 1228 995
rect 1286 999 1292 1000
rect 1286 995 1287 999
rect 1291 995 1292 999
rect 1286 994 1292 995
rect 1342 999 1348 1000
rect 1342 995 1343 999
rect 1347 995 1348 999
rect 1342 994 1348 995
rect 1398 999 1404 1000
rect 1398 995 1399 999
rect 1403 995 1404 999
rect 1398 994 1404 995
rect 1446 999 1452 1000
rect 1446 995 1447 999
rect 1451 995 1452 999
rect 1446 994 1452 995
rect 1494 999 1500 1000
rect 1494 995 1495 999
rect 1499 995 1500 999
rect 1494 994 1500 995
rect 1542 999 1548 1000
rect 1542 995 1543 999
rect 1547 995 1548 999
rect 1542 994 1548 995
rect 1590 999 1596 1000
rect 1590 995 1591 999
rect 1595 995 1596 999
rect 1590 994 1596 995
rect 1622 999 1628 1000
rect 1622 995 1623 999
rect 1627 995 1628 999
rect 1622 994 1628 995
rect 1662 997 1668 998
rect 110 992 116 993
rect 1662 993 1663 997
rect 1667 993 1668 997
rect 1662 992 1668 993
rect 246 982 252 983
rect 110 980 116 981
rect 110 976 111 980
rect 115 976 116 980
rect 246 978 247 982
rect 251 978 252 982
rect 246 977 252 978
rect 278 982 284 983
rect 278 978 279 982
rect 283 978 284 982
rect 278 977 284 978
rect 310 982 316 983
rect 310 978 311 982
rect 315 978 316 982
rect 310 977 316 978
rect 342 982 348 983
rect 342 978 343 982
rect 347 978 348 982
rect 342 977 348 978
rect 382 982 388 983
rect 382 978 383 982
rect 387 978 388 982
rect 382 977 388 978
rect 422 982 428 983
rect 422 978 423 982
rect 427 978 428 982
rect 422 977 428 978
rect 478 982 484 983
rect 478 978 479 982
rect 483 978 484 982
rect 478 977 484 978
rect 542 982 548 983
rect 542 978 543 982
rect 547 978 548 982
rect 542 977 548 978
rect 614 982 620 983
rect 614 978 615 982
rect 619 978 620 982
rect 614 977 620 978
rect 686 982 692 983
rect 686 978 687 982
rect 691 978 692 982
rect 686 977 692 978
rect 758 982 764 983
rect 758 978 759 982
rect 763 978 764 982
rect 758 977 764 978
rect 830 982 836 983
rect 830 978 831 982
rect 835 978 836 982
rect 830 977 836 978
rect 902 982 908 983
rect 902 978 903 982
rect 907 978 908 982
rect 902 977 908 978
rect 966 982 972 983
rect 966 978 967 982
rect 971 978 972 982
rect 966 977 972 978
rect 1030 982 1036 983
rect 1030 978 1031 982
rect 1035 978 1036 982
rect 1030 977 1036 978
rect 1094 982 1100 983
rect 1094 978 1095 982
rect 1099 978 1100 982
rect 1094 977 1100 978
rect 1158 982 1164 983
rect 1158 978 1159 982
rect 1163 978 1164 982
rect 1158 977 1164 978
rect 1222 982 1228 983
rect 1222 978 1223 982
rect 1227 978 1228 982
rect 1222 977 1228 978
rect 1286 982 1292 983
rect 1286 978 1287 982
rect 1291 978 1292 982
rect 1286 977 1292 978
rect 1342 982 1348 983
rect 1342 978 1343 982
rect 1347 978 1348 982
rect 1342 977 1348 978
rect 1398 982 1404 983
rect 1398 978 1399 982
rect 1403 978 1404 982
rect 1398 977 1404 978
rect 1446 982 1452 983
rect 1446 978 1447 982
rect 1451 978 1452 982
rect 1446 977 1452 978
rect 1494 982 1500 983
rect 1494 978 1495 982
rect 1499 978 1500 982
rect 1494 977 1500 978
rect 1542 982 1548 983
rect 1542 978 1543 982
rect 1547 978 1548 982
rect 1542 977 1548 978
rect 1590 982 1596 983
rect 1590 978 1591 982
rect 1595 978 1596 982
rect 1590 977 1596 978
rect 1622 982 1628 983
rect 1622 978 1623 982
rect 1627 978 1628 982
rect 1622 977 1628 978
rect 1662 980 1668 981
rect 110 975 116 976
rect 1662 976 1663 980
rect 1667 976 1668 980
rect 1662 975 1668 976
rect 110 952 116 953
rect 110 948 111 952
rect 115 948 116 952
rect 1662 952 1668 953
rect 110 947 116 948
rect 166 950 172 951
rect 166 946 167 950
rect 171 946 172 950
rect 166 945 172 946
rect 198 950 204 951
rect 198 946 199 950
rect 203 946 204 950
rect 198 945 204 946
rect 238 950 244 951
rect 238 946 239 950
rect 243 946 244 950
rect 238 945 244 946
rect 286 950 292 951
rect 286 946 287 950
rect 291 946 292 950
rect 286 945 292 946
rect 342 950 348 951
rect 342 946 343 950
rect 347 946 348 950
rect 342 945 348 946
rect 406 950 412 951
rect 406 946 407 950
rect 411 946 412 950
rect 406 945 412 946
rect 470 950 476 951
rect 470 946 471 950
rect 475 946 476 950
rect 470 945 476 946
rect 534 950 540 951
rect 534 946 535 950
rect 539 946 540 950
rect 534 945 540 946
rect 598 950 604 951
rect 598 946 599 950
rect 603 946 604 950
rect 598 945 604 946
rect 662 950 668 951
rect 662 946 663 950
rect 667 946 668 950
rect 662 945 668 946
rect 726 950 732 951
rect 726 946 727 950
rect 731 946 732 950
rect 726 945 732 946
rect 790 950 796 951
rect 790 946 791 950
rect 795 946 796 950
rect 790 945 796 946
rect 846 950 852 951
rect 846 946 847 950
rect 851 946 852 950
rect 846 945 852 946
rect 910 950 916 951
rect 910 946 911 950
rect 915 946 916 950
rect 910 945 916 946
rect 974 950 980 951
rect 974 946 975 950
rect 979 946 980 950
rect 974 945 980 946
rect 1038 950 1044 951
rect 1038 946 1039 950
rect 1043 946 1044 950
rect 1038 945 1044 946
rect 1102 950 1108 951
rect 1102 946 1103 950
rect 1107 946 1108 950
rect 1102 945 1108 946
rect 1166 950 1172 951
rect 1166 946 1167 950
rect 1171 946 1172 950
rect 1166 945 1172 946
rect 1230 950 1236 951
rect 1230 946 1231 950
rect 1235 946 1236 950
rect 1230 945 1236 946
rect 1286 950 1292 951
rect 1286 946 1287 950
rect 1291 946 1292 950
rect 1286 945 1292 946
rect 1342 950 1348 951
rect 1342 946 1343 950
rect 1347 946 1348 950
rect 1342 945 1348 946
rect 1390 950 1396 951
rect 1390 946 1391 950
rect 1395 946 1396 950
rect 1390 945 1396 946
rect 1430 950 1436 951
rect 1430 946 1431 950
rect 1435 946 1436 950
rect 1430 945 1436 946
rect 1470 950 1476 951
rect 1470 946 1471 950
rect 1475 946 1476 950
rect 1470 945 1476 946
rect 1510 950 1516 951
rect 1510 946 1511 950
rect 1515 946 1516 950
rect 1510 945 1516 946
rect 1550 950 1556 951
rect 1550 946 1551 950
rect 1555 946 1556 950
rect 1550 945 1556 946
rect 1590 950 1596 951
rect 1590 946 1591 950
rect 1595 946 1596 950
rect 1590 945 1596 946
rect 1622 950 1628 951
rect 1622 946 1623 950
rect 1627 946 1628 950
rect 1662 948 1663 952
rect 1667 948 1668 952
rect 1662 947 1668 948
rect 1622 945 1628 946
rect 110 935 116 936
rect 110 931 111 935
rect 115 931 116 935
rect 1662 935 1668 936
rect 110 930 116 931
rect 166 933 172 934
rect 166 929 167 933
rect 171 929 172 933
rect 166 928 172 929
rect 198 933 204 934
rect 198 929 199 933
rect 203 929 204 933
rect 198 928 204 929
rect 238 933 244 934
rect 238 929 239 933
rect 243 929 244 933
rect 238 928 244 929
rect 286 933 292 934
rect 286 929 287 933
rect 291 929 292 933
rect 286 928 292 929
rect 342 933 348 934
rect 342 929 343 933
rect 347 929 348 933
rect 342 928 348 929
rect 406 933 412 934
rect 406 929 407 933
rect 411 929 412 933
rect 406 928 412 929
rect 470 933 476 934
rect 470 929 471 933
rect 475 929 476 933
rect 470 928 476 929
rect 534 933 540 934
rect 534 929 535 933
rect 539 929 540 933
rect 534 928 540 929
rect 598 933 604 934
rect 598 929 599 933
rect 603 929 604 933
rect 598 928 604 929
rect 662 933 668 934
rect 662 929 663 933
rect 667 929 668 933
rect 662 928 668 929
rect 726 933 732 934
rect 726 929 727 933
rect 731 929 732 933
rect 726 928 732 929
rect 790 933 796 934
rect 790 929 791 933
rect 795 929 796 933
rect 790 928 796 929
rect 846 933 852 934
rect 846 929 847 933
rect 851 929 852 933
rect 846 928 852 929
rect 910 933 916 934
rect 910 929 911 933
rect 915 929 916 933
rect 910 928 916 929
rect 974 933 980 934
rect 974 929 975 933
rect 979 929 980 933
rect 974 928 980 929
rect 1038 933 1044 934
rect 1038 929 1039 933
rect 1043 929 1044 933
rect 1038 928 1044 929
rect 1102 933 1108 934
rect 1102 929 1103 933
rect 1107 929 1108 933
rect 1102 928 1108 929
rect 1166 933 1172 934
rect 1166 929 1167 933
rect 1171 929 1172 933
rect 1166 928 1172 929
rect 1230 933 1236 934
rect 1230 929 1231 933
rect 1235 929 1236 933
rect 1230 928 1236 929
rect 1286 933 1292 934
rect 1286 929 1287 933
rect 1291 929 1292 933
rect 1286 928 1292 929
rect 1342 933 1348 934
rect 1342 929 1343 933
rect 1347 929 1348 933
rect 1342 928 1348 929
rect 1390 933 1396 934
rect 1390 929 1391 933
rect 1395 929 1396 933
rect 1390 928 1396 929
rect 1430 933 1436 934
rect 1430 929 1431 933
rect 1435 929 1436 933
rect 1430 928 1436 929
rect 1470 933 1476 934
rect 1470 929 1471 933
rect 1475 929 1476 933
rect 1470 928 1476 929
rect 1510 933 1516 934
rect 1510 929 1511 933
rect 1515 929 1516 933
rect 1510 928 1516 929
rect 1550 933 1556 934
rect 1550 929 1551 933
rect 1555 929 1556 933
rect 1550 928 1556 929
rect 1590 933 1596 934
rect 1590 929 1591 933
rect 1595 929 1596 933
rect 1590 928 1596 929
rect 1622 933 1628 934
rect 1622 929 1623 933
rect 1627 929 1628 933
rect 1662 931 1663 935
rect 1667 931 1668 935
rect 1662 930 1668 931
rect 1622 928 1628 929
rect 134 915 140 916
rect 110 913 116 914
rect 110 909 111 913
rect 115 909 116 913
rect 134 911 135 915
rect 139 911 140 915
rect 134 910 140 911
rect 166 915 172 916
rect 166 911 167 915
rect 171 911 172 915
rect 166 910 172 911
rect 206 915 212 916
rect 206 911 207 915
rect 211 911 212 915
rect 206 910 212 911
rect 270 915 276 916
rect 270 911 271 915
rect 275 911 276 915
rect 270 910 276 911
rect 334 915 340 916
rect 334 911 335 915
rect 339 911 340 915
rect 334 910 340 911
rect 406 915 412 916
rect 406 911 407 915
rect 411 911 412 915
rect 406 910 412 911
rect 470 915 476 916
rect 470 911 471 915
rect 475 911 476 915
rect 470 910 476 911
rect 534 915 540 916
rect 534 911 535 915
rect 539 911 540 915
rect 534 910 540 911
rect 590 915 596 916
rect 590 911 591 915
rect 595 911 596 915
rect 590 910 596 911
rect 646 915 652 916
rect 646 911 647 915
rect 651 911 652 915
rect 646 910 652 911
rect 702 915 708 916
rect 702 911 703 915
rect 707 911 708 915
rect 702 910 708 911
rect 750 915 756 916
rect 750 911 751 915
rect 755 911 756 915
rect 750 910 756 911
rect 798 915 804 916
rect 798 911 799 915
rect 803 911 804 915
rect 798 910 804 911
rect 846 915 852 916
rect 846 911 847 915
rect 851 911 852 915
rect 846 910 852 911
rect 902 915 908 916
rect 902 911 903 915
rect 907 911 908 915
rect 902 910 908 911
rect 958 915 964 916
rect 958 911 959 915
rect 963 911 964 915
rect 958 910 964 911
rect 1022 915 1028 916
rect 1022 911 1023 915
rect 1027 911 1028 915
rect 1022 910 1028 911
rect 1086 915 1092 916
rect 1086 911 1087 915
rect 1091 911 1092 915
rect 1086 910 1092 911
rect 1142 915 1148 916
rect 1142 911 1143 915
rect 1147 911 1148 915
rect 1142 910 1148 911
rect 1198 915 1204 916
rect 1198 911 1199 915
rect 1203 911 1204 915
rect 1198 910 1204 911
rect 1254 915 1260 916
rect 1254 911 1255 915
rect 1259 911 1260 915
rect 1254 910 1260 911
rect 1318 915 1324 916
rect 1318 911 1319 915
rect 1323 911 1324 915
rect 1318 910 1324 911
rect 1382 915 1388 916
rect 1382 911 1383 915
rect 1387 911 1388 915
rect 1382 910 1388 911
rect 1662 913 1668 914
rect 110 908 116 909
rect 1662 909 1663 913
rect 1667 909 1668 913
rect 1662 908 1668 909
rect 134 898 140 899
rect 110 896 116 897
rect 110 892 111 896
rect 115 892 116 896
rect 134 894 135 898
rect 139 894 140 898
rect 134 893 140 894
rect 166 898 172 899
rect 166 894 167 898
rect 171 894 172 898
rect 166 893 172 894
rect 206 898 212 899
rect 206 894 207 898
rect 211 894 212 898
rect 206 893 212 894
rect 270 898 276 899
rect 270 894 271 898
rect 275 894 276 898
rect 270 893 276 894
rect 334 898 340 899
rect 334 894 335 898
rect 339 894 340 898
rect 334 893 340 894
rect 406 898 412 899
rect 406 894 407 898
rect 411 894 412 898
rect 406 893 412 894
rect 470 898 476 899
rect 470 894 471 898
rect 475 894 476 898
rect 470 893 476 894
rect 534 898 540 899
rect 534 894 535 898
rect 539 894 540 898
rect 534 893 540 894
rect 590 898 596 899
rect 590 894 591 898
rect 595 894 596 898
rect 590 893 596 894
rect 646 898 652 899
rect 646 894 647 898
rect 651 894 652 898
rect 646 893 652 894
rect 702 898 708 899
rect 702 894 703 898
rect 707 894 708 898
rect 702 893 708 894
rect 750 898 756 899
rect 750 894 751 898
rect 755 894 756 898
rect 750 893 756 894
rect 798 898 804 899
rect 798 894 799 898
rect 803 894 804 898
rect 798 893 804 894
rect 846 898 852 899
rect 846 894 847 898
rect 851 894 852 898
rect 846 893 852 894
rect 902 898 908 899
rect 902 894 903 898
rect 907 894 908 898
rect 902 893 908 894
rect 958 898 964 899
rect 958 894 959 898
rect 963 894 964 898
rect 958 893 964 894
rect 1022 898 1028 899
rect 1022 894 1023 898
rect 1027 894 1028 898
rect 1022 893 1028 894
rect 1086 898 1092 899
rect 1086 894 1087 898
rect 1091 894 1092 898
rect 1086 893 1092 894
rect 1142 898 1148 899
rect 1142 894 1143 898
rect 1147 894 1148 898
rect 1142 893 1148 894
rect 1198 898 1204 899
rect 1198 894 1199 898
rect 1203 894 1204 898
rect 1198 893 1204 894
rect 1254 898 1260 899
rect 1254 894 1255 898
rect 1259 894 1260 898
rect 1254 893 1260 894
rect 1318 898 1324 899
rect 1318 894 1319 898
rect 1323 894 1324 898
rect 1318 893 1324 894
rect 1382 898 1388 899
rect 1382 894 1383 898
rect 1387 894 1388 898
rect 1382 893 1388 894
rect 1662 896 1668 897
rect 110 891 116 892
rect 1662 892 1663 896
rect 1667 892 1668 896
rect 1662 891 1668 892
rect 110 864 116 865
rect 110 860 111 864
rect 115 860 116 864
rect 1662 864 1668 865
rect 110 859 116 860
rect 134 862 140 863
rect 134 858 135 862
rect 139 858 140 862
rect 134 857 140 858
rect 166 862 172 863
rect 166 858 167 862
rect 171 858 172 862
rect 166 857 172 858
rect 206 862 212 863
rect 206 858 207 862
rect 211 858 212 862
rect 206 857 212 858
rect 270 862 276 863
rect 270 858 271 862
rect 275 858 276 862
rect 270 857 276 858
rect 334 862 340 863
rect 334 858 335 862
rect 339 858 340 862
rect 334 857 340 858
rect 406 862 412 863
rect 406 858 407 862
rect 411 858 412 862
rect 406 857 412 858
rect 470 862 476 863
rect 470 858 471 862
rect 475 858 476 862
rect 470 857 476 858
rect 534 862 540 863
rect 534 858 535 862
rect 539 858 540 862
rect 534 857 540 858
rect 598 862 604 863
rect 598 858 599 862
rect 603 858 604 862
rect 598 857 604 858
rect 654 862 660 863
rect 654 858 655 862
rect 659 858 660 862
rect 654 857 660 858
rect 702 862 708 863
rect 702 858 703 862
rect 707 858 708 862
rect 702 857 708 858
rect 750 862 756 863
rect 750 858 751 862
rect 755 858 756 862
rect 750 857 756 858
rect 798 862 804 863
rect 798 858 799 862
rect 803 858 804 862
rect 798 857 804 858
rect 846 862 852 863
rect 846 858 847 862
rect 851 858 852 862
rect 846 857 852 858
rect 902 862 908 863
rect 902 858 903 862
rect 907 858 908 862
rect 902 857 908 858
rect 966 862 972 863
rect 966 858 967 862
rect 971 858 972 862
rect 966 857 972 858
rect 1038 862 1044 863
rect 1038 858 1039 862
rect 1043 858 1044 862
rect 1038 857 1044 858
rect 1102 862 1108 863
rect 1102 858 1103 862
rect 1107 858 1108 862
rect 1102 857 1108 858
rect 1166 862 1172 863
rect 1166 858 1167 862
rect 1171 858 1172 862
rect 1166 857 1172 858
rect 1230 862 1236 863
rect 1230 858 1231 862
rect 1235 858 1236 862
rect 1230 857 1236 858
rect 1286 862 1292 863
rect 1286 858 1287 862
rect 1291 858 1292 862
rect 1286 857 1292 858
rect 1342 862 1348 863
rect 1342 858 1343 862
rect 1347 858 1348 862
rect 1342 857 1348 858
rect 1398 862 1404 863
rect 1398 858 1399 862
rect 1403 858 1404 862
rect 1398 857 1404 858
rect 1462 862 1468 863
rect 1462 858 1463 862
rect 1467 858 1468 862
rect 1662 860 1663 864
rect 1667 860 1668 864
rect 1662 859 1668 860
rect 1462 857 1468 858
rect 110 847 116 848
rect 110 843 111 847
rect 115 843 116 847
rect 1662 847 1668 848
rect 110 842 116 843
rect 134 845 140 846
rect 134 841 135 845
rect 139 841 140 845
rect 134 840 140 841
rect 166 845 172 846
rect 166 841 167 845
rect 171 841 172 845
rect 166 840 172 841
rect 206 845 212 846
rect 206 841 207 845
rect 211 841 212 845
rect 206 840 212 841
rect 270 845 276 846
rect 270 841 271 845
rect 275 841 276 845
rect 270 840 276 841
rect 334 845 340 846
rect 334 841 335 845
rect 339 841 340 845
rect 334 840 340 841
rect 406 845 412 846
rect 406 841 407 845
rect 411 841 412 845
rect 406 840 412 841
rect 470 845 476 846
rect 470 841 471 845
rect 475 841 476 845
rect 470 840 476 841
rect 534 845 540 846
rect 534 841 535 845
rect 539 841 540 845
rect 534 840 540 841
rect 598 845 604 846
rect 598 841 599 845
rect 603 841 604 845
rect 598 840 604 841
rect 654 845 660 846
rect 654 841 655 845
rect 659 841 660 845
rect 654 840 660 841
rect 702 845 708 846
rect 702 841 703 845
rect 707 841 708 845
rect 702 840 708 841
rect 750 845 756 846
rect 750 841 751 845
rect 755 841 756 845
rect 750 840 756 841
rect 798 845 804 846
rect 798 841 799 845
rect 803 841 804 845
rect 798 840 804 841
rect 846 845 852 846
rect 846 841 847 845
rect 851 841 852 845
rect 846 840 852 841
rect 902 845 908 846
rect 902 841 903 845
rect 907 841 908 845
rect 902 840 908 841
rect 966 845 972 846
rect 966 841 967 845
rect 971 841 972 845
rect 966 840 972 841
rect 1038 845 1044 846
rect 1038 841 1039 845
rect 1043 841 1044 845
rect 1038 840 1044 841
rect 1102 845 1108 846
rect 1102 841 1103 845
rect 1107 841 1108 845
rect 1102 840 1108 841
rect 1166 845 1172 846
rect 1166 841 1167 845
rect 1171 841 1172 845
rect 1166 840 1172 841
rect 1230 845 1236 846
rect 1230 841 1231 845
rect 1235 841 1236 845
rect 1230 840 1236 841
rect 1286 845 1292 846
rect 1286 841 1287 845
rect 1291 841 1292 845
rect 1286 840 1292 841
rect 1342 845 1348 846
rect 1342 841 1343 845
rect 1347 841 1348 845
rect 1342 840 1348 841
rect 1398 845 1404 846
rect 1398 841 1399 845
rect 1403 841 1404 845
rect 1398 840 1404 841
rect 1462 845 1468 846
rect 1462 841 1463 845
rect 1467 841 1468 845
rect 1662 843 1663 847
rect 1667 843 1668 847
rect 1662 842 1668 843
rect 1462 840 1468 841
rect 134 831 140 832
rect 110 829 116 830
rect 110 825 111 829
rect 115 825 116 829
rect 134 827 135 831
rect 139 827 140 831
rect 134 826 140 827
rect 166 831 172 832
rect 166 827 167 831
rect 171 827 172 831
rect 166 826 172 827
rect 214 831 220 832
rect 214 827 215 831
rect 219 827 220 831
rect 214 826 220 827
rect 278 831 284 832
rect 278 827 279 831
rect 283 827 284 831
rect 278 826 284 827
rect 342 831 348 832
rect 342 827 343 831
rect 347 827 348 831
rect 342 826 348 827
rect 414 831 420 832
rect 414 827 415 831
rect 419 827 420 831
rect 414 826 420 827
rect 478 831 484 832
rect 478 827 479 831
rect 483 827 484 831
rect 478 826 484 827
rect 542 831 548 832
rect 542 827 543 831
rect 547 827 548 831
rect 542 826 548 827
rect 606 831 612 832
rect 606 827 607 831
rect 611 827 612 831
rect 606 826 612 827
rect 670 831 676 832
rect 670 827 671 831
rect 675 827 676 831
rect 670 826 676 827
rect 734 831 740 832
rect 734 827 735 831
rect 739 827 740 831
rect 734 826 740 827
rect 790 831 796 832
rect 790 827 791 831
rect 795 827 796 831
rect 790 826 796 827
rect 846 831 852 832
rect 846 827 847 831
rect 851 827 852 831
rect 846 826 852 827
rect 910 831 916 832
rect 910 827 911 831
rect 915 827 916 831
rect 910 826 916 827
rect 974 831 980 832
rect 974 827 975 831
rect 979 827 980 831
rect 974 826 980 827
rect 1038 831 1044 832
rect 1038 827 1039 831
rect 1043 827 1044 831
rect 1038 826 1044 827
rect 1110 831 1116 832
rect 1110 827 1111 831
rect 1115 827 1116 831
rect 1110 826 1116 827
rect 1182 831 1188 832
rect 1182 827 1183 831
rect 1187 827 1188 831
rect 1182 826 1188 827
rect 1246 831 1252 832
rect 1246 827 1247 831
rect 1251 827 1252 831
rect 1246 826 1252 827
rect 1310 831 1316 832
rect 1310 827 1311 831
rect 1315 827 1316 831
rect 1310 826 1316 827
rect 1366 831 1372 832
rect 1366 827 1367 831
rect 1371 827 1372 831
rect 1366 826 1372 827
rect 1422 831 1428 832
rect 1422 827 1423 831
rect 1427 827 1428 831
rect 1422 826 1428 827
rect 1478 831 1484 832
rect 1478 827 1479 831
rect 1483 827 1484 831
rect 1478 826 1484 827
rect 1534 831 1540 832
rect 1534 827 1535 831
rect 1539 827 1540 831
rect 1534 826 1540 827
rect 1590 831 1596 832
rect 1590 827 1591 831
rect 1595 827 1596 831
rect 1590 826 1596 827
rect 1662 829 1668 830
rect 110 824 116 825
rect 1662 825 1663 829
rect 1667 825 1668 829
rect 1662 824 1668 825
rect 134 814 140 815
rect 110 812 116 813
rect 110 808 111 812
rect 115 808 116 812
rect 134 810 135 814
rect 139 810 140 814
rect 134 809 140 810
rect 166 814 172 815
rect 166 810 167 814
rect 171 810 172 814
rect 166 809 172 810
rect 214 814 220 815
rect 214 810 215 814
rect 219 810 220 814
rect 214 809 220 810
rect 278 814 284 815
rect 278 810 279 814
rect 283 810 284 814
rect 278 809 284 810
rect 342 814 348 815
rect 342 810 343 814
rect 347 810 348 814
rect 342 809 348 810
rect 414 814 420 815
rect 414 810 415 814
rect 419 810 420 814
rect 414 809 420 810
rect 478 814 484 815
rect 478 810 479 814
rect 483 810 484 814
rect 478 809 484 810
rect 542 814 548 815
rect 542 810 543 814
rect 547 810 548 814
rect 542 809 548 810
rect 606 814 612 815
rect 606 810 607 814
rect 611 810 612 814
rect 606 809 612 810
rect 670 814 676 815
rect 670 810 671 814
rect 675 810 676 814
rect 670 809 676 810
rect 734 814 740 815
rect 734 810 735 814
rect 739 810 740 814
rect 734 809 740 810
rect 790 814 796 815
rect 790 810 791 814
rect 795 810 796 814
rect 790 809 796 810
rect 846 814 852 815
rect 846 810 847 814
rect 851 810 852 814
rect 846 809 852 810
rect 910 814 916 815
rect 910 810 911 814
rect 915 810 916 814
rect 910 809 916 810
rect 974 814 980 815
rect 974 810 975 814
rect 979 810 980 814
rect 974 809 980 810
rect 1038 814 1044 815
rect 1038 810 1039 814
rect 1043 810 1044 814
rect 1038 809 1044 810
rect 1110 814 1116 815
rect 1110 810 1111 814
rect 1115 810 1116 814
rect 1110 809 1116 810
rect 1182 814 1188 815
rect 1182 810 1183 814
rect 1187 810 1188 814
rect 1182 809 1188 810
rect 1246 814 1252 815
rect 1246 810 1247 814
rect 1251 810 1252 814
rect 1246 809 1252 810
rect 1310 814 1316 815
rect 1310 810 1311 814
rect 1315 810 1316 814
rect 1310 809 1316 810
rect 1366 814 1372 815
rect 1366 810 1367 814
rect 1371 810 1372 814
rect 1366 809 1372 810
rect 1422 814 1428 815
rect 1422 810 1423 814
rect 1427 810 1428 814
rect 1422 809 1428 810
rect 1478 814 1484 815
rect 1478 810 1479 814
rect 1483 810 1484 814
rect 1478 809 1484 810
rect 1534 814 1540 815
rect 1534 810 1535 814
rect 1539 810 1540 814
rect 1534 809 1540 810
rect 1590 814 1596 815
rect 1590 810 1591 814
rect 1595 810 1596 814
rect 1590 809 1596 810
rect 1662 812 1668 813
rect 110 807 116 808
rect 1662 808 1663 812
rect 1667 808 1668 812
rect 1662 807 1668 808
rect 110 780 116 781
rect 110 776 111 780
rect 115 776 116 780
rect 1662 780 1668 781
rect 110 775 116 776
rect 134 778 140 779
rect 134 774 135 778
rect 139 774 140 778
rect 134 773 140 774
rect 174 778 180 779
rect 174 774 175 778
rect 179 774 180 778
rect 174 773 180 774
rect 230 778 236 779
rect 230 774 231 778
rect 235 774 236 778
rect 230 773 236 774
rect 294 778 300 779
rect 294 774 295 778
rect 299 774 300 778
rect 294 773 300 774
rect 366 778 372 779
rect 366 774 367 778
rect 371 774 372 778
rect 366 773 372 774
rect 446 778 452 779
rect 446 774 447 778
rect 451 774 452 778
rect 446 773 452 774
rect 526 778 532 779
rect 526 774 527 778
rect 531 774 532 778
rect 526 773 532 774
rect 614 778 620 779
rect 614 774 615 778
rect 619 774 620 778
rect 614 773 620 774
rect 702 778 708 779
rect 702 774 703 778
rect 707 774 708 778
rect 702 773 708 774
rect 790 778 796 779
rect 790 774 791 778
rect 795 774 796 778
rect 790 773 796 774
rect 870 778 876 779
rect 870 774 871 778
rect 875 774 876 778
rect 870 773 876 774
rect 950 778 956 779
rect 950 774 951 778
rect 955 774 956 778
rect 950 773 956 774
rect 1022 778 1028 779
rect 1022 774 1023 778
rect 1027 774 1028 778
rect 1022 773 1028 774
rect 1094 778 1100 779
rect 1094 774 1095 778
rect 1099 774 1100 778
rect 1094 773 1100 774
rect 1166 778 1172 779
rect 1166 774 1167 778
rect 1171 774 1172 778
rect 1166 773 1172 774
rect 1230 778 1236 779
rect 1230 774 1231 778
rect 1235 774 1236 778
rect 1230 773 1236 774
rect 1294 778 1300 779
rect 1294 774 1295 778
rect 1299 774 1300 778
rect 1294 773 1300 774
rect 1358 778 1364 779
rect 1358 774 1359 778
rect 1363 774 1364 778
rect 1358 773 1364 774
rect 1414 778 1420 779
rect 1414 774 1415 778
rect 1419 774 1420 778
rect 1414 773 1420 774
rect 1470 778 1476 779
rect 1470 774 1471 778
rect 1475 774 1476 778
rect 1470 773 1476 774
rect 1526 778 1532 779
rect 1526 774 1527 778
rect 1531 774 1532 778
rect 1526 773 1532 774
rect 1590 778 1596 779
rect 1590 774 1591 778
rect 1595 774 1596 778
rect 1662 776 1663 780
rect 1667 776 1668 780
rect 1662 775 1668 776
rect 1590 773 1596 774
rect 110 763 116 764
rect 110 759 111 763
rect 115 759 116 763
rect 1662 763 1668 764
rect 110 758 116 759
rect 134 761 140 762
rect 134 757 135 761
rect 139 757 140 761
rect 134 756 140 757
rect 174 761 180 762
rect 174 757 175 761
rect 179 757 180 761
rect 174 756 180 757
rect 230 761 236 762
rect 230 757 231 761
rect 235 757 236 761
rect 230 756 236 757
rect 294 761 300 762
rect 294 757 295 761
rect 299 757 300 761
rect 294 756 300 757
rect 366 761 372 762
rect 366 757 367 761
rect 371 757 372 761
rect 366 756 372 757
rect 446 761 452 762
rect 446 757 447 761
rect 451 757 452 761
rect 446 756 452 757
rect 526 761 532 762
rect 526 757 527 761
rect 531 757 532 761
rect 526 756 532 757
rect 614 761 620 762
rect 614 757 615 761
rect 619 757 620 761
rect 614 756 620 757
rect 702 761 708 762
rect 702 757 703 761
rect 707 757 708 761
rect 702 756 708 757
rect 790 761 796 762
rect 790 757 791 761
rect 795 757 796 761
rect 790 756 796 757
rect 870 761 876 762
rect 870 757 871 761
rect 875 757 876 761
rect 870 756 876 757
rect 950 761 956 762
rect 950 757 951 761
rect 955 757 956 761
rect 950 756 956 757
rect 1022 761 1028 762
rect 1022 757 1023 761
rect 1027 757 1028 761
rect 1022 756 1028 757
rect 1094 761 1100 762
rect 1094 757 1095 761
rect 1099 757 1100 761
rect 1094 756 1100 757
rect 1166 761 1172 762
rect 1166 757 1167 761
rect 1171 757 1172 761
rect 1166 756 1172 757
rect 1230 761 1236 762
rect 1230 757 1231 761
rect 1235 757 1236 761
rect 1230 756 1236 757
rect 1294 761 1300 762
rect 1294 757 1295 761
rect 1299 757 1300 761
rect 1294 756 1300 757
rect 1358 761 1364 762
rect 1358 757 1359 761
rect 1363 757 1364 761
rect 1358 756 1364 757
rect 1414 761 1420 762
rect 1414 757 1415 761
rect 1419 757 1420 761
rect 1414 756 1420 757
rect 1470 761 1476 762
rect 1470 757 1471 761
rect 1475 757 1476 761
rect 1470 756 1476 757
rect 1526 761 1532 762
rect 1526 757 1527 761
rect 1531 757 1532 761
rect 1526 756 1532 757
rect 1590 761 1596 762
rect 1590 757 1591 761
rect 1595 757 1596 761
rect 1662 759 1663 763
rect 1667 759 1668 763
rect 1662 758 1668 759
rect 1590 756 1596 757
rect 214 747 220 748
rect 110 745 116 746
rect 110 741 111 745
rect 115 741 116 745
rect 214 743 215 747
rect 219 743 220 747
rect 214 742 220 743
rect 246 747 252 748
rect 246 743 247 747
rect 251 743 252 747
rect 246 742 252 743
rect 278 747 284 748
rect 278 743 279 747
rect 283 743 284 747
rect 278 742 284 743
rect 318 747 324 748
rect 318 743 319 747
rect 323 743 324 747
rect 318 742 324 743
rect 358 747 364 748
rect 358 743 359 747
rect 363 743 364 747
rect 358 742 364 743
rect 398 747 404 748
rect 398 743 399 747
rect 403 743 404 747
rect 398 742 404 743
rect 438 747 444 748
rect 438 743 439 747
rect 443 743 444 747
rect 438 742 444 743
rect 486 747 492 748
rect 486 743 487 747
rect 491 743 492 747
rect 486 742 492 743
rect 542 747 548 748
rect 542 743 543 747
rect 547 743 548 747
rect 542 742 548 743
rect 606 747 612 748
rect 606 743 607 747
rect 611 743 612 747
rect 606 742 612 743
rect 670 747 676 748
rect 670 743 671 747
rect 675 743 676 747
rect 670 742 676 743
rect 734 747 740 748
rect 734 743 735 747
rect 739 743 740 747
rect 734 742 740 743
rect 798 747 804 748
rect 798 743 799 747
rect 803 743 804 747
rect 798 742 804 743
rect 862 747 868 748
rect 862 743 863 747
rect 867 743 868 747
rect 862 742 868 743
rect 926 747 932 748
rect 926 743 927 747
rect 931 743 932 747
rect 926 742 932 743
rect 990 747 996 748
rect 990 743 991 747
rect 995 743 996 747
rect 990 742 996 743
rect 1054 747 1060 748
rect 1054 743 1055 747
rect 1059 743 1060 747
rect 1054 742 1060 743
rect 1118 747 1124 748
rect 1118 743 1119 747
rect 1123 743 1124 747
rect 1118 742 1124 743
rect 1182 747 1188 748
rect 1182 743 1183 747
rect 1187 743 1188 747
rect 1182 742 1188 743
rect 1238 747 1244 748
rect 1238 743 1239 747
rect 1243 743 1244 747
rect 1238 742 1244 743
rect 1294 747 1300 748
rect 1294 743 1295 747
rect 1299 743 1300 747
rect 1294 742 1300 743
rect 1350 747 1356 748
rect 1350 743 1351 747
rect 1355 743 1356 747
rect 1350 742 1356 743
rect 1406 747 1412 748
rect 1406 743 1407 747
rect 1411 743 1412 747
rect 1406 742 1412 743
rect 1462 747 1468 748
rect 1462 743 1463 747
rect 1467 743 1468 747
rect 1462 742 1468 743
rect 1518 747 1524 748
rect 1518 743 1519 747
rect 1523 743 1524 747
rect 1518 742 1524 743
rect 1582 747 1588 748
rect 1582 743 1583 747
rect 1587 743 1588 747
rect 1582 742 1588 743
rect 1622 747 1628 748
rect 1622 743 1623 747
rect 1627 743 1628 747
rect 1622 742 1628 743
rect 1662 745 1668 746
rect 110 740 116 741
rect 1662 741 1663 745
rect 1667 741 1668 745
rect 1662 740 1668 741
rect 214 730 220 731
rect 110 728 116 729
rect 110 724 111 728
rect 115 724 116 728
rect 214 726 215 730
rect 219 726 220 730
rect 214 725 220 726
rect 246 730 252 731
rect 246 726 247 730
rect 251 726 252 730
rect 246 725 252 726
rect 278 730 284 731
rect 278 726 279 730
rect 283 726 284 730
rect 278 725 284 726
rect 318 730 324 731
rect 318 726 319 730
rect 323 726 324 730
rect 318 725 324 726
rect 358 730 364 731
rect 358 726 359 730
rect 363 726 364 730
rect 358 725 364 726
rect 398 730 404 731
rect 398 726 399 730
rect 403 726 404 730
rect 398 725 404 726
rect 438 730 444 731
rect 438 726 439 730
rect 443 726 444 730
rect 438 725 444 726
rect 486 730 492 731
rect 486 726 487 730
rect 491 726 492 730
rect 486 725 492 726
rect 542 730 548 731
rect 542 726 543 730
rect 547 726 548 730
rect 542 725 548 726
rect 606 730 612 731
rect 606 726 607 730
rect 611 726 612 730
rect 606 725 612 726
rect 670 730 676 731
rect 670 726 671 730
rect 675 726 676 730
rect 670 725 676 726
rect 734 730 740 731
rect 734 726 735 730
rect 739 726 740 730
rect 734 725 740 726
rect 798 730 804 731
rect 798 726 799 730
rect 803 726 804 730
rect 798 725 804 726
rect 862 730 868 731
rect 862 726 863 730
rect 867 726 868 730
rect 862 725 868 726
rect 926 730 932 731
rect 926 726 927 730
rect 931 726 932 730
rect 926 725 932 726
rect 990 730 996 731
rect 990 726 991 730
rect 995 726 996 730
rect 990 725 996 726
rect 1054 730 1060 731
rect 1054 726 1055 730
rect 1059 726 1060 730
rect 1054 725 1060 726
rect 1118 730 1124 731
rect 1118 726 1119 730
rect 1123 726 1124 730
rect 1118 725 1124 726
rect 1182 730 1188 731
rect 1182 726 1183 730
rect 1187 726 1188 730
rect 1182 725 1188 726
rect 1238 730 1244 731
rect 1238 726 1239 730
rect 1243 726 1244 730
rect 1238 725 1244 726
rect 1294 730 1300 731
rect 1294 726 1295 730
rect 1299 726 1300 730
rect 1294 725 1300 726
rect 1350 730 1356 731
rect 1350 726 1351 730
rect 1355 726 1356 730
rect 1350 725 1356 726
rect 1406 730 1412 731
rect 1406 726 1407 730
rect 1411 726 1412 730
rect 1406 725 1412 726
rect 1462 730 1468 731
rect 1462 726 1463 730
rect 1467 726 1468 730
rect 1462 725 1468 726
rect 1518 730 1524 731
rect 1518 726 1519 730
rect 1523 726 1524 730
rect 1518 725 1524 726
rect 1582 730 1588 731
rect 1582 726 1583 730
rect 1587 726 1588 730
rect 1582 725 1588 726
rect 1622 730 1628 731
rect 1622 726 1623 730
rect 1627 726 1628 730
rect 1622 725 1628 726
rect 1662 728 1668 729
rect 110 723 116 724
rect 1662 724 1663 728
rect 1667 724 1668 728
rect 1662 723 1668 724
rect 110 696 116 697
rect 110 692 111 696
rect 115 692 116 696
rect 1662 696 1668 697
rect 110 691 116 692
rect 278 694 284 695
rect 278 690 279 694
rect 283 690 284 694
rect 278 689 284 690
rect 310 694 316 695
rect 310 690 311 694
rect 315 690 316 694
rect 310 689 316 690
rect 342 694 348 695
rect 342 690 343 694
rect 347 690 348 694
rect 342 689 348 690
rect 374 694 380 695
rect 374 690 375 694
rect 379 690 380 694
rect 374 689 380 690
rect 406 694 412 695
rect 406 690 407 694
rect 411 690 412 694
rect 406 689 412 690
rect 438 694 444 695
rect 438 690 439 694
rect 443 690 444 694
rect 438 689 444 690
rect 470 694 476 695
rect 470 690 471 694
rect 475 690 476 694
rect 470 689 476 690
rect 502 694 508 695
rect 502 690 503 694
rect 507 690 508 694
rect 502 689 508 690
rect 542 694 548 695
rect 542 690 543 694
rect 547 690 548 694
rect 542 689 548 690
rect 590 694 596 695
rect 590 690 591 694
rect 595 690 596 694
rect 590 689 596 690
rect 646 694 652 695
rect 646 690 647 694
rect 651 690 652 694
rect 646 689 652 690
rect 702 694 708 695
rect 702 690 703 694
rect 707 690 708 694
rect 702 689 708 690
rect 758 694 764 695
rect 758 690 759 694
rect 763 690 764 694
rect 758 689 764 690
rect 822 694 828 695
rect 822 690 823 694
rect 827 690 828 694
rect 822 689 828 690
rect 886 694 892 695
rect 886 690 887 694
rect 891 690 892 694
rect 886 689 892 690
rect 958 694 964 695
rect 958 690 959 694
rect 963 690 964 694
rect 958 689 964 690
rect 1022 694 1028 695
rect 1022 690 1023 694
rect 1027 690 1028 694
rect 1022 689 1028 690
rect 1086 694 1092 695
rect 1086 690 1087 694
rect 1091 690 1092 694
rect 1086 689 1092 690
rect 1158 694 1164 695
rect 1158 690 1159 694
rect 1163 690 1164 694
rect 1158 689 1164 690
rect 1222 694 1228 695
rect 1222 690 1223 694
rect 1227 690 1228 694
rect 1222 689 1228 690
rect 1286 694 1292 695
rect 1286 690 1287 694
rect 1291 690 1292 694
rect 1286 689 1292 690
rect 1350 694 1356 695
rect 1350 690 1351 694
rect 1355 690 1356 694
rect 1350 689 1356 690
rect 1414 694 1420 695
rect 1414 690 1415 694
rect 1419 690 1420 694
rect 1414 689 1420 690
rect 1470 694 1476 695
rect 1470 690 1471 694
rect 1475 690 1476 694
rect 1470 689 1476 690
rect 1526 694 1532 695
rect 1526 690 1527 694
rect 1531 690 1532 694
rect 1526 689 1532 690
rect 1582 694 1588 695
rect 1582 690 1583 694
rect 1587 690 1588 694
rect 1582 689 1588 690
rect 1622 694 1628 695
rect 1622 690 1623 694
rect 1627 690 1628 694
rect 1662 692 1663 696
rect 1667 692 1668 696
rect 1662 691 1668 692
rect 1622 689 1628 690
rect 110 679 116 680
rect 110 675 111 679
rect 115 675 116 679
rect 1662 679 1668 680
rect 110 674 116 675
rect 278 677 284 678
rect 278 673 279 677
rect 283 673 284 677
rect 278 672 284 673
rect 310 677 316 678
rect 310 673 311 677
rect 315 673 316 677
rect 310 672 316 673
rect 342 677 348 678
rect 342 673 343 677
rect 347 673 348 677
rect 342 672 348 673
rect 374 677 380 678
rect 374 673 375 677
rect 379 673 380 677
rect 374 672 380 673
rect 406 677 412 678
rect 406 673 407 677
rect 411 673 412 677
rect 406 672 412 673
rect 438 677 444 678
rect 438 673 439 677
rect 443 673 444 677
rect 438 672 444 673
rect 470 677 476 678
rect 470 673 471 677
rect 475 673 476 677
rect 470 672 476 673
rect 502 677 508 678
rect 502 673 503 677
rect 507 673 508 677
rect 502 672 508 673
rect 542 677 548 678
rect 542 673 543 677
rect 547 673 548 677
rect 542 672 548 673
rect 590 677 596 678
rect 590 673 591 677
rect 595 673 596 677
rect 590 672 596 673
rect 646 677 652 678
rect 646 673 647 677
rect 651 673 652 677
rect 646 672 652 673
rect 702 677 708 678
rect 702 673 703 677
rect 707 673 708 677
rect 702 672 708 673
rect 758 677 764 678
rect 758 673 759 677
rect 763 673 764 677
rect 758 672 764 673
rect 822 677 828 678
rect 822 673 823 677
rect 827 673 828 677
rect 822 672 828 673
rect 886 677 892 678
rect 886 673 887 677
rect 891 673 892 677
rect 886 672 892 673
rect 958 677 964 678
rect 958 673 959 677
rect 963 673 964 677
rect 958 672 964 673
rect 1022 677 1028 678
rect 1022 673 1023 677
rect 1027 673 1028 677
rect 1022 672 1028 673
rect 1086 677 1092 678
rect 1086 673 1087 677
rect 1091 673 1092 677
rect 1086 672 1092 673
rect 1158 677 1164 678
rect 1158 673 1159 677
rect 1163 673 1164 677
rect 1158 672 1164 673
rect 1222 677 1228 678
rect 1222 673 1223 677
rect 1227 673 1228 677
rect 1222 672 1228 673
rect 1286 677 1292 678
rect 1286 673 1287 677
rect 1291 673 1292 677
rect 1286 672 1292 673
rect 1350 677 1356 678
rect 1350 673 1351 677
rect 1355 673 1356 677
rect 1350 672 1356 673
rect 1414 677 1420 678
rect 1414 673 1415 677
rect 1419 673 1420 677
rect 1414 672 1420 673
rect 1470 677 1476 678
rect 1470 673 1471 677
rect 1475 673 1476 677
rect 1470 672 1476 673
rect 1526 677 1532 678
rect 1526 673 1527 677
rect 1531 673 1532 677
rect 1526 672 1532 673
rect 1582 677 1588 678
rect 1582 673 1583 677
rect 1587 673 1588 677
rect 1582 672 1588 673
rect 1622 677 1628 678
rect 1622 673 1623 677
rect 1627 673 1628 677
rect 1662 675 1663 679
rect 1667 675 1668 679
rect 1662 674 1668 675
rect 1622 672 1628 673
rect 294 663 300 664
rect 110 661 116 662
rect 110 657 111 661
rect 115 657 116 661
rect 294 659 295 663
rect 299 659 300 663
rect 294 658 300 659
rect 326 663 332 664
rect 326 659 327 663
rect 331 659 332 663
rect 326 658 332 659
rect 358 663 364 664
rect 358 659 359 663
rect 363 659 364 663
rect 358 658 364 659
rect 390 663 396 664
rect 390 659 391 663
rect 395 659 396 663
rect 390 658 396 659
rect 422 663 428 664
rect 422 659 423 663
rect 427 659 428 663
rect 422 658 428 659
rect 454 663 460 664
rect 454 659 455 663
rect 459 659 460 663
rect 454 658 460 659
rect 486 663 492 664
rect 486 659 487 663
rect 491 659 492 663
rect 486 658 492 659
rect 518 663 524 664
rect 518 659 519 663
rect 523 659 524 663
rect 518 658 524 659
rect 550 663 556 664
rect 550 659 551 663
rect 555 659 556 663
rect 550 658 556 659
rect 590 663 596 664
rect 590 659 591 663
rect 595 659 596 663
rect 590 658 596 659
rect 638 663 644 664
rect 638 659 639 663
rect 643 659 644 663
rect 638 658 644 659
rect 686 663 692 664
rect 686 659 687 663
rect 691 659 692 663
rect 686 658 692 659
rect 734 663 740 664
rect 734 659 735 663
rect 739 659 740 663
rect 734 658 740 659
rect 790 663 796 664
rect 790 659 791 663
rect 795 659 796 663
rect 790 658 796 659
rect 846 663 852 664
rect 846 659 847 663
rect 851 659 852 663
rect 846 658 852 659
rect 910 663 916 664
rect 910 659 911 663
rect 915 659 916 663
rect 910 658 916 659
rect 974 663 980 664
rect 974 659 975 663
rect 979 659 980 663
rect 974 658 980 659
rect 1046 663 1052 664
rect 1046 659 1047 663
rect 1051 659 1052 663
rect 1046 658 1052 659
rect 1126 663 1132 664
rect 1126 659 1127 663
rect 1131 659 1132 663
rect 1126 658 1132 659
rect 1214 663 1220 664
rect 1214 659 1215 663
rect 1219 659 1220 663
rect 1214 658 1220 659
rect 1294 663 1300 664
rect 1294 659 1295 663
rect 1299 659 1300 663
rect 1294 658 1300 659
rect 1382 663 1388 664
rect 1382 659 1383 663
rect 1387 659 1388 663
rect 1382 658 1388 659
rect 1470 663 1476 664
rect 1470 659 1471 663
rect 1475 659 1476 663
rect 1470 658 1476 659
rect 1558 663 1564 664
rect 1558 659 1559 663
rect 1563 659 1564 663
rect 1558 658 1564 659
rect 1622 663 1628 664
rect 1622 659 1623 663
rect 1627 659 1628 663
rect 1622 658 1628 659
rect 1662 661 1668 662
rect 110 656 116 657
rect 1662 657 1663 661
rect 1667 657 1668 661
rect 1662 656 1668 657
rect 294 646 300 647
rect 110 644 116 645
rect 110 640 111 644
rect 115 640 116 644
rect 294 642 295 646
rect 299 642 300 646
rect 294 641 300 642
rect 326 646 332 647
rect 326 642 327 646
rect 331 642 332 646
rect 326 641 332 642
rect 358 646 364 647
rect 358 642 359 646
rect 363 642 364 646
rect 358 641 364 642
rect 390 646 396 647
rect 390 642 391 646
rect 395 642 396 646
rect 390 641 396 642
rect 422 646 428 647
rect 422 642 423 646
rect 427 642 428 646
rect 422 641 428 642
rect 454 646 460 647
rect 454 642 455 646
rect 459 642 460 646
rect 454 641 460 642
rect 486 646 492 647
rect 486 642 487 646
rect 491 642 492 646
rect 486 641 492 642
rect 518 646 524 647
rect 518 642 519 646
rect 523 642 524 646
rect 518 641 524 642
rect 550 646 556 647
rect 550 642 551 646
rect 555 642 556 646
rect 550 641 556 642
rect 590 646 596 647
rect 590 642 591 646
rect 595 642 596 646
rect 590 641 596 642
rect 638 646 644 647
rect 638 642 639 646
rect 643 642 644 646
rect 638 641 644 642
rect 686 646 692 647
rect 686 642 687 646
rect 691 642 692 646
rect 686 641 692 642
rect 734 646 740 647
rect 734 642 735 646
rect 739 642 740 646
rect 734 641 740 642
rect 790 646 796 647
rect 790 642 791 646
rect 795 642 796 646
rect 790 641 796 642
rect 846 646 852 647
rect 846 642 847 646
rect 851 642 852 646
rect 846 641 852 642
rect 910 646 916 647
rect 910 642 911 646
rect 915 642 916 646
rect 910 641 916 642
rect 974 646 980 647
rect 974 642 975 646
rect 979 642 980 646
rect 974 641 980 642
rect 1046 646 1052 647
rect 1046 642 1047 646
rect 1051 642 1052 646
rect 1046 641 1052 642
rect 1126 646 1132 647
rect 1126 642 1127 646
rect 1131 642 1132 646
rect 1126 641 1132 642
rect 1214 646 1220 647
rect 1214 642 1215 646
rect 1219 642 1220 646
rect 1214 641 1220 642
rect 1294 646 1300 647
rect 1294 642 1295 646
rect 1299 642 1300 646
rect 1294 641 1300 642
rect 1382 646 1388 647
rect 1382 642 1383 646
rect 1387 642 1388 646
rect 1382 641 1388 642
rect 1470 646 1476 647
rect 1470 642 1471 646
rect 1475 642 1476 646
rect 1470 641 1476 642
rect 1558 646 1564 647
rect 1558 642 1559 646
rect 1563 642 1564 646
rect 1558 641 1564 642
rect 1622 646 1628 647
rect 1622 642 1623 646
rect 1627 642 1628 646
rect 1622 641 1628 642
rect 1662 644 1668 645
rect 110 639 116 640
rect 1662 640 1663 644
rect 1667 640 1668 644
rect 1662 639 1668 640
rect 110 616 116 617
rect 110 612 111 616
rect 115 612 116 616
rect 1662 616 1668 617
rect 110 611 116 612
rect 246 614 252 615
rect 246 610 247 614
rect 251 610 252 614
rect 246 609 252 610
rect 278 614 284 615
rect 278 610 279 614
rect 283 610 284 614
rect 278 609 284 610
rect 318 614 324 615
rect 318 610 319 614
rect 323 610 324 614
rect 318 609 324 610
rect 366 614 372 615
rect 366 610 367 614
rect 371 610 372 614
rect 366 609 372 610
rect 422 614 428 615
rect 422 610 423 614
rect 427 610 428 614
rect 422 609 428 610
rect 470 614 476 615
rect 470 610 471 614
rect 475 610 476 614
rect 470 609 476 610
rect 518 614 524 615
rect 518 610 519 614
rect 523 610 524 614
rect 518 609 524 610
rect 566 614 572 615
rect 566 610 567 614
rect 571 610 572 614
rect 566 609 572 610
rect 614 614 620 615
rect 614 610 615 614
rect 619 610 620 614
rect 614 609 620 610
rect 662 614 668 615
rect 662 610 663 614
rect 667 610 668 614
rect 662 609 668 610
rect 718 614 724 615
rect 718 610 719 614
rect 723 610 724 614
rect 718 609 724 610
rect 774 614 780 615
rect 774 610 775 614
rect 779 610 780 614
rect 774 609 780 610
rect 830 614 836 615
rect 830 610 831 614
rect 835 610 836 614
rect 830 609 836 610
rect 894 614 900 615
rect 894 610 895 614
rect 899 610 900 614
rect 894 609 900 610
rect 966 614 972 615
rect 966 610 967 614
rect 971 610 972 614
rect 966 609 972 610
rect 1046 614 1052 615
rect 1046 610 1047 614
rect 1051 610 1052 614
rect 1046 609 1052 610
rect 1126 614 1132 615
rect 1126 610 1127 614
rect 1131 610 1132 614
rect 1126 609 1132 610
rect 1206 614 1212 615
rect 1206 610 1207 614
rect 1211 610 1212 614
rect 1206 609 1212 610
rect 1286 614 1292 615
rect 1286 610 1287 614
rect 1291 610 1292 614
rect 1286 609 1292 610
rect 1358 614 1364 615
rect 1358 610 1359 614
rect 1363 610 1364 614
rect 1358 609 1364 610
rect 1430 614 1436 615
rect 1430 610 1431 614
rect 1435 610 1436 614
rect 1430 609 1436 610
rect 1502 614 1508 615
rect 1502 610 1503 614
rect 1507 610 1508 614
rect 1502 609 1508 610
rect 1574 614 1580 615
rect 1574 610 1575 614
rect 1579 610 1580 614
rect 1574 609 1580 610
rect 1622 614 1628 615
rect 1622 610 1623 614
rect 1627 610 1628 614
rect 1662 612 1663 616
rect 1667 612 1668 616
rect 1662 611 1668 612
rect 1622 609 1628 610
rect 110 599 116 600
rect 110 595 111 599
rect 115 595 116 599
rect 1662 599 1668 600
rect 110 594 116 595
rect 246 597 252 598
rect 246 593 247 597
rect 251 593 252 597
rect 246 592 252 593
rect 278 597 284 598
rect 278 593 279 597
rect 283 593 284 597
rect 278 592 284 593
rect 318 597 324 598
rect 318 593 319 597
rect 323 593 324 597
rect 318 592 324 593
rect 366 597 372 598
rect 366 593 367 597
rect 371 593 372 597
rect 366 592 372 593
rect 422 597 428 598
rect 422 593 423 597
rect 427 593 428 597
rect 422 592 428 593
rect 470 597 476 598
rect 470 593 471 597
rect 475 593 476 597
rect 470 592 476 593
rect 518 597 524 598
rect 518 593 519 597
rect 523 593 524 597
rect 518 592 524 593
rect 566 597 572 598
rect 566 593 567 597
rect 571 593 572 597
rect 566 592 572 593
rect 614 597 620 598
rect 614 593 615 597
rect 619 593 620 597
rect 614 592 620 593
rect 662 597 668 598
rect 662 593 663 597
rect 667 593 668 597
rect 662 592 668 593
rect 718 597 724 598
rect 718 593 719 597
rect 723 593 724 597
rect 718 592 724 593
rect 774 597 780 598
rect 774 593 775 597
rect 779 593 780 597
rect 774 592 780 593
rect 830 597 836 598
rect 830 593 831 597
rect 835 593 836 597
rect 830 592 836 593
rect 894 597 900 598
rect 894 593 895 597
rect 899 593 900 597
rect 894 592 900 593
rect 966 597 972 598
rect 966 593 967 597
rect 971 593 972 597
rect 966 592 972 593
rect 1046 597 1052 598
rect 1046 593 1047 597
rect 1051 593 1052 597
rect 1046 592 1052 593
rect 1126 597 1132 598
rect 1126 593 1127 597
rect 1131 593 1132 597
rect 1126 592 1132 593
rect 1206 597 1212 598
rect 1206 593 1207 597
rect 1211 593 1212 597
rect 1206 592 1212 593
rect 1286 597 1292 598
rect 1286 593 1287 597
rect 1291 593 1292 597
rect 1286 592 1292 593
rect 1358 597 1364 598
rect 1358 593 1359 597
rect 1363 593 1364 597
rect 1358 592 1364 593
rect 1430 597 1436 598
rect 1430 593 1431 597
rect 1435 593 1436 597
rect 1430 592 1436 593
rect 1502 597 1508 598
rect 1502 593 1503 597
rect 1507 593 1508 597
rect 1502 592 1508 593
rect 1574 597 1580 598
rect 1574 593 1575 597
rect 1579 593 1580 597
rect 1574 592 1580 593
rect 1622 597 1628 598
rect 1622 593 1623 597
rect 1627 593 1628 597
rect 1662 595 1663 599
rect 1667 595 1668 599
rect 1662 594 1668 595
rect 1622 592 1628 593
rect 166 583 172 584
rect 110 581 116 582
rect 110 577 111 581
rect 115 577 116 581
rect 166 579 167 583
rect 171 579 172 583
rect 166 578 172 579
rect 214 583 220 584
rect 214 579 215 583
rect 219 579 220 583
rect 214 578 220 579
rect 270 583 276 584
rect 270 579 271 583
rect 275 579 276 583
rect 270 578 276 579
rect 334 583 340 584
rect 334 579 335 583
rect 339 579 340 583
rect 334 578 340 579
rect 406 583 412 584
rect 406 579 407 583
rect 411 579 412 583
rect 406 578 412 579
rect 486 583 492 584
rect 486 579 487 583
rect 491 579 492 583
rect 486 578 492 579
rect 558 583 564 584
rect 558 579 559 583
rect 563 579 564 583
rect 558 578 564 579
rect 630 583 636 584
rect 630 579 631 583
rect 635 579 636 583
rect 630 578 636 579
rect 702 583 708 584
rect 702 579 703 583
rect 707 579 708 583
rect 702 578 708 579
rect 766 583 772 584
rect 766 579 767 583
rect 771 579 772 583
rect 766 578 772 579
rect 822 583 828 584
rect 822 579 823 583
rect 827 579 828 583
rect 822 578 828 579
rect 878 583 884 584
rect 878 579 879 583
rect 883 579 884 583
rect 878 578 884 579
rect 934 583 940 584
rect 934 579 935 583
rect 939 579 940 583
rect 934 578 940 579
rect 990 583 996 584
rect 990 579 991 583
rect 995 579 996 583
rect 990 578 996 579
rect 1046 583 1052 584
rect 1046 579 1047 583
rect 1051 579 1052 583
rect 1046 578 1052 579
rect 1102 583 1108 584
rect 1102 579 1103 583
rect 1107 579 1108 583
rect 1102 578 1108 579
rect 1158 583 1164 584
rect 1158 579 1159 583
rect 1163 579 1164 583
rect 1158 578 1164 579
rect 1214 583 1220 584
rect 1214 579 1215 583
rect 1219 579 1220 583
rect 1214 578 1220 579
rect 1270 583 1276 584
rect 1270 579 1271 583
rect 1275 579 1276 583
rect 1270 578 1276 579
rect 1326 583 1332 584
rect 1326 579 1327 583
rect 1331 579 1332 583
rect 1326 578 1332 579
rect 1382 583 1388 584
rect 1382 579 1383 583
rect 1387 579 1388 583
rect 1382 578 1388 579
rect 1446 583 1452 584
rect 1446 579 1447 583
rect 1451 579 1452 583
rect 1446 578 1452 579
rect 1510 583 1516 584
rect 1510 579 1511 583
rect 1515 579 1516 583
rect 1510 578 1516 579
rect 1574 583 1580 584
rect 1574 579 1575 583
rect 1579 579 1580 583
rect 1574 578 1580 579
rect 1622 583 1628 584
rect 1622 579 1623 583
rect 1627 579 1628 583
rect 1622 578 1628 579
rect 1662 581 1668 582
rect 110 576 116 577
rect 1662 577 1663 581
rect 1667 577 1668 581
rect 1662 576 1668 577
rect 166 566 172 567
rect 110 564 116 565
rect 110 560 111 564
rect 115 560 116 564
rect 166 562 167 566
rect 171 562 172 566
rect 166 561 172 562
rect 214 566 220 567
rect 214 562 215 566
rect 219 562 220 566
rect 214 561 220 562
rect 270 566 276 567
rect 270 562 271 566
rect 275 562 276 566
rect 270 561 276 562
rect 334 566 340 567
rect 334 562 335 566
rect 339 562 340 566
rect 334 561 340 562
rect 406 566 412 567
rect 406 562 407 566
rect 411 562 412 566
rect 406 561 412 562
rect 486 566 492 567
rect 486 562 487 566
rect 491 562 492 566
rect 486 561 492 562
rect 558 566 564 567
rect 558 562 559 566
rect 563 562 564 566
rect 558 561 564 562
rect 630 566 636 567
rect 630 562 631 566
rect 635 562 636 566
rect 630 561 636 562
rect 702 566 708 567
rect 702 562 703 566
rect 707 562 708 566
rect 702 561 708 562
rect 766 566 772 567
rect 766 562 767 566
rect 771 562 772 566
rect 766 561 772 562
rect 822 566 828 567
rect 822 562 823 566
rect 827 562 828 566
rect 822 561 828 562
rect 878 566 884 567
rect 878 562 879 566
rect 883 562 884 566
rect 878 561 884 562
rect 934 566 940 567
rect 934 562 935 566
rect 939 562 940 566
rect 934 561 940 562
rect 990 566 996 567
rect 990 562 991 566
rect 995 562 996 566
rect 990 561 996 562
rect 1046 566 1052 567
rect 1046 562 1047 566
rect 1051 562 1052 566
rect 1046 561 1052 562
rect 1102 566 1108 567
rect 1102 562 1103 566
rect 1107 562 1108 566
rect 1102 561 1108 562
rect 1158 566 1164 567
rect 1158 562 1159 566
rect 1163 562 1164 566
rect 1158 561 1164 562
rect 1214 566 1220 567
rect 1214 562 1215 566
rect 1219 562 1220 566
rect 1214 561 1220 562
rect 1270 566 1276 567
rect 1270 562 1271 566
rect 1275 562 1276 566
rect 1270 561 1276 562
rect 1326 566 1332 567
rect 1326 562 1327 566
rect 1331 562 1332 566
rect 1326 561 1332 562
rect 1382 566 1388 567
rect 1382 562 1383 566
rect 1387 562 1388 566
rect 1382 561 1388 562
rect 1446 566 1452 567
rect 1446 562 1447 566
rect 1451 562 1452 566
rect 1446 561 1452 562
rect 1510 566 1516 567
rect 1510 562 1511 566
rect 1515 562 1516 566
rect 1510 561 1516 562
rect 1574 566 1580 567
rect 1574 562 1575 566
rect 1579 562 1580 566
rect 1574 561 1580 562
rect 1622 566 1628 567
rect 1622 562 1623 566
rect 1627 562 1628 566
rect 1622 561 1628 562
rect 1662 564 1668 565
rect 110 559 116 560
rect 1662 560 1663 564
rect 1667 560 1668 564
rect 1662 559 1668 560
rect 110 532 116 533
rect 110 528 111 532
rect 115 528 116 532
rect 1662 532 1668 533
rect 110 527 116 528
rect 134 530 140 531
rect 134 526 135 530
rect 139 526 140 530
rect 134 525 140 526
rect 166 530 172 531
rect 166 526 167 530
rect 171 526 172 530
rect 166 525 172 526
rect 198 530 204 531
rect 198 526 199 530
rect 203 526 204 530
rect 198 525 204 526
rect 230 530 236 531
rect 230 526 231 530
rect 235 526 236 530
rect 230 525 236 526
rect 278 530 284 531
rect 278 526 279 530
rect 283 526 284 530
rect 278 525 284 526
rect 326 530 332 531
rect 326 526 327 530
rect 331 526 332 530
rect 326 525 332 526
rect 374 530 380 531
rect 374 526 375 530
rect 379 526 380 530
rect 374 525 380 526
rect 430 530 436 531
rect 430 526 431 530
rect 435 526 436 530
rect 430 525 436 526
rect 494 530 500 531
rect 494 526 495 530
rect 499 526 500 530
rect 494 525 500 526
rect 558 530 564 531
rect 558 526 559 530
rect 563 526 564 530
rect 558 525 564 526
rect 622 530 628 531
rect 622 526 623 530
rect 627 526 628 530
rect 622 525 628 526
rect 686 530 692 531
rect 686 526 687 530
rect 691 526 692 530
rect 686 525 692 526
rect 750 530 756 531
rect 750 526 751 530
rect 755 526 756 530
rect 750 525 756 526
rect 814 530 820 531
rect 814 526 815 530
rect 819 526 820 530
rect 814 525 820 526
rect 878 530 884 531
rect 878 526 879 530
rect 883 526 884 530
rect 878 525 884 526
rect 942 530 948 531
rect 942 526 943 530
rect 947 526 948 530
rect 942 525 948 526
rect 1006 530 1012 531
rect 1006 526 1007 530
rect 1011 526 1012 530
rect 1006 525 1012 526
rect 1070 530 1076 531
rect 1070 526 1071 530
rect 1075 526 1076 530
rect 1070 525 1076 526
rect 1126 530 1132 531
rect 1126 526 1127 530
rect 1131 526 1132 530
rect 1126 525 1132 526
rect 1182 530 1188 531
rect 1182 526 1183 530
rect 1187 526 1188 530
rect 1182 525 1188 526
rect 1230 530 1236 531
rect 1230 526 1231 530
rect 1235 526 1236 530
rect 1230 525 1236 526
rect 1278 530 1284 531
rect 1278 526 1279 530
rect 1283 526 1284 530
rect 1278 525 1284 526
rect 1334 530 1340 531
rect 1334 526 1335 530
rect 1339 526 1340 530
rect 1334 525 1340 526
rect 1390 530 1396 531
rect 1390 526 1391 530
rect 1395 526 1396 530
rect 1390 525 1396 526
rect 1446 530 1452 531
rect 1446 526 1447 530
rect 1451 526 1452 530
rect 1446 525 1452 526
rect 1510 530 1516 531
rect 1510 526 1511 530
rect 1515 526 1516 530
rect 1510 525 1516 526
rect 1574 530 1580 531
rect 1574 526 1575 530
rect 1579 526 1580 530
rect 1574 525 1580 526
rect 1622 530 1628 531
rect 1622 526 1623 530
rect 1627 526 1628 530
rect 1662 528 1663 532
rect 1667 528 1668 532
rect 1662 527 1668 528
rect 1622 525 1628 526
rect 110 515 116 516
rect 110 511 111 515
rect 115 511 116 515
rect 1662 515 1668 516
rect 110 510 116 511
rect 134 513 140 514
rect 134 509 135 513
rect 139 509 140 513
rect 134 508 140 509
rect 166 513 172 514
rect 166 509 167 513
rect 171 509 172 513
rect 166 508 172 509
rect 198 513 204 514
rect 198 509 199 513
rect 203 509 204 513
rect 198 508 204 509
rect 230 513 236 514
rect 230 509 231 513
rect 235 509 236 513
rect 230 508 236 509
rect 278 513 284 514
rect 278 509 279 513
rect 283 509 284 513
rect 278 508 284 509
rect 326 513 332 514
rect 326 509 327 513
rect 331 509 332 513
rect 326 508 332 509
rect 374 513 380 514
rect 374 509 375 513
rect 379 509 380 513
rect 374 508 380 509
rect 430 513 436 514
rect 430 509 431 513
rect 435 509 436 513
rect 430 508 436 509
rect 494 513 500 514
rect 494 509 495 513
rect 499 509 500 513
rect 494 508 500 509
rect 558 513 564 514
rect 558 509 559 513
rect 563 509 564 513
rect 558 508 564 509
rect 622 513 628 514
rect 622 509 623 513
rect 627 509 628 513
rect 622 508 628 509
rect 686 513 692 514
rect 686 509 687 513
rect 691 509 692 513
rect 686 508 692 509
rect 750 513 756 514
rect 750 509 751 513
rect 755 509 756 513
rect 750 508 756 509
rect 814 513 820 514
rect 814 509 815 513
rect 819 509 820 513
rect 814 508 820 509
rect 878 513 884 514
rect 878 509 879 513
rect 883 509 884 513
rect 878 508 884 509
rect 942 513 948 514
rect 942 509 943 513
rect 947 509 948 513
rect 942 508 948 509
rect 1006 513 1012 514
rect 1006 509 1007 513
rect 1011 509 1012 513
rect 1006 508 1012 509
rect 1070 513 1076 514
rect 1070 509 1071 513
rect 1075 509 1076 513
rect 1070 508 1076 509
rect 1126 513 1132 514
rect 1126 509 1127 513
rect 1131 509 1132 513
rect 1126 508 1132 509
rect 1182 513 1188 514
rect 1182 509 1183 513
rect 1187 509 1188 513
rect 1182 508 1188 509
rect 1230 513 1236 514
rect 1230 509 1231 513
rect 1235 509 1236 513
rect 1230 508 1236 509
rect 1278 513 1284 514
rect 1278 509 1279 513
rect 1283 509 1284 513
rect 1278 508 1284 509
rect 1334 513 1340 514
rect 1334 509 1335 513
rect 1339 509 1340 513
rect 1334 508 1340 509
rect 1390 513 1396 514
rect 1390 509 1391 513
rect 1395 509 1396 513
rect 1390 508 1396 509
rect 1446 513 1452 514
rect 1446 509 1447 513
rect 1451 509 1452 513
rect 1446 508 1452 509
rect 1510 513 1516 514
rect 1510 509 1511 513
rect 1515 509 1516 513
rect 1510 508 1516 509
rect 1574 513 1580 514
rect 1574 509 1575 513
rect 1579 509 1580 513
rect 1574 508 1580 509
rect 1622 513 1628 514
rect 1622 509 1623 513
rect 1627 509 1628 513
rect 1662 511 1663 515
rect 1667 511 1668 515
rect 1662 510 1668 511
rect 1622 508 1628 509
rect 134 499 140 500
rect 110 497 116 498
rect 110 493 111 497
rect 115 493 116 497
rect 134 495 135 499
rect 139 495 140 499
rect 134 494 140 495
rect 166 499 172 500
rect 166 495 167 499
rect 171 495 172 499
rect 166 494 172 495
rect 198 499 204 500
rect 198 495 199 499
rect 203 495 204 499
rect 198 494 204 495
rect 238 499 244 500
rect 238 495 239 499
rect 243 495 244 499
rect 238 494 244 495
rect 286 499 292 500
rect 286 495 287 499
rect 291 495 292 499
rect 286 494 292 495
rect 326 499 332 500
rect 326 495 327 499
rect 331 495 332 499
rect 326 494 332 495
rect 374 499 380 500
rect 374 495 375 499
rect 379 495 380 499
rect 374 494 380 495
rect 422 499 428 500
rect 422 495 423 499
rect 427 495 428 499
rect 422 494 428 495
rect 478 499 484 500
rect 478 495 479 499
rect 483 495 484 499
rect 478 494 484 495
rect 542 499 548 500
rect 542 495 543 499
rect 547 495 548 499
rect 542 494 548 495
rect 614 499 620 500
rect 614 495 615 499
rect 619 495 620 499
rect 614 494 620 495
rect 694 499 700 500
rect 694 495 695 499
rect 699 495 700 499
rect 694 494 700 495
rect 774 499 780 500
rect 774 495 775 499
rect 779 495 780 499
rect 774 494 780 495
rect 846 499 852 500
rect 846 495 847 499
rect 851 495 852 499
rect 846 494 852 495
rect 918 499 924 500
rect 918 495 919 499
rect 923 495 924 499
rect 918 494 924 495
rect 982 499 988 500
rect 982 495 983 499
rect 987 495 988 499
rect 982 494 988 495
rect 1038 499 1044 500
rect 1038 495 1039 499
rect 1043 495 1044 499
rect 1038 494 1044 495
rect 1094 499 1100 500
rect 1094 495 1095 499
rect 1099 495 1100 499
rect 1094 494 1100 495
rect 1142 499 1148 500
rect 1142 495 1143 499
rect 1147 495 1148 499
rect 1142 494 1148 495
rect 1190 499 1196 500
rect 1190 495 1191 499
rect 1195 495 1196 499
rect 1190 494 1196 495
rect 1238 499 1244 500
rect 1238 495 1239 499
rect 1243 495 1244 499
rect 1238 494 1244 495
rect 1286 499 1292 500
rect 1286 495 1287 499
rect 1291 495 1292 499
rect 1286 494 1292 495
rect 1334 499 1340 500
rect 1334 495 1335 499
rect 1339 495 1340 499
rect 1334 494 1340 495
rect 1382 499 1388 500
rect 1382 495 1383 499
rect 1387 495 1388 499
rect 1382 494 1388 495
rect 1430 499 1436 500
rect 1430 495 1431 499
rect 1435 495 1436 499
rect 1430 494 1436 495
rect 1478 499 1484 500
rect 1478 495 1479 499
rect 1483 495 1484 499
rect 1478 494 1484 495
rect 1534 499 1540 500
rect 1534 495 1535 499
rect 1539 495 1540 499
rect 1534 494 1540 495
rect 1590 499 1596 500
rect 1590 495 1591 499
rect 1595 495 1596 499
rect 1590 494 1596 495
rect 1622 499 1628 500
rect 1622 495 1623 499
rect 1627 495 1628 499
rect 1622 494 1628 495
rect 1662 497 1668 498
rect 110 492 116 493
rect 1662 493 1663 497
rect 1667 493 1668 497
rect 1662 492 1668 493
rect 134 482 140 483
rect 110 480 116 481
rect 110 476 111 480
rect 115 476 116 480
rect 134 478 135 482
rect 139 478 140 482
rect 134 477 140 478
rect 166 482 172 483
rect 166 478 167 482
rect 171 478 172 482
rect 166 477 172 478
rect 198 482 204 483
rect 198 478 199 482
rect 203 478 204 482
rect 198 477 204 478
rect 238 482 244 483
rect 238 478 239 482
rect 243 478 244 482
rect 238 477 244 478
rect 286 482 292 483
rect 286 478 287 482
rect 291 478 292 482
rect 286 477 292 478
rect 326 482 332 483
rect 326 478 327 482
rect 331 478 332 482
rect 326 477 332 478
rect 374 482 380 483
rect 374 478 375 482
rect 379 478 380 482
rect 374 477 380 478
rect 422 482 428 483
rect 422 478 423 482
rect 427 478 428 482
rect 422 477 428 478
rect 478 482 484 483
rect 478 478 479 482
rect 483 478 484 482
rect 478 477 484 478
rect 542 482 548 483
rect 542 478 543 482
rect 547 478 548 482
rect 542 477 548 478
rect 614 482 620 483
rect 614 478 615 482
rect 619 478 620 482
rect 614 477 620 478
rect 694 482 700 483
rect 694 478 695 482
rect 699 478 700 482
rect 694 477 700 478
rect 774 482 780 483
rect 774 478 775 482
rect 779 478 780 482
rect 774 477 780 478
rect 846 482 852 483
rect 846 478 847 482
rect 851 478 852 482
rect 846 477 852 478
rect 918 482 924 483
rect 918 478 919 482
rect 923 478 924 482
rect 918 477 924 478
rect 982 482 988 483
rect 982 478 983 482
rect 987 478 988 482
rect 982 477 988 478
rect 1038 482 1044 483
rect 1038 478 1039 482
rect 1043 478 1044 482
rect 1038 477 1044 478
rect 1094 482 1100 483
rect 1094 478 1095 482
rect 1099 478 1100 482
rect 1094 477 1100 478
rect 1142 482 1148 483
rect 1142 478 1143 482
rect 1147 478 1148 482
rect 1142 477 1148 478
rect 1190 482 1196 483
rect 1190 478 1191 482
rect 1195 478 1196 482
rect 1190 477 1196 478
rect 1238 482 1244 483
rect 1238 478 1239 482
rect 1243 478 1244 482
rect 1238 477 1244 478
rect 1286 482 1292 483
rect 1286 478 1287 482
rect 1291 478 1292 482
rect 1286 477 1292 478
rect 1334 482 1340 483
rect 1334 478 1335 482
rect 1339 478 1340 482
rect 1334 477 1340 478
rect 1382 482 1388 483
rect 1382 478 1383 482
rect 1387 478 1388 482
rect 1382 477 1388 478
rect 1430 482 1436 483
rect 1430 478 1431 482
rect 1435 478 1436 482
rect 1430 477 1436 478
rect 1478 482 1484 483
rect 1478 478 1479 482
rect 1483 478 1484 482
rect 1478 477 1484 478
rect 1534 482 1540 483
rect 1534 478 1535 482
rect 1539 478 1540 482
rect 1534 477 1540 478
rect 1590 482 1596 483
rect 1590 478 1591 482
rect 1595 478 1596 482
rect 1590 477 1596 478
rect 1622 482 1628 483
rect 1622 478 1623 482
rect 1627 478 1628 482
rect 1622 477 1628 478
rect 1662 480 1668 481
rect 110 475 116 476
rect 1662 476 1663 480
rect 1667 476 1668 480
rect 1662 475 1668 476
rect 110 452 116 453
rect 110 448 111 452
rect 115 448 116 452
rect 1662 452 1668 453
rect 110 447 116 448
rect 150 450 156 451
rect 150 446 151 450
rect 155 446 156 450
rect 150 445 156 446
rect 206 450 212 451
rect 206 446 207 450
rect 211 446 212 450
rect 206 445 212 446
rect 254 450 260 451
rect 254 446 255 450
rect 259 446 260 450
rect 254 445 260 446
rect 310 450 316 451
rect 310 446 311 450
rect 315 446 316 450
rect 310 445 316 446
rect 366 450 372 451
rect 366 446 367 450
rect 371 446 372 450
rect 366 445 372 446
rect 438 450 444 451
rect 438 446 439 450
rect 443 446 444 450
rect 438 445 444 446
rect 518 450 524 451
rect 518 446 519 450
rect 523 446 524 450
rect 518 445 524 446
rect 598 450 604 451
rect 598 446 599 450
rect 603 446 604 450
rect 598 445 604 446
rect 678 450 684 451
rect 678 446 679 450
rect 683 446 684 450
rect 678 445 684 446
rect 758 450 764 451
rect 758 446 759 450
rect 763 446 764 450
rect 758 445 764 446
rect 838 450 844 451
rect 838 446 839 450
rect 843 446 844 450
rect 838 445 844 446
rect 910 450 916 451
rect 910 446 911 450
rect 915 446 916 450
rect 910 445 916 446
rect 982 450 988 451
rect 982 446 983 450
rect 987 446 988 450
rect 982 445 988 446
rect 1054 450 1060 451
rect 1054 446 1055 450
rect 1059 446 1060 450
rect 1054 445 1060 446
rect 1126 450 1132 451
rect 1126 446 1127 450
rect 1131 446 1132 450
rect 1126 445 1132 446
rect 1198 450 1204 451
rect 1198 446 1199 450
rect 1203 446 1204 450
rect 1198 445 1204 446
rect 1262 450 1268 451
rect 1262 446 1263 450
rect 1267 446 1268 450
rect 1262 445 1268 446
rect 1318 450 1324 451
rect 1318 446 1319 450
rect 1323 446 1324 450
rect 1318 445 1324 446
rect 1374 450 1380 451
rect 1374 446 1375 450
rect 1379 446 1380 450
rect 1374 445 1380 446
rect 1430 450 1436 451
rect 1430 446 1431 450
rect 1435 446 1436 450
rect 1430 445 1436 446
rect 1494 450 1500 451
rect 1494 446 1495 450
rect 1499 446 1500 450
rect 1662 448 1663 452
rect 1667 448 1668 452
rect 1662 447 1668 448
rect 1494 445 1500 446
rect 110 435 116 436
rect 110 431 111 435
rect 115 431 116 435
rect 1662 435 1668 436
rect 110 430 116 431
rect 150 433 156 434
rect 150 429 151 433
rect 155 429 156 433
rect 150 428 156 429
rect 206 433 212 434
rect 206 429 207 433
rect 211 429 212 433
rect 206 428 212 429
rect 254 433 260 434
rect 254 429 255 433
rect 259 429 260 433
rect 254 428 260 429
rect 310 433 316 434
rect 310 429 311 433
rect 315 429 316 433
rect 310 428 316 429
rect 366 433 372 434
rect 366 429 367 433
rect 371 429 372 433
rect 366 428 372 429
rect 438 433 444 434
rect 438 429 439 433
rect 443 429 444 433
rect 438 428 444 429
rect 518 433 524 434
rect 518 429 519 433
rect 523 429 524 433
rect 518 428 524 429
rect 598 433 604 434
rect 598 429 599 433
rect 603 429 604 433
rect 598 428 604 429
rect 678 433 684 434
rect 678 429 679 433
rect 683 429 684 433
rect 678 428 684 429
rect 758 433 764 434
rect 758 429 759 433
rect 763 429 764 433
rect 758 428 764 429
rect 838 433 844 434
rect 838 429 839 433
rect 843 429 844 433
rect 838 428 844 429
rect 910 433 916 434
rect 910 429 911 433
rect 915 429 916 433
rect 910 428 916 429
rect 982 433 988 434
rect 982 429 983 433
rect 987 429 988 433
rect 982 428 988 429
rect 1054 433 1060 434
rect 1054 429 1055 433
rect 1059 429 1060 433
rect 1054 428 1060 429
rect 1126 433 1132 434
rect 1126 429 1127 433
rect 1131 429 1132 433
rect 1126 428 1132 429
rect 1198 433 1204 434
rect 1198 429 1199 433
rect 1203 429 1204 433
rect 1198 428 1204 429
rect 1262 433 1268 434
rect 1262 429 1263 433
rect 1267 429 1268 433
rect 1262 428 1268 429
rect 1318 433 1324 434
rect 1318 429 1319 433
rect 1323 429 1324 433
rect 1318 428 1324 429
rect 1374 433 1380 434
rect 1374 429 1375 433
rect 1379 429 1380 433
rect 1374 428 1380 429
rect 1430 433 1436 434
rect 1430 429 1431 433
rect 1435 429 1436 433
rect 1430 428 1436 429
rect 1494 433 1500 434
rect 1494 429 1495 433
rect 1499 429 1500 433
rect 1662 431 1663 435
rect 1667 431 1668 435
rect 1662 430 1668 431
rect 1494 428 1500 429
rect 174 419 180 420
rect 110 417 116 418
rect 110 413 111 417
rect 115 413 116 417
rect 174 415 175 419
rect 179 415 180 419
rect 174 414 180 415
rect 222 419 228 420
rect 222 415 223 419
rect 227 415 228 419
rect 222 414 228 415
rect 270 419 276 420
rect 270 415 271 419
rect 275 415 276 419
rect 270 414 276 415
rect 318 419 324 420
rect 318 415 319 419
rect 323 415 324 419
rect 318 414 324 415
rect 366 419 372 420
rect 366 415 367 419
rect 371 415 372 419
rect 366 414 372 415
rect 414 419 420 420
rect 414 415 415 419
rect 419 415 420 419
rect 414 414 420 415
rect 470 419 476 420
rect 470 415 471 419
rect 475 415 476 419
rect 470 414 476 415
rect 526 419 532 420
rect 526 415 527 419
rect 531 415 532 419
rect 526 414 532 415
rect 590 419 596 420
rect 590 415 591 419
rect 595 415 596 419
rect 590 414 596 415
rect 662 419 668 420
rect 662 415 663 419
rect 667 415 668 419
rect 662 414 668 415
rect 734 419 740 420
rect 734 415 735 419
rect 739 415 740 419
rect 734 414 740 415
rect 806 419 812 420
rect 806 415 807 419
rect 811 415 812 419
rect 806 414 812 415
rect 870 419 876 420
rect 870 415 871 419
rect 875 415 876 419
rect 870 414 876 415
rect 934 419 940 420
rect 934 415 935 419
rect 939 415 940 419
rect 934 414 940 415
rect 990 419 996 420
rect 990 415 991 419
rect 995 415 996 419
rect 990 414 996 415
rect 1038 419 1044 420
rect 1038 415 1039 419
rect 1043 415 1044 419
rect 1038 414 1044 415
rect 1086 419 1092 420
rect 1086 415 1087 419
rect 1091 415 1092 419
rect 1086 414 1092 415
rect 1126 419 1132 420
rect 1126 415 1127 419
rect 1131 415 1132 419
rect 1126 414 1132 415
rect 1166 419 1172 420
rect 1166 415 1167 419
rect 1171 415 1172 419
rect 1166 414 1172 415
rect 1206 419 1212 420
rect 1206 415 1207 419
rect 1211 415 1212 419
rect 1206 414 1212 415
rect 1246 419 1252 420
rect 1246 415 1247 419
rect 1251 415 1252 419
rect 1246 414 1252 415
rect 1286 419 1292 420
rect 1286 415 1287 419
rect 1291 415 1292 419
rect 1286 414 1292 415
rect 1334 419 1340 420
rect 1334 415 1335 419
rect 1339 415 1340 419
rect 1334 414 1340 415
rect 1382 419 1388 420
rect 1382 415 1383 419
rect 1387 415 1388 419
rect 1382 414 1388 415
rect 1662 417 1668 418
rect 110 412 116 413
rect 1662 413 1663 417
rect 1667 413 1668 417
rect 1662 412 1668 413
rect 174 402 180 403
rect 110 400 116 401
rect 110 396 111 400
rect 115 396 116 400
rect 174 398 175 402
rect 179 398 180 402
rect 174 397 180 398
rect 222 402 228 403
rect 222 398 223 402
rect 227 398 228 402
rect 222 397 228 398
rect 270 402 276 403
rect 270 398 271 402
rect 275 398 276 402
rect 270 397 276 398
rect 318 402 324 403
rect 318 398 319 402
rect 323 398 324 402
rect 318 397 324 398
rect 366 402 372 403
rect 366 398 367 402
rect 371 398 372 402
rect 366 397 372 398
rect 414 402 420 403
rect 414 398 415 402
rect 419 398 420 402
rect 414 397 420 398
rect 470 402 476 403
rect 470 398 471 402
rect 475 398 476 402
rect 470 397 476 398
rect 526 402 532 403
rect 526 398 527 402
rect 531 398 532 402
rect 526 397 532 398
rect 590 402 596 403
rect 590 398 591 402
rect 595 398 596 402
rect 590 397 596 398
rect 662 402 668 403
rect 662 398 663 402
rect 667 398 668 402
rect 662 397 668 398
rect 734 402 740 403
rect 734 398 735 402
rect 739 398 740 402
rect 734 397 740 398
rect 806 402 812 403
rect 806 398 807 402
rect 811 398 812 402
rect 806 397 812 398
rect 870 402 876 403
rect 870 398 871 402
rect 875 398 876 402
rect 870 397 876 398
rect 934 402 940 403
rect 934 398 935 402
rect 939 398 940 402
rect 934 397 940 398
rect 990 402 996 403
rect 990 398 991 402
rect 995 398 996 402
rect 990 397 996 398
rect 1038 402 1044 403
rect 1038 398 1039 402
rect 1043 398 1044 402
rect 1038 397 1044 398
rect 1086 402 1092 403
rect 1086 398 1087 402
rect 1091 398 1092 402
rect 1086 397 1092 398
rect 1126 402 1132 403
rect 1126 398 1127 402
rect 1131 398 1132 402
rect 1126 397 1132 398
rect 1166 402 1172 403
rect 1166 398 1167 402
rect 1171 398 1172 402
rect 1166 397 1172 398
rect 1206 402 1212 403
rect 1206 398 1207 402
rect 1211 398 1212 402
rect 1206 397 1212 398
rect 1246 402 1252 403
rect 1246 398 1247 402
rect 1251 398 1252 402
rect 1246 397 1252 398
rect 1286 402 1292 403
rect 1286 398 1287 402
rect 1291 398 1292 402
rect 1286 397 1292 398
rect 1334 402 1340 403
rect 1334 398 1335 402
rect 1339 398 1340 402
rect 1334 397 1340 398
rect 1382 402 1388 403
rect 1382 398 1383 402
rect 1387 398 1388 402
rect 1382 397 1388 398
rect 1662 400 1668 401
rect 110 395 116 396
rect 1662 396 1663 400
rect 1667 396 1668 400
rect 1662 395 1668 396
rect 110 368 116 369
rect 110 364 111 368
rect 115 364 116 368
rect 1662 368 1668 369
rect 110 363 116 364
rect 134 366 140 367
rect 134 362 135 366
rect 139 362 140 366
rect 134 361 140 362
rect 166 366 172 367
rect 166 362 167 366
rect 171 362 172 366
rect 166 361 172 362
rect 198 366 204 367
rect 198 362 199 366
rect 203 362 204 366
rect 198 361 204 362
rect 238 366 244 367
rect 238 362 239 366
rect 243 362 244 366
rect 238 361 244 362
rect 294 366 300 367
rect 294 362 295 366
rect 299 362 300 366
rect 294 361 300 362
rect 350 366 356 367
rect 350 362 351 366
rect 355 362 356 366
rect 350 361 356 362
rect 406 366 412 367
rect 406 362 407 366
rect 411 362 412 366
rect 406 361 412 362
rect 462 366 468 367
rect 462 362 463 366
rect 467 362 468 366
rect 462 361 468 362
rect 518 366 524 367
rect 518 362 519 366
rect 523 362 524 366
rect 518 361 524 362
rect 574 366 580 367
rect 574 362 575 366
rect 579 362 580 366
rect 574 361 580 362
rect 630 366 636 367
rect 630 362 631 366
rect 635 362 636 366
rect 630 361 636 362
rect 686 366 692 367
rect 686 362 687 366
rect 691 362 692 366
rect 686 361 692 362
rect 742 366 748 367
rect 742 362 743 366
rect 747 362 748 366
rect 742 361 748 362
rect 798 366 804 367
rect 798 362 799 366
rect 803 362 804 366
rect 798 361 804 362
rect 854 366 860 367
rect 854 362 855 366
rect 859 362 860 366
rect 854 361 860 362
rect 918 366 924 367
rect 918 362 919 366
rect 923 362 924 366
rect 918 361 924 362
rect 982 366 988 367
rect 982 362 983 366
rect 987 362 988 366
rect 982 361 988 362
rect 1038 366 1044 367
rect 1038 362 1039 366
rect 1043 362 1044 366
rect 1038 361 1044 362
rect 1094 366 1100 367
rect 1094 362 1095 366
rect 1099 362 1100 366
rect 1094 361 1100 362
rect 1150 366 1156 367
rect 1150 362 1151 366
rect 1155 362 1156 366
rect 1150 361 1156 362
rect 1206 366 1212 367
rect 1206 362 1207 366
rect 1211 362 1212 366
rect 1206 361 1212 362
rect 1254 366 1260 367
rect 1254 362 1255 366
rect 1259 362 1260 366
rect 1254 361 1260 362
rect 1302 366 1308 367
rect 1302 362 1303 366
rect 1307 362 1308 366
rect 1302 361 1308 362
rect 1350 366 1356 367
rect 1350 362 1351 366
rect 1355 362 1356 366
rect 1350 361 1356 362
rect 1398 366 1404 367
rect 1398 362 1399 366
rect 1403 362 1404 366
rect 1398 361 1404 362
rect 1446 366 1452 367
rect 1446 362 1447 366
rect 1451 362 1452 366
rect 1446 361 1452 362
rect 1494 366 1500 367
rect 1494 362 1495 366
rect 1499 362 1500 366
rect 1494 361 1500 362
rect 1542 366 1548 367
rect 1542 362 1543 366
rect 1547 362 1548 366
rect 1542 361 1548 362
rect 1590 366 1596 367
rect 1590 362 1591 366
rect 1595 362 1596 366
rect 1590 361 1596 362
rect 1622 366 1628 367
rect 1622 362 1623 366
rect 1627 362 1628 366
rect 1662 364 1663 368
rect 1667 364 1668 368
rect 1662 363 1668 364
rect 1622 361 1628 362
rect 110 351 116 352
rect 110 347 111 351
rect 115 347 116 351
rect 1662 351 1668 352
rect 110 346 116 347
rect 134 349 140 350
rect 134 345 135 349
rect 139 345 140 349
rect 134 344 140 345
rect 166 349 172 350
rect 166 345 167 349
rect 171 345 172 349
rect 166 344 172 345
rect 198 349 204 350
rect 198 345 199 349
rect 203 345 204 349
rect 198 344 204 345
rect 238 349 244 350
rect 238 345 239 349
rect 243 345 244 349
rect 238 344 244 345
rect 294 349 300 350
rect 294 345 295 349
rect 299 345 300 349
rect 294 344 300 345
rect 350 349 356 350
rect 350 345 351 349
rect 355 345 356 349
rect 350 344 356 345
rect 406 349 412 350
rect 406 345 407 349
rect 411 345 412 349
rect 406 344 412 345
rect 462 349 468 350
rect 462 345 463 349
rect 467 345 468 349
rect 462 344 468 345
rect 518 349 524 350
rect 518 345 519 349
rect 523 345 524 349
rect 518 344 524 345
rect 574 349 580 350
rect 574 345 575 349
rect 579 345 580 349
rect 574 344 580 345
rect 630 349 636 350
rect 630 345 631 349
rect 635 345 636 349
rect 630 344 636 345
rect 686 349 692 350
rect 686 345 687 349
rect 691 345 692 349
rect 686 344 692 345
rect 742 349 748 350
rect 742 345 743 349
rect 747 345 748 349
rect 742 344 748 345
rect 798 349 804 350
rect 798 345 799 349
rect 803 345 804 349
rect 798 344 804 345
rect 854 349 860 350
rect 854 345 855 349
rect 859 345 860 349
rect 854 344 860 345
rect 918 349 924 350
rect 918 345 919 349
rect 923 345 924 349
rect 918 344 924 345
rect 982 349 988 350
rect 982 345 983 349
rect 987 345 988 349
rect 982 344 988 345
rect 1038 349 1044 350
rect 1038 345 1039 349
rect 1043 345 1044 349
rect 1038 344 1044 345
rect 1094 349 1100 350
rect 1094 345 1095 349
rect 1099 345 1100 349
rect 1094 344 1100 345
rect 1150 349 1156 350
rect 1150 345 1151 349
rect 1155 345 1156 349
rect 1150 344 1156 345
rect 1206 349 1212 350
rect 1206 345 1207 349
rect 1211 345 1212 349
rect 1206 344 1212 345
rect 1254 349 1260 350
rect 1254 345 1255 349
rect 1259 345 1260 349
rect 1254 344 1260 345
rect 1302 349 1308 350
rect 1302 345 1303 349
rect 1307 345 1308 349
rect 1302 344 1308 345
rect 1350 349 1356 350
rect 1350 345 1351 349
rect 1355 345 1356 349
rect 1350 344 1356 345
rect 1398 349 1404 350
rect 1398 345 1399 349
rect 1403 345 1404 349
rect 1398 344 1404 345
rect 1446 349 1452 350
rect 1446 345 1447 349
rect 1451 345 1452 349
rect 1446 344 1452 345
rect 1494 349 1500 350
rect 1494 345 1495 349
rect 1499 345 1500 349
rect 1494 344 1500 345
rect 1542 349 1548 350
rect 1542 345 1543 349
rect 1547 345 1548 349
rect 1542 344 1548 345
rect 1590 349 1596 350
rect 1590 345 1591 349
rect 1595 345 1596 349
rect 1590 344 1596 345
rect 1622 349 1628 350
rect 1622 345 1623 349
rect 1627 345 1628 349
rect 1662 347 1663 351
rect 1667 347 1668 351
rect 1662 346 1668 347
rect 1622 344 1628 345
rect 134 335 140 336
rect 110 333 116 334
rect 110 329 111 333
rect 115 329 116 333
rect 134 331 135 335
rect 139 331 140 335
rect 134 330 140 331
rect 166 335 172 336
rect 166 331 167 335
rect 171 331 172 335
rect 166 330 172 331
rect 206 335 212 336
rect 206 331 207 335
rect 211 331 212 335
rect 206 330 212 331
rect 262 335 268 336
rect 262 331 263 335
rect 267 331 268 335
rect 262 330 268 331
rect 326 335 332 336
rect 326 331 327 335
rect 331 331 332 335
rect 326 330 332 331
rect 390 335 396 336
rect 390 331 391 335
rect 395 331 396 335
rect 390 330 396 331
rect 454 335 460 336
rect 454 331 455 335
rect 459 331 460 335
rect 454 330 460 331
rect 518 335 524 336
rect 518 331 519 335
rect 523 331 524 335
rect 518 330 524 331
rect 574 335 580 336
rect 574 331 575 335
rect 579 331 580 335
rect 574 330 580 331
rect 630 335 636 336
rect 630 331 631 335
rect 635 331 636 335
rect 630 330 636 331
rect 686 335 692 336
rect 686 331 687 335
rect 691 331 692 335
rect 686 330 692 331
rect 750 335 756 336
rect 750 331 751 335
rect 755 331 756 335
rect 750 330 756 331
rect 814 335 820 336
rect 814 331 815 335
rect 819 331 820 335
rect 814 330 820 331
rect 878 335 884 336
rect 878 331 879 335
rect 883 331 884 335
rect 878 330 884 331
rect 950 335 956 336
rect 950 331 951 335
rect 955 331 956 335
rect 950 330 956 331
rect 1030 335 1036 336
rect 1030 331 1031 335
rect 1035 331 1036 335
rect 1030 330 1036 331
rect 1110 335 1116 336
rect 1110 331 1111 335
rect 1115 331 1116 335
rect 1110 330 1116 331
rect 1190 335 1196 336
rect 1190 331 1191 335
rect 1195 331 1196 335
rect 1190 330 1196 331
rect 1270 335 1276 336
rect 1270 331 1271 335
rect 1275 331 1276 335
rect 1270 330 1276 331
rect 1342 335 1348 336
rect 1342 331 1343 335
rect 1347 331 1348 335
rect 1342 330 1348 331
rect 1406 335 1412 336
rect 1406 331 1407 335
rect 1411 331 1412 335
rect 1406 330 1412 331
rect 1462 335 1468 336
rect 1462 331 1463 335
rect 1467 331 1468 335
rect 1462 330 1468 331
rect 1518 335 1524 336
rect 1518 331 1519 335
rect 1523 331 1524 335
rect 1518 330 1524 331
rect 1582 335 1588 336
rect 1582 331 1583 335
rect 1587 331 1588 335
rect 1582 330 1588 331
rect 1622 335 1628 336
rect 1622 331 1623 335
rect 1627 331 1628 335
rect 1622 330 1628 331
rect 1662 333 1668 334
rect 110 328 116 329
rect 1662 329 1663 333
rect 1667 329 1668 333
rect 1662 328 1668 329
rect 134 318 140 319
rect 110 316 116 317
rect 110 312 111 316
rect 115 312 116 316
rect 134 314 135 318
rect 139 314 140 318
rect 134 313 140 314
rect 166 318 172 319
rect 166 314 167 318
rect 171 314 172 318
rect 166 313 172 314
rect 206 318 212 319
rect 206 314 207 318
rect 211 314 212 318
rect 206 313 212 314
rect 262 318 268 319
rect 262 314 263 318
rect 267 314 268 318
rect 262 313 268 314
rect 326 318 332 319
rect 326 314 327 318
rect 331 314 332 318
rect 326 313 332 314
rect 390 318 396 319
rect 390 314 391 318
rect 395 314 396 318
rect 390 313 396 314
rect 454 318 460 319
rect 454 314 455 318
rect 459 314 460 318
rect 454 313 460 314
rect 518 318 524 319
rect 518 314 519 318
rect 523 314 524 318
rect 518 313 524 314
rect 574 318 580 319
rect 574 314 575 318
rect 579 314 580 318
rect 574 313 580 314
rect 630 318 636 319
rect 630 314 631 318
rect 635 314 636 318
rect 630 313 636 314
rect 686 318 692 319
rect 686 314 687 318
rect 691 314 692 318
rect 686 313 692 314
rect 750 318 756 319
rect 750 314 751 318
rect 755 314 756 318
rect 750 313 756 314
rect 814 318 820 319
rect 814 314 815 318
rect 819 314 820 318
rect 814 313 820 314
rect 878 318 884 319
rect 878 314 879 318
rect 883 314 884 318
rect 878 313 884 314
rect 950 318 956 319
rect 950 314 951 318
rect 955 314 956 318
rect 950 313 956 314
rect 1030 318 1036 319
rect 1030 314 1031 318
rect 1035 314 1036 318
rect 1030 313 1036 314
rect 1110 318 1116 319
rect 1110 314 1111 318
rect 1115 314 1116 318
rect 1110 313 1116 314
rect 1190 318 1196 319
rect 1190 314 1191 318
rect 1195 314 1196 318
rect 1190 313 1196 314
rect 1270 318 1276 319
rect 1270 314 1271 318
rect 1275 314 1276 318
rect 1270 313 1276 314
rect 1342 318 1348 319
rect 1342 314 1343 318
rect 1347 314 1348 318
rect 1342 313 1348 314
rect 1406 318 1412 319
rect 1406 314 1407 318
rect 1411 314 1412 318
rect 1406 313 1412 314
rect 1462 318 1468 319
rect 1462 314 1463 318
rect 1467 314 1468 318
rect 1462 313 1468 314
rect 1518 318 1524 319
rect 1518 314 1519 318
rect 1523 314 1524 318
rect 1518 313 1524 314
rect 1582 318 1588 319
rect 1582 314 1583 318
rect 1587 314 1588 318
rect 1582 313 1588 314
rect 1622 318 1628 319
rect 1622 314 1623 318
rect 1627 314 1628 318
rect 1622 313 1628 314
rect 1662 316 1668 317
rect 110 311 116 312
rect 1662 312 1663 316
rect 1667 312 1668 316
rect 1662 311 1668 312
rect 110 288 116 289
rect 110 284 111 288
rect 115 284 116 288
rect 1662 288 1668 289
rect 110 283 116 284
rect 134 286 140 287
rect 134 282 135 286
rect 139 282 140 286
rect 134 281 140 282
rect 166 286 172 287
rect 166 282 167 286
rect 171 282 172 286
rect 166 281 172 282
rect 230 286 236 287
rect 230 282 231 286
rect 235 282 236 286
rect 230 281 236 282
rect 294 286 300 287
rect 294 282 295 286
rect 299 282 300 286
rect 294 281 300 282
rect 366 286 372 287
rect 366 282 367 286
rect 371 282 372 286
rect 366 281 372 282
rect 438 286 444 287
rect 438 282 439 286
rect 443 282 444 286
rect 438 281 444 282
rect 502 286 508 287
rect 502 282 503 286
rect 507 282 508 286
rect 502 281 508 282
rect 566 286 572 287
rect 566 282 567 286
rect 571 282 572 286
rect 566 281 572 282
rect 630 286 636 287
rect 630 282 631 286
rect 635 282 636 286
rect 630 281 636 282
rect 686 286 692 287
rect 686 282 687 286
rect 691 282 692 286
rect 686 281 692 282
rect 742 286 748 287
rect 742 282 743 286
rect 747 282 748 286
rect 742 281 748 282
rect 806 286 812 287
rect 806 282 807 286
rect 811 282 812 286
rect 806 281 812 282
rect 878 286 884 287
rect 878 282 879 286
rect 883 282 884 286
rect 878 281 884 282
rect 950 286 956 287
rect 950 282 951 286
rect 955 282 956 286
rect 950 281 956 282
rect 1030 286 1036 287
rect 1030 282 1031 286
rect 1035 282 1036 286
rect 1030 281 1036 282
rect 1110 286 1116 287
rect 1110 282 1111 286
rect 1115 282 1116 286
rect 1110 281 1116 282
rect 1190 286 1196 287
rect 1190 282 1191 286
rect 1195 282 1196 286
rect 1190 281 1196 282
rect 1262 286 1268 287
rect 1262 282 1263 286
rect 1267 282 1268 286
rect 1262 281 1268 282
rect 1326 286 1332 287
rect 1326 282 1327 286
rect 1331 282 1332 286
rect 1326 281 1332 282
rect 1390 286 1396 287
rect 1390 282 1391 286
rect 1395 282 1396 286
rect 1390 281 1396 282
rect 1446 286 1452 287
rect 1446 282 1447 286
rect 1451 282 1452 286
rect 1446 281 1452 282
rect 1494 286 1500 287
rect 1494 282 1495 286
rect 1499 282 1500 286
rect 1494 281 1500 282
rect 1542 286 1548 287
rect 1542 282 1543 286
rect 1547 282 1548 286
rect 1542 281 1548 282
rect 1590 286 1596 287
rect 1590 282 1591 286
rect 1595 282 1596 286
rect 1590 281 1596 282
rect 1622 286 1628 287
rect 1622 282 1623 286
rect 1627 282 1628 286
rect 1662 284 1663 288
rect 1667 284 1668 288
rect 1662 283 1668 284
rect 1622 281 1628 282
rect 110 271 116 272
rect 110 267 111 271
rect 115 267 116 271
rect 1662 271 1668 272
rect 110 266 116 267
rect 134 269 140 270
rect 134 265 135 269
rect 139 265 140 269
rect 134 264 140 265
rect 166 269 172 270
rect 166 265 167 269
rect 171 265 172 269
rect 166 264 172 265
rect 230 269 236 270
rect 230 265 231 269
rect 235 265 236 269
rect 230 264 236 265
rect 294 269 300 270
rect 294 265 295 269
rect 299 265 300 269
rect 294 264 300 265
rect 366 269 372 270
rect 366 265 367 269
rect 371 265 372 269
rect 366 264 372 265
rect 438 269 444 270
rect 438 265 439 269
rect 443 265 444 269
rect 438 264 444 265
rect 502 269 508 270
rect 502 265 503 269
rect 507 265 508 269
rect 502 264 508 265
rect 566 269 572 270
rect 566 265 567 269
rect 571 265 572 269
rect 566 264 572 265
rect 630 269 636 270
rect 630 265 631 269
rect 635 265 636 269
rect 630 264 636 265
rect 686 269 692 270
rect 686 265 687 269
rect 691 265 692 269
rect 686 264 692 265
rect 742 269 748 270
rect 742 265 743 269
rect 747 265 748 269
rect 742 264 748 265
rect 806 269 812 270
rect 806 265 807 269
rect 811 265 812 269
rect 806 264 812 265
rect 878 269 884 270
rect 878 265 879 269
rect 883 265 884 269
rect 878 264 884 265
rect 950 269 956 270
rect 950 265 951 269
rect 955 265 956 269
rect 950 264 956 265
rect 1030 269 1036 270
rect 1030 265 1031 269
rect 1035 265 1036 269
rect 1030 264 1036 265
rect 1110 269 1116 270
rect 1110 265 1111 269
rect 1115 265 1116 269
rect 1110 264 1116 265
rect 1190 269 1196 270
rect 1190 265 1191 269
rect 1195 265 1196 269
rect 1190 264 1196 265
rect 1262 269 1268 270
rect 1262 265 1263 269
rect 1267 265 1268 269
rect 1262 264 1268 265
rect 1326 269 1332 270
rect 1326 265 1327 269
rect 1331 265 1332 269
rect 1326 264 1332 265
rect 1390 269 1396 270
rect 1390 265 1391 269
rect 1395 265 1396 269
rect 1390 264 1396 265
rect 1446 269 1452 270
rect 1446 265 1447 269
rect 1451 265 1452 269
rect 1446 264 1452 265
rect 1494 269 1500 270
rect 1494 265 1495 269
rect 1499 265 1500 269
rect 1494 264 1500 265
rect 1542 269 1548 270
rect 1542 265 1543 269
rect 1547 265 1548 269
rect 1542 264 1548 265
rect 1590 269 1596 270
rect 1590 265 1591 269
rect 1595 265 1596 269
rect 1590 264 1596 265
rect 1622 269 1628 270
rect 1622 265 1623 269
rect 1627 265 1628 269
rect 1662 267 1663 271
rect 1667 267 1668 271
rect 1662 266 1668 267
rect 1622 264 1628 265
rect 134 251 140 252
rect 110 249 116 250
rect 110 245 111 249
rect 115 245 116 249
rect 134 247 135 251
rect 139 247 140 251
rect 134 246 140 247
rect 174 251 180 252
rect 174 247 175 251
rect 179 247 180 251
rect 174 246 180 247
rect 246 251 252 252
rect 246 247 247 251
rect 251 247 252 251
rect 246 246 252 247
rect 318 251 324 252
rect 318 247 319 251
rect 323 247 324 251
rect 318 246 324 247
rect 382 251 388 252
rect 382 247 383 251
rect 387 247 388 251
rect 382 246 388 247
rect 446 251 452 252
rect 446 247 447 251
rect 451 247 452 251
rect 446 246 452 247
rect 518 251 524 252
rect 518 247 519 251
rect 523 247 524 251
rect 518 246 524 247
rect 590 251 596 252
rect 590 247 591 251
rect 595 247 596 251
rect 590 246 596 247
rect 662 251 668 252
rect 662 247 663 251
rect 667 247 668 251
rect 662 246 668 247
rect 742 251 748 252
rect 742 247 743 251
rect 747 247 748 251
rect 742 246 748 247
rect 822 251 828 252
rect 822 247 823 251
rect 827 247 828 251
rect 822 246 828 247
rect 894 251 900 252
rect 894 247 895 251
rect 899 247 900 251
rect 894 246 900 247
rect 966 251 972 252
rect 966 247 967 251
rect 971 247 972 251
rect 966 246 972 247
rect 1030 251 1036 252
rect 1030 247 1031 251
rect 1035 247 1036 251
rect 1030 246 1036 247
rect 1086 251 1092 252
rect 1086 247 1087 251
rect 1091 247 1092 251
rect 1086 246 1092 247
rect 1142 251 1148 252
rect 1142 247 1143 251
rect 1147 247 1148 251
rect 1142 246 1148 247
rect 1198 251 1204 252
rect 1198 247 1199 251
rect 1203 247 1204 251
rect 1198 246 1204 247
rect 1254 251 1260 252
rect 1254 247 1255 251
rect 1259 247 1260 251
rect 1254 246 1260 247
rect 1310 251 1316 252
rect 1310 247 1311 251
rect 1315 247 1316 251
rect 1310 246 1316 247
rect 1366 251 1372 252
rect 1366 247 1367 251
rect 1371 247 1372 251
rect 1366 246 1372 247
rect 1414 251 1420 252
rect 1414 247 1415 251
rect 1419 247 1420 251
rect 1414 246 1420 247
rect 1462 251 1468 252
rect 1462 247 1463 251
rect 1467 247 1468 251
rect 1462 246 1468 247
rect 1518 251 1524 252
rect 1518 247 1519 251
rect 1523 247 1524 251
rect 1518 246 1524 247
rect 1574 251 1580 252
rect 1574 247 1575 251
rect 1579 247 1580 251
rect 1574 246 1580 247
rect 1622 251 1628 252
rect 1622 247 1623 251
rect 1627 247 1628 251
rect 1622 246 1628 247
rect 1662 249 1668 250
rect 110 244 116 245
rect 1662 245 1663 249
rect 1667 245 1668 249
rect 1662 244 1668 245
rect 134 234 140 235
rect 110 232 116 233
rect 110 228 111 232
rect 115 228 116 232
rect 134 230 135 234
rect 139 230 140 234
rect 134 229 140 230
rect 174 234 180 235
rect 174 230 175 234
rect 179 230 180 234
rect 174 229 180 230
rect 246 234 252 235
rect 246 230 247 234
rect 251 230 252 234
rect 246 229 252 230
rect 318 234 324 235
rect 318 230 319 234
rect 323 230 324 234
rect 318 229 324 230
rect 382 234 388 235
rect 382 230 383 234
rect 387 230 388 234
rect 382 229 388 230
rect 446 234 452 235
rect 446 230 447 234
rect 451 230 452 234
rect 446 229 452 230
rect 518 234 524 235
rect 518 230 519 234
rect 523 230 524 234
rect 518 229 524 230
rect 590 234 596 235
rect 590 230 591 234
rect 595 230 596 234
rect 590 229 596 230
rect 662 234 668 235
rect 662 230 663 234
rect 667 230 668 234
rect 662 229 668 230
rect 742 234 748 235
rect 742 230 743 234
rect 747 230 748 234
rect 742 229 748 230
rect 822 234 828 235
rect 822 230 823 234
rect 827 230 828 234
rect 822 229 828 230
rect 894 234 900 235
rect 894 230 895 234
rect 899 230 900 234
rect 894 229 900 230
rect 966 234 972 235
rect 966 230 967 234
rect 971 230 972 234
rect 966 229 972 230
rect 1030 234 1036 235
rect 1030 230 1031 234
rect 1035 230 1036 234
rect 1030 229 1036 230
rect 1086 234 1092 235
rect 1086 230 1087 234
rect 1091 230 1092 234
rect 1086 229 1092 230
rect 1142 234 1148 235
rect 1142 230 1143 234
rect 1147 230 1148 234
rect 1142 229 1148 230
rect 1198 234 1204 235
rect 1198 230 1199 234
rect 1203 230 1204 234
rect 1198 229 1204 230
rect 1254 234 1260 235
rect 1254 230 1255 234
rect 1259 230 1260 234
rect 1254 229 1260 230
rect 1310 234 1316 235
rect 1310 230 1311 234
rect 1315 230 1316 234
rect 1310 229 1316 230
rect 1366 234 1372 235
rect 1366 230 1367 234
rect 1371 230 1372 234
rect 1366 229 1372 230
rect 1414 234 1420 235
rect 1414 230 1415 234
rect 1419 230 1420 234
rect 1414 229 1420 230
rect 1462 234 1468 235
rect 1462 230 1463 234
rect 1467 230 1468 234
rect 1462 229 1468 230
rect 1518 234 1524 235
rect 1518 230 1519 234
rect 1523 230 1524 234
rect 1518 229 1524 230
rect 1574 234 1580 235
rect 1574 230 1575 234
rect 1579 230 1580 234
rect 1574 229 1580 230
rect 1622 234 1628 235
rect 1622 230 1623 234
rect 1627 230 1628 234
rect 1622 229 1628 230
rect 1662 232 1668 233
rect 110 227 116 228
rect 1662 228 1663 232
rect 1667 228 1668 232
rect 1662 227 1668 228
rect 110 204 116 205
rect 110 200 111 204
rect 115 200 116 204
rect 1662 204 1668 205
rect 110 199 116 200
rect 134 202 140 203
rect 134 198 135 202
rect 139 198 140 202
rect 134 197 140 198
rect 166 202 172 203
rect 166 198 167 202
rect 171 198 172 202
rect 166 197 172 198
rect 206 202 212 203
rect 206 198 207 202
rect 211 198 212 202
rect 206 197 212 198
rect 254 202 260 203
rect 254 198 255 202
rect 259 198 260 202
rect 254 197 260 198
rect 302 202 308 203
rect 302 198 303 202
rect 307 198 308 202
rect 302 197 308 198
rect 342 202 348 203
rect 342 198 343 202
rect 347 198 348 202
rect 342 197 348 198
rect 374 202 380 203
rect 374 198 375 202
rect 379 198 380 202
rect 374 197 380 198
rect 414 202 420 203
rect 414 198 415 202
rect 419 198 420 202
rect 414 197 420 198
rect 470 202 476 203
rect 470 198 471 202
rect 475 198 476 202
rect 470 197 476 198
rect 534 202 540 203
rect 534 198 535 202
rect 539 198 540 202
rect 534 197 540 198
rect 614 202 620 203
rect 614 198 615 202
rect 619 198 620 202
rect 614 197 620 198
rect 694 202 700 203
rect 694 198 695 202
rect 699 198 700 202
rect 694 197 700 198
rect 774 202 780 203
rect 774 198 775 202
rect 779 198 780 202
rect 774 197 780 198
rect 854 202 860 203
rect 854 198 855 202
rect 859 198 860 202
rect 854 197 860 198
rect 926 202 932 203
rect 926 198 927 202
rect 931 198 932 202
rect 926 197 932 198
rect 998 202 1004 203
rect 998 198 999 202
rect 1003 198 1004 202
rect 998 197 1004 198
rect 1070 202 1076 203
rect 1070 198 1071 202
rect 1075 198 1076 202
rect 1070 197 1076 198
rect 1142 202 1148 203
rect 1142 198 1143 202
rect 1147 198 1148 202
rect 1142 197 1148 198
rect 1214 202 1220 203
rect 1214 198 1215 202
rect 1219 198 1220 202
rect 1214 197 1220 198
rect 1286 202 1292 203
rect 1286 198 1287 202
rect 1291 198 1292 202
rect 1286 197 1292 198
rect 1350 202 1356 203
rect 1350 198 1351 202
rect 1355 198 1356 202
rect 1350 197 1356 198
rect 1414 202 1420 203
rect 1414 198 1415 202
rect 1419 198 1420 202
rect 1414 197 1420 198
rect 1470 202 1476 203
rect 1470 198 1471 202
rect 1475 198 1476 202
rect 1470 197 1476 198
rect 1526 202 1532 203
rect 1526 198 1527 202
rect 1531 198 1532 202
rect 1526 197 1532 198
rect 1582 202 1588 203
rect 1582 198 1583 202
rect 1587 198 1588 202
rect 1582 197 1588 198
rect 1622 202 1628 203
rect 1622 198 1623 202
rect 1627 198 1628 202
rect 1662 200 1663 204
rect 1667 200 1668 204
rect 1662 199 1668 200
rect 1622 197 1628 198
rect 110 187 116 188
rect 110 183 111 187
rect 115 183 116 187
rect 1662 187 1668 188
rect 110 182 116 183
rect 134 185 140 186
rect 134 181 135 185
rect 139 181 140 185
rect 134 180 140 181
rect 166 185 172 186
rect 166 181 167 185
rect 171 181 172 185
rect 166 180 172 181
rect 206 185 212 186
rect 206 181 207 185
rect 211 181 212 185
rect 206 180 212 181
rect 254 185 260 186
rect 254 181 255 185
rect 259 181 260 185
rect 254 180 260 181
rect 302 185 308 186
rect 302 181 303 185
rect 307 181 308 185
rect 302 180 308 181
rect 342 185 348 186
rect 342 181 343 185
rect 347 181 348 185
rect 342 180 348 181
rect 374 185 380 186
rect 374 181 375 185
rect 379 181 380 185
rect 374 180 380 181
rect 414 185 420 186
rect 414 181 415 185
rect 419 181 420 185
rect 414 180 420 181
rect 470 185 476 186
rect 470 181 471 185
rect 475 181 476 185
rect 470 180 476 181
rect 534 185 540 186
rect 534 181 535 185
rect 539 181 540 185
rect 534 180 540 181
rect 614 185 620 186
rect 614 181 615 185
rect 619 181 620 185
rect 614 180 620 181
rect 694 185 700 186
rect 694 181 695 185
rect 699 181 700 185
rect 694 180 700 181
rect 774 185 780 186
rect 774 181 775 185
rect 779 181 780 185
rect 774 180 780 181
rect 854 185 860 186
rect 854 181 855 185
rect 859 181 860 185
rect 854 180 860 181
rect 926 185 932 186
rect 926 181 927 185
rect 931 181 932 185
rect 926 180 932 181
rect 998 185 1004 186
rect 998 181 999 185
rect 1003 181 1004 185
rect 998 180 1004 181
rect 1070 185 1076 186
rect 1070 181 1071 185
rect 1075 181 1076 185
rect 1070 180 1076 181
rect 1142 185 1148 186
rect 1142 181 1143 185
rect 1147 181 1148 185
rect 1142 180 1148 181
rect 1214 185 1220 186
rect 1214 181 1215 185
rect 1219 181 1220 185
rect 1214 180 1220 181
rect 1286 185 1292 186
rect 1286 181 1287 185
rect 1291 181 1292 185
rect 1286 180 1292 181
rect 1350 185 1356 186
rect 1350 181 1351 185
rect 1355 181 1356 185
rect 1350 180 1356 181
rect 1414 185 1420 186
rect 1414 181 1415 185
rect 1419 181 1420 185
rect 1414 180 1420 181
rect 1470 185 1476 186
rect 1470 181 1471 185
rect 1475 181 1476 185
rect 1470 180 1476 181
rect 1526 185 1532 186
rect 1526 181 1527 185
rect 1531 181 1532 185
rect 1526 180 1532 181
rect 1582 185 1588 186
rect 1582 181 1583 185
rect 1587 181 1588 185
rect 1582 180 1588 181
rect 1622 185 1628 186
rect 1622 181 1623 185
rect 1627 181 1628 185
rect 1662 183 1663 187
rect 1667 183 1668 187
rect 1662 182 1668 183
rect 1622 180 1628 181
rect 134 171 140 172
rect 110 169 116 170
rect 110 165 111 169
rect 115 165 116 169
rect 134 167 135 171
rect 139 167 140 171
rect 134 166 140 167
rect 174 171 180 172
rect 174 167 175 171
rect 179 167 180 171
rect 174 166 180 167
rect 230 171 236 172
rect 230 167 231 171
rect 235 167 236 171
rect 230 166 236 167
rect 286 171 292 172
rect 286 167 287 171
rect 291 167 292 171
rect 286 166 292 167
rect 342 171 348 172
rect 342 167 343 171
rect 347 167 348 171
rect 342 166 348 167
rect 398 171 404 172
rect 398 167 399 171
rect 403 167 404 171
rect 398 166 404 167
rect 454 171 460 172
rect 454 167 455 171
rect 459 167 460 171
rect 454 166 460 167
rect 510 171 516 172
rect 510 167 511 171
rect 515 167 516 171
rect 510 166 516 167
rect 574 171 580 172
rect 574 167 575 171
rect 579 167 580 171
rect 574 166 580 167
rect 638 171 644 172
rect 638 167 639 171
rect 643 167 644 171
rect 638 166 644 167
rect 702 171 708 172
rect 702 167 703 171
rect 707 167 708 171
rect 702 166 708 167
rect 766 171 772 172
rect 766 167 767 171
rect 771 167 772 171
rect 766 166 772 167
rect 830 171 836 172
rect 830 167 831 171
rect 835 167 836 171
rect 830 166 836 167
rect 894 171 900 172
rect 894 167 895 171
rect 899 167 900 171
rect 894 166 900 167
rect 950 171 956 172
rect 950 167 951 171
rect 955 167 956 171
rect 950 166 956 167
rect 1014 171 1020 172
rect 1014 167 1015 171
rect 1019 167 1020 171
rect 1014 166 1020 167
rect 1078 171 1084 172
rect 1078 167 1079 171
rect 1083 167 1084 171
rect 1078 166 1084 167
rect 1142 171 1148 172
rect 1142 167 1143 171
rect 1147 167 1148 171
rect 1142 166 1148 167
rect 1206 171 1212 172
rect 1206 167 1207 171
rect 1211 167 1212 171
rect 1206 166 1212 167
rect 1278 171 1284 172
rect 1278 167 1279 171
rect 1283 167 1284 171
rect 1278 166 1284 167
rect 1350 171 1356 172
rect 1350 167 1351 171
rect 1355 167 1356 171
rect 1350 166 1356 167
rect 1422 171 1428 172
rect 1422 167 1423 171
rect 1427 167 1428 171
rect 1422 166 1428 167
rect 1494 171 1500 172
rect 1494 167 1495 171
rect 1499 167 1500 171
rect 1494 166 1500 167
rect 1566 171 1572 172
rect 1566 167 1567 171
rect 1571 167 1572 171
rect 1566 166 1572 167
rect 1622 171 1628 172
rect 1622 167 1623 171
rect 1627 167 1628 171
rect 1622 166 1628 167
rect 1662 169 1668 170
rect 110 164 116 165
rect 1662 165 1663 169
rect 1667 165 1668 169
rect 1662 164 1668 165
rect 134 154 140 155
rect 110 152 116 153
rect 110 148 111 152
rect 115 148 116 152
rect 134 150 135 154
rect 139 150 140 154
rect 134 149 140 150
rect 174 154 180 155
rect 174 150 175 154
rect 179 150 180 154
rect 174 149 180 150
rect 230 154 236 155
rect 230 150 231 154
rect 235 150 236 154
rect 230 149 236 150
rect 286 154 292 155
rect 286 150 287 154
rect 291 150 292 154
rect 286 149 292 150
rect 342 154 348 155
rect 342 150 343 154
rect 347 150 348 154
rect 342 149 348 150
rect 398 154 404 155
rect 398 150 399 154
rect 403 150 404 154
rect 398 149 404 150
rect 454 154 460 155
rect 454 150 455 154
rect 459 150 460 154
rect 454 149 460 150
rect 510 154 516 155
rect 510 150 511 154
rect 515 150 516 154
rect 510 149 516 150
rect 574 154 580 155
rect 574 150 575 154
rect 579 150 580 154
rect 574 149 580 150
rect 638 154 644 155
rect 638 150 639 154
rect 643 150 644 154
rect 638 149 644 150
rect 702 154 708 155
rect 702 150 703 154
rect 707 150 708 154
rect 702 149 708 150
rect 766 154 772 155
rect 766 150 767 154
rect 771 150 772 154
rect 766 149 772 150
rect 830 154 836 155
rect 830 150 831 154
rect 835 150 836 154
rect 830 149 836 150
rect 894 154 900 155
rect 894 150 895 154
rect 899 150 900 154
rect 894 149 900 150
rect 950 154 956 155
rect 950 150 951 154
rect 955 150 956 154
rect 950 149 956 150
rect 1014 154 1020 155
rect 1014 150 1015 154
rect 1019 150 1020 154
rect 1014 149 1020 150
rect 1078 154 1084 155
rect 1078 150 1079 154
rect 1083 150 1084 154
rect 1078 149 1084 150
rect 1142 154 1148 155
rect 1142 150 1143 154
rect 1147 150 1148 154
rect 1142 149 1148 150
rect 1206 154 1212 155
rect 1206 150 1207 154
rect 1211 150 1212 154
rect 1206 149 1212 150
rect 1278 154 1284 155
rect 1278 150 1279 154
rect 1283 150 1284 154
rect 1278 149 1284 150
rect 1350 154 1356 155
rect 1350 150 1351 154
rect 1355 150 1356 154
rect 1350 149 1356 150
rect 1422 154 1428 155
rect 1422 150 1423 154
rect 1427 150 1428 154
rect 1422 149 1428 150
rect 1494 154 1500 155
rect 1494 150 1495 154
rect 1499 150 1500 154
rect 1494 149 1500 150
rect 1566 154 1572 155
rect 1566 150 1567 154
rect 1571 150 1572 154
rect 1566 149 1572 150
rect 1622 154 1628 155
rect 1622 150 1623 154
rect 1627 150 1628 154
rect 1622 149 1628 150
rect 1662 152 1668 153
rect 110 147 116 148
rect 1662 148 1663 152
rect 1667 148 1668 152
rect 1662 147 1668 148
rect 110 108 116 109
rect 110 104 111 108
rect 115 104 116 108
rect 1662 108 1668 109
rect 110 103 116 104
rect 134 106 140 107
rect 134 102 135 106
rect 139 102 140 106
rect 134 101 140 102
rect 166 106 172 107
rect 166 102 167 106
rect 171 102 172 106
rect 166 101 172 102
rect 198 106 204 107
rect 198 102 199 106
rect 203 102 204 106
rect 198 101 204 102
rect 230 106 236 107
rect 230 102 231 106
rect 235 102 236 106
rect 230 101 236 102
rect 262 106 268 107
rect 262 102 263 106
rect 267 102 268 106
rect 262 101 268 102
rect 294 106 300 107
rect 294 102 295 106
rect 299 102 300 106
rect 294 101 300 102
rect 326 106 332 107
rect 326 102 327 106
rect 331 102 332 106
rect 326 101 332 102
rect 358 106 364 107
rect 358 102 359 106
rect 363 102 364 106
rect 358 101 364 102
rect 390 106 396 107
rect 390 102 391 106
rect 395 102 396 106
rect 390 101 396 102
rect 422 106 428 107
rect 422 102 423 106
rect 427 102 428 106
rect 422 101 428 102
rect 462 106 468 107
rect 462 102 463 106
rect 467 102 468 106
rect 462 101 468 102
rect 502 106 508 107
rect 502 102 503 106
rect 507 102 508 106
rect 502 101 508 102
rect 542 106 548 107
rect 542 102 543 106
rect 547 102 548 106
rect 542 101 548 102
rect 574 106 580 107
rect 574 102 575 106
rect 579 102 580 106
rect 574 101 580 102
rect 606 106 612 107
rect 606 102 607 106
rect 611 102 612 106
rect 606 101 612 102
rect 638 106 644 107
rect 638 102 639 106
rect 643 102 644 106
rect 638 101 644 102
rect 670 106 676 107
rect 670 102 671 106
rect 675 102 676 106
rect 670 101 676 102
rect 702 106 708 107
rect 702 102 703 106
rect 707 102 708 106
rect 702 101 708 102
rect 734 106 740 107
rect 734 102 735 106
rect 739 102 740 106
rect 734 101 740 102
rect 766 106 772 107
rect 766 102 767 106
rect 771 102 772 106
rect 766 101 772 102
rect 798 106 804 107
rect 798 102 799 106
rect 803 102 804 106
rect 798 101 804 102
rect 830 106 836 107
rect 830 102 831 106
rect 835 102 836 106
rect 830 101 836 102
rect 862 106 868 107
rect 862 102 863 106
rect 867 102 868 106
rect 862 101 868 102
rect 894 106 900 107
rect 894 102 895 106
rect 899 102 900 106
rect 894 101 900 102
rect 934 106 940 107
rect 934 102 935 106
rect 939 102 940 106
rect 934 101 940 102
rect 974 106 980 107
rect 974 102 975 106
rect 979 102 980 106
rect 974 101 980 102
rect 1014 106 1020 107
rect 1014 102 1015 106
rect 1019 102 1020 106
rect 1014 101 1020 102
rect 1062 106 1068 107
rect 1062 102 1063 106
rect 1067 102 1068 106
rect 1062 101 1068 102
rect 1102 106 1108 107
rect 1102 102 1103 106
rect 1107 102 1108 106
rect 1102 101 1108 102
rect 1142 106 1148 107
rect 1142 102 1143 106
rect 1147 102 1148 106
rect 1142 101 1148 102
rect 1182 106 1188 107
rect 1182 102 1183 106
rect 1187 102 1188 106
rect 1182 101 1188 102
rect 1222 106 1228 107
rect 1222 102 1223 106
rect 1227 102 1228 106
rect 1222 101 1228 102
rect 1262 106 1268 107
rect 1262 102 1263 106
rect 1267 102 1268 106
rect 1262 101 1268 102
rect 1294 106 1300 107
rect 1294 102 1295 106
rect 1299 102 1300 106
rect 1294 101 1300 102
rect 1334 106 1340 107
rect 1334 102 1335 106
rect 1339 102 1340 106
rect 1334 101 1340 102
rect 1374 106 1380 107
rect 1374 102 1375 106
rect 1379 102 1380 106
rect 1374 101 1380 102
rect 1414 106 1420 107
rect 1414 102 1415 106
rect 1419 102 1420 106
rect 1414 101 1420 102
rect 1454 106 1460 107
rect 1454 102 1455 106
rect 1459 102 1460 106
rect 1454 101 1460 102
rect 1502 106 1508 107
rect 1502 102 1503 106
rect 1507 102 1508 106
rect 1502 101 1508 102
rect 1550 106 1556 107
rect 1550 102 1551 106
rect 1555 102 1556 106
rect 1550 101 1556 102
rect 1590 106 1596 107
rect 1590 102 1591 106
rect 1595 102 1596 106
rect 1590 101 1596 102
rect 1622 106 1628 107
rect 1622 102 1623 106
rect 1627 102 1628 106
rect 1662 104 1663 108
rect 1667 104 1668 108
rect 1662 103 1668 104
rect 1622 101 1628 102
rect 110 91 116 92
rect 110 87 111 91
rect 115 87 116 91
rect 1662 91 1668 92
rect 110 86 116 87
rect 134 89 140 90
rect 134 85 135 89
rect 139 85 140 89
rect 134 84 140 85
rect 166 89 172 90
rect 166 85 167 89
rect 171 85 172 89
rect 166 84 172 85
rect 198 89 204 90
rect 198 85 199 89
rect 203 85 204 89
rect 198 84 204 85
rect 230 89 236 90
rect 230 85 231 89
rect 235 85 236 89
rect 230 84 236 85
rect 262 89 268 90
rect 262 85 263 89
rect 267 85 268 89
rect 262 84 268 85
rect 294 89 300 90
rect 294 85 295 89
rect 299 85 300 89
rect 294 84 300 85
rect 326 89 332 90
rect 326 85 327 89
rect 331 85 332 89
rect 326 84 332 85
rect 358 89 364 90
rect 358 85 359 89
rect 363 85 364 89
rect 358 84 364 85
rect 390 89 396 90
rect 390 85 391 89
rect 395 85 396 89
rect 390 84 396 85
rect 422 89 428 90
rect 422 85 423 89
rect 427 85 428 89
rect 422 84 428 85
rect 462 89 468 90
rect 462 85 463 89
rect 467 85 468 89
rect 462 84 468 85
rect 502 89 508 90
rect 502 85 503 89
rect 507 85 508 89
rect 502 84 508 85
rect 542 89 548 90
rect 542 85 543 89
rect 547 85 548 89
rect 542 84 548 85
rect 574 89 580 90
rect 574 85 575 89
rect 579 85 580 89
rect 574 84 580 85
rect 606 89 612 90
rect 606 85 607 89
rect 611 85 612 89
rect 606 84 612 85
rect 638 89 644 90
rect 638 85 639 89
rect 643 85 644 89
rect 638 84 644 85
rect 670 89 676 90
rect 670 85 671 89
rect 675 85 676 89
rect 670 84 676 85
rect 702 89 708 90
rect 702 85 703 89
rect 707 85 708 89
rect 702 84 708 85
rect 734 89 740 90
rect 734 85 735 89
rect 739 85 740 89
rect 734 84 740 85
rect 766 89 772 90
rect 766 85 767 89
rect 771 85 772 89
rect 766 84 772 85
rect 798 89 804 90
rect 798 85 799 89
rect 803 85 804 89
rect 798 84 804 85
rect 830 89 836 90
rect 830 85 831 89
rect 835 85 836 89
rect 830 84 836 85
rect 862 89 868 90
rect 862 85 863 89
rect 867 85 868 89
rect 862 84 868 85
rect 894 89 900 90
rect 894 85 895 89
rect 899 85 900 89
rect 894 84 900 85
rect 934 89 940 90
rect 934 85 935 89
rect 939 85 940 89
rect 934 84 940 85
rect 974 89 980 90
rect 974 85 975 89
rect 979 85 980 89
rect 974 84 980 85
rect 1014 89 1020 90
rect 1014 85 1015 89
rect 1019 85 1020 89
rect 1014 84 1020 85
rect 1062 89 1068 90
rect 1062 85 1063 89
rect 1067 85 1068 89
rect 1062 84 1068 85
rect 1102 89 1108 90
rect 1102 85 1103 89
rect 1107 85 1108 89
rect 1102 84 1108 85
rect 1142 89 1148 90
rect 1142 85 1143 89
rect 1147 85 1148 89
rect 1142 84 1148 85
rect 1182 89 1188 90
rect 1182 85 1183 89
rect 1187 85 1188 89
rect 1182 84 1188 85
rect 1222 89 1228 90
rect 1222 85 1223 89
rect 1227 85 1228 89
rect 1222 84 1228 85
rect 1262 89 1268 90
rect 1262 85 1263 89
rect 1267 85 1268 89
rect 1262 84 1268 85
rect 1294 89 1300 90
rect 1294 85 1295 89
rect 1299 85 1300 89
rect 1294 84 1300 85
rect 1334 89 1340 90
rect 1334 85 1335 89
rect 1339 85 1340 89
rect 1334 84 1340 85
rect 1374 89 1380 90
rect 1374 85 1375 89
rect 1379 85 1380 89
rect 1374 84 1380 85
rect 1414 89 1420 90
rect 1414 85 1415 89
rect 1419 85 1420 89
rect 1414 84 1420 85
rect 1454 89 1460 90
rect 1454 85 1455 89
rect 1459 85 1460 89
rect 1454 84 1460 85
rect 1502 89 1508 90
rect 1502 85 1503 89
rect 1507 85 1508 89
rect 1502 84 1508 85
rect 1550 89 1556 90
rect 1550 85 1551 89
rect 1555 85 1556 89
rect 1550 84 1556 85
rect 1590 89 1596 90
rect 1590 85 1591 89
rect 1595 85 1596 89
rect 1590 84 1596 85
rect 1622 89 1628 90
rect 1622 85 1623 89
rect 1627 85 1628 89
rect 1662 87 1663 91
rect 1667 87 1668 91
rect 1662 86 1668 87
rect 1622 84 1628 85
<< m3c >>
rect 111 1700 115 1704
rect 255 1698 259 1702
rect 287 1698 291 1702
rect 319 1698 323 1702
rect 359 1698 363 1702
rect 407 1698 411 1702
rect 455 1698 459 1702
rect 503 1698 507 1702
rect 551 1698 555 1702
rect 607 1698 611 1702
rect 663 1698 667 1702
rect 727 1698 731 1702
rect 783 1698 787 1702
rect 839 1698 843 1702
rect 895 1698 899 1702
rect 951 1698 955 1702
rect 1007 1698 1011 1702
rect 1063 1698 1067 1702
rect 1119 1698 1123 1702
rect 1175 1698 1179 1702
rect 1231 1698 1235 1702
rect 1287 1698 1291 1702
rect 1335 1698 1339 1702
rect 1375 1698 1379 1702
rect 1423 1698 1427 1702
rect 1471 1698 1475 1702
rect 1519 1698 1523 1702
rect 1663 1700 1667 1704
rect 111 1683 115 1687
rect 255 1681 259 1685
rect 287 1681 291 1685
rect 319 1681 323 1685
rect 359 1681 363 1685
rect 407 1681 411 1685
rect 455 1681 459 1685
rect 503 1681 507 1685
rect 551 1681 555 1685
rect 607 1681 611 1685
rect 663 1681 667 1685
rect 727 1681 731 1685
rect 783 1681 787 1685
rect 839 1681 843 1685
rect 895 1681 899 1685
rect 951 1681 955 1685
rect 1007 1681 1011 1685
rect 1063 1681 1067 1685
rect 1119 1681 1123 1685
rect 1175 1681 1179 1685
rect 1231 1681 1235 1685
rect 1287 1681 1291 1685
rect 1335 1681 1339 1685
rect 1375 1681 1379 1685
rect 1423 1681 1427 1685
rect 1471 1681 1475 1685
rect 1519 1681 1523 1685
rect 1663 1683 1667 1687
rect 111 1665 115 1669
rect 135 1667 139 1671
rect 167 1667 171 1671
rect 215 1667 219 1671
rect 279 1667 283 1671
rect 343 1667 347 1671
rect 415 1667 419 1671
rect 487 1667 491 1671
rect 559 1667 563 1671
rect 631 1667 635 1671
rect 711 1667 715 1671
rect 791 1667 795 1671
rect 871 1667 875 1671
rect 951 1667 955 1671
rect 1031 1667 1035 1671
rect 1103 1667 1107 1671
rect 1175 1667 1179 1671
rect 1247 1667 1251 1671
rect 1319 1667 1323 1671
rect 1391 1667 1395 1671
rect 1455 1667 1459 1671
rect 1519 1667 1523 1671
rect 1583 1667 1587 1671
rect 1623 1667 1627 1671
rect 1663 1665 1667 1669
rect 111 1648 115 1652
rect 135 1650 139 1654
rect 167 1650 171 1654
rect 215 1650 219 1654
rect 279 1650 283 1654
rect 343 1650 347 1654
rect 415 1650 419 1654
rect 487 1650 491 1654
rect 559 1650 563 1654
rect 631 1650 635 1654
rect 711 1650 715 1654
rect 791 1650 795 1654
rect 871 1650 875 1654
rect 951 1650 955 1654
rect 1031 1650 1035 1654
rect 1103 1650 1107 1654
rect 1175 1650 1179 1654
rect 1247 1650 1251 1654
rect 1319 1650 1323 1654
rect 1391 1650 1395 1654
rect 1455 1650 1459 1654
rect 1519 1650 1523 1654
rect 1583 1650 1587 1654
rect 1623 1650 1627 1654
rect 1663 1648 1667 1652
rect 111 1620 115 1624
rect 135 1618 139 1622
rect 183 1618 187 1622
rect 247 1618 251 1622
rect 303 1618 307 1622
rect 359 1618 363 1622
rect 415 1618 419 1622
rect 471 1618 475 1622
rect 535 1618 539 1622
rect 599 1618 603 1622
rect 663 1618 667 1622
rect 727 1618 731 1622
rect 799 1618 803 1622
rect 871 1618 875 1622
rect 943 1618 947 1622
rect 1023 1618 1027 1622
rect 1103 1618 1107 1622
rect 1175 1618 1179 1622
rect 1247 1618 1251 1622
rect 1319 1618 1323 1622
rect 1399 1618 1403 1622
rect 1479 1618 1483 1622
rect 1559 1618 1563 1622
rect 1623 1618 1627 1622
rect 1663 1620 1667 1624
rect 111 1603 115 1607
rect 135 1601 139 1605
rect 183 1601 187 1605
rect 247 1601 251 1605
rect 303 1601 307 1605
rect 359 1601 363 1605
rect 415 1601 419 1605
rect 471 1601 475 1605
rect 535 1601 539 1605
rect 599 1601 603 1605
rect 663 1601 667 1605
rect 727 1601 731 1605
rect 799 1601 803 1605
rect 871 1601 875 1605
rect 943 1601 947 1605
rect 1023 1601 1027 1605
rect 1103 1601 1107 1605
rect 1175 1601 1179 1605
rect 1247 1601 1251 1605
rect 1319 1601 1323 1605
rect 1399 1601 1403 1605
rect 1479 1601 1483 1605
rect 1559 1601 1563 1605
rect 1623 1601 1627 1605
rect 1663 1603 1667 1607
rect 111 1585 115 1589
rect 135 1587 139 1591
rect 167 1587 171 1591
rect 223 1587 227 1591
rect 279 1587 283 1591
rect 335 1587 339 1591
rect 383 1587 387 1591
rect 431 1587 435 1591
rect 479 1587 483 1591
rect 535 1587 539 1591
rect 599 1587 603 1591
rect 663 1587 667 1591
rect 727 1587 731 1591
rect 799 1587 803 1591
rect 871 1587 875 1591
rect 951 1587 955 1591
rect 1039 1587 1043 1591
rect 1119 1587 1123 1591
rect 1199 1587 1203 1591
rect 1279 1587 1283 1591
rect 1351 1587 1355 1591
rect 1415 1587 1419 1591
rect 1471 1587 1475 1591
rect 1527 1587 1531 1591
rect 1583 1587 1587 1591
rect 1623 1587 1627 1591
rect 1663 1585 1667 1589
rect 111 1568 115 1572
rect 135 1570 139 1574
rect 167 1570 171 1574
rect 223 1570 227 1574
rect 279 1570 283 1574
rect 335 1570 339 1574
rect 383 1570 387 1574
rect 431 1570 435 1574
rect 479 1570 483 1574
rect 535 1570 539 1574
rect 599 1570 603 1574
rect 663 1570 667 1574
rect 727 1570 731 1574
rect 799 1570 803 1574
rect 871 1570 875 1574
rect 951 1570 955 1574
rect 1039 1570 1043 1574
rect 1119 1570 1123 1574
rect 1199 1570 1203 1574
rect 1279 1570 1283 1574
rect 1351 1570 1355 1574
rect 1415 1570 1419 1574
rect 1471 1570 1475 1574
rect 1527 1570 1531 1574
rect 1583 1570 1587 1574
rect 1623 1570 1627 1574
rect 1663 1568 1667 1572
rect 111 1540 115 1544
rect 135 1538 139 1542
rect 167 1538 171 1542
rect 215 1538 219 1542
rect 263 1538 267 1542
rect 311 1538 315 1542
rect 359 1538 363 1542
rect 407 1538 411 1542
rect 455 1538 459 1542
rect 511 1538 515 1542
rect 567 1538 571 1542
rect 631 1538 635 1542
rect 695 1538 699 1542
rect 759 1538 763 1542
rect 831 1538 835 1542
rect 919 1538 923 1542
rect 1007 1538 1011 1542
rect 1095 1538 1099 1542
rect 1183 1538 1187 1542
rect 1263 1538 1267 1542
rect 1335 1538 1339 1542
rect 1407 1538 1411 1542
rect 1471 1538 1475 1542
rect 1527 1538 1531 1542
rect 1583 1538 1587 1542
rect 1623 1538 1627 1542
rect 1663 1540 1667 1544
rect 111 1523 115 1527
rect 135 1521 139 1525
rect 167 1521 171 1525
rect 215 1521 219 1525
rect 263 1521 267 1525
rect 311 1521 315 1525
rect 359 1521 363 1525
rect 407 1521 411 1525
rect 455 1521 459 1525
rect 511 1521 515 1525
rect 567 1521 571 1525
rect 631 1521 635 1525
rect 695 1521 699 1525
rect 759 1521 763 1525
rect 831 1521 835 1525
rect 919 1521 923 1525
rect 1007 1521 1011 1525
rect 1095 1521 1099 1525
rect 1183 1521 1187 1525
rect 1263 1521 1267 1525
rect 1335 1521 1339 1525
rect 1407 1521 1411 1525
rect 1471 1521 1475 1525
rect 1527 1521 1531 1525
rect 1583 1521 1587 1525
rect 1623 1521 1627 1525
rect 1663 1523 1667 1527
rect 111 1501 115 1505
rect 135 1503 139 1507
rect 167 1503 171 1507
rect 223 1503 227 1507
rect 295 1503 299 1507
rect 375 1503 379 1507
rect 455 1503 459 1507
rect 527 1503 531 1507
rect 599 1503 603 1507
rect 671 1503 675 1507
rect 743 1503 747 1507
rect 815 1503 819 1507
rect 879 1503 883 1507
rect 943 1503 947 1507
rect 1007 1503 1011 1507
rect 1063 1503 1067 1507
rect 1111 1503 1115 1507
rect 1151 1503 1155 1507
rect 1183 1503 1187 1507
rect 1215 1503 1219 1507
rect 1255 1503 1259 1507
rect 1295 1503 1299 1507
rect 1351 1503 1355 1507
rect 1415 1503 1419 1507
rect 1487 1503 1491 1507
rect 1567 1503 1571 1507
rect 1623 1503 1627 1507
rect 1663 1501 1667 1505
rect 111 1484 115 1488
rect 135 1486 139 1490
rect 167 1486 171 1490
rect 223 1486 227 1490
rect 295 1486 299 1490
rect 375 1486 379 1490
rect 455 1486 459 1490
rect 527 1486 531 1490
rect 599 1486 603 1490
rect 671 1486 675 1490
rect 743 1486 747 1490
rect 815 1486 819 1490
rect 879 1486 883 1490
rect 943 1486 947 1490
rect 1007 1486 1011 1490
rect 1063 1486 1067 1490
rect 1111 1486 1115 1490
rect 1151 1486 1155 1490
rect 1183 1486 1187 1490
rect 1215 1486 1219 1490
rect 1255 1486 1259 1490
rect 1295 1486 1299 1490
rect 1351 1486 1355 1490
rect 1415 1486 1419 1490
rect 1487 1486 1491 1490
rect 1567 1486 1571 1490
rect 1623 1486 1627 1490
rect 1663 1484 1667 1488
rect 111 1456 115 1460
rect 135 1454 139 1458
rect 167 1454 171 1458
rect 223 1454 227 1458
rect 295 1454 299 1458
rect 375 1454 379 1458
rect 455 1454 459 1458
rect 527 1454 531 1458
rect 599 1454 603 1458
rect 663 1454 667 1458
rect 719 1454 723 1458
rect 783 1454 787 1458
rect 847 1454 851 1458
rect 903 1454 907 1458
rect 959 1454 963 1458
rect 1015 1454 1019 1458
rect 1071 1454 1075 1458
rect 1119 1454 1123 1458
rect 1159 1454 1163 1458
rect 1207 1454 1211 1458
rect 1263 1454 1267 1458
rect 1327 1454 1331 1458
rect 1399 1454 1403 1458
rect 1479 1454 1483 1458
rect 1559 1454 1563 1458
rect 1623 1454 1627 1458
rect 1663 1456 1667 1460
rect 111 1439 115 1443
rect 135 1437 139 1441
rect 167 1437 171 1441
rect 223 1437 227 1441
rect 295 1437 299 1441
rect 375 1437 379 1441
rect 455 1437 459 1441
rect 527 1437 531 1441
rect 599 1437 603 1441
rect 663 1437 667 1441
rect 719 1437 723 1441
rect 783 1437 787 1441
rect 847 1437 851 1441
rect 903 1437 907 1441
rect 959 1437 963 1441
rect 1015 1437 1019 1441
rect 1071 1437 1075 1441
rect 1119 1437 1123 1441
rect 1159 1437 1163 1441
rect 1207 1437 1211 1441
rect 1263 1437 1267 1441
rect 1327 1437 1331 1441
rect 1399 1437 1403 1441
rect 1479 1437 1483 1441
rect 1559 1437 1563 1441
rect 1623 1437 1627 1441
rect 1663 1439 1667 1443
rect 111 1417 115 1421
rect 135 1419 139 1423
rect 167 1419 171 1423
rect 215 1419 219 1423
rect 287 1419 291 1423
rect 359 1419 363 1423
rect 439 1419 443 1423
rect 519 1419 523 1423
rect 599 1419 603 1423
rect 679 1419 683 1423
rect 759 1419 763 1423
rect 831 1419 835 1423
rect 903 1419 907 1423
rect 967 1419 971 1423
rect 1031 1419 1035 1423
rect 1103 1419 1107 1423
rect 1167 1419 1171 1423
rect 1231 1419 1235 1423
rect 1295 1419 1299 1423
rect 1359 1419 1363 1423
rect 1415 1419 1419 1423
rect 1463 1419 1467 1423
rect 1503 1419 1507 1423
rect 1551 1419 1555 1423
rect 1591 1419 1595 1423
rect 1623 1419 1627 1423
rect 1663 1417 1667 1421
rect 111 1400 115 1404
rect 135 1402 139 1406
rect 167 1402 171 1406
rect 215 1402 219 1406
rect 287 1402 291 1406
rect 359 1402 363 1406
rect 439 1402 443 1406
rect 519 1402 523 1406
rect 599 1402 603 1406
rect 679 1402 683 1406
rect 759 1402 763 1406
rect 831 1402 835 1406
rect 903 1402 907 1406
rect 967 1402 971 1406
rect 1031 1402 1035 1406
rect 1103 1402 1107 1406
rect 1167 1402 1171 1406
rect 1231 1402 1235 1406
rect 1295 1402 1299 1406
rect 1359 1402 1363 1406
rect 1415 1402 1419 1406
rect 1463 1402 1467 1406
rect 1503 1402 1507 1406
rect 1551 1402 1555 1406
rect 1591 1402 1595 1406
rect 1623 1402 1627 1406
rect 1663 1400 1667 1404
rect 111 1372 115 1376
rect 135 1370 139 1374
rect 167 1370 171 1374
rect 223 1370 227 1374
rect 287 1370 291 1374
rect 359 1370 363 1374
rect 431 1370 435 1374
rect 503 1370 507 1374
rect 583 1370 587 1374
rect 663 1370 667 1374
rect 743 1370 747 1374
rect 815 1370 819 1374
rect 887 1370 891 1374
rect 959 1370 963 1374
rect 1031 1370 1035 1374
rect 1103 1370 1107 1374
rect 1175 1370 1179 1374
rect 1239 1370 1243 1374
rect 1303 1370 1307 1374
rect 1367 1370 1371 1374
rect 1431 1370 1435 1374
rect 1495 1370 1499 1374
rect 1567 1370 1571 1374
rect 1623 1370 1627 1374
rect 1663 1372 1667 1376
rect 111 1355 115 1359
rect 135 1353 139 1357
rect 167 1353 171 1357
rect 223 1353 227 1357
rect 287 1353 291 1357
rect 359 1353 363 1357
rect 431 1353 435 1357
rect 503 1353 507 1357
rect 583 1353 587 1357
rect 663 1353 667 1357
rect 743 1353 747 1357
rect 815 1353 819 1357
rect 887 1353 891 1357
rect 959 1353 963 1357
rect 1031 1353 1035 1357
rect 1103 1353 1107 1357
rect 1175 1353 1179 1357
rect 1239 1353 1243 1357
rect 1303 1353 1307 1357
rect 1367 1353 1371 1357
rect 1431 1353 1435 1357
rect 1495 1353 1499 1357
rect 1567 1353 1571 1357
rect 1623 1353 1627 1357
rect 1663 1355 1667 1359
rect 111 1337 115 1341
rect 135 1339 139 1343
rect 183 1339 187 1343
rect 239 1339 243 1343
rect 295 1339 299 1343
rect 351 1339 355 1343
rect 399 1339 403 1343
rect 455 1339 459 1343
rect 511 1339 515 1343
rect 567 1339 571 1343
rect 631 1339 635 1343
rect 695 1339 699 1343
rect 759 1339 763 1343
rect 823 1339 827 1343
rect 887 1339 891 1343
rect 959 1339 963 1343
rect 1023 1339 1027 1343
rect 1087 1339 1091 1343
rect 1151 1339 1155 1343
rect 1215 1339 1219 1343
rect 1279 1339 1283 1343
rect 1343 1339 1347 1343
rect 1407 1339 1411 1343
rect 1479 1339 1483 1343
rect 1559 1339 1563 1343
rect 1623 1339 1627 1343
rect 1663 1337 1667 1341
rect 111 1320 115 1324
rect 135 1322 139 1326
rect 183 1322 187 1326
rect 239 1322 243 1326
rect 295 1322 299 1326
rect 351 1322 355 1326
rect 399 1322 403 1326
rect 455 1322 459 1326
rect 511 1322 515 1326
rect 567 1322 571 1326
rect 631 1322 635 1326
rect 695 1322 699 1326
rect 759 1322 763 1326
rect 823 1322 827 1326
rect 887 1322 891 1326
rect 959 1322 963 1326
rect 1023 1322 1027 1326
rect 1087 1322 1091 1326
rect 1151 1322 1155 1326
rect 1215 1322 1219 1326
rect 1279 1322 1283 1326
rect 1343 1322 1347 1326
rect 1407 1322 1411 1326
rect 1479 1322 1483 1326
rect 1559 1322 1563 1326
rect 1623 1322 1627 1326
rect 1663 1320 1667 1324
rect 111 1288 115 1292
rect 135 1286 139 1290
rect 183 1286 187 1290
rect 231 1286 235 1290
rect 279 1286 283 1290
rect 327 1286 331 1290
rect 375 1286 379 1290
rect 431 1286 435 1290
rect 487 1286 491 1290
rect 543 1286 547 1290
rect 607 1286 611 1290
rect 663 1286 667 1290
rect 719 1286 723 1290
rect 775 1286 779 1290
rect 831 1286 835 1290
rect 895 1286 899 1290
rect 959 1286 963 1290
rect 1023 1286 1027 1290
rect 1079 1286 1083 1290
rect 1143 1286 1147 1290
rect 1207 1286 1211 1290
rect 1279 1286 1283 1290
rect 1359 1286 1363 1290
rect 1447 1286 1451 1290
rect 1543 1286 1547 1290
rect 1623 1286 1627 1290
rect 1663 1288 1667 1292
rect 111 1271 115 1275
rect 135 1269 139 1273
rect 183 1269 187 1273
rect 231 1269 235 1273
rect 279 1269 283 1273
rect 327 1269 331 1273
rect 375 1269 379 1273
rect 431 1269 435 1273
rect 487 1269 491 1273
rect 543 1269 547 1273
rect 607 1269 611 1273
rect 663 1269 667 1273
rect 719 1269 723 1273
rect 775 1269 779 1273
rect 831 1269 835 1273
rect 895 1269 899 1273
rect 959 1269 963 1273
rect 1023 1269 1027 1273
rect 1079 1269 1083 1273
rect 1143 1269 1147 1273
rect 1207 1269 1211 1273
rect 1279 1269 1283 1273
rect 1359 1269 1363 1273
rect 1447 1269 1451 1273
rect 1543 1269 1547 1273
rect 1623 1269 1627 1273
rect 1663 1271 1667 1275
rect 111 1253 115 1257
rect 135 1255 139 1259
rect 167 1255 171 1259
rect 223 1255 227 1259
rect 279 1255 283 1259
rect 327 1255 331 1259
rect 383 1255 387 1259
rect 439 1255 443 1259
rect 495 1255 499 1259
rect 551 1255 555 1259
rect 607 1255 611 1259
rect 663 1255 667 1259
rect 719 1255 723 1259
rect 767 1255 771 1259
rect 815 1255 819 1259
rect 871 1255 875 1259
rect 927 1255 931 1259
rect 983 1255 987 1259
rect 1039 1255 1043 1259
rect 1095 1255 1099 1259
rect 1159 1255 1163 1259
rect 1231 1255 1235 1259
rect 1319 1255 1323 1259
rect 1423 1255 1427 1259
rect 1535 1255 1539 1259
rect 1623 1255 1627 1259
rect 1663 1253 1667 1257
rect 111 1236 115 1240
rect 135 1238 139 1242
rect 167 1238 171 1242
rect 223 1238 227 1242
rect 279 1238 283 1242
rect 327 1238 331 1242
rect 383 1238 387 1242
rect 439 1238 443 1242
rect 495 1238 499 1242
rect 551 1238 555 1242
rect 607 1238 611 1242
rect 663 1238 667 1242
rect 719 1238 723 1242
rect 767 1238 771 1242
rect 815 1238 819 1242
rect 871 1238 875 1242
rect 927 1238 931 1242
rect 983 1238 987 1242
rect 1039 1238 1043 1242
rect 1095 1238 1099 1242
rect 1159 1238 1163 1242
rect 1231 1238 1235 1242
rect 1319 1238 1323 1242
rect 1423 1238 1427 1242
rect 1535 1238 1539 1242
rect 1623 1238 1627 1242
rect 1663 1236 1667 1240
rect 111 1204 115 1208
rect 135 1202 139 1206
rect 167 1202 171 1206
rect 223 1202 227 1206
rect 279 1202 283 1206
rect 335 1202 339 1206
rect 383 1202 387 1206
rect 431 1202 435 1206
rect 487 1202 491 1206
rect 543 1202 547 1206
rect 599 1202 603 1206
rect 655 1202 659 1206
rect 711 1202 715 1206
rect 767 1202 771 1206
rect 823 1202 827 1206
rect 887 1202 891 1206
rect 951 1202 955 1206
rect 1015 1202 1019 1206
rect 1079 1202 1083 1206
rect 1143 1202 1147 1206
rect 1207 1202 1211 1206
rect 1279 1202 1283 1206
rect 1359 1202 1363 1206
rect 1447 1202 1451 1206
rect 1543 1202 1547 1206
rect 1623 1202 1627 1206
rect 1663 1204 1667 1208
rect 111 1187 115 1191
rect 135 1185 139 1189
rect 167 1185 171 1189
rect 223 1185 227 1189
rect 279 1185 283 1189
rect 335 1185 339 1189
rect 383 1185 387 1189
rect 431 1185 435 1189
rect 487 1185 491 1189
rect 543 1185 547 1189
rect 599 1185 603 1189
rect 655 1185 659 1189
rect 711 1185 715 1189
rect 767 1185 771 1189
rect 823 1185 827 1189
rect 887 1185 891 1189
rect 951 1185 955 1189
rect 1015 1185 1019 1189
rect 1079 1185 1083 1189
rect 1143 1185 1147 1189
rect 1207 1185 1211 1189
rect 1279 1185 1283 1189
rect 1359 1185 1363 1189
rect 1447 1185 1451 1189
rect 1543 1185 1547 1189
rect 1623 1185 1627 1189
rect 1663 1187 1667 1191
rect 111 1165 115 1169
rect 135 1167 139 1171
rect 167 1167 171 1171
rect 223 1167 227 1171
rect 287 1167 291 1171
rect 351 1167 355 1171
rect 415 1167 419 1171
rect 471 1167 475 1171
rect 535 1167 539 1171
rect 599 1167 603 1171
rect 663 1167 667 1171
rect 727 1167 731 1171
rect 783 1167 787 1171
rect 839 1167 843 1171
rect 903 1167 907 1171
rect 967 1167 971 1171
rect 1031 1167 1035 1171
rect 1095 1167 1099 1171
rect 1159 1167 1163 1171
rect 1215 1167 1219 1171
rect 1279 1167 1283 1171
rect 1343 1167 1347 1171
rect 1407 1167 1411 1171
rect 1479 1167 1483 1171
rect 1559 1167 1563 1171
rect 1623 1167 1627 1171
rect 1663 1165 1667 1169
rect 111 1148 115 1152
rect 135 1150 139 1154
rect 167 1150 171 1154
rect 223 1150 227 1154
rect 287 1150 291 1154
rect 351 1150 355 1154
rect 415 1150 419 1154
rect 471 1150 475 1154
rect 535 1150 539 1154
rect 599 1150 603 1154
rect 663 1150 667 1154
rect 727 1150 731 1154
rect 783 1150 787 1154
rect 839 1150 843 1154
rect 903 1150 907 1154
rect 967 1150 971 1154
rect 1031 1150 1035 1154
rect 1095 1150 1099 1154
rect 1159 1150 1163 1154
rect 1215 1150 1219 1154
rect 1279 1150 1283 1154
rect 1343 1150 1347 1154
rect 1407 1150 1411 1154
rect 1479 1150 1483 1154
rect 1559 1150 1563 1154
rect 1623 1150 1627 1154
rect 1663 1148 1667 1152
rect 111 1116 115 1120
rect 143 1114 147 1118
rect 175 1114 179 1118
rect 215 1114 219 1118
rect 271 1114 275 1118
rect 335 1114 339 1118
rect 399 1114 403 1118
rect 463 1114 467 1118
rect 527 1114 531 1118
rect 599 1114 603 1118
rect 663 1114 667 1118
rect 727 1114 731 1118
rect 791 1114 795 1118
rect 855 1114 859 1118
rect 911 1114 915 1118
rect 967 1114 971 1118
rect 1023 1114 1027 1118
rect 1087 1114 1091 1118
rect 1151 1114 1155 1118
rect 1215 1114 1219 1118
rect 1279 1114 1283 1118
rect 1335 1114 1339 1118
rect 1391 1114 1395 1118
rect 1447 1114 1451 1118
rect 1495 1114 1499 1118
rect 1543 1114 1547 1118
rect 1591 1114 1595 1118
rect 1623 1114 1627 1118
rect 1663 1116 1667 1120
rect 111 1099 115 1103
rect 143 1097 147 1101
rect 175 1097 179 1101
rect 215 1097 219 1101
rect 271 1097 275 1101
rect 335 1097 339 1101
rect 399 1097 403 1101
rect 463 1097 467 1101
rect 527 1097 531 1101
rect 599 1097 603 1101
rect 663 1097 667 1101
rect 727 1097 731 1101
rect 791 1097 795 1101
rect 855 1097 859 1101
rect 911 1097 915 1101
rect 967 1097 971 1101
rect 1023 1097 1027 1101
rect 1087 1097 1091 1101
rect 1151 1097 1155 1101
rect 1215 1097 1219 1101
rect 1279 1097 1283 1101
rect 1335 1097 1339 1101
rect 1391 1097 1395 1101
rect 1447 1097 1451 1101
rect 1495 1097 1499 1101
rect 1543 1097 1547 1101
rect 1591 1097 1595 1101
rect 1623 1097 1627 1101
rect 1663 1099 1667 1103
rect 111 1077 115 1081
rect 215 1079 219 1083
rect 247 1079 251 1083
rect 279 1079 283 1083
rect 311 1079 315 1083
rect 351 1079 355 1083
rect 391 1079 395 1083
rect 439 1079 443 1083
rect 503 1079 507 1083
rect 575 1079 579 1083
rect 655 1079 659 1083
rect 735 1079 739 1083
rect 815 1079 819 1083
rect 895 1079 899 1083
rect 967 1079 971 1083
rect 1039 1079 1043 1083
rect 1111 1079 1115 1083
rect 1175 1079 1179 1083
rect 1239 1079 1243 1083
rect 1303 1079 1307 1083
rect 1359 1079 1363 1083
rect 1415 1079 1419 1083
rect 1463 1079 1467 1083
rect 1503 1079 1507 1083
rect 1551 1079 1555 1083
rect 1591 1079 1595 1083
rect 1623 1079 1627 1083
rect 1663 1077 1667 1081
rect 111 1060 115 1064
rect 215 1062 219 1066
rect 247 1062 251 1066
rect 279 1062 283 1066
rect 311 1062 315 1066
rect 351 1062 355 1066
rect 391 1062 395 1066
rect 439 1062 443 1066
rect 503 1062 507 1066
rect 575 1062 579 1066
rect 655 1062 659 1066
rect 735 1062 739 1066
rect 815 1062 819 1066
rect 895 1062 899 1066
rect 967 1062 971 1066
rect 1039 1062 1043 1066
rect 1111 1062 1115 1066
rect 1175 1062 1179 1066
rect 1239 1062 1243 1066
rect 1303 1062 1307 1066
rect 1359 1062 1363 1066
rect 1415 1062 1419 1066
rect 1463 1062 1467 1066
rect 1503 1062 1507 1066
rect 1551 1062 1555 1066
rect 1591 1062 1595 1066
rect 1623 1062 1627 1066
rect 1663 1060 1667 1064
rect 111 1028 115 1032
rect 295 1026 299 1030
rect 327 1026 331 1030
rect 359 1026 363 1030
rect 391 1026 395 1030
rect 423 1026 427 1030
rect 455 1026 459 1030
rect 503 1026 507 1030
rect 559 1026 563 1030
rect 631 1026 635 1030
rect 711 1026 715 1030
rect 799 1026 803 1030
rect 879 1026 883 1030
rect 959 1026 963 1030
rect 1031 1026 1035 1030
rect 1095 1026 1099 1030
rect 1159 1026 1163 1030
rect 1223 1026 1227 1030
rect 1279 1026 1283 1030
rect 1335 1026 1339 1030
rect 1383 1026 1387 1030
rect 1431 1026 1435 1030
rect 1479 1026 1483 1030
rect 1535 1026 1539 1030
rect 1591 1026 1595 1030
rect 1623 1026 1627 1030
rect 1663 1028 1667 1032
rect 111 1011 115 1015
rect 295 1009 299 1013
rect 327 1009 331 1013
rect 359 1009 363 1013
rect 391 1009 395 1013
rect 423 1009 427 1013
rect 455 1009 459 1013
rect 503 1009 507 1013
rect 559 1009 563 1013
rect 631 1009 635 1013
rect 711 1009 715 1013
rect 799 1009 803 1013
rect 879 1009 883 1013
rect 959 1009 963 1013
rect 1031 1009 1035 1013
rect 1095 1009 1099 1013
rect 1159 1009 1163 1013
rect 1223 1009 1227 1013
rect 1279 1009 1283 1013
rect 1335 1009 1339 1013
rect 1383 1009 1387 1013
rect 1431 1009 1435 1013
rect 1479 1009 1483 1013
rect 1535 1009 1539 1013
rect 1591 1009 1595 1013
rect 1623 1009 1627 1013
rect 1663 1011 1667 1015
rect 111 993 115 997
rect 247 995 251 999
rect 279 995 283 999
rect 311 995 315 999
rect 343 995 347 999
rect 383 995 387 999
rect 423 995 427 999
rect 479 995 483 999
rect 543 995 547 999
rect 615 995 619 999
rect 687 995 691 999
rect 759 995 763 999
rect 831 995 835 999
rect 903 995 907 999
rect 967 995 971 999
rect 1031 995 1035 999
rect 1095 995 1099 999
rect 1159 995 1163 999
rect 1223 995 1227 999
rect 1287 995 1291 999
rect 1343 995 1347 999
rect 1399 995 1403 999
rect 1447 995 1451 999
rect 1495 995 1499 999
rect 1543 995 1547 999
rect 1591 995 1595 999
rect 1623 995 1627 999
rect 1663 993 1667 997
rect 111 976 115 980
rect 247 978 251 982
rect 279 978 283 982
rect 311 978 315 982
rect 343 978 347 982
rect 383 978 387 982
rect 423 978 427 982
rect 479 978 483 982
rect 543 978 547 982
rect 615 978 619 982
rect 687 978 691 982
rect 759 978 763 982
rect 831 978 835 982
rect 903 978 907 982
rect 967 978 971 982
rect 1031 978 1035 982
rect 1095 978 1099 982
rect 1159 978 1163 982
rect 1223 978 1227 982
rect 1287 978 1291 982
rect 1343 978 1347 982
rect 1399 978 1403 982
rect 1447 978 1451 982
rect 1495 978 1499 982
rect 1543 978 1547 982
rect 1591 978 1595 982
rect 1623 978 1627 982
rect 1663 976 1667 980
rect 111 948 115 952
rect 167 946 171 950
rect 199 946 203 950
rect 239 946 243 950
rect 287 946 291 950
rect 343 946 347 950
rect 407 946 411 950
rect 471 946 475 950
rect 535 946 539 950
rect 599 946 603 950
rect 663 946 667 950
rect 727 946 731 950
rect 791 946 795 950
rect 847 946 851 950
rect 911 946 915 950
rect 975 946 979 950
rect 1039 946 1043 950
rect 1103 946 1107 950
rect 1167 946 1171 950
rect 1231 946 1235 950
rect 1287 946 1291 950
rect 1343 946 1347 950
rect 1391 946 1395 950
rect 1431 946 1435 950
rect 1471 946 1475 950
rect 1511 946 1515 950
rect 1551 946 1555 950
rect 1591 946 1595 950
rect 1623 946 1627 950
rect 1663 948 1667 952
rect 111 931 115 935
rect 167 929 171 933
rect 199 929 203 933
rect 239 929 243 933
rect 287 929 291 933
rect 343 929 347 933
rect 407 929 411 933
rect 471 929 475 933
rect 535 929 539 933
rect 599 929 603 933
rect 663 929 667 933
rect 727 929 731 933
rect 791 929 795 933
rect 847 929 851 933
rect 911 929 915 933
rect 975 929 979 933
rect 1039 929 1043 933
rect 1103 929 1107 933
rect 1167 929 1171 933
rect 1231 929 1235 933
rect 1287 929 1291 933
rect 1343 929 1347 933
rect 1391 929 1395 933
rect 1431 929 1435 933
rect 1471 929 1475 933
rect 1511 929 1515 933
rect 1551 929 1555 933
rect 1591 929 1595 933
rect 1623 929 1627 933
rect 1663 931 1667 935
rect 111 909 115 913
rect 135 911 139 915
rect 167 911 171 915
rect 207 911 211 915
rect 271 911 275 915
rect 335 911 339 915
rect 407 911 411 915
rect 471 911 475 915
rect 535 911 539 915
rect 591 911 595 915
rect 647 911 651 915
rect 703 911 707 915
rect 751 911 755 915
rect 799 911 803 915
rect 847 911 851 915
rect 903 911 907 915
rect 959 911 963 915
rect 1023 911 1027 915
rect 1087 911 1091 915
rect 1143 911 1147 915
rect 1199 911 1203 915
rect 1255 911 1259 915
rect 1319 911 1323 915
rect 1383 911 1387 915
rect 1663 909 1667 913
rect 111 892 115 896
rect 135 894 139 898
rect 167 894 171 898
rect 207 894 211 898
rect 271 894 275 898
rect 335 894 339 898
rect 407 894 411 898
rect 471 894 475 898
rect 535 894 539 898
rect 591 894 595 898
rect 647 894 651 898
rect 703 894 707 898
rect 751 894 755 898
rect 799 894 803 898
rect 847 894 851 898
rect 903 894 907 898
rect 959 894 963 898
rect 1023 894 1027 898
rect 1087 894 1091 898
rect 1143 894 1147 898
rect 1199 894 1203 898
rect 1255 894 1259 898
rect 1319 894 1323 898
rect 1383 894 1387 898
rect 1663 892 1667 896
rect 111 860 115 864
rect 135 858 139 862
rect 167 858 171 862
rect 207 858 211 862
rect 271 858 275 862
rect 335 858 339 862
rect 407 858 411 862
rect 471 858 475 862
rect 535 858 539 862
rect 599 858 603 862
rect 655 858 659 862
rect 703 858 707 862
rect 751 858 755 862
rect 799 858 803 862
rect 847 858 851 862
rect 903 858 907 862
rect 967 858 971 862
rect 1039 858 1043 862
rect 1103 858 1107 862
rect 1167 858 1171 862
rect 1231 858 1235 862
rect 1287 858 1291 862
rect 1343 858 1347 862
rect 1399 858 1403 862
rect 1463 858 1467 862
rect 1663 860 1667 864
rect 111 843 115 847
rect 135 841 139 845
rect 167 841 171 845
rect 207 841 211 845
rect 271 841 275 845
rect 335 841 339 845
rect 407 841 411 845
rect 471 841 475 845
rect 535 841 539 845
rect 599 841 603 845
rect 655 841 659 845
rect 703 841 707 845
rect 751 841 755 845
rect 799 841 803 845
rect 847 841 851 845
rect 903 841 907 845
rect 967 841 971 845
rect 1039 841 1043 845
rect 1103 841 1107 845
rect 1167 841 1171 845
rect 1231 841 1235 845
rect 1287 841 1291 845
rect 1343 841 1347 845
rect 1399 841 1403 845
rect 1463 841 1467 845
rect 1663 843 1667 847
rect 111 825 115 829
rect 135 827 139 831
rect 167 827 171 831
rect 215 827 219 831
rect 279 827 283 831
rect 343 827 347 831
rect 415 827 419 831
rect 479 827 483 831
rect 543 827 547 831
rect 607 827 611 831
rect 671 827 675 831
rect 735 827 739 831
rect 791 827 795 831
rect 847 827 851 831
rect 911 827 915 831
rect 975 827 979 831
rect 1039 827 1043 831
rect 1111 827 1115 831
rect 1183 827 1187 831
rect 1247 827 1251 831
rect 1311 827 1315 831
rect 1367 827 1371 831
rect 1423 827 1427 831
rect 1479 827 1483 831
rect 1535 827 1539 831
rect 1591 827 1595 831
rect 1663 825 1667 829
rect 111 808 115 812
rect 135 810 139 814
rect 167 810 171 814
rect 215 810 219 814
rect 279 810 283 814
rect 343 810 347 814
rect 415 810 419 814
rect 479 810 483 814
rect 543 810 547 814
rect 607 810 611 814
rect 671 810 675 814
rect 735 810 739 814
rect 791 810 795 814
rect 847 810 851 814
rect 911 810 915 814
rect 975 810 979 814
rect 1039 810 1043 814
rect 1111 810 1115 814
rect 1183 810 1187 814
rect 1247 810 1251 814
rect 1311 810 1315 814
rect 1367 810 1371 814
rect 1423 810 1427 814
rect 1479 810 1483 814
rect 1535 810 1539 814
rect 1591 810 1595 814
rect 1663 808 1667 812
rect 111 776 115 780
rect 135 774 139 778
rect 175 774 179 778
rect 231 774 235 778
rect 295 774 299 778
rect 367 774 371 778
rect 447 774 451 778
rect 527 774 531 778
rect 615 774 619 778
rect 703 774 707 778
rect 791 774 795 778
rect 871 774 875 778
rect 951 774 955 778
rect 1023 774 1027 778
rect 1095 774 1099 778
rect 1167 774 1171 778
rect 1231 774 1235 778
rect 1295 774 1299 778
rect 1359 774 1363 778
rect 1415 774 1419 778
rect 1471 774 1475 778
rect 1527 774 1531 778
rect 1591 774 1595 778
rect 1663 776 1667 780
rect 111 759 115 763
rect 135 757 139 761
rect 175 757 179 761
rect 231 757 235 761
rect 295 757 299 761
rect 367 757 371 761
rect 447 757 451 761
rect 527 757 531 761
rect 615 757 619 761
rect 703 757 707 761
rect 791 757 795 761
rect 871 757 875 761
rect 951 757 955 761
rect 1023 757 1027 761
rect 1095 757 1099 761
rect 1167 757 1171 761
rect 1231 757 1235 761
rect 1295 757 1299 761
rect 1359 757 1363 761
rect 1415 757 1419 761
rect 1471 757 1475 761
rect 1527 757 1531 761
rect 1591 757 1595 761
rect 1663 759 1667 763
rect 111 741 115 745
rect 215 743 219 747
rect 247 743 251 747
rect 279 743 283 747
rect 319 743 323 747
rect 359 743 363 747
rect 399 743 403 747
rect 439 743 443 747
rect 487 743 491 747
rect 543 743 547 747
rect 607 743 611 747
rect 671 743 675 747
rect 735 743 739 747
rect 799 743 803 747
rect 863 743 867 747
rect 927 743 931 747
rect 991 743 995 747
rect 1055 743 1059 747
rect 1119 743 1123 747
rect 1183 743 1187 747
rect 1239 743 1243 747
rect 1295 743 1299 747
rect 1351 743 1355 747
rect 1407 743 1411 747
rect 1463 743 1467 747
rect 1519 743 1523 747
rect 1583 743 1587 747
rect 1623 743 1627 747
rect 1663 741 1667 745
rect 111 724 115 728
rect 215 726 219 730
rect 247 726 251 730
rect 279 726 283 730
rect 319 726 323 730
rect 359 726 363 730
rect 399 726 403 730
rect 439 726 443 730
rect 487 726 491 730
rect 543 726 547 730
rect 607 726 611 730
rect 671 726 675 730
rect 735 726 739 730
rect 799 726 803 730
rect 863 726 867 730
rect 927 726 931 730
rect 991 726 995 730
rect 1055 726 1059 730
rect 1119 726 1123 730
rect 1183 726 1187 730
rect 1239 726 1243 730
rect 1295 726 1299 730
rect 1351 726 1355 730
rect 1407 726 1411 730
rect 1463 726 1467 730
rect 1519 726 1523 730
rect 1583 726 1587 730
rect 1623 726 1627 730
rect 1663 724 1667 728
rect 111 692 115 696
rect 279 690 283 694
rect 311 690 315 694
rect 343 690 347 694
rect 375 690 379 694
rect 407 690 411 694
rect 439 690 443 694
rect 471 690 475 694
rect 503 690 507 694
rect 543 690 547 694
rect 591 690 595 694
rect 647 690 651 694
rect 703 690 707 694
rect 759 690 763 694
rect 823 690 827 694
rect 887 690 891 694
rect 959 690 963 694
rect 1023 690 1027 694
rect 1087 690 1091 694
rect 1159 690 1163 694
rect 1223 690 1227 694
rect 1287 690 1291 694
rect 1351 690 1355 694
rect 1415 690 1419 694
rect 1471 690 1475 694
rect 1527 690 1531 694
rect 1583 690 1587 694
rect 1623 690 1627 694
rect 1663 692 1667 696
rect 111 675 115 679
rect 279 673 283 677
rect 311 673 315 677
rect 343 673 347 677
rect 375 673 379 677
rect 407 673 411 677
rect 439 673 443 677
rect 471 673 475 677
rect 503 673 507 677
rect 543 673 547 677
rect 591 673 595 677
rect 647 673 651 677
rect 703 673 707 677
rect 759 673 763 677
rect 823 673 827 677
rect 887 673 891 677
rect 959 673 963 677
rect 1023 673 1027 677
rect 1087 673 1091 677
rect 1159 673 1163 677
rect 1223 673 1227 677
rect 1287 673 1291 677
rect 1351 673 1355 677
rect 1415 673 1419 677
rect 1471 673 1475 677
rect 1527 673 1531 677
rect 1583 673 1587 677
rect 1623 673 1627 677
rect 1663 675 1667 679
rect 111 657 115 661
rect 295 659 299 663
rect 327 659 331 663
rect 359 659 363 663
rect 391 659 395 663
rect 423 659 427 663
rect 455 659 459 663
rect 487 659 491 663
rect 519 659 523 663
rect 551 659 555 663
rect 591 659 595 663
rect 639 659 643 663
rect 687 659 691 663
rect 735 659 739 663
rect 791 659 795 663
rect 847 659 851 663
rect 911 659 915 663
rect 975 659 979 663
rect 1047 659 1051 663
rect 1127 659 1131 663
rect 1215 659 1219 663
rect 1295 659 1299 663
rect 1383 659 1387 663
rect 1471 659 1475 663
rect 1559 659 1563 663
rect 1623 659 1627 663
rect 1663 657 1667 661
rect 111 640 115 644
rect 295 642 299 646
rect 327 642 331 646
rect 359 642 363 646
rect 391 642 395 646
rect 423 642 427 646
rect 455 642 459 646
rect 487 642 491 646
rect 519 642 523 646
rect 551 642 555 646
rect 591 642 595 646
rect 639 642 643 646
rect 687 642 691 646
rect 735 642 739 646
rect 791 642 795 646
rect 847 642 851 646
rect 911 642 915 646
rect 975 642 979 646
rect 1047 642 1051 646
rect 1127 642 1131 646
rect 1215 642 1219 646
rect 1295 642 1299 646
rect 1383 642 1387 646
rect 1471 642 1475 646
rect 1559 642 1563 646
rect 1623 642 1627 646
rect 1663 640 1667 644
rect 111 612 115 616
rect 247 610 251 614
rect 279 610 283 614
rect 319 610 323 614
rect 367 610 371 614
rect 423 610 427 614
rect 471 610 475 614
rect 519 610 523 614
rect 567 610 571 614
rect 615 610 619 614
rect 663 610 667 614
rect 719 610 723 614
rect 775 610 779 614
rect 831 610 835 614
rect 895 610 899 614
rect 967 610 971 614
rect 1047 610 1051 614
rect 1127 610 1131 614
rect 1207 610 1211 614
rect 1287 610 1291 614
rect 1359 610 1363 614
rect 1431 610 1435 614
rect 1503 610 1507 614
rect 1575 610 1579 614
rect 1623 610 1627 614
rect 1663 612 1667 616
rect 111 595 115 599
rect 247 593 251 597
rect 279 593 283 597
rect 319 593 323 597
rect 367 593 371 597
rect 423 593 427 597
rect 471 593 475 597
rect 519 593 523 597
rect 567 593 571 597
rect 615 593 619 597
rect 663 593 667 597
rect 719 593 723 597
rect 775 593 779 597
rect 831 593 835 597
rect 895 593 899 597
rect 967 593 971 597
rect 1047 593 1051 597
rect 1127 593 1131 597
rect 1207 593 1211 597
rect 1287 593 1291 597
rect 1359 593 1363 597
rect 1431 593 1435 597
rect 1503 593 1507 597
rect 1575 593 1579 597
rect 1623 593 1627 597
rect 1663 595 1667 599
rect 111 577 115 581
rect 167 579 171 583
rect 215 579 219 583
rect 271 579 275 583
rect 335 579 339 583
rect 407 579 411 583
rect 487 579 491 583
rect 559 579 563 583
rect 631 579 635 583
rect 703 579 707 583
rect 767 579 771 583
rect 823 579 827 583
rect 879 579 883 583
rect 935 579 939 583
rect 991 579 995 583
rect 1047 579 1051 583
rect 1103 579 1107 583
rect 1159 579 1163 583
rect 1215 579 1219 583
rect 1271 579 1275 583
rect 1327 579 1331 583
rect 1383 579 1387 583
rect 1447 579 1451 583
rect 1511 579 1515 583
rect 1575 579 1579 583
rect 1623 579 1627 583
rect 1663 577 1667 581
rect 111 560 115 564
rect 167 562 171 566
rect 215 562 219 566
rect 271 562 275 566
rect 335 562 339 566
rect 407 562 411 566
rect 487 562 491 566
rect 559 562 563 566
rect 631 562 635 566
rect 703 562 707 566
rect 767 562 771 566
rect 823 562 827 566
rect 879 562 883 566
rect 935 562 939 566
rect 991 562 995 566
rect 1047 562 1051 566
rect 1103 562 1107 566
rect 1159 562 1163 566
rect 1215 562 1219 566
rect 1271 562 1275 566
rect 1327 562 1331 566
rect 1383 562 1387 566
rect 1447 562 1451 566
rect 1511 562 1515 566
rect 1575 562 1579 566
rect 1623 562 1627 566
rect 1663 560 1667 564
rect 111 528 115 532
rect 135 526 139 530
rect 167 526 171 530
rect 199 526 203 530
rect 231 526 235 530
rect 279 526 283 530
rect 327 526 331 530
rect 375 526 379 530
rect 431 526 435 530
rect 495 526 499 530
rect 559 526 563 530
rect 623 526 627 530
rect 687 526 691 530
rect 751 526 755 530
rect 815 526 819 530
rect 879 526 883 530
rect 943 526 947 530
rect 1007 526 1011 530
rect 1071 526 1075 530
rect 1127 526 1131 530
rect 1183 526 1187 530
rect 1231 526 1235 530
rect 1279 526 1283 530
rect 1335 526 1339 530
rect 1391 526 1395 530
rect 1447 526 1451 530
rect 1511 526 1515 530
rect 1575 526 1579 530
rect 1623 526 1627 530
rect 1663 528 1667 532
rect 111 511 115 515
rect 135 509 139 513
rect 167 509 171 513
rect 199 509 203 513
rect 231 509 235 513
rect 279 509 283 513
rect 327 509 331 513
rect 375 509 379 513
rect 431 509 435 513
rect 495 509 499 513
rect 559 509 563 513
rect 623 509 627 513
rect 687 509 691 513
rect 751 509 755 513
rect 815 509 819 513
rect 879 509 883 513
rect 943 509 947 513
rect 1007 509 1011 513
rect 1071 509 1075 513
rect 1127 509 1131 513
rect 1183 509 1187 513
rect 1231 509 1235 513
rect 1279 509 1283 513
rect 1335 509 1339 513
rect 1391 509 1395 513
rect 1447 509 1451 513
rect 1511 509 1515 513
rect 1575 509 1579 513
rect 1623 509 1627 513
rect 1663 511 1667 515
rect 111 493 115 497
rect 135 495 139 499
rect 167 495 171 499
rect 199 495 203 499
rect 239 495 243 499
rect 287 495 291 499
rect 327 495 331 499
rect 375 495 379 499
rect 423 495 427 499
rect 479 495 483 499
rect 543 495 547 499
rect 615 495 619 499
rect 695 495 699 499
rect 775 495 779 499
rect 847 495 851 499
rect 919 495 923 499
rect 983 495 987 499
rect 1039 495 1043 499
rect 1095 495 1099 499
rect 1143 495 1147 499
rect 1191 495 1195 499
rect 1239 495 1243 499
rect 1287 495 1291 499
rect 1335 495 1339 499
rect 1383 495 1387 499
rect 1431 495 1435 499
rect 1479 495 1483 499
rect 1535 495 1539 499
rect 1591 495 1595 499
rect 1623 495 1627 499
rect 1663 493 1667 497
rect 111 476 115 480
rect 135 478 139 482
rect 167 478 171 482
rect 199 478 203 482
rect 239 478 243 482
rect 287 478 291 482
rect 327 478 331 482
rect 375 478 379 482
rect 423 478 427 482
rect 479 478 483 482
rect 543 478 547 482
rect 615 478 619 482
rect 695 478 699 482
rect 775 478 779 482
rect 847 478 851 482
rect 919 478 923 482
rect 983 478 987 482
rect 1039 478 1043 482
rect 1095 478 1099 482
rect 1143 478 1147 482
rect 1191 478 1195 482
rect 1239 478 1243 482
rect 1287 478 1291 482
rect 1335 478 1339 482
rect 1383 478 1387 482
rect 1431 478 1435 482
rect 1479 478 1483 482
rect 1535 478 1539 482
rect 1591 478 1595 482
rect 1623 478 1627 482
rect 1663 476 1667 480
rect 111 448 115 452
rect 151 446 155 450
rect 207 446 211 450
rect 255 446 259 450
rect 311 446 315 450
rect 367 446 371 450
rect 439 446 443 450
rect 519 446 523 450
rect 599 446 603 450
rect 679 446 683 450
rect 759 446 763 450
rect 839 446 843 450
rect 911 446 915 450
rect 983 446 987 450
rect 1055 446 1059 450
rect 1127 446 1131 450
rect 1199 446 1203 450
rect 1263 446 1267 450
rect 1319 446 1323 450
rect 1375 446 1379 450
rect 1431 446 1435 450
rect 1495 446 1499 450
rect 1663 448 1667 452
rect 111 431 115 435
rect 151 429 155 433
rect 207 429 211 433
rect 255 429 259 433
rect 311 429 315 433
rect 367 429 371 433
rect 439 429 443 433
rect 519 429 523 433
rect 599 429 603 433
rect 679 429 683 433
rect 759 429 763 433
rect 839 429 843 433
rect 911 429 915 433
rect 983 429 987 433
rect 1055 429 1059 433
rect 1127 429 1131 433
rect 1199 429 1203 433
rect 1263 429 1267 433
rect 1319 429 1323 433
rect 1375 429 1379 433
rect 1431 429 1435 433
rect 1495 429 1499 433
rect 1663 431 1667 435
rect 111 413 115 417
rect 175 415 179 419
rect 223 415 227 419
rect 271 415 275 419
rect 319 415 323 419
rect 367 415 371 419
rect 415 415 419 419
rect 471 415 475 419
rect 527 415 531 419
rect 591 415 595 419
rect 663 415 667 419
rect 735 415 739 419
rect 807 415 811 419
rect 871 415 875 419
rect 935 415 939 419
rect 991 415 995 419
rect 1039 415 1043 419
rect 1087 415 1091 419
rect 1127 415 1131 419
rect 1167 415 1171 419
rect 1207 415 1211 419
rect 1247 415 1251 419
rect 1287 415 1291 419
rect 1335 415 1339 419
rect 1383 415 1387 419
rect 1663 413 1667 417
rect 111 396 115 400
rect 175 398 179 402
rect 223 398 227 402
rect 271 398 275 402
rect 319 398 323 402
rect 367 398 371 402
rect 415 398 419 402
rect 471 398 475 402
rect 527 398 531 402
rect 591 398 595 402
rect 663 398 667 402
rect 735 398 739 402
rect 807 398 811 402
rect 871 398 875 402
rect 935 398 939 402
rect 991 398 995 402
rect 1039 398 1043 402
rect 1087 398 1091 402
rect 1127 398 1131 402
rect 1167 398 1171 402
rect 1207 398 1211 402
rect 1247 398 1251 402
rect 1287 398 1291 402
rect 1335 398 1339 402
rect 1383 398 1387 402
rect 1663 396 1667 400
rect 111 364 115 368
rect 135 362 139 366
rect 167 362 171 366
rect 199 362 203 366
rect 239 362 243 366
rect 295 362 299 366
rect 351 362 355 366
rect 407 362 411 366
rect 463 362 467 366
rect 519 362 523 366
rect 575 362 579 366
rect 631 362 635 366
rect 687 362 691 366
rect 743 362 747 366
rect 799 362 803 366
rect 855 362 859 366
rect 919 362 923 366
rect 983 362 987 366
rect 1039 362 1043 366
rect 1095 362 1099 366
rect 1151 362 1155 366
rect 1207 362 1211 366
rect 1255 362 1259 366
rect 1303 362 1307 366
rect 1351 362 1355 366
rect 1399 362 1403 366
rect 1447 362 1451 366
rect 1495 362 1499 366
rect 1543 362 1547 366
rect 1591 362 1595 366
rect 1623 362 1627 366
rect 1663 364 1667 368
rect 111 347 115 351
rect 135 345 139 349
rect 167 345 171 349
rect 199 345 203 349
rect 239 345 243 349
rect 295 345 299 349
rect 351 345 355 349
rect 407 345 411 349
rect 463 345 467 349
rect 519 345 523 349
rect 575 345 579 349
rect 631 345 635 349
rect 687 345 691 349
rect 743 345 747 349
rect 799 345 803 349
rect 855 345 859 349
rect 919 345 923 349
rect 983 345 987 349
rect 1039 345 1043 349
rect 1095 345 1099 349
rect 1151 345 1155 349
rect 1207 345 1211 349
rect 1255 345 1259 349
rect 1303 345 1307 349
rect 1351 345 1355 349
rect 1399 345 1403 349
rect 1447 345 1451 349
rect 1495 345 1499 349
rect 1543 345 1547 349
rect 1591 345 1595 349
rect 1623 345 1627 349
rect 1663 347 1667 351
rect 111 329 115 333
rect 135 331 139 335
rect 167 331 171 335
rect 207 331 211 335
rect 263 331 267 335
rect 327 331 331 335
rect 391 331 395 335
rect 455 331 459 335
rect 519 331 523 335
rect 575 331 579 335
rect 631 331 635 335
rect 687 331 691 335
rect 751 331 755 335
rect 815 331 819 335
rect 879 331 883 335
rect 951 331 955 335
rect 1031 331 1035 335
rect 1111 331 1115 335
rect 1191 331 1195 335
rect 1271 331 1275 335
rect 1343 331 1347 335
rect 1407 331 1411 335
rect 1463 331 1467 335
rect 1519 331 1523 335
rect 1583 331 1587 335
rect 1623 331 1627 335
rect 1663 329 1667 333
rect 111 312 115 316
rect 135 314 139 318
rect 167 314 171 318
rect 207 314 211 318
rect 263 314 267 318
rect 327 314 331 318
rect 391 314 395 318
rect 455 314 459 318
rect 519 314 523 318
rect 575 314 579 318
rect 631 314 635 318
rect 687 314 691 318
rect 751 314 755 318
rect 815 314 819 318
rect 879 314 883 318
rect 951 314 955 318
rect 1031 314 1035 318
rect 1111 314 1115 318
rect 1191 314 1195 318
rect 1271 314 1275 318
rect 1343 314 1347 318
rect 1407 314 1411 318
rect 1463 314 1467 318
rect 1519 314 1523 318
rect 1583 314 1587 318
rect 1623 314 1627 318
rect 1663 312 1667 316
rect 111 284 115 288
rect 135 282 139 286
rect 167 282 171 286
rect 231 282 235 286
rect 295 282 299 286
rect 367 282 371 286
rect 439 282 443 286
rect 503 282 507 286
rect 567 282 571 286
rect 631 282 635 286
rect 687 282 691 286
rect 743 282 747 286
rect 807 282 811 286
rect 879 282 883 286
rect 951 282 955 286
rect 1031 282 1035 286
rect 1111 282 1115 286
rect 1191 282 1195 286
rect 1263 282 1267 286
rect 1327 282 1331 286
rect 1391 282 1395 286
rect 1447 282 1451 286
rect 1495 282 1499 286
rect 1543 282 1547 286
rect 1591 282 1595 286
rect 1623 282 1627 286
rect 1663 284 1667 288
rect 111 267 115 271
rect 135 265 139 269
rect 167 265 171 269
rect 231 265 235 269
rect 295 265 299 269
rect 367 265 371 269
rect 439 265 443 269
rect 503 265 507 269
rect 567 265 571 269
rect 631 265 635 269
rect 687 265 691 269
rect 743 265 747 269
rect 807 265 811 269
rect 879 265 883 269
rect 951 265 955 269
rect 1031 265 1035 269
rect 1111 265 1115 269
rect 1191 265 1195 269
rect 1263 265 1267 269
rect 1327 265 1331 269
rect 1391 265 1395 269
rect 1447 265 1451 269
rect 1495 265 1499 269
rect 1543 265 1547 269
rect 1591 265 1595 269
rect 1623 265 1627 269
rect 1663 267 1667 271
rect 111 245 115 249
rect 135 247 139 251
rect 175 247 179 251
rect 247 247 251 251
rect 319 247 323 251
rect 383 247 387 251
rect 447 247 451 251
rect 519 247 523 251
rect 591 247 595 251
rect 663 247 667 251
rect 743 247 747 251
rect 823 247 827 251
rect 895 247 899 251
rect 967 247 971 251
rect 1031 247 1035 251
rect 1087 247 1091 251
rect 1143 247 1147 251
rect 1199 247 1203 251
rect 1255 247 1259 251
rect 1311 247 1315 251
rect 1367 247 1371 251
rect 1415 247 1419 251
rect 1463 247 1467 251
rect 1519 247 1523 251
rect 1575 247 1579 251
rect 1623 247 1627 251
rect 1663 245 1667 249
rect 111 228 115 232
rect 135 230 139 234
rect 175 230 179 234
rect 247 230 251 234
rect 319 230 323 234
rect 383 230 387 234
rect 447 230 451 234
rect 519 230 523 234
rect 591 230 595 234
rect 663 230 667 234
rect 743 230 747 234
rect 823 230 827 234
rect 895 230 899 234
rect 967 230 971 234
rect 1031 230 1035 234
rect 1087 230 1091 234
rect 1143 230 1147 234
rect 1199 230 1203 234
rect 1255 230 1259 234
rect 1311 230 1315 234
rect 1367 230 1371 234
rect 1415 230 1419 234
rect 1463 230 1467 234
rect 1519 230 1523 234
rect 1575 230 1579 234
rect 1623 230 1627 234
rect 1663 228 1667 232
rect 111 200 115 204
rect 135 198 139 202
rect 167 198 171 202
rect 207 198 211 202
rect 255 198 259 202
rect 303 198 307 202
rect 343 198 347 202
rect 375 198 379 202
rect 415 198 419 202
rect 471 198 475 202
rect 535 198 539 202
rect 615 198 619 202
rect 695 198 699 202
rect 775 198 779 202
rect 855 198 859 202
rect 927 198 931 202
rect 999 198 1003 202
rect 1071 198 1075 202
rect 1143 198 1147 202
rect 1215 198 1219 202
rect 1287 198 1291 202
rect 1351 198 1355 202
rect 1415 198 1419 202
rect 1471 198 1475 202
rect 1527 198 1531 202
rect 1583 198 1587 202
rect 1623 198 1627 202
rect 1663 200 1667 204
rect 111 183 115 187
rect 135 181 139 185
rect 167 181 171 185
rect 207 181 211 185
rect 255 181 259 185
rect 303 181 307 185
rect 343 181 347 185
rect 375 181 379 185
rect 415 181 419 185
rect 471 181 475 185
rect 535 181 539 185
rect 615 181 619 185
rect 695 181 699 185
rect 775 181 779 185
rect 855 181 859 185
rect 927 181 931 185
rect 999 181 1003 185
rect 1071 181 1075 185
rect 1143 181 1147 185
rect 1215 181 1219 185
rect 1287 181 1291 185
rect 1351 181 1355 185
rect 1415 181 1419 185
rect 1471 181 1475 185
rect 1527 181 1531 185
rect 1583 181 1587 185
rect 1623 181 1627 185
rect 1663 183 1667 187
rect 111 165 115 169
rect 135 167 139 171
rect 175 167 179 171
rect 231 167 235 171
rect 287 167 291 171
rect 343 167 347 171
rect 399 167 403 171
rect 455 167 459 171
rect 511 167 515 171
rect 575 167 579 171
rect 639 167 643 171
rect 703 167 707 171
rect 767 167 771 171
rect 831 167 835 171
rect 895 167 899 171
rect 951 167 955 171
rect 1015 167 1019 171
rect 1079 167 1083 171
rect 1143 167 1147 171
rect 1207 167 1211 171
rect 1279 167 1283 171
rect 1351 167 1355 171
rect 1423 167 1427 171
rect 1495 167 1499 171
rect 1567 167 1571 171
rect 1623 167 1627 171
rect 1663 165 1667 169
rect 111 148 115 152
rect 135 150 139 154
rect 175 150 179 154
rect 231 150 235 154
rect 287 150 291 154
rect 343 150 347 154
rect 399 150 403 154
rect 455 150 459 154
rect 511 150 515 154
rect 575 150 579 154
rect 639 150 643 154
rect 703 150 707 154
rect 767 150 771 154
rect 831 150 835 154
rect 895 150 899 154
rect 951 150 955 154
rect 1015 150 1019 154
rect 1079 150 1083 154
rect 1143 150 1147 154
rect 1207 150 1211 154
rect 1279 150 1283 154
rect 1351 150 1355 154
rect 1423 150 1427 154
rect 1495 150 1499 154
rect 1567 150 1571 154
rect 1623 150 1627 154
rect 1663 148 1667 152
rect 111 104 115 108
rect 135 102 139 106
rect 167 102 171 106
rect 199 102 203 106
rect 231 102 235 106
rect 263 102 267 106
rect 295 102 299 106
rect 327 102 331 106
rect 359 102 363 106
rect 391 102 395 106
rect 423 102 427 106
rect 463 102 467 106
rect 503 102 507 106
rect 543 102 547 106
rect 575 102 579 106
rect 607 102 611 106
rect 639 102 643 106
rect 671 102 675 106
rect 703 102 707 106
rect 735 102 739 106
rect 767 102 771 106
rect 799 102 803 106
rect 831 102 835 106
rect 863 102 867 106
rect 895 102 899 106
rect 935 102 939 106
rect 975 102 979 106
rect 1015 102 1019 106
rect 1063 102 1067 106
rect 1103 102 1107 106
rect 1143 102 1147 106
rect 1183 102 1187 106
rect 1223 102 1227 106
rect 1263 102 1267 106
rect 1295 102 1299 106
rect 1335 102 1339 106
rect 1375 102 1379 106
rect 1415 102 1419 106
rect 1455 102 1459 106
rect 1503 102 1507 106
rect 1551 102 1555 106
rect 1591 102 1595 106
rect 1623 102 1627 106
rect 1663 104 1667 108
rect 111 87 115 91
rect 135 85 139 89
rect 167 85 171 89
rect 199 85 203 89
rect 231 85 235 89
rect 263 85 267 89
rect 295 85 299 89
rect 327 85 331 89
rect 359 85 363 89
rect 391 85 395 89
rect 423 85 427 89
rect 463 85 467 89
rect 503 85 507 89
rect 543 85 547 89
rect 575 85 579 89
rect 607 85 611 89
rect 639 85 643 89
rect 671 85 675 89
rect 703 85 707 89
rect 735 85 739 89
rect 767 85 771 89
rect 799 85 803 89
rect 831 85 835 89
rect 863 85 867 89
rect 895 85 899 89
rect 935 85 939 89
rect 975 85 979 89
rect 1015 85 1019 89
rect 1063 85 1067 89
rect 1103 85 1107 89
rect 1143 85 1147 89
rect 1183 85 1187 89
rect 1223 85 1227 89
rect 1263 85 1267 89
rect 1295 85 1299 89
rect 1335 85 1339 89
rect 1375 85 1379 89
rect 1415 85 1419 89
rect 1455 85 1459 89
rect 1503 85 1507 89
rect 1551 85 1555 89
rect 1591 85 1595 89
rect 1623 85 1627 89
rect 1663 87 1667 91
<< m3 >>
rect 111 1718 115 1719
rect 111 1713 115 1714
rect 255 1718 259 1719
rect 255 1713 259 1714
rect 287 1718 291 1719
rect 287 1713 291 1714
rect 319 1718 323 1719
rect 319 1713 323 1714
rect 359 1718 363 1719
rect 359 1713 363 1714
rect 407 1718 411 1719
rect 407 1713 411 1714
rect 455 1718 459 1719
rect 455 1713 459 1714
rect 503 1718 507 1719
rect 503 1713 507 1714
rect 551 1718 555 1719
rect 551 1713 555 1714
rect 607 1718 611 1719
rect 607 1713 611 1714
rect 663 1718 667 1719
rect 663 1713 667 1714
rect 727 1718 731 1719
rect 727 1713 731 1714
rect 783 1718 787 1719
rect 783 1713 787 1714
rect 839 1718 843 1719
rect 839 1713 843 1714
rect 895 1718 899 1719
rect 895 1713 899 1714
rect 951 1718 955 1719
rect 951 1713 955 1714
rect 1007 1718 1011 1719
rect 1007 1713 1011 1714
rect 1063 1718 1067 1719
rect 1063 1713 1067 1714
rect 1119 1718 1123 1719
rect 1119 1713 1123 1714
rect 1175 1718 1179 1719
rect 1175 1713 1179 1714
rect 1231 1718 1235 1719
rect 1231 1713 1235 1714
rect 1287 1718 1291 1719
rect 1287 1713 1291 1714
rect 1335 1718 1339 1719
rect 1335 1713 1339 1714
rect 1375 1718 1379 1719
rect 1375 1713 1379 1714
rect 1423 1718 1427 1719
rect 1423 1713 1427 1714
rect 1471 1718 1475 1719
rect 1471 1713 1475 1714
rect 1519 1718 1523 1719
rect 1519 1713 1523 1714
rect 1663 1718 1667 1719
rect 1663 1713 1667 1714
rect 112 1705 114 1713
rect 110 1704 116 1705
rect 110 1700 111 1704
rect 115 1700 116 1704
rect 256 1703 258 1713
rect 288 1703 290 1713
rect 320 1703 322 1713
rect 360 1703 362 1713
rect 408 1703 410 1713
rect 456 1703 458 1713
rect 504 1703 506 1713
rect 552 1703 554 1713
rect 608 1703 610 1713
rect 664 1703 666 1713
rect 728 1703 730 1713
rect 784 1703 786 1713
rect 840 1703 842 1713
rect 896 1703 898 1713
rect 952 1703 954 1713
rect 1008 1703 1010 1713
rect 1064 1703 1066 1713
rect 1120 1703 1122 1713
rect 1176 1703 1178 1713
rect 1232 1703 1234 1713
rect 1288 1703 1290 1713
rect 1336 1703 1338 1713
rect 1376 1703 1378 1713
rect 1424 1703 1426 1713
rect 1472 1703 1474 1713
rect 1520 1703 1522 1713
rect 1664 1705 1666 1713
rect 1662 1704 1668 1705
rect 110 1699 116 1700
rect 254 1702 260 1703
rect 254 1698 255 1702
rect 259 1698 260 1702
rect 254 1697 260 1698
rect 286 1702 292 1703
rect 286 1698 287 1702
rect 291 1698 292 1702
rect 286 1697 292 1698
rect 318 1702 324 1703
rect 318 1698 319 1702
rect 323 1698 324 1702
rect 318 1697 324 1698
rect 358 1702 364 1703
rect 358 1698 359 1702
rect 363 1698 364 1702
rect 358 1697 364 1698
rect 406 1702 412 1703
rect 406 1698 407 1702
rect 411 1698 412 1702
rect 406 1697 412 1698
rect 454 1702 460 1703
rect 454 1698 455 1702
rect 459 1698 460 1702
rect 454 1697 460 1698
rect 502 1702 508 1703
rect 502 1698 503 1702
rect 507 1698 508 1702
rect 502 1697 508 1698
rect 550 1702 556 1703
rect 550 1698 551 1702
rect 555 1698 556 1702
rect 550 1697 556 1698
rect 606 1702 612 1703
rect 606 1698 607 1702
rect 611 1698 612 1702
rect 606 1697 612 1698
rect 662 1702 668 1703
rect 662 1698 663 1702
rect 667 1698 668 1702
rect 662 1697 668 1698
rect 726 1702 732 1703
rect 726 1698 727 1702
rect 731 1698 732 1702
rect 726 1697 732 1698
rect 782 1702 788 1703
rect 782 1698 783 1702
rect 787 1698 788 1702
rect 782 1697 788 1698
rect 838 1702 844 1703
rect 838 1698 839 1702
rect 843 1698 844 1702
rect 838 1697 844 1698
rect 894 1702 900 1703
rect 894 1698 895 1702
rect 899 1698 900 1702
rect 894 1697 900 1698
rect 950 1702 956 1703
rect 950 1698 951 1702
rect 955 1698 956 1702
rect 950 1697 956 1698
rect 1006 1702 1012 1703
rect 1006 1698 1007 1702
rect 1011 1698 1012 1702
rect 1006 1697 1012 1698
rect 1062 1702 1068 1703
rect 1062 1698 1063 1702
rect 1067 1698 1068 1702
rect 1062 1697 1068 1698
rect 1118 1702 1124 1703
rect 1118 1698 1119 1702
rect 1123 1698 1124 1702
rect 1118 1697 1124 1698
rect 1174 1702 1180 1703
rect 1174 1698 1175 1702
rect 1179 1698 1180 1702
rect 1174 1697 1180 1698
rect 1230 1702 1236 1703
rect 1230 1698 1231 1702
rect 1235 1698 1236 1702
rect 1230 1697 1236 1698
rect 1286 1702 1292 1703
rect 1286 1698 1287 1702
rect 1291 1698 1292 1702
rect 1286 1697 1292 1698
rect 1334 1702 1340 1703
rect 1334 1698 1335 1702
rect 1339 1698 1340 1702
rect 1334 1697 1340 1698
rect 1374 1702 1380 1703
rect 1374 1698 1375 1702
rect 1379 1698 1380 1702
rect 1374 1697 1380 1698
rect 1422 1702 1428 1703
rect 1422 1698 1423 1702
rect 1427 1698 1428 1702
rect 1422 1697 1428 1698
rect 1470 1702 1476 1703
rect 1470 1698 1471 1702
rect 1475 1698 1476 1702
rect 1470 1697 1476 1698
rect 1518 1702 1524 1703
rect 1518 1698 1519 1702
rect 1523 1698 1524 1702
rect 1662 1700 1663 1704
rect 1667 1700 1668 1704
rect 1662 1699 1668 1700
rect 1518 1697 1524 1698
rect 110 1687 116 1688
rect 110 1683 111 1687
rect 115 1683 116 1687
rect 1662 1687 1668 1688
rect 110 1682 116 1683
rect 254 1685 260 1686
rect 112 1679 114 1682
rect 254 1681 255 1685
rect 259 1681 260 1685
rect 254 1680 260 1681
rect 286 1685 292 1686
rect 286 1681 287 1685
rect 291 1681 292 1685
rect 286 1680 292 1681
rect 318 1685 324 1686
rect 318 1681 319 1685
rect 323 1681 324 1685
rect 318 1680 324 1681
rect 358 1685 364 1686
rect 358 1681 359 1685
rect 363 1681 364 1685
rect 358 1680 364 1681
rect 406 1685 412 1686
rect 406 1681 407 1685
rect 411 1681 412 1685
rect 406 1680 412 1681
rect 454 1685 460 1686
rect 454 1681 455 1685
rect 459 1681 460 1685
rect 454 1680 460 1681
rect 502 1685 508 1686
rect 502 1681 503 1685
rect 507 1681 508 1685
rect 502 1680 508 1681
rect 550 1685 556 1686
rect 550 1681 551 1685
rect 555 1681 556 1685
rect 550 1680 556 1681
rect 606 1685 612 1686
rect 606 1681 607 1685
rect 611 1681 612 1685
rect 606 1680 612 1681
rect 662 1685 668 1686
rect 662 1681 663 1685
rect 667 1681 668 1685
rect 662 1680 668 1681
rect 726 1685 732 1686
rect 726 1681 727 1685
rect 731 1681 732 1685
rect 726 1680 732 1681
rect 782 1685 788 1686
rect 782 1681 783 1685
rect 787 1681 788 1685
rect 782 1680 788 1681
rect 838 1685 844 1686
rect 838 1681 839 1685
rect 843 1681 844 1685
rect 838 1680 844 1681
rect 894 1685 900 1686
rect 894 1681 895 1685
rect 899 1681 900 1685
rect 894 1680 900 1681
rect 950 1685 956 1686
rect 950 1681 951 1685
rect 955 1681 956 1685
rect 950 1680 956 1681
rect 1006 1685 1012 1686
rect 1006 1681 1007 1685
rect 1011 1681 1012 1685
rect 1006 1680 1012 1681
rect 1062 1685 1068 1686
rect 1062 1681 1063 1685
rect 1067 1681 1068 1685
rect 1062 1680 1068 1681
rect 1118 1685 1124 1686
rect 1118 1681 1119 1685
rect 1123 1681 1124 1685
rect 1118 1680 1124 1681
rect 1174 1685 1180 1686
rect 1174 1681 1175 1685
rect 1179 1681 1180 1685
rect 1174 1680 1180 1681
rect 1230 1685 1236 1686
rect 1230 1681 1231 1685
rect 1235 1681 1236 1685
rect 1230 1680 1236 1681
rect 1286 1685 1292 1686
rect 1286 1681 1287 1685
rect 1291 1681 1292 1685
rect 1286 1680 1292 1681
rect 1334 1685 1340 1686
rect 1334 1681 1335 1685
rect 1339 1681 1340 1685
rect 1334 1680 1340 1681
rect 1374 1685 1380 1686
rect 1374 1681 1375 1685
rect 1379 1681 1380 1685
rect 1374 1680 1380 1681
rect 1422 1685 1428 1686
rect 1422 1681 1423 1685
rect 1427 1681 1428 1685
rect 1422 1680 1428 1681
rect 1470 1685 1476 1686
rect 1470 1681 1471 1685
rect 1475 1681 1476 1685
rect 1470 1680 1476 1681
rect 1518 1685 1524 1686
rect 1518 1681 1519 1685
rect 1523 1681 1524 1685
rect 1662 1683 1663 1687
rect 1667 1683 1668 1687
rect 1662 1682 1668 1683
rect 1518 1680 1524 1681
rect 111 1678 115 1679
rect 111 1673 115 1674
rect 135 1678 139 1679
rect 112 1670 114 1673
rect 135 1672 139 1674
rect 167 1678 171 1679
rect 167 1672 171 1674
rect 215 1678 219 1679
rect 215 1672 219 1674
rect 255 1678 259 1680
rect 255 1673 259 1674
rect 279 1678 283 1679
rect 279 1672 283 1674
rect 287 1678 291 1680
rect 287 1673 291 1674
rect 319 1678 323 1680
rect 319 1673 323 1674
rect 343 1678 347 1679
rect 343 1672 347 1674
rect 359 1678 363 1680
rect 359 1673 363 1674
rect 407 1678 411 1680
rect 407 1673 411 1674
rect 415 1678 419 1679
rect 415 1672 419 1674
rect 455 1678 459 1680
rect 455 1673 459 1674
rect 487 1678 491 1679
rect 487 1672 491 1674
rect 503 1678 507 1680
rect 503 1673 507 1674
rect 551 1678 555 1680
rect 551 1673 555 1674
rect 559 1678 563 1679
rect 559 1672 563 1674
rect 607 1678 611 1680
rect 607 1673 611 1674
rect 631 1678 635 1679
rect 631 1672 635 1674
rect 663 1678 667 1680
rect 663 1673 667 1674
rect 711 1678 715 1679
rect 711 1672 715 1674
rect 727 1678 731 1680
rect 727 1673 731 1674
rect 783 1678 787 1680
rect 783 1673 787 1674
rect 791 1678 795 1679
rect 791 1672 795 1674
rect 839 1678 843 1680
rect 839 1673 843 1674
rect 871 1678 875 1679
rect 871 1672 875 1674
rect 895 1678 899 1680
rect 895 1673 899 1674
rect 951 1678 955 1680
rect 951 1672 955 1674
rect 1007 1678 1011 1680
rect 1007 1673 1011 1674
rect 1031 1678 1035 1679
rect 1031 1672 1035 1674
rect 1063 1678 1067 1680
rect 1063 1673 1067 1674
rect 1103 1678 1107 1679
rect 1103 1672 1107 1674
rect 1119 1678 1123 1680
rect 1119 1673 1123 1674
rect 1175 1678 1179 1680
rect 1175 1672 1179 1674
rect 1231 1678 1235 1680
rect 1231 1673 1235 1674
rect 1247 1678 1251 1679
rect 1247 1672 1251 1674
rect 1287 1678 1291 1680
rect 1287 1673 1291 1674
rect 1319 1678 1323 1679
rect 1319 1672 1323 1674
rect 1335 1678 1339 1680
rect 1335 1673 1339 1674
rect 1375 1678 1379 1680
rect 1375 1673 1379 1674
rect 1391 1678 1395 1679
rect 1391 1672 1395 1674
rect 1423 1678 1427 1680
rect 1423 1673 1427 1674
rect 1455 1678 1459 1679
rect 1455 1672 1459 1674
rect 1471 1678 1475 1680
rect 1471 1673 1475 1674
rect 1519 1678 1523 1680
rect 1664 1679 1666 1682
rect 1519 1672 1523 1674
rect 1583 1678 1587 1679
rect 1583 1672 1587 1674
rect 1623 1678 1627 1679
rect 1623 1672 1627 1674
rect 1663 1678 1667 1679
rect 1663 1673 1667 1674
rect 134 1671 140 1672
rect 110 1669 116 1670
rect 110 1665 111 1669
rect 115 1665 116 1669
rect 134 1667 135 1671
rect 139 1667 140 1671
rect 134 1666 140 1667
rect 166 1671 172 1672
rect 166 1667 167 1671
rect 171 1667 172 1671
rect 166 1666 172 1667
rect 214 1671 220 1672
rect 214 1667 215 1671
rect 219 1667 220 1671
rect 214 1666 220 1667
rect 278 1671 284 1672
rect 278 1667 279 1671
rect 283 1667 284 1671
rect 278 1666 284 1667
rect 342 1671 348 1672
rect 342 1667 343 1671
rect 347 1667 348 1671
rect 342 1666 348 1667
rect 414 1671 420 1672
rect 414 1667 415 1671
rect 419 1667 420 1671
rect 414 1666 420 1667
rect 486 1671 492 1672
rect 486 1667 487 1671
rect 491 1667 492 1671
rect 486 1666 492 1667
rect 558 1671 564 1672
rect 558 1667 559 1671
rect 563 1667 564 1671
rect 558 1666 564 1667
rect 630 1671 636 1672
rect 630 1667 631 1671
rect 635 1667 636 1671
rect 630 1666 636 1667
rect 710 1671 716 1672
rect 710 1667 711 1671
rect 715 1667 716 1671
rect 710 1666 716 1667
rect 790 1671 796 1672
rect 790 1667 791 1671
rect 795 1667 796 1671
rect 790 1666 796 1667
rect 870 1671 876 1672
rect 870 1667 871 1671
rect 875 1667 876 1671
rect 870 1666 876 1667
rect 950 1671 956 1672
rect 950 1667 951 1671
rect 955 1667 956 1671
rect 950 1666 956 1667
rect 1030 1671 1036 1672
rect 1030 1667 1031 1671
rect 1035 1667 1036 1671
rect 1030 1666 1036 1667
rect 1102 1671 1108 1672
rect 1102 1667 1103 1671
rect 1107 1667 1108 1671
rect 1102 1666 1108 1667
rect 1174 1671 1180 1672
rect 1174 1667 1175 1671
rect 1179 1667 1180 1671
rect 1174 1666 1180 1667
rect 1246 1671 1252 1672
rect 1246 1667 1247 1671
rect 1251 1667 1252 1671
rect 1246 1666 1252 1667
rect 1318 1671 1324 1672
rect 1318 1667 1319 1671
rect 1323 1667 1324 1671
rect 1318 1666 1324 1667
rect 1390 1671 1396 1672
rect 1390 1667 1391 1671
rect 1395 1667 1396 1671
rect 1390 1666 1396 1667
rect 1454 1671 1460 1672
rect 1454 1667 1455 1671
rect 1459 1667 1460 1671
rect 1454 1666 1460 1667
rect 1518 1671 1524 1672
rect 1518 1667 1519 1671
rect 1523 1667 1524 1671
rect 1518 1666 1524 1667
rect 1582 1671 1588 1672
rect 1582 1667 1583 1671
rect 1587 1667 1588 1671
rect 1582 1666 1588 1667
rect 1622 1671 1628 1672
rect 1622 1667 1623 1671
rect 1627 1667 1628 1671
rect 1664 1670 1666 1673
rect 1622 1666 1628 1667
rect 1662 1669 1668 1670
rect 110 1664 116 1665
rect 1662 1665 1663 1669
rect 1667 1665 1668 1669
rect 1662 1664 1668 1665
rect 134 1654 140 1655
rect 110 1652 116 1653
rect 110 1648 111 1652
rect 115 1648 116 1652
rect 134 1650 135 1654
rect 139 1650 140 1654
rect 134 1649 140 1650
rect 166 1654 172 1655
rect 166 1650 167 1654
rect 171 1650 172 1654
rect 166 1649 172 1650
rect 214 1654 220 1655
rect 214 1650 215 1654
rect 219 1650 220 1654
rect 214 1649 220 1650
rect 278 1654 284 1655
rect 278 1650 279 1654
rect 283 1650 284 1654
rect 278 1649 284 1650
rect 342 1654 348 1655
rect 342 1650 343 1654
rect 347 1650 348 1654
rect 342 1649 348 1650
rect 414 1654 420 1655
rect 414 1650 415 1654
rect 419 1650 420 1654
rect 414 1649 420 1650
rect 486 1654 492 1655
rect 486 1650 487 1654
rect 491 1650 492 1654
rect 486 1649 492 1650
rect 558 1654 564 1655
rect 558 1650 559 1654
rect 563 1650 564 1654
rect 558 1649 564 1650
rect 630 1654 636 1655
rect 630 1650 631 1654
rect 635 1650 636 1654
rect 630 1649 636 1650
rect 710 1654 716 1655
rect 710 1650 711 1654
rect 715 1650 716 1654
rect 710 1649 716 1650
rect 790 1654 796 1655
rect 790 1650 791 1654
rect 795 1650 796 1654
rect 790 1649 796 1650
rect 870 1654 876 1655
rect 870 1650 871 1654
rect 875 1650 876 1654
rect 870 1649 876 1650
rect 950 1654 956 1655
rect 950 1650 951 1654
rect 955 1650 956 1654
rect 950 1649 956 1650
rect 1030 1654 1036 1655
rect 1030 1650 1031 1654
rect 1035 1650 1036 1654
rect 1030 1649 1036 1650
rect 1102 1654 1108 1655
rect 1102 1650 1103 1654
rect 1107 1650 1108 1654
rect 1102 1649 1108 1650
rect 1174 1654 1180 1655
rect 1174 1650 1175 1654
rect 1179 1650 1180 1654
rect 1174 1649 1180 1650
rect 1246 1654 1252 1655
rect 1246 1650 1247 1654
rect 1251 1650 1252 1654
rect 1246 1649 1252 1650
rect 1318 1654 1324 1655
rect 1318 1650 1319 1654
rect 1323 1650 1324 1654
rect 1318 1649 1324 1650
rect 1390 1654 1396 1655
rect 1390 1650 1391 1654
rect 1395 1650 1396 1654
rect 1390 1649 1396 1650
rect 1454 1654 1460 1655
rect 1454 1650 1455 1654
rect 1459 1650 1460 1654
rect 1454 1649 1460 1650
rect 1518 1654 1524 1655
rect 1518 1650 1519 1654
rect 1523 1650 1524 1654
rect 1518 1649 1524 1650
rect 1582 1654 1588 1655
rect 1582 1650 1583 1654
rect 1587 1650 1588 1654
rect 1582 1649 1588 1650
rect 1622 1654 1628 1655
rect 1622 1650 1623 1654
rect 1627 1650 1628 1654
rect 1622 1649 1628 1650
rect 1662 1652 1668 1653
rect 110 1647 116 1648
rect 112 1639 114 1647
rect 136 1639 138 1649
rect 168 1639 170 1649
rect 216 1639 218 1649
rect 280 1639 282 1649
rect 344 1639 346 1649
rect 416 1639 418 1649
rect 488 1639 490 1649
rect 560 1639 562 1649
rect 632 1639 634 1649
rect 712 1639 714 1649
rect 792 1639 794 1649
rect 872 1639 874 1649
rect 952 1639 954 1649
rect 1032 1639 1034 1649
rect 1104 1639 1106 1649
rect 1176 1639 1178 1649
rect 1248 1639 1250 1649
rect 1320 1639 1322 1649
rect 1392 1639 1394 1649
rect 1456 1639 1458 1649
rect 1520 1639 1522 1649
rect 1584 1639 1586 1649
rect 1624 1639 1626 1649
rect 1662 1648 1663 1652
rect 1667 1648 1668 1652
rect 1662 1647 1668 1648
rect 1664 1639 1666 1647
rect 111 1638 115 1639
rect 111 1633 115 1634
rect 135 1638 139 1639
rect 135 1633 139 1634
rect 167 1638 171 1639
rect 167 1633 171 1634
rect 183 1638 187 1639
rect 183 1633 187 1634
rect 215 1638 219 1639
rect 215 1633 219 1634
rect 247 1638 251 1639
rect 247 1633 251 1634
rect 279 1638 283 1639
rect 279 1633 283 1634
rect 303 1638 307 1639
rect 303 1633 307 1634
rect 343 1638 347 1639
rect 343 1633 347 1634
rect 359 1638 363 1639
rect 359 1633 363 1634
rect 415 1638 419 1639
rect 415 1633 419 1634
rect 471 1638 475 1639
rect 471 1633 475 1634
rect 487 1638 491 1639
rect 487 1633 491 1634
rect 535 1638 539 1639
rect 535 1633 539 1634
rect 559 1638 563 1639
rect 559 1633 563 1634
rect 599 1638 603 1639
rect 599 1633 603 1634
rect 631 1638 635 1639
rect 631 1633 635 1634
rect 663 1638 667 1639
rect 663 1633 667 1634
rect 711 1638 715 1639
rect 711 1633 715 1634
rect 727 1638 731 1639
rect 727 1633 731 1634
rect 791 1638 795 1639
rect 791 1633 795 1634
rect 799 1638 803 1639
rect 799 1633 803 1634
rect 871 1638 875 1639
rect 871 1633 875 1634
rect 943 1638 947 1639
rect 943 1633 947 1634
rect 951 1638 955 1639
rect 951 1633 955 1634
rect 1023 1638 1027 1639
rect 1023 1633 1027 1634
rect 1031 1638 1035 1639
rect 1031 1633 1035 1634
rect 1103 1638 1107 1639
rect 1103 1633 1107 1634
rect 1175 1638 1179 1639
rect 1175 1633 1179 1634
rect 1247 1638 1251 1639
rect 1247 1633 1251 1634
rect 1319 1638 1323 1639
rect 1319 1633 1323 1634
rect 1391 1638 1395 1639
rect 1391 1633 1395 1634
rect 1399 1638 1403 1639
rect 1399 1633 1403 1634
rect 1455 1638 1459 1639
rect 1455 1633 1459 1634
rect 1479 1638 1483 1639
rect 1479 1633 1483 1634
rect 1519 1638 1523 1639
rect 1519 1633 1523 1634
rect 1559 1638 1563 1639
rect 1559 1633 1563 1634
rect 1583 1638 1587 1639
rect 1583 1633 1587 1634
rect 1623 1638 1627 1639
rect 1623 1633 1627 1634
rect 1663 1638 1667 1639
rect 1663 1633 1667 1634
rect 112 1625 114 1633
rect 110 1624 116 1625
rect 110 1620 111 1624
rect 115 1620 116 1624
rect 136 1623 138 1633
rect 184 1623 186 1633
rect 248 1623 250 1633
rect 304 1623 306 1633
rect 360 1623 362 1633
rect 416 1623 418 1633
rect 472 1623 474 1633
rect 536 1623 538 1633
rect 600 1623 602 1633
rect 664 1623 666 1633
rect 728 1623 730 1633
rect 800 1623 802 1633
rect 872 1623 874 1633
rect 944 1623 946 1633
rect 1024 1623 1026 1633
rect 1104 1623 1106 1633
rect 1176 1623 1178 1633
rect 1248 1623 1250 1633
rect 1320 1623 1322 1633
rect 1400 1623 1402 1633
rect 1480 1623 1482 1633
rect 1560 1623 1562 1633
rect 1624 1623 1626 1633
rect 1664 1625 1666 1633
rect 1662 1624 1668 1625
rect 110 1619 116 1620
rect 134 1622 140 1623
rect 134 1618 135 1622
rect 139 1618 140 1622
rect 134 1617 140 1618
rect 182 1622 188 1623
rect 182 1618 183 1622
rect 187 1618 188 1622
rect 182 1617 188 1618
rect 246 1622 252 1623
rect 246 1618 247 1622
rect 251 1618 252 1622
rect 246 1617 252 1618
rect 302 1622 308 1623
rect 302 1618 303 1622
rect 307 1618 308 1622
rect 302 1617 308 1618
rect 358 1622 364 1623
rect 358 1618 359 1622
rect 363 1618 364 1622
rect 358 1617 364 1618
rect 414 1622 420 1623
rect 414 1618 415 1622
rect 419 1618 420 1622
rect 414 1617 420 1618
rect 470 1622 476 1623
rect 470 1618 471 1622
rect 475 1618 476 1622
rect 470 1617 476 1618
rect 534 1622 540 1623
rect 534 1618 535 1622
rect 539 1618 540 1622
rect 534 1617 540 1618
rect 598 1622 604 1623
rect 598 1618 599 1622
rect 603 1618 604 1622
rect 598 1617 604 1618
rect 662 1622 668 1623
rect 662 1618 663 1622
rect 667 1618 668 1622
rect 662 1617 668 1618
rect 726 1622 732 1623
rect 726 1618 727 1622
rect 731 1618 732 1622
rect 726 1617 732 1618
rect 798 1622 804 1623
rect 798 1618 799 1622
rect 803 1618 804 1622
rect 798 1617 804 1618
rect 870 1622 876 1623
rect 870 1618 871 1622
rect 875 1618 876 1622
rect 870 1617 876 1618
rect 942 1622 948 1623
rect 942 1618 943 1622
rect 947 1618 948 1622
rect 942 1617 948 1618
rect 1022 1622 1028 1623
rect 1022 1618 1023 1622
rect 1027 1618 1028 1622
rect 1022 1617 1028 1618
rect 1102 1622 1108 1623
rect 1102 1618 1103 1622
rect 1107 1618 1108 1622
rect 1102 1617 1108 1618
rect 1174 1622 1180 1623
rect 1174 1618 1175 1622
rect 1179 1618 1180 1622
rect 1174 1617 1180 1618
rect 1246 1622 1252 1623
rect 1246 1618 1247 1622
rect 1251 1618 1252 1622
rect 1246 1617 1252 1618
rect 1318 1622 1324 1623
rect 1318 1618 1319 1622
rect 1323 1618 1324 1622
rect 1318 1617 1324 1618
rect 1398 1622 1404 1623
rect 1398 1618 1399 1622
rect 1403 1618 1404 1622
rect 1398 1617 1404 1618
rect 1478 1622 1484 1623
rect 1478 1618 1479 1622
rect 1483 1618 1484 1622
rect 1478 1617 1484 1618
rect 1558 1622 1564 1623
rect 1558 1618 1559 1622
rect 1563 1618 1564 1622
rect 1558 1617 1564 1618
rect 1622 1622 1628 1623
rect 1622 1618 1623 1622
rect 1627 1618 1628 1622
rect 1662 1620 1663 1624
rect 1667 1620 1668 1624
rect 1662 1619 1668 1620
rect 1622 1617 1628 1618
rect 110 1607 116 1608
rect 110 1603 111 1607
rect 115 1603 116 1607
rect 1662 1607 1668 1608
rect 110 1602 116 1603
rect 134 1605 140 1606
rect 112 1599 114 1602
rect 134 1601 135 1605
rect 139 1601 140 1605
rect 134 1600 140 1601
rect 182 1605 188 1606
rect 182 1601 183 1605
rect 187 1601 188 1605
rect 182 1600 188 1601
rect 246 1605 252 1606
rect 246 1601 247 1605
rect 251 1601 252 1605
rect 246 1600 252 1601
rect 302 1605 308 1606
rect 302 1601 303 1605
rect 307 1601 308 1605
rect 302 1600 308 1601
rect 358 1605 364 1606
rect 358 1601 359 1605
rect 363 1601 364 1605
rect 358 1600 364 1601
rect 414 1605 420 1606
rect 414 1601 415 1605
rect 419 1601 420 1605
rect 414 1600 420 1601
rect 470 1605 476 1606
rect 470 1601 471 1605
rect 475 1601 476 1605
rect 470 1600 476 1601
rect 534 1605 540 1606
rect 534 1601 535 1605
rect 539 1601 540 1605
rect 534 1600 540 1601
rect 598 1605 604 1606
rect 598 1601 599 1605
rect 603 1601 604 1605
rect 598 1600 604 1601
rect 662 1605 668 1606
rect 662 1601 663 1605
rect 667 1601 668 1605
rect 662 1600 668 1601
rect 726 1605 732 1606
rect 726 1601 727 1605
rect 731 1601 732 1605
rect 726 1600 732 1601
rect 798 1605 804 1606
rect 798 1601 799 1605
rect 803 1601 804 1605
rect 798 1600 804 1601
rect 870 1605 876 1606
rect 870 1601 871 1605
rect 875 1601 876 1605
rect 870 1600 876 1601
rect 942 1605 948 1606
rect 942 1601 943 1605
rect 947 1601 948 1605
rect 942 1600 948 1601
rect 1022 1605 1028 1606
rect 1022 1601 1023 1605
rect 1027 1601 1028 1605
rect 1022 1600 1028 1601
rect 1102 1605 1108 1606
rect 1102 1601 1103 1605
rect 1107 1601 1108 1605
rect 1102 1600 1108 1601
rect 1174 1605 1180 1606
rect 1174 1601 1175 1605
rect 1179 1601 1180 1605
rect 1174 1600 1180 1601
rect 1246 1605 1252 1606
rect 1246 1601 1247 1605
rect 1251 1601 1252 1605
rect 1246 1600 1252 1601
rect 1318 1605 1324 1606
rect 1318 1601 1319 1605
rect 1323 1601 1324 1605
rect 1318 1600 1324 1601
rect 1398 1605 1404 1606
rect 1398 1601 1399 1605
rect 1403 1601 1404 1605
rect 1398 1600 1404 1601
rect 1478 1605 1484 1606
rect 1478 1601 1479 1605
rect 1483 1601 1484 1605
rect 1478 1600 1484 1601
rect 1558 1605 1564 1606
rect 1558 1601 1559 1605
rect 1563 1601 1564 1605
rect 1558 1600 1564 1601
rect 1622 1605 1628 1606
rect 1622 1601 1623 1605
rect 1627 1601 1628 1605
rect 1662 1603 1663 1607
rect 1667 1603 1668 1607
rect 1662 1602 1668 1603
rect 1622 1600 1628 1601
rect 111 1598 115 1599
rect 111 1593 115 1594
rect 135 1598 139 1600
rect 112 1590 114 1593
rect 135 1592 139 1594
rect 167 1598 171 1599
rect 167 1592 171 1594
rect 183 1598 187 1600
rect 183 1593 187 1594
rect 223 1598 227 1599
rect 223 1592 227 1594
rect 247 1598 251 1600
rect 247 1593 251 1594
rect 279 1598 283 1599
rect 279 1592 283 1594
rect 303 1598 307 1600
rect 303 1593 307 1594
rect 335 1598 339 1599
rect 335 1592 339 1594
rect 359 1598 363 1600
rect 359 1593 363 1594
rect 383 1598 387 1599
rect 383 1592 387 1594
rect 415 1598 419 1600
rect 415 1593 419 1594
rect 431 1598 435 1599
rect 431 1592 435 1594
rect 471 1598 475 1600
rect 471 1593 475 1594
rect 479 1598 483 1599
rect 479 1592 483 1594
rect 535 1598 539 1600
rect 535 1592 539 1594
rect 599 1598 603 1600
rect 599 1592 603 1594
rect 663 1598 667 1600
rect 663 1592 667 1594
rect 727 1598 731 1600
rect 727 1592 731 1594
rect 799 1598 803 1600
rect 799 1592 803 1594
rect 871 1598 875 1600
rect 871 1592 875 1594
rect 943 1598 947 1600
rect 943 1593 947 1594
rect 951 1598 955 1599
rect 951 1592 955 1594
rect 1023 1598 1027 1600
rect 1023 1593 1027 1594
rect 1039 1598 1043 1599
rect 1039 1592 1043 1594
rect 1103 1598 1107 1600
rect 1103 1593 1107 1594
rect 1119 1598 1123 1599
rect 1119 1592 1123 1594
rect 1175 1598 1179 1600
rect 1175 1593 1179 1594
rect 1199 1598 1203 1599
rect 1199 1592 1203 1594
rect 1247 1598 1251 1600
rect 1247 1593 1251 1594
rect 1279 1598 1283 1599
rect 1279 1592 1283 1594
rect 1319 1598 1323 1600
rect 1319 1593 1323 1594
rect 1351 1598 1355 1599
rect 1351 1592 1355 1594
rect 1399 1598 1403 1600
rect 1399 1593 1403 1594
rect 1415 1598 1419 1599
rect 1415 1592 1419 1594
rect 1471 1598 1475 1599
rect 1471 1592 1475 1594
rect 1479 1598 1483 1600
rect 1479 1593 1483 1594
rect 1527 1598 1531 1599
rect 1527 1592 1531 1594
rect 1559 1598 1563 1600
rect 1559 1593 1563 1594
rect 1583 1598 1587 1599
rect 1583 1592 1587 1594
rect 1623 1598 1627 1600
rect 1664 1599 1666 1602
rect 1623 1592 1627 1594
rect 1663 1598 1667 1599
rect 1663 1593 1667 1594
rect 134 1591 140 1592
rect 110 1589 116 1590
rect 110 1585 111 1589
rect 115 1585 116 1589
rect 134 1587 135 1591
rect 139 1587 140 1591
rect 134 1586 140 1587
rect 166 1591 172 1592
rect 166 1587 167 1591
rect 171 1587 172 1591
rect 166 1586 172 1587
rect 222 1591 228 1592
rect 222 1587 223 1591
rect 227 1587 228 1591
rect 222 1586 228 1587
rect 278 1591 284 1592
rect 278 1587 279 1591
rect 283 1587 284 1591
rect 278 1586 284 1587
rect 334 1591 340 1592
rect 334 1587 335 1591
rect 339 1587 340 1591
rect 334 1586 340 1587
rect 382 1591 388 1592
rect 382 1587 383 1591
rect 387 1587 388 1591
rect 382 1586 388 1587
rect 430 1591 436 1592
rect 430 1587 431 1591
rect 435 1587 436 1591
rect 430 1586 436 1587
rect 478 1591 484 1592
rect 478 1587 479 1591
rect 483 1587 484 1591
rect 478 1586 484 1587
rect 534 1591 540 1592
rect 534 1587 535 1591
rect 539 1587 540 1591
rect 534 1586 540 1587
rect 598 1591 604 1592
rect 598 1587 599 1591
rect 603 1587 604 1591
rect 598 1586 604 1587
rect 662 1591 668 1592
rect 662 1587 663 1591
rect 667 1587 668 1591
rect 662 1586 668 1587
rect 726 1591 732 1592
rect 726 1587 727 1591
rect 731 1587 732 1591
rect 726 1586 732 1587
rect 798 1591 804 1592
rect 798 1587 799 1591
rect 803 1587 804 1591
rect 798 1586 804 1587
rect 870 1591 876 1592
rect 870 1587 871 1591
rect 875 1587 876 1591
rect 870 1586 876 1587
rect 950 1591 956 1592
rect 950 1587 951 1591
rect 955 1587 956 1591
rect 950 1586 956 1587
rect 1038 1591 1044 1592
rect 1038 1587 1039 1591
rect 1043 1587 1044 1591
rect 1038 1586 1044 1587
rect 1118 1591 1124 1592
rect 1118 1587 1119 1591
rect 1123 1587 1124 1591
rect 1118 1586 1124 1587
rect 1198 1591 1204 1592
rect 1198 1587 1199 1591
rect 1203 1587 1204 1591
rect 1198 1586 1204 1587
rect 1278 1591 1284 1592
rect 1278 1587 1279 1591
rect 1283 1587 1284 1591
rect 1278 1586 1284 1587
rect 1350 1591 1356 1592
rect 1350 1587 1351 1591
rect 1355 1587 1356 1591
rect 1350 1586 1356 1587
rect 1414 1591 1420 1592
rect 1414 1587 1415 1591
rect 1419 1587 1420 1591
rect 1414 1586 1420 1587
rect 1470 1591 1476 1592
rect 1470 1587 1471 1591
rect 1475 1587 1476 1591
rect 1470 1586 1476 1587
rect 1526 1591 1532 1592
rect 1526 1587 1527 1591
rect 1531 1587 1532 1591
rect 1526 1586 1532 1587
rect 1582 1591 1588 1592
rect 1582 1587 1583 1591
rect 1587 1587 1588 1591
rect 1582 1586 1588 1587
rect 1622 1591 1628 1592
rect 1622 1587 1623 1591
rect 1627 1587 1628 1591
rect 1664 1590 1666 1593
rect 1622 1586 1628 1587
rect 1662 1589 1668 1590
rect 110 1584 116 1585
rect 1662 1585 1663 1589
rect 1667 1585 1668 1589
rect 1662 1584 1668 1585
rect 134 1574 140 1575
rect 110 1572 116 1573
rect 110 1568 111 1572
rect 115 1568 116 1572
rect 134 1570 135 1574
rect 139 1570 140 1574
rect 134 1569 140 1570
rect 166 1574 172 1575
rect 166 1570 167 1574
rect 171 1570 172 1574
rect 166 1569 172 1570
rect 222 1574 228 1575
rect 222 1570 223 1574
rect 227 1570 228 1574
rect 222 1569 228 1570
rect 278 1574 284 1575
rect 278 1570 279 1574
rect 283 1570 284 1574
rect 278 1569 284 1570
rect 334 1574 340 1575
rect 334 1570 335 1574
rect 339 1570 340 1574
rect 334 1569 340 1570
rect 382 1574 388 1575
rect 382 1570 383 1574
rect 387 1570 388 1574
rect 382 1569 388 1570
rect 430 1574 436 1575
rect 430 1570 431 1574
rect 435 1570 436 1574
rect 430 1569 436 1570
rect 478 1574 484 1575
rect 478 1570 479 1574
rect 483 1570 484 1574
rect 478 1569 484 1570
rect 534 1574 540 1575
rect 534 1570 535 1574
rect 539 1570 540 1574
rect 534 1569 540 1570
rect 598 1574 604 1575
rect 598 1570 599 1574
rect 603 1570 604 1574
rect 598 1569 604 1570
rect 662 1574 668 1575
rect 662 1570 663 1574
rect 667 1570 668 1574
rect 662 1569 668 1570
rect 726 1574 732 1575
rect 726 1570 727 1574
rect 731 1570 732 1574
rect 726 1569 732 1570
rect 798 1574 804 1575
rect 798 1570 799 1574
rect 803 1570 804 1574
rect 798 1569 804 1570
rect 870 1574 876 1575
rect 870 1570 871 1574
rect 875 1570 876 1574
rect 870 1569 876 1570
rect 950 1574 956 1575
rect 950 1570 951 1574
rect 955 1570 956 1574
rect 950 1569 956 1570
rect 1038 1574 1044 1575
rect 1038 1570 1039 1574
rect 1043 1570 1044 1574
rect 1038 1569 1044 1570
rect 1118 1574 1124 1575
rect 1118 1570 1119 1574
rect 1123 1570 1124 1574
rect 1118 1569 1124 1570
rect 1198 1574 1204 1575
rect 1198 1570 1199 1574
rect 1203 1570 1204 1574
rect 1198 1569 1204 1570
rect 1278 1574 1284 1575
rect 1278 1570 1279 1574
rect 1283 1570 1284 1574
rect 1278 1569 1284 1570
rect 1350 1574 1356 1575
rect 1350 1570 1351 1574
rect 1355 1570 1356 1574
rect 1350 1569 1356 1570
rect 1414 1574 1420 1575
rect 1414 1570 1415 1574
rect 1419 1570 1420 1574
rect 1414 1569 1420 1570
rect 1470 1574 1476 1575
rect 1470 1570 1471 1574
rect 1475 1570 1476 1574
rect 1470 1569 1476 1570
rect 1526 1574 1532 1575
rect 1526 1570 1527 1574
rect 1531 1570 1532 1574
rect 1526 1569 1532 1570
rect 1582 1574 1588 1575
rect 1582 1570 1583 1574
rect 1587 1570 1588 1574
rect 1582 1569 1588 1570
rect 1622 1574 1628 1575
rect 1622 1570 1623 1574
rect 1627 1570 1628 1574
rect 1622 1569 1628 1570
rect 1662 1572 1668 1573
rect 110 1567 116 1568
rect 112 1559 114 1567
rect 136 1559 138 1569
rect 168 1559 170 1569
rect 224 1559 226 1569
rect 280 1559 282 1569
rect 336 1559 338 1569
rect 384 1559 386 1569
rect 432 1559 434 1569
rect 480 1559 482 1569
rect 536 1559 538 1569
rect 600 1559 602 1569
rect 664 1559 666 1569
rect 728 1559 730 1569
rect 800 1559 802 1569
rect 872 1559 874 1569
rect 952 1559 954 1569
rect 1040 1559 1042 1569
rect 1120 1559 1122 1569
rect 1200 1559 1202 1569
rect 1280 1559 1282 1569
rect 1352 1559 1354 1569
rect 1416 1559 1418 1569
rect 1472 1559 1474 1569
rect 1528 1559 1530 1569
rect 1584 1559 1586 1569
rect 1624 1559 1626 1569
rect 1662 1568 1663 1572
rect 1667 1568 1668 1572
rect 1662 1567 1668 1568
rect 1664 1559 1666 1567
rect 111 1558 115 1559
rect 111 1553 115 1554
rect 135 1558 139 1559
rect 135 1553 139 1554
rect 167 1558 171 1559
rect 167 1553 171 1554
rect 215 1558 219 1559
rect 215 1553 219 1554
rect 223 1558 227 1559
rect 223 1553 227 1554
rect 263 1558 267 1559
rect 263 1553 267 1554
rect 279 1558 283 1559
rect 279 1553 283 1554
rect 311 1558 315 1559
rect 311 1553 315 1554
rect 335 1558 339 1559
rect 335 1553 339 1554
rect 359 1558 363 1559
rect 359 1553 363 1554
rect 383 1558 387 1559
rect 383 1553 387 1554
rect 407 1558 411 1559
rect 407 1553 411 1554
rect 431 1558 435 1559
rect 431 1553 435 1554
rect 455 1558 459 1559
rect 455 1553 459 1554
rect 479 1558 483 1559
rect 479 1553 483 1554
rect 511 1558 515 1559
rect 511 1553 515 1554
rect 535 1558 539 1559
rect 535 1553 539 1554
rect 567 1558 571 1559
rect 567 1553 571 1554
rect 599 1558 603 1559
rect 599 1553 603 1554
rect 631 1558 635 1559
rect 631 1553 635 1554
rect 663 1558 667 1559
rect 663 1553 667 1554
rect 695 1558 699 1559
rect 695 1553 699 1554
rect 727 1558 731 1559
rect 727 1553 731 1554
rect 759 1558 763 1559
rect 759 1553 763 1554
rect 799 1558 803 1559
rect 799 1553 803 1554
rect 831 1558 835 1559
rect 831 1553 835 1554
rect 871 1558 875 1559
rect 871 1553 875 1554
rect 919 1558 923 1559
rect 919 1553 923 1554
rect 951 1558 955 1559
rect 951 1553 955 1554
rect 1007 1558 1011 1559
rect 1007 1553 1011 1554
rect 1039 1558 1043 1559
rect 1039 1553 1043 1554
rect 1095 1558 1099 1559
rect 1095 1553 1099 1554
rect 1119 1558 1123 1559
rect 1119 1553 1123 1554
rect 1183 1558 1187 1559
rect 1183 1553 1187 1554
rect 1199 1558 1203 1559
rect 1199 1553 1203 1554
rect 1263 1558 1267 1559
rect 1263 1553 1267 1554
rect 1279 1558 1283 1559
rect 1279 1553 1283 1554
rect 1335 1558 1339 1559
rect 1335 1553 1339 1554
rect 1351 1558 1355 1559
rect 1351 1553 1355 1554
rect 1407 1558 1411 1559
rect 1407 1553 1411 1554
rect 1415 1558 1419 1559
rect 1415 1553 1419 1554
rect 1471 1558 1475 1559
rect 1471 1553 1475 1554
rect 1527 1558 1531 1559
rect 1527 1553 1531 1554
rect 1583 1558 1587 1559
rect 1583 1553 1587 1554
rect 1623 1558 1627 1559
rect 1623 1553 1627 1554
rect 1663 1558 1667 1559
rect 1663 1553 1667 1554
rect 112 1545 114 1553
rect 110 1544 116 1545
rect 110 1540 111 1544
rect 115 1540 116 1544
rect 136 1543 138 1553
rect 168 1543 170 1553
rect 216 1543 218 1553
rect 264 1543 266 1553
rect 312 1543 314 1553
rect 360 1543 362 1553
rect 408 1543 410 1553
rect 456 1543 458 1553
rect 512 1543 514 1553
rect 568 1543 570 1553
rect 632 1543 634 1553
rect 696 1543 698 1553
rect 760 1543 762 1553
rect 832 1543 834 1553
rect 920 1543 922 1553
rect 1008 1543 1010 1553
rect 1096 1543 1098 1553
rect 1184 1543 1186 1553
rect 1264 1543 1266 1553
rect 1336 1543 1338 1553
rect 1408 1543 1410 1553
rect 1472 1543 1474 1553
rect 1528 1543 1530 1553
rect 1584 1543 1586 1553
rect 1624 1543 1626 1553
rect 1664 1545 1666 1553
rect 1662 1544 1668 1545
rect 110 1539 116 1540
rect 134 1542 140 1543
rect 134 1538 135 1542
rect 139 1538 140 1542
rect 134 1537 140 1538
rect 166 1542 172 1543
rect 166 1538 167 1542
rect 171 1538 172 1542
rect 166 1537 172 1538
rect 214 1542 220 1543
rect 214 1538 215 1542
rect 219 1538 220 1542
rect 214 1537 220 1538
rect 262 1542 268 1543
rect 262 1538 263 1542
rect 267 1538 268 1542
rect 262 1537 268 1538
rect 310 1542 316 1543
rect 310 1538 311 1542
rect 315 1538 316 1542
rect 310 1537 316 1538
rect 358 1542 364 1543
rect 358 1538 359 1542
rect 363 1538 364 1542
rect 358 1537 364 1538
rect 406 1542 412 1543
rect 406 1538 407 1542
rect 411 1538 412 1542
rect 406 1537 412 1538
rect 454 1542 460 1543
rect 454 1538 455 1542
rect 459 1538 460 1542
rect 454 1537 460 1538
rect 510 1542 516 1543
rect 510 1538 511 1542
rect 515 1538 516 1542
rect 510 1537 516 1538
rect 566 1542 572 1543
rect 566 1538 567 1542
rect 571 1538 572 1542
rect 566 1537 572 1538
rect 630 1542 636 1543
rect 630 1538 631 1542
rect 635 1538 636 1542
rect 630 1537 636 1538
rect 694 1542 700 1543
rect 694 1538 695 1542
rect 699 1538 700 1542
rect 694 1537 700 1538
rect 758 1542 764 1543
rect 758 1538 759 1542
rect 763 1538 764 1542
rect 758 1537 764 1538
rect 830 1542 836 1543
rect 830 1538 831 1542
rect 835 1538 836 1542
rect 830 1537 836 1538
rect 918 1542 924 1543
rect 918 1538 919 1542
rect 923 1538 924 1542
rect 918 1537 924 1538
rect 1006 1542 1012 1543
rect 1006 1538 1007 1542
rect 1011 1538 1012 1542
rect 1006 1537 1012 1538
rect 1094 1542 1100 1543
rect 1094 1538 1095 1542
rect 1099 1538 1100 1542
rect 1094 1537 1100 1538
rect 1182 1542 1188 1543
rect 1182 1538 1183 1542
rect 1187 1538 1188 1542
rect 1182 1537 1188 1538
rect 1262 1542 1268 1543
rect 1262 1538 1263 1542
rect 1267 1538 1268 1542
rect 1262 1537 1268 1538
rect 1334 1542 1340 1543
rect 1334 1538 1335 1542
rect 1339 1538 1340 1542
rect 1334 1537 1340 1538
rect 1406 1542 1412 1543
rect 1406 1538 1407 1542
rect 1411 1538 1412 1542
rect 1406 1537 1412 1538
rect 1470 1542 1476 1543
rect 1470 1538 1471 1542
rect 1475 1538 1476 1542
rect 1470 1537 1476 1538
rect 1526 1542 1532 1543
rect 1526 1538 1527 1542
rect 1531 1538 1532 1542
rect 1526 1537 1532 1538
rect 1582 1542 1588 1543
rect 1582 1538 1583 1542
rect 1587 1538 1588 1542
rect 1582 1537 1588 1538
rect 1622 1542 1628 1543
rect 1622 1538 1623 1542
rect 1627 1538 1628 1542
rect 1662 1540 1663 1544
rect 1667 1540 1668 1544
rect 1662 1539 1668 1540
rect 1622 1537 1628 1538
rect 110 1527 116 1528
rect 110 1523 111 1527
rect 115 1523 116 1527
rect 1662 1527 1668 1528
rect 110 1522 116 1523
rect 134 1525 140 1526
rect 112 1515 114 1522
rect 134 1521 135 1525
rect 139 1521 140 1525
rect 134 1520 140 1521
rect 166 1525 172 1526
rect 166 1521 167 1525
rect 171 1521 172 1525
rect 166 1520 172 1521
rect 214 1525 220 1526
rect 214 1521 215 1525
rect 219 1521 220 1525
rect 214 1520 220 1521
rect 262 1525 268 1526
rect 262 1521 263 1525
rect 267 1521 268 1525
rect 262 1520 268 1521
rect 310 1525 316 1526
rect 310 1521 311 1525
rect 315 1521 316 1525
rect 310 1520 316 1521
rect 358 1525 364 1526
rect 358 1521 359 1525
rect 363 1521 364 1525
rect 358 1520 364 1521
rect 406 1525 412 1526
rect 406 1521 407 1525
rect 411 1521 412 1525
rect 406 1520 412 1521
rect 454 1525 460 1526
rect 454 1521 455 1525
rect 459 1521 460 1525
rect 454 1520 460 1521
rect 510 1525 516 1526
rect 510 1521 511 1525
rect 515 1521 516 1525
rect 510 1520 516 1521
rect 566 1525 572 1526
rect 566 1521 567 1525
rect 571 1521 572 1525
rect 566 1520 572 1521
rect 630 1525 636 1526
rect 630 1521 631 1525
rect 635 1521 636 1525
rect 630 1520 636 1521
rect 694 1525 700 1526
rect 694 1521 695 1525
rect 699 1521 700 1525
rect 694 1520 700 1521
rect 758 1525 764 1526
rect 758 1521 759 1525
rect 763 1521 764 1525
rect 758 1520 764 1521
rect 830 1525 836 1526
rect 830 1521 831 1525
rect 835 1521 836 1525
rect 830 1520 836 1521
rect 918 1525 924 1526
rect 918 1521 919 1525
rect 923 1521 924 1525
rect 918 1520 924 1521
rect 1006 1525 1012 1526
rect 1006 1521 1007 1525
rect 1011 1521 1012 1525
rect 1006 1520 1012 1521
rect 1094 1525 1100 1526
rect 1094 1521 1095 1525
rect 1099 1521 1100 1525
rect 1094 1520 1100 1521
rect 1182 1525 1188 1526
rect 1182 1521 1183 1525
rect 1187 1521 1188 1525
rect 1182 1520 1188 1521
rect 1262 1525 1268 1526
rect 1262 1521 1263 1525
rect 1267 1521 1268 1525
rect 1262 1520 1268 1521
rect 1334 1525 1340 1526
rect 1334 1521 1335 1525
rect 1339 1521 1340 1525
rect 1334 1520 1340 1521
rect 1406 1525 1412 1526
rect 1406 1521 1407 1525
rect 1411 1521 1412 1525
rect 1406 1520 1412 1521
rect 1470 1525 1476 1526
rect 1470 1521 1471 1525
rect 1475 1521 1476 1525
rect 1470 1520 1476 1521
rect 1526 1525 1532 1526
rect 1526 1521 1527 1525
rect 1531 1521 1532 1525
rect 1526 1520 1532 1521
rect 1582 1525 1588 1526
rect 1582 1521 1583 1525
rect 1587 1521 1588 1525
rect 1582 1520 1588 1521
rect 1622 1525 1628 1526
rect 1622 1521 1623 1525
rect 1627 1521 1628 1525
rect 1662 1523 1663 1527
rect 1667 1523 1668 1527
rect 1662 1522 1668 1523
rect 1622 1520 1628 1521
rect 136 1515 138 1520
rect 168 1515 170 1520
rect 216 1515 218 1520
rect 264 1515 266 1520
rect 312 1515 314 1520
rect 360 1515 362 1520
rect 408 1515 410 1520
rect 456 1515 458 1520
rect 512 1515 514 1520
rect 568 1515 570 1520
rect 632 1515 634 1520
rect 696 1515 698 1520
rect 760 1515 762 1520
rect 832 1515 834 1520
rect 920 1515 922 1520
rect 1008 1515 1010 1520
rect 1096 1515 1098 1520
rect 1184 1515 1186 1520
rect 1264 1515 1266 1520
rect 1336 1515 1338 1520
rect 1408 1515 1410 1520
rect 1472 1515 1474 1520
rect 1528 1515 1530 1520
rect 1584 1515 1586 1520
rect 1624 1515 1626 1520
rect 1664 1515 1666 1522
rect 111 1514 115 1515
rect 111 1509 115 1510
rect 135 1514 139 1515
rect 112 1506 114 1509
rect 135 1508 139 1510
rect 167 1514 171 1515
rect 167 1508 171 1510
rect 215 1514 219 1515
rect 215 1509 219 1510
rect 223 1514 227 1515
rect 223 1508 227 1510
rect 263 1514 267 1515
rect 263 1509 267 1510
rect 295 1514 299 1515
rect 295 1508 299 1510
rect 311 1514 315 1515
rect 311 1509 315 1510
rect 359 1514 363 1515
rect 359 1509 363 1510
rect 375 1514 379 1515
rect 375 1508 379 1510
rect 407 1514 411 1515
rect 407 1509 411 1510
rect 455 1514 459 1515
rect 455 1508 459 1510
rect 511 1514 515 1515
rect 511 1509 515 1510
rect 527 1514 531 1515
rect 527 1508 531 1510
rect 567 1514 571 1515
rect 567 1509 571 1510
rect 599 1514 603 1515
rect 599 1508 603 1510
rect 631 1514 635 1515
rect 631 1509 635 1510
rect 671 1514 675 1515
rect 671 1508 675 1510
rect 695 1514 699 1515
rect 695 1509 699 1510
rect 743 1514 747 1515
rect 743 1508 747 1510
rect 759 1514 763 1515
rect 759 1509 763 1510
rect 815 1514 819 1515
rect 815 1508 819 1510
rect 831 1514 835 1515
rect 831 1509 835 1510
rect 879 1514 883 1515
rect 879 1508 883 1510
rect 919 1514 923 1515
rect 919 1509 923 1510
rect 943 1514 947 1515
rect 943 1508 947 1510
rect 1007 1514 1011 1515
rect 1007 1508 1011 1510
rect 1063 1514 1067 1515
rect 1063 1508 1067 1510
rect 1095 1514 1099 1515
rect 1095 1509 1099 1510
rect 1111 1514 1115 1515
rect 1111 1508 1115 1510
rect 1151 1514 1155 1515
rect 1151 1508 1155 1510
rect 1183 1514 1187 1515
rect 1183 1508 1187 1510
rect 1215 1514 1219 1515
rect 1215 1508 1219 1510
rect 1255 1514 1259 1515
rect 1255 1508 1259 1510
rect 1263 1514 1267 1515
rect 1263 1509 1267 1510
rect 1295 1514 1299 1515
rect 1295 1508 1299 1510
rect 1335 1514 1339 1515
rect 1335 1509 1339 1510
rect 1351 1514 1355 1515
rect 1351 1508 1355 1510
rect 1407 1514 1411 1515
rect 1407 1509 1411 1510
rect 1415 1514 1419 1515
rect 1415 1508 1419 1510
rect 1471 1514 1475 1515
rect 1471 1509 1475 1510
rect 1487 1514 1491 1515
rect 1487 1508 1491 1510
rect 1527 1514 1531 1515
rect 1527 1509 1531 1510
rect 1567 1514 1571 1515
rect 1567 1508 1571 1510
rect 1583 1514 1587 1515
rect 1583 1509 1587 1510
rect 1623 1514 1627 1515
rect 1623 1508 1627 1510
rect 1663 1514 1667 1515
rect 1663 1509 1667 1510
rect 134 1507 140 1508
rect 110 1505 116 1506
rect 110 1501 111 1505
rect 115 1501 116 1505
rect 134 1503 135 1507
rect 139 1503 140 1507
rect 134 1502 140 1503
rect 166 1507 172 1508
rect 166 1503 167 1507
rect 171 1503 172 1507
rect 166 1502 172 1503
rect 222 1507 228 1508
rect 222 1503 223 1507
rect 227 1503 228 1507
rect 222 1502 228 1503
rect 294 1507 300 1508
rect 294 1503 295 1507
rect 299 1503 300 1507
rect 294 1502 300 1503
rect 374 1507 380 1508
rect 374 1503 375 1507
rect 379 1503 380 1507
rect 374 1502 380 1503
rect 454 1507 460 1508
rect 454 1503 455 1507
rect 459 1503 460 1507
rect 454 1502 460 1503
rect 526 1507 532 1508
rect 526 1503 527 1507
rect 531 1503 532 1507
rect 526 1502 532 1503
rect 598 1507 604 1508
rect 598 1503 599 1507
rect 603 1503 604 1507
rect 598 1502 604 1503
rect 670 1507 676 1508
rect 670 1503 671 1507
rect 675 1503 676 1507
rect 670 1502 676 1503
rect 742 1507 748 1508
rect 742 1503 743 1507
rect 747 1503 748 1507
rect 742 1502 748 1503
rect 814 1507 820 1508
rect 814 1503 815 1507
rect 819 1503 820 1507
rect 814 1502 820 1503
rect 878 1507 884 1508
rect 878 1503 879 1507
rect 883 1503 884 1507
rect 878 1502 884 1503
rect 942 1507 948 1508
rect 942 1503 943 1507
rect 947 1503 948 1507
rect 942 1502 948 1503
rect 1006 1507 1012 1508
rect 1006 1503 1007 1507
rect 1011 1503 1012 1507
rect 1006 1502 1012 1503
rect 1062 1507 1068 1508
rect 1062 1503 1063 1507
rect 1067 1503 1068 1507
rect 1062 1502 1068 1503
rect 1110 1507 1116 1508
rect 1110 1503 1111 1507
rect 1115 1503 1116 1507
rect 1110 1502 1116 1503
rect 1150 1507 1156 1508
rect 1150 1503 1151 1507
rect 1155 1503 1156 1507
rect 1150 1502 1156 1503
rect 1182 1507 1188 1508
rect 1182 1503 1183 1507
rect 1187 1503 1188 1507
rect 1182 1502 1188 1503
rect 1214 1507 1220 1508
rect 1214 1503 1215 1507
rect 1219 1503 1220 1507
rect 1214 1502 1220 1503
rect 1254 1507 1260 1508
rect 1254 1503 1255 1507
rect 1259 1503 1260 1507
rect 1254 1502 1260 1503
rect 1294 1507 1300 1508
rect 1294 1503 1295 1507
rect 1299 1503 1300 1507
rect 1294 1502 1300 1503
rect 1350 1507 1356 1508
rect 1350 1503 1351 1507
rect 1355 1503 1356 1507
rect 1350 1502 1356 1503
rect 1414 1507 1420 1508
rect 1414 1503 1415 1507
rect 1419 1503 1420 1507
rect 1414 1502 1420 1503
rect 1486 1507 1492 1508
rect 1486 1503 1487 1507
rect 1491 1503 1492 1507
rect 1486 1502 1492 1503
rect 1566 1507 1572 1508
rect 1566 1503 1567 1507
rect 1571 1503 1572 1507
rect 1566 1502 1572 1503
rect 1622 1507 1628 1508
rect 1622 1503 1623 1507
rect 1627 1503 1628 1507
rect 1664 1506 1666 1509
rect 1622 1502 1628 1503
rect 1662 1505 1668 1506
rect 110 1500 116 1501
rect 1662 1501 1663 1505
rect 1667 1501 1668 1505
rect 1662 1500 1668 1501
rect 134 1490 140 1491
rect 110 1488 116 1489
rect 110 1484 111 1488
rect 115 1484 116 1488
rect 134 1486 135 1490
rect 139 1486 140 1490
rect 134 1485 140 1486
rect 166 1490 172 1491
rect 166 1486 167 1490
rect 171 1486 172 1490
rect 166 1485 172 1486
rect 222 1490 228 1491
rect 222 1486 223 1490
rect 227 1486 228 1490
rect 222 1485 228 1486
rect 294 1490 300 1491
rect 294 1486 295 1490
rect 299 1486 300 1490
rect 294 1485 300 1486
rect 374 1490 380 1491
rect 374 1486 375 1490
rect 379 1486 380 1490
rect 374 1485 380 1486
rect 454 1490 460 1491
rect 454 1486 455 1490
rect 459 1486 460 1490
rect 454 1485 460 1486
rect 526 1490 532 1491
rect 526 1486 527 1490
rect 531 1486 532 1490
rect 526 1485 532 1486
rect 598 1490 604 1491
rect 598 1486 599 1490
rect 603 1486 604 1490
rect 598 1485 604 1486
rect 670 1490 676 1491
rect 670 1486 671 1490
rect 675 1486 676 1490
rect 670 1485 676 1486
rect 742 1490 748 1491
rect 742 1486 743 1490
rect 747 1486 748 1490
rect 742 1485 748 1486
rect 814 1490 820 1491
rect 814 1486 815 1490
rect 819 1486 820 1490
rect 814 1485 820 1486
rect 878 1490 884 1491
rect 878 1486 879 1490
rect 883 1486 884 1490
rect 878 1485 884 1486
rect 942 1490 948 1491
rect 942 1486 943 1490
rect 947 1486 948 1490
rect 942 1485 948 1486
rect 1006 1490 1012 1491
rect 1006 1486 1007 1490
rect 1011 1486 1012 1490
rect 1006 1485 1012 1486
rect 1062 1490 1068 1491
rect 1062 1486 1063 1490
rect 1067 1486 1068 1490
rect 1062 1485 1068 1486
rect 1110 1490 1116 1491
rect 1110 1486 1111 1490
rect 1115 1486 1116 1490
rect 1110 1485 1116 1486
rect 1150 1490 1156 1491
rect 1150 1486 1151 1490
rect 1155 1486 1156 1490
rect 1150 1485 1156 1486
rect 1182 1490 1188 1491
rect 1182 1486 1183 1490
rect 1187 1486 1188 1490
rect 1182 1485 1188 1486
rect 1214 1490 1220 1491
rect 1214 1486 1215 1490
rect 1219 1486 1220 1490
rect 1214 1485 1220 1486
rect 1254 1490 1260 1491
rect 1254 1486 1255 1490
rect 1259 1486 1260 1490
rect 1254 1485 1260 1486
rect 1294 1490 1300 1491
rect 1294 1486 1295 1490
rect 1299 1486 1300 1490
rect 1294 1485 1300 1486
rect 1350 1490 1356 1491
rect 1350 1486 1351 1490
rect 1355 1486 1356 1490
rect 1350 1485 1356 1486
rect 1414 1490 1420 1491
rect 1414 1486 1415 1490
rect 1419 1486 1420 1490
rect 1414 1485 1420 1486
rect 1486 1490 1492 1491
rect 1486 1486 1487 1490
rect 1491 1486 1492 1490
rect 1486 1485 1492 1486
rect 1566 1490 1572 1491
rect 1566 1486 1567 1490
rect 1571 1486 1572 1490
rect 1566 1485 1572 1486
rect 1622 1490 1628 1491
rect 1622 1486 1623 1490
rect 1627 1486 1628 1490
rect 1622 1485 1628 1486
rect 1662 1488 1668 1489
rect 110 1483 116 1484
rect 112 1475 114 1483
rect 136 1475 138 1485
rect 168 1475 170 1485
rect 224 1475 226 1485
rect 296 1475 298 1485
rect 376 1475 378 1485
rect 456 1475 458 1485
rect 528 1475 530 1485
rect 600 1475 602 1485
rect 672 1475 674 1485
rect 744 1475 746 1485
rect 816 1475 818 1485
rect 880 1475 882 1485
rect 944 1475 946 1485
rect 1008 1475 1010 1485
rect 1064 1475 1066 1485
rect 1112 1475 1114 1485
rect 1152 1475 1154 1485
rect 1184 1475 1186 1485
rect 1216 1475 1218 1485
rect 1256 1475 1258 1485
rect 1296 1475 1298 1485
rect 1352 1475 1354 1485
rect 1416 1475 1418 1485
rect 1488 1475 1490 1485
rect 1568 1475 1570 1485
rect 1624 1475 1626 1485
rect 1662 1484 1663 1488
rect 1667 1484 1668 1488
rect 1662 1483 1668 1484
rect 1664 1475 1666 1483
rect 111 1474 115 1475
rect 111 1469 115 1470
rect 135 1474 139 1475
rect 135 1469 139 1470
rect 167 1474 171 1475
rect 167 1469 171 1470
rect 223 1474 227 1475
rect 223 1469 227 1470
rect 295 1474 299 1475
rect 295 1469 299 1470
rect 375 1474 379 1475
rect 375 1469 379 1470
rect 455 1474 459 1475
rect 455 1469 459 1470
rect 527 1474 531 1475
rect 527 1469 531 1470
rect 599 1474 603 1475
rect 599 1469 603 1470
rect 663 1474 667 1475
rect 663 1469 667 1470
rect 671 1474 675 1475
rect 671 1469 675 1470
rect 719 1474 723 1475
rect 719 1469 723 1470
rect 743 1474 747 1475
rect 743 1469 747 1470
rect 783 1474 787 1475
rect 783 1469 787 1470
rect 815 1474 819 1475
rect 815 1469 819 1470
rect 847 1474 851 1475
rect 847 1469 851 1470
rect 879 1474 883 1475
rect 879 1469 883 1470
rect 903 1474 907 1475
rect 903 1469 907 1470
rect 943 1474 947 1475
rect 943 1469 947 1470
rect 959 1474 963 1475
rect 959 1469 963 1470
rect 1007 1474 1011 1475
rect 1007 1469 1011 1470
rect 1015 1474 1019 1475
rect 1015 1469 1019 1470
rect 1063 1474 1067 1475
rect 1063 1469 1067 1470
rect 1071 1474 1075 1475
rect 1071 1469 1075 1470
rect 1111 1474 1115 1475
rect 1111 1469 1115 1470
rect 1119 1474 1123 1475
rect 1119 1469 1123 1470
rect 1151 1474 1155 1475
rect 1151 1469 1155 1470
rect 1159 1474 1163 1475
rect 1159 1469 1163 1470
rect 1183 1474 1187 1475
rect 1183 1469 1187 1470
rect 1207 1474 1211 1475
rect 1207 1469 1211 1470
rect 1215 1474 1219 1475
rect 1215 1469 1219 1470
rect 1255 1474 1259 1475
rect 1255 1469 1259 1470
rect 1263 1474 1267 1475
rect 1263 1469 1267 1470
rect 1295 1474 1299 1475
rect 1295 1469 1299 1470
rect 1327 1474 1331 1475
rect 1327 1469 1331 1470
rect 1351 1474 1355 1475
rect 1351 1469 1355 1470
rect 1399 1474 1403 1475
rect 1399 1469 1403 1470
rect 1415 1474 1419 1475
rect 1415 1469 1419 1470
rect 1479 1474 1483 1475
rect 1479 1469 1483 1470
rect 1487 1474 1491 1475
rect 1487 1469 1491 1470
rect 1559 1474 1563 1475
rect 1559 1469 1563 1470
rect 1567 1474 1571 1475
rect 1567 1469 1571 1470
rect 1623 1474 1627 1475
rect 1623 1469 1627 1470
rect 1663 1474 1667 1475
rect 1663 1469 1667 1470
rect 112 1461 114 1469
rect 110 1460 116 1461
rect 110 1456 111 1460
rect 115 1456 116 1460
rect 136 1459 138 1469
rect 168 1459 170 1469
rect 224 1459 226 1469
rect 296 1459 298 1469
rect 376 1459 378 1469
rect 456 1459 458 1469
rect 528 1459 530 1469
rect 600 1459 602 1469
rect 664 1459 666 1469
rect 720 1459 722 1469
rect 784 1459 786 1469
rect 848 1459 850 1469
rect 904 1459 906 1469
rect 960 1459 962 1469
rect 1016 1459 1018 1469
rect 1072 1459 1074 1469
rect 1120 1459 1122 1469
rect 1160 1459 1162 1469
rect 1208 1459 1210 1469
rect 1264 1459 1266 1469
rect 1328 1459 1330 1469
rect 1400 1459 1402 1469
rect 1480 1459 1482 1469
rect 1560 1459 1562 1469
rect 1624 1459 1626 1469
rect 1664 1461 1666 1469
rect 1662 1460 1668 1461
rect 110 1455 116 1456
rect 134 1458 140 1459
rect 134 1454 135 1458
rect 139 1454 140 1458
rect 134 1453 140 1454
rect 166 1458 172 1459
rect 166 1454 167 1458
rect 171 1454 172 1458
rect 166 1453 172 1454
rect 222 1458 228 1459
rect 222 1454 223 1458
rect 227 1454 228 1458
rect 222 1453 228 1454
rect 294 1458 300 1459
rect 294 1454 295 1458
rect 299 1454 300 1458
rect 294 1453 300 1454
rect 374 1458 380 1459
rect 374 1454 375 1458
rect 379 1454 380 1458
rect 374 1453 380 1454
rect 454 1458 460 1459
rect 454 1454 455 1458
rect 459 1454 460 1458
rect 454 1453 460 1454
rect 526 1458 532 1459
rect 526 1454 527 1458
rect 531 1454 532 1458
rect 526 1453 532 1454
rect 598 1458 604 1459
rect 598 1454 599 1458
rect 603 1454 604 1458
rect 598 1453 604 1454
rect 662 1458 668 1459
rect 662 1454 663 1458
rect 667 1454 668 1458
rect 662 1453 668 1454
rect 718 1458 724 1459
rect 718 1454 719 1458
rect 723 1454 724 1458
rect 718 1453 724 1454
rect 782 1458 788 1459
rect 782 1454 783 1458
rect 787 1454 788 1458
rect 782 1453 788 1454
rect 846 1458 852 1459
rect 846 1454 847 1458
rect 851 1454 852 1458
rect 846 1453 852 1454
rect 902 1458 908 1459
rect 902 1454 903 1458
rect 907 1454 908 1458
rect 902 1453 908 1454
rect 958 1458 964 1459
rect 958 1454 959 1458
rect 963 1454 964 1458
rect 958 1453 964 1454
rect 1014 1458 1020 1459
rect 1014 1454 1015 1458
rect 1019 1454 1020 1458
rect 1014 1453 1020 1454
rect 1070 1458 1076 1459
rect 1070 1454 1071 1458
rect 1075 1454 1076 1458
rect 1070 1453 1076 1454
rect 1118 1458 1124 1459
rect 1118 1454 1119 1458
rect 1123 1454 1124 1458
rect 1118 1453 1124 1454
rect 1158 1458 1164 1459
rect 1158 1454 1159 1458
rect 1163 1454 1164 1458
rect 1158 1453 1164 1454
rect 1206 1458 1212 1459
rect 1206 1454 1207 1458
rect 1211 1454 1212 1458
rect 1206 1453 1212 1454
rect 1262 1458 1268 1459
rect 1262 1454 1263 1458
rect 1267 1454 1268 1458
rect 1262 1453 1268 1454
rect 1326 1458 1332 1459
rect 1326 1454 1327 1458
rect 1331 1454 1332 1458
rect 1326 1453 1332 1454
rect 1398 1458 1404 1459
rect 1398 1454 1399 1458
rect 1403 1454 1404 1458
rect 1398 1453 1404 1454
rect 1478 1458 1484 1459
rect 1478 1454 1479 1458
rect 1483 1454 1484 1458
rect 1478 1453 1484 1454
rect 1558 1458 1564 1459
rect 1558 1454 1559 1458
rect 1563 1454 1564 1458
rect 1558 1453 1564 1454
rect 1622 1458 1628 1459
rect 1622 1454 1623 1458
rect 1627 1454 1628 1458
rect 1662 1456 1663 1460
rect 1667 1456 1668 1460
rect 1662 1455 1668 1456
rect 1622 1453 1628 1454
rect 110 1443 116 1444
rect 110 1439 111 1443
rect 115 1439 116 1443
rect 1662 1443 1668 1444
rect 110 1438 116 1439
rect 134 1441 140 1442
rect 112 1431 114 1438
rect 134 1437 135 1441
rect 139 1437 140 1441
rect 134 1436 140 1437
rect 166 1441 172 1442
rect 166 1437 167 1441
rect 171 1437 172 1441
rect 166 1436 172 1437
rect 222 1441 228 1442
rect 222 1437 223 1441
rect 227 1437 228 1441
rect 222 1436 228 1437
rect 294 1441 300 1442
rect 294 1437 295 1441
rect 299 1437 300 1441
rect 294 1436 300 1437
rect 374 1441 380 1442
rect 374 1437 375 1441
rect 379 1437 380 1441
rect 374 1436 380 1437
rect 454 1441 460 1442
rect 454 1437 455 1441
rect 459 1437 460 1441
rect 454 1436 460 1437
rect 526 1441 532 1442
rect 526 1437 527 1441
rect 531 1437 532 1441
rect 526 1436 532 1437
rect 598 1441 604 1442
rect 598 1437 599 1441
rect 603 1437 604 1441
rect 598 1436 604 1437
rect 662 1441 668 1442
rect 662 1437 663 1441
rect 667 1437 668 1441
rect 662 1436 668 1437
rect 718 1441 724 1442
rect 718 1437 719 1441
rect 723 1437 724 1441
rect 718 1436 724 1437
rect 782 1441 788 1442
rect 782 1437 783 1441
rect 787 1437 788 1441
rect 782 1436 788 1437
rect 846 1441 852 1442
rect 846 1437 847 1441
rect 851 1437 852 1441
rect 846 1436 852 1437
rect 902 1441 908 1442
rect 902 1437 903 1441
rect 907 1437 908 1441
rect 902 1436 908 1437
rect 958 1441 964 1442
rect 958 1437 959 1441
rect 963 1437 964 1441
rect 958 1436 964 1437
rect 1014 1441 1020 1442
rect 1014 1437 1015 1441
rect 1019 1437 1020 1441
rect 1014 1436 1020 1437
rect 1070 1441 1076 1442
rect 1070 1437 1071 1441
rect 1075 1437 1076 1441
rect 1070 1436 1076 1437
rect 1118 1441 1124 1442
rect 1118 1437 1119 1441
rect 1123 1437 1124 1441
rect 1118 1436 1124 1437
rect 1158 1441 1164 1442
rect 1158 1437 1159 1441
rect 1163 1437 1164 1441
rect 1158 1436 1164 1437
rect 1206 1441 1212 1442
rect 1206 1437 1207 1441
rect 1211 1437 1212 1441
rect 1206 1436 1212 1437
rect 1262 1441 1268 1442
rect 1262 1437 1263 1441
rect 1267 1437 1268 1441
rect 1262 1436 1268 1437
rect 1326 1441 1332 1442
rect 1326 1437 1327 1441
rect 1331 1437 1332 1441
rect 1326 1436 1332 1437
rect 1398 1441 1404 1442
rect 1398 1437 1399 1441
rect 1403 1437 1404 1441
rect 1398 1436 1404 1437
rect 1478 1441 1484 1442
rect 1478 1437 1479 1441
rect 1483 1437 1484 1441
rect 1478 1436 1484 1437
rect 1558 1441 1564 1442
rect 1558 1437 1559 1441
rect 1563 1437 1564 1441
rect 1558 1436 1564 1437
rect 1622 1441 1628 1442
rect 1622 1437 1623 1441
rect 1627 1437 1628 1441
rect 1662 1439 1663 1443
rect 1667 1439 1668 1443
rect 1662 1438 1668 1439
rect 1622 1436 1628 1437
rect 136 1431 138 1436
rect 168 1431 170 1436
rect 224 1431 226 1436
rect 296 1431 298 1436
rect 376 1431 378 1436
rect 456 1431 458 1436
rect 528 1431 530 1436
rect 600 1431 602 1436
rect 664 1431 666 1436
rect 720 1431 722 1436
rect 784 1431 786 1436
rect 848 1431 850 1436
rect 904 1431 906 1436
rect 960 1431 962 1436
rect 1016 1431 1018 1436
rect 1072 1431 1074 1436
rect 1120 1431 1122 1436
rect 1160 1431 1162 1436
rect 1208 1431 1210 1436
rect 1264 1431 1266 1436
rect 1328 1431 1330 1436
rect 1400 1431 1402 1436
rect 1480 1431 1482 1436
rect 1560 1431 1562 1436
rect 1624 1431 1626 1436
rect 1664 1431 1666 1438
rect 111 1430 115 1431
rect 111 1425 115 1426
rect 135 1430 139 1431
rect 112 1422 114 1425
rect 135 1424 139 1426
rect 167 1430 171 1431
rect 167 1424 171 1426
rect 215 1430 219 1431
rect 215 1424 219 1426
rect 223 1430 227 1431
rect 223 1425 227 1426
rect 287 1430 291 1431
rect 287 1424 291 1426
rect 295 1430 299 1431
rect 295 1425 299 1426
rect 359 1430 363 1431
rect 359 1424 363 1426
rect 375 1430 379 1431
rect 375 1425 379 1426
rect 439 1430 443 1431
rect 439 1424 443 1426
rect 455 1430 459 1431
rect 455 1425 459 1426
rect 519 1430 523 1431
rect 519 1424 523 1426
rect 527 1430 531 1431
rect 527 1425 531 1426
rect 599 1430 603 1431
rect 599 1424 603 1426
rect 663 1430 667 1431
rect 663 1425 667 1426
rect 679 1430 683 1431
rect 679 1424 683 1426
rect 719 1430 723 1431
rect 719 1425 723 1426
rect 759 1430 763 1431
rect 759 1424 763 1426
rect 783 1430 787 1431
rect 783 1425 787 1426
rect 831 1430 835 1431
rect 831 1424 835 1426
rect 847 1430 851 1431
rect 847 1425 851 1426
rect 903 1430 907 1431
rect 903 1424 907 1426
rect 959 1430 963 1431
rect 959 1425 963 1426
rect 967 1430 971 1431
rect 967 1424 971 1426
rect 1015 1430 1019 1431
rect 1015 1425 1019 1426
rect 1031 1430 1035 1431
rect 1031 1424 1035 1426
rect 1071 1430 1075 1431
rect 1071 1425 1075 1426
rect 1103 1430 1107 1431
rect 1103 1424 1107 1426
rect 1119 1430 1123 1431
rect 1119 1425 1123 1426
rect 1159 1430 1163 1431
rect 1159 1425 1163 1426
rect 1167 1430 1171 1431
rect 1167 1424 1171 1426
rect 1207 1430 1211 1431
rect 1207 1425 1211 1426
rect 1231 1430 1235 1431
rect 1231 1424 1235 1426
rect 1263 1430 1267 1431
rect 1263 1425 1267 1426
rect 1295 1430 1299 1431
rect 1295 1424 1299 1426
rect 1327 1430 1331 1431
rect 1327 1425 1331 1426
rect 1359 1430 1363 1431
rect 1359 1424 1363 1426
rect 1399 1430 1403 1431
rect 1399 1425 1403 1426
rect 1415 1430 1419 1431
rect 1415 1424 1419 1426
rect 1463 1430 1467 1431
rect 1463 1424 1467 1426
rect 1479 1430 1483 1431
rect 1479 1425 1483 1426
rect 1503 1430 1507 1431
rect 1503 1424 1507 1426
rect 1551 1430 1555 1431
rect 1551 1424 1555 1426
rect 1559 1430 1563 1431
rect 1559 1425 1563 1426
rect 1591 1430 1595 1431
rect 1591 1424 1595 1426
rect 1623 1430 1627 1431
rect 1623 1424 1627 1426
rect 1663 1430 1667 1431
rect 1663 1425 1667 1426
rect 134 1423 140 1424
rect 110 1421 116 1422
rect 110 1417 111 1421
rect 115 1417 116 1421
rect 134 1419 135 1423
rect 139 1419 140 1423
rect 134 1418 140 1419
rect 166 1423 172 1424
rect 166 1419 167 1423
rect 171 1419 172 1423
rect 166 1418 172 1419
rect 214 1423 220 1424
rect 214 1419 215 1423
rect 219 1419 220 1423
rect 214 1418 220 1419
rect 286 1423 292 1424
rect 286 1419 287 1423
rect 291 1419 292 1423
rect 286 1418 292 1419
rect 358 1423 364 1424
rect 358 1419 359 1423
rect 363 1419 364 1423
rect 358 1418 364 1419
rect 438 1423 444 1424
rect 438 1419 439 1423
rect 443 1419 444 1423
rect 438 1418 444 1419
rect 518 1423 524 1424
rect 518 1419 519 1423
rect 523 1419 524 1423
rect 518 1418 524 1419
rect 598 1423 604 1424
rect 598 1419 599 1423
rect 603 1419 604 1423
rect 598 1418 604 1419
rect 678 1423 684 1424
rect 678 1419 679 1423
rect 683 1419 684 1423
rect 678 1418 684 1419
rect 758 1423 764 1424
rect 758 1419 759 1423
rect 763 1419 764 1423
rect 758 1418 764 1419
rect 830 1423 836 1424
rect 830 1419 831 1423
rect 835 1419 836 1423
rect 830 1418 836 1419
rect 902 1423 908 1424
rect 902 1419 903 1423
rect 907 1419 908 1423
rect 902 1418 908 1419
rect 966 1423 972 1424
rect 966 1419 967 1423
rect 971 1419 972 1423
rect 966 1418 972 1419
rect 1030 1423 1036 1424
rect 1030 1419 1031 1423
rect 1035 1419 1036 1423
rect 1030 1418 1036 1419
rect 1102 1423 1108 1424
rect 1102 1419 1103 1423
rect 1107 1419 1108 1423
rect 1102 1418 1108 1419
rect 1166 1423 1172 1424
rect 1166 1419 1167 1423
rect 1171 1419 1172 1423
rect 1166 1418 1172 1419
rect 1230 1423 1236 1424
rect 1230 1419 1231 1423
rect 1235 1419 1236 1423
rect 1230 1418 1236 1419
rect 1294 1423 1300 1424
rect 1294 1419 1295 1423
rect 1299 1419 1300 1423
rect 1294 1418 1300 1419
rect 1358 1423 1364 1424
rect 1358 1419 1359 1423
rect 1363 1419 1364 1423
rect 1358 1418 1364 1419
rect 1414 1423 1420 1424
rect 1414 1419 1415 1423
rect 1419 1419 1420 1423
rect 1414 1418 1420 1419
rect 1462 1423 1468 1424
rect 1462 1419 1463 1423
rect 1467 1419 1468 1423
rect 1462 1418 1468 1419
rect 1502 1423 1508 1424
rect 1502 1419 1503 1423
rect 1507 1419 1508 1423
rect 1502 1418 1508 1419
rect 1550 1423 1556 1424
rect 1550 1419 1551 1423
rect 1555 1419 1556 1423
rect 1550 1418 1556 1419
rect 1590 1423 1596 1424
rect 1590 1419 1591 1423
rect 1595 1419 1596 1423
rect 1590 1418 1596 1419
rect 1622 1423 1628 1424
rect 1622 1419 1623 1423
rect 1627 1419 1628 1423
rect 1664 1422 1666 1425
rect 1622 1418 1628 1419
rect 1662 1421 1668 1422
rect 110 1416 116 1417
rect 1662 1417 1663 1421
rect 1667 1417 1668 1421
rect 1662 1416 1668 1417
rect 134 1406 140 1407
rect 110 1404 116 1405
rect 110 1400 111 1404
rect 115 1400 116 1404
rect 134 1402 135 1406
rect 139 1402 140 1406
rect 134 1401 140 1402
rect 166 1406 172 1407
rect 166 1402 167 1406
rect 171 1402 172 1406
rect 166 1401 172 1402
rect 214 1406 220 1407
rect 214 1402 215 1406
rect 219 1402 220 1406
rect 214 1401 220 1402
rect 286 1406 292 1407
rect 286 1402 287 1406
rect 291 1402 292 1406
rect 286 1401 292 1402
rect 358 1406 364 1407
rect 358 1402 359 1406
rect 363 1402 364 1406
rect 358 1401 364 1402
rect 438 1406 444 1407
rect 438 1402 439 1406
rect 443 1402 444 1406
rect 438 1401 444 1402
rect 518 1406 524 1407
rect 518 1402 519 1406
rect 523 1402 524 1406
rect 518 1401 524 1402
rect 598 1406 604 1407
rect 598 1402 599 1406
rect 603 1402 604 1406
rect 598 1401 604 1402
rect 678 1406 684 1407
rect 678 1402 679 1406
rect 683 1402 684 1406
rect 678 1401 684 1402
rect 758 1406 764 1407
rect 758 1402 759 1406
rect 763 1402 764 1406
rect 758 1401 764 1402
rect 830 1406 836 1407
rect 830 1402 831 1406
rect 835 1402 836 1406
rect 830 1401 836 1402
rect 902 1406 908 1407
rect 902 1402 903 1406
rect 907 1402 908 1406
rect 902 1401 908 1402
rect 966 1406 972 1407
rect 966 1402 967 1406
rect 971 1402 972 1406
rect 966 1401 972 1402
rect 1030 1406 1036 1407
rect 1030 1402 1031 1406
rect 1035 1402 1036 1406
rect 1030 1401 1036 1402
rect 1102 1406 1108 1407
rect 1102 1402 1103 1406
rect 1107 1402 1108 1406
rect 1102 1401 1108 1402
rect 1166 1406 1172 1407
rect 1166 1402 1167 1406
rect 1171 1402 1172 1406
rect 1166 1401 1172 1402
rect 1230 1406 1236 1407
rect 1230 1402 1231 1406
rect 1235 1402 1236 1406
rect 1230 1401 1236 1402
rect 1294 1406 1300 1407
rect 1294 1402 1295 1406
rect 1299 1402 1300 1406
rect 1294 1401 1300 1402
rect 1358 1406 1364 1407
rect 1358 1402 1359 1406
rect 1363 1402 1364 1406
rect 1358 1401 1364 1402
rect 1414 1406 1420 1407
rect 1414 1402 1415 1406
rect 1419 1402 1420 1406
rect 1414 1401 1420 1402
rect 1462 1406 1468 1407
rect 1462 1402 1463 1406
rect 1467 1402 1468 1406
rect 1462 1401 1468 1402
rect 1502 1406 1508 1407
rect 1502 1402 1503 1406
rect 1507 1402 1508 1406
rect 1502 1401 1508 1402
rect 1550 1406 1556 1407
rect 1550 1402 1551 1406
rect 1555 1402 1556 1406
rect 1550 1401 1556 1402
rect 1590 1406 1596 1407
rect 1590 1402 1591 1406
rect 1595 1402 1596 1406
rect 1590 1401 1596 1402
rect 1622 1406 1628 1407
rect 1622 1402 1623 1406
rect 1627 1402 1628 1406
rect 1622 1401 1628 1402
rect 1662 1404 1668 1405
rect 110 1399 116 1400
rect 112 1391 114 1399
rect 136 1391 138 1401
rect 168 1391 170 1401
rect 216 1391 218 1401
rect 288 1391 290 1401
rect 360 1391 362 1401
rect 440 1391 442 1401
rect 520 1391 522 1401
rect 600 1391 602 1401
rect 680 1391 682 1401
rect 760 1391 762 1401
rect 832 1391 834 1401
rect 904 1391 906 1401
rect 968 1391 970 1401
rect 1032 1391 1034 1401
rect 1104 1391 1106 1401
rect 1168 1391 1170 1401
rect 1232 1391 1234 1401
rect 1296 1391 1298 1401
rect 1360 1391 1362 1401
rect 1416 1391 1418 1401
rect 1464 1391 1466 1401
rect 1504 1391 1506 1401
rect 1552 1391 1554 1401
rect 1592 1391 1594 1401
rect 1624 1391 1626 1401
rect 1662 1400 1663 1404
rect 1667 1400 1668 1404
rect 1662 1399 1668 1400
rect 1664 1391 1666 1399
rect 111 1390 115 1391
rect 111 1385 115 1386
rect 135 1390 139 1391
rect 135 1385 139 1386
rect 167 1390 171 1391
rect 167 1385 171 1386
rect 215 1390 219 1391
rect 215 1385 219 1386
rect 223 1390 227 1391
rect 223 1385 227 1386
rect 287 1390 291 1391
rect 287 1385 291 1386
rect 359 1390 363 1391
rect 359 1385 363 1386
rect 431 1390 435 1391
rect 431 1385 435 1386
rect 439 1390 443 1391
rect 439 1385 443 1386
rect 503 1390 507 1391
rect 503 1385 507 1386
rect 519 1390 523 1391
rect 519 1385 523 1386
rect 583 1390 587 1391
rect 583 1385 587 1386
rect 599 1390 603 1391
rect 599 1385 603 1386
rect 663 1390 667 1391
rect 663 1385 667 1386
rect 679 1390 683 1391
rect 679 1385 683 1386
rect 743 1390 747 1391
rect 743 1385 747 1386
rect 759 1390 763 1391
rect 759 1385 763 1386
rect 815 1390 819 1391
rect 815 1385 819 1386
rect 831 1390 835 1391
rect 831 1385 835 1386
rect 887 1390 891 1391
rect 887 1385 891 1386
rect 903 1390 907 1391
rect 903 1385 907 1386
rect 959 1390 963 1391
rect 959 1385 963 1386
rect 967 1390 971 1391
rect 967 1385 971 1386
rect 1031 1390 1035 1391
rect 1031 1385 1035 1386
rect 1103 1390 1107 1391
rect 1103 1385 1107 1386
rect 1167 1390 1171 1391
rect 1167 1385 1171 1386
rect 1175 1390 1179 1391
rect 1175 1385 1179 1386
rect 1231 1390 1235 1391
rect 1231 1385 1235 1386
rect 1239 1390 1243 1391
rect 1239 1385 1243 1386
rect 1295 1390 1299 1391
rect 1295 1385 1299 1386
rect 1303 1390 1307 1391
rect 1303 1385 1307 1386
rect 1359 1390 1363 1391
rect 1359 1385 1363 1386
rect 1367 1390 1371 1391
rect 1367 1385 1371 1386
rect 1415 1390 1419 1391
rect 1415 1385 1419 1386
rect 1431 1390 1435 1391
rect 1431 1385 1435 1386
rect 1463 1390 1467 1391
rect 1463 1385 1467 1386
rect 1495 1390 1499 1391
rect 1495 1385 1499 1386
rect 1503 1390 1507 1391
rect 1503 1385 1507 1386
rect 1551 1390 1555 1391
rect 1551 1385 1555 1386
rect 1567 1390 1571 1391
rect 1567 1385 1571 1386
rect 1591 1390 1595 1391
rect 1591 1385 1595 1386
rect 1623 1390 1627 1391
rect 1623 1385 1627 1386
rect 1663 1390 1667 1391
rect 1663 1385 1667 1386
rect 112 1377 114 1385
rect 110 1376 116 1377
rect 110 1372 111 1376
rect 115 1372 116 1376
rect 136 1375 138 1385
rect 168 1375 170 1385
rect 224 1375 226 1385
rect 288 1375 290 1385
rect 360 1375 362 1385
rect 432 1375 434 1385
rect 504 1375 506 1385
rect 584 1375 586 1385
rect 664 1375 666 1385
rect 744 1375 746 1385
rect 816 1375 818 1385
rect 888 1375 890 1385
rect 960 1375 962 1385
rect 1032 1375 1034 1385
rect 1104 1375 1106 1385
rect 1176 1375 1178 1385
rect 1240 1375 1242 1385
rect 1304 1375 1306 1385
rect 1368 1375 1370 1385
rect 1432 1375 1434 1385
rect 1496 1375 1498 1385
rect 1568 1375 1570 1385
rect 1624 1375 1626 1385
rect 1664 1377 1666 1385
rect 1662 1376 1668 1377
rect 110 1371 116 1372
rect 134 1374 140 1375
rect 134 1370 135 1374
rect 139 1370 140 1374
rect 134 1369 140 1370
rect 166 1374 172 1375
rect 166 1370 167 1374
rect 171 1370 172 1374
rect 166 1369 172 1370
rect 222 1374 228 1375
rect 222 1370 223 1374
rect 227 1370 228 1374
rect 222 1369 228 1370
rect 286 1374 292 1375
rect 286 1370 287 1374
rect 291 1370 292 1374
rect 286 1369 292 1370
rect 358 1374 364 1375
rect 358 1370 359 1374
rect 363 1370 364 1374
rect 358 1369 364 1370
rect 430 1374 436 1375
rect 430 1370 431 1374
rect 435 1370 436 1374
rect 430 1369 436 1370
rect 502 1374 508 1375
rect 502 1370 503 1374
rect 507 1370 508 1374
rect 502 1369 508 1370
rect 582 1374 588 1375
rect 582 1370 583 1374
rect 587 1370 588 1374
rect 582 1369 588 1370
rect 662 1374 668 1375
rect 662 1370 663 1374
rect 667 1370 668 1374
rect 662 1369 668 1370
rect 742 1374 748 1375
rect 742 1370 743 1374
rect 747 1370 748 1374
rect 742 1369 748 1370
rect 814 1374 820 1375
rect 814 1370 815 1374
rect 819 1370 820 1374
rect 814 1369 820 1370
rect 886 1374 892 1375
rect 886 1370 887 1374
rect 891 1370 892 1374
rect 886 1369 892 1370
rect 958 1374 964 1375
rect 958 1370 959 1374
rect 963 1370 964 1374
rect 958 1369 964 1370
rect 1030 1374 1036 1375
rect 1030 1370 1031 1374
rect 1035 1370 1036 1374
rect 1030 1369 1036 1370
rect 1102 1374 1108 1375
rect 1102 1370 1103 1374
rect 1107 1370 1108 1374
rect 1102 1369 1108 1370
rect 1174 1374 1180 1375
rect 1174 1370 1175 1374
rect 1179 1370 1180 1374
rect 1174 1369 1180 1370
rect 1238 1374 1244 1375
rect 1238 1370 1239 1374
rect 1243 1370 1244 1374
rect 1238 1369 1244 1370
rect 1302 1374 1308 1375
rect 1302 1370 1303 1374
rect 1307 1370 1308 1374
rect 1302 1369 1308 1370
rect 1366 1374 1372 1375
rect 1366 1370 1367 1374
rect 1371 1370 1372 1374
rect 1366 1369 1372 1370
rect 1430 1374 1436 1375
rect 1430 1370 1431 1374
rect 1435 1370 1436 1374
rect 1430 1369 1436 1370
rect 1494 1374 1500 1375
rect 1494 1370 1495 1374
rect 1499 1370 1500 1374
rect 1494 1369 1500 1370
rect 1566 1374 1572 1375
rect 1566 1370 1567 1374
rect 1571 1370 1572 1374
rect 1566 1369 1572 1370
rect 1622 1374 1628 1375
rect 1622 1370 1623 1374
rect 1627 1370 1628 1374
rect 1662 1372 1663 1376
rect 1667 1372 1668 1376
rect 1662 1371 1668 1372
rect 1622 1369 1628 1370
rect 110 1359 116 1360
rect 110 1355 111 1359
rect 115 1355 116 1359
rect 1662 1359 1668 1360
rect 110 1354 116 1355
rect 134 1357 140 1358
rect 112 1351 114 1354
rect 134 1353 135 1357
rect 139 1353 140 1357
rect 134 1352 140 1353
rect 166 1357 172 1358
rect 166 1353 167 1357
rect 171 1353 172 1357
rect 166 1352 172 1353
rect 222 1357 228 1358
rect 222 1353 223 1357
rect 227 1353 228 1357
rect 222 1352 228 1353
rect 286 1357 292 1358
rect 286 1353 287 1357
rect 291 1353 292 1357
rect 286 1352 292 1353
rect 358 1357 364 1358
rect 358 1353 359 1357
rect 363 1353 364 1357
rect 358 1352 364 1353
rect 430 1357 436 1358
rect 430 1353 431 1357
rect 435 1353 436 1357
rect 430 1352 436 1353
rect 502 1357 508 1358
rect 502 1353 503 1357
rect 507 1353 508 1357
rect 502 1352 508 1353
rect 582 1357 588 1358
rect 582 1353 583 1357
rect 587 1353 588 1357
rect 582 1352 588 1353
rect 662 1357 668 1358
rect 662 1353 663 1357
rect 667 1353 668 1357
rect 662 1352 668 1353
rect 742 1357 748 1358
rect 742 1353 743 1357
rect 747 1353 748 1357
rect 742 1352 748 1353
rect 814 1357 820 1358
rect 814 1353 815 1357
rect 819 1353 820 1357
rect 814 1352 820 1353
rect 886 1357 892 1358
rect 886 1353 887 1357
rect 891 1353 892 1357
rect 886 1352 892 1353
rect 958 1357 964 1358
rect 958 1353 959 1357
rect 963 1353 964 1357
rect 958 1352 964 1353
rect 1030 1357 1036 1358
rect 1030 1353 1031 1357
rect 1035 1353 1036 1357
rect 1030 1352 1036 1353
rect 1102 1357 1108 1358
rect 1102 1353 1103 1357
rect 1107 1353 1108 1357
rect 1102 1352 1108 1353
rect 1174 1357 1180 1358
rect 1174 1353 1175 1357
rect 1179 1353 1180 1357
rect 1174 1352 1180 1353
rect 1238 1357 1244 1358
rect 1238 1353 1239 1357
rect 1243 1353 1244 1357
rect 1238 1352 1244 1353
rect 1302 1357 1308 1358
rect 1302 1353 1303 1357
rect 1307 1353 1308 1357
rect 1302 1352 1308 1353
rect 1366 1357 1372 1358
rect 1366 1353 1367 1357
rect 1371 1353 1372 1357
rect 1366 1352 1372 1353
rect 1430 1357 1436 1358
rect 1430 1353 1431 1357
rect 1435 1353 1436 1357
rect 1430 1352 1436 1353
rect 1494 1357 1500 1358
rect 1494 1353 1495 1357
rect 1499 1353 1500 1357
rect 1494 1352 1500 1353
rect 1566 1357 1572 1358
rect 1566 1353 1567 1357
rect 1571 1353 1572 1357
rect 1566 1352 1572 1353
rect 1622 1357 1628 1358
rect 1622 1353 1623 1357
rect 1627 1353 1628 1357
rect 1662 1355 1663 1359
rect 1667 1355 1668 1359
rect 1662 1354 1668 1355
rect 1622 1352 1628 1353
rect 111 1350 115 1351
rect 111 1345 115 1346
rect 135 1350 139 1352
rect 112 1342 114 1345
rect 135 1344 139 1346
rect 167 1350 171 1352
rect 167 1345 171 1346
rect 183 1350 187 1351
rect 183 1344 187 1346
rect 223 1350 227 1352
rect 223 1345 227 1346
rect 239 1350 243 1351
rect 239 1344 243 1346
rect 287 1350 291 1352
rect 287 1345 291 1346
rect 295 1350 299 1351
rect 295 1344 299 1346
rect 351 1350 355 1351
rect 351 1344 355 1346
rect 359 1350 363 1352
rect 359 1345 363 1346
rect 399 1350 403 1351
rect 399 1344 403 1346
rect 431 1350 435 1352
rect 431 1345 435 1346
rect 455 1350 459 1351
rect 455 1344 459 1346
rect 503 1350 507 1352
rect 503 1345 507 1346
rect 511 1350 515 1351
rect 511 1344 515 1346
rect 567 1350 571 1351
rect 567 1344 571 1346
rect 583 1350 587 1352
rect 583 1345 587 1346
rect 631 1350 635 1351
rect 631 1344 635 1346
rect 663 1350 667 1352
rect 663 1345 667 1346
rect 695 1350 699 1351
rect 695 1344 699 1346
rect 743 1350 747 1352
rect 743 1345 747 1346
rect 759 1350 763 1351
rect 759 1344 763 1346
rect 815 1350 819 1352
rect 815 1345 819 1346
rect 823 1350 827 1351
rect 823 1344 827 1346
rect 887 1350 891 1352
rect 887 1344 891 1346
rect 959 1350 963 1352
rect 959 1344 963 1346
rect 1023 1350 1027 1351
rect 1023 1344 1027 1346
rect 1031 1350 1035 1352
rect 1031 1345 1035 1346
rect 1087 1350 1091 1351
rect 1087 1344 1091 1346
rect 1103 1350 1107 1352
rect 1103 1345 1107 1346
rect 1151 1350 1155 1351
rect 1151 1344 1155 1346
rect 1175 1350 1179 1352
rect 1175 1345 1179 1346
rect 1215 1350 1219 1351
rect 1215 1344 1219 1346
rect 1239 1350 1243 1352
rect 1239 1345 1243 1346
rect 1279 1350 1283 1351
rect 1279 1344 1283 1346
rect 1303 1350 1307 1352
rect 1303 1345 1307 1346
rect 1343 1350 1347 1351
rect 1343 1344 1347 1346
rect 1367 1350 1371 1352
rect 1367 1345 1371 1346
rect 1407 1350 1411 1351
rect 1407 1344 1411 1346
rect 1431 1350 1435 1352
rect 1431 1345 1435 1346
rect 1479 1350 1483 1351
rect 1479 1344 1483 1346
rect 1495 1350 1499 1352
rect 1495 1345 1499 1346
rect 1559 1350 1563 1351
rect 1559 1344 1563 1346
rect 1567 1350 1571 1352
rect 1567 1345 1571 1346
rect 1623 1350 1627 1352
rect 1664 1351 1666 1354
rect 1623 1344 1627 1346
rect 1663 1350 1667 1351
rect 1663 1345 1667 1346
rect 134 1343 140 1344
rect 110 1341 116 1342
rect 110 1337 111 1341
rect 115 1337 116 1341
rect 134 1339 135 1343
rect 139 1339 140 1343
rect 134 1338 140 1339
rect 182 1343 188 1344
rect 182 1339 183 1343
rect 187 1339 188 1343
rect 182 1338 188 1339
rect 238 1343 244 1344
rect 238 1339 239 1343
rect 243 1339 244 1343
rect 238 1338 244 1339
rect 294 1343 300 1344
rect 294 1339 295 1343
rect 299 1339 300 1343
rect 294 1338 300 1339
rect 350 1343 356 1344
rect 350 1339 351 1343
rect 355 1339 356 1343
rect 350 1338 356 1339
rect 398 1343 404 1344
rect 398 1339 399 1343
rect 403 1339 404 1343
rect 398 1338 404 1339
rect 454 1343 460 1344
rect 454 1339 455 1343
rect 459 1339 460 1343
rect 454 1338 460 1339
rect 510 1343 516 1344
rect 510 1339 511 1343
rect 515 1339 516 1343
rect 510 1338 516 1339
rect 566 1343 572 1344
rect 566 1339 567 1343
rect 571 1339 572 1343
rect 566 1338 572 1339
rect 630 1343 636 1344
rect 630 1339 631 1343
rect 635 1339 636 1343
rect 630 1338 636 1339
rect 694 1343 700 1344
rect 694 1339 695 1343
rect 699 1339 700 1343
rect 694 1338 700 1339
rect 758 1343 764 1344
rect 758 1339 759 1343
rect 763 1339 764 1343
rect 758 1338 764 1339
rect 822 1343 828 1344
rect 822 1339 823 1343
rect 827 1339 828 1343
rect 822 1338 828 1339
rect 886 1343 892 1344
rect 886 1339 887 1343
rect 891 1339 892 1343
rect 886 1338 892 1339
rect 958 1343 964 1344
rect 958 1339 959 1343
rect 963 1339 964 1343
rect 958 1338 964 1339
rect 1022 1343 1028 1344
rect 1022 1339 1023 1343
rect 1027 1339 1028 1343
rect 1022 1338 1028 1339
rect 1086 1343 1092 1344
rect 1086 1339 1087 1343
rect 1091 1339 1092 1343
rect 1086 1338 1092 1339
rect 1150 1343 1156 1344
rect 1150 1339 1151 1343
rect 1155 1339 1156 1343
rect 1150 1338 1156 1339
rect 1214 1343 1220 1344
rect 1214 1339 1215 1343
rect 1219 1339 1220 1343
rect 1214 1338 1220 1339
rect 1278 1343 1284 1344
rect 1278 1339 1279 1343
rect 1283 1339 1284 1343
rect 1278 1338 1284 1339
rect 1342 1343 1348 1344
rect 1342 1339 1343 1343
rect 1347 1339 1348 1343
rect 1342 1338 1348 1339
rect 1406 1343 1412 1344
rect 1406 1339 1407 1343
rect 1411 1339 1412 1343
rect 1406 1338 1412 1339
rect 1478 1343 1484 1344
rect 1478 1339 1479 1343
rect 1483 1339 1484 1343
rect 1478 1338 1484 1339
rect 1558 1343 1564 1344
rect 1558 1339 1559 1343
rect 1563 1339 1564 1343
rect 1558 1338 1564 1339
rect 1622 1343 1628 1344
rect 1622 1339 1623 1343
rect 1627 1339 1628 1343
rect 1664 1342 1666 1345
rect 1622 1338 1628 1339
rect 1662 1341 1668 1342
rect 110 1336 116 1337
rect 1662 1337 1663 1341
rect 1667 1337 1668 1341
rect 1662 1336 1668 1337
rect 134 1326 140 1327
rect 110 1324 116 1325
rect 110 1320 111 1324
rect 115 1320 116 1324
rect 134 1322 135 1326
rect 139 1322 140 1326
rect 134 1321 140 1322
rect 182 1326 188 1327
rect 182 1322 183 1326
rect 187 1322 188 1326
rect 182 1321 188 1322
rect 238 1326 244 1327
rect 238 1322 239 1326
rect 243 1322 244 1326
rect 238 1321 244 1322
rect 294 1326 300 1327
rect 294 1322 295 1326
rect 299 1322 300 1326
rect 294 1321 300 1322
rect 350 1326 356 1327
rect 350 1322 351 1326
rect 355 1322 356 1326
rect 350 1321 356 1322
rect 398 1326 404 1327
rect 398 1322 399 1326
rect 403 1322 404 1326
rect 398 1321 404 1322
rect 454 1326 460 1327
rect 454 1322 455 1326
rect 459 1322 460 1326
rect 454 1321 460 1322
rect 510 1326 516 1327
rect 510 1322 511 1326
rect 515 1322 516 1326
rect 510 1321 516 1322
rect 566 1326 572 1327
rect 566 1322 567 1326
rect 571 1322 572 1326
rect 566 1321 572 1322
rect 630 1326 636 1327
rect 630 1322 631 1326
rect 635 1322 636 1326
rect 630 1321 636 1322
rect 694 1326 700 1327
rect 694 1322 695 1326
rect 699 1322 700 1326
rect 694 1321 700 1322
rect 758 1326 764 1327
rect 758 1322 759 1326
rect 763 1322 764 1326
rect 758 1321 764 1322
rect 822 1326 828 1327
rect 822 1322 823 1326
rect 827 1322 828 1326
rect 822 1321 828 1322
rect 886 1326 892 1327
rect 886 1322 887 1326
rect 891 1322 892 1326
rect 886 1321 892 1322
rect 958 1326 964 1327
rect 958 1322 959 1326
rect 963 1322 964 1326
rect 958 1321 964 1322
rect 1022 1326 1028 1327
rect 1022 1322 1023 1326
rect 1027 1322 1028 1326
rect 1022 1321 1028 1322
rect 1086 1326 1092 1327
rect 1086 1322 1087 1326
rect 1091 1322 1092 1326
rect 1086 1321 1092 1322
rect 1150 1326 1156 1327
rect 1150 1322 1151 1326
rect 1155 1322 1156 1326
rect 1150 1321 1156 1322
rect 1214 1326 1220 1327
rect 1214 1322 1215 1326
rect 1219 1322 1220 1326
rect 1214 1321 1220 1322
rect 1278 1326 1284 1327
rect 1278 1322 1279 1326
rect 1283 1322 1284 1326
rect 1278 1321 1284 1322
rect 1342 1326 1348 1327
rect 1342 1322 1343 1326
rect 1347 1322 1348 1326
rect 1342 1321 1348 1322
rect 1406 1326 1412 1327
rect 1406 1322 1407 1326
rect 1411 1322 1412 1326
rect 1406 1321 1412 1322
rect 1478 1326 1484 1327
rect 1478 1322 1479 1326
rect 1483 1322 1484 1326
rect 1478 1321 1484 1322
rect 1558 1326 1564 1327
rect 1558 1322 1559 1326
rect 1563 1322 1564 1326
rect 1558 1321 1564 1322
rect 1622 1326 1628 1327
rect 1622 1322 1623 1326
rect 1627 1322 1628 1326
rect 1622 1321 1628 1322
rect 1662 1324 1668 1325
rect 110 1319 116 1320
rect 112 1307 114 1319
rect 136 1307 138 1321
rect 184 1307 186 1321
rect 240 1307 242 1321
rect 296 1307 298 1321
rect 352 1307 354 1321
rect 400 1307 402 1321
rect 456 1307 458 1321
rect 512 1307 514 1321
rect 568 1307 570 1321
rect 632 1307 634 1321
rect 696 1307 698 1321
rect 760 1307 762 1321
rect 824 1307 826 1321
rect 888 1307 890 1321
rect 960 1307 962 1321
rect 1024 1307 1026 1321
rect 1088 1307 1090 1321
rect 1152 1307 1154 1321
rect 1216 1307 1218 1321
rect 1280 1307 1282 1321
rect 1344 1307 1346 1321
rect 1408 1307 1410 1321
rect 1480 1307 1482 1321
rect 1560 1307 1562 1321
rect 1624 1307 1626 1321
rect 1662 1320 1663 1324
rect 1667 1320 1668 1324
rect 1662 1319 1668 1320
rect 1664 1307 1666 1319
rect 111 1306 115 1307
rect 111 1301 115 1302
rect 135 1306 139 1307
rect 135 1301 139 1302
rect 183 1306 187 1307
rect 183 1301 187 1302
rect 231 1306 235 1307
rect 231 1301 235 1302
rect 239 1306 243 1307
rect 239 1301 243 1302
rect 279 1306 283 1307
rect 279 1301 283 1302
rect 295 1306 299 1307
rect 295 1301 299 1302
rect 327 1306 331 1307
rect 327 1301 331 1302
rect 351 1306 355 1307
rect 351 1301 355 1302
rect 375 1306 379 1307
rect 375 1301 379 1302
rect 399 1306 403 1307
rect 399 1301 403 1302
rect 431 1306 435 1307
rect 431 1301 435 1302
rect 455 1306 459 1307
rect 455 1301 459 1302
rect 487 1306 491 1307
rect 487 1301 491 1302
rect 511 1306 515 1307
rect 511 1301 515 1302
rect 543 1306 547 1307
rect 543 1301 547 1302
rect 567 1306 571 1307
rect 567 1301 571 1302
rect 607 1306 611 1307
rect 607 1301 611 1302
rect 631 1306 635 1307
rect 631 1301 635 1302
rect 663 1306 667 1307
rect 663 1301 667 1302
rect 695 1306 699 1307
rect 695 1301 699 1302
rect 719 1306 723 1307
rect 719 1301 723 1302
rect 759 1306 763 1307
rect 759 1301 763 1302
rect 775 1306 779 1307
rect 775 1301 779 1302
rect 823 1306 827 1307
rect 823 1301 827 1302
rect 831 1306 835 1307
rect 831 1301 835 1302
rect 887 1306 891 1307
rect 887 1301 891 1302
rect 895 1306 899 1307
rect 895 1301 899 1302
rect 959 1306 963 1307
rect 959 1301 963 1302
rect 1023 1306 1027 1307
rect 1023 1301 1027 1302
rect 1079 1306 1083 1307
rect 1079 1301 1083 1302
rect 1087 1306 1091 1307
rect 1087 1301 1091 1302
rect 1143 1306 1147 1307
rect 1143 1301 1147 1302
rect 1151 1306 1155 1307
rect 1151 1301 1155 1302
rect 1207 1306 1211 1307
rect 1207 1301 1211 1302
rect 1215 1306 1219 1307
rect 1215 1301 1219 1302
rect 1279 1306 1283 1307
rect 1279 1301 1283 1302
rect 1343 1306 1347 1307
rect 1343 1301 1347 1302
rect 1359 1306 1363 1307
rect 1359 1301 1363 1302
rect 1407 1306 1411 1307
rect 1407 1301 1411 1302
rect 1447 1306 1451 1307
rect 1447 1301 1451 1302
rect 1479 1306 1483 1307
rect 1479 1301 1483 1302
rect 1543 1306 1547 1307
rect 1543 1301 1547 1302
rect 1559 1306 1563 1307
rect 1559 1301 1563 1302
rect 1623 1306 1627 1307
rect 1623 1301 1627 1302
rect 1663 1306 1667 1307
rect 1663 1301 1667 1302
rect 112 1293 114 1301
rect 110 1292 116 1293
rect 110 1288 111 1292
rect 115 1288 116 1292
rect 136 1291 138 1301
rect 184 1291 186 1301
rect 232 1291 234 1301
rect 280 1291 282 1301
rect 328 1291 330 1301
rect 376 1291 378 1301
rect 432 1291 434 1301
rect 488 1291 490 1301
rect 544 1291 546 1301
rect 608 1291 610 1301
rect 664 1291 666 1301
rect 720 1291 722 1301
rect 776 1291 778 1301
rect 832 1291 834 1301
rect 896 1291 898 1301
rect 960 1291 962 1301
rect 1024 1291 1026 1301
rect 1080 1291 1082 1301
rect 1144 1291 1146 1301
rect 1208 1291 1210 1301
rect 1280 1291 1282 1301
rect 1360 1291 1362 1301
rect 1448 1291 1450 1301
rect 1544 1291 1546 1301
rect 1624 1291 1626 1301
rect 1664 1293 1666 1301
rect 1662 1292 1668 1293
rect 110 1287 116 1288
rect 134 1290 140 1291
rect 134 1286 135 1290
rect 139 1286 140 1290
rect 134 1285 140 1286
rect 182 1290 188 1291
rect 182 1286 183 1290
rect 187 1286 188 1290
rect 182 1285 188 1286
rect 230 1290 236 1291
rect 230 1286 231 1290
rect 235 1286 236 1290
rect 230 1285 236 1286
rect 278 1290 284 1291
rect 278 1286 279 1290
rect 283 1286 284 1290
rect 278 1285 284 1286
rect 326 1290 332 1291
rect 326 1286 327 1290
rect 331 1286 332 1290
rect 326 1285 332 1286
rect 374 1290 380 1291
rect 374 1286 375 1290
rect 379 1286 380 1290
rect 374 1285 380 1286
rect 430 1290 436 1291
rect 430 1286 431 1290
rect 435 1286 436 1290
rect 430 1285 436 1286
rect 486 1290 492 1291
rect 486 1286 487 1290
rect 491 1286 492 1290
rect 486 1285 492 1286
rect 542 1290 548 1291
rect 542 1286 543 1290
rect 547 1286 548 1290
rect 542 1285 548 1286
rect 606 1290 612 1291
rect 606 1286 607 1290
rect 611 1286 612 1290
rect 606 1285 612 1286
rect 662 1290 668 1291
rect 662 1286 663 1290
rect 667 1286 668 1290
rect 662 1285 668 1286
rect 718 1290 724 1291
rect 718 1286 719 1290
rect 723 1286 724 1290
rect 718 1285 724 1286
rect 774 1290 780 1291
rect 774 1286 775 1290
rect 779 1286 780 1290
rect 774 1285 780 1286
rect 830 1290 836 1291
rect 830 1286 831 1290
rect 835 1286 836 1290
rect 830 1285 836 1286
rect 894 1290 900 1291
rect 894 1286 895 1290
rect 899 1286 900 1290
rect 894 1285 900 1286
rect 958 1290 964 1291
rect 958 1286 959 1290
rect 963 1286 964 1290
rect 958 1285 964 1286
rect 1022 1290 1028 1291
rect 1022 1286 1023 1290
rect 1027 1286 1028 1290
rect 1022 1285 1028 1286
rect 1078 1290 1084 1291
rect 1078 1286 1079 1290
rect 1083 1286 1084 1290
rect 1078 1285 1084 1286
rect 1142 1290 1148 1291
rect 1142 1286 1143 1290
rect 1147 1286 1148 1290
rect 1142 1285 1148 1286
rect 1206 1290 1212 1291
rect 1206 1286 1207 1290
rect 1211 1286 1212 1290
rect 1206 1285 1212 1286
rect 1278 1290 1284 1291
rect 1278 1286 1279 1290
rect 1283 1286 1284 1290
rect 1278 1285 1284 1286
rect 1358 1290 1364 1291
rect 1358 1286 1359 1290
rect 1363 1286 1364 1290
rect 1358 1285 1364 1286
rect 1446 1290 1452 1291
rect 1446 1286 1447 1290
rect 1451 1286 1452 1290
rect 1446 1285 1452 1286
rect 1542 1290 1548 1291
rect 1542 1286 1543 1290
rect 1547 1286 1548 1290
rect 1542 1285 1548 1286
rect 1622 1290 1628 1291
rect 1622 1286 1623 1290
rect 1627 1286 1628 1290
rect 1662 1288 1663 1292
rect 1667 1288 1668 1292
rect 1662 1287 1668 1288
rect 1622 1285 1628 1286
rect 110 1275 116 1276
rect 110 1271 111 1275
rect 115 1271 116 1275
rect 1662 1275 1668 1276
rect 110 1270 116 1271
rect 134 1273 140 1274
rect 112 1267 114 1270
rect 134 1269 135 1273
rect 139 1269 140 1273
rect 134 1268 140 1269
rect 182 1273 188 1274
rect 182 1269 183 1273
rect 187 1269 188 1273
rect 182 1268 188 1269
rect 230 1273 236 1274
rect 230 1269 231 1273
rect 235 1269 236 1273
rect 230 1268 236 1269
rect 278 1273 284 1274
rect 278 1269 279 1273
rect 283 1269 284 1273
rect 278 1268 284 1269
rect 326 1273 332 1274
rect 326 1269 327 1273
rect 331 1269 332 1273
rect 326 1268 332 1269
rect 374 1273 380 1274
rect 374 1269 375 1273
rect 379 1269 380 1273
rect 374 1268 380 1269
rect 430 1273 436 1274
rect 430 1269 431 1273
rect 435 1269 436 1273
rect 430 1268 436 1269
rect 486 1273 492 1274
rect 486 1269 487 1273
rect 491 1269 492 1273
rect 486 1268 492 1269
rect 542 1273 548 1274
rect 542 1269 543 1273
rect 547 1269 548 1273
rect 542 1268 548 1269
rect 606 1273 612 1274
rect 606 1269 607 1273
rect 611 1269 612 1273
rect 606 1268 612 1269
rect 662 1273 668 1274
rect 662 1269 663 1273
rect 667 1269 668 1273
rect 662 1268 668 1269
rect 718 1273 724 1274
rect 718 1269 719 1273
rect 723 1269 724 1273
rect 718 1268 724 1269
rect 774 1273 780 1274
rect 774 1269 775 1273
rect 779 1269 780 1273
rect 774 1268 780 1269
rect 830 1273 836 1274
rect 830 1269 831 1273
rect 835 1269 836 1273
rect 830 1268 836 1269
rect 894 1273 900 1274
rect 894 1269 895 1273
rect 899 1269 900 1273
rect 894 1268 900 1269
rect 958 1273 964 1274
rect 958 1269 959 1273
rect 963 1269 964 1273
rect 958 1268 964 1269
rect 1022 1273 1028 1274
rect 1022 1269 1023 1273
rect 1027 1269 1028 1273
rect 1022 1268 1028 1269
rect 1078 1273 1084 1274
rect 1078 1269 1079 1273
rect 1083 1269 1084 1273
rect 1078 1268 1084 1269
rect 1142 1273 1148 1274
rect 1142 1269 1143 1273
rect 1147 1269 1148 1273
rect 1142 1268 1148 1269
rect 1206 1273 1212 1274
rect 1206 1269 1207 1273
rect 1211 1269 1212 1273
rect 1206 1268 1212 1269
rect 1278 1273 1284 1274
rect 1278 1269 1279 1273
rect 1283 1269 1284 1273
rect 1278 1268 1284 1269
rect 1358 1273 1364 1274
rect 1358 1269 1359 1273
rect 1363 1269 1364 1273
rect 1358 1268 1364 1269
rect 1446 1273 1452 1274
rect 1446 1269 1447 1273
rect 1451 1269 1452 1273
rect 1446 1268 1452 1269
rect 1542 1273 1548 1274
rect 1542 1269 1543 1273
rect 1547 1269 1548 1273
rect 1542 1268 1548 1269
rect 1622 1273 1628 1274
rect 1622 1269 1623 1273
rect 1627 1269 1628 1273
rect 1662 1271 1663 1275
rect 1667 1271 1668 1275
rect 1662 1270 1668 1271
rect 1622 1268 1628 1269
rect 111 1266 115 1267
rect 111 1261 115 1262
rect 135 1266 139 1268
rect 112 1258 114 1261
rect 135 1260 139 1262
rect 167 1266 171 1267
rect 167 1260 171 1262
rect 183 1266 187 1268
rect 183 1261 187 1262
rect 223 1266 227 1267
rect 223 1260 227 1262
rect 231 1266 235 1268
rect 231 1261 235 1262
rect 279 1266 283 1268
rect 279 1260 283 1262
rect 327 1266 331 1268
rect 327 1260 331 1262
rect 375 1266 379 1268
rect 375 1261 379 1262
rect 383 1266 387 1267
rect 383 1260 387 1262
rect 431 1266 435 1268
rect 431 1261 435 1262
rect 439 1266 443 1267
rect 439 1260 443 1262
rect 487 1266 491 1268
rect 487 1261 491 1262
rect 495 1266 499 1267
rect 495 1260 499 1262
rect 543 1266 547 1268
rect 543 1261 547 1262
rect 551 1266 555 1267
rect 551 1260 555 1262
rect 607 1266 611 1268
rect 607 1260 611 1262
rect 663 1266 667 1268
rect 663 1260 667 1262
rect 719 1266 723 1268
rect 719 1260 723 1262
rect 767 1266 771 1267
rect 767 1260 771 1262
rect 775 1266 779 1268
rect 775 1261 779 1262
rect 815 1266 819 1267
rect 815 1260 819 1262
rect 831 1266 835 1268
rect 831 1261 835 1262
rect 871 1266 875 1267
rect 871 1260 875 1262
rect 895 1266 899 1268
rect 895 1261 899 1262
rect 927 1266 931 1267
rect 927 1260 931 1262
rect 959 1266 963 1268
rect 959 1261 963 1262
rect 983 1266 987 1267
rect 983 1260 987 1262
rect 1023 1266 1027 1268
rect 1023 1261 1027 1262
rect 1039 1266 1043 1267
rect 1039 1260 1043 1262
rect 1079 1266 1083 1268
rect 1079 1261 1083 1262
rect 1095 1266 1099 1267
rect 1095 1260 1099 1262
rect 1143 1266 1147 1268
rect 1143 1261 1147 1262
rect 1159 1266 1163 1267
rect 1159 1260 1163 1262
rect 1207 1266 1211 1268
rect 1207 1261 1211 1262
rect 1231 1266 1235 1267
rect 1231 1260 1235 1262
rect 1279 1266 1283 1268
rect 1279 1261 1283 1262
rect 1319 1266 1323 1267
rect 1319 1260 1323 1262
rect 1359 1266 1363 1268
rect 1359 1261 1363 1262
rect 1423 1266 1427 1267
rect 1423 1260 1427 1262
rect 1447 1266 1451 1268
rect 1447 1261 1451 1262
rect 1535 1266 1539 1267
rect 1535 1260 1539 1262
rect 1543 1266 1547 1268
rect 1543 1261 1547 1262
rect 1623 1266 1627 1268
rect 1664 1267 1666 1270
rect 1623 1260 1627 1262
rect 1663 1266 1667 1267
rect 1663 1261 1667 1262
rect 134 1259 140 1260
rect 110 1257 116 1258
rect 110 1253 111 1257
rect 115 1253 116 1257
rect 134 1255 135 1259
rect 139 1255 140 1259
rect 134 1254 140 1255
rect 166 1259 172 1260
rect 166 1255 167 1259
rect 171 1255 172 1259
rect 166 1254 172 1255
rect 222 1259 228 1260
rect 222 1255 223 1259
rect 227 1255 228 1259
rect 222 1254 228 1255
rect 278 1259 284 1260
rect 278 1255 279 1259
rect 283 1255 284 1259
rect 278 1254 284 1255
rect 326 1259 332 1260
rect 326 1255 327 1259
rect 331 1255 332 1259
rect 326 1254 332 1255
rect 382 1259 388 1260
rect 382 1255 383 1259
rect 387 1255 388 1259
rect 382 1254 388 1255
rect 438 1259 444 1260
rect 438 1255 439 1259
rect 443 1255 444 1259
rect 438 1254 444 1255
rect 494 1259 500 1260
rect 494 1255 495 1259
rect 499 1255 500 1259
rect 494 1254 500 1255
rect 550 1259 556 1260
rect 550 1255 551 1259
rect 555 1255 556 1259
rect 550 1254 556 1255
rect 606 1259 612 1260
rect 606 1255 607 1259
rect 611 1255 612 1259
rect 606 1254 612 1255
rect 662 1259 668 1260
rect 662 1255 663 1259
rect 667 1255 668 1259
rect 662 1254 668 1255
rect 718 1259 724 1260
rect 718 1255 719 1259
rect 723 1255 724 1259
rect 718 1254 724 1255
rect 766 1259 772 1260
rect 766 1255 767 1259
rect 771 1255 772 1259
rect 766 1254 772 1255
rect 814 1259 820 1260
rect 814 1255 815 1259
rect 819 1255 820 1259
rect 814 1254 820 1255
rect 870 1259 876 1260
rect 870 1255 871 1259
rect 875 1255 876 1259
rect 870 1254 876 1255
rect 926 1259 932 1260
rect 926 1255 927 1259
rect 931 1255 932 1259
rect 926 1254 932 1255
rect 982 1259 988 1260
rect 982 1255 983 1259
rect 987 1255 988 1259
rect 982 1254 988 1255
rect 1038 1259 1044 1260
rect 1038 1255 1039 1259
rect 1043 1255 1044 1259
rect 1038 1254 1044 1255
rect 1094 1259 1100 1260
rect 1094 1255 1095 1259
rect 1099 1255 1100 1259
rect 1094 1254 1100 1255
rect 1158 1259 1164 1260
rect 1158 1255 1159 1259
rect 1163 1255 1164 1259
rect 1158 1254 1164 1255
rect 1230 1259 1236 1260
rect 1230 1255 1231 1259
rect 1235 1255 1236 1259
rect 1230 1254 1236 1255
rect 1318 1259 1324 1260
rect 1318 1255 1319 1259
rect 1323 1255 1324 1259
rect 1318 1254 1324 1255
rect 1422 1259 1428 1260
rect 1422 1255 1423 1259
rect 1427 1255 1428 1259
rect 1422 1254 1428 1255
rect 1534 1259 1540 1260
rect 1534 1255 1535 1259
rect 1539 1255 1540 1259
rect 1534 1254 1540 1255
rect 1622 1259 1628 1260
rect 1622 1255 1623 1259
rect 1627 1255 1628 1259
rect 1664 1258 1666 1261
rect 1622 1254 1628 1255
rect 1662 1257 1668 1258
rect 110 1252 116 1253
rect 1662 1253 1663 1257
rect 1667 1253 1668 1257
rect 1662 1252 1668 1253
rect 134 1242 140 1243
rect 110 1240 116 1241
rect 110 1236 111 1240
rect 115 1236 116 1240
rect 134 1238 135 1242
rect 139 1238 140 1242
rect 134 1237 140 1238
rect 166 1242 172 1243
rect 166 1238 167 1242
rect 171 1238 172 1242
rect 166 1237 172 1238
rect 222 1242 228 1243
rect 222 1238 223 1242
rect 227 1238 228 1242
rect 222 1237 228 1238
rect 278 1242 284 1243
rect 278 1238 279 1242
rect 283 1238 284 1242
rect 278 1237 284 1238
rect 326 1242 332 1243
rect 326 1238 327 1242
rect 331 1238 332 1242
rect 326 1237 332 1238
rect 382 1242 388 1243
rect 382 1238 383 1242
rect 387 1238 388 1242
rect 382 1237 388 1238
rect 438 1242 444 1243
rect 438 1238 439 1242
rect 443 1238 444 1242
rect 438 1237 444 1238
rect 494 1242 500 1243
rect 494 1238 495 1242
rect 499 1238 500 1242
rect 494 1237 500 1238
rect 550 1242 556 1243
rect 550 1238 551 1242
rect 555 1238 556 1242
rect 550 1237 556 1238
rect 606 1242 612 1243
rect 606 1238 607 1242
rect 611 1238 612 1242
rect 606 1237 612 1238
rect 662 1242 668 1243
rect 662 1238 663 1242
rect 667 1238 668 1242
rect 662 1237 668 1238
rect 718 1242 724 1243
rect 718 1238 719 1242
rect 723 1238 724 1242
rect 718 1237 724 1238
rect 766 1242 772 1243
rect 766 1238 767 1242
rect 771 1238 772 1242
rect 766 1237 772 1238
rect 814 1242 820 1243
rect 814 1238 815 1242
rect 819 1238 820 1242
rect 814 1237 820 1238
rect 870 1242 876 1243
rect 870 1238 871 1242
rect 875 1238 876 1242
rect 870 1237 876 1238
rect 926 1242 932 1243
rect 926 1238 927 1242
rect 931 1238 932 1242
rect 926 1237 932 1238
rect 982 1242 988 1243
rect 982 1238 983 1242
rect 987 1238 988 1242
rect 982 1237 988 1238
rect 1038 1242 1044 1243
rect 1038 1238 1039 1242
rect 1043 1238 1044 1242
rect 1038 1237 1044 1238
rect 1094 1242 1100 1243
rect 1094 1238 1095 1242
rect 1099 1238 1100 1242
rect 1094 1237 1100 1238
rect 1158 1242 1164 1243
rect 1158 1238 1159 1242
rect 1163 1238 1164 1242
rect 1158 1237 1164 1238
rect 1230 1242 1236 1243
rect 1230 1238 1231 1242
rect 1235 1238 1236 1242
rect 1230 1237 1236 1238
rect 1318 1242 1324 1243
rect 1318 1238 1319 1242
rect 1323 1238 1324 1242
rect 1318 1237 1324 1238
rect 1422 1242 1428 1243
rect 1422 1238 1423 1242
rect 1427 1238 1428 1242
rect 1422 1237 1428 1238
rect 1534 1242 1540 1243
rect 1534 1238 1535 1242
rect 1539 1238 1540 1242
rect 1534 1237 1540 1238
rect 1622 1242 1628 1243
rect 1622 1238 1623 1242
rect 1627 1238 1628 1242
rect 1622 1237 1628 1238
rect 1662 1240 1668 1241
rect 110 1235 116 1236
rect 112 1223 114 1235
rect 136 1223 138 1237
rect 168 1223 170 1237
rect 224 1223 226 1237
rect 280 1223 282 1237
rect 328 1223 330 1237
rect 384 1223 386 1237
rect 440 1223 442 1237
rect 496 1223 498 1237
rect 552 1223 554 1237
rect 608 1223 610 1237
rect 664 1223 666 1237
rect 720 1223 722 1237
rect 768 1223 770 1237
rect 816 1223 818 1237
rect 872 1223 874 1237
rect 928 1223 930 1237
rect 984 1223 986 1237
rect 1040 1223 1042 1237
rect 1096 1223 1098 1237
rect 1160 1223 1162 1237
rect 1232 1223 1234 1237
rect 1320 1223 1322 1237
rect 1424 1223 1426 1237
rect 1536 1223 1538 1237
rect 1624 1223 1626 1237
rect 1662 1236 1663 1240
rect 1667 1236 1668 1240
rect 1662 1235 1668 1236
rect 1664 1223 1666 1235
rect 111 1222 115 1223
rect 111 1217 115 1218
rect 135 1222 139 1223
rect 135 1217 139 1218
rect 167 1222 171 1223
rect 167 1217 171 1218
rect 223 1222 227 1223
rect 223 1217 227 1218
rect 279 1222 283 1223
rect 279 1217 283 1218
rect 327 1222 331 1223
rect 327 1217 331 1218
rect 335 1222 339 1223
rect 335 1217 339 1218
rect 383 1222 387 1223
rect 383 1217 387 1218
rect 431 1222 435 1223
rect 431 1217 435 1218
rect 439 1222 443 1223
rect 439 1217 443 1218
rect 487 1222 491 1223
rect 487 1217 491 1218
rect 495 1222 499 1223
rect 495 1217 499 1218
rect 543 1222 547 1223
rect 543 1217 547 1218
rect 551 1222 555 1223
rect 551 1217 555 1218
rect 599 1222 603 1223
rect 599 1217 603 1218
rect 607 1222 611 1223
rect 607 1217 611 1218
rect 655 1222 659 1223
rect 655 1217 659 1218
rect 663 1222 667 1223
rect 663 1217 667 1218
rect 711 1222 715 1223
rect 711 1217 715 1218
rect 719 1222 723 1223
rect 719 1217 723 1218
rect 767 1222 771 1223
rect 767 1217 771 1218
rect 815 1222 819 1223
rect 815 1217 819 1218
rect 823 1222 827 1223
rect 823 1217 827 1218
rect 871 1222 875 1223
rect 871 1217 875 1218
rect 887 1222 891 1223
rect 887 1217 891 1218
rect 927 1222 931 1223
rect 927 1217 931 1218
rect 951 1222 955 1223
rect 951 1217 955 1218
rect 983 1222 987 1223
rect 983 1217 987 1218
rect 1015 1222 1019 1223
rect 1015 1217 1019 1218
rect 1039 1222 1043 1223
rect 1039 1217 1043 1218
rect 1079 1222 1083 1223
rect 1079 1217 1083 1218
rect 1095 1222 1099 1223
rect 1095 1217 1099 1218
rect 1143 1222 1147 1223
rect 1143 1217 1147 1218
rect 1159 1222 1163 1223
rect 1159 1217 1163 1218
rect 1207 1222 1211 1223
rect 1207 1217 1211 1218
rect 1231 1222 1235 1223
rect 1231 1217 1235 1218
rect 1279 1222 1283 1223
rect 1279 1217 1283 1218
rect 1319 1222 1323 1223
rect 1319 1217 1323 1218
rect 1359 1222 1363 1223
rect 1359 1217 1363 1218
rect 1423 1222 1427 1223
rect 1423 1217 1427 1218
rect 1447 1222 1451 1223
rect 1447 1217 1451 1218
rect 1535 1222 1539 1223
rect 1535 1217 1539 1218
rect 1543 1222 1547 1223
rect 1543 1217 1547 1218
rect 1623 1222 1627 1223
rect 1623 1217 1627 1218
rect 1663 1222 1667 1223
rect 1663 1217 1667 1218
rect 112 1209 114 1217
rect 110 1208 116 1209
rect 110 1204 111 1208
rect 115 1204 116 1208
rect 136 1207 138 1217
rect 168 1207 170 1217
rect 224 1207 226 1217
rect 280 1207 282 1217
rect 336 1207 338 1217
rect 384 1207 386 1217
rect 432 1207 434 1217
rect 488 1207 490 1217
rect 544 1207 546 1217
rect 600 1207 602 1217
rect 656 1207 658 1217
rect 712 1207 714 1217
rect 768 1207 770 1217
rect 824 1207 826 1217
rect 888 1207 890 1217
rect 952 1207 954 1217
rect 1016 1207 1018 1217
rect 1080 1207 1082 1217
rect 1144 1207 1146 1217
rect 1208 1207 1210 1217
rect 1280 1207 1282 1217
rect 1360 1207 1362 1217
rect 1448 1207 1450 1217
rect 1544 1207 1546 1217
rect 1624 1207 1626 1217
rect 1664 1209 1666 1217
rect 1662 1208 1668 1209
rect 110 1203 116 1204
rect 134 1206 140 1207
rect 134 1202 135 1206
rect 139 1202 140 1206
rect 134 1201 140 1202
rect 166 1206 172 1207
rect 166 1202 167 1206
rect 171 1202 172 1206
rect 166 1201 172 1202
rect 222 1206 228 1207
rect 222 1202 223 1206
rect 227 1202 228 1206
rect 222 1201 228 1202
rect 278 1206 284 1207
rect 278 1202 279 1206
rect 283 1202 284 1206
rect 278 1201 284 1202
rect 334 1206 340 1207
rect 334 1202 335 1206
rect 339 1202 340 1206
rect 334 1201 340 1202
rect 382 1206 388 1207
rect 382 1202 383 1206
rect 387 1202 388 1206
rect 382 1201 388 1202
rect 430 1206 436 1207
rect 430 1202 431 1206
rect 435 1202 436 1206
rect 430 1201 436 1202
rect 486 1206 492 1207
rect 486 1202 487 1206
rect 491 1202 492 1206
rect 486 1201 492 1202
rect 542 1206 548 1207
rect 542 1202 543 1206
rect 547 1202 548 1206
rect 542 1201 548 1202
rect 598 1206 604 1207
rect 598 1202 599 1206
rect 603 1202 604 1206
rect 598 1201 604 1202
rect 654 1206 660 1207
rect 654 1202 655 1206
rect 659 1202 660 1206
rect 654 1201 660 1202
rect 710 1206 716 1207
rect 710 1202 711 1206
rect 715 1202 716 1206
rect 710 1201 716 1202
rect 766 1206 772 1207
rect 766 1202 767 1206
rect 771 1202 772 1206
rect 766 1201 772 1202
rect 822 1206 828 1207
rect 822 1202 823 1206
rect 827 1202 828 1206
rect 822 1201 828 1202
rect 886 1206 892 1207
rect 886 1202 887 1206
rect 891 1202 892 1206
rect 886 1201 892 1202
rect 950 1206 956 1207
rect 950 1202 951 1206
rect 955 1202 956 1206
rect 950 1201 956 1202
rect 1014 1206 1020 1207
rect 1014 1202 1015 1206
rect 1019 1202 1020 1206
rect 1014 1201 1020 1202
rect 1078 1206 1084 1207
rect 1078 1202 1079 1206
rect 1083 1202 1084 1206
rect 1078 1201 1084 1202
rect 1142 1206 1148 1207
rect 1142 1202 1143 1206
rect 1147 1202 1148 1206
rect 1142 1201 1148 1202
rect 1206 1206 1212 1207
rect 1206 1202 1207 1206
rect 1211 1202 1212 1206
rect 1206 1201 1212 1202
rect 1278 1206 1284 1207
rect 1278 1202 1279 1206
rect 1283 1202 1284 1206
rect 1278 1201 1284 1202
rect 1358 1206 1364 1207
rect 1358 1202 1359 1206
rect 1363 1202 1364 1206
rect 1358 1201 1364 1202
rect 1446 1206 1452 1207
rect 1446 1202 1447 1206
rect 1451 1202 1452 1206
rect 1446 1201 1452 1202
rect 1542 1206 1548 1207
rect 1542 1202 1543 1206
rect 1547 1202 1548 1206
rect 1542 1201 1548 1202
rect 1622 1206 1628 1207
rect 1622 1202 1623 1206
rect 1627 1202 1628 1206
rect 1662 1204 1663 1208
rect 1667 1204 1668 1208
rect 1662 1203 1668 1204
rect 1622 1201 1628 1202
rect 110 1191 116 1192
rect 110 1187 111 1191
rect 115 1187 116 1191
rect 1662 1191 1668 1192
rect 110 1186 116 1187
rect 134 1189 140 1190
rect 112 1179 114 1186
rect 134 1185 135 1189
rect 139 1185 140 1189
rect 134 1184 140 1185
rect 166 1189 172 1190
rect 166 1185 167 1189
rect 171 1185 172 1189
rect 166 1184 172 1185
rect 222 1189 228 1190
rect 222 1185 223 1189
rect 227 1185 228 1189
rect 222 1184 228 1185
rect 278 1189 284 1190
rect 278 1185 279 1189
rect 283 1185 284 1189
rect 278 1184 284 1185
rect 334 1189 340 1190
rect 334 1185 335 1189
rect 339 1185 340 1189
rect 334 1184 340 1185
rect 382 1189 388 1190
rect 382 1185 383 1189
rect 387 1185 388 1189
rect 382 1184 388 1185
rect 430 1189 436 1190
rect 430 1185 431 1189
rect 435 1185 436 1189
rect 430 1184 436 1185
rect 486 1189 492 1190
rect 486 1185 487 1189
rect 491 1185 492 1189
rect 486 1184 492 1185
rect 542 1189 548 1190
rect 542 1185 543 1189
rect 547 1185 548 1189
rect 542 1184 548 1185
rect 598 1189 604 1190
rect 598 1185 599 1189
rect 603 1185 604 1189
rect 598 1184 604 1185
rect 654 1189 660 1190
rect 654 1185 655 1189
rect 659 1185 660 1189
rect 654 1184 660 1185
rect 710 1189 716 1190
rect 710 1185 711 1189
rect 715 1185 716 1189
rect 710 1184 716 1185
rect 766 1189 772 1190
rect 766 1185 767 1189
rect 771 1185 772 1189
rect 766 1184 772 1185
rect 822 1189 828 1190
rect 822 1185 823 1189
rect 827 1185 828 1189
rect 822 1184 828 1185
rect 886 1189 892 1190
rect 886 1185 887 1189
rect 891 1185 892 1189
rect 886 1184 892 1185
rect 950 1189 956 1190
rect 950 1185 951 1189
rect 955 1185 956 1189
rect 950 1184 956 1185
rect 1014 1189 1020 1190
rect 1014 1185 1015 1189
rect 1019 1185 1020 1189
rect 1014 1184 1020 1185
rect 1078 1189 1084 1190
rect 1078 1185 1079 1189
rect 1083 1185 1084 1189
rect 1078 1184 1084 1185
rect 1142 1189 1148 1190
rect 1142 1185 1143 1189
rect 1147 1185 1148 1189
rect 1142 1184 1148 1185
rect 1206 1189 1212 1190
rect 1206 1185 1207 1189
rect 1211 1185 1212 1189
rect 1206 1184 1212 1185
rect 1278 1189 1284 1190
rect 1278 1185 1279 1189
rect 1283 1185 1284 1189
rect 1278 1184 1284 1185
rect 1358 1189 1364 1190
rect 1358 1185 1359 1189
rect 1363 1185 1364 1189
rect 1358 1184 1364 1185
rect 1446 1189 1452 1190
rect 1446 1185 1447 1189
rect 1451 1185 1452 1189
rect 1446 1184 1452 1185
rect 1542 1189 1548 1190
rect 1542 1185 1543 1189
rect 1547 1185 1548 1189
rect 1542 1184 1548 1185
rect 1622 1189 1628 1190
rect 1622 1185 1623 1189
rect 1627 1185 1628 1189
rect 1662 1187 1663 1191
rect 1667 1187 1668 1191
rect 1662 1186 1668 1187
rect 1622 1184 1628 1185
rect 136 1179 138 1184
rect 168 1179 170 1184
rect 224 1179 226 1184
rect 280 1179 282 1184
rect 336 1179 338 1184
rect 384 1179 386 1184
rect 432 1179 434 1184
rect 488 1179 490 1184
rect 544 1179 546 1184
rect 600 1179 602 1184
rect 656 1179 658 1184
rect 712 1179 714 1184
rect 768 1179 770 1184
rect 824 1179 826 1184
rect 888 1179 890 1184
rect 952 1179 954 1184
rect 1016 1179 1018 1184
rect 1080 1179 1082 1184
rect 1144 1179 1146 1184
rect 1208 1179 1210 1184
rect 1280 1179 1282 1184
rect 1360 1179 1362 1184
rect 1448 1179 1450 1184
rect 1544 1179 1546 1184
rect 1624 1179 1626 1184
rect 1664 1179 1666 1186
rect 111 1178 115 1179
rect 111 1173 115 1174
rect 135 1178 139 1179
rect 112 1170 114 1173
rect 135 1172 139 1174
rect 167 1178 171 1179
rect 167 1172 171 1174
rect 223 1178 227 1179
rect 223 1172 227 1174
rect 279 1178 283 1179
rect 279 1173 283 1174
rect 287 1178 291 1179
rect 287 1172 291 1174
rect 335 1178 339 1179
rect 335 1173 339 1174
rect 351 1178 355 1179
rect 351 1172 355 1174
rect 383 1178 387 1179
rect 383 1173 387 1174
rect 415 1178 419 1179
rect 415 1172 419 1174
rect 431 1178 435 1179
rect 431 1173 435 1174
rect 471 1178 475 1179
rect 471 1172 475 1174
rect 487 1178 491 1179
rect 487 1173 491 1174
rect 535 1178 539 1179
rect 535 1172 539 1174
rect 543 1178 547 1179
rect 543 1173 547 1174
rect 599 1178 603 1179
rect 599 1172 603 1174
rect 655 1178 659 1179
rect 655 1173 659 1174
rect 663 1178 667 1179
rect 663 1172 667 1174
rect 711 1178 715 1179
rect 711 1173 715 1174
rect 727 1178 731 1179
rect 727 1172 731 1174
rect 767 1178 771 1179
rect 767 1173 771 1174
rect 783 1178 787 1179
rect 783 1172 787 1174
rect 823 1178 827 1179
rect 823 1173 827 1174
rect 839 1178 843 1179
rect 839 1172 843 1174
rect 887 1178 891 1179
rect 887 1173 891 1174
rect 903 1178 907 1179
rect 903 1172 907 1174
rect 951 1178 955 1179
rect 951 1173 955 1174
rect 967 1178 971 1179
rect 967 1172 971 1174
rect 1015 1178 1019 1179
rect 1015 1173 1019 1174
rect 1031 1178 1035 1179
rect 1031 1172 1035 1174
rect 1079 1178 1083 1179
rect 1079 1173 1083 1174
rect 1095 1178 1099 1179
rect 1095 1172 1099 1174
rect 1143 1178 1147 1179
rect 1143 1173 1147 1174
rect 1159 1178 1163 1179
rect 1159 1172 1163 1174
rect 1207 1178 1211 1179
rect 1207 1173 1211 1174
rect 1215 1178 1219 1179
rect 1215 1172 1219 1174
rect 1279 1178 1283 1179
rect 1279 1172 1283 1174
rect 1343 1178 1347 1179
rect 1343 1172 1347 1174
rect 1359 1178 1363 1179
rect 1359 1173 1363 1174
rect 1407 1178 1411 1179
rect 1407 1172 1411 1174
rect 1447 1178 1451 1179
rect 1447 1173 1451 1174
rect 1479 1178 1483 1179
rect 1479 1172 1483 1174
rect 1543 1178 1547 1179
rect 1543 1173 1547 1174
rect 1559 1178 1563 1179
rect 1559 1172 1563 1174
rect 1623 1178 1627 1179
rect 1623 1172 1627 1174
rect 1663 1178 1667 1179
rect 1663 1173 1667 1174
rect 134 1171 140 1172
rect 110 1169 116 1170
rect 110 1165 111 1169
rect 115 1165 116 1169
rect 134 1167 135 1171
rect 139 1167 140 1171
rect 134 1166 140 1167
rect 166 1171 172 1172
rect 166 1167 167 1171
rect 171 1167 172 1171
rect 166 1166 172 1167
rect 222 1171 228 1172
rect 222 1167 223 1171
rect 227 1167 228 1171
rect 222 1166 228 1167
rect 286 1171 292 1172
rect 286 1167 287 1171
rect 291 1167 292 1171
rect 286 1166 292 1167
rect 350 1171 356 1172
rect 350 1167 351 1171
rect 355 1167 356 1171
rect 350 1166 356 1167
rect 414 1171 420 1172
rect 414 1167 415 1171
rect 419 1167 420 1171
rect 414 1166 420 1167
rect 470 1171 476 1172
rect 470 1167 471 1171
rect 475 1167 476 1171
rect 470 1166 476 1167
rect 534 1171 540 1172
rect 534 1167 535 1171
rect 539 1167 540 1171
rect 534 1166 540 1167
rect 598 1171 604 1172
rect 598 1167 599 1171
rect 603 1167 604 1171
rect 598 1166 604 1167
rect 662 1171 668 1172
rect 662 1167 663 1171
rect 667 1167 668 1171
rect 662 1166 668 1167
rect 726 1171 732 1172
rect 726 1167 727 1171
rect 731 1167 732 1171
rect 726 1166 732 1167
rect 782 1171 788 1172
rect 782 1167 783 1171
rect 787 1167 788 1171
rect 782 1166 788 1167
rect 838 1171 844 1172
rect 838 1167 839 1171
rect 843 1167 844 1171
rect 838 1166 844 1167
rect 902 1171 908 1172
rect 902 1167 903 1171
rect 907 1167 908 1171
rect 902 1166 908 1167
rect 966 1171 972 1172
rect 966 1167 967 1171
rect 971 1167 972 1171
rect 966 1166 972 1167
rect 1030 1171 1036 1172
rect 1030 1167 1031 1171
rect 1035 1167 1036 1171
rect 1030 1166 1036 1167
rect 1094 1171 1100 1172
rect 1094 1167 1095 1171
rect 1099 1167 1100 1171
rect 1094 1166 1100 1167
rect 1158 1171 1164 1172
rect 1158 1167 1159 1171
rect 1163 1167 1164 1171
rect 1158 1166 1164 1167
rect 1214 1171 1220 1172
rect 1214 1167 1215 1171
rect 1219 1167 1220 1171
rect 1214 1166 1220 1167
rect 1278 1171 1284 1172
rect 1278 1167 1279 1171
rect 1283 1167 1284 1171
rect 1278 1166 1284 1167
rect 1342 1171 1348 1172
rect 1342 1167 1343 1171
rect 1347 1167 1348 1171
rect 1342 1166 1348 1167
rect 1406 1171 1412 1172
rect 1406 1167 1407 1171
rect 1411 1167 1412 1171
rect 1406 1166 1412 1167
rect 1478 1171 1484 1172
rect 1478 1167 1479 1171
rect 1483 1167 1484 1171
rect 1478 1166 1484 1167
rect 1558 1171 1564 1172
rect 1558 1167 1559 1171
rect 1563 1167 1564 1171
rect 1558 1166 1564 1167
rect 1622 1171 1628 1172
rect 1622 1167 1623 1171
rect 1627 1167 1628 1171
rect 1664 1170 1666 1173
rect 1622 1166 1628 1167
rect 1662 1169 1668 1170
rect 110 1164 116 1165
rect 1662 1165 1663 1169
rect 1667 1165 1668 1169
rect 1662 1164 1668 1165
rect 134 1154 140 1155
rect 110 1152 116 1153
rect 110 1148 111 1152
rect 115 1148 116 1152
rect 134 1150 135 1154
rect 139 1150 140 1154
rect 134 1149 140 1150
rect 166 1154 172 1155
rect 166 1150 167 1154
rect 171 1150 172 1154
rect 166 1149 172 1150
rect 222 1154 228 1155
rect 222 1150 223 1154
rect 227 1150 228 1154
rect 222 1149 228 1150
rect 286 1154 292 1155
rect 286 1150 287 1154
rect 291 1150 292 1154
rect 286 1149 292 1150
rect 350 1154 356 1155
rect 350 1150 351 1154
rect 355 1150 356 1154
rect 350 1149 356 1150
rect 414 1154 420 1155
rect 414 1150 415 1154
rect 419 1150 420 1154
rect 414 1149 420 1150
rect 470 1154 476 1155
rect 470 1150 471 1154
rect 475 1150 476 1154
rect 470 1149 476 1150
rect 534 1154 540 1155
rect 534 1150 535 1154
rect 539 1150 540 1154
rect 534 1149 540 1150
rect 598 1154 604 1155
rect 598 1150 599 1154
rect 603 1150 604 1154
rect 598 1149 604 1150
rect 662 1154 668 1155
rect 662 1150 663 1154
rect 667 1150 668 1154
rect 662 1149 668 1150
rect 726 1154 732 1155
rect 726 1150 727 1154
rect 731 1150 732 1154
rect 726 1149 732 1150
rect 782 1154 788 1155
rect 782 1150 783 1154
rect 787 1150 788 1154
rect 782 1149 788 1150
rect 838 1154 844 1155
rect 838 1150 839 1154
rect 843 1150 844 1154
rect 838 1149 844 1150
rect 902 1154 908 1155
rect 902 1150 903 1154
rect 907 1150 908 1154
rect 902 1149 908 1150
rect 966 1154 972 1155
rect 966 1150 967 1154
rect 971 1150 972 1154
rect 966 1149 972 1150
rect 1030 1154 1036 1155
rect 1030 1150 1031 1154
rect 1035 1150 1036 1154
rect 1030 1149 1036 1150
rect 1094 1154 1100 1155
rect 1094 1150 1095 1154
rect 1099 1150 1100 1154
rect 1094 1149 1100 1150
rect 1158 1154 1164 1155
rect 1158 1150 1159 1154
rect 1163 1150 1164 1154
rect 1158 1149 1164 1150
rect 1214 1154 1220 1155
rect 1214 1150 1215 1154
rect 1219 1150 1220 1154
rect 1214 1149 1220 1150
rect 1278 1154 1284 1155
rect 1278 1150 1279 1154
rect 1283 1150 1284 1154
rect 1278 1149 1284 1150
rect 1342 1154 1348 1155
rect 1342 1150 1343 1154
rect 1347 1150 1348 1154
rect 1342 1149 1348 1150
rect 1406 1154 1412 1155
rect 1406 1150 1407 1154
rect 1411 1150 1412 1154
rect 1406 1149 1412 1150
rect 1478 1154 1484 1155
rect 1478 1150 1479 1154
rect 1483 1150 1484 1154
rect 1478 1149 1484 1150
rect 1558 1154 1564 1155
rect 1558 1150 1559 1154
rect 1563 1150 1564 1154
rect 1558 1149 1564 1150
rect 1622 1154 1628 1155
rect 1622 1150 1623 1154
rect 1627 1150 1628 1154
rect 1622 1149 1628 1150
rect 1662 1152 1668 1153
rect 110 1147 116 1148
rect 112 1135 114 1147
rect 136 1135 138 1149
rect 168 1135 170 1149
rect 224 1135 226 1149
rect 288 1135 290 1149
rect 352 1135 354 1149
rect 416 1135 418 1149
rect 472 1135 474 1149
rect 536 1135 538 1149
rect 600 1135 602 1149
rect 664 1135 666 1149
rect 728 1135 730 1149
rect 784 1135 786 1149
rect 840 1135 842 1149
rect 904 1135 906 1149
rect 968 1135 970 1149
rect 1032 1135 1034 1149
rect 1096 1135 1098 1149
rect 1160 1135 1162 1149
rect 1216 1135 1218 1149
rect 1280 1135 1282 1149
rect 1344 1135 1346 1149
rect 1408 1135 1410 1149
rect 1480 1135 1482 1149
rect 1560 1135 1562 1149
rect 1624 1135 1626 1149
rect 1662 1148 1663 1152
rect 1667 1148 1668 1152
rect 1662 1147 1668 1148
rect 1664 1135 1666 1147
rect 111 1134 115 1135
rect 111 1129 115 1130
rect 135 1134 139 1135
rect 135 1129 139 1130
rect 143 1134 147 1135
rect 143 1129 147 1130
rect 167 1134 171 1135
rect 167 1129 171 1130
rect 175 1134 179 1135
rect 175 1129 179 1130
rect 215 1134 219 1135
rect 215 1129 219 1130
rect 223 1134 227 1135
rect 223 1129 227 1130
rect 271 1134 275 1135
rect 271 1129 275 1130
rect 287 1134 291 1135
rect 287 1129 291 1130
rect 335 1134 339 1135
rect 335 1129 339 1130
rect 351 1134 355 1135
rect 351 1129 355 1130
rect 399 1134 403 1135
rect 399 1129 403 1130
rect 415 1134 419 1135
rect 415 1129 419 1130
rect 463 1134 467 1135
rect 463 1129 467 1130
rect 471 1134 475 1135
rect 471 1129 475 1130
rect 527 1134 531 1135
rect 527 1129 531 1130
rect 535 1134 539 1135
rect 535 1129 539 1130
rect 599 1134 603 1135
rect 599 1129 603 1130
rect 663 1134 667 1135
rect 663 1129 667 1130
rect 727 1134 731 1135
rect 727 1129 731 1130
rect 783 1134 787 1135
rect 783 1129 787 1130
rect 791 1134 795 1135
rect 791 1129 795 1130
rect 839 1134 843 1135
rect 839 1129 843 1130
rect 855 1134 859 1135
rect 855 1129 859 1130
rect 903 1134 907 1135
rect 903 1129 907 1130
rect 911 1134 915 1135
rect 911 1129 915 1130
rect 967 1134 971 1135
rect 967 1129 971 1130
rect 1023 1134 1027 1135
rect 1023 1129 1027 1130
rect 1031 1134 1035 1135
rect 1031 1129 1035 1130
rect 1087 1134 1091 1135
rect 1087 1129 1091 1130
rect 1095 1134 1099 1135
rect 1095 1129 1099 1130
rect 1151 1134 1155 1135
rect 1151 1129 1155 1130
rect 1159 1134 1163 1135
rect 1159 1129 1163 1130
rect 1215 1134 1219 1135
rect 1215 1129 1219 1130
rect 1279 1134 1283 1135
rect 1279 1129 1283 1130
rect 1335 1134 1339 1135
rect 1335 1129 1339 1130
rect 1343 1134 1347 1135
rect 1343 1129 1347 1130
rect 1391 1134 1395 1135
rect 1391 1129 1395 1130
rect 1407 1134 1411 1135
rect 1407 1129 1411 1130
rect 1447 1134 1451 1135
rect 1447 1129 1451 1130
rect 1479 1134 1483 1135
rect 1479 1129 1483 1130
rect 1495 1134 1499 1135
rect 1495 1129 1499 1130
rect 1543 1134 1547 1135
rect 1543 1129 1547 1130
rect 1559 1134 1563 1135
rect 1559 1129 1563 1130
rect 1591 1134 1595 1135
rect 1591 1129 1595 1130
rect 1623 1134 1627 1135
rect 1623 1129 1627 1130
rect 1663 1134 1667 1135
rect 1663 1129 1667 1130
rect 112 1121 114 1129
rect 110 1120 116 1121
rect 110 1116 111 1120
rect 115 1116 116 1120
rect 144 1119 146 1129
rect 176 1119 178 1129
rect 216 1119 218 1129
rect 272 1119 274 1129
rect 336 1119 338 1129
rect 400 1119 402 1129
rect 464 1119 466 1129
rect 528 1119 530 1129
rect 600 1119 602 1129
rect 664 1119 666 1129
rect 728 1119 730 1129
rect 792 1119 794 1129
rect 856 1119 858 1129
rect 912 1119 914 1129
rect 968 1119 970 1129
rect 1024 1119 1026 1129
rect 1088 1119 1090 1129
rect 1152 1119 1154 1129
rect 1216 1119 1218 1129
rect 1280 1119 1282 1129
rect 1336 1119 1338 1129
rect 1392 1119 1394 1129
rect 1448 1119 1450 1129
rect 1496 1119 1498 1129
rect 1544 1119 1546 1129
rect 1592 1119 1594 1129
rect 1624 1119 1626 1129
rect 1664 1121 1666 1129
rect 1662 1120 1668 1121
rect 110 1115 116 1116
rect 142 1118 148 1119
rect 142 1114 143 1118
rect 147 1114 148 1118
rect 142 1113 148 1114
rect 174 1118 180 1119
rect 174 1114 175 1118
rect 179 1114 180 1118
rect 174 1113 180 1114
rect 214 1118 220 1119
rect 214 1114 215 1118
rect 219 1114 220 1118
rect 214 1113 220 1114
rect 270 1118 276 1119
rect 270 1114 271 1118
rect 275 1114 276 1118
rect 270 1113 276 1114
rect 334 1118 340 1119
rect 334 1114 335 1118
rect 339 1114 340 1118
rect 334 1113 340 1114
rect 398 1118 404 1119
rect 398 1114 399 1118
rect 403 1114 404 1118
rect 398 1113 404 1114
rect 462 1118 468 1119
rect 462 1114 463 1118
rect 467 1114 468 1118
rect 462 1113 468 1114
rect 526 1118 532 1119
rect 526 1114 527 1118
rect 531 1114 532 1118
rect 526 1113 532 1114
rect 598 1118 604 1119
rect 598 1114 599 1118
rect 603 1114 604 1118
rect 598 1113 604 1114
rect 662 1118 668 1119
rect 662 1114 663 1118
rect 667 1114 668 1118
rect 662 1113 668 1114
rect 726 1118 732 1119
rect 726 1114 727 1118
rect 731 1114 732 1118
rect 726 1113 732 1114
rect 790 1118 796 1119
rect 790 1114 791 1118
rect 795 1114 796 1118
rect 790 1113 796 1114
rect 854 1118 860 1119
rect 854 1114 855 1118
rect 859 1114 860 1118
rect 854 1113 860 1114
rect 910 1118 916 1119
rect 910 1114 911 1118
rect 915 1114 916 1118
rect 910 1113 916 1114
rect 966 1118 972 1119
rect 966 1114 967 1118
rect 971 1114 972 1118
rect 966 1113 972 1114
rect 1022 1118 1028 1119
rect 1022 1114 1023 1118
rect 1027 1114 1028 1118
rect 1022 1113 1028 1114
rect 1086 1118 1092 1119
rect 1086 1114 1087 1118
rect 1091 1114 1092 1118
rect 1086 1113 1092 1114
rect 1150 1118 1156 1119
rect 1150 1114 1151 1118
rect 1155 1114 1156 1118
rect 1150 1113 1156 1114
rect 1214 1118 1220 1119
rect 1214 1114 1215 1118
rect 1219 1114 1220 1118
rect 1214 1113 1220 1114
rect 1278 1118 1284 1119
rect 1278 1114 1279 1118
rect 1283 1114 1284 1118
rect 1278 1113 1284 1114
rect 1334 1118 1340 1119
rect 1334 1114 1335 1118
rect 1339 1114 1340 1118
rect 1334 1113 1340 1114
rect 1390 1118 1396 1119
rect 1390 1114 1391 1118
rect 1395 1114 1396 1118
rect 1390 1113 1396 1114
rect 1446 1118 1452 1119
rect 1446 1114 1447 1118
rect 1451 1114 1452 1118
rect 1446 1113 1452 1114
rect 1494 1118 1500 1119
rect 1494 1114 1495 1118
rect 1499 1114 1500 1118
rect 1494 1113 1500 1114
rect 1542 1118 1548 1119
rect 1542 1114 1543 1118
rect 1547 1114 1548 1118
rect 1542 1113 1548 1114
rect 1590 1118 1596 1119
rect 1590 1114 1591 1118
rect 1595 1114 1596 1118
rect 1590 1113 1596 1114
rect 1622 1118 1628 1119
rect 1622 1114 1623 1118
rect 1627 1114 1628 1118
rect 1662 1116 1663 1120
rect 1667 1116 1668 1120
rect 1662 1115 1668 1116
rect 1622 1113 1628 1114
rect 110 1103 116 1104
rect 110 1099 111 1103
rect 115 1099 116 1103
rect 1662 1103 1668 1104
rect 110 1098 116 1099
rect 142 1101 148 1102
rect 112 1091 114 1098
rect 142 1097 143 1101
rect 147 1097 148 1101
rect 142 1096 148 1097
rect 174 1101 180 1102
rect 174 1097 175 1101
rect 179 1097 180 1101
rect 174 1096 180 1097
rect 214 1101 220 1102
rect 214 1097 215 1101
rect 219 1097 220 1101
rect 214 1096 220 1097
rect 270 1101 276 1102
rect 270 1097 271 1101
rect 275 1097 276 1101
rect 270 1096 276 1097
rect 334 1101 340 1102
rect 334 1097 335 1101
rect 339 1097 340 1101
rect 334 1096 340 1097
rect 398 1101 404 1102
rect 398 1097 399 1101
rect 403 1097 404 1101
rect 398 1096 404 1097
rect 462 1101 468 1102
rect 462 1097 463 1101
rect 467 1097 468 1101
rect 462 1096 468 1097
rect 526 1101 532 1102
rect 526 1097 527 1101
rect 531 1097 532 1101
rect 526 1096 532 1097
rect 598 1101 604 1102
rect 598 1097 599 1101
rect 603 1097 604 1101
rect 598 1096 604 1097
rect 662 1101 668 1102
rect 662 1097 663 1101
rect 667 1097 668 1101
rect 662 1096 668 1097
rect 726 1101 732 1102
rect 726 1097 727 1101
rect 731 1097 732 1101
rect 726 1096 732 1097
rect 790 1101 796 1102
rect 790 1097 791 1101
rect 795 1097 796 1101
rect 790 1096 796 1097
rect 854 1101 860 1102
rect 854 1097 855 1101
rect 859 1097 860 1101
rect 854 1096 860 1097
rect 910 1101 916 1102
rect 910 1097 911 1101
rect 915 1097 916 1101
rect 910 1096 916 1097
rect 966 1101 972 1102
rect 966 1097 967 1101
rect 971 1097 972 1101
rect 966 1096 972 1097
rect 1022 1101 1028 1102
rect 1022 1097 1023 1101
rect 1027 1097 1028 1101
rect 1022 1096 1028 1097
rect 1086 1101 1092 1102
rect 1086 1097 1087 1101
rect 1091 1097 1092 1101
rect 1086 1096 1092 1097
rect 1150 1101 1156 1102
rect 1150 1097 1151 1101
rect 1155 1097 1156 1101
rect 1150 1096 1156 1097
rect 1214 1101 1220 1102
rect 1214 1097 1215 1101
rect 1219 1097 1220 1101
rect 1214 1096 1220 1097
rect 1278 1101 1284 1102
rect 1278 1097 1279 1101
rect 1283 1097 1284 1101
rect 1278 1096 1284 1097
rect 1334 1101 1340 1102
rect 1334 1097 1335 1101
rect 1339 1097 1340 1101
rect 1334 1096 1340 1097
rect 1390 1101 1396 1102
rect 1390 1097 1391 1101
rect 1395 1097 1396 1101
rect 1390 1096 1396 1097
rect 1446 1101 1452 1102
rect 1446 1097 1447 1101
rect 1451 1097 1452 1101
rect 1446 1096 1452 1097
rect 1494 1101 1500 1102
rect 1494 1097 1495 1101
rect 1499 1097 1500 1101
rect 1494 1096 1500 1097
rect 1542 1101 1548 1102
rect 1542 1097 1543 1101
rect 1547 1097 1548 1101
rect 1542 1096 1548 1097
rect 1590 1101 1596 1102
rect 1590 1097 1591 1101
rect 1595 1097 1596 1101
rect 1590 1096 1596 1097
rect 1622 1101 1628 1102
rect 1622 1097 1623 1101
rect 1627 1097 1628 1101
rect 1662 1099 1663 1103
rect 1667 1099 1668 1103
rect 1662 1098 1668 1099
rect 1622 1096 1628 1097
rect 144 1091 146 1096
rect 176 1091 178 1096
rect 216 1091 218 1096
rect 272 1091 274 1096
rect 336 1091 338 1096
rect 400 1091 402 1096
rect 464 1091 466 1096
rect 528 1091 530 1096
rect 600 1091 602 1096
rect 664 1091 666 1096
rect 728 1091 730 1096
rect 792 1091 794 1096
rect 856 1091 858 1096
rect 912 1091 914 1096
rect 968 1091 970 1096
rect 1024 1091 1026 1096
rect 1088 1091 1090 1096
rect 1152 1091 1154 1096
rect 1216 1091 1218 1096
rect 1280 1091 1282 1096
rect 1336 1091 1338 1096
rect 1392 1091 1394 1096
rect 1448 1091 1450 1096
rect 1496 1091 1498 1096
rect 1544 1091 1546 1096
rect 1592 1091 1594 1096
rect 1624 1091 1626 1096
rect 1664 1091 1666 1098
rect 111 1090 115 1091
rect 111 1085 115 1086
rect 143 1090 147 1091
rect 143 1085 147 1086
rect 175 1090 179 1091
rect 175 1085 179 1086
rect 215 1090 219 1091
rect 112 1082 114 1085
rect 215 1084 219 1086
rect 247 1090 251 1091
rect 247 1084 251 1086
rect 271 1090 275 1091
rect 271 1085 275 1086
rect 279 1090 283 1091
rect 279 1084 283 1086
rect 311 1090 315 1091
rect 311 1084 315 1086
rect 335 1090 339 1091
rect 335 1085 339 1086
rect 351 1090 355 1091
rect 351 1084 355 1086
rect 391 1090 395 1091
rect 391 1084 395 1086
rect 399 1090 403 1091
rect 399 1085 403 1086
rect 439 1090 443 1091
rect 439 1084 443 1086
rect 463 1090 467 1091
rect 463 1085 467 1086
rect 503 1090 507 1091
rect 503 1084 507 1086
rect 527 1090 531 1091
rect 527 1085 531 1086
rect 575 1090 579 1091
rect 575 1084 579 1086
rect 599 1090 603 1091
rect 599 1085 603 1086
rect 655 1090 659 1091
rect 655 1084 659 1086
rect 663 1090 667 1091
rect 663 1085 667 1086
rect 727 1090 731 1091
rect 727 1085 731 1086
rect 735 1090 739 1091
rect 735 1084 739 1086
rect 791 1090 795 1091
rect 791 1085 795 1086
rect 815 1090 819 1091
rect 815 1084 819 1086
rect 855 1090 859 1091
rect 855 1085 859 1086
rect 895 1090 899 1091
rect 895 1084 899 1086
rect 911 1090 915 1091
rect 911 1085 915 1086
rect 967 1090 971 1091
rect 967 1084 971 1086
rect 1023 1090 1027 1091
rect 1023 1085 1027 1086
rect 1039 1090 1043 1091
rect 1039 1084 1043 1086
rect 1087 1090 1091 1091
rect 1087 1085 1091 1086
rect 1111 1090 1115 1091
rect 1111 1084 1115 1086
rect 1151 1090 1155 1091
rect 1151 1085 1155 1086
rect 1175 1090 1179 1091
rect 1175 1084 1179 1086
rect 1215 1090 1219 1091
rect 1215 1085 1219 1086
rect 1239 1090 1243 1091
rect 1239 1084 1243 1086
rect 1279 1090 1283 1091
rect 1279 1085 1283 1086
rect 1303 1090 1307 1091
rect 1303 1084 1307 1086
rect 1335 1090 1339 1091
rect 1335 1085 1339 1086
rect 1359 1090 1363 1091
rect 1359 1084 1363 1086
rect 1391 1090 1395 1091
rect 1391 1085 1395 1086
rect 1415 1090 1419 1091
rect 1415 1084 1419 1086
rect 1447 1090 1451 1091
rect 1447 1085 1451 1086
rect 1463 1090 1467 1091
rect 1463 1084 1467 1086
rect 1495 1090 1499 1091
rect 1495 1085 1499 1086
rect 1503 1090 1507 1091
rect 1503 1084 1507 1086
rect 1543 1090 1547 1091
rect 1543 1085 1547 1086
rect 1551 1090 1555 1091
rect 1551 1084 1555 1086
rect 1591 1090 1595 1091
rect 1591 1084 1595 1086
rect 1623 1090 1627 1091
rect 1623 1084 1627 1086
rect 1663 1090 1667 1091
rect 1663 1085 1667 1086
rect 214 1083 220 1084
rect 110 1081 116 1082
rect 110 1077 111 1081
rect 115 1077 116 1081
rect 214 1079 215 1083
rect 219 1079 220 1083
rect 214 1078 220 1079
rect 246 1083 252 1084
rect 246 1079 247 1083
rect 251 1079 252 1083
rect 246 1078 252 1079
rect 278 1083 284 1084
rect 278 1079 279 1083
rect 283 1079 284 1083
rect 278 1078 284 1079
rect 310 1083 316 1084
rect 310 1079 311 1083
rect 315 1079 316 1083
rect 310 1078 316 1079
rect 350 1083 356 1084
rect 350 1079 351 1083
rect 355 1079 356 1083
rect 350 1078 356 1079
rect 390 1083 396 1084
rect 390 1079 391 1083
rect 395 1079 396 1083
rect 390 1078 396 1079
rect 438 1083 444 1084
rect 438 1079 439 1083
rect 443 1079 444 1083
rect 438 1078 444 1079
rect 502 1083 508 1084
rect 502 1079 503 1083
rect 507 1079 508 1083
rect 502 1078 508 1079
rect 574 1083 580 1084
rect 574 1079 575 1083
rect 579 1079 580 1083
rect 574 1078 580 1079
rect 654 1083 660 1084
rect 654 1079 655 1083
rect 659 1079 660 1083
rect 654 1078 660 1079
rect 734 1083 740 1084
rect 734 1079 735 1083
rect 739 1079 740 1083
rect 734 1078 740 1079
rect 814 1083 820 1084
rect 814 1079 815 1083
rect 819 1079 820 1083
rect 814 1078 820 1079
rect 894 1083 900 1084
rect 894 1079 895 1083
rect 899 1079 900 1083
rect 894 1078 900 1079
rect 966 1083 972 1084
rect 966 1079 967 1083
rect 971 1079 972 1083
rect 966 1078 972 1079
rect 1038 1083 1044 1084
rect 1038 1079 1039 1083
rect 1043 1079 1044 1083
rect 1038 1078 1044 1079
rect 1110 1083 1116 1084
rect 1110 1079 1111 1083
rect 1115 1079 1116 1083
rect 1110 1078 1116 1079
rect 1174 1083 1180 1084
rect 1174 1079 1175 1083
rect 1179 1079 1180 1083
rect 1174 1078 1180 1079
rect 1238 1083 1244 1084
rect 1238 1079 1239 1083
rect 1243 1079 1244 1083
rect 1238 1078 1244 1079
rect 1302 1083 1308 1084
rect 1302 1079 1303 1083
rect 1307 1079 1308 1083
rect 1302 1078 1308 1079
rect 1358 1083 1364 1084
rect 1358 1079 1359 1083
rect 1363 1079 1364 1083
rect 1358 1078 1364 1079
rect 1414 1083 1420 1084
rect 1414 1079 1415 1083
rect 1419 1079 1420 1083
rect 1414 1078 1420 1079
rect 1462 1083 1468 1084
rect 1462 1079 1463 1083
rect 1467 1079 1468 1083
rect 1462 1078 1468 1079
rect 1502 1083 1508 1084
rect 1502 1079 1503 1083
rect 1507 1079 1508 1083
rect 1502 1078 1508 1079
rect 1550 1083 1556 1084
rect 1550 1079 1551 1083
rect 1555 1079 1556 1083
rect 1550 1078 1556 1079
rect 1590 1083 1596 1084
rect 1590 1079 1591 1083
rect 1595 1079 1596 1083
rect 1590 1078 1596 1079
rect 1622 1083 1628 1084
rect 1622 1079 1623 1083
rect 1627 1079 1628 1083
rect 1664 1082 1666 1085
rect 1622 1078 1628 1079
rect 1662 1081 1668 1082
rect 110 1076 116 1077
rect 1662 1077 1663 1081
rect 1667 1077 1668 1081
rect 1662 1076 1668 1077
rect 214 1066 220 1067
rect 110 1064 116 1065
rect 110 1060 111 1064
rect 115 1060 116 1064
rect 214 1062 215 1066
rect 219 1062 220 1066
rect 214 1061 220 1062
rect 246 1066 252 1067
rect 246 1062 247 1066
rect 251 1062 252 1066
rect 246 1061 252 1062
rect 278 1066 284 1067
rect 278 1062 279 1066
rect 283 1062 284 1066
rect 278 1061 284 1062
rect 310 1066 316 1067
rect 310 1062 311 1066
rect 315 1062 316 1066
rect 310 1061 316 1062
rect 350 1066 356 1067
rect 350 1062 351 1066
rect 355 1062 356 1066
rect 350 1061 356 1062
rect 390 1066 396 1067
rect 390 1062 391 1066
rect 395 1062 396 1066
rect 390 1061 396 1062
rect 438 1066 444 1067
rect 438 1062 439 1066
rect 443 1062 444 1066
rect 438 1061 444 1062
rect 502 1066 508 1067
rect 502 1062 503 1066
rect 507 1062 508 1066
rect 502 1061 508 1062
rect 574 1066 580 1067
rect 574 1062 575 1066
rect 579 1062 580 1066
rect 574 1061 580 1062
rect 654 1066 660 1067
rect 654 1062 655 1066
rect 659 1062 660 1066
rect 654 1061 660 1062
rect 734 1066 740 1067
rect 734 1062 735 1066
rect 739 1062 740 1066
rect 734 1061 740 1062
rect 814 1066 820 1067
rect 814 1062 815 1066
rect 819 1062 820 1066
rect 814 1061 820 1062
rect 894 1066 900 1067
rect 894 1062 895 1066
rect 899 1062 900 1066
rect 894 1061 900 1062
rect 966 1066 972 1067
rect 966 1062 967 1066
rect 971 1062 972 1066
rect 966 1061 972 1062
rect 1038 1066 1044 1067
rect 1038 1062 1039 1066
rect 1043 1062 1044 1066
rect 1038 1061 1044 1062
rect 1110 1066 1116 1067
rect 1110 1062 1111 1066
rect 1115 1062 1116 1066
rect 1110 1061 1116 1062
rect 1174 1066 1180 1067
rect 1174 1062 1175 1066
rect 1179 1062 1180 1066
rect 1174 1061 1180 1062
rect 1238 1066 1244 1067
rect 1238 1062 1239 1066
rect 1243 1062 1244 1066
rect 1238 1061 1244 1062
rect 1302 1066 1308 1067
rect 1302 1062 1303 1066
rect 1307 1062 1308 1066
rect 1302 1061 1308 1062
rect 1358 1066 1364 1067
rect 1358 1062 1359 1066
rect 1363 1062 1364 1066
rect 1358 1061 1364 1062
rect 1414 1066 1420 1067
rect 1414 1062 1415 1066
rect 1419 1062 1420 1066
rect 1414 1061 1420 1062
rect 1462 1066 1468 1067
rect 1462 1062 1463 1066
rect 1467 1062 1468 1066
rect 1462 1061 1468 1062
rect 1502 1066 1508 1067
rect 1502 1062 1503 1066
rect 1507 1062 1508 1066
rect 1502 1061 1508 1062
rect 1550 1066 1556 1067
rect 1550 1062 1551 1066
rect 1555 1062 1556 1066
rect 1550 1061 1556 1062
rect 1590 1066 1596 1067
rect 1590 1062 1591 1066
rect 1595 1062 1596 1066
rect 1590 1061 1596 1062
rect 1622 1066 1628 1067
rect 1622 1062 1623 1066
rect 1627 1062 1628 1066
rect 1622 1061 1628 1062
rect 1662 1064 1668 1065
rect 110 1059 116 1060
rect 112 1047 114 1059
rect 216 1047 218 1061
rect 248 1047 250 1061
rect 280 1047 282 1061
rect 312 1047 314 1061
rect 352 1047 354 1061
rect 392 1047 394 1061
rect 440 1047 442 1061
rect 504 1047 506 1061
rect 576 1047 578 1061
rect 656 1047 658 1061
rect 736 1047 738 1061
rect 816 1047 818 1061
rect 896 1047 898 1061
rect 968 1047 970 1061
rect 1040 1047 1042 1061
rect 1112 1047 1114 1061
rect 1176 1047 1178 1061
rect 1240 1047 1242 1061
rect 1304 1047 1306 1061
rect 1360 1047 1362 1061
rect 1416 1047 1418 1061
rect 1464 1047 1466 1061
rect 1504 1047 1506 1061
rect 1552 1047 1554 1061
rect 1592 1047 1594 1061
rect 1624 1047 1626 1061
rect 1662 1060 1663 1064
rect 1667 1060 1668 1064
rect 1662 1059 1668 1060
rect 1664 1047 1666 1059
rect 111 1046 115 1047
rect 111 1041 115 1042
rect 215 1046 219 1047
rect 215 1041 219 1042
rect 247 1046 251 1047
rect 247 1041 251 1042
rect 279 1046 283 1047
rect 279 1041 283 1042
rect 295 1046 299 1047
rect 295 1041 299 1042
rect 311 1046 315 1047
rect 311 1041 315 1042
rect 327 1046 331 1047
rect 327 1041 331 1042
rect 351 1046 355 1047
rect 351 1041 355 1042
rect 359 1046 363 1047
rect 359 1041 363 1042
rect 391 1046 395 1047
rect 391 1041 395 1042
rect 423 1046 427 1047
rect 423 1041 427 1042
rect 439 1046 443 1047
rect 439 1041 443 1042
rect 455 1046 459 1047
rect 455 1041 459 1042
rect 503 1046 507 1047
rect 503 1041 507 1042
rect 559 1046 563 1047
rect 559 1041 563 1042
rect 575 1046 579 1047
rect 575 1041 579 1042
rect 631 1046 635 1047
rect 631 1041 635 1042
rect 655 1046 659 1047
rect 655 1041 659 1042
rect 711 1046 715 1047
rect 711 1041 715 1042
rect 735 1046 739 1047
rect 735 1041 739 1042
rect 799 1046 803 1047
rect 799 1041 803 1042
rect 815 1046 819 1047
rect 815 1041 819 1042
rect 879 1046 883 1047
rect 879 1041 883 1042
rect 895 1046 899 1047
rect 895 1041 899 1042
rect 959 1046 963 1047
rect 959 1041 963 1042
rect 967 1046 971 1047
rect 967 1041 971 1042
rect 1031 1046 1035 1047
rect 1031 1041 1035 1042
rect 1039 1046 1043 1047
rect 1039 1041 1043 1042
rect 1095 1046 1099 1047
rect 1095 1041 1099 1042
rect 1111 1046 1115 1047
rect 1111 1041 1115 1042
rect 1159 1046 1163 1047
rect 1159 1041 1163 1042
rect 1175 1046 1179 1047
rect 1175 1041 1179 1042
rect 1223 1046 1227 1047
rect 1223 1041 1227 1042
rect 1239 1046 1243 1047
rect 1239 1041 1243 1042
rect 1279 1046 1283 1047
rect 1279 1041 1283 1042
rect 1303 1046 1307 1047
rect 1303 1041 1307 1042
rect 1335 1046 1339 1047
rect 1335 1041 1339 1042
rect 1359 1046 1363 1047
rect 1359 1041 1363 1042
rect 1383 1046 1387 1047
rect 1383 1041 1387 1042
rect 1415 1046 1419 1047
rect 1415 1041 1419 1042
rect 1431 1046 1435 1047
rect 1431 1041 1435 1042
rect 1463 1046 1467 1047
rect 1463 1041 1467 1042
rect 1479 1046 1483 1047
rect 1479 1041 1483 1042
rect 1503 1046 1507 1047
rect 1503 1041 1507 1042
rect 1535 1046 1539 1047
rect 1535 1041 1539 1042
rect 1551 1046 1555 1047
rect 1551 1041 1555 1042
rect 1591 1046 1595 1047
rect 1591 1041 1595 1042
rect 1623 1046 1627 1047
rect 1623 1041 1627 1042
rect 1663 1046 1667 1047
rect 1663 1041 1667 1042
rect 112 1033 114 1041
rect 110 1032 116 1033
rect 110 1028 111 1032
rect 115 1028 116 1032
rect 296 1031 298 1041
rect 328 1031 330 1041
rect 360 1031 362 1041
rect 392 1031 394 1041
rect 424 1031 426 1041
rect 456 1031 458 1041
rect 504 1031 506 1041
rect 560 1031 562 1041
rect 632 1031 634 1041
rect 712 1031 714 1041
rect 800 1031 802 1041
rect 880 1031 882 1041
rect 960 1031 962 1041
rect 1032 1031 1034 1041
rect 1096 1031 1098 1041
rect 1160 1031 1162 1041
rect 1224 1031 1226 1041
rect 1280 1031 1282 1041
rect 1336 1031 1338 1041
rect 1384 1031 1386 1041
rect 1432 1031 1434 1041
rect 1480 1031 1482 1041
rect 1536 1031 1538 1041
rect 1592 1031 1594 1041
rect 1624 1031 1626 1041
rect 1664 1033 1666 1041
rect 1662 1032 1668 1033
rect 110 1027 116 1028
rect 294 1030 300 1031
rect 294 1026 295 1030
rect 299 1026 300 1030
rect 294 1025 300 1026
rect 326 1030 332 1031
rect 326 1026 327 1030
rect 331 1026 332 1030
rect 326 1025 332 1026
rect 358 1030 364 1031
rect 358 1026 359 1030
rect 363 1026 364 1030
rect 358 1025 364 1026
rect 390 1030 396 1031
rect 390 1026 391 1030
rect 395 1026 396 1030
rect 390 1025 396 1026
rect 422 1030 428 1031
rect 422 1026 423 1030
rect 427 1026 428 1030
rect 422 1025 428 1026
rect 454 1030 460 1031
rect 454 1026 455 1030
rect 459 1026 460 1030
rect 454 1025 460 1026
rect 502 1030 508 1031
rect 502 1026 503 1030
rect 507 1026 508 1030
rect 502 1025 508 1026
rect 558 1030 564 1031
rect 558 1026 559 1030
rect 563 1026 564 1030
rect 558 1025 564 1026
rect 630 1030 636 1031
rect 630 1026 631 1030
rect 635 1026 636 1030
rect 630 1025 636 1026
rect 710 1030 716 1031
rect 710 1026 711 1030
rect 715 1026 716 1030
rect 710 1025 716 1026
rect 798 1030 804 1031
rect 798 1026 799 1030
rect 803 1026 804 1030
rect 798 1025 804 1026
rect 878 1030 884 1031
rect 878 1026 879 1030
rect 883 1026 884 1030
rect 878 1025 884 1026
rect 958 1030 964 1031
rect 958 1026 959 1030
rect 963 1026 964 1030
rect 958 1025 964 1026
rect 1030 1030 1036 1031
rect 1030 1026 1031 1030
rect 1035 1026 1036 1030
rect 1030 1025 1036 1026
rect 1094 1030 1100 1031
rect 1094 1026 1095 1030
rect 1099 1026 1100 1030
rect 1094 1025 1100 1026
rect 1158 1030 1164 1031
rect 1158 1026 1159 1030
rect 1163 1026 1164 1030
rect 1158 1025 1164 1026
rect 1222 1030 1228 1031
rect 1222 1026 1223 1030
rect 1227 1026 1228 1030
rect 1222 1025 1228 1026
rect 1278 1030 1284 1031
rect 1278 1026 1279 1030
rect 1283 1026 1284 1030
rect 1278 1025 1284 1026
rect 1334 1030 1340 1031
rect 1334 1026 1335 1030
rect 1339 1026 1340 1030
rect 1334 1025 1340 1026
rect 1382 1030 1388 1031
rect 1382 1026 1383 1030
rect 1387 1026 1388 1030
rect 1382 1025 1388 1026
rect 1430 1030 1436 1031
rect 1430 1026 1431 1030
rect 1435 1026 1436 1030
rect 1430 1025 1436 1026
rect 1478 1030 1484 1031
rect 1478 1026 1479 1030
rect 1483 1026 1484 1030
rect 1478 1025 1484 1026
rect 1534 1030 1540 1031
rect 1534 1026 1535 1030
rect 1539 1026 1540 1030
rect 1534 1025 1540 1026
rect 1590 1030 1596 1031
rect 1590 1026 1591 1030
rect 1595 1026 1596 1030
rect 1590 1025 1596 1026
rect 1622 1030 1628 1031
rect 1622 1026 1623 1030
rect 1627 1026 1628 1030
rect 1662 1028 1663 1032
rect 1667 1028 1668 1032
rect 1662 1027 1668 1028
rect 1622 1025 1628 1026
rect 110 1015 116 1016
rect 110 1011 111 1015
rect 115 1011 116 1015
rect 1662 1015 1668 1016
rect 110 1010 116 1011
rect 294 1013 300 1014
rect 112 1007 114 1010
rect 294 1009 295 1013
rect 299 1009 300 1013
rect 294 1008 300 1009
rect 326 1013 332 1014
rect 326 1009 327 1013
rect 331 1009 332 1013
rect 326 1008 332 1009
rect 358 1013 364 1014
rect 358 1009 359 1013
rect 363 1009 364 1013
rect 358 1008 364 1009
rect 390 1013 396 1014
rect 390 1009 391 1013
rect 395 1009 396 1013
rect 390 1008 396 1009
rect 422 1013 428 1014
rect 422 1009 423 1013
rect 427 1009 428 1013
rect 422 1008 428 1009
rect 454 1013 460 1014
rect 454 1009 455 1013
rect 459 1009 460 1013
rect 454 1008 460 1009
rect 502 1013 508 1014
rect 502 1009 503 1013
rect 507 1009 508 1013
rect 502 1008 508 1009
rect 558 1013 564 1014
rect 558 1009 559 1013
rect 563 1009 564 1013
rect 558 1008 564 1009
rect 630 1013 636 1014
rect 630 1009 631 1013
rect 635 1009 636 1013
rect 630 1008 636 1009
rect 710 1013 716 1014
rect 710 1009 711 1013
rect 715 1009 716 1013
rect 710 1008 716 1009
rect 798 1013 804 1014
rect 798 1009 799 1013
rect 803 1009 804 1013
rect 798 1008 804 1009
rect 878 1013 884 1014
rect 878 1009 879 1013
rect 883 1009 884 1013
rect 878 1008 884 1009
rect 958 1013 964 1014
rect 958 1009 959 1013
rect 963 1009 964 1013
rect 958 1008 964 1009
rect 1030 1013 1036 1014
rect 1030 1009 1031 1013
rect 1035 1009 1036 1013
rect 1030 1008 1036 1009
rect 1094 1013 1100 1014
rect 1094 1009 1095 1013
rect 1099 1009 1100 1013
rect 1094 1008 1100 1009
rect 1158 1013 1164 1014
rect 1158 1009 1159 1013
rect 1163 1009 1164 1013
rect 1158 1008 1164 1009
rect 1222 1013 1228 1014
rect 1222 1009 1223 1013
rect 1227 1009 1228 1013
rect 1222 1008 1228 1009
rect 1278 1013 1284 1014
rect 1278 1009 1279 1013
rect 1283 1009 1284 1013
rect 1278 1008 1284 1009
rect 1334 1013 1340 1014
rect 1334 1009 1335 1013
rect 1339 1009 1340 1013
rect 1334 1008 1340 1009
rect 1382 1013 1388 1014
rect 1382 1009 1383 1013
rect 1387 1009 1388 1013
rect 1382 1008 1388 1009
rect 1430 1013 1436 1014
rect 1430 1009 1431 1013
rect 1435 1009 1436 1013
rect 1430 1008 1436 1009
rect 1478 1013 1484 1014
rect 1478 1009 1479 1013
rect 1483 1009 1484 1013
rect 1478 1008 1484 1009
rect 1534 1013 1540 1014
rect 1534 1009 1535 1013
rect 1539 1009 1540 1013
rect 1534 1008 1540 1009
rect 1590 1013 1596 1014
rect 1590 1009 1591 1013
rect 1595 1009 1596 1013
rect 1590 1008 1596 1009
rect 1622 1013 1628 1014
rect 1622 1009 1623 1013
rect 1627 1009 1628 1013
rect 1662 1011 1663 1015
rect 1667 1011 1668 1015
rect 1662 1010 1668 1011
rect 1622 1008 1628 1009
rect 111 1006 115 1007
rect 111 1001 115 1002
rect 247 1006 251 1007
rect 112 998 114 1001
rect 247 1000 251 1002
rect 279 1006 283 1007
rect 279 1000 283 1002
rect 295 1006 299 1008
rect 295 1001 299 1002
rect 311 1006 315 1007
rect 311 1000 315 1002
rect 327 1006 331 1008
rect 327 1001 331 1002
rect 343 1006 347 1007
rect 343 1000 347 1002
rect 359 1006 363 1008
rect 359 1001 363 1002
rect 383 1006 387 1007
rect 383 1000 387 1002
rect 391 1006 395 1008
rect 391 1001 395 1002
rect 423 1006 427 1008
rect 423 1000 427 1002
rect 455 1006 459 1008
rect 455 1001 459 1002
rect 479 1006 483 1007
rect 479 1000 483 1002
rect 503 1006 507 1008
rect 503 1001 507 1002
rect 543 1006 547 1007
rect 543 1000 547 1002
rect 559 1006 563 1008
rect 559 1001 563 1002
rect 615 1006 619 1007
rect 615 1000 619 1002
rect 631 1006 635 1008
rect 631 1001 635 1002
rect 687 1006 691 1007
rect 687 1000 691 1002
rect 711 1006 715 1008
rect 711 1001 715 1002
rect 759 1006 763 1007
rect 759 1000 763 1002
rect 799 1006 803 1008
rect 799 1001 803 1002
rect 831 1006 835 1007
rect 831 1000 835 1002
rect 879 1006 883 1008
rect 879 1001 883 1002
rect 903 1006 907 1007
rect 903 1000 907 1002
rect 959 1006 963 1008
rect 959 1001 963 1002
rect 967 1006 971 1007
rect 967 1000 971 1002
rect 1031 1006 1035 1008
rect 1031 1000 1035 1002
rect 1095 1006 1099 1008
rect 1095 1000 1099 1002
rect 1159 1006 1163 1008
rect 1159 1000 1163 1002
rect 1223 1006 1227 1008
rect 1223 1000 1227 1002
rect 1279 1006 1283 1008
rect 1279 1001 1283 1002
rect 1287 1006 1291 1007
rect 1287 1000 1291 1002
rect 1335 1006 1339 1008
rect 1335 1001 1339 1002
rect 1343 1006 1347 1007
rect 1343 1000 1347 1002
rect 1383 1006 1387 1008
rect 1383 1001 1387 1002
rect 1399 1006 1403 1007
rect 1399 1000 1403 1002
rect 1431 1006 1435 1008
rect 1431 1001 1435 1002
rect 1447 1006 1451 1007
rect 1447 1000 1451 1002
rect 1479 1006 1483 1008
rect 1479 1001 1483 1002
rect 1495 1006 1499 1007
rect 1495 1000 1499 1002
rect 1535 1006 1539 1008
rect 1535 1001 1539 1002
rect 1543 1006 1547 1007
rect 1543 1000 1547 1002
rect 1591 1006 1595 1008
rect 1591 1000 1595 1002
rect 1623 1006 1627 1008
rect 1664 1007 1666 1010
rect 1623 1000 1627 1002
rect 1663 1006 1667 1007
rect 1663 1001 1667 1002
rect 246 999 252 1000
rect 110 997 116 998
rect 110 993 111 997
rect 115 993 116 997
rect 246 995 247 999
rect 251 995 252 999
rect 246 994 252 995
rect 278 999 284 1000
rect 278 995 279 999
rect 283 995 284 999
rect 278 994 284 995
rect 310 999 316 1000
rect 310 995 311 999
rect 315 995 316 999
rect 310 994 316 995
rect 342 999 348 1000
rect 342 995 343 999
rect 347 995 348 999
rect 342 994 348 995
rect 382 999 388 1000
rect 382 995 383 999
rect 387 995 388 999
rect 382 994 388 995
rect 422 999 428 1000
rect 422 995 423 999
rect 427 995 428 999
rect 422 994 428 995
rect 478 999 484 1000
rect 478 995 479 999
rect 483 995 484 999
rect 478 994 484 995
rect 542 999 548 1000
rect 542 995 543 999
rect 547 995 548 999
rect 542 994 548 995
rect 614 999 620 1000
rect 614 995 615 999
rect 619 995 620 999
rect 614 994 620 995
rect 686 999 692 1000
rect 686 995 687 999
rect 691 995 692 999
rect 686 994 692 995
rect 758 999 764 1000
rect 758 995 759 999
rect 763 995 764 999
rect 758 994 764 995
rect 830 999 836 1000
rect 830 995 831 999
rect 835 995 836 999
rect 830 994 836 995
rect 902 999 908 1000
rect 902 995 903 999
rect 907 995 908 999
rect 902 994 908 995
rect 966 999 972 1000
rect 966 995 967 999
rect 971 995 972 999
rect 966 994 972 995
rect 1030 999 1036 1000
rect 1030 995 1031 999
rect 1035 995 1036 999
rect 1030 994 1036 995
rect 1094 999 1100 1000
rect 1094 995 1095 999
rect 1099 995 1100 999
rect 1094 994 1100 995
rect 1158 999 1164 1000
rect 1158 995 1159 999
rect 1163 995 1164 999
rect 1158 994 1164 995
rect 1222 999 1228 1000
rect 1222 995 1223 999
rect 1227 995 1228 999
rect 1222 994 1228 995
rect 1286 999 1292 1000
rect 1286 995 1287 999
rect 1291 995 1292 999
rect 1286 994 1292 995
rect 1342 999 1348 1000
rect 1342 995 1343 999
rect 1347 995 1348 999
rect 1342 994 1348 995
rect 1398 999 1404 1000
rect 1398 995 1399 999
rect 1403 995 1404 999
rect 1398 994 1404 995
rect 1446 999 1452 1000
rect 1446 995 1447 999
rect 1451 995 1452 999
rect 1446 994 1452 995
rect 1494 999 1500 1000
rect 1494 995 1495 999
rect 1499 995 1500 999
rect 1494 994 1500 995
rect 1542 999 1548 1000
rect 1542 995 1543 999
rect 1547 995 1548 999
rect 1542 994 1548 995
rect 1590 999 1596 1000
rect 1590 995 1591 999
rect 1595 995 1596 999
rect 1590 994 1596 995
rect 1622 999 1628 1000
rect 1622 995 1623 999
rect 1627 995 1628 999
rect 1664 998 1666 1001
rect 1622 994 1628 995
rect 1662 997 1668 998
rect 110 992 116 993
rect 1662 993 1663 997
rect 1667 993 1668 997
rect 1662 992 1668 993
rect 246 982 252 983
rect 110 980 116 981
rect 110 976 111 980
rect 115 976 116 980
rect 246 978 247 982
rect 251 978 252 982
rect 246 977 252 978
rect 278 982 284 983
rect 278 978 279 982
rect 283 978 284 982
rect 278 977 284 978
rect 310 982 316 983
rect 310 978 311 982
rect 315 978 316 982
rect 310 977 316 978
rect 342 982 348 983
rect 342 978 343 982
rect 347 978 348 982
rect 342 977 348 978
rect 382 982 388 983
rect 382 978 383 982
rect 387 978 388 982
rect 382 977 388 978
rect 422 982 428 983
rect 422 978 423 982
rect 427 978 428 982
rect 422 977 428 978
rect 478 982 484 983
rect 478 978 479 982
rect 483 978 484 982
rect 478 977 484 978
rect 542 982 548 983
rect 542 978 543 982
rect 547 978 548 982
rect 542 977 548 978
rect 614 982 620 983
rect 614 978 615 982
rect 619 978 620 982
rect 614 977 620 978
rect 686 982 692 983
rect 686 978 687 982
rect 691 978 692 982
rect 686 977 692 978
rect 758 982 764 983
rect 758 978 759 982
rect 763 978 764 982
rect 758 977 764 978
rect 830 982 836 983
rect 830 978 831 982
rect 835 978 836 982
rect 830 977 836 978
rect 902 982 908 983
rect 902 978 903 982
rect 907 978 908 982
rect 902 977 908 978
rect 966 982 972 983
rect 966 978 967 982
rect 971 978 972 982
rect 966 977 972 978
rect 1030 982 1036 983
rect 1030 978 1031 982
rect 1035 978 1036 982
rect 1030 977 1036 978
rect 1094 982 1100 983
rect 1094 978 1095 982
rect 1099 978 1100 982
rect 1094 977 1100 978
rect 1158 982 1164 983
rect 1158 978 1159 982
rect 1163 978 1164 982
rect 1158 977 1164 978
rect 1222 982 1228 983
rect 1222 978 1223 982
rect 1227 978 1228 982
rect 1222 977 1228 978
rect 1286 982 1292 983
rect 1286 978 1287 982
rect 1291 978 1292 982
rect 1286 977 1292 978
rect 1342 982 1348 983
rect 1342 978 1343 982
rect 1347 978 1348 982
rect 1342 977 1348 978
rect 1398 982 1404 983
rect 1398 978 1399 982
rect 1403 978 1404 982
rect 1398 977 1404 978
rect 1446 982 1452 983
rect 1446 978 1447 982
rect 1451 978 1452 982
rect 1446 977 1452 978
rect 1494 982 1500 983
rect 1494 978 1495 982
rect 1499 978 1500 982
rect 1494 977 1500 978
rect 1542 982 1548 983
rect 1542 978 1543 982
rect 1547 978 1548 982
rect 1542 977 1548 978
rect 1590 982 1596 983
rect 1590 978 1591 982
rect 1595 978 1596 982
rect 1590 977 1596 978
rect 1622 982 1628 983
rect 1622 978 1623 982
rect 1627 978 1628 982
rect 1622 977 1628 978
rect 1662 980 1668 981
rect 110 975 116 976
rect 112 967 114 975
rect 248 967 250 977
rect 280 967 282 977
rect 312 967 314 977
rect 344 967 346 977
rect 384 967 386 977
rect 424 967 426 977
rect 480 967 482 977
rect 544 967 546 977
rect 616 967 618 977
rect 688 967 690 977
rect 760 967 762 977
rect 832 967 834 977
rect 904 967 906 977
rect 968 967 970 977
rect 1032 967 1034 977
rect 1096 967 1098 977
rect 1160 967 1162 977
rect 1224 967 1226 977
rect 1288 967 1290 977
rect 1344 967 1346 977
rect 1400 967 1402 977
rect 1448 967 1450 977
rect 1496 967 1498 977
rect 1544 967 1546 977
rect 1592 967 1594 977
rect 1624 967 1626 977
rect 1662 976 1663 980
rect 1667 976 1668 980
rect 1662 975 1668 976
rect 1664 967 1666 975
rect 111 966 115 967
rect 111 961 115 962
rect 167 966 171 967
rect 167 961 171 962
rect 199 966 203 967
rect 199 961 203 962
rect 239 966 243 967
rect 239 961 243 962
rect 247 966 251 967
rect 247 961 251 962
rect 279 966 283 967
rect 279 961 283 962
rect 287 966 291 967
rect 287 961 291 962
rect 311 966 315 967
rect 311 961 315 962
rect 343 966 347 967
rect 343 961 347 962
rect 383 966 387 967
rect 383 961 387 962
rect 407 966 411 967
rect 407 961 411 962
rect 423 966 427 967
rect 423 961 427 962
rect 471 966 475 967
rect 471 961 475 962
rect 479 966 483 967
rect 479 961 483 962
rect 535 966 539 967
rect 535 961 539 962
rect 543 966 547 967
rect 543 961 547 962
rect 599 966 603 967
rect 599 961 603 962
rect 615 966 619 967
rect 615 961 619 962
rect 663 966 667 967
rect 663 961 667 962
rect 687 966 691 967
rect 687 961 691 962
rect 727 966 731 967
rect 727 961 731 962
rect 759 966 763 967
rect 759 961 763 962
rect 791 966 795 967
rect 791 961 795 962
rect 831 966 835 967
rect 831 961 835 962
rect 847 966 851 967
rect 847 961 851 962
rect 903 966 907 967
rect 903 961 907 962
rect 911 966 915 967
rect 911 961 915 962
rect 967 966 971 967
rect 967 961 971 962
rect 975 966 979 967
rect 975 961 979 962
rect 1031 966 1035 967
rect 1031 961 1035 962
rect 1039 966 1043 967
rect 1039 961 1043 962
rect 1095 966 1099 967
rect 1095 961 1099 962
rect 1103 966 1107 967
rect 1103 961 1107 962
rect 1159 966 1163 967
rect 1159 961 1163 962
rect 1167 966 1171 967
rect 1167 961 1171 962
rect 1223 966 1227 967
rect 1223 961 1227 962
rect 1231 966 1235 967
rect 1231 961 1235 962
rect 1287 966 1291 967
rect 1287 961 1291 962
rect 1343 966 1347 967
rect 1343 961 1347 962
rect 1391 966 1395 967
rect 1391 961 1395 962
rect 1399 966 1403 967
rect 1399 961 1403 962
rect 1431 966 1435 967
rect 1431 961 1435 962
rect 1447 966 1451 967
rect 1447 961 1451 962
rect 1471 966 1475 967
rect 1471 961 1475 962
rect 1495 966 1499 967
rect 1495 961 1499 962
rect 1511 966 1515 967
rect 1511 961 1515 962
rect 1543 966 1547 967
rect 1543 961 1547 962
rect 1551 966 1555 967
rect 1551 961 1555 962
rect 1591 966 1595 967
rect 1591 961 1595 962
rect 1623 966 1627 967
rect 1623 961 1627 962
rect 1663 966 1667 967
rect 1663 961 1667 962
rect 112 953 114 961
rect 110 952 116 953
rect 110 948 111 952
rect 115 948 116 952
rect 168 951 170 961
rect 200 951 202 961
rect 240 951 242 961
rect 288 951 290 961
rect 344 951 346 961
rect 408 951 410 961
rect 472 951 474 961
rect 536 951 538 961
rect 600 951 602 961
rect 664 951 666 961
rect 728 951 730 961
rect 792 951 794 961
rect 848 951 850 961
rect 912 951 914 961
rect 976 951 978 961
rect 1040 951 1042 961
rect 1104 951 1106 961
rect 1168 951 1170 961
rect 1232 951 1234 961
rect 1288 951 1290 961
rect 1344 951 1346 961
rect 1392 951 1394 961
rect 1432 951 1434 961
rect 1472 951 1474 961
rect 1512 951 1514 961
rect 1552 951 1554 961
rect 1592 951 1594 961
rect 1624 951 1626 961
rect 1664 953 1666 961
rect 1662 952 1668 953
rect 110 947 116 948
rect 166 950 172 951
rect 166 946 167 950
rect 171 946 172 950
rect 166 945 172 946
rect 198 950 204 951
rect 198 946 199 950
rect 203 946 204 950
rect 198 945 204 946
rect 238 950 244 951
rect 238 946 239 950
rect 243 946 244 950
rect 238 945 244 946
rect 286 950 292 951
rect 286 946 287 950
rect 291 946 292 950
rect 286 945 292 946
rect 342 950 348 951
rect 342 946 343 950
rect 347 946 348 950
rect 342 945 348 946
rect 406 950 412 951
rect 406 946 407 950
rect 411 946 412 950
rect 406 945 412 946
rect 470 950 476 951
rect 470 946 471 950
rect 475 946 476 950
rect 470 945 476 946
rect 534 950 540 951
rect 534 946 535 950
rect 539 946 540 950
rect 534 945 540 946
rect 598 950 604 951
rect 598 946 599 950
rect 603 946 604 950
rect 598 945 604 946
rect 662 950 668 951
rect 662 946 663 950
rect 667 946 668 950
rect 662 945 668 946
rect 726 950 732 951
rect 726 946 727 950
rect 731 946 732 950
rect 726 945 732 946
rect 790 950 796 951
rect 790 946 791 950
rect 795 946 796 950
rect 790 945 796 946
rect 846 950 852 951
rect 846 946 847 950
rect 851 946 852 950
rect 846 945 852 946
rect 910 950 916 951
rect 910 946 911 950
rect 915 946 916 950
rect 910 945 916 946
rect 974 950 980 951
rect 974 946 975 950
rect 979 946 980 950
rect 974 945 980 946
rect 1038 950 1044 951
rect 1038 946 1039 950
rect 1043 946 1044 950
rect 1038 945 1044 946
rect 1102 950 1108 951
rect 1102 946 1103 950
rect 1107 946 1108 950
rect 1102 945 1108 946
rect 1166 950 1172 951
rect 1166 946 1167 950
rect 1171 946 1172 950
rect 1166 945 1172 946
rect 1230 950 1236 951
rect 1230 946 1231 950
rect 1235 946 1236 950
rect 1230 945 1236 946
rect 1286 950 1292 951
rect 1286 946 1287 950
rect 1291 946 1292 950
rect 1286 945 1292 946
rect 1342 950 1348 951
rect 1342 946 1343 950
rect 1347 946 1348 950
rect 1342 945 1348 946
rect 1390 950 1396 951
rect 1390 946 1391 950
rect 1395 946 1396 950
rect 1390 945 1396 946
rect 1430 950 1436 951
rect 1430 946 1431 950
rect 1435 946 1436 950
rect 1430 945 1436 946
rect 1470 950 1476 951
rect 1470 946 1471 950
rect 1475 946 1476 950
rect 1470 945 1476 946
rect 1510 950 1516 951
rect 1510 946 1511 950
rect 1515 946 1516 950
rect 1510 945 1516 946
rect 1550 950 1556 951
rect 1550 946 1551 950
rect 1555 946 1556 950
rect 1550 945 1556 946
rect 1590 950 1596 951
rect 1590 946 1591 950
rect 1595 946 1596 950
rect 1590 945 1596 946
rect 1622 950 1628 951
rect 1622 946 1623 950
rect 1627 946 1628 950
rect 1662 948 1663 952
rect 1667 948 1668 952
rect 1662 947 1668 948
rect 1622 945 1628 946
rect 110 935 116 936
rect 110 931 111 935
rect 115 931 116 935
rect 1662 935 1668 936
rect 110 930 116 931
rect 166 933 172 934
rect 112 923 114 930
rect 166 929 167 933
rect 171 929 172 933
rect 166 928 172 929
rect 198 933 204 934
rect 198 929 199 933
rect 203 929 204 933
rect 198 928 204 929
rect 238 933 244 934
rect 238 929 239 933
rect 243 929 244 933
rect 238 928 244 929
rect 286 933 292 934
rect 286 929 287 933
rect 291 929 292 933
rect 286 928 292 929
rect 342 933 348 934
rect 342 929 343 933
rect 347 929 348 933
rect 342 928 348 929
rect 406 933 412 934
rect 406 929 407 933
rect 411 929 412 933
rect 406 928 412 929
rect 470 933 476 934
rect 470 929 471 933
rect 475 929 476 933
rect 470 928 476 929
rect 534 933 540 934
rect 534 929 535 933
rect 539 929 540 933
rect 534 928 540 929
rect 598 933 604 934
rect 598 929 599 933
rect 603 929 604 933
rect 598 928 604 929
rect 662 933 668 934
rect 662 929 663 933
rect 667 929 668 933
rect 662 928 668 929
rect 726 933 732 934
rect 726 929 727 933
rect 731 929 732 933
rect 726 928 732 929
rect 790 933 796 934
rect 790 929 791 933
rect 795 929 796 933
rect 790 928 796 929
rect 846 933 852 934
rect 846 929 847 933
rect 851 929 852 933
rect 846 928 852 929
rect 910 933 916 934
rect 910 929 911 933
rect 915 929 916 933
rect 910 928 916 929
rect 974 933 980 934
rect 974 929 975 933
rect 979 929 980 933
rect 974 928 980 929
rect 1038 933 1044 934
rect 1038 929 1039 933
rect 1043 929 1044 933
rect 1038 928 1044 929
rect 1102 933 1108 934
rect 1102 929 1103 933
rect 1107 929 1108 933
rect 1102 928 1108 929
rect 1166 933 1172 934
rect 1166 929 1167 933
rect 1171 929 1172 933
rect 1166 928 1172 929
rect 1230 933 1236 934
rect 1230 929 1231 933
rect 1235 929 1236 933
rect 1230 928 1236 929
rect 1286 933 1292 934
rect 1286 929 1287 933
rect 1291 929 1292 933
rect 1286 928 1292 929
rect 1342 933 1348 934
rect 1342 929 1343 933
rect 1347 929 1348 933
rect 1342 928 1348 929
rect 1390 933 1396 934
rect 1390 929 1391 933
rect 1395 929 1396 933
rect 1390 928 1396 929
rect 1430 933 1436 934
rect 1430 929 1431 933
rect 1435 929 1436 933
rect 1430 928 1436 929
rect 1470 933 1476 934
rect 1470 929 1471 933
rect 1475 929 1476 933
rect 1470 928 1476 929
rect 1510 933 1516 934
rect 1510 929 1511 933
rect 1515 929 1516 933
rect 1510 928 1516 929
rect 1550 933 1556 934
rect 1550 929 1551 933
rect 1555 929 1556 933
rect 1550 928 1556 929
rect 1590 933 1596 934
rect 1590 929 1591 933
rect 1595 929 1596 933
rect 1590 928 1596 929
rect 1622 933 1628 934
rect 1622 929 1623 933
rect 1627 929 1628 933
rect 1662 931 1663 935
rect 1667 931 1668 935
rect 1662 930 1668 931
rect 1622 928 1628 929
rect 168 923 170 928
rect 200 923 202 928
rect 240 923 242 928
rect 288 923 290 928
rect 344 923 346 928
rect 408 923 410 928
rect 472 923 474 928
rect 536 923 538 928
rect 600 923 602 928
rect 664 923 666 928
rect 728 923 730 928
rect 792 923 794 928
rect 848 923 850 928
rect 912 923 914 928
rect 976 923 978 928
rect 1040 923 1042 928
rect 1104 923 1106 928
rect 1168 923 1170 928
rect 1232 923 1234 928
rect 1288 923 1290 928
rect 1344 923 1346 928
rect 1392 923 1394 928
rect 1432 923 1434 928
rect 1472 923 1474 928
rect 1512 923 1514 928
rect 1552 923 1554 928
rect 1592 923 1594 928
rect 1624 923 1626 928
rect 1664 923 1666 930
rect 111 922 115 923
rect 111 917 115 918
rect 135 922 139 923
rect 112 914 114 917
rect 135 916 139 918
rect 167 922 171 923
rect 167 916 171 918
rect 199 922 203 923
rect 199 917 203 918
rect 207 922 211 923
rect 207 916 211 918
rect 239 922 243 923
rect 239 917 243 918
rect 271 922 275 923
rect 271 916 275 918
rect 287 922 291 923
rect 287 917 291 918
rect 335 922 339 923
rect 335 916 339 918
rect 343 922 347 923
rect 343 917 347 918
rect 407 922 411 923
rect 407 916 411 918
rect 471 922 475 923
rect 471 916 475 918
rect 535 922 539 923
rect 535 916 539 918
rect 591 922 595 923
rect 591 916 595 918
rect 599 922 603 923
rect 599 917 603 918
rect 647 922 651 923
rect 647 916 651 918
rect 663 922 667 923
rect 663 917 667 918
rect 703 922 707 923
rect 703 916 707 918
rect 727 922 731 923
rect 727 917 731 918
rect 751 922 755 923
rect 751 916 755 918
rect 791 922 795 923
rect 791 917 795 918
rect 799 922 803 923
rect 799 916 803 918
rect 847 922 851 923
rect 847 916 851 918
rect 903 922 907 923
rect 903 916 907 918
rect 911 922 915 923
rect 911 917 915 918
rect 959 922 963 923
rect 959 916 963 918
rect 975 922 979 923
rect 975 917 979 918
rect 1023 922 1027 923
rect 1023 916 1027 918
rect 1039 922 1043 923
rect 1039 917 1043 918
rect 1087 922 1091 923
rect 1087 916 1091 918
rect 1103 922 1107 923
rect 1103 917 1107 918
rect 1143 922 1147 923
rect 1143 916 1147 918
rect 1167 922 1171 923
rect 1167 917 1171 918
rect 1199 922 1203 923
rect 1199 916 1203 918
rect 1231 922 1235 923
rect 1231 917 1235 918
rect 1255 922 1259 923
rect 1255 916 1259 918
rect 1287 922 1291 923
rect 1287 917 1291 918
rect 1319 922 1323 923
rect 1319 916 1323 918
rect 1343 922 1347 923
rect 1343 917 1347 918
rect 1383 922 1387 923
rect 1383 916 1387 918
rect 1391 922 1395 923
rect 1391 917 1395 918
rect 1431 922 1435 923
rect 1431 917 1435 918
rect 1471 922 1475 923
rect 1471 917 1475 918
rect 1511 922 1515 923
rect 1511 917 1515 918
rect 1551 922 1555 923
rect 1551 917 1555 918
rect 1591 922 1595 923
rect 1591 917 1595 918
rect 1623 922 1627 923
rect 1623 917 1627 918
rect 1663 922 1667 923
rect 1663 917 1667 918
rect 134 915 140 916
rect 110 913 116 914
rect 110 909 111 913
rect 115 909 116 913
rect 134 911 135 915
rect 139 911 140 915
rect 134 910 140 911
rect 166 915 172 916
rect 166 911 167 915
rect 171 911 172 915
rect 166 910 172 911
rect 206 915 212 916
rect 206 911 207 915
rect 211 911 212 915
rect 206 910 212 911
rect 270 915 276 916
rect 270 911 271 915
rect 275 911 276 915
rect 270 910 276 911
rect 334 915 340 916
rect 334 911 335 915
rect 339 911 340 915
rect 334 910 340 911
rect 406 915 412 916
rect 406 911 407 915
rect 411 911 412 915
rect 406 910 412 911
rect 470 915 476 916
rect 470 911 471 915
rect 475 911 476 915
rect 470 910 476 911
rect 534 915 540 916
rect 534 911 535 915
rect 539 911 540 915
rect 534 910 540 911
rect 590 915 596 916
rect 590 911 591 915
rect 595 911 596 915
rect 590 910 596 911
rect 646 915 652 916
rect 646 911 647 915
rect 651 911 652 915
rect 646 910 652 911
rect 702 915 708 916
rect 702 911 703 915
rect 707 911 708 915
rect 702 910 708 911
rect 750 915 756 916
rect 750 911 751 915
rect 755 911 756 915
rect 750 910 756 911
rect 798 915 804 916
rect 798 911 799 915
rect 803 911 804 915
rect 798 910 804 911
rect 846 915 852 916
rect 846 911 847 915
rect 851 911 852 915
rect 846 910 852 911
rect 902 915 908 916
rect 902 911 903 915
rect 907 911 908 915
rect 902 910 908 911
rect 958 915 964 916
rect 958 911 959 915
rect 963 911 964 915
rect 958 910 964 911
rect 1022 915 1028 916
rect 1022 911 1023 915
rect 1027 911 1028 915
rect 1022 910 1028 911
rect 1086 915 1092 916
rect 1086 911 1087 915
rect 1091 911 1092 915
rect 1086 910 1092 911
rect 1142 915 1148 916
rect 1142 911 1143 915
rect 1147 911 1148 915
rect 1142 910 1148 911
rect 1198 915 1204 916
rect 1198 911 1199 915
rect 1203 911 1204 915
rect 1198 910 1204 911
rect 1254 915 1260 916
rect 1254 911 1255 915
rect 1259 911 1260 915
rect 1254 910 1260 911
rect 1318 915 1324 916
rect 1318 911 1319 915
rect 1323 911 1324 915
rect 1318 910 1324 911
rect 1382 915 1388 916
rect 1382 911 1383 915
rect 1387 911 1388 915
rect 1664 914 1666 917
rect 1382 910 1388 911
rect 1662 913 1668 914
rect 110 908 116 909
rect 1662 909 1663 913
rect 1667 909 1668 913
rect 1662 908 1668 909
rect 134 898 140 899
rect 110 896 116 897
rect 110 892 111 896
rect 115 892 116 896
rect 134 894 135 898
rect 139 894 140 898
rect 134 893 140 894
rect 166 898 172 899
rect 166 894 167 898
rect 171 894 172 898
rect 166 893 172 894
rect 206 898 212 899
rect 206 894 207 898
rect 211 894 212 898
rect 206 893 212 894
rect 270 898 276 899
rect 270 894 271 898
rect 275 894 276 898
rect 270 893 276 894
rect 334 898 340 899
rect 334 894 335 898
rect 339 894 340 898
rect 334 893 340 894
rect 406 898 412 899
rect 406 894 407 898
rect 411 894 412 898
rect 406 893 412 894
rect 470 898 476 899
rect 470 894 471 898
rect 475 894 476 898
rect 470 893 476 894
rect 534 898 540 899
rect 534 894 535 898
rect 539 894 540 898
rect 534 893 540 894
rect 590 898 596 899
rect 590 894 591 898
rect 595 894 596 898
rect 590 893 596 894
rect 646 898 652 899
rect 646 894 647 898
rect 651 894 652 898
rect 646 893 652 894
rect 702 898 708 899
rect 702 894 703 898
rect 707 894 708 898
rect 702 893 708 894
rect 750 898 756 899
rect 750 894 751 898
rect 755 894 756 898
rect 750 893 756 894
rect 798 898 804 899
rect 798 894 799 898
rect 803 894 804 898
rect 798 893 804 894
rect 846 898 852 899
rect 846 894 847 898
rect 851 894 852 898
rect 846 893 852 894
rect 902 898 908 899
rect 902 894 903 898
rect 907 894 908 898
rect 902 893 908 894
rect 958 898 964 899
rect 958 894 959 898
rect 963 894 964 898
rect 958 893 964 894
rect 1022 898 1028 899
rect 1022 894 1023 898
rect 1027 894 1028 898
rect 1022 893 1028 894
rect 1086 898 1092 899
rect 1086 894 1087 898
rect 1091 894 1092 898
rect 1086 893 1092 894
rect 1142 898 1148 899
rect 1142 894 1143 898
rect 1147 894 1148 898
rect 1142 893 1148 894
rect 1198 898 1204 899
rect 1198 894 1199 898
rect 1203 894 1204 898
rect 1198 893 1204 894
rect 1254 898 1260 899
rect 1254 894 1255 898
rect 1259 894 1260 898
rect 1254 893 1260 894
rect 1318 898 1324 899
rect 1318 894 1319 898
rect 1323 894 1324 898
rect 1318 893 1324 894
rect 1382 898 1388 899
rect 1382 894 1383 898
rect 1387 894 1388 898
rect 1382 893 1388 894
rect 1662 896 1668 897
rect 110 891 116 892
rect 112 879 114 891
rect 136 879 138 893
rect 168 879 170 893
rect 208 879 210 893
rect 272 879 274 893
rect 336 879 338 893
rect 408 879 410 893
rect 472 879 474 893
rect 536 879 538 893
rect 592 879 594 893
rect 648 879 650 893
rect 704 879 706 893
rect 752 879 754 893
rect 800 879 802 893
rect 848 879 850 893
rect 904 879 906 893
rect 960 879 962 893
rect 1024 879 1026 893
rect 1088 879 1090 893
rect 1144 879 1146 893
rect 1200 879 1202 893
rect 1256 879 1258 893
rect 1320 879 1322 893
rect 1384 879 1386 893
rect 1662 892 1663 896
rect 1667 892 1668 896
rect 1662 891 1668 892
rect 1664 879 1666 891
rect 111 878 115 879
rect 111 873 115 874
rect 135 878 139 879
rect 135 873 139 874
rect 167 878 171 879
rect 167 873 171 874
rect 207 878 211 879
rect 207 873 211 874
rect 271 878 275 879
rect 271 873 275 874
rect 335 878 339 879
rect 335 873 339 874
rect 407 878 411 879
rect 407 873 411 874
rect 471 878 475 879
rect 471 873 475 874
rect 535 878 539 879
rect 535 873 539 874
rect 591 878 595 879
rect 591 873 595 874
rect 599 878 603 879
rect 599 873 603 874
rect 647 878 651 879
rect 647 873 651 874
rect 655 878 659 879
rect 655 873 659 874
rect 703 878 707 879
rect 703 873 707 874
rect 751 878 755 879
rect 751 873 755 874
rect 799 878 803 879
rect 799 873 803 874
rect 847 878 851 879
rect 847 873 851 874
rect 903 878 907 879
rect 903 873 907 874
rect 959 878 963 879
rect 959 873 963 874
rect 967 878 971 879
rect 967 873 971 874
rect 1023 878 1027 879
rect 1023 873 1027 874
rect 1039 878 1043 879
rect 1039 873 1043 874
rect 1087 878 1091 879
rect 1087 873 1091 874
rect 1103 878 1107 879
rect 1103 873 1107 874
rect 1143 878 1147 879
rect 1143 873 1147 874
rect 1167 878 1171 879
rect 1167 873 1171 874
rect 1199 878 1203 879
rect 1199 873 1203 874
rect 1231 878 1235 879
rect 1231 873 1235 874
rect 1255 878 1259 879
rect 1255 873 1259 874
rect 1287 878 1291 879
rect 1287 873 1291 874
rect 1319 878 1323 879
rect 1319 873 1323 874
rect 1343 878 1347 879
rect 1343 873 1347 874
rect 1383 878 1387 879
rect 1383 873 1387 874
rect 1399 878 1403 879
rect 1399 873 1403 874
rect 1463 878 1467 879
rect 1463 873 1467 874
rect 1663 878 1667 879
rect 1663 873 1667 874
rect 112 865 114 873
rect 110 864 116 865
rect 110 860 111 864
rect 115 860 116 864
rect 136 863 138 873
rect 168 863 170 873
rect 208 863 210 873
rect 272 863 274 873
rect 336 863 338 873
rect 408 863 410 873
rect 472 863 474 873
rect 536 863 538 873
rect 600 863 602 873
rect 656 863 658 873
rect 704 863 706 873
rect 752 863 754 873
rect 800 863 802 873
rect 848 863 850 873
rect 904 863 906 873
rect 968 863 970 873
rect 1040 863 1042 873
rect 1104 863 1106 873
rect 1168 863 1170 873
rect 1232 863 1234 873
rect 1288 863 1290 873
rect 1344 863 1346 873
rect 1400 863 1402 873
rect 1464 863 1466 873
rect 1664 865 1666 873
rect 1662 864 1668 865
rect 110 859 116 860
rect 134 862 140 863
rect 134 858 135 862
rect 139 858 140 862
rect 134 857 140 858
rect 166 862 172 863
rect 166 858 167 862
rect 171 858 172 862
rect 166 857 172 858
rect 206 862 212 863
rect 206 858 207 862
rect 211 858 212 862
rect 206 857 212 858
rect 270 862 276 863
rect 270 858 271 862
rect 275 858 276 862
rect 270 857 276 858
rect 334 862 340 863
rect 334 858 335 862
rect 339 858 340 862
rect 334 857 340 858
rect 406 862 412 863
rect 406 858 407 862
rect 411 858 412 862
rect 406 857 412 858
rect 470 862 476 863
rect 470 858 471 862
rect 475 858 476 862
rect 470 857 476 858
rect 534 862 540 863
rect 534 858 535 862
rect 539 858 540 862
rect 534 857 540 858
rect 598 862 604 863
rect 598 858 599 862
rect 603 858 604 862
rect 598 857 604 858
rect 654 862 660 863
rect 654 858 655 862
rect 659 858 660 862
rect 654 857 660 858
rect 702 862 708 863
rect 702 858 703 862
rect 707 858 708 862
rect 702 857 708 858
rect 750 862 756 863
rect 750 858 751 862
rect 755 858 756 862
rect 750 857 756 858
rect 798 862 804 863
rect 798 858 799 862
rect 803 858 804 862
rect 798 857 804 858
rect 846 862 852 863
rect 846 858 847 862
rect 851 858 852 862
rect 846 857 852 858
rect 902 862 908 863
rect 902 858 903 862
rect 907 858 908 862
rect 902 857 908 858
rect 966 862 972 863
rect 966 858 967 862
rect 971 858 972 862
rect 966 857 972 858
rect 1038 862 1044 863
rect 1038 858 1039 862
rect 1043 858 1044 862
rect 1038 857 1044 858
rect 1102 862 1108 863
rect 1102 858 1103 862
rect 1107 858 1108 862
rect 1102 857 1108 858
rect 1166 862 1172 863
rect 1166 858 1167 862
rect 1171 858 1172 862
rect 1166 857 1172 858
rect 1230 862 1236 863
rect 1230 858 1231 862
rect 1235 858 1236 862
rect 1230 857 1236 858
rect 1286 862 1292 863
rect 1286 858 1287 862
rect 1291 858 1292 862
rect 1286 857 1292 858
rect 1342 862 1348 863
rect 1342 858 1343 862
rect 1347 858 1348 862
rect 1342 857 1348 858
rect 1398 862 1404 863
rect 1398 858 1399 862
rect 1403 858 1404 862
rect 1398 857 1404 858
rect 1462 862 1468 863
rect 1462 858 1463 862
rect 1467 858 1468 862
rect 1662 860 1663 864
rect 1667 860 1668 864
rect 1662 859 1668 860
rect 1462 857 1468 858
rect 110 847 116 848
rect 110 843 111 847
rect 115 843 116 847
rect 1662 847 1668 848
rect 110 842 116 843
rect 134 845 140 846
rect 112 839 114 842
rect 134 841 135 845
rect 139 841 140 845
rect 134 840 140 841
rect 166 845 172 846
rect 166 841 167 845
rect 171 841 172 845
rect 166 840 172 841
rect 206 845 212 846
rect 206 841 207 845
rect 211 841 212 845
rect 206 840 212 841
rect 270 845 276 846
rect 270 841 271 845
rect 275 841 276 845
rect 270 840 276 841
rect 334 845 340 846
rect 334 841 335 845
rect 339 841 340 845
rect 334 840 340 841
rect 406 845 412 846
rect 406 841 407 845
rect 411 841 412 845
rect 406 840 412 841
rect 470 845 476 846
rect 470 841 471 845
rect 475 841 476 845
rect 470 840 476 841
rect 534 845 540 846
rect 534 841 535 845
rect 539 841 540 845
rect 534 840 540 841
rect 598 845 604 846
rect 598 841 599 845
rect 603 841 604 845
rect 598 840 604 841
rect 654 845 660 846
rect 654 841 655 845
rect 659 841 660 845
rect 654 840 660 841
rect 702 845 708 846
rect 702 841 703 845
rect 707 841 708 845
rect 702 840 708 841
rect 750 845 756 846
rect 750 841 751 845
rect 755 841 756 845
rect 750 840 756 841
rect 798 845 804 846
rect 798 841 799 845
rect 803 841 804 845
rect 798 840 804 841
rect 846 845 852 846
rect 846 841 847 845
rect 851 841 852 845
rect 846 840 852 841
rect 902 845 908 846
rect 902 841 903 845
rect 907 841 908 845
rect 902 840 908 841
rect 966 845 972 846
rect 966 841 967 845
rect 971 841 972 845
rect 966 840 972 841
rect 1038 845 1044 846
rect 1038 841 1039 845
rect 1043 841 1044 845
rect 1038 840 1044 841
rect 1102 845 1108 846
rect 1102 841 1103 845
rect 1107 841 1108 845
rect 1102 840 1108 841
rect 1166 845 1172 846
rect 1166 841 1167 845
rect 1171 841 1172 845
rect 1166 840 1172 841
rect 1230 845 1236 846
rect 1230 841 1231 845
rect 1235 841 1236 845
rect 1230 840 1236 841
rect 1286 845 1292 846
rect 1286 841 1287 845
rect 1291 841 1292 845
rect 1286 840 1292 841
rect 1342 845 1348 846
rect 1342 841 1343 845
rect 1347 841 1348 845
rect 1342 840 1348 841
rect 1398 845 1404 846
rect 1398 841 1399 845
rect 1403 841 1404 845
rect 1398 840 1404 841
rect 1462 845 1468 846
rect 1462 841 1463 845
rect 1467 841 1468 845
rect 1662 843 1663 847
rect 1667 843 1668 847
rect 1662 842 1668 843
rect 1462 840 1468 841
rect 111 838 115 839
rect 111 833 115 834
rect 135 838 139 840
rect 112 830 114 833
rect 135 832 139 834
rect 167 838 171 840
rect 167 832 171 834
rect 207 838 211 840
rect 207 833 211 834
rect 215 838 219 839
rect 215 832 219 834
rect 271 838 275 840
rect 271 833 275 834
rect 279 838 283 839
rect 279 832 283 834
rect 335 838 339 840
rect 335 833 339 834
rect 343 838 347 839
rect 343 832 347 834
rect 407 838 411 840
rect 407 833 411 834
rect 415 838 419 839
rect 415 832 419 834
rect 471 838 475 840
rect 471 833 475 834
rect 479 838 483 839
rect 479 832 483 834
rect 535 838 539 840
rect 535 833 539 834
rect 543 838 547 839
rect 543 832 547 834
rect 599 838 603 840
rect 599 833 603 834
rect 607 838 611 839
rect 607 832 611 834
rect 655 838 659 840
rect 655 833 659 834
rect 671 838 675 839
rect 671 832 675 834
rect 703 838 707 840
rect 703 833 707 834
rect 735 838 739 839
rect 735 832 739 834
rect 751 838 755 840
rect 751 833 755 834
rect 791 838 795 839
rect 791 832 795 834
rect 799 838 803 840
rect 799 833 803 834
rect 847 838 851 840
rect 847 832 851 834
rect 903 838 907 840
rect 903 833 907 834
rect 911 838 915 839
rect 911 832 915 834
rect 967 838 971 840
rect 967 833 971 834
rect 975 838 979 839
rect 975 832 979 834
rect 1039 838 1043 840
rect 1039 832 1043 834
rect 1103 838 1107 840
rect 1103 833 1107 834
rect 1111 838 1115 839
rect 1111 832 1115 834
rect 1167 838 1171 840
rect 1167 833 1171 834
rect 1183 838 1187 839
rect 1183 832 1187 834
rect 1231 838 1235 840
rect 1231 833 1235 834
rect 1247 838 1251 839
rect 1247 832 1251 834
rect 1287 838 1291 840
rect 1287 833 1291 834
rect 1311 838 1315 839
rect 1311 832 1315 834
rect 1343 838 1347 840
rect 1343 833 1347 834
rect 1367 838 1371 839
rect 1367 832 1371 834
rect 1399 838 1403 840
rect 1399 833 1403 834
rect 1423 838 1427 839
rect 1423 832 1427 834
rect 1463 838 1467 840
rect 1664 839 1666 842
rect 1463 833 1467 834
rect 1479 838 1483 839
rect 1479 832 1483 834
rect 1535 838 1539 839
rect 1535 832 1539 834
rect 1591 838 1595 839
rect 1591 832 1595 834
rect 1663 838 1667 839
rect 1663 833 1667 834
rect 134 831 140 832
rect 110 829 116 830
rect 110 825 111 829
rect 115 825 116 829
rect 134 827 135 831
rect 139 827 140 831
rect 134 826 140 827
rect 166 831 172 832
rect 166 827 167 831
rect 171 827 172 831
rect 166 826 172 827
rect 214 831 220 832
rect 214 827 215 831
rect 219 827 220 831
rect 214 826 220 827
rect 278 831 284 832
rect 278 827 279 831
rect 283 827 284 831
rect 278 826 284 827
rect 342 831 348 832
rect 342 827 343 831
rect 347 827 348 831
rect 342 826 348 827
rect 414 831 420 832
rect 414 827 415 831
rect 419 827 420 831
rect 414 826 420 827
rect 478 831 484 832
rect 478 827 479 831
rect 483 827 484 831
rect 478 826 484 827
rect 542 831 548 832
rect 542 827 543 831
rect 547 827 548 831
rect 542 826 548 827
rect 606 831 612 832
rect 606 827 607 831
rect 611 827 612 831
rect 606 826 612 827
rect 670 831 676 832
rect 670 827 671 831
rect 675 827 676 831
rect 670 826 676 827
rect 734 831 740 832
rect 734 827 735 831
rect 739 827 740 831
rect 734 826 740 827
rect 790 831 796 832
rect 790 827 791 831
rect 795 827 796 831
rect 790 826 796 827
rect 846 831 852 832
rect 846 827 847 831
rect 851 827 852 831
rect 846 826 852 827
rect 910 831 916 832
rect 910 827 911 831
rect 915 827 916 831
rect 910 826 916 827
rect 974 831 980 832
rect 974 827 975 831
rect 979 827 980 831
rect 974 826 980 827
rect 1038 831 1044 832
rect 1038 827 1039 831
rect 1043 827 1044 831
rect 1038 826 1044 827
rect 1110 831 1116 832
rect 1110 827 1111 831
rect 1115 827 1116 831
rect 1110 826 1116 827
rect 1182 831 1188 832
rect 1182 827 1183 831
rect 1187 827 1188 831
rect 1182 826 1188 827
rect 1246 831 1252 832
rect 1246 827 1247 831
rect 1251 827 1252 831
rect 1246 826 1252 827
rect 1310 831 1316 832
rect 1310 827 1311 831
rect 1315 827 1316 831
rect 1310 826 1316 827
rect 1366 831 1372 832
rect 1366 827 1367 831
rect 1371 827 1372 831
rect 1366 826 1372 827
rect 1422 831 1428 832
rect 1422 827 1423 831
rect 1427 827 1428 831
rect 1422 826 1428 827
rect 1478 831 1484 832
rect 1478 827 1479 831
rect 1483 827 1484 831
rect 1478 826 1484 827
rect 1534 831 1540 832
rect 1534 827 1535 831
rect 1539 827 1540 831
rect 1534 826 1540 827
rect 1590 831 1596 832
rect 1590 827 1591 831
rect 1595 827 1596 831
rect 1664 830 1666 833
rect 1590 826 1596 827
rect 1662 829 1668 830
rect 110 824 116 825
rect 1662 825 1663 829
rect 1667 825 1668 829
rect 1662 824 1668 825
rect 134 814 140 815
rect 110 812 116 813
rect 110 808 111 812
rect 115 808 116 812
rect 134 810 135 814
rect 139 810 140 814
rect 134 809 140 810
rect 166 814 172 815
rect 166 810 167 814
rect 171 810 172 814
rect 166 809 172 810
rect 214 814 220 815
rect 214 810 215 814
rect 219 810 220 814
rect 214 809 220 810
rect 278 814 284 815
rect 278 810 279 814
rect 283 810 284 814
rect 278 809 284 810
rect 342 814 348 815
rect 342 810 343 814
rect 347 810 348 814
rect 342 809 348 810
rect 414 814 420 815
rect 414 810 415 814
rect 419 810 420 814
rect 414 809 420 810
rect 478 814 484 815
rect 478 810 479 814
rect 483 810 484 814
rect 478 809 484 810
rect 542 814 548 815
rect 542 810 543 814
rect 547 810 548 814
rect 542 809 548 810
rect 606 814 612 815
rect 606 810 607 814
rect 611 810 612 814
rect 606 809 612 810
rect 670 814 676 815
rect 670 810 671 814
rect 675 810 676 814
rect 670 809 676 810
rect 734 814 740 815
rect 734 810 735 814
rect 739 810 740 814
rect 734 809 740 810
rect 790 814 796 815
rect 790 810 791 814
rect 795 810 796 814
rect 790 809 796 810
rect 846 814 852 815
rect 846 810 847 814
rect 851 810 852 814
rect 846 809 852 810
rect 910 814 916 815
rect 910 810 911 814
rect 915 810 916 814
rect 910 809 916 810
rect 974 814 980 815
rect 974 810 975 814
rect 979 810 980 814
rect 974 809 980 810
rect 1038 814 1044 815
rect 1038 810 1039 814
rect 1043 810 1044 814
rect 1038 809 1044 810
rect 1110 814 1116 815
rect 1110 810 1111 814
rect 1115 810 1116 814
rect 1110 809 1116 810
rect 1182 814 1188 815
rect 1182 810 1183 814
rect 1187 810 1188 814
rect 1182 809 1188 810
rect 1246 814 1252 815
rect 1246 810 1247 814
rect 1251 810 1252 814
rect 1246 809 1252 810
rect 1310 814 1316 815
rect 1310 810 1311 814
rect 1315 810 1316 814
rect 1310 809 1316 810
rect 1366 814 1372 815
rect 1366 810 1367 814
rect 1371 810 1372 814
rect 1366 809 1372 810
rect 1422 814 1428 815
rect 1422 810 1423 814
rect 1427 810 1428 814
rect 1422 809 1428 810
rect 1478 814 1484 815
rect 1478 810 1479 814
rect 1483 810 1484 814
rect 1478 809 1484 810
rect 1534 814 1540 815
rect 1534 810 1535 814
rect 1539 810 1540 814
rect 1534 809 1540 810
rect 1590 814 1596 815
rect 1590 810 1591 814
rect 1595 810 1596 814
rect 1590 809 1596 810
rect 1662 812 1668 813
rect 110 807 116 808
rect 112 795 114 807
rect 136 795 138 809
rect 168 795 170 809
rect 216 795 218 809
rect 280 795 282 809
rect 344 795 346 809
rect 416 795 418 809
rect 480 795 482 809
rect 544 795 546 809
rect 608 795 610 809
rect 672 795 674 809
rect 736 795 738 809
rect 792 795 794 809
rect 848 795 850 809
rect 912 795 914 809
rect 976 795 978 809
rect 1040 795 1042 809
rect 1112 795 1114 809
rect 1184 795 1186 809
rect 1248 795 1250 809
rect 1312 795 1314 809
rect 1368 795 1370 809
rect 1424 795 1426 809
rect 1480 795 1482 809
rect 1536 795 1538 809
rect 1592 795 1594 809
rect 1662 808 1663 812
rect 1667 808 1668 812
rect 1662 807 1668 808
rect 1664 795 1666 807
rect 111 794 115 795
rect 111 789 115 790
rect 135 794 139 795
rect 135 789 139 790
rect 167 794 171 795
rect 167 789 171 790
rect 175 794 179 795
rect 175 789 179 790
rect 215 794 219 795
rect 215 789 219 790
rect 231 794 235 795
rect 231 789 235 790
rect 279 794 283 795
rect 279 789 283 790
rect 295 794 299 795
rect 295 789 299 790
rect 343 794 347 795
rect 343 789 347 790
rect 367 794 371 795
rect 367 789 371 790
rect 415 794 419 795
rect 415 789 419 790
rect 447 794 451 795
rect 447 789 451 790
rect 479 794 483 795
rect 479 789 483 790
rect 527 794 531 795
rect 527 789 531 790
rect 543 794 547 795
rect 543 789 547 790
rect 607 794 611 795
rect 607 789 611 790
rect 615 794 619 795
rect 615 789 619 790
rect 671 794 675 795
rect 671 789 675 790
rect 703 794 707 795
rect 703 789 707 790
rect 735 794 739 795
rect 735 789 739 790
rect 791 794 795 795
rect 791 789 795 790
rect 847 794 851 795
rect 847 789 851 790
rect 871 794 875 795
rect 871 789 875 790
rect 911 794 915 795
rect 911 789 915 790
rect 951 794 955 795
rect 951 789 955 790
rect 975 794 979 795
rect 975 789 979 790
rect 1023 794 1027 795
rect 1023 789 1027 790
rect 1039 794 1043 795
rect 1039 789 1043 790
rect 1095 794 1099 795
rect 1095 789 1099 790
rect 1111 794 1115 795
rect 1111 789 1115 790
rect 1167 794 1171 795
rect 1167 789 1171 790
rect 1183 794 1187 795
rect 1183 789 1187 790
rect 1231 794 1235 795
rect 1231 789 1235 790
rect 1247 794 1251 795
rect 1247 789 1251 790
rect 1295 794 1299 795
rect 1295 789 1299 790
rect 1311 794 1315 795
rect 1311 789 1315 790
rect 1359 794 1363 795
rect 1359 789 1363 790
rect 1367 794 1371 795
rect 1367 789 1371 790
rect 1415 794 1419 795
rect 1415 789 1419 790
rect 1423 794 1427 795
rect 1423 789 1427 790
rect 1471 794 1475 795
rect 1471 789 1475 790
rect 1479 794 1483 795
rect 1479 789 1483 790
rect 1527 794 1531 795
rect 1527 789 1531 790
rect 1535 794 1539 795
rect 1535 789 1539 790
rect 1591 794 1595 795
rect 1591 789 1595 790
rect 1663 794 1667 795
rect 1663 789 1667 790
rect 112 781 114 789
rect 110 780 116 781
rect 110 776 111 780
rect 115 776 116 780
rect 136 779 138 789
rect 176 779 178 789
rect 232 779 234 789
rect 296 779 298 789
rect 368 779 370 789
rect 448 779 450 789
rect 528 779 530 789
rect 616 779 618 789
rect 704 779 706 789
rect 792 779 794 789
rect 872 779 874 789
rect 952 779 954 789
rect 1024 779 1026 789
rect 1096 779 1098 789
rect 1168 779 1170 789
rect 1232 779 1234 789
rect 1296 779 1298 789
rect 1360 779 1362 789
rect 1416 779 1418 789
rect 1472 779 1474 789
rect 1528 779 1530 789
rect 1592 779 1594 789
rect 1664 781 1666 789
rect 1662 780 1668 781
rect 110 775 116 776
rect 134 778 140 779
rect 134 774 135 778
rect 139 774 140 778
rect 134 773 140 774
rect 174 778 180 779
rect 174 774 175 778
rect 179 774 180 778
rect 174 773 180 774
rect 230 778 236 779
rect 230 774 231 778
rect 235 774 236 778
rect 230 773 236 774
rect 294 778 300 779
rect 294 774 295 778
rect 299 774 300 778
rect 294 773 300 774
rect 366 778 372 779
rect 366 774 367 778
rect 371 774 372 778
rect 366 773 372 774
rect 446 778 452 779
rect 446 774 447 778
rect 451 774 452 778
rect 446 773 452 774
rect 526 778 532 779
rect 526 774 527 778
rect 531 774 532 778
rect 526 773 532 774
rect 614 778 620 779
rect 614 774 615 778
rect 619 774 620 778
rect 614 773 620 774
rect 702 778 708 779
rect 702 774 703 778
rect 707 774 708 778
rect 702 773 708 774
rect 790 778 796 779
rect 790 774 791 778
rect 795 774 796 778
rect 790 773 796 774
rect 870 778 876 779
rect 870 774 871 778
rect 875 774 876 778
rect 870 773 876 774
rect 950 778 956 779
rect 950 774 951 778
rect 955 774 956 778
rect 950 773 956 774
rect 1022 778 1028 779
rect 1022 774 1023 778
rect 1027 774 1028 778
rect 1022 773 1028 774
rect 1094 778 1100 779
rect 1094 774 1095 778
rect 1099 774 1100 778
rect 1094 773 1100 774
rect 1166 778 1172 779
rect 1166 774 1167 778
rect 1171 774 1172 778
rect 1166 773 1172 774
rect 1230 778 1236 779
rect 1230 774 1231 778
rect 1235 774 1236 778
rect 1230 773 1236 774
rect 1294 778 1300 779
rect 1294 774 1295 778
rect 1299 774 1300 778
rect 1294 773 1300 774
rect 1358 778 1364 779
rect 1358 774 1359 778
rect 1363 774 1364 778
rect 1358 773 1364 774
rect 1414 778 1420 779
rect 1414 774 1415 778
rect 1419 774 1420 778
rect 1414 773 1420 774
rect 1470 778 1476 779
rect 1470 774 1471 778
rect 1475 774 1476 778
rect 1470 773 1476 774
rect 1526 778 1532 779
rect 1526 774 1527 778
rect 1531 774 1532 778
rect 1526 773 1532 774
rect 1590 778 1596 779
rect 1590 774 1591 778
rect 1595 774 1596 778
rect 1662 776 1663 780
rect 1667 776 1668 780
rect 1662 775 1668 776
rect 1590 773 1596 774
rect 110 763 116 764
rect 110 759 111 763
rect 115 759 116 763
rect 1662 763 1668 764
rect 110 758 116 759
rect 134 761 140 762
rect 112 755 114 758
rect 134 757 135 761
rect 139 757 140 761
rect 134 756 140 757
rect 174 761 180 762
rect 174 757 175 761
rect 179 757 180 761
rect 174 756 180 757
rect 230 761 236 762
rect 230 757 231 761
rect 235 757 236 761
rect 230 756 236 757
rect 294 761 300 762
rect 294 757 295 761
rect 299 757 300 761
rect 294 756 300 757
rect 366 761 372 762
rect 366 757 367 761
rect 371 757 372 761
rect 366 756 372 757
rect 446 761 452 762
rect 446 757 447 761
rect 451 757 452 761
rect 446 756 452 757
rect 526 761 532 762
rect 526 757 527 761
rect 531 757 532 761
rect 526 756 532 757
rect 614 761 620 762
rect 614 757 615 761
rect 619 757 620 761
rect 614 756 620 757
rect 702 761 708 762
rect 702 757 703 761
rect 707 757 708 761
rect 702 756 708 757
rect 790 761 796 762
rect 790 757 791 761
rect 795 757 796 761
rect 790 756 796 757
rect 870 761 876 762
rect 870 757 871 761
rect 875 757 876 761
rect 870 756 876 757
rect 950 761 956 762
rect 950 757 951 761
rect 955 757 956 761
rect 950 756 956 757
rect 1022 761 1028 762
rect 1022 757 1023 761
rect 1027 757 1028 761
rect 1022 756 1028 757
rect 1094 761 1100 762
rect 1094 757 1095 761
rect 1099 757 1100 761
rect 1094 756 1100 757
rect 1166 761 1172 762
rect 1166 757 1167 761
rect 1171 757 1172 761
rect 1166 756 1172 757
rect 1230 761 1236 762
rect 1230 757 1231 761
rect 1235 757 1236 761
rect 1230 756 1236 757
rect 1294 761 1300 762
rect 1294 757 1295 761
rect 1299 757 1300 761
rect 1294 756 1300 757
rect 1358 761 1364 762
rect 1358 757 1359 761
rect 1363 757 1364 761
rect 1358 756 1364 757
rect 1414 761 1420 762
rect 1414 757 1415 761
rect 1419 757 1420 761
rect 1414 756 1420 757
rect 1470 761 1476 762
rect 1470 757 1471 761
rect 1475 757 1476 761
rect 1470 756 1476 757
rect 1526 761 1532 762
rect 1526 757 1527 761
rect 1531 757 1532 761
rect 1526 756 1532 757
rect 1590 761 1596 762
rect 1590 757 1591 761
rect 1595 757 1596 761
rect 1662 759 1663 763
rect 1667 759 1668 763
rect 1662 758 1668 759
rect 1590 756 1596 757
rect 111 754 115 755
rect 111 749 115 750
rect 135 754 139 756
rect 135 749 139 750
rect 175 754 179 756
rect 175 749 179 750
rect 215 754 219 755
rect 112 746 114 749
rect 215 748 219 750
rect 231 754 235 756
rect 231 749 235 750
rect 247 754 251 755
rect 247 748 251 750
rect 279 754 283 755
rect 279 748 283 750
rect 295 754 299 756
rect 295 749 299 750
rect 319 754 323 755
rect 319 748 323 750
rect 359 754 363 755
rect 359 748 363 750
rect 367 754 371 756
rect 367 749 371 750
rect 399 754 403 755
rect 399 748 403 750
rect 439 754 443 755
rect 439 748 443 750
rect 447 754 451 756
rect 447 749 451 750
rect 487 754 491 755
rect 487 748 491 750
rect 527 754 531 756
rect 527 749 531 750
rect 543 754 547 755
rect 543 748 547 750
rect 607 754 611 755
rect 607 748 611 750
rect 615 754 619 756
rect 615 749 619 750
rect 671 754 675 755
rect 671 748 675 750
rect 703 754 707 756
rect 703 749 707 750
rect 735 754 739 755
rect 735 748 739 750
rect 791 754 795 756
rect 791 749 795 750
rect 799 754 803 755
rect 799 748 803 750
rect 863 754 867 755
rect 863 748 867 750
rect 871 754 875 756
rect 871 749 875 750
rect 927 754 931 755
rect 927 748 931 750
rect 951 754 955 756
rect 951 749 955 750
rect 991 754 995 755
rect 991 748 995 750
rect 1023 754 1027 756
rect 1023 749 1027 750
rect 1055 754 1059 755
rect 1055 748 1059 750
rect 1095 754 1099 756
rect 1095 749 1099 750
rect 1119 754 1123 755
rect 1119 748 1123 750
rect 1167 754 1171 756
rect 1167 749 1171 750
rect 1183 754 1187 755
rect 1183 748 1187 750
rect 1231 754 1235 756
rect 1231 749 1235 750
rect 1239 754 1243 755
rect 1239 748 1243 750
rect 1295 754 1299 756
rect 1295 748 1299 750
rect 1351 754 1355 755
rect 1351 748 1355 750
rect 1359 754 1363 756
rect 1359 749 1363 750
rect 1407 754 1411 755
rect 1407 748 1411 750
rect 1415 754 1419 756
rect 1415 749 1419 750
rect 1463 754 1467 755
rect 1463 748 1467 750
rect 1471 754 1475 756
rect 1471 749 1475 750
rect 1519 754 1523 755
rect 1519 748 1523 750
rect 1527 754 1531 756
rect 1527 749 1531 750
rect 1583 754 1587 755
rect 1583 748 1587 750
rect 1591 754 1595 756
rect 1664 755 1666 758
rect 1591 749 1595 750
rect 1623 754 1627 755
rect 1623 748 1627 750
rect 1663 754 1667 755
rect 1663 749 1667 750
rect 214 747 220 748
rect 110 745 116 746
rect 110 741 111 745
rect 115 741 116 745
rect 214 743 215 747
rect 219 743 220 747
rect 214 742 220 743
rect 246 747 252 748
rect 246 743 247 747
rect 251 743 252 747
rect 246 742 252 743
rect 278 747 284 748
rect 278 743 279 747
rect 283 743 284 747
rect 278 742 284 743
rect 318 747 324 748
rect 318 743 319 747
rect 323 743 324 747
rect 318 742 324 743
rect 358 747 364 748
rect 358 743 359 747
rect 363 743 364 747
rect 358 742 364 743
rect 398 747 404 748
rect 398 743 399 747
rect 403 743 404 747
rect 398 742 404 743
rect 438 747 444 748
rect 438 743 439 747
rect 443 743 444 747
rect 438 742 444 743
rect 486 747 492 748
rect 486 743 487 747
rect 491 743 492 747
rect 486 742 492 743
rect 542 747 548 748
rect 542 743 543 747
rect 547 743 548 747
rect 542 742 548 743
rect 606 747 612 748
rect 606 743 607 747
rect 611 743 612 747
rect 606 742 612 743
rect 670 747 676 748
rect 670 743 671 747
rect 675 743 676 747
rect 670 742 676 743
rect 734 747 740 748
rect 734 743 735 747
rect 739 743 740 747
rect 734 742 740 743
rect 798 747 804 748
rect 798 743 799 747
rect 803 743 804 747
rect 798 742 804 743
rect 862 747 868 748
rect 862 743 863 747
rect 867 743 868 747
rect 862 742 868 743
rect 926 747 932 748
rect 926 743 927 747
rect 931 743 932 747
rect 926 742 932 743
rect 990 747 996 748
rect 990 743 991 747
rect 995 743 996 747
rect 990 742 996 743
rect 1054 747 1060 748
rect 1054 743 1055 747
rect 1059 743 1060 747
rect 1054 742 1060 743
rect 1118 747 1124 748
rect 1118 743 1119 747
rect 1123 743 1124 747
rect 1118 742 1124 743
rect 1182 747 1188 748
rect 1182 743 1183 747
rect 1187 743 1188 747
rect 1182 742 1188 743
rect 1238 747 1244 748
rect 1238 743 1239 747
rect 1243 743 1244 747
rect 1238 742 1244 743
rect 1294 747 1300 748
rect 1294 743 1295 747
rect 1299 743 1300 747
rect 1294 742 1300 743
rect 1350 747 1356 748
rect 1350 743 1351 747
rect 1355 743 1356 747
rect 1350 742 1356 743
rect 1406 747 1412 748
rect 1406 743 1407 747
rect 1411 743 1412 747
rect 1406 742 1412 743
rect 1462 747 1468 748
rect 1462 743 1463 747
rect 1467 743 1468 747
rect 1462 742 1468 743
rect 1518 747 1524 748
rect 1518 743 1519 747
rect 1523 743 1524 747
rect 1518 742 1524 743
rect 1582 747 1588 748
rect 1582 743 1583 747
rect 1587 743 1588 747
rect 1582 742 1588 743
rect 1622 747 1628 748
rect 1622 743 1623 747
rect 1627 743 1628 747
rect 1664 746 1666 749
rect 1622 742 1628 743
rect 1662 745 1668 746
rect 110 740 116 741
rect 1662 741 1663 745
rect 1667 741 1668 745
rect 1662 740 1668 741
rect 214 730 220 731
rect 110 728 116 729
rect 110 724 111 728
rect 115 724 116 728
rect 214 726 215 730
rect 219 726 220 730
rect 214 725 220 726
rect 246 730 252 731
rect 246 726 247 730
rect 251 726 252 730
rect 246 725 252 726
rect 278 730 284 731
rect 278 726 279 730
rect 283 726 284 730
rect 278 725 284 726
rect 318 730 324 731
rect 318 726 319 730
rect 323 726 324 730
rect 318 725 324 726
rect 358 730 364 731
rect 358 726 359 730
rect 363 726 364 730
rect 358 725 364 726
rect 398 730 404 731
rect 398 726 399 730
rect 403 726 404 730
rect 398 725 404 726
rect 438 730 444 731
rect 438 726 439 730
rect 443 726 444 730
rect 438 725 444 726
rect 486 730 492 731
rect 486 726 487 730
rect 491 726 492 730
rect 486 725 492 726
rect 542 730 548 731
rect 542 726 543 730
rect 547 726 548 730
rect 542 725 548 726
rect 606 730 612 731
rect 606 726 607 730
rect 611 726 612 730
rect 606 725 612 726
rect 670 730 676 731
rect 670 726 671 730
rect 675 726 676 730
rect 670 725 676 726
rect 734 730 740 731
rect 734 726 735 730
rect 739 726 740 730
rect 734 725 740 726
rect 798 730 804 731
rect 798 726 799 730
rect 803 726 804 730
rect 798 725 804 726
rect 862 730 868 731
rect 862 726 863 730
rect 867 726 868 730
rect 862 725 868 726
rect 926 730 932 731
rect 926 726 927 730
rect 931 726 932 730
rect 926 725 932 726
rect 990 730 996 731
rect 990 726 991 730
rect 995 726 996 730
rect 990 725 996 726
rect 1054 730 1060 731
rect 1054 726 1055 730
rect 1059 726 1060 730
rect 1054 725 1060 726
rect 1118 730 1124 731
rect 1118 726 1119 730
rect 1123 726 1124 730
rect 1118 725 1124 726
rect 1182 730 1188 731
rect 1182 726 1183 730
rect 1187 726 1188 730
rect 1182 725 1188 726
rect 1238 730 1244 731
rect 1238 726 1239 730
rect 1243 726 1244 730
rect 1238 725 1244 726
rect 1294 730 1300 731
rect 1294 726 1295 730
rect 1299 726 1300 730
rect 1294 725 1300 726
rect 1350 730 1356 731
rect 1350 726 1351 730
rect 1355 726 1356 730
rect 1350 725 1356 726
rect 1406 730 1412 731
rect 1406 726 1407 730
rect 1411 726 1412 730
rect 1406 725 1412 726
rect 1462 730 1468 731
rect 1462 726 1463 730
rect 1467 726 1468 730
rect 1462 725 1468 726
rect 1518 730 1524 731
rect 1518 726 1519 730
rect 1523 726 1524 730
rect 1518 725 1524 726
rect 1582 730 1588 731
rect 1582 726 1583 730
rect 1587 726 1588 730
rect 1582 725 1588 726
rect 1622 730 1628 731
rect 1622 726 1623 730
rect 1627 726 1628 730
rect 1622 725 1628 726
rect 1662 728 1668 729
rect 110 723 116 724
rect 112 711 114 723
rect 216 711 218 725
rect 248 711 250 725
rect 280 711 282 725
rect 320 711 322 725
rect 360 711 362 725
rect 400 711 402 725
rect 440 711 442 725
rect 488 711 490 725
rect 544 711 546 725
rect 608 711 610 725
rect 672 711 674 725
rect 736 711 738 725
rect 800 711 802 725
rect 864 711 866 725
rect 928 711 930 725
rect 992 711 994 725
rect 1056 711 1058 725
rect 1120 711 1122 725
rect 1184 711 1186 725
rect 1240 711 1242 725
rect 1296 711 1298 725
rect 1352 711 1354 725
rect 1408 711 1410 725
rect 1464 711 1466 725
rect 1520 711 1522 725
rect 1584 711 1586 725
rect 1624 711 1626 725
rect 1662 724 1663 728
rect 1667 724 1668 728
rect 1662 723 1668 724
rect 1664 711 1666 723
rect 111 710 115 711
rect 111 705 115 706
rect 215 710 219 711
rect 215 705 219 706
rect 247 710 251 711
rect 247 705 251 706
rect 279 710 283 711
rect 279 705 283 706
rect 311 710 315 711
rect 311 705 315 706
rect 319 710 323 711
rect 319 705 323 706
rect 343 710 347 711
rect 343 705 347 706
rect 359 710 363 711
rect 359 705 363 706
rect 375 710 379 711
rect 375 705 379 706
rect 399 710 403 711
rect 399 705 403 706
rect 407 710 411 711
rect 407 705 411 706
rect 439 710 443 711
rect 439 705 443 706
rect 471 710 475 711
rect 471 705 475 706
rect 487 710 491 711
rect 487 705 491 706
rect 503 710 507 711
rect 503 705 507 706
rect 543 710 547 711
rect 543 705 547 706
rect 591 710 595 711
rect 591 705 595 706
rect 607 710 611 711
rect 607 705 611 706
rect 647 710 651 711
rect 647 705 651 706
rect 671 710 675 711
rect 671 705 675 706
rect 703 710 707 711
rect 703 705 707 706
rect 735 710 739 711
rect 735 705 739 706
rect 759 710 763 711
rect 759 705 763 706
rect 799 710 803 711
rect 799 705 803 706
rect 823 710 827 711
rect 823 705 827 706
rect 863 710 867 711
rect 863 705 867 706
rect 887 710 891 711
rect 887 705 891 706
rect 927 710 931 711
rect 927 705 931 706
rect 959 710 963 711
rect 959 705 963 706
rect 991 710 995 711
rect 991 705 995 706
rect 1023 710 1027 711
rect 1023 705 1027 706
rect 1055 710 1059 711
rect 1055 705 1059 706
rect 1087 710 1091 711
rect 1087 705 1091 706
rect 1119 710 1123 711
rect 1119 705 1123 706
rect 1159 710 1163 711
rect 1159 705 1163 706
rect 1183 710 1187 711
rect 1183 705 1187 706
rect 1223 710 1227 711
rect 1223 705 1227 706
rect 1239 710 1243 711
rect 1239 705 1243 706
rect 1287 710 1291 711
rect 1287 705 1291 706
rect 1295 710 1299 711
rect 1295 705 1299 706
rect 1351 710 1355 711
rect 1351 705 1355 706
rect 1407 710 1411 711
rect 1407 705 1411 706
rect 1415 710 1419 711
rect 1415 705 1419 706
rect 1463 710 1467 711
rect 1463 705 1467 706
rect 1471 710 1475 711
rect 1471 705 1475 706
rect 1519 710 1523 711
rect 1519 705 1523 706
rect 1527 710 1531 711
rect 1527 705 1531 706
rect 1583 710 1587 711
rect 1583 705 1587 706
rect 1623 710 1627 711
rect 1623 705 1627 706
rect 1663 710 1667 711
rect 1663 705 1667 706
rect 112 697 114 705
rect 110 696 116 697
rect 110 692 111 696
rect 115 692 116 696
rect 280 695 282 705
rect 312 695 314 705
rect 344 695 346 705
rect 376 695 378 705
rect 408 695 410 705
rect 440 695 442 705
rect 472 695 474 705
rect 504 695 506 705
rect 544 695 546 705
rect 592 695 594 705
rect 648 695 650 705
rect 704 695 706 705
rect 760 695 762 705
rect 824 695 826 705
rect 888 695 890 705
rect 960 695 962 705
rect 1024 695 1026 705
rect 1088 695 1090 705
rect 1160 695 1162 705
rect 1224 695 1226 705
rect 1288 695 1290 705
rect 1352 695 1354 705
rect 1416 695 1418 705
rect 1472 695 1474 705
rect 1528 695 1530 705
rect 1584 695 1586 705
rect 1624 695 1626 705
rect 1664 697 1666 705
rect 1662 696 1668 697
rect 110 691 116 692
rect 278 694 284 695
rect 278 690 279 694
rect 283 690 284 694
rect 278 689 284 690
rect 310 694 316 695
rect 310 690 311 694
rect 315 690 316 694
rect 310 689 316 690
rect 342 694 348 695
rect 342 690 343 694
rect 347 690 348 694
rect 342 689 348 690
rect 374 694 380 695
rect 374 690 375 694
rect 379 690 380 694
rect 374 689 380 690
rect 406 694 412 695
rect 406 690 407 694
rect 411 690 412 694
rect 406 689 412 690
rect 438 694 444 695
rect 438 690 439 694
rect 443 690 444 694
rect 438 689 444 690
rect 470 694 476 695
rect 470 690 471 694
rect 475 690 476 694
rect 470 689 476 690
rect 502 694 508 695
rect 502 690 503 694
rect 507 690 508 694
rect 502 689 508 690
rect 542 694 548 695
rect 542 690 543 694
rect 547 690 548 694
rect 542 689 548 690
rect 590 694 596 695
rect 590 690 591 694
rect 595 690 596 694
rect 590 689 596 690
rect 646 694 652 695
rect 646 690 647 694
rect 651 690 652 694
rect 646 689 652 690
rect 702 694 708 695
rect 702 690 703 694
rect 707 690 708 694
rect 702 689 708 690
rect 758 694 764 695
rect 758 690 759 694
rect 763 690 764 694
rect 758 689 764 690
rect 822 694 828 695
rect 822 690 823 694
rect 827 690 828 694
rect 822 689 828 690
rect 886 694 892 695
rect 886 690 887 694
rect 891 690 892 694
rect 886 689 892 690
rect 958 694 964 695
rect 958 690 959 694
rect 963 690 964 694
rect 958 689 964 690
rect 1022 694 1028 695
rect 1022 690 1023 694
rect 1027 690 1028 694
rect 1022 689 1028 690
rect 1086 694 1092 695
rect 1086 690 1087 694
rect 1091 690 1092 694
rect 1086 689 1092 690
rect 1158 694 1164 695
rect 1158 690 1159 694
rect 1163 690 1164 694
rect 1158 689 1164 690
rect 1222 694 1228 695
rect 1222 690 1223 694
rect 1227 690 1228 694
rect 1222 689 1228 690
rect 1286 694 1292 695
rect 1286 690 1287 694
rect 1291 690 1292 694
rect 1286 689 1292 690
rect 1350 694 1356 695
rect 1350 690 1351 694
rect 1355 690 1356 694
rect 1350 689 1356 690
rect 1414 694 1420 695
rect 1414 690 1415 694
rect 1419 690 1420 694
rect 1414 689 1420 690
rect 1470 694 1476 695
rect 1470 690 1471 694
rect 1475 690 1476 694
rect 1470 689 1476 690
rect 1526 694 1532 695
rect 1526 690 1527 694
rect 1531 690 1532 694
rect 1526 689 1532 690
rect 1582 694 1588 695
rect 1582 690 1583 694
rect 1587 690 1588 694
rect 1582 689 1588 690
rect 1622 694 1628 695
rect 1622 690 1623 694
rect 1627 690 1628 694
rect 1662 692 1663 696
rect 1667 692 1668 696
rect 1662 691 1668 692
rect 1622 689 1628 690
rect 110 679 116 680
rect 110 675 111 679
rect 115 675 116 679
rect 1662 679 1668 680
rect 110 674 116 675
rect 278 677 284 678
rect 112 671 114 674
rect 278 673 279 677
rect 283 673 284 677
rect 278 672 284 673
rect 310 677 316 678
rect 310 673 311 677
rect 315 673 316 677
rect 310 672 316 673
rect 342 677 348 678
rect 342 673 343 677
rect 347 673 348 677
rect 342 672 348 673
rect 374 677 380 678
rect 374 673 375 677
rect 379 673 380 677
rect 374 672 380 673
rect 406 677 412 678
rect 406 673 407 677
rect 411 673 412 677
rect 406 672 412 673
rect 438 677 444 678
rect 438 673 439 677
rect 443 673 444 677
rect 438 672 444 673
rect 470 677 476 678
rect 470 673 471 677
rect 475 673 476 677
rect 470 672 476 673
rect 502 677 508 678
rect 502 673 503 677
rect 507 673 508 677
rect 502 672 508 673
rect 542 677 548 678
rect 542 673 543 677
rect 547 673 548 677
rect 542 672 548 673
rect 590 677 596 678
rect 590 673 591 677
rect 595 673 596 677
rect 590 672 596 673
rect 646 677 652 678
rect 646 673 647 677
rect 651 673 652 677
rect 646 672 652 673
rect 702 677 708 678
rect 702 673 703 677
rect 707 673 708 677
rect 702 672 708 673
rect 758 677 764 678
rect 758 673 759 677
rect 763 673 764 677
rect 758 672 764 673
rect 822 677 828 678
rect 822 673 823 677
rect 827 673 828 677
rect 822 672 828 673
rect 886 677 892 678
rect 886 673 887 677
rect 891 673 892 677
rect 886 672 892 673
rect 958 677 964 678
rect 958 673 959 677
rect 963 673 964 677
rect 958 672 964 673
rect 1022 677 1028 678
rect 1022 673 1023 677
rect 1027 673 1028 677
rect 1022 672 1028 673
rect 1086 677 1092 678
rect 1086 673 1087 677
rect 1091 673 1092 677
rect 1086 672 1092 673
rect 1158 677 1164 678
rect 1158 673 1159 677
rect 1163 673 1164 677
rect 1158 672 1164 673
rect 1222 677 1228 678
rect 1222 673 1223 677
rect 1227 673 1228 677
rect 1222 672 1228 673
rect 1286 677 1292 678
rect 1286 673 1287 677
rect 1291 673 1292 677
rect 1286 672 1292 673
rect 1350 677 1356 678
rect 1350 673 1351 677
rect 1355 673 1356 677
rect 1350 672 1356 673
rect 1414 677 1420 678
rect 1414 673 1415 677
rect 1419 673 1420 677
rect 1414 672 1420 673
rect 1470 677 1476 678
rect 1470 673 1471 677
rect 1475 673 1476 677
rect 1470 672 1476 673
rect 1526 677 1532 678
rect 1526 673 1527 677
rect 1531 673 1532 677
rect 1526 672 1532 673
rect 1582 677 1588 678
rect 1582 673 1583 677
rect 1587 673 1588 677
rect 1582 672 1588 673
rect 1622 677 1628 678
rect 1622 673 1623 677
rect 1627 673 1628 677
rect 1662 675 1663 679
rect 1667 675 1668 679
rect 1662 674 1668 675
rect 1622 672 1628 673
rect 111 670 115 671
rect 111 665 115 666
rect 279 670 283 672
rect 279 665 283 666
rect 295 670 299 671
rect 112 662 114 665
rect 295 664 299 666
rect 311 670 315 672
rect 311 665 315 666
rect 327 670 331 671
rect 327 664 331 666
rect 343 670 347 672
rect 343 665 347 666
rect 359 670 363 671
rect 359 664 363 666
rect 375 670 379 672
rect 375 665 379 666
rect 391 670 395 671
rect 391 664 395 666
rect 407 670 411 672
rect 407 665 411 666
rect 423 670 427 671
rect 423 664 427 666
rect 439 670 443 672
rect 439 665 443 666
rect 455 670 459 671
rect 455 664 459 666
rect 471 670 475 672
rect 471 665 475 666
rect 487 670 491 671
rect 487 664 491 666
rect 503 670 507 672
rect 503 665 507 666
rect 519 670 523 671
rect 519 664 523 666
rect 543 670 547 672
rect 543 665 547 666
rect 551 670 555 671
rect 551 664 555 666
rect 591 670 595 672
rect 591 664 595 666
rect 639 670 643 671
rect 639 664 643 666
rect 647 670 651 672
rect 647 665 651 666
rect 687 670 691 671
rect 687 664 691 666
rect 703 670 707 672
rect 703 665 707 666
rect 735 670 739 671
rect 735 664 739 666
rect 759 670 763 672
rect 759 665 763 666
rect 791 670 795 671
rect 791 664 795 666
rect 823 670 827 672
rect 823 665 827 666
rect 847 670 851 671
rect 847 664 851 666
rect 887 670 891 672
rect 887 665 891 666
rect 911 670 915 671
rect 911 664 915 666
rect 959 670 963 672
rect 959 665 963 666
rect 975 670 979 671
rect 975 664 979 666
rect 1023 670 1027 672
rect 1023 665 1027 666
rect 1047 670 1051 671
rect 1047 664 1051 666
rect 1087 670 1091 672
rect 1087 665 1091 666
rect 1127 670 1131 671
rect 1127 664 1131 666
rect 1159 670 1163 672
rect 1159 665 1163 666
rect 1215 670 1219 671
rect 1215 664 1219 666
rect 1223 670 1227 672
rect 1223 665 1227 666
rect 1287 670 1291 672
rect 1287 665 1291 666
rect 1295 670 1299 671
rect 1295 664 1299 666
rect 1351 670 1355 672
rect 1351 665 1355 666
rect 1383 670 1387 671
rect 1383 664 1387 666
rect 1415 670 1419 672
rect 1415 665 1419 666
rect 1471 670 1475 672
rect 1471 664 1475 666
rect 1527 670 1531 672
rect 1527 665 1531 666
rect 1559 670 1563 671
rect 1559 664 1563 666
rect 1583 670 1587 672
rect 1583 665 1587 666
rect 1623 670 1627 672
rect 1664 671 1666 674
rect 1623 664 1627 666
rect 1663 670 1667 671
rect 1663 665 1667 666
rect 294 663 300 664
rect 110 661 116 662
rect 110 657 111 661
rect 115 657 116 661
rect 294 659 295 663
rect 299 659 300 663
rect 294 658 300 659
rect 326 663 332 664
rect 326 659 327 663
rect 331 659 332 663
rect 326 658 332 659
rect 358 663 364 664
rect 358 659 359 663
rect 363 659 364 663
rect 358 658 364 659
rect 390 663 396 664
rect 390 659 391 663
rect 395 659 396 663
rect 390 658 396 659
rect 422 663 428 664
rect 422 659 423 663
rect 427 659 428 663
rect 422 658 428 659
rect 454 663 460 664
rect 454 659 455 663
rect 459 659 460 663
rect 454 658 460 659
rect 486 663 492 664
rect 486 659 487 663
rect 491 659 492 663
rect 486 658 492 659
rect 518 663 524 664
rect 518 659 519 663
rect 523 659 524 663
rect 518 658 524 659
rect 550 663 556 664
rect 550 659 551 663
rect 555 659 556 663
rect 550 658 556 659
rect 590 663 596 664
rect 590 659 591 663
rect 595 659 596 663
rect 590 658 596 659
rect 638 663 644 664
rect 638 659 639 663
rect 643 659 644 663
rect 638 658 644 659
rect 686 663 692 664
rect 686 659 687 663
rect 691 659 692 663
rect 686 658 692 659
rect 734 663 740 664
rect 734 659 735 663
rect 739 659 740 663
rect 734 658 740 659
rect 790 663 796 664
rect 790 659 791 663
rect 795 659 796 663
rect 790 658 796 659
rect 846 663 852 664
rect 846 659 847 663
rect 851 659 852 663
rect 846 658 852 659
rect 910 663 916 664
rect 910 659 911 663
rect 915 659 916 663
rect 910 658 916 659
rect 974 663 980 664
rect 974 659 975 663
rect 979 659 980 663
rect 974 658 980 659
rect 1046 663 1052 664
rect 1046 659 1047 663
rect 1051 659 1052 663
rect 1046 658 1052 659
rect 1126 663 1132 664
rect 1126 659 1127 663
rect 1131 659 1132 663
rect 1126 658 1132 659
rect 1214 663 1220 664
rect 1214 659 1215 663
rect 1219 659 1220 663
rect 1214 658 1220 659
rect 1294 663 1300 664
rect 1294 659 1295 663
rect 1299 659 1300 663
rect 1294 658 1300 659
rect 1382 663 1388 664
rect 1382 659 1383 663
rect 1387 659 1388 663
rect 1382 658 1388 659
rect 1470 663 1476 664
rect 1470 659 1471 663
rect 1475 659 1476 663
rect 1470 658 1476 659
rect 1558 663 1564 664
rect 1558 659 1559 663
rect 1563 659 1564 663
rect 1558 658 1564 659
rect 1622 663 1628 664
rect 1622 659 1623 663
rect 1627 659 1628 663
rect 1664 662 1666 665
rect 1622 658 1628 659
rect 1662 661 1668 662
rect 110 656 116 657
rect 1662 657 1663 661
rect 1667 657 1668 661
rect 1662 656 1668 657
rect 294 646 300 647
rect 110 644 116 645
rect 110 640 111 644
rect 115 640 116 644
rect 294 642 295 646
rect 299 642 300 646
rect 294 641 300 642
rect 326 646 332 647
rect 326 642 327 646
rect 331 642 332 646
rect 326 641 332 642
rect 358 646 364 647
rect 358 642 359 646
rect 363 642 364 646
rect 358 641 364 642
rect 390 646 396 647
rect 390 642 391 646
rect 395 642 396 646
rect 390 641 396 642
rect 422 646 428 647
rect 422 642 423 646
rect 427 642 428 646
rect 422 641 428 642
rect 454 646 460 647
rect 454 642 455 646
rect 459 642 460 646
rect 454 641 460 642
rect 486 646 492 647
rect 486 642 487 646
rect 491 642 492 646
rect 486 641 492 642
rect 518 646 524 647
rect 518 642 519 646
rect 523 642 524 646
rect 518 641 524 642
rect 550 646 556 647
rect 550 642 551 646
rect 555 642 556 646
rect 550 641 556 642
rect 590 646 596 647
rect 590 642 591 646
rect 595 642 596 646
rect 590 641 596 642
rect 638 646 644 647
rect 638 642 639 646
rect 643 642 644 646
rect 638 641 644 642
rect 686 646 692 647
rect 686 642 687 646
rect 691 642 692 646
rect 686 641 692 642
rect 734 646 740 647
rect 734 642 735 646
rect 739 642 740 646
rect 734 641 740 642
rect 790 646 796 647
rect 790 642 791 646
rect 795 642 796 646
rect 790 641 796 642
rect 846 646 852 647
rect 846 642 847 646
rect 851 642 852 646
rect 846 641 852 642
rect 910 646 916 647
rect 910 642 911 646
rect 915 642 916 646
rect 910 641 916 642
rect 974 646 980 647
rect 974 642 975 646
rect 979 642 980 646
rect 974 641 980 642
rect 1046 646 1052 647
rect 1046 642 1047 646
rect 1051 642 1052 646
rect 1046 641 1052 642
rect 1126 646 1132 647
rect 1126 642 1127 646
rect 1131 642 1132 646
rect 1126 641 1132 642
rect 1214 646 1220 647
rect 1214 642 1215 646
rect 1219 642 1220 646
rect 1214 641 1220 642
rect 1294 646 1300 647
rect 1294 642 1295 646
rect 1299 642 1300 646
rect 1294 641 1300 642
rect 1382 646 1388 647
rect 1382 642 1383 646
rect 1387 642 1388 646
rect 1382 641 1388 642
rect 1470 646 1476 647
rect 1470 642 1471 646
rect 1475 642 1476 646
rect 1470 641 1476 642
rect 1558 646 1564 647
rect 1558 642 1559 646
rect 1563 642 1564 646
rect 1558 641 1564 642
rect 1622 646 1628 647
rect 1622 642 1623 646
rect 1627 642 1628 646
rect 1622 641 1628 642
rect 1662 644 1668 645
rect 110 639 116 640
rect 112 631 114 639
rect 296 631 298 641
rect 328 631 330 641
rect 360 631 362 641
rect 392 631 394 641
rect 424 631 426 641
rect 456 631 458 641
rect 488 631 490 641
rect 520 631 522 641
rect 552 631 554 641
rect 592 631 594 641
rect 640 631 642 641
rect 688 631 690 641
rect 736 631 738 641
rect 792 631 794 641
rect 848 631 850 641
rect 912 631 914 641
rect 976 631 978 641
rect 1048 631 1050 641
rect 1128 631 1130 641
rect 1216 631 1218 641
rect 1296 631 1298 641
rect 1384 631 1386 641
rect 1472 631 1474 641
rect 1560 631 1562 641
rect 1624 631 1626 641
rect 1662 640 1663 644
rect 1667 640 1668 644
rect 1662 639 1668 640
rect 1664 631 1666 639
rect 111 630 115 631
rect 111 625 115 626
rect 247 630 251 631
rect 247 625 251 626
rect 279 630 283 631
rect 279 625 283 626
rect 295 630 299 631
rect 295 625 299 626
rect 319 630 323 631
rect 319 625 323 626
rect 327 630 331 631
rect 327 625 331 626
rect 359 630 363 631
rect 359 625 363 626
rect 367 630 371 631
rect 367 625 371 626
rect 391 630 395 631
rect 391 625 395 626
rect 423 630 427 631
rect 423 625 427 626
rect 455 630 459 631
rect 455 625 459 626
rect 471 630 475 631
rect 471 625 475 626
rect 487 630 491 631
rect 487 625 491 626
rect 519 630 523 631
rect 519 625 523 626
rect 551 630 555 631
rect 551 625 555 626
rect 567 630 571 631
rect 567 625 571 626
rect 591 630 595 631
rect 591 625 595 626
rect 615 630 619 631
rect 615 625 619 626
rect 639 630 643 631
rect 639 625 643 626
rect 663 630 667 631
rect 663 625 667 626
rect 687 630 691 631
rect 687 625 691 626
rect 719 630 723 631
rect 719 625 723 626
rect 735 630 739 631
rect 735 625 739 626
rect 775 630 779 631
rect 775 625 779 626
rect 791 630 795 631
rect 791 625 795 626
rect 831 630 835 631
rect 831 625 835 626
rect 847 630 851 631
rect 847 625 851 626
rect 895 630 899 631
rect 895 625 899 626
rect 911 630 915 631
rect 911 625 915 626
rect 967 630 971 631
rect 967 625 971 626
rect 975 630 979 631
rect 975 625 979 626
rect 1047 630 1051 631
rect 1047 625 1051 626
rect 1127 630 1131 631
rect 1127 625 1131 626
rect 1207 630 1211 631
rect 1207 625 1211 626
rect 1215 630 1219 631
rect 1215 625 1219 626
rect 1287 630 1291 631
rect 1287 625 1291 626
rect 1295 630 1299 631
rect 1295 625 1299 626
rect 1359 630 1363 631
rect 1359 625 1363 626
rect 1383 630 1387 631
rect 1383 625 1387 626
rect 1431 630 1435 631
rect 1431 625 1435 626
rect 1471 630 1475 631
rect 1471 625 1475 626
rect 1503 630 1507 631
rect 1503 625 1507 626
rect 1559 630 1563 631
rect 1559 625 1563 626
rect 1575 630 1579 631
rect 1575 625 1579 626
rect 1623 630 1627 631
rect 1623 625 1627 626
rect 1663 630 1667 631
rect 1663 625 1667 626
rect 112 617 114 625
rect 110 616 116 617
rect 110 612 111 616
rect 115 612 116 616
rect 248 615 250 625
rect 280 615 282 625
rect 320 615 322 625
rect 368 615 370 625
rect 424 615 426 625
rect 472 615 474 625
rect 520 615 522 625
rect 568 615 570 625
rect 616 615 618 625
rect 664 615 666 625
rect 720 615 722 625
rect 776 615 778 625
rect 832 615 834 625
rect 896 615 898 625
rect 968 615 970 625
rect 1048 615 1050 625
rect 1128 615 1130 625
rect 1208 615 1210 625
rect 1288 615 1290 625
rect 1360 615 1362 625
rect 1432 615 1434 625
rect 1504 615 1506 625
rect 1576 615 1578 625
rect 1624 615 1626 625
rect 1664 617 1666 625
rect 1662 616 1668 617
rect 110 611 116 612
rect 246 614 252 615
rect 246 610 247 614
rect 251 610 252 614
rect 246 609 252 610
rect 278 614 284 615
rect 278 610 279 614
rect 283 610 284 614
rect 278 609 284 610
rect 318 614 324 615
rect 318 610 319 614
rect 323 610 324 614
rect 318 609 324 610
rect 366 614 372 615
rect 366 610 367 614
rect 371 610 372 614
rect 366 609 372 610
rect 422 614 428 615
rect 422 610 423 614
rect 427 610 428 614
rect 422 609 428 610
rect 470 614 476 615
rect 470 610 471 614
rect 475 610 476 614
rect 470 609 476 610
rect 518 614 524 615
rect 518 610 519 614
rect 523 610 524 614
rect 518 609 524 610
rect 566 614 572 615
rect 566 610 567 614
rect 571 610 572 614
rect 566 609 572 610
rect 614 614 620 615
rect 614 610 615 614
rect 619 610 620 614
rect 614 609 620 610
rect 662 614 668 615
rect 662 610 663 614
rect 667 610 668 614
rect 662 609 668 610
rect 718 614 724 615
rect 718 610 719 614
rect 723 610 724 614
rect 718 609 724 610
rect 774 614 780 615
rect 774 610 775 614
rect 779 610 780 614
rect 774 609 780 610
rect 830 614 836 615
rect 830 610 831 614
rect 835 610 836 614
rect 830 609 836 610
rect 894 614 900 615
rect 894 610 895 614
rect 899 610 900 614
rect 894 609 900 610
rect 966 614 972 615
rect 966 610 967 614
rect 971 610 972 614
rect 966 609 972 610
rect 1046 614 1052 615
rect 1046 610 1047 614
rect 1051 610 1052 614
rect 1046 609 1052 610
rect 1126 614 1132 615
rect 1126 610 1127 614
rect 1131 610 1132 614
rect 1126 609 1132 610
rect 1206 614 1212 615
rect 1206 610 1207 614
rect 1211 610 1212 614
rect 1206 609 1212 610
rect 1286 614 1292 615
rect 1286 610 1287 614
rect 1291 610 1292 614
rect 1286 609 1292 610
rect 1358 614 1364 615
rect 1358 610 1359 614
rect 1363 610 1364 614
rect 1358 609 1364 610
rect 1430 614 1436 615
rect 1430 610 1431 614
rect 1435 610 1436 614
rect 1430 609 1436 610
rect 1502 614 1508 615
rect 1502 610 1503 614
rect 1507 610 1508 614
rect 1502 609 1508 610
rect 1574 614 1580 615
rect 1574 610 1575 614
rect 1579 610 1580 614
rect 1574 609 1580 610
rect 1622 614 1628 615
rect 1622 610 1623 614
rect 1627 610 1628 614
rect 1662 612 1663 616
rect 1667 612 1668 616
rect 1662 611 1668 612
rect 1622 609 1628 610
rect 110 599 116 600
rect 110 595 111 599
rect 115 595 116 599
rect 1662 599 1668 600
rect 110 594 116 595
rect 246 597 252 598
rect 112 591 114 594
rect 246 593 247 597
rect 251 593 252 597
rect 246 592 252 593
rect 278 597 284 598
rect 278 593 279 597
rect 283 593 284 597
rect 278 592 284 593
rect 318 597 324 598
rect 318 593 319 597
rect 323 593 324 597
rect 318 592 324 593
rect 366 597 372 598
rect 366 593 367 597
rect 371 593 372 597
rect 366 592 372 593
rect 422 597 428 598
rect 422 593 423 597
rect 427 593 428 597
rect 422 592 428 593
rect 470 597 476 598
rect 470 593 471 597
rect 475 593 476 597
rect 470 592 476 593
rect 518 597 524 598
rect 518 593 519 597
rect 523 593 524 597
rect 518 592 524 593
rect 566 597 572 598
rect 566 593 567 597
rect 571 593 572 597
rect 566 592 572 593
rect 614 597 620 598
rect 614 593 615 597
rect 619 593 620 597
rect 614 592 620 593
rect 662 597 668 598
rect 662 593 663 597
rect 667 593 668 597
rect 662 592 668 593
rect 718 597 724 598
rect 718 593 719 597
rect 723 593 724 597
rect 718 592 724 593
rect 774 597 780 598
rect 774 593 775 597
rect 779 593 780 597
rect 774 592 780 593
rect 830 597 836 598
rect 830 593 831 597
rect 835 593 836 597
rect 830 592 836 593
rect 894 597 900 598
rect 894 593 895 597
rect 899 593 900 597
rect 894 592 900 593
rect 966 597 972 598
rect 966 593 967 597
rect 971 593 972 597
rect 966 592 972 593
rect 1046 597 1052 598
rect 1046 593 1047 597
rect 1051 593 1052 597
rect 1046 592 1052 593
rect 1126 597 1132 598
rect 1126 593 1127 597
rect 1131 593 1132 597
rect 1126 592 1132 593
rect 1206 597 1212 598
rect 1206 593 1207 597
rect 1211 593 1212 597
rect 1206 592 1212 593
rect 1286 597 1292 598
rect 1286 593 1287 597
rect 1291 593 1292 597
rect 1286 592 1292 593
rect 1358 597 1364 598
rect 1358 593 1359 597
rect 1363 593 1364 597
rect 1358 592 1364 593
rect 1430 597 1436 598
rect 1430 593 1431 597
rect 1435 593 1436 597
rect 1430 592 1436 593
rect 1502 597 1508 598
rect 1502 593 1503 597
rect 1507 593 1508 597
rect 1502 592 1508 593
rect 1574 597 1580 598
rect 1574 593 1575 597
rect 1579 593 1580 597
rect 1574 592 1580 593
rect 1622 597 1628 598
rect 1622 593 1623 597
rect 1627 593 1628 597
rect 1662 595 1663 599
rect 1667 595 1668 599
rect 1662 594 1668 595
rect 1622 592 1628 593
rect 111 590 115 591
rect 111 585 115 586
rect 167 590 171 591
rect 112 582 114 585
rect 167 584 171 586
rect 215 590 219 591
rect 215 584 219 586
rect 247 590 251 592
rect 247 585 251 586
rect 271 590 275 591
rect 271 584 275 586
rect 279 590 283 592
rect 279 585 283 586
rect 319 590 323 592
rect 319 585 323 586
rect 335 590 339 591
rect 335 584 339 586
rect 367 590 371 592
rect 367 585 371 586
rect 407 590 411 591
rect 407 584 411 586
rect 423 590 427 592
rect 423 585 427 586
rect 471 590 475 592
rect 471 585 475 586
rect 487 590 491 591
rect 487 584 491 586
rect 519 590 523 592
rect 519 585 523 586
rect 559 590 563 591
rect 559 584 563 586
rect 567 590 571 592
rect 567 585 571 586
rect 615 590 619 592
rect 615 585 619 586
rect 631 590 635 591
rect 631 584 635 586
rect 663 590 667 592
rect 663 585 667 586
rect 703 590 707 591
rect 703 584 707 586
rect 719 590 723 592
rect 719 585 723 586
rect 767 590 771 591
rect 767 584 771 586
rect 775 590 779 592
rect 775 585 779 586
rect 823 590 827 591
rect 823 584 827 586
rect 831 590 835 592
rect 831 585 835 586
rect 879 590 883 591
rect 879 584 883 586
rect 895 590 899 592
rect 895 585 899 586
rect 935 590 939 591
rect 935 584 939 586
rect 967 590 971 592
rect 967 585 971 586
rect 991 590 995 591
rect 991 584 995 586
rect 1047 590 1051 592
rect 1047 584 1051 586
rect 1103 590 1107 591
rect 1103 584 1107 586
rect 1127 590 1131 592
rect 1127 585 1131 586
rect 1159 590 1163 591
rect 1159 584 1163 586
rect 1207 590 1211 592
rect 1207 585 1211 586
rect 1215 590 1219 591
rect 1215 584 1219 586
rect 1271 590 1275 591
rect 1271 584 1275 586
rect 1287 590 1291 592
rect 1287 585 1291 586
rect 1327 590 1331 591
rect 1327 584 1331 586
rect 1359 590 1363 592
rect 1359 585 1363 586
rect 1383 590 1387 591
rect 1383 584 1387 586
rect 1431 590 1435 592
rect 1431 585 1435 586
rect 1447 590 1451 591
rect 1447 584 1451 586
rect 1503 590 1507 592
rect 1503 585 1507 586
rect 1511 590 1515 591
rect 1511 584 1515 586
rect 1575 590 1579 592
rect 1575 584 1579 586
rect 1623 590 1627 592
rect 1664 591 1666 594
rect 1623 584 1627 586
rect 1663 590 1667 591
rect 1663 585 1667 586
rect 166 583 172 584
rect 110 581 116 582
rect 110 577 111 581
rect 115 577 116 581
rect 166 579 167 583
rect 171 579 172 583
rect 166 578 172 579
rect 214 583 220 584
rect 214 579 215 583
rect 219 579 220 583
rect 214 578 220 579
rect 270 583 276 584
rect 270 579 271 583
rect 275 579 276 583
rect 270 578 276 579
rect 334 583 340 584
rect 334 579 335 583
rect 339 579 340 583
rect 334 578 340 579
rect 406 583 412 584
rect 406 579 407 583
rect 411 579 412 583
rect 406 578 412 579
rect 486 583 492 584
rect 486 579 487 583
rect 491 579 492 583
rect 486 578 492 579
rect 558 583 564 584
rect 558 579 559 583
rect 563 579 564 583
rect 558 578 564 579
rect 630 583 636 584
rect 630 579 631 583
rect 635 579 636 583
rect 630 578 636 579
rect 702 583 708 584
rect 702 579 703 583
rect 707 579 708 583
rect 702 578 708 579
rect 766 583 772 584
rect 766 579 767 583
rect 771 579 772 583
rect 766 578 772 579
rect 822 583 828 584
rect 822 579 823 583
rect 827 579 828 583
rect 822 578 828 579
rect 878 583 884 584
rect 878 579 879 583
rect 883 579 884 583
rect 878 578 884 579
rect 934 583 940 584
rect 934 579 935 583
rect 939 579 940 583
rect 934 578 940 579
rect 990 583 996 584
rect 990 579 991 583
rect 995 579 996 583
rect 990 578 996 579
rect 1046 583 1052 584
rect 1046 579 1047 583
rect 1051 579 1052 583
rect 1046 578 1052 579
rect 1102 583 1108 584
rect 1102 579 1103 583
rect 1107 579 1108 583
rect 1102 578 1108 579
rect 1158 583 1164 584
rect 1158 579 1159 583
rect 1163 579 1164 583
rect 1158 578 1164 579
rect 1214 583 1220 584
rect 1214 579 1215 583
rect 1219 579 1220 583
rect 1214 578 1220 579
rect 1270 583 1276 584
rect 1270 579 1271 583
rect 1275 579 1276 583
rect 1270 578 1276 579
rect 1326 583 1332 584
rect 1326 579 1327 583
rect 1331 579 1332 583
rect 1326 578 1332 579
rect 1382 583 1388 584
rect 1382 579 1383 583
rect 1387 579 1388 583
rect 1382 578 1388 579
rect 1446 583 1452 584
rect 1446 579 1447 583
rect 1451 579 1452 583
rect 1446 578 1452 579
rect 1510 583 1516 584
rect 1510 579 1511 583
rect 1515 579 1516 583
rect 1510 578 1516 579
rect 1574 583 1580 584
rect 1574 579 1575 583
rect 1579 579 1580 583
rect 1574 578 1580 579
rect 1622 583 1628 584
rect 1622 579 1623 583
rect 1627 579 1628 583
rect 1664 582 1666 585
rect 1622 578 1628 579
rect 1662 581 1668 582
rect 110 576 116 577
rect 1662 577 1663 581
rect 1667 577 1668 581
rect 1662 576 1668 577
rect 166 566 172 567
rect 110 564 116 565
rect 110 560 111 564
rect 115 560 116 564
rect 166 562 167 566
rect 171 562 172 566
rect 166 561 172 562
rect 214 566 220 567
rect 214 562 215 566
rect 219 562 220 566
rect 214 561 220 562
rect 270 566 276 567
rect 270 562 271 566
rect 275 562 276 566
rect 270 561 276 562
rect 334 566 340 567
rect 334 562 335 566
rect 339 562 340 566
rect 334 561 340 562
rect 406 566 412 567
rect 406 562 407 566
rect 411 562 412 566
rect 406 561 412 562
rect 486 566 492 567
rect 486 562 487 566
rect 491 562 492 566
rect 486 561 492 562
rect 558 566 564 567
rect 558 562 559 566
rect 563 562 564 566
rect 558 561 564 562
rect 630 566 636 567
rect 630 562 631 566
rect 635 562 636 566
rect 630 561 636 562
rect 702 566 708 567
rect 702 562 703 566
rect 707 562 708 566
rect 702 561 708 562
rect 766 566 772 567
rect 766 562 767 566
rect 771 562 772 566
rect 766 561 772 562
rect 822 566 828 567
rect 822 562 823 566
rect 827 562 828 566
rect 822 561 828 562
rect 878 566 884 567
rect 878 562 879 566
rect 883 562 884 566
rect 878 561 884 562
rect 934 566 940 567
rect 934 562 935 566
rect 939 562 940 566
rect 934 561 940 562
rect 990 566 996 567
rect 990 562 991 566
rect 995 562 996 566
rect 990 561 996 562
rect 1046 566 1052 567
rect 1046 562 1047 566
rect 1051 562 1052 566
rect 1046 561 1052 562
rect 1102 566 1108 567
rect 1102 562 1103 566
rect 1107 562 1108 566
rect 1102 561 1108 562
rect 1158 566 1164 567
rect 1158 562 1159 566
rect 1163 562 1164 566
rect 1158 561 1164 562
rect 1214 566 1220 567
rect 1214 562 1215 566
rect 1219 562 1220 566
rect 1214 561 1220 562
rect 1270 566 1276 567
rect 1270 562 1271 566
rect 1275 562 1276 566
rect 1270 561 1276 562
rect 1326 566 1332 567
rect 1326 562 1327 566
rect 1331 562 1332 566
rect 1326 561 1332 562
rect 1382 566 1388 567
rect 1382 562 1383 566
rect 1387 562 1388 566
rect 1382 561 1388 562
rect 1446 566 1452 567
rect 1446 562 1447 566
rect 1451 562 1452 566
rect 1446 561 1452 562
rect 1510 566 1516 567
rect 1510 562 1511 566
rect 1515 562 1516 566
rect 1510 561 1516 562
rect 1574 566 1580 567
rect 1574 562 1575 566
rect 1579 562 1580 566
rect 1574 561 1580 562
rect 1622 566 1628 567
rect 1622 562 1623 566
rect 1627 562 1628 566
rect 1622 561 1628 562
rect 1662 564 1668 565
rect 110 559 116 560
rect 112 547 114 559
rect 168 547 170 561
rect 216 547 218 561
rect 272 547 274 561
rect 336 547 338 561
rect 408 547 410 561
rect 488 547 490 561
rect 560 547 562 561
rect 632 547 634 561
rect 704 547 706 561
rect 768 547 770 561
rect 824 547 826 561
rect 880 547 882 561
rect 936 547 938 561
rect 992 547 994 561
rect 1048 547 1050 561
rect 1104 547 1106 561
rect 1160 547 1162 561
rect 1216 547 1218 561
rect 1272 547 1274 561
rect 1328 547 1330 561
rect 1384 547 1386 561
rect 1448 547 1450 561
rect 1512 547 1514 561
rect 1576 547 1578 561
rect 1624 547 1626 561
rect 1662 560 1663 564
rect 1667 560 1668 564
rect 1662 559 1668 560
rect 1664 547 1666 559
rect 111 546 115 547
rect 111 541 115 542
rect 135 546 139 547
rect 135 541 139 542
rect 167 546 171 547
rect 167 541 171 542
rect 199 546 203 547
rect 199 541 203 542
rect 215 546 219 547
rect 215 541 219 542
rect 231 546 235 547
rect 231 541 235 542
rect 271 546 275 547
rect 271 541 275 542
rect 279 546 283 547
rect 279 541 283 542
rect 327 546 331 547
rect 327 541 331 542
rect 335 546 339 547
rect 335 541 339 542
rect 375 546 379 547
rect 375 541 379 542
rect 407 546 411 547
rect 407 541 411 542
rect 431 546 435 547
rect 431 541 435 542
rect 487 546 491 547
rect 487 541 491 542
rect 495 546 499 547
rect 495 541 499 542
rect 559 546 563 547
rect 559 541 563 542
rect 623 546 627 547
rect 623 541 627 542
rect 631 546 635 547
rect 631 541 635 542
rect 687 546 691 547
rect 687 541 691 542
rect 703 546 707 547
rect 703 541 707 542
rect 751 546 755 547
rect 751 541 755 542
rect 767 546 771 547
rect 767 541 771 542
rect 815 546 819 547
rect 815 541 819 542
rect 823 546 827 547
rect 823 541 827 542
rect 879 546 883 547
rect 879 541 883 542
rect 935 546 939 547
rect 935 541 939 542
rect 943 546 947 547
rect 943 541 947 542
rect 991 546 995 547
rect 991 541 995 542
rect 1007 546 1011 547
rect 1007 541 1011 542
rect 1047 546 1051 547
rect 1047 541 1051 542
rect 1071 546 1075 547
rect 1071 541 1075 542
rect 1103 546 1107 547
rect 1103 541 1107 542
rect 1127 546 1131 547
rect 1127 541 1131 542
rect 1159 546 1163 547
rect 1159 541 1163 542
rect 1183 546 1187 547
rect 1183 541 1187 542
rect 1215 546 1219 547
rect 1215 541 1219 542
rect 1231 546 1235 547
rect 1231 541 1235 542
rect 1271 546 1275 547
rect 1271 541 1275 542
rect 1279 546 1283 547
rect 1279 541 1283 542
rect 1327 546 1331 547
rect 1327 541 1331 542
rect 1335 546 1339 547
rect 1335 541 1339 542
rect 1383 546 1387 547
rect 1383 541 1387 542
rect 1391 546 1395 547
rect 1391 541 1395 542
rect 1447 546 1451 547
rect 1447 541 1451 542
rect 1511 546 1515 547
rect 1511 541 1515 542
rect 1575 546 1579 547
rect 1575 541 1579 542
rect 1623 546 1627 547
rect 1623 541 1627 542
rect 1663 546 1667 547
rect 1663 541 1667 542
rect 112 533 114 541
rect 110 532 116 533
rect 110 528 111 532
rect 115 528 116 532
rect 136 531 138 541
rect 168 531 170 541
rect 200 531 202 541
rect 232 531 234 541
rect 280 531 282 541
rect 328 531 330 541
rect 376 531 378 541
rect 432 531 434 541
rect 496 531 498 541
rect 560 531 562 541
rect 624 531 626 541
rect 688 531 690 541
rect 752 531 754 541
rect 816 531 818 541
rect 880 531 882 541
rect 944 531 946 541
rect 1008 531 1010 541
rect 1072 531 1074 541
rect 1128 531 1130 541
rect 1184 531 1186 541
rect 1232 531 1234 541
rect 1280 531 1282 541
rect 1336 531 1338 541
rect 1392 531 1394 541
rect 1448 531 1450 541
rect 1512 531 1514 541
rect 1576 531 1578 541
rect 1624 531 1626 541
rect 1664 533 1666 541
rect 1662 532 1668 533
rect 110 527 116 528
rect 134 530 140 531
rect 134 526 135 530
rect 139 526 140 530
rect 134 525 140 526
rect 166 530 172 531
rect 166 526 167 530
rect 171 526 172 530
rect 166 525 172 526
rect 198 530 204 531
rect 198 526 199 530
rect 203 526 204 530
rect 198 525 204 526
rect 230 530 236 531
rect 230 526 231 530
rect 235 526 236 530
rect 230 525 236 526
rect 278 530 284 531
rect 278 526 279 530
rect 283 526 284 530
rect 278 525 284 526
rect 326 530 332 531
rect 326 526 327 530
rect 331 526 332 530
rect 326 525 332 526
rect 374 530 380 531
rect 374 526 375 530
rect 379 526 380 530
rect 374 525 380 526
rect 430 530 436 531
rect 430 526 431 530
rect 435 526 436 530
rect 430 525 436 526
rect 494 530 500 531
rect 494 526 495 530
rect 499 526 500 530
rect 494 525 500 526
rect 558 530 564 531
rect 558 526 559 530
rect 563 526 564 530
rect 558 525 564 526
rect 622 530 628 531
rect 622 526 623 530
rect 627 526 628 530
rect 622 525 628 526
rect 686 530 692 531
rect 686 526 687 530
rect 691 526 692 530
rect 686 525 692 526
rect 750 530 756 531
rect 750 526 751 530
rect 755 526 756 530
rect 750 525 756 526
rect 814 530 820 531
rect 814 526 815 530
rect 819 526 820 530
rect 814 525 820 526
rect 878 530 884 531
rect 878 526 879 530
rect 883 526 884 530
rect 878 525 884 526
rect 942 530 948 531
rect 942 526 943 530
rect 947 526 948 530
rect 942 525 948 526
rect 1006 530 1012 531
rect 1006 526 1007 530
rect 1011 526 1012 530
rect 1006 525 1012 526
rect 1070 530 1076 531
rect 1070 526 1071 530
rect 1075 526 1076 530
rect 1070 525 1076 526
rect 1126 530 1132 531
rect 1126 526 1127 530
rect 1131 526 1132 530
rect 1126 525 1132 526
rect 1182 530 1188 531
rect 1182 526 1183 530
rect 1187 526 1188 530
rect 1182 525 1188 526
rect 1230 530 1236 531
rect 1230 526 1231 530
rect 1235 526 1236 530
rect 1230 525 1236 526
rect 1278 530 1284 531
rect 1278 526 1279 530
rect 1283 526 1284 530
rect 1278 525 1284 526
rect 1334 530 1340 531
rect 1334 526 1335 530
rect 1339 526 1340 530
rect 1334 525 1340 526
rect 1390 530 1396 531
rect 1390 526 1391 530
rect 1395 526 1396 530
rect 1390 525 1396 526
rect 1446 530 1452 531
rect 1446 526 1447 530
rect 1451 526 1452 530
rect 1446 525 1452 526
rect 1510 530 1516 531
rect 1510 526 1511 530
rect 1515 526 1516 530
rect 1510 525 1516 526
rect 1574 530 1580 531
rect 1574 526 1575 530
rect 1579 526 1580 530
rect 1574 525 1580 526
rect 1622 530 1628 531
rect 1622 526 1623 530
rect 1627 526 1628 530
rect 1662 528 1663 532
rect 1667 528 1668 532
rect 1662 527 1668 528
rect 1622 525 1628 526
rect 110 515 116 516
rect 110 511 111 515
rect 115 511 116 515
rect 1662 515 1668 516
rect 110 510 116 511
rect 134 513 140 514
rect 112 507 114 510
rect 134 509 135 513
rect 139 509 140 513
rect 134 508 140 509
rect 166 513 172 514
rect 166 509 167 513
rect 171 509 172 513
rect 166 508 172 509
rect 198 513 204 514
rect 198 509 199 513
rect 203 509 204 513
rect 198 508 204 509
rect 230 513 236 514
rect 230 509 231 513
rect 235 509 236 513
rect 230 508 236 509
rect 278 513 284 514
rect 278 509 279 513
rect 283 509 284 513
rect 278 508 284 509
rect 326 513 332 514
rect 326 509 327 513
rect 331 509 332 513
rect 326 508 332 509
rect 374 513 380 514
rect 374 509 375 513
rect 379 509 380 513
rect 374 508 380 509
rect 430 513 436 514
rect 430 509 431 513
rect 435 509 436 513
rect 430 508 436 509
rect 494 513 500 514
rect 494 509 495 513
rect 499 509 500 513
rect 494 508 500 509
rect 558 513 564 514
rect 558 509 559 513
rect 563 509 564 513
rect 558 508 564 509
rect 622 513 628 514
rect 622 509 623 513
rect 627 509 628 513
rect 622 508 628 509
rect 686 513 692 514
rect 686 509 687 513
rect 691 509 692 513
rect 686 508 692 509
rect 750 513 756 514
rect 750 509 751 513
rect 755 509 756 513
rect 750 508 756 509
rect 814 513 820 514
rect 814 509 815 513
rect 819 509 820 513
rect 814 508 820 509
rect 878 513 884 514
rect 878 509 879 513
rect 883 509 884 513
rect 878 508 884 509
rect 942 513 948 514
rect 942 509 943 513
rect 947 509 948 513
rect 942 508 948 509
rect 1006 513 1012 514
rect 1006 509 1007 513
rect 1011 509 1012 513
rect 1006 508 1012 509
rect 1070 513 1076 514
rect 1070 509 1071 513
rect 1075 509 1076 513
rect 1070 508 1076 509
rect 1126 513 1132 514
rect 1126 509 1127 513
rect 1131 509 1132 513
rect 1126 508 1132 509
rect 1182 513 1188 514
rect 1182 509 1183 513
rect 1187 509 1188 513
rect 1182 508 1188 509
rect 1230 513 1236 514
rect 1230 509 1231 513
rect 1235 509 1236 513
rect 1230 508 1236 509
rect 1278 513 1284 514
rect 1278 509 1279 513
rect 1283 509 1284 513
rect 1278 508 1284 509
rect 1334 513 1340 514
rect 1334 509 1335 513
rect 1339 509 1340 513
rect 1334 508 1340 509
rect 1390 513 1396 514
rect 1390 509 1391 513
rect 1395 509 1396 513
rect 1390 508 1396 509
rect 1446 513 1452 514
rect 1446 509 1447 513
rect 1451 509 1452 513
rect 1446 508 1452 509
rect 1510 513 1516 514
rect 1510 509 1511 513
rect 1515 509 1516 513
rect 1510 508 1516 509
rect 1574 513 1580 514
rect 1574 509 1575 513
rect 1579 509 1580 513
rect 1574 508 1580 509
rect 1622 513 1628 514
rect 1622 509 1623 513
rect 1627 509 1628 513
rect 1662 511 1663 515
rect 1667 511 1668 515
rect 1662 510 1668 511
rect 1622 508 1628 509
rect 111 506 115 507
rect 111 501 115 502
rect 135 506 139 508
rect 112 498 114 501
rect 135 500 139 502
rect 167 506 171 508
rect 167 500 171 502
rect 199 506 203 508
rect 199 500 203 502
rect 231 506 235 508
rect 231 501 235 502
rect 239 506 243 507
rect 239 500 243 502
rect 279 506 283 508
rect 279 501 283 502
rect 287 506 291 507
rect 287 500 291 502
rect 327 506 331 508
rect 327 500 331 502
rect 375 506 379 508
rect 375 500 379 502
rect 423 506 427 507
rect 423 500 427 502
rect 431 506 435 508
rect 431 501 435 502
rect 479 506 483 507
rect 479 500 483 502
rect 495 506 499 508
rect 495 501 499 502
rect 543 506 547 507
rect 543 500 547 502
rect 559 506 563 508
rect 559 501 563 502
rect 615 506 619 507
rect 615 500 619 502
rect 623 506 627 508
rect 623 501 627 502
rect 687 506 691 508
rect 687 501 691 502
rect 695 506 699 507
rect 695 500 699 502
rect 751 506 755 508
rect 751 501 755 502
rect 775 506 779 507
rect 775 500 779 502
rect 815 506 819 508
rect 815 501 819 502
rect 847 506 851 507
rect 847 500 851 502
rect 879 506 883 508
rect 879 501 883 502
rect 919 506 923 507
rect 919 500 923 502
rect 943 506 947 508
rect 943 501 947 502
rect 983 506 987 507
rect 983 500 987 502
rect 1007 506 1011 508
rect 1007 501 1011 502
rect 1039 506 1043 507
rect 1039 500 1043 502
rect 1071 506 1075 508
rect 1071 501 1075 502
rect 1095 506 1099 507
rect 1095 500 1099 502
rect 1127 506 1131 508
rect 1127 501 1131 502
rect 1143 506 1147 507
rect 1143 500 1147 502
rect 1183 506 1187 508
rect 1183 501 1187 502
rect 1191 506 1195 507
rect 1191 500 1195 502
rect 1231 506 1235 508
rect 1231 501 1235 502
rect 1239 506 1243 507
rect 1239 500 1243 502
rect 1279 506 1283 508
rect 1279 501 1283 502
rect 1287 506 1291 507
rect 1287 500 1291 502
rect 1335 506 1339 508
rect 1335 500 1339 502
rect 1383 506 1387 507
rect 1383 500 1387 502
rect 1391 506 1395 508
rect 1391 501 1395 502
rect 1431 506 1435 507
rect 1431 500 1435 502
rect 1447 506 1451 508
rect 1447 501 1451 502
rect 1479 506 1483 507
rect 1479 500 1483 502
rect 1511 506 1515 508
rect 1511 501 1515 502
rect 1535 506 1539 507
rect 1535 500 1539 502
rect 1575 506 1579 508
rect 1575 501 1579 502
rect 1591 506 1595 507
rect 1591 500 1595 502
rect 1623 506 1627 508
rect 1664 507 1666 510
rect 1623 500 1627 502
rect 1663 506 1667 507
rect 1663 501 1667 502
rect 134 499 140 500
rect 110 497 116 498
rect 110 493 111 497
rect 115 493 116 497
rect 134 495 135 499
rect 139 495 140 499
rect 134 494 140 495
rect 166 499 172 500
rect 166 495 167 499
rect 171 495 172 499
rect 166 494 172 495
rect 198 499 204 500
rect 198 495 199 499
rect 203 495 204 499
rect 198 494 204 495
rect 238 499 244 500
rect 238 495 239 499
rect 243 495 244 499
rect 238 494 244 495
rect 286 499 292 500
rect 286 495 287 499
rect 291 495 292 499
rect 286 494 292 495
rect 326 499 332 500
rect 326 495 327 499
rect 331 495 332 499
rect 326 494 332 495
rect 374 499 380 500
rect 374 495 375 499
rect 379 495 380 499
rect 374 494 380 495
rect 422 499 428 500
rect 422 495 423 499
rect 427 495 428 499
rect 422 494 428 495
rect 478 499 484 500
rect 478 495 479 499
rect 483 495 484 499
rect 478 494 484 495
rect 542 499 548 500
rect 542 495 543 499
rect 547 495 548 499
rect 542 494 548 495
rect 614 499 620 500
rect 614 495 615 499
rect 619 495 620 499
rect 614 494 620 495
rect 694 499 700 500
rect 694 495 695 499
rect 699 495 700 499
rect 694 494 700 495
rect 774 499 780 500
rect 774 495 775 499
rect 779 495 780 499
rect 774 494 780 495
rect 846 499 852 500
rect 846 495 847 499
rect 851 495 852 499
rect 846 494 852 495
rect 918 499 924 500
rect 918 495 919 499
rect 923 495 924 499
rect 918 494 924 495
rect 982 499 988 500
rect 982 495 983 499
rect 987 495 988 499
rect 982 494 988 495
rect 1038 499 1044 500
rect 1038 495 1039 499
rect 1043 495 1044 499
rect 1038 494 1044 495
rect 1094 499 1100 500
rect 1094 495 1095 499
rect 1099 495 1100 499
rect 1094 494 1100 495
rect 1142 499 1148 500
rect 1142 495 1143 499
rect 1147 495 1148 499
rect 1142 494 1148 495
rect 1190 499 1196 500
rect 1190 495 1191 499
rect 1195 495 1196 499
rect 1190 494 1196 495
rect 1238 499 1244 500
rect 1238 495 1239 499
rect 1243 495 1244 499
rect 1238 494 1244 495
rect 1286 499 1292 500
rect 1286 495 1287 499
rect 1291 495 1292 499
rect 1286 494 1292 495
rect 1334 499 1340 500
rect 1334 495 1335 499
rect 1339 495 1340 499
rect 1334 494 1340 495
rect 1382 499 1388 500
rect 1382 495 1383 499
rect 1387 495 1388 499
rect 1382 494 1388 495
rect 1430 499 1436 500
rect 1430 495 1431 499
rect 1435 495 1436 499
rect 1430 494 1436 495
rect 1478 499 1484 500
rect 1478 495 1479 499
rect 1483 495 1484 499
rect 1478 494 1484 495
rect 1534 499 1540 500
rect 1534 495 1535 499
rect 1539 495 1540 499
rect 1534 494 1540 495
rect 1590 499 1596 500
rect 1590 495 1591 499
rect 1595 495 1596 499
rect 1590 494 1596 495
rect 1622 499 1628 500
rect 1622 495 1623 499
rect 1627 495 1628 499
rect 1664 498 1666 501
rect 1622 494 1628 495
rect 1662 497 1668 498
rect 110 492 116 493
rect 1662 493 1663 497
rect 1667 493 1668 497
rect 1662 492 1668 493
rect 134 482 140 483
rect 110 480 116 481
rect 110 476 111 480
rect 115 476 116 480
rect 134 478 135 482
rect 139 478 140 482
rect 134 477 140 478
rect 166 482 172 483
rect 166 478 167 482
rect 171 478 172 482
rect 166 477 172 478
rect 198 482 204 483
rect 198 478 199 482
rect 203 478 204 482
rect 198 477 204 478
rect 238 482 244 483
rect 238 478 239 482
rect 243 478 244 482
rect 238 477 244 478
rect 286 482 292 483
rect 286 478 287 482
rect 291 478 292 482
rect 286 477 292 478
rect 326 482 332 483
rect 326 478 327 482
rect 331 478 332 482
rect 326 477 332 478
rect 374 482 380 483
rect 374 478 375 482
rect 379 478 380 482
rect 374 477 380 478
rect 422 482 428 483
rect 422 478 423 482
rect 427 478 428 482
rect 422 477 428 478
rect 478 482 484 483
rect 478 478 479 482
rect 483 478 484 482
rect 478 477 484 478
rect 542 482 548 483
rect 542 478 543 482
rect 547 478 548 482
rect 542 477 548 478
rect 614 482 620 483
rect 614 478 615 482
rect 619 478 620 482
rect 614 477 620 478
rect 694 482 700 483
rect 694 478 695 482
rect 699 478 700 482
rect 694 477 700 478
rect 774 482 780 483
rect 774 478 775 482
rect 779 478 780 482
rect 774 477 780 478
rect 846 482 852 483
rect 846 478 847 482
rect 851 478 852 482
rect 846 477 852 478
rect 918 482 924 483
rect 918 478 919 482
rect 923 478 924 482
rect 918 477 924 478
rect 982 482 988 483
rect 982 478 983 482
rect 987 478 988 482
rect 982 477 988 478
rect 1038 482 1044 483
rect 1038 478 1039 482
rect 1043 478 1044 482
rect 1038 477 1044 478
rect 1094 482 1100 483
rect 1094 478 1095 482
rect 1099 478 1100 482
rect 1094 477 1100 478
rect 1142 482 1148 483
rect 1142 478 1143 482
rect 1147 478 1148 482
rect 1142 477 1148 478
rect 1190 482 1196 483
rect 1190 478 1191 482
rect 1195 478 1196 482
rect 1190 477 1196 478
rect 1238 482 1244 483
rect 1238 478 1239 482
rect 1243 478 1244 482
rect 1238 477 1244 478
rect 1286 482 1292 483
rect 1286 478 1287 482
rect 1291 478 1292 482
rect 1286 477 1292 478
rect 1334 482 1340 483
rect 1334 478 1335 482
rect 1339 478 1340 482
rect 1334 477 1340 478
rect 1382 482 1388 483
rect 1382 478 1383 482
rect 1387 478 1388 482
rect 1382 477 1388 478
rect 1430 482 1436 483
rect 1430 478 1431 482
rect 1435 478 1436 482
rect 1430 477 1436 478
rect 1478 482 1484 483
rect 1478 478 1479 482
rect 1483 478 1484 482
rect 1478 477 1484 478
rect 1534 482 1540 483
rect 1534 478 1535 482
rect 1539 478 1540 482
rect 1534 477 1540 478
rect 1590 482 1596 483
rect 1590 478 1591 482
rect 1595 478 1596 482
rect 1590 477 1596 478
rect 1622 482 1628 483
rect 1622 478 1623 482
rect 1627 478 1628 482
rect 1622 477 1628 478
rect 1662 480 1668 481
rect 110 475 116 476
rect 112 467 114 475
rect 136 467 138 477
rect 168 467 170 477
rect 200 467 202 477
rect 240 467 242 477
rect 288 467 290 477
rect 328 467 330 477
rect 376 467 378 477
rect 424 467 426 477
rect 480 467 482 477
rect 544 467 546 477
rect 616 467 618 477
rect 696 467 698 477
rect 776 467 778 477
rect 848 467 850 477
rect 920 467 922 477
rect 984 467 986 477
rect 1040 467 1042 477
rect 1096 467 1098 477
rect 1144 467 1146 477
rect 1192 467 1194 477
rect 1240 467 1242 477
rect 1288 467 1290 477
rect 1336 467 1338 477
rect 1384 467 1386 477
rect 1432 467 1434 477
rect 1480 467 1482 477
rect 1536 467 1538 477
rect 1592 467 1594 477
rect 1624 467 1626 477
rect 1662 476 1663 480
rect 1667 476 1668 480
rect 1662 475 1668 476
rect 1664 467 1666 475
rect 111 466 115 467
rect 111 461 115 462
rect 135 466 139 467
rect 135 461 139 462
rect 151 466 155 467
rect 151 461 155 462
rect 167 466 171 467
rect 167 461 171 462
rect 199 466 203 467
rect 199 461 203 462
rect 207 466 211 467
rect 207 461 211 462
rect 239 466 243 467
rect 239 461 243 462
rect 255 466 259 467
rect 255 461 259 462
rect 287 466 291 467
rect 287 461 291 462
rect 311 466 315 467
rect 311 461 315 462
rect 327 466 331 467
rect 327 461 331 462
rect 367 466 371 467
rect 367 461 371 462
rect 375 466 379 467
rect 375 461 379 462
rect 423 466 427 467
rect 423 461 427 462
rect 439 466 443 467
rect 439 461 443 462
rect 479 466 483 467
rect 479 461 483 462
rect 519 466 523 467
rect 519 461 523 462
rect 543 466 547 467
rect 543 461 547 462
rect 599 466 603 467
rect 599 461 603 462
rect 615 466 619 467
rect 615 461 619 462
rect 679 466 683 467
rect 679 461 683 462
rect 695 466 699 467
rect 695 461 699 462
rect 759 466 763 467
rect 759 461 763 462
rect 775 466 779 467
rect 775 461 779 462
rect 839 466 843 467
rect 839 461 843 462
rect 847 466 851 467
rect 847 461 851 462
rect 911 466 915 467
rect 911 461 915 462
rect 919 466 923 467
rect 919 461 923 462
rect 983 466 987 467
rect 983 461 987 462
rect 1039 466 1043 467
rect 1039 461 1043 462
rect 1055 466 1059 467
rect 1055 461 1059 462
rect 1095 466 1099 467
rect 1095 461 1099 462
rect 1127 466 1131 467
rect 1127 461 1131 462
rect 1143 466 1147 467
rect 1143 461 1147 462
rect 1191 466 1195 467
rect 1191 461 1195 462
rect 1199 466 1203 467
rect 1199 461 1203 462
rect 1239 466 1243 467
rect 1239 461 1243 462
rect 1263 466 1267 467
rect 1263 461 1267 462
rect 1287 466 1291 467
rect 1287 461 1291 462
rect 1319 466 1323 467
rect 1319 461 1323 462
rect 1335 466 1339 467
rect 1335 461 1339 462
rect 1375 466 1379 467
rect 1375 461 1379 462
rect 1383 466 1387 467
rect 1383 461 1387 462
rect 1431 466 1435 467
rect 1431 461 1435 462
rect 1479 466 1483 467
rect 1479 461 1483 462
rect 1495 466 1499 467
rect 1495 461 1499 462
rect 1535 466 1539 467
rect 1535 461 1539 462
rect 1591 466 1595 467
rect 1591 461 1595 462
rect 1623 466 1627 467
rect 1623 461 1627 462
rect 1663 466 1667 467
rect 1663 461 1667 462
rect 112 453 114 461
rect 110 452 116 453
rect 110 448 111 452
rect 115 448 116 452
rect 152 451 154 461
rect 208 451 210 461
rect 256 451 258 461
rect 312 451 314 461
rect 368 451 370 461
rect 440 451 442 461
rect 520 451 522 461
rect 600 451 602 461
rect 680 451 682 461
rect 760 451 762 461
rect 840 451 842 461
rect 912 451 914 461
rect 984 451 986 461
rect 1056 451 1058 461
rect 1128 451 1130 461
rect 1200 451 1202 461
rect 1264 451 1266 461
rect 1320 451 1322 461
rect 1376 451 1378 461
rect 1432 451 1434 461
rect 1496 451 1498 461
rect 1664 453 1666 461
rect 1662 452 1668 453
rect 110 447 116 448
rect 150 450 156 451
rect 150 446 151 450
rect 155 446 156 450
rect 150 445 156 446
rect 206 450 212 451
rect 206 446 207 450
rect 211 446 212 450
rect 206 445 212 446
rect 254 450 260 451
rect 254 446 255 450
rect 259 446 260 450
rect 254 445 260 446
rect 310 450 316 451
rect 310 446 311 450
rect 315 446 316 450
rect 310 445 316 446
rect 366 450 372 451
rect 366 446 367 450
rect 371 446 372 450
rect 366 445 372 446
rect 438 450 444 451
rect 438 446 439 450
rect 443 446 444 450
rect 438 445 444 446
rect 518 450 524 451
rect 518 446 519 450
rect 523 446 524 450
rect 518 445 524 446
rect 598 450 604 451
rect 598 446 599 450
rect 603 446 604 450
rect 598 445 604 446
rect 678 450 684 451
rect 678 446 679 450
rect 683 446 684 450
rect 678 445 684 446
rect 758 450 764 451
rect 758 446 759 450
rect 763 446 764 450
rect 758 445 764 446
rect 838 450 844 451
rect 838 446 839 450
rect 843 446 844 450
rect 838 445 844 446
rect 910 450 916 451
rect 910 446 911 450
rect 915 446 916 450
rect 910 445 916 446
rect 982 450 988 451
rect 982 446 983 450
rect 987 446 988 450
rect 982 445 988 446
rect 1054 450 1060 451
rect 1054 446 1055 450
rect 1059 446 1060 450
rect 1054 445 1060 446
rect 1126 450 1132 451
rect 1126 446 1127 450
rect 1131 446 1132 450
rect 1126 445 1132 446
rect 1198 450 1204 451
rect 1198 446 1199 450
rect 1203 446 1204 450
rect 1198 445 1204 446
rect 1262 450 1268 451
rect 1262 446 1263 450
rect 1267 446 1268 450
rect 1262 445 1268 446
rect 1318 450 1324 451
rect 1318 446 1319 450
rect 1323 446 1324 450
rect 1318 445 1324 446
rect 1374 450 1380 451
rect 1374 446 1375 450
rect 1379 446 1380 450
rect 1374 445 1380 446
rect 1430 450 1436 451
rect 1430 446 1431 450
rect 1435 446 1436 450
rect 1430 445 1436 446
rect 1494 450 1500 451
rect 1494 446 1495 450
rect 1499 446 1500 450
rect 1662 448 1663 452
rect 1667 448 1668 452
rect 1662 447 1668 448
rect 1494 445 1500 446
rect 110 435 116 436
rect 110 431 111 435
rect 115 431 116 435
rect 1662 435 1668 436
rect 110 430 116 431
rect 150 433 156 434
rect 112 427 114 430
rect 150 429 151 433
rect 155 429 156 433
rect 150 428 156 429
rect 206 433 212 434
rect 206 429 207 433
rect 211 429 212 433
rect 206 428 212 429
rect 254 433 260 434
rect 254 429 255 433
rect 259 429 260 433
rect 254 428 260 429
rect 310 433 316 434
rect 310 429 311 433
rect 315 429 316 433
rect 310 428 316 429
rect 366 433 372 434
rect 366 429 367 433
rect 371 429 372 433
rect 366 428 372 429
rect 438 433 444 434
rect 438 429 439 433
rect 443 429 444 433
rect 438 428 444 429
rect 518 433 524 434
rect 518 429 519 433
rect 523 429 524 433
rect 518 428 524 429
rect 598 433 604 434
rect 598 429 599 433
rect 603 429 604 433
rect 598 428 604 429
rect 678 433 684 434
rect 678 429 679 433
rect 683 429 684 433
rect 678 428 684 429
rect 758 433 764 434
rect 758 429 759 433
rect 763 429 764 433
rect 758 428 764 429
rect 838 433 844 434
rect 838 429 839 433
rect 843 429 844 433
rect 838 428 844 429
rect 910 433 916 434
rect 910 429 911 433
rect 915 429 916 433
rect 910 428 916 429
rect 982 433 988 434
rect 982 429 983 433
rect 987 429 988 433
rect 982 428 988 429
rect 1054 433 1060 434
rect 1054 429 1055 433
rect 1059 429 1060 433
rect 1054 428 1060 429
rect 1126 433 1132 434
rect 1126 429 1127 433
rect 1131 429 1132 433
rect 1126 428 1132 429
rect 1198 433 1204 434
rect 1198 429 1199 433
rect 1203 429 1204 433
rect 1198 428 1204 429
rect 1262 433 1268 434
rect 1262 429 1263 433
rect 1267 429 1268 433
rect 1262 428 1268 429
rect 1318 433 1324 434
rect 1318 429 1319 433
rect 1323 429 1324 433
rect 1318 428 1324 429
rect 1374 433 1380 434
rect 1374 429 1375 433
rect 1379 429 1380 433
rect 1374 428 1380 429
rect 1430 433 1436 434
rect 1430 429 1431 433
rect 1435 429 1436 433
rect 1430 428 1436 429
rect 1494 433 1500 434
rect 1494 429 1495 433
rect 1499 429 1500 433
rect 1662 431 1663 435
rect 1667 431 1668 435
rect 1662 430 1668 431
rect 1494 428 1500 429
rect 111 426 115 427
rect 111 421 115 422
rect 151 426 155 428
rect 151 421 155 422
rect 175 426 179 427
rect 112 418 114 421
rect 175 420 179 422
rect 207 426 211 428
rect 207 421 211 422
rect 223 426 227 427
rect 223 420 227 422
rect 255 426 259 428
rect 255 421 259 422
rect 271 426 275 427
rect 271 420 275 422
rect 311 426 315 428
rect 311 421 315 422
rect 319 426 323 427
rect 319 420 323 422
rect 367 426 371 428
rect 367 420 371 422
rect 415 426 419 427
rect 415 420 419 422
rect 439 426 443 428
rect 439 421 443 422
rect 471 426 475 427
rect 471 420 475 422
rect 519 426 523 428
rect 519 421 523 422
rect 527 426 531 427
rect 527 420 531 422
rect 591 426 595 427
rect 591 420 595 422
rect 599 426 603 428
rect 599 421 603 422
rect 663 426 667 427
rect 663 420 667 422
rect 679 426 683 428
rect 679 421 683 422
rect 735 426 739 427
rect 735 420 739 422
rect 759 426 763 428
rect 759 421 763 422
rect 807 426 811 427
rect 807 420 811 422
rect 839 426 843 428
rect 839 421 843 422
rect 871 426 875 427
rect 871 420 875 422
rect 911 426 915 428
rect 911 421 915 422
rect 935 426 939 427
rect 935 420 939 422
rect 983 426 987 428
rect 983 421 987 422
rect 991 426 995 427
rect 991 420 995 422
rect 1039 426 1043 427
rect 1039 420 1043 422
rect 1055 426 1059 428
rect 1055 421 1059 422
rect 1087 426 1091 427
rect 1087 420 1091 422
rect 1127 426 1131 428
rect 1127 420 1131 422
rect 1167 426 1171 427
rect 1167 420 1171 422
rect 1199 426 1203 428
rect 1199 421 1203 422
rect 1207 426 1211 427
rect 1207 420 1211 422
rect 1247 426 1251 427
rect 1247 420 1251 422
rect 1263 426 1267 428
rect 1263 421 1267 422
rect 1287 426 1291 427
rect 1287 420 1291 422
rect 1319 426 1323 428
rect 1319 421 1323 422
rect 1335 426 1339 427
rect 1335 420 1339 422
rect 1375 426 1379 428
rect 1375 421 1379 422
rect 1383 426 1387 427
rect 1383 420 1387 422
rect 1431 426 1435 428
rect 1431 421 1435 422
rect 1495 426 1499 428
rect 1664 427 1666 430
rect 1495 421 1499 422
rect 1663 426 1667 427
rect 1663 421 1667 422
rect 174 419 180 420
rect 110 417 116 418
rect 110 413 111 417
rect 115 413 116 417
rect 174 415 175 419
rect 179 415 180 419
rect 174 414 180 415
rect 222 419 228 420
rect 222 415 223 419
rect 227 415 228 419
rect 222 414 228 415
rect 270 419 276 420
rect 270 415 271 419
rect 275 415 276 419
rect 270 414 276 415
rect 318 419 324 420
rect 318 415 319 419
rect 323 415 324 419
rect 318 414 324 415
rect 366 419 372 420
rect 366 415 367 419
rect 371 415 372 419
rect 366 414 372 415
rect 414 419 420 420
rect 414 415 415 419
rect 419 415 420 419
rect 414 414 420 415
rect 470 419 476 420
rect 470 415 471 419
rect 475 415 476 419
rect 470 414 476 415
rect 526 419 532 420
rect 526 415 527 419
rect 531 415 532 419
rect 526 414 532 415
rect 590 419 596 420
rect 590 415 591 419
rect 595 415 596 419
rect 590 414 596 415
rect 662 419 668 420
rect 662 415 663 419
rect 667 415 668 419
rect 662 414 668 415
rect 734 419 740 420
rect 734 415 735 419
rect 739 415 740 419
rect 734 414 740 415
rect 806 419 812 420
rect 806 415 807 419
rect 811 415 812 419
rect 806 414 812 415
rect 870 419 876 420
rect 870 415 871 419
rect 875 415 876 419
rect 870 414 876 415
rect 934 419 940 420
rect 934 415 935 419
rect 939 415 940 419
rect 934 414 940 415
rect 990 419 996 420
rect 990 415 991 419
rect 995 415 996 419
rect 990 414 996 415
rect 1038 419 1044 420
rect 1038 415 1039 419
rect 1043 415 1044 419
rect 1038 414 1044 415
rect 1086 419 1092 420
rect 1086 415 1087 419
rect 1091 415 1092 419
rect 1086 414 1092 415
rect 1126 419 1132 420
rect 1126 415 1127 419
rect 1131 415 1132 419
rect 1126 414 1132 415
rect 1166 419 1172 420
rect 1166 415 1167 419
rect 1171 415 1172 419
rect 1166 414 1172 415
rect 1206 419 1212 420
rect 1206 415 1207 419
rect 1211 415 1212 419
rect 1206 414 1212 415
rect 1246 419 1252 420
rect 1246 415 1247 419
rect 1251 415 1252 419
rect 1246 414 1252 415
rect 1286 419 1292 420
rect 1286 415 1287 419
rect 1291 415 1292 419
rect 1286 414 1292 415
rect 1334 419 1340 420
rect 1334 415 1335 419
rect 1339 415 1340 419
rect 1334 414 1340 415
rect 1382 419 1388 420
rect 1382 415 1383 419
rect 1387 415 1388 419
rect 1664 418 1666 421
rect 1382 414 1388 415
rect 1662 417 1668 418
rect 110 412 116 413
rect 1662 413 1663 417
rect 1667 413 1668 417
rect 1662 412 1668 413
rect 174 402 180 403
rect 110 400 116 401
rect 110 396 111 400
rect 115 396 116 400
rect 174 398 175 402
rect 179 398 180 402
rect 174 397 180 398
rect 222 402 228 403
rect 222 398 223 402
rect 227 398 228 402
rect 222 397 228 398
rect 270 402 276 403
rect 270 398 271 402
rect 275 398 276 402
rect 270 397 276 398
rect 318 402 324 403
rect 318 398 319 402
rect 323 398 324 402
rect 318 397 324 398
rect 366 402 372 403
rect 366 398 367 402
rect 371 398 372 402
rect 366 397 372 398
rect 414 402 420 403
rect 414 398 415 402
rect 419 398 420 402
rect 414 397 420 398
rect 470 402 476 403
rect 470 398 471 402
rect 475 398 476 402
rect 470 397 476 398
rect 526 402 532 403
rect 526 398 527 402
rect 531 398 532 402
rect 526 397 532 398
rect 590 402 596 403
rect 590 398 591 402
rect 595 398 596 402
rect 590 397 596 398
rect 662 402 668 403
rect 662 398 663 402
rect 667 398 668 402
rect 662 397 668 398
rect 734 402 740 403
rect 734 398 735 402
rect 739 398 740 402
rect 734 397 740 398
rect 806 402 812 403
rect 806 398 807 402
rect 811 398 812 402
rect 806 397 812 398
rect 870 402 876 403
rect 870 398 871 402
rect 875 398 876 402
rect 870 397 876 398
rect 934 402 940 403
rect 934 398 935 402
rect 939 398 940 402
rect 934 397 940 398
rect 990 402 996 403
rect 990 398 991 402
rect 995 398 996 402
rect 990 397 996 398
rect 1038 402 1044 403
rect 1038 398 1039 402
rect 1043 398 1044 402
rect 1038 397 1044 398
rect 1086 402 1092 403
rect 1086 398 1087 402
rect 1091 398 1092 402
rect 1086 397 1092 398
rect 1126 402 1132 403
rect 1126 398 1127 402
rect 1131 398 1132 402
rect 1126 397 1132 398
rect 1166 402 1172 403
rect 1166 398 1167 402
rect 1171 398 1172 402
rect 1166 397 1172 398
rect 1206 402 1212 403
rect 1206 398 1207 402
rect 1211 398 1212 402
rect 1206 397 1212 398
rect 1246 402 1252 403
rect 1246 398 1247 402
rect 1251 398 1252 402
rect 1246 397 1252 398
rect 1286 402 1292 403
rect 1286 398 1287 402
rect 1291 398 1292 402
rect 1286 397 1292 398
rect 1334 402 1340 403
rect 1334 398 1335 402
rect 1339 398 1340 402
rect 1334 397 1340 398
rect 1382 402 1388 403
rect 1382 398 1383 402
rect 1387 398 1388 402
rect 1382 397 1388 398
rect 1662 400 1668 401
rect 110 395 116 396
rect 112 383 114 395
rect 176 383 178 397
rect 224 383 226 397
rect 272 383 274 397
rect 320 383 322 397
rect 368 383 370 397
rect 416 383 418 397
rect 472 383 474 397
rect 528 383 530 397
rect 592 383 594 397
rect 664 383 666 397
rect 736 383 738 397
rect 808 383 810 397
rect 872 383 874 397
rect 936 383 938 397
rect 992 383 994 397
rect 1040 383 1042 397
rect 1088 383 1090 397
rect 1128 383 1130 397
rect 1168 383 1170 397
rect 1208 383 1210 397
rect 1248 383 1250 397
rect 1288 383 1290 397
rect 1336 383 1338 397
rect 1384 383 1386 397
rect 1662 396 1663 400
rect 1667 396 1668 400
rect 1662 395 1668 396
rect 1664 383 1666 395
rect 111 382 115 383
rect 111 377 115 378
rect 135 382 139 383
rect 135 377 139 378
rect 167 382 171 383
rect 167 377 171 378
rect 175 382 179 383
rect 175 377 179 378
rect 199 382 203 383
rect 199 377 203 378
rect 223 382 227 383
rect 223 377 227 378
rect 239 382 243 383
rect 239 377 243 378
rect 271 382 275 383
rect 271 377 275 378
rect 295 382 299 383
rect 295 377 299 378
rect 319 382 323 383
rect 319 377 323 378
rect 351 382 355 383
rect 351 377 355 378
rect 367 382 371 383
rect 367 377 371 378
rect 407 382 411 383
rect 407 377 411 378
rect 415 382 419 383
rect 415 377 419 378
rect 463 382 467 383
rect 463 377 467 378
rect 471 382 475 383
rect 471 377 475 378
rect 519 382 523 383
rect 519 377 523 378
rect 527 382 531 383
rect 527 377 531 378
rect 575 382 579 383
rect 575 377 579 378
rect 591 382 595 383
rect 591 377 595 378
rect 631 382 635 383
rect 631 377 635 378
rect 663 382 667 383
rect 663 377 667 378
rect 687 382 691 383
rect 687 377 691 378
rect 735 382 739 383
rect 735 377 739 378
rect 743 382 747 383
rect 743 377 747 378
rect 799 382 803 383
rect 799 377 803 378
rect 807 382 811 383
rect 807 377 811 378
rect 855 382 859 383
rect 855 377 859 378
rect 871 382 875 383
rect 871 377 875 378
rect 919 382 923 383
rect 919 377 923 378
rect 935 382 939 383
rect 935 377 939 378
rect 983 382 987 383
rect 983 377 987 378
rect 991 382 995 383
rect 991 377 995 378
rect 1039 382 1043 383
rect 1039 377 1043 378
rect 1087 382 1091 383
rect 1087 377 1091 378
rect 1095 382 1099 383
rect 1095 377 1099 378
rect 1127 382 1131 383
rect 1127 377 1131 378
rect 1151 382 1155 383
rect 1151 377 1155 378
rect 1167 382 1171 383
rect 1167 377 1171 378
rect 1207 382 1211 383
rect 1207 377 1211 378
rect 1247 382 1251 383
rect 1247 377 1251 378
rect 1255 382 1259 383
rect 1255 377 1259 378
rect 1287 382 1291 383
rect 1287 377 1291 378
rect 1303 382 1307 383
rect 1303 377 1307 378
rect 1335 382 1339 383
rect 1335 377 1339 378
rect 1351 382 1355 383
rect 1351 377 1355 378
rect 1383 382 1387 383
rect 1383 377 1387 378
rect 1399 382 1403 383
rect 1399 377 1403 378
rect 1447 382 1451 383
rect 1447 377 1451 378
rect 1495 382 1499 383
rect 1495 377 1499 378
rect 1543 382 1547 383
rect 1543 377 1547 378
rect 1591 382 1595 383
rect 1591 377 1595 378
rect 1623 382 1627 383
rect 1623 377 1627 378
rect 1663 382 1667 383
rect 1663 377 1667 378
rect 112 369 114 377
rect 110 368 116 369
rect 110 364 111 368
rect 115 364 116 368
rect 136 367 138 377
rect 168 367 170 377
rect 200 367 202 377
rect 240 367 242 377
rect 296 367 298 377
rect 352 367 354 377
rect 408 367 410 377
rect 464 367 466 377
rect 520 367 522 377
rect 576 367 578 377
rect 632 367 634 377
rect 688 367 690 377
rect 744 367 746 377
rect 800 367 802 377
rect 856 367 858 377
rect 920 367 922 377
rect 984 367 986 377
rect 1040 367 1042 377
rect 1096 367 1098 377
rect 1152 367 1154 377
rect 1208 367 1210 377
rect 1256 367 1258 377
rect 1304 367 1306 377
rect 1352 367 1354 377
rect 1400 367 1402 377
rect 1448 367 1450 377
rect 1496 367 1498 377
rect 1544 367 1546 377
rect 1592 367 1594 377
rect 1624 367 1626 377
rect 1664 369 1666 377
rect 1662 368 1668 369
rect 110 363 116 364
rect 134 366 140 367
rect 134 362 135 366
rect 139 362 140 366
rect 134 361 140 362
rect 166 366 172 367
rect 166 362 167 366
rect 171 362 172 366
rect 166 361 172 362
rect 198 366 204 367
rect 198 362 199 366
rect 203 362 204 366
rect 198 361 204 362
rect 238 366 244 367
rect 238 362 239 366
rect 243 362 244 366
rect 238 361 244 362
rect 294 366 300 367
rect 294 362 295 366
rect 299 362 300 366
rect 294 361 300 362
rect 350 366 356 367
rect 350 362 351 366
rect 355 362 356 366
rect 350 361 356 362
rect 406 366 412 367
rect 406 362 407 366
rect 411 362 412 366
rect 406 361 412 362
rect 462 366 468 367
rect 462 362 463 366
rect 467 362 468 366
rect 462 361 468 362
rect 518 366 524 367
rect 518 362 519 366
rect 523 362 524 366
rect 518 361 524 362
rect 574 366 580 367
rect 574 362 575 366
rect 579 362 580 366
rect 574 361 580 362
rect 630 366 636 367
rect 630 362 631 366
rect 635 362 636 366
rect 630 361 636 362
rect 686 366 692 367
rect 686 362 687 366
rect 691 362 692 366
rect 686 361 692 362
rect 742 366 748 367
rect 742 362 743 366
rect 747 362 748 366
rect 742 361 748 362
rect 798 366 804 367
rect 798 362 799 366
rect 803 362 804 366
rect 798 361 804 362
rect 854 366 860 367
rect 854 362 855 366
rect 859 362 860 366
rect 854 361 860 362
rect 918 366 924 367
rect 918 362 919 366
rect 923 362 924 366
rect 918 361 924 362
rect 982 366 988 367
rect 982 362 983 366
rect 987 362 988 366
rect 982 361 988 362
rect 1038 366 1044 367
rect 1038 362 1039 366
rect 1043 362 1044 366
rect 1038 361 1044 362
rect 1094 366 1100 367
rect 1094 362 1095 366
rect 1099 362 1100 366
rect 1094 361 1100 362
rect 1150 366 1156 367
rect 1150 362 1151 366
rect 1155 362 1156 366
rect 1150 361 1156 362
rect 1206 366 1212 367
rect 1206 362 1207 366
rect 1211 362 1212 366
rect 1206 361 1212 362
rect 1254 366 1260 367
rect 1254 362 1255 366
rect 1259 362 1260 366
rect 1254 361 1260 362
rect 1302 366 1308 367
rect 1302 362 1303 366
rect 1307 362 1308 366
rect 1302 361 1308 362
rect 1350 366 1356 367
rect 1350 362 1351 366
rect 1355 362 1356 366
rect 1350 361 1356 362
rect 1398 366 1404 367
rect 1398 362 1399 366
rect 1403 362 1404 366
rect 1398 361 1404 362
rect 1446 366 1452 367
rect 1446 362 1447 366
rect 1451 362 1452 366
rect 1446 361 1452 362
rect 1494 366 1500 367
rect 1494 362 1495 366
rect 1499 362 1500 366
rect 1494 361 1500 362
rect 1542 366 1548 367
rect 1542 362 1543 366
rect 1547 362 1548 366
rect 1542 361 1548 362
rect 1590 366 1596 367
rect 1590 362 1591 366
rect 1595 362 1596 366
rect 1590 361 1596 362
rect 1622 366 1628 367
rect 1622 362 1623 366
rect 1627 362 1628 366
rect 1662 364 1663 368
rect 1667 364 1668 368
rect 1662 363 1668 364
rect 1622 361 1628 362
rect 110 351 116 352
rect 110 347 111 351
rect 115 347 116 351
rect 1662 351 1668 352
rect 110 346 116 347
rect 134 349 140 350
rect 112 343 114 346
rect 134 345 135 349
rect 139 345 140 349
rect 134 344 140 345
rect 166 349 172 350
rect 166 345 167 349
rect 171 345 172 349
rect 166 344 172 345
rect 198 349 204 350
rect 198 345 199 349
rect 203 345 204 349
rect 198 344 204 345
rect 238 349 244 350
rect 238 345 239 349
rect 243 345 244 349
rect 238 344 244 345
rect 294 349 300 350
rect 294 345 295 349
rect 299 345 300 349
rect 294 344 300 345
rect 350 349 356 350
rect 350 345 351 349
rect 355 345 356 349
rect 350 344 356 345
rect 406 349 412 350
rect 406 345 407 349
rect 411 345 412 349
rect 406 344 412 345
rect 462 349 468 350
rect 462 345 463 349
rect 467 345 468 349
rect 462 344 468 345
rect 518 349 524 350
rect 518 345 519 349
rect 523 345 524 349
rect 518 344 524 345
rect 574 349 580 350
rect 574 345 575 349
rect 579 345 580 349
rect 574 344 580 345
rect 630 349 636 350
rect 630 345 631 349
rect 635 345 636 349
rect 630 344 636 345
rect 686 349 692 350
rect 686 345 687 349
rect 691 345 692 349
rect 686 344 692 345
rect 742 349 748 350
rect 742 345 743 349
rect 747 345 748 349
rect 742 344 748 345
rect 798 349 804 350
rect 798 345 799 349
rect 803 345 804 349
rect 798 344 804 345
rect 854 349 860 350
rect 854 345 855 349
rect 859 345 860 349
rect 854 344 860 345
rect 918 349 924 350
rect 918 345 919 349
rect 923 345 924 349
rect 918 344 924 345
rect 982 349 988 350
rect 982 345 983 349
rect 987 345 988 349
rect 982 344 988 345
rect 1038 349 1044 350
rect 1038 345 1039 349
rect 1043 345 1044 349
rect 1038 344 1044 345
rect 1094 349 1100 350
rect 1094 345 1095 349
rect 1099 345 1100 349
rect 1094 344 1100 345
rect 1150 349 1156 350
rect 1150 345 1151 349
rect 1155 345 1156 349
rect 1150 344 1156 345
rect 1206 349 1212 350
rect 1206 345 1207 349
rect 1211 345 1212 349
rect 1206 344 1212 345
rect 1254 349 1260 350
rect 1254 345 1255 349
rect 1259 345 1260 349
rect 1254 344 1260 345
rect 1302 349 1308 350
rect 1302 345 1303 349
rect 1307 345 1308 349
rect 1302 344 1308 345
rect 1350 349 1356 350
rect 1350 345 1351 349
rect 1355 345 1356 349
rect 1350 344 1356 345
rect 1398 349 1404 350
rect 1398 345 1399 349
rect 1403 345 1404 349
rect 1398 344 1404 345
rect 1446 349 1452 350
rect 1446 345 1447 349
rect 1451 345 1452 349
rect 1446 344 1452 345
rect 1494 349 1500 350
rect 1494 345 1495 349
rect 1499 345 1500 349
rect 1494 344 1500 345
rect 1542 349 1548 350
rect 1542 345 1543 349
rect 1547 345 1548 349
rect 1542 344 1548 345
rect 1590 349 1596 350
rect 1590 345 1591 349
rect 1595 345 1596 349
rect 1590 344 1596 345
rect 1622 349 1628 350
rect 1622 345 1623 349
rect 1627 345 1628 349
rect 1662 347 1663 351
rect 1667 347 1668 351
rect 1662 346 1668 347
rect 1622 344 1628 345
rect 111 342 115 343
rect 111 337 115 338
rect 135 342 139 344
rect 112 334 114 337
rect 135 336 139 338
rect 167 342 171 344
rect 167 336 171 338
rect 199 342 203 344
rect 199 337 203 338
rect 207 342 211 343
rect 207 336 211 338
rect 239 342 243 344
rect 239 337 243 338
rect 263 342 267 343
rect 263 336 267 338
rect 295 342 299 344
rect 295 337 299 338
rect 327 342 331 343
rect 327 336 331 338
rect 351 342 355 344
rect 351 337 355 338
rect 391 342 395 343
rect 391 336 395 338
rect 407 342 411 344
rect 407 337 411 338
rect 455 342 459 343
rect 455 336 459 338
rect 463 342 467 344
rect 463 337 467 338
rect 519 342 523 344
rect 519 336 523 338
rect 575 342 579 344
rect 575 336 579 338
rect 631 342 635 344
rect 631 336 635 338
rect 687 342 691 344
rect 687 336 691 338
rect 743 342 747 344
rect 743 337 747 338
rect 751 342 755 343
rect 751 336 755 338
rect 799 342 803 344
rect 799 337 803 338
rect 815 342 819 343
rect 815 336 819 338
rect 855 342 859 344
rect 855 337 859 338
rect 879 342 883 343
rect 879 336 883 338
rect 919 342 923 344
rect 919 337 923 338
rect 951 342 955 343
rect 951 336 955 338
rect 983 342 987 344
rect 983 337 987 338
rect 1031 342 1035 343
rect 1031 336 1035 338
rect 1039 342 1043 344
rect 1039 337 1043 338
rect 1095 342 1099 344
rect 1095 337 1099 338
rect 1111 342 1115 343
rect 1111 336 1115 338
rect 1151 342 1155 344
rect 1151 337 1155 338
rect 1191 342 1195 343
rect 1191 336 1195 338
rect 1207 342 1211 344
rect 1207 337 1211 338
rect 1255 342 1259 344
rect 1255 337 1259 338
rect 1271 342 1275 343
rect 1271 336 1275 338
rect 1303 342 1307 344
rect 1303 337 1307 338
rect 1343 342 1347 343
rect 1343 336 1347 338
rect 1351 342 1355 344
rect 1351 337 1355 338
rect 1399 342 1403 344
rect 1399 337 1403 338
rect 1407 342 1411 343
rect 1407 336 1411 338
rect 1447 342 1451 344
rect 1447 337 1451 338
rect 1463 342 1467 343
rect 1463 336 1467 338
rect 1495 342 1499 344
rect 1495 337 1499 338
rect 1519 342 1523 343
rect 1519 336 1523 338
rect 1543 342 1547 344
rect 1543 337 1547 338
rect 1583 342 1587 343
rect 1583 336 1587 338
rect 1591 342 1595 344
rect 1591 337 1595 338
rect 1623 342 1627 344
rect 1664 343 1666 346
rect 1623 336 1627 338
rect 1663 342 1667 343
rect 1663 337 1667 338
rect 134 335 140 336
rect 110 333 116 334
rect 110 329 111 333
rect 115 329 116 333
rect 134 331 135 335
rect 139 331 140 335
rect 134 330 140 331
rect 166 335 172 336
rect 166 331 167 335
rect 171 331 172 335
rect 166 330 172 331
rect 206 335 212 336
rect 206 331 207 335
rect 211 331 212 335
rect 206 330 212 331
rect 262 335 268 336
rect 262 331 263 335
rect 267 331 268 335
rect 262 330 268 331
rect 326 335 332 336
rect 326 331 327 335
rect 331 331 332 335
rect 326 330 332 331
rect 390 335 396 336
rect 390 331 391 335
rect 395 331 396 335
rect 390 330 396 331
rect 454 335 460 336
rect 454 331 455 335
rect 459 331 460 335
rect 454 330 460 331
rect 518 335 524 336
rect 518 331 519 335
rect 523 331 524 335
rect 518 330 524 331
rect 574 335 580 336
rect 574 331 575 335
rect 579 331 580 335
rect 574 330 580 331
rect 630 335 636 336
rect 630 331 631 335
rect 635 331 636 335
rect 630 330 636 331
rect 686 335 692 336
rect 686 331 687 335
rect 691 331 692 335
rect 686 330 692 331
rect 750 335 756 336
rect 750 331 751 335
rect 755 331 756 335
rect 750 330 756 331
rect 814 335 820 336
rect 814 331 815 335
rect 819 331 820 335
rect 814 330 820 331
rect 878 335 884 336
rect 878 331 879 335
rect 883 331 884 335
rect 878 330 884 331
rect 950 335 956 336
rect 950 331 951 335
rect 955 331 956 335
rect 950 330 956 331
rect 1030 335 1036 336
rect 1030 331 1031 335
rect 1035 331 1036 335
rect 1030 330 1036 331
rect 1110 335 1116 336
rect 1110 331 1111 335
rect 1115 331 1116 335
rect 1110 330 1116 331
rect 1190 335 1196 336
rect 1190 331 1191 335
rect 1195 331 1196 335
rect 1190 330 1196 331
rect 1270 335 1276 336
rect 1270 331 1271 335
rect 1275 331 1276 335
rect 1270 330 1276 331
rect 1342 335 1348 336
rect 1342 331 1343 335
rect 1347 331 1348 335
rect 1342 330 1348 331
rect 1406 335 1412 336
rect 1406 331 1407 335
rect 1411 331 1412 335
rect 1406 330 1412 331
rect 1462 335 1468 336
rect 1462 331 1463 335
rect 1467 331 1468 335
rect 1462 330 1468 331
rect 1518 335 1524 336
rect 1518 331 1519 335
rect 1523 331 1524 335
rect 1518 330 1524 331
rect 1582 335 1588 336
rect 1582 331 1583 335
rect 1587 331 1588 335
rect 1582 330 1588 331
rect 1622 335 1628 336
rect 1622 331 1623 335
rect 1627 331 1628 335
rect 1664 334 1666 337
rect 1622 330 1628 331
rect 1662 333 1668 334
rect 110 328 116 329
rect 1662 329 1663 333
rect 1667 329 1668 333
rect 1662 328 1668 329
rect 134 318 140 319
rect 110 316 116 317
rect 110 312 111 316
rect 115 312 116 316
rect 134 314 135 318
rect 139 314 140 318
rect 134 313 140 314
rect 166 318 172 319
rect 166 314 167 318
rect 171 314 172 318
rect 166 313 172 314
rect 206 318 212 319
rect 206 314 207 318
rect 211 314 212 318
rect 206 313 212 314
rect 262 318 268 319
rect 262 314 263 318
rect 267 314 268 318
rect 262 313 268 314
rect 326 318 332 319
rect 326 314 327 318
rect 331 314 332 318
rect 326 313 332 314
rect 390 318 396 319
rect 390 314 391 318
rect 395 314 396 318
rect 390 313 396 314
rect 454 318 460 319
rect 454 314 455 318
rect 459 314 460 318
rect 454 313 460 314
rect 518 318 524 319
rect 518 314 519 318
rect 523 314 524 318
rect 518 313 524 314
rect 574 318 580 319
rect 574 314 575 318
rect 579 314 580 318
rect 574 313 580 314
rect 630 318 636 319
rect 630 314 631 318
rect 635 314 636 318
rect 630 313 636 314
rect 686 318 692 319
rect 686 314 687 318
rect 691 314 692 318
rect 686 313 692 314
rect 750 318 756 319
rect 750 314 751 318
rect 755 314 756 318
rect 750 313 756 314
rect 814 318 820 319
rect 814 314 815 318
rect 819 314 820 318
rect 814 313 820 314
rect 878 318 884 319
rect 878 314 879 318
rect 883 314 884 318
rect 878 313 884 314
rect 950 318 956 319
rect 950 314 951 318
rect 955 314 956 318
rect 950 313 956 314
rect 1030 318 1036 319
rect 1030 314 1031 318
rect 1035 314 1036 318
rect 1030 313 1036 314
rect 1110 318 1116 319
rect 1110 314 1111 318
rect 1115 314 1116 318
rect 1110 313 1116 314
rect 1190 318 1196 319
rect 1190 314 1191 318
rect 1195 314 1196 318
rect 1190 313 1196 314
rect 1270 318 1276 319
rect 1270 314 1271 318
rect 1275 314 1276 318
rect 1270 313 1276 314
rect 1342 318 1348 319
rect 1342 314 1343 318
rect 1347 314 1348 318
rect 1342 313 1348 314
rect 1406 318 1412 319
rect 1406 314 1407 318
rect 1411 314 1412 318
rect 1406 313 1412 314
rect 1462 318 1468 319
rect 1462 314 1463 318
rect 1467 314 1468 318
rect 1462 313 1468 314
rect 1518 318 1524 319
rect 1518 314 1519 318
rect 1523 314 1524 318
rect 1518 313 1524 314
rect 1582 318 1588 319
rect 1582 314 1583 318
rect 1587 314 1588 318
rect 1582 313 1588 314
rect 1622 318 1628 319
rect 1622 314 1623 318
rect 1627 314 1628 318
rect 1622 313 1628 314
rect 1662 316 1668 317
rect 110 311 116 312
rect 112 303 114 311
rect 136 303 138 313
rect 168 303 170 313
rect 208 303 210 313
rect 264 303 266 313
rect 328 303 330 313
rect 392 303 394 313
rect 456 303 458 313
rect 520 303 522 313
rect 576 303 578 313
rect 632 303 634 313
rect 688 303 690 313
rect 752 303 754 313
rect 816 303 818 313
rect 880 303 882 313
rect 952 303 954 313
rect 1032 303 1034 313
rect 1112 303 1114 313
rect 1192 303 1194 313
rect 1272 303 1274 313
rect 1344 303 1346 313
rect 1408 303 1410 313
rect 1464 303 1466 313
rect 1520 303 1522 313
rect 1584 303 1586 313
rect 1624 303 1626 313
rect 1662 312 1663 316
rect 1667 312 1668 316
rect 1662 311 1668 312
rect 1664 303 1666 311
rect 111 302 115 303
rect 111 297 115 298
rect 135 302 139 303
rect 135 297 139 298
rect 167 302 171 303
rect 167 297 171 298
rect 207 302 211 303
rect 207 297 211 298
rect 231 302 235 303
rect 231 297 235 298
rect 263 302 267 303
rect 263 297 267 298
rect 295 302 299 303
rect 295 297 299 298
rect 327 302 331 303
rect 327 297 331 298
rect 367 302 371 303
rect 367 297 371 298
rect 391 302 395 303
rect 391 297 395 298
rect 439 302 443 303
rect 439 297 443 298
rect 455 302 459 303
rect 455 297 459 298
rect 503 302 507 303
rect 503 297 507 298
rect 519 302 523 303
rect 519 297 523 298
rect 567 302 571 303
rect 567 297 571 298
rect 575 302 579 303
rect 575 297 579 298
rect 631 302 635 303
rect 631 297 635 298
rect 687 302 691 303
rect 687 297 691 298
rect 743 302 747 303
rect 743 297 747 298
rect 751 302 755 303
rect 751 297 755 298
rect 807 302 811 303
rect 807 297 811 298
rect 815 302 819 303
rect 815 297 819 298
rect 879 302 883 303
rect 879 297 883 298
rect 951 302 955 303
rect 951 297 955 298
rect 1031 302 1035 303
rect 1031 297 1035 298
rect 1111 302 1115 303
rect 1111 297 1115 298
rect 1191 302 1195 303
rect 1191 297 1195 298
rect 1263 302 1267 303
rect 1263 297 1267 298
rect 1271 302 1275 303
rect 1271 297 1275 298
rect 1327 302 1331 303
rect 1327 297 1331 298
rect 1343 302 1347 303
rect 1343 297 1347 298
rect 1391 302 1395 303
rect 1391 297 1395 298
rect 1407 302 1411 303
rect 1407 297 1411 298
rect 1447 302 1451 303
rect 1447 297 1451 298
rect 1463 302 1467 303
rect 1463 297 1467 298
rect 1495 302 1499 303
rect 1495 297 1499 298
rect 1519 302 1523 303
rect 1519 297 1523 298
rect 1543 302 1547 303
rect 1543 297 1547 298
rect 1583 302 1587 303
rect 1583 297 1587 298
rect 1591 302 1595 303
rect 1591 297 1595 298
rect 1623 302 1627 303
rect 1623 297 1627 298
rect 1663 302 1667 303
rect 1663 297 1667 298
rect 112 289 114 297
rect 110 288 116 289
rect 110 284 111 288
rect 115 284 116 288
rect 136 287 138 297
rect 168 287 170 297
rect 232 287 234 297
rect 296 287 298 297
rect 368 287 370 297
rect 440 287 442 297
rect 504 287 506 297
rect 568 287 570 297
rect 632 287 634 297
rect 688 287 690 297
rect 744 287 746 297
rect 808 287 810 297
rect 880 287 882 297
rect 952 287 954 297
rect 1032 287 1034 297
rect 1112 287 1114 297
rect 1192 287 1194 297
rect 1264 287 1266 297
rect 1328 287 1330 297
rect 1392 287 1394 297
rect 1448 287 1450 297
rect 1496 287 1498 297
rect 1544 287 1546 297
rect 1592 287 1594 297
rect 1624 287 1626 297
rect 1664 289 1666 297
rect 1662 288 1668 289
rect 110 283 116 284
rect 134 286 140 287
rect 134 282 135 286
rect 139 282 140 286
rect 134 281 140 282
rect 166 286 172 287
rect 166 282 167 286
rect 171 282 172 286
rect 166 281 172 282
rect 230 286 236 287
rect 230 282 231 286
rect 235 282 236 286
rect 230 281 236 282
rect 294 286 300 287
rect 294 282 295 286
rect 299 282 300 286
rect 294 281 300 282
rect 366 286 372 287
rect 366 282 367 286
rect 371 282 372 286
rect 366 281 372 282
rect 438 286 444 287
rect 438 282 439 286
rect 443 282 444 286
rect 438 281 444 282
rect 502 286 508 287
rect 502 282 503 286
rect 507 282 508 286
rect 502 281 508 282
rect 566 286 572 287
rect 566 282 567 286
rect 571 282 572 286
rect 566 281 572 282
rect 630 286 636 287
rect 630 282 631 286
rect 635 282 636 286
rect 630 281 636 282
rect 686 286 692 287
rect 686 282 687 286
rect 691 282 692 286
rect 686 281 692 282
rect 742 286 748 287
rect 742 282 743 286
rect 747 282 748 286
rect 742 281 748 282
rect 806 286 812 287
rect 806 282 807 286
rect 811 282 812 286
rect 806 281 812 282
rect 878 286 884 287
rect 878 282 879 286
rect 883 282 884 286
rect 878 281 884 282
rect 950 286 956 287
rect 950 282 951 286
rect 955 282 956 286
rect 950 281 956 282
rect 1030 286 1036 287
rect 1030 282 1031 286
rect 1035 282 1036 286
rect 1030 281 1036 282
rect 1110 286 1116 287
rect 1110 282 1111 286
rect 1115 282 1116 286
rect 1110 281 1116 282
rect 1190 286 1196 287
rect 1190 282 1191 286
rect 1195 282 1196 286
rect 1190 281 1196 282
rect 1262 286 1268 287
rect 1262 282 1263 286
rect 1267 282 1268 286
rect 1262 281 1268 282
rect 1326 286 1332 287
rect 1326 282 1327 286
rect 1331 282 1332 286
rect 1326 281 1332 282
rect 1390 286 1396 287
rect 1390 282 1391 286
rect 1395 282 1396 286
rect 1390 281 1396 282
rect 1446 286 1452 287
rect 1446 282 1447 286
rect 1451 282 1452 286
rect 1446 281 1452 282
rect 1494 286 1500 287
rect 1494 282 1495 286
rect 1499 282 1500 286
rect 1494 281 1500 282
rect 1542 286 1548 287
rect 1542 282 1543 286
rect 1547 282 1548 286
rect 1542 281 1548 282
rect 1590 286 1596 287
rect 1590 282 1591 286
rect 1595 282 1596 286
rect 1590 281 1596 282
rect 1622 286 1628 287
rect 1622 282 1623 286
rect 1627 282 1628 286
rect 1662 284 1663 288
rect 1667 284 1668 288
rect 1662 283 1668 284
rect 1622 281 1628 282
rect 110 271 116 272
rect 110 267 111 271
rect 115 267 116 271
rect 1662 271 1668 272
rect 110 266 116 267
rect 134 269 140 270
rect 112 259 114 266
rect 134 265 135 269
rect 139 265 140 269
rect 134 264 140 265
rect 166 269 172 270
rect 166 265 167 269
rect 171 265 172 269
rect 166 264 172 265
rect 230 269 236 270
rect 230 265 231 269
rect 235 265 236 269
rect 230 264 236 265
rect 294 269 300 270
rect 294 265 295 269
rect 299 265 300 269
rect 294 264 300 265
rect 366 269 372 270
rect 366 265 367 269
rect 371 265 372 269
rect 366 264 372 265
rect 438 269 444 270
rect 438 265 439 269
rect 443 265 444 269
rect 438 264 444 265
rect 502 269 508 270
rect 502 265 503 269
rect 507 265 508 269
rect 502 264 508 265
rect 566 269 572 270
rect 566 265 567 269
rect 571 265 572 269
rect 566 264 572 265
rect 630 269 636 270
rect 630 265 631 269
rect 635 265 636 269
rect 630 264 636 265
rect 686 269 692 270
rect 686 265 687 269
rect 691 265 692 269
rect 686 264 692 265
rect 742 269 748 270
rect 742 265 743 269
rect 747 265 748 269
rect 742 264 748 265
rect 806 269 812 270
rect 806 265 807 269
rect 811 265 812 269
rect 806 264 812 265
rect 878 269 884 270
rect 878 265 879 269
rect 883 265 884 269
rect 878 264 884 265
rect 950 269 956 270
rect 950 265 951 269
rect 955 265 956 269
rect 950 264 956 265
rect 1030 269 1036 270
rect 1030 265 1031 269
rect 1035 265 1036 269
rect 1030 264 1036 265
rect 1110 269 1116 270
rect 1110 265 1111 269
rect 1115 265 1116 269
rect 1110 264 1116 265
rect 1190 269 1196 270
rect 1190 265 1191 269
rect 1195 265 1196 269
rect 1190 264 1196 265
rect 1262 269 1268 270
rect 1262 265 1263 269
rect 1267 265 1268 269
rect 1262 264 1268 265
rect 1326 269 1332 270
rect 1326 265 1327 269
rect 1331 265 1332 269
rect 1326 264 1332 265
rect 1390 269 1396 270
rect 1390 265 1391 269
rect 1395 265 1396 269
rect 1390 264 1396 265
rect 1446 269 1452 270
rect 1446 265 1447 269
rect 1451 265 1452 269
rect 1446 264 1452 265
rect 1494 269 1500 270
rect 1494 265 1495 269
rect 1499 265 1500 269
rect 1494 264 1500 265
rect 1542 269 1548 270
rect 1542 265 1543 269
rect 1547 265 1548 269
rect 1542 264 1548 265
rect 1590 269 1596 270
rect 1590 265 1591 269
rect 1595 265 1596 269
rect 1590 264 1596 265
rect 1622 269 1628 270
rect 1622 265 1623 269
rect 1627 265 1628 269
rect 1662 267 1663 271
rect 1667 267 1668 271
rect 1662 266 1668 267
rect 1622 264 1628 265
rect 136 259 138 264
rect 168 259 170 264
rect 232 259 234 264
rect 296 259 298 264
rect 368 259 370 264
rect 440 259 442 264
rect 504 259 506 264
rect 568 259 570 264
rect 632 259 634 264
rect 688 259 690 264
rect 744 259 746 264
rect 808 259 810 264
rect 880 259 882 264
rect 952 259 954 264
rect 1032 259 1034 264
rect 1112 259 1114 264
rect 1192 259 1194 264
rect 1264 259 1266 264
rect 1328 259 1330 264
rect 1392 259 1394 264
rect 1448 259 1450 264
rect 1496 259 1498 264
rect 1544 259 1546 264
rect 1592 259 1594 264
rect 1624 259 1626 264
rect 1664 259 1666 266
rect 111 258 115 259
rect 111 253 115 254
rect 135 258 139 259
rect 112 250 114 253
rect 135 252 139 254
rect 167 258 171 259
rect 167 253 171 254
rect 175 258 179 259
rect 175 252 179 254
rect 231 258 235 259
rect 231 253 235 254
rect 247 258 251 259
rect 247 252 251 254
rect 295 258 299 259
rect 295 253 299 254
rect 319 258 323 259
rect 319 252 323 254
rect 367 258 371 259
rect 367 253 371 254
rect 383 258 387 259
rect 383 252 387 254
rect 439 258 443 259
rect 439 253 443 254
rect 447 258 451 259
rect 447 252 451 254
rect 503 258 507 259
rect 503 253 507 254
rect 519 258 523 259
rect 519 252 523 254
rect 567 258 571 259
rect 567 253 571 254
rect 591 258 595 259
rect 591 252 595 254
rect 631 258 635 259
rect 631 253 635 254
rect 663 258 667 259
rect 663 252 667 254
rect 687 258 691 259
rect 687 253 691 254
rect 743 258 747 259
rect 743 252 747 254
rect 807 258 811 259
rect 807 253 811 254
rect 823 258 827 259
rect 823 252 827 254
rect 879 258 883 259
rect 879 253 883 254
rect 895 258 899 259
rect 895 252 899 254
rect 951 258 955 259
rect 951 253 955 254
rect 967 258 971 259
rect 967 252 971 254
rect 1031 258 1035 259
rect 1031 252 1035 254
rect 1087 258 1091 259
rect 1087 252 1091 254
rect 1111 258 1115 259
rect 1111 253 1115 254
rect 1143 258 1147 259
rect 1143 252 1147 254
rect 1191 258 1195 259
rect 1191 253 1195 254
rect 1199 258 1203 259
rect 1199 252 1203 254
rect 1255 258 1259 259
rect 1255 252 1259 254
rect 1263 258 1267 259
rect 1263 253 1267 254
rect 1311 258 1315 259
rect 1311 252 1315 254
rect 1327 258 1331 259
rect 1327 253 1331 254
rect 1367 258 1371 259
rect 1367 252 1371 254
rect 1391 258 1395 259
rect 1391 253 1395 254
rect 1415 258 1419 259
rect 1415 252 1419 254
rect 1447 258 1451 259
rect 1447 253 1451 254
rect 1463 258 1467 259
rect 1463 252 1467 254
rect 1495 258 1499 259
rect 1495 253 1499 254
rect 1519 258 1523 259
rect 1519 252 1523 254
rect 1543 258 1547 259
rect 1543 253 1547 254
rect 1575 258 1579 259
rect 1575 252 1579 254
rect 1591 258 1595 259
rect 1591 253 1595 254
rect 1623 258 1627 259
rect 1623 252 1627 254
rect 1663 258 1667 259
rect 1663 253 1667 254
rect 134 251 140 252
rect 110 249 116 250
rect 110 245 111 249
rect 115 245 116 249
rect 134 247 135 251
rect 139 247 140 251
rect 134 246 140 247
rect 174 251 180 252
rect 174 247 175 251
rect 179 247 180 251
rect 174 246 180 247
rect 246 251 252 252
rect 246 247 247 251
rect 251 247 252 251
rect 246 246 252 247
rect 318 251 324 252
rect 318 247 319 251
rect 323 247 324 251
rect 318 246 324 247
rect 382 251 388 252
rect 382 247 383 251
rect 387 247 388 251
rect 382 246 388 247
rect 446 251 452 252
rect 446 247 447 251
rect 451 247 452 251
rect 446 246 452 247
rect 518 251 524 252
rect 518 247 519 251
rect 523 247 524 251
rect 518 246 524 247
rect 590 251 596 252
rect 590 247 591 251
rect 595 247 596 251
rect 590 246 596 247
rect 662 251 668 252
rect 662 247 663 251
rect 667 247 668 251
rect 662 246 668 247
rect 742 251 748 252
rect 742 247 743 251
rect 747 247 748 251
rect 742 246 748 247
rect 822 251 828 252
rect 822 247 823 251
rect 827 247 828 251
rect 822 246 828 247
rect 894 251 900 252
rect 894 247 895 251
rect 899 247 900 251
rect 894 246 900 247
rect 966 251 972 252
rect 966 247 967 251
rect 971 247 972 251
rect 966 246 972 247
rect 1030 251 1036 252
rect 1030 247 1031 251
rect 1035 247 1036 251
rect 1030 246 1036 247
rect 1086 251 1092 252
rect 1086 247 1087 251
rect 1091 247 1092 251
rect 1086 246 1092 247
rect 1142 251 1148 252
rect 1142 247 1143 251
rect 1147 247 1148 251
rect 1142 246 1148 247
rect 1198 251 1204 252
rect 1198 247 1199 251
rect 1203 247 1204 251
rect 1198 246 1204 247
rect 1254 251 1260 252
rect 1254 247 1255 251
rect 1259 247 1260 251
rect 1254 246 1260 247
rect 1310 251 1316 252
rect 1310 247 1311 251
rect 1315 247 1316 251
rect 1310 246 1316 247
rect 1366 251 1372 252
rect 1366 247 1367 251
rect 1371 247 1372 251
rect 1366 246 1372 247
rect 1414 251 1420 252
rect 1414 247 1415 251
rect 1419 247 1420 251
rect 1414 246 1420 247
rect 1462 251 1468 252
rect 1462 247 1463 251
rect 1467 247 1468 251
rect 1462 246 1468 247
rect 1518 251 1524 252
rect 1518 247 1519 251
rect 1523 247 1524 251
rect 1518 246 1524 247
rect 1574 251 1580 252
rect 1574 247 1575 251
rect 1579 247 1580 251
rect 1574 246 1580 247
rect 1622 251 1628 252
rect 1622 247 1623 251
rect 1627 247 1628 251
rect 1664 250 1666 253
rect 1622 246 1628 247
rect 1662 249 1668 250
rect 110 244 116 245
rect 1662 245 1663 249
rect 1667 245 1668 249
rect 1662 244 1668 245
rect 134 234 140 235
rect 110 232 116 233
rect 110 228 111 232
rect 115 228 116 232
rect 134 230 135 234
rect 139 230 140 234
rect 134 229 140 230
rect 174 234 180 235
rect 174 230 175 234
rect 179 230 180 234
rect 174 229 180 230
rect 246 234 252 235
rect 246 230 247 234
rect 251 230 252 234
rect 246 229 252 230
rect 318 234 324 235
rect 318 230 319 234
rect 323 230 324 234
rect 318 229 324 230
rect 382 234 388 235
rect 382 230 383 234
rect 387 230 388 234
rect 382 229 388 230
rect 446 234 452 235
rect 446 230 447 234
rect 451 230 452 234
rect 446 229 452 230
rect 518 234 524 235
rect 518 230 519 234
rect 523 230 524 234
rect 518 229 524 230
rect 590 234 596 235
rect 590 230 591 234
rect 595 230 596 234
rect 590 229 596 230
rect 662 234 668 235
rect 662 230 663 234
rect 667 230 668 234
rect 662 229 668 230
rect 742 234 748 235
rect 742 230 743 234
rect 747 230 748 234
rect 742 229 748 230
rect 822 234 828 235
rect 822 230 823 234
rect 827 230 828 234
rect 822 229 828 230
rect 894 234 900 235
rect 894 230 895 234
rect 899 230 900 234
rect 894 229 900 230
rect 966 234 972 235
rect 966 230 967 234
rect 971 230 972 234
rect 966 229 972 230
rect 1030 234 1036 235
rect 1030 230 1031 234
rect 1035 230 1036 234
rect 1030 229 1036 230
rect 1086 234 1092 235
rect 1086 230 1087 234
rect 1091 230 1092 234
rect 1086 229 1092 230
rect 1142 234 1148 235
rect 1142 230 1143 234
rect 1147 230 1148 234
rect 1142 229 1148 230
rect 1198 234 1204 235
rect 1198 230 1199 234
rect 1203 230 1204 234
rect 1198 229 1204 230
rect 1254 234 1260 235
rect 1254 230 1255 234
rect 1259 230 1260 234
rect 1254 229 1260 230
rect 1310 234 1316 235
rect 1310 230 1311 234
rect 1315 230 1316 234
rect 1310 229 1316 230
rect 1366 234 1372 235
rect 1366 230 1367 234
rect 1371 230 1372 234
rect 1366 229 1372 230
rect 1414 234 1420 235
rect 1414 230 1415 234
rect 1419 230 1420 234
rect 1414 229 1420 230
rect 1462 234 1468 235
rect 1462 230 1463 234
rect 1467 230 1468 234
rect 1462 229 1468 230
rect 1518 234 1524 235
rect 1518 230 1519 234
rect 1523 230 1524 234
rect 1518 229 1524 230
rect 1574 234 1580 235
rect 1574 230 1575 234
rect 1579 230 1580 234
rect 1574 229 1580 230
rect 1622 234 1628 235
rect 1622 230 1623 234
rect 1627 230 1628 234
rect 1622 229 1628 230
rect 1662 232 1668 233
rect 110 227 116 228
rect 112 219 114 227
rect 136 219 138 229
rect 176 219 178 229
rect 248 219 250 229
rect 320 219 322 229
rect 384 219 386 229
rect 448 219 450 229
rect 520 219 522 229
rect 592 219 594 229
rect 664 219 666 229
rect 744 219 746 229
rect 824 219 826 229
rect 896 219 898 229
rect 968 219 970 229
rect 1032 219 1034 229
rect 1088 219 1090 229
rect 1144 219 1146 229
rect 1200 219 1202 229
rect 1256 219 1258 229
rect 1312 219 1314 229
rect 1368 219 1370 229
rect 1416 219 1418 229
rect 1464 219 1466 229
rect 1520 219 1522 229
rect 1576 219 1578 229
rect 1624 219 1626 229
rect 1662 228 1663 232
rect 1667 228 1668 232
rect 1662 227 1668 228
rect 1664 219 1666 227
rect 111 218 115 219
rect 111 213 115 214
rect 135 218 139 219
rect 135 213 139 214
rect 167 218 171 219
rect 167 213 171 214
rect 175 218 179 219
rect 175 213 179 214
rect 207 218 211 219
rect 207 213 211 214
rect 247 218 251 219
rect 247 213 251 214
rect 255 218 259 219
rect 255 213 259 214
rect 303 218 307 219
rect 303 213 307 214
rect 319 218 323 219
rect 319 213 323 214
rect 343 218 347 219
rect 343 213 347 214
rect 375 218 379 219
rect 375 213 379 214
rect 383 218 387 219
rect 383 213 387 214
rect 415 218 419 219
rect 415 213 419 214
rect 447 218 451 219
rect 447 213 451 214
rect 471 218 475 219
rect 471 213 475 214
rect 519 218 523 219
rect 519 213 523 214
rect 535 218 539 219
rect 535 213 539 214
rect 591 218 595 219
rect 591 213 595 214
rect 615 218 619 219
rect 615 213 619 214
rect 663 218 667 219
rect 663 213 667 214
rect 695 218 699 219
rect 695 213 699 214
rect 743 218 747 219
rect 743 213 747 214
rect 775 218 779 219
rect 775 213 779 214
rect 823 218 827 219
rect 823 213 827 214
rect 855 218 859 219
rect 855 213 859 214
rect 895 218 899 219
rect 895 213 899 214
rect 927 218 931 219
rect 927 213 931 214
rect 967 218 971 219
rect 967 213 971 214
rect 999 218 1003 219
rect 999 213 1003 214
rect 1031 218 1035 219
rect 1031 213 1035 214
rect 1071 218 1075 219
rect 1071 213 1075 214
rect 1087 218 1091 219
rect 1087 213 1091 214
rect 1143 218 1147 219
rect 1143 213 1147 214
rect 1199 218 1203 219
rect 1199 213 1203 214
rect 1215 218 1219 219
rect 1215 213 1219 214
rect 1255 218 1259 219
rect 1255 213 1259 214
rect 1287 218 1291 219
rect 1287 213 1291 214
rect 1311 218 1315 219
rect 1311 213 1315 214
rect 1351 218 1355 219
rect 1351 213 1355 214
rect 1367 218 1371 219
rect 1367 213 1371 214
rect 1415 218 1419 219
rect 1415 213 1419 214
rect 1463 218 1467 219
rect 1463 213 1467 214
rect 1471 218 1475 219
rect 1471 213 1475 214
rect 1519 218 1523 219
rect 1519 213 1523 214
rect 1527 218 1531 219
rect 1527 213 1531 214
rect 1575 218 1579 219
rect 1575 213 1579 214
rect 1583 218 1587 219
rect 1583 213 1587 214
rect 1623 218 1627 219
rect 1623 213 1627 214
rect 1663 218 1667 219
rect 1663 213 1667 214
rect 112 205 114 213
rect 110 204 116 205
rect 110 200 111 204
rect 115 200 116 204
rect 136 203 138 213
rect 168 203 170 213
rect 208 203 210 213
rect 256 203 258 213
rect 304 203 306 213
rect 344 203 346 213
rect 376 203 378 213
rect 416 203 418 213
rect 472 203 474 213
rect 536 203 538 213
rect 616 203 618 213
rect 696 203 698 213
rect 776 203 778 213
rect 856 203 858 213
rect 928 203 930 213
rect 1000 203 1002 213
rect 1072 203 1074 213
rect 1144 203 1146 213
rect 1216 203 1218 213
rect 1288 203 1290 213
rect 1352 203 1354 213
rect 1416 203 1418 213
rect 1472 203 1474 213
rect 1528 203 1530 213
rect 1584 203 1586 213
rect 1624 203 1626 213
rect 1664 205 1666 213
rect 1662 204 1668 205
rect 110 199 116 200
rect 134 202 140 203
rect 134 198 135 202
rect 139 198 140 202
rect 134 197 140 198
rect 166 202 172 203
rect 166 198 167 202
rect 171 198 172 202
rect 166 197 172 198
rect 206 202 212 203
rect 206 198 207 202
rect 211 198 212 202
rect 206 197 212 198
rect 254 202 260 203
rect 254 198 255 202
rect 259 198 260 202
rect 254 197 260 198
rect 302 202 308 203
rect 302 198 303 202
rect 307 198 308 202
rect 302 197 308 198
rect 342 202 348 203
rect 342 198 343 202
rect 347 198 348 202
rect 342 197 348 198
rect 374 202 380 203
rect 374 198 375 202
rect 379 198 380 202
rect 374 197 380 198
rect 414 202 420 203
rect 414 198 415 202
rect 419 198 420 202
rect 414 197 420 198
rect 470 202 476 203
rect 470 198 471 202
rect 475 198 476 202
rect 470 197 476 198
rect 534 202 540 203
rect 534 198 535 202
rect 539 198 540 202
rect 534 197 540 198
rect 614 202 620 203
rect 614 198 615 202
rect 619 198 620 202
rect 614 197 620 198
rect 694 202 700 203
rect 694 198 695 202
rect 699 198 700 202
rect 694 197 700 198
rect 774 202 780 203
rect 774 198 775 202
rect 779 198 780 202
rect 774 197 780 198
rect 854 202 860 203
rect 854 198 855 202
rect 859 198 860 202
rect 854 197 860 198
rect 926 202 932 203
rect 926 198 927 202
rect 931 198 932 202
rect 926 197 932 198
rect 998 202 1004 203
rect 998 198 999 202
rect 1003 198 1004 202
rect 998 197 1004 198
rect 1070 202 1076 203
rect 1070 198 1071 202
rect 1075 198 1076 202
rect 1070 197 1076 198
rect 1142 202 1148 203
rect 1142 198 1143 202
rect 1147 198 1148 202
rect 1142 197 1148 198
rect 1214 202 1220 203
rect 1214 198 1215 202
rect 1219 198 1220 202
rect 1214 197 1220 198
rect 1286 202 1292 203
rect 1286 198 1287 202
rect 1291 198 1292 202
rect 1286 197 1292 198
rect 1350 202 1356 203
rect 1350 198 1351 202
rect 1355 198 1356 202
rect 1350 197 1356 198
rect 1414 202 1420 203
rect 1414 198 1415 202
rect 1419 198 1420 202
rect 1414 197 1420 198
rect 1470 202 1476 203
rect 1470 198 1471 202
rect 1475 198 1476 202
rect 1470 197 1476 198
rect 1526 202 1532 203
rect 1526 198 1527 202
rect 1531 198 1532 202
rect 1526 197 1532 198
rect 1582 202 1588 203
rect 1582 198 1583 202
rect 1587 198 1588 202
rect 1582 197 1588 198
rect 1622 202 1628 203
rect 1622 198 1623 202
rect 1627 198 1628 202
rect 1662 200 1663 204
rect 1667 200 1668 204
rect 1662 199 1668 200
rect 1622 197 1628 198
rect 110 187 116 188
rect 110 183 111 187
rect 115 183 116 187
rect 1662 187 1668 188
rect 110 182 116 183
rect 134 185 140 186
rect 112 179 114 182
rect 134 181 135 185
rect 139 181 140 185
rect 134 180 140 181
rect 166 185 172 186
rect 166 181 167 185
rect 171 181 172 185
rect 166 180 172 181
rect 206 185 212 186
rect 206 181 207 185
rect 211 181 212 185
rect 206 180 212 181
rect 254 185 260 186
rect 254 181 255 185
rect 259 181 260 185
rect 254 180 260 181
rect 302 185 308 186
rect 302 181 303 185
rect 307 181 308 185
rect 302 180 308 181
rect 342 185 348 186
rect 342 181 343 185
rect 347 181 348 185
rect 342 180 348 181
rect 374 185 380 186
rect 374 181 375 185
rect 379 181 380 185
rect 374 180 380 181
rect 414 185 420 186
rect 414 181 415 185
rect 419 181 420 185
rect 414 180 420 181
rect 470 185 476 186
rect 470 181 471 185
rect 475 181 476 185
rect 470 180 476 181
rect 534 185 540 186
rect 534 181 535 185
rect 539 181 540 185
rect 534 180 540 181
rect 614 185 620 186
rect 614 181 615 185
rect 619 181 620 185
rect 614 180 620 181
rect 694 185 700 186
rect 694 181 695 185
rect 699 181 700 185
rect 694 180 700 181
rect 774 185 780 186
rect 774 181 775 185
rect 779 181 780 185
rect 774 180 780 181
rect 854 185 860 186
rect 854 181 855 185
rect 859 181 860 185
rect 854 180 860 181
rect 926 185 932 186
rect 926 181 927 185
rect 931 181 932 185
rect 926 180 932 181
rect 998 185 1004 186
rect 998 181 999 185
rect 1003 181 1004 185
rect 998 180 1004 181
rect 1070 185 1076 186
rect 1070 181 1071 185
rect 1075 181 1076 185
rect 1070 180 1076 181
rect 1142 185 1148 186
rect 1142 181 1143 185
rect 1147 181 1148 185
rect 1142 180 1148 181
rect 1214 185 1220 186
rect 1214 181 1215 185
rect 1219 181 1220 185
rect 1214 180 1220 181
rect 1286 185 1292 186
rect 1286 181 1287 185
rect 1291 181 1292 185
rect 1286 180 1292 181
rect 1350 185 1356 186
rect 1350 181 1351 185
rect 1355 181 1356 185
rect 1350 180 1356 181
rect 1414 185 1420 186
rect 1414 181 1415 185
rect 1419 181 1420 185
rect 1414 180 1420 181
rect 1470 185 1476 186
rect 1470 181 1471 185
rect 1475 181 1476 185
rect 1470 180 1476 181
rect 1526 185 1532 186
rect 1526 181 1527 185
rect 1531 181 1532 185
rect 1526 180 1532 181
rect 1582 185 1588 186
rect 1582 181 1583 185
rect 1587 181 1588 185
rect 1582 180 1588 181
rect 1622 185 1628 186
rect 1622 181 1623 185
rect 1627 181 1628 185
rect 1662 183 1663 187
rect 1667 183 1668 187
rect 1662 182 1668 183
rect 1622 180 1628 181
rect 111 178 115 179
rect 111 173 115 174
rect 135 178 139 180
rect 112 170 114 173
rect 135 172 139 174
rect 167 178 171 180
rect 167 173 171 174
rect 175 178 179 179
rect 175 172 179 174
rect 207 178 211 180
rect 207 173 211 174
rect 231 178 235 179
rect 231 172 235 174
rect 255 178 259 180
rect 255 173 259 174
rect 287 178 291 179
rect 287 172 291 174
rect 303 178 307 180
rect 303 173 307 174
rect 343 178 347 180
rect 343 172 347 174
rect 375 178 379 180
rect 375 173 379 174
rect 399 178 403 179
rect 399 172 403 174
rect 415 178 419 180
rect 415 173 419 174
rect 455 178 459 179
rect 455 172 459 174
rect 471 178 475 180
rect 471 173 475 174
rect 511 178 515 179
rect 511 172 515 174
rect 535 178 539 180
rect 535 173 539 174
rect 575 178 579 179
rect 575 172 579 174
rect 615 178 619 180
rect 615 173 619 174
rect 639 178 643 179
rect 639 172 643 174
rect 695 178 699 180
rect 695 173 699 174
rect 703 178 707 179
rect 703 172 707 174
rect 767 178 771 179
rect 767 172 771 174
rect 775 178 779 180
rect 775 173 779 174
rect 831 178 835 179
rect 831 172 835 174
rect 855 178 859 180
rect 855 173 859 174
rect 895 178 899 179
rect 895 172 899 174
rect 927 178 931 180
rect 927 173 931 174
rect 951 178 955 179
rect 951 172 955 174
rect 999 178 1003 180
rect 999 173 1003 174
rect 1015 178 1019 179
rect 1015 172 1019 174
rect 1071 178 1075 180
rect 1071 173 1075 174
rect 1079 178 1083 179
rect 1079 172 1083 174
rect 1143 178 1147 180
rect 1143 172 1147 174
rect 1207 178 1211 179
rect 1207 172 1211 174
rect 1215 178 1219 180
rect 1215 173 1219 174
rect 1279 178 1283 179
rect 1279 172 1283 174
rect 1287 178 1291 180
rect 1287 173 1291 174
rect 1351 178 1355 180
rect 1351 172 1355 174
rect 1415 178 1419 180
rect 1415 173 1419 174
rect 1423 178 1427 179
rect 1423 172 1427 174
rect 1471 178 1475 180
rect 1471 173 1475 174
rect 1495 178 1499 179
rect 1495 172 1499 174
rect 1527 178 1531 180
rect 1527 173 1531 174
rect 1567 178 1571 179
rect 1567 172 1571 174
rect 1583 178 1587 180
rect 1583 173 1587 174
rect 1623 178 1627 180
rect 1664 179 1666 182
rect 1623 172 1627 174
rect 1663 178 1667 179
rect 1663 173 1667 174
rect 134 171 140 172
rect 110 169 116 170
rect 110 165 111 169
rect 115 165 116 169
rect 134 167 135 171
rect 139 167 140 171
rect 134 166 140 167
rect 174 171 180 172
rect 174 167 175 171
rect 179 167 180 171
rect 174 166 180 167
rect 230 171 236 172
rect 230 167 231 171
rect 235 167 236 171
rect 230 166 236 167
rect 286 171 292 172
rect 286 167 287 171
rect 291 167 292 171
rect 286 166 292 167
rect 342 171 348 172
rect 342 167 343 171
rect 347 167 348 171
rect 342 166 348 167
rect 398 171 404 172
rect 398 167 399 171
rect 403 167 404 171
rect 398 166 404 167
rect 454 171 460 172
rect 454 167 455 171
rect 459 167 460 171
rect 454 166 460 167
rect 510 171 516 172
rect 510 167 511 171
rect 515 167 516 171
rect 510 166 516 167
rect 574 171 580 172
rect 574 167 575 171
rect 579 167 580 171
rect 574 166 580 167
rect 638 171 644 172
rect 638 167 639 171
rect 643 167 644 171
rect 638 166 644 167
rect 702 171 708 172
rect 702 167 703 171
rect 707 167 708 171
rect 702 166 708 167
rect 766 171 772 172
rect 766 167 767 171
rect 771 167 772 171
rect 766 166 772 167
rect 830 171 836 172
rect 830 167 831 171
rect 835 167 836 171
rect 830 166 836 167
rect 894 171 900 172
rect 894 167 895 171
rect 899 167 900 171
rect 894 166 900 167
rect 950 171 956 172
rect 950 167 951 171
rect 955 167 956 171
rect 950 166 956 167
rect 1014 171 1020 172
rect 1014 167 1015 171
rect 1019 167 1020 171
rect 1014 166 1020 167
rect 1078 171 1084 172
rect 1078 167 1079 171
rect 1083 167 1084 171
rect 1078 166 1084 167
rect 1142 171 1148 172
rect 1142 167 1143 171
rect 1147 167 1148 171
rect 1142 166 1148 167
rect 1206 171 1212 172
rect 1206 167 1207 171
rect 1211 167 1212 171
rect 1206 166 1212 167
rect 1278 171 1284 172
rect 1278 167 1279 171
rect 1283 167 1284 171
rect 1278 166 1284 167
rect 1350 171 1356 172
rect 1350 167 1351 171
rect 1355 167 1356 171
rect 1350 166 1356 167
rect 1422 171 1428 172
rect 1422 167 1423 171
rect 1427 167 1428 171
rect 1422 166 1428 167
rect 1494 171 1500 172
rect 1494 167 1495 171
rect 1499 167 1500 171
rect 1494 166 1500 167
rect 1566 171 1572 172
rect 1566 167 1567 171
rect 1571 167 1572 171
rect 1566 166 1572 167
rect 1622 171 1628 172
rect 1622 167 1623 171
rect 1627 167 1628 171
rect 1664 170 1666 173
rect 1622 166 1628 167
rect 1662 169 1668 170
rect 110 164 116 165
rect 1662 165 1663 169
rect 1667 165 1668 169
rect 1662 164 1668 165
rect 134 154 140 155
rect 110 152 116 153
rect 110 148 111 152
rect 115 148 116 152
rect 134 150 135 154
rect 139 150 140 154
rect 134 149 140 150
rect 174 154 180 155
rect 174 150 175 154
rect 179 150 180 154
rect 174 149 180 150
rect 230 154 236 155
rect 230 150 231 154
rect 235 150 236 154
rect 230 149 236 150
rect 286 154 292 155
rect 286 150 287 154
rect 291 150 292 154
rect 286 149 292 150
rect 342 154 348 155
rect 342 150 343 154
rect 347 150 348 154
rect 342 149 348 150
rect 398 154 404 155
rect 398 150 399 154
rect 403 150 404 154
rect 398 149 404 150
rect 454 154 460 155
rect 454 150 455 154
rect 459 150 460 154
rect 454 149 460 150
rect 510 154 516 155
rect 510 150 511 154
rect 515 150 516 154
rect 510 149 516 150
rect 574 154 580 155
rect 574 150 575 154
rect 579 150 580 154
rect 574 149 580 150
rect 638 154 644 155
rect 638 150 639 154
rect 643 150 644 154
rect 638 149 644 150
rect 702 154 708 155
rect 702 150 703 154
rect 707 150 708 154
rect 702 149 708 150
rect 766 154 772 155
rect 766 150 767 154
rect 771 150 772 154
rect 766 149 772 150
rect 830 154 836 155
rect 830 150 831 154
rect 835 150 836 154
rect 830 149 836 150
rect 894 154 900 155
rect 894 150 895 154
rect 899 150 900 154
rect 894 149 900 150
rect 950 154 956 155
rect 950 150 951 154
rect 955 150 956 154
rect 950 149 956 150
rect 1014 154 1020 155
rect 1014 150 1015 154
rect 1019 150 1020 154
rect 1014 149 1020 150
rect 1078 154 1084 155
rect 1078 150 1079 154
rect 1083 150 1084 154
rect 1078 149 1084 150
rect 1142 154 1148 155
rect 1142 150 1143 154
rect 1147 150 1148 154
rect 1142 149 1148 150
rect 1206 154 1212 155
rect 1206 150 1207 154
rect 1211 150 1212 154
rect 1206 149 1212 150
rect 1278 154 1284 155
rect 1278 150 1279 154
rect 1283 150 1284 154
rect 1278 149 1284 150
rect 1350 154 1356 155
rect 1350 150 1351 154
rect 1355 150 1356 154
rect 1350 149 1356 150
rect 1422 154 1428 155
rect 1422 150 1423 154
rect 1427 150 1428 154
rect 1422 149 1428 150
rect 1494 154 1500 155
rect 1494 150 1495 154
rect 1499 150 1500 154
rect 1494 149 1500 150
rect 1566 154 1572 155
rect 1566 150 1567 154
rect 1571 150 1572 154
rect 1566 149 1572 150
rect 1622 154 1628 155
rect 1622 150 1623 154
rect 1627 150 1628 154
rect 1622 149 1628 150
rect 1662 152 1668 153
rect 110 147 116 148
rect 112 123 114 147
rect 136 123 138 149
rect 176 123 178 149
rect 232 123 234 149
rect 288 123 290 149
rect 344 123 346 149
rect 400 123 402 149
rect 456 123 458 149
rect 512 123 514 149
rect 576 123 578 149
rect 640 123 642 149
rect 704 123 706 149
rect 768 123 770 149
rect 832 123 834 149
rect 896 123 898 149
rect 952 123 954 149
rect 1016 123 1018 149
rect 1080 123 1082 149
rect 1144 123 1146 149
rect 1208 123 1210 149
rect 1280 123 1282 149
rect 1352 123 1354 149
rect 1424 123 1426 149
rect 1496 123 1498 149
rect 1568 123 1570 149
rect 1624 123 1626 149
rect 1662 148 1663 152
rect 1667 148 1668 152
rect 1662 147 1668 148
rect 1664 123 1666 147
rect 111 122 115 123
rect 111 117 115 118
rect 135 122 139 123
rect 135 117 139 118
rect 167 122 171 123
rect 167 117 171 118
rect 175 122 179 123
rect 175 117 179 118
rect 199 122 203 123
rect 199 117 203 118
rect 231 122 235 123
rect 231 117 235 118
rect 263 122 267 123
rect 263 117 267 118
rect 287 122 291 123
rect 287 117 291 118
rect 295 122 299 123
rect 295 117 299 118
rect 327 122 331 123
rect 327 117 331 118
rect 343 122 347 123
rect 343 117 347 118
rect 359 122 363 123
rect 359 117 363 118
rect 391 122 395 123
rect 391 117 395 118
rect 399 122 403 123
rect 399 117 403 118
rect 423 122 427 123
rect 423 117 427 118
rect 455 122 459 123
rect 455 117 459 118
rect 463 122 467 123
rect 463 117 467 118
rect 503 122 507 123
rect 503 117 507 118
rect 511 122 515 123
rect 511 117 515 118
rect 543 122 547 123
rect 543 117 547 118
rect 575 122 579 123
rect 575 117 579 118
rect 607 122 611 123
rect 607 117 611 118
rect 639 122 643 123
rect 639 117 643 118
rect 671 122 675 123
rect 671 117 675 118
rect 703 122 707 123
rect 703 117 707 118
rect 735 122 739 123
rect 735 117 739 118
rect 767 122 771 123
rect 767 117 771 118
rect 799 122 803 123
rect 799 117 803 118
rect 831 122 835 123
rect 831 117 835 118
rect 863 122 867 123
rect 863 117 867 118
rect 895 122 899 123
rect 895 117 899 118
rect 935 122 939 123
rect 935 117 939 118
rect 951 122 955 123
rect 951 117 955 118
rect 975 122 979 123
rect 975 117 979 118
rect 1015 122 1019 123
rect 1015 117 1019 118
rect 1063 122 1067 123
rect 1063 117 1067 118
rect 1079 122 1083 123
rect 1079 117 1083 118
rect 1103 122 1107 123
rect 1103 117 1107 118
rect 1143 122 1147 123
rect 1143 117 1147 118
rect 1183 122 1187 123
rect 1183 117 1187 118
rect 1207 122 1211 123
rect 1207 117 1211 118
rect 1223 122 1227 123
rect 1223 117 1227 118
rect 1263 122 1267 123
rect 1263 117 1267 118
rect 1279 122 1283 123
rect 1279 117 1283 118
rect 1295 122 1299 123
rect 1295 117 1299 118
rect 1335 122 1339 123
rect 1335 117 1339 118
rect 1351 122 1355 123
rect 1351 117 1355 118
rect 1375 122 1379 123
rect 1375 117 1379 118
rect 1415 122 1419 123
rect 1415 117 1419 118
rect 1423 122 1427 123
rect 1423 117 1427 118
rect 1455 122 1459 123
rect 1455 117 1459 118
rect 1495 122 1499 123
rect 1495 117 1499 118
rect 1503 122 1507 123
rect 1503 117 1507 118
rect 1551 122 1555 123
rect 1551 117 1555 118
rect 1567 122 1571 123
rect 1567 117 1571 118
rect 1591 122 1595 123
rect 1591 117 1595 118
rect 1623 122 1627 123
rect 1623 117 1627 118
rect 1663 122 1667 123
rect 1663 117 1667 118
rect 112 109 114 117
rect 110 108 116 109
rect 110 104 111 108
rect 115 104 116 108
rect 136 107 138 117
rect 168 107 170 117
rect 200 107 202 117
rect 232 107 234 117
rect 264 107 266 117
rect 296 107 298 117
rect 328 107 330 117
rect 360 107 362 117
rect 392 107 394 117
rect 424 107 426 117
rect 464 107 466 117
rect 504 107 506 117
rect 544 107 546 117
rect 576 107 578 117
rect 608 107 610 117
rect 640 107 642 117
rect 672 107 674 117
rect 704 107 706 117
rect 736 107 738 117
rect 768 107 770 117
rect 800 107 802 117
rect 832 107 834 117
rect 864 107 866 117
rect 896 107 898 117
rect 936 107 938 117
rect 976 107 978 117
rect 1016 107 1018 117
rect 1064 107 1066 117
rect 1104 107 1106 117
rect 1144 107 1146 117
rect 1184 107 1186 117
rect 1224 107 1226 117
rect 1264 107 1266 117
rect 1296 107 1298 117
rect 1336 107 1338 117
rect 1376 107 1378 117
rect 1416 107 1418 117
rect 1456 107 1458 117
rect 1504 107 1506 117
rect 1552 107 1554 117
rect 1592 107 1594 117
rect 1624 107 1626 117
rect 1664 109 1666 117
rect 1662 108 1668 109
rect 110 103 116 104
rect 134 106 140 107
rect 134 102 135 106
rect 139 102 140 106
rect 134 101 140 102
rect 166 106 172 107
rect 166 102 167 106
rect 171 102 172 106
rect 166 101 172 102
rect 198 106 204 107
rect 198 102 199 106
rect 203 102 204 106
rect 198 101 204 102
rect 230 106 236 107
rect 230 102 231 106
rect 235 102 236 106
rect 230 101 236 102
rect 262 106 268 107
rect 262 102 263 106
rect 267 102 268 106
rect 262 101 268 102
rect 294 106 300 107
rect 294 102 295 106
rect 299 102 300 106
rect 294 101 300 102
rect 326 106 332 107
rect 326 102 327 106
rect 331 102 332 106
rect 326 101 332 102
rect 358 106 364 107
rect 358 102 359 106
rect 363 102 364 106
rect 358 101 364 102
rect 390 106 396 107
rect 390 102 391 106
rect 395 102 396 106
rect 390 101 396 102
rect 422 106 428 107
rect 422 102 423 106
rect 427 102 428 106
rect 422 101 428 102
rect 462 106 468 107
rect 462 102 463 106
rect 467 102 468 106
rect 462 101 468 102
rect 502 106 508 107
rect 502 102 503 106
rect 507 102 508 106
rect 502 101 508 102
rect 542 106 548 107
rect 542 102 543 106
rect 547 102 548 106
rect 542 101 548 102
rect 574 106 580 107
rect 574 102 575 106
rect 579 102 580 106
rect 574 101 580 102
rect 606 106 612 107
rect 606 102 607 106
rect 611 102 612 106
rect 606 101 612 102
rect 638 106 644 107
rect 638 102 639 106
rect 643 102 644 106
rect 638 101 644 102
rect 670 106 676 107
rect 670 102 671 106
rect 675 102 676 106
rect 670 101 676 102
rect 702 106 708 107
rect 702 102 703 106
rect 707 102 708 106
rect 702 101 708 102
rect 734 106 740 107
rect 734 102 735 106
rect 739 102 740 106
rect 734 101 740 102
rect 766 106 772 107
rect 766 102 767 106
rect 771 102 772 106
rect 766 101 772 102
rect 798 106 804 107
rect 798 102 799 106
rect 803 102 804 106
rect 798 101 804 102
rect 830 106 836 107
rect 830 102 831 106
rect 835 102 836 106
rect 830 101 836 102
rect 862 106 868 107
rect 862 102 863 106
rect 867 102 868 106
rect 862 101 868 102
rect 894 106 900 107
rect 894 102 895 106
rect 899 102 900 106
rect 894 101 900 102
rect 934 106 940 107
rect 934 102 935 106
rect 939 102 940 106
rect 934 101 940 102
rect 974 106 980 107
rect 974 102 975 106
rect 979 102 980 106
rect 974 101 980 102
rect 1014 106 1020 107
rect 1014 102 1015 106
rect 1019 102 1020 106
rect 1014 101 1020 102
rect 1062 106 1068 107
rect 1062 102 1063 106
rect 1067 102 1068 106
rect 1062 101 1068 102
rect 1102 106 1108 107
rect 1102 102 1103 106
rect 1107 102 1108 106
rect 1102 101 1108 102
rect 1142 106 1148 107
rect 1142 102 1143 106
rect 1147 102 1148 106
rect 1142 101 1148 102
rect 1182 106 1188 107
rect 1182 102 1183 106
rect 1187 102 1188 106
rect 1182 101 1188 102
rect 1222 106 1228 107
rect 1222 102 1223 106
rect 1227 102 1228 106
rect 1222 101 1228 102
rect 1262 106 1268 107
rect 1262 102 1263 106
rect 1267 102 1268 106
rect 1262 101 1268 102
rect 1294 106 1300 107
rect 1294 102 1295 106
rect 1299 102 1300 106
rect 1294 101 1300 102
rect 1334 106 1340 107
rect 1334 102 1335 106
rect 1339 102 1340 106
rect 1334 101 1340 102
rect 1374 106 1380 107
rect 1374 102 1375 106
rect 1379 102 1380 106
rect 1374 101 1380 102
rect 1414 106 1420 107
rect 1414 102 1415 106
rect 1419 102 1420 106
rect 1414 101 1420 102
rect 1454 106 1460 107
rect 1454 102 1455 106
rect 1459 102 1460 106
rect 1454 101 1460 102
rect 1502 106 1508 107
rect 1502 102 1503 106
rect 1507 102 1508 106
rect 1502 101 1508 102
rect 1550 106 1556 107
rect 1550 102 1551 106
rect 1555 102 1556 106
rect 1550 101 1556 102
rect 1590 106 1596 107
rect 1590 102 1591 106
rect 1595 102 1596 106
rect 1590 101 1596 102
rect 1622 106 1628 107
rect 1622 102 1623 106
rect 1627 102 1628 106
rect 1662 104 1663 108
rect 1667 104 1668 108
rect 1662 103 1668 104
rect 1622 101 1628 102
rect 110 91 116 92
rect 110 87 111 91
rect 115 87 116 91
rect 1662 91 1668 92
rect 110 86 116 87
rect 134 89 140 90
rect 112 83 114 86
rect 134 85 135 89
rect 139 85 140 89
rect 134 84 140 85
rect 166 89 172 90
rect 166 85 167 89
rect 171 85 172 89
rect 166 84 172 85
rect 198 89 204 90
rect 198 85 199 89
rect 203 85 204 89
rect 198 84 204 85
rect 230 89 236 90
rect 230 85 231 89
rect 235 85 236 89
rect 230 84 236 85
rect 262 89 268 90
rect 262 85 263 89
rect 267 85 268 89
rect 262 84 268 85
rect 294 89 300 90
rect 294 85 295 89
rect 299 85 300 89
rect 294 84 300 85
rect 326 89 332 90
rect 326 85 327 89
rect 331 85 332 89
rect 326 84 332 85
rect 358 89 364 90
rect 358 85 359 89
rect 363 85 364 89
rect 358 84 364 85
rect 390 89 396 90
rect 390 85 391 89
rect 395 85 396 89
rect 390 84 396 85
rect 422 89 428 90
rect 422 85 423 89
rect 427 85 428 89
rect 422 84 428 85
rect 462 89 468 90
rect 462 85 463 89
rect 467 85 468 89
rect 462 84 468 85
rect 502 89 508 90
rect 502 85 503 89
rect 507 85 508 89
rect 502 84 508 85
rect 542 89 548 90
rect 542 85 543 89
rect 547 85 548 89
rect 542 84 548 85
rect 574 89 580 90
rect 574 85 575 89
rect 579 85 580 89
rect 574 84 580 85
rect 606 89 612 90
rect 606 85 607 89
rect 611 85 612 89
rect 606 84 612 85
rect 638 89 644 90
rect 638 85 639 89
rect 643 85 644 89
rect 638 84 644 85
rect 670 89 676 90
rect 670 85 671 89
rect 675 85 676 89
rect 670 84 676 85
rect 702 89 708 90
rect 702 85 703 89
rect 707 85 708 89
rect 702 84 708 85
rect 734 89 740 90
rect 734 85 735 89
rect 739 85 740 89
rect 734 84 740 85
rect 766 89 772 90
rect 766 85 767 89
rect 771 85 772 89
rect 766 84 772 85
rect 798 89 804 90
rect 798 85 799 89
rect 803 85 804 89
rect 798 84 804 85
rect 830 89 836 90
rect 830 85 831 89
rect 835 85 836 89
rect 830 84 836 85
rect 862 89 868 90
rect 862 85 863 89
rect 867 85 868 89
rect 862 84 868 85
rect 894 89 900 90
rect 894 85 895 89
rect 899 85 900 89
rect 894 84 900 85
rect 934 89 940 90
rect 934 85 935 89
rect 939 85 940 89
rect 934 84 940 85
rect 974 89 980 90
rect 974 85 975 89
rect 979 85 980 89
rect 974 84 980 85
rect 1014 89 1020 90
rect 1014 85 1015 89
rect 1019 85 1020 89
rect 1014 84 1020 85
rect 1062 89 1068 90
rect 1062 85 1063 89
rect 1067 85 1068 89
rect 1062 84 1068 85
rect 1102 89 1108 90
rect 1102 85 1103 89
rect 1107 85 1108 89
rect 1102 84 1108 85
rect 1142 89 1148 90
rect 1142 85 1143 89
rect 1147 85 1148 89
rect 1142 84 1148 85
rect 1182 89 1188 90
rect 1182 85 1183 89
rect 1187 85 1188 89
rect 1182 84 1188 85
rect 1222 89 1228 90
rect 1222 85 1223 89
rect 1227 85 1228 89
rect 1222 84 1228 85
rect 1262 89 1268 90
rect 1262 85 1263 89
rect 1267 85 1268 89
rect 1262 84 1268 85
rect 1294 89 1300 90
rect 1294 85 1295 89
rect 1299 85 1300 89
rect 1294 84 1300 85
rect 1334 89 1340 90
rect 1334 85 1335 89
rect 1339 85 1340 89
rect 1334 84 1340 85
rect 1374 89 1380 90
rect 1374 85 1375 89
rect 1379 85 1380 89
rect 1374 84 1380 85
rect 1414 89 1420 90
rect 1414 85 1415 89
rect 1419 85 1420 89
rect 1414 84 1420 85
rect 1454 89 1460 90
rect 1454 85 1455 89
rect 1459 85 1460 89
rect 1454 84 1460 85
rect 1502 89 1508 90
rect 1502 85 1503 89
rect 1507 85 1508 89
rect 1502 84 1508 85
rect 1550 89 1556 90
rect 1550 85 1551 89
rect 1555 85 1556 89
rect 1550 84 1556 85
rect 1590 89 1596 90
rect 1590 85 1591 89
rect 1595 85 1596 89
rect 1590 84 1596 85
rect 1622 89 1628 90
rect 1622 85 1623 89
rect 1627 85 1628 89
rect 1662 87 1663 91
rect 1667 87 1668 91
rect 1662 86 1668 87
rect 1622 84 1628 85
rect 111 82 115 83
rect 111 77 115 78
rect 135 82 139 84
rect 135 77 139 78
rect 167 82 171 84
rect 167 77 171 78
rect 199 82 203 84
rect 199 77 203 78
rect 231 82 235 84
rect 231 77 235 78
rect 263 82 267 84
rect 263 77 267 78
rect 295 82 299 84
rect 295 77 299 78
rect 327 82 331 84
rect 327 77 331 78
rect 359 82 363 84
rect 359 77 363 78
rect 391 82 395 84
rect 391 77 395 78
rect 423 82 427 84
rect 423 77 427 78
rect 463 82 467 84
rect 463 77 467 78
rect 503 82 507 84
rect 503 77 507 78
rect 543 82 547 84
rect 543 77 547 78
rect 575 82 579 84
rect 575 77 579 78
rect 607 82 611 84
rect 607 77 611 78
rect 639 82 643 84
rect 639 77 643 78
rect 671 82 675 84
rect 671 77 675 78
rect 703 82 707 84
rect 703 77 707 78
rect 735 82 739 84
rect 735 77 739 78
rect 767 82 771 84
rect 767 77 771 78
rect 799 82 803 84
rect 799 77 803 78
rect 831 82 835 84
rect 831 77 835 78
rect 863 82 867 84
rect 863 77 867 78
rect 895 82 899 84
rect 895 77 899 78
rect 935 82 939 84
rect 935 77 939 78
rect 975 82 979 84
rect 975 77 979 78
rect 1015 82 1019 84
rect 1015 77 1019 78
rect 1063 82 1067 84
rect 1063 77 1067 78
rect 1103 82 1107 84
rect 1103 77 1107 78
rect 1143 82 1147 84
rect 1143 77 1147 78
rect 1183 82 1187 84
rect 1183 77 1187 78
rect 1223 82 1227 84
rect 1223 77 1227 78
rect 1263 82 1267 84
rect 1263 77 1267 78
rect 1295 82 1299 84
rect 1295 77 1299 78
rect 1335 82 1339 84
rect 1335 77 1339 78
rect 1375 82 1379 84
rect 1375 77 1379 78
rect 1415 82 1419 84
rect 1415 77 1419 78
rect 1455 82 1459 84
rect 1455 77 1459 78
rect 1503 82 1507 84
rect 1503 77 1507 78
rect 1551 82 1555 84
rect 1551 77 1555 78
rect 1591 82 1595 84
rect 1591 77 1595 78
rect 1623 82 1627 84
rect 1664 83 1666 86
rect 1623 77 1627 78
rect 1663 82 1667 83
rect 1663 77 1667 78
<< m4c >>
rect 111 1714 115 1718
rect 255 1714 259 1718
rect 287 1714 291 1718
rect 319 1714 323 1718
rect 359 1714 363 1718
rect 407 1714 411 1718
rect 455 1714 459 1718
rect 503 1714 507 1718
rect 551 1714 555 1718
rect 607 1714 611 1718
rect 663 1714 667 1718
rect 727 1714 731 1718
rect 783 1714 787 1718
rect 839 1714 843 1718
rect 895 1714 899 1718
rect 951 1714 955 1718
rect 1007 1714 1011 1718
rect 1063 1714 1067 1718
rect 1119 1714 1123 1718
rect 1175 1714 1179 1718
rect 1231 1714 1235 1718
rect 1287 1714 1291 1718
rect 1335 1714 1339 1718
rect 1375 1714 1379 1718
rect 1423 1714 1427 1718
rect 1471 1714 1475 1718
rect 1519 1714 1523 1718
rect 1663 1714 1667 1718
rect 111 1674 115 1678
rect 135 1674 139 1678
rect 167 1674 171 1678
rect 215 1674 219 1678
rect 255 1674 259 1678
rect 279 1674 283 1678
rect 287 1674 291 1678
rect 319 1674 323 1678
rect 343 1674 347 1678
rect 359 1674 363 1678
rect 407 1674 411 1678
rect 415 1674 419 1678
rect 455 1674 459 1678
rect 487 1674 491 1678
rect 503 1674 507 1678
rect 551 1674 555 1678
rect 559 1674 563 1678
rect 607 1674 611 1678
rect 631 1674 635 1678
rect 663 1674 667 1678
rect 711 1674 715 1678
rect 727 1674 731 1678
rect 783 1674 787 1678
rect 791 1674 795 1678
rect 839 1674 843 1678
rect 871 1674 875 1678
rect 895 1674 899 1678
rect 951 1674 955 1678
rect 1007 1674 1011 1678
rect 1031 1674 1035 1678
rect 1063 1674 1067 1678
rect 1103 1674 1107 1678
rect 1119 1674 1123 1678
rect 1175 1674 1179 1678
rect 1231 1674 1235 1678
rect 1247 1674 1251 1678
rect 1287 1674 1291 1678
rect 1319 1674 1323 1678
rect 1335 1674 1339 1678
rect 1375 1674 1379 1678
rect 1391 1674 1395 1678
rect 1423 1674 1427 1678
rect 1455 1674 1459 1678
rect 1471 1674 1475 1678
rect 1519 1674 1523 1678
rect 1583 1674 1587 1678
rect 1623 1674 1627 1678
rect 1663 1674 1667 1678
rect 111 1634 115 1638
rect 135 1634 139 1638
rect 167 1634 171 1638
rect 183 1634 187 1638
rect 215 1634 219 1638
rect 247 1634 251 1638
rect 279 1634 283 1638
rect 303 1634 307 1638
rect 343 1634 347 1638
rect 359 1634 363 1638
rect 415 1634 419 1638
rect 471 1634 475 1638
rect 487 1634 491 1638
rect 535 1634 539 1638
rect 559 1634 563 1638
rect 599 1634 603 1638
rect 631 1634 635 1638
rect 663 1634 667 1638
rect 711 1634 715 1638
rect 727 1634 731 1638
rect 791 1634 795 1638
rect 799 1634 803 1638
rect 871 1634 875 1638
rect 943 1634 947 1638
rect 951 1634 955 1638
rect 1023 1634 1027 1638
rect 1031 1634 1035 1638
rect 1103 1634 1107 1638
rect 1175 1634 1179 1638
rect 1247 1634 1251 1638
rect 1319 1634 1323 1638
rect 1391 1634 1395 1638
rect 1399 1634 1403 1638
rect 1455 1634 1459 1638
rect 1479 1634 1483 1638
rect 1519 1634 1523 1638
rect 1559 1634 1563 1638
rect 1583 1634 1587 1638
rect 1623 1634 1627 1638
rect 1663 1634 1667 1638
rect 111 1594 115 1598
rect 135 1594 139 1598
rect 167 1594 171 1598
rect 183 1594 187 1598
rect 223 1594 227 1598
rect 247 1594 251 1598
rect 279 1594 283 1598
rect 303 1594 307 1598
rect 335 1594 339 1598
rect 359 1594 363 1598
rect 383 1594 387 1598
rect 415 1594 419 1598
rect 431 1594 435 1598
rect 471 1594 475 1598
rect 479 1594 483 1598
rect 535 1594 539 1598
rect 599 1594 603 1598
rect 663 1594 667 1598
rect 727 1594 731 1598
rect 799 1594 803 1598
rect 871 1594 875 1598
rect 943 1594 947 1598
rect 951 1594 955 1598
rect 1023 1594 1027 1598
rect 1039 1594 1043 1598
rect 1103 1594 1107 1598
rect 1119 1594 1123 1598
rect 1175 1594 1179 1598
rect 1199 1594 1203 1598
rect 1247 1594 1251 1598
rect 1279 1594 1283 1598
rect 1319 1594 1323 1598
rect 1351 1594 1355 1598
rect 1399 1594 1403 1598
rect 1415 1594 1419 1598
rect 1471 1594 1475 1598
rect 1479 1594 1483 1598
rect 1527 1594 1531 1598
rect 1559 1594 1563 1598
rect 1583 1594 1587 1598
rect 1623 1594 1627 1598
rect 1663 1594 1667 1598
rect 111 1554 115 1558
rect 135 1554 139 1558
rect 167 1554 171 1558
rect 215 1554 219 1558
rect 223 1554 227 1558
rect 263 1554 267 1558
rect 279 1554 283 1558
rect 311 1554 315 1558
rect 335 1554 339 1558
rect 359 1554 363 1558
rect 383 1554 387 1558
rect 407 1554 411 1558
rect 431 1554 435 1558
rect 455 1554 459 1558
rect 479 1554 483 1558
rect 511 1554 515 1558
rect 535 1554 539 1558
rect 567 1554 571 1558
rect 599 1554 603 1558
rect 631 1554 635 1558
rect 663 1554 667 1558
rect 695 1554 699 1558
rect 727 1554 731 1558
rect 759 1554 763 1558
rect 799 1554 803 1558
rect 831 1554 835 1558
rect 871 1554 875 1558
rect 919 1554 923 1558
rect 951 1554 955 1558
rect 1007 1554 1011 1558
rect 1039 1554 1043 1558
rect 1095 1554 1099 1558
rect 1119 1554 1123 1558
rect 1183 1554 1187 1558
rect 1199 1554 1203 1558
rect 1263 1554 1267 1558
rect 1279 1554 1283 1558
rect 1335 1554 1339 1558
rect 1351 1554 1355 1558
rect 1407 1554 1411 1558
rect 1415 1554 1419 1558
rect 1471 1554 1475 1558
rect 1527 1554 1531 1558
rect 1583 1554 1587 1558
rect 1623 1554 1627 1558
rect 1663 1554 1667 1558
rect 111 1510 115 1514
rect 135 1510 139 1514
rect 167 1510 171 1514
rect 215 1510 219 1514
rect 223 1510 227 1514
rect 263 1510 267 1514
rect 295 1510 299 1514
rect 311 1510 315 1514
rect 359 1510 363 1514
rect 375 1510 379 1514
rect 407 1510 411 1514
rect 455 1510 459 1514
rect 511 1510 515 1514
rect 527 1510 531 1514
rect 567 1510 571 1514
rect 599 1510 603 1514
rect 631 1510 635 1514
rect 671 1510 675 1514
rect 695 1510 699 1514
rect 743 1510 747 1514
rect 759 1510 763 1514
rect 815 1510 819 1514
rect 831 1510 835 1514
rect 879 1510 883 1514
rect 919 1510 923 1514
rect 943 1510 947 1514
rect 1007 1510 1011 1514
rect 1063 1510 1067 1514
rect 1095 1510 1099 1514
rect 1111 1510 1115 1514
rect 1151 1510 1155 1514
rect 1183 1510 1187 1514
rect 1215 1510 1219 1514
rect 1255 1510 1259 1514
rect 1263 1510 1267 1514
rect 1295 1510 1299 1514
rect 1335 1510 1339 1514
rect 1351 1510 1355 1514
rect 1407 1510 1411 1514
rect 1415 1510 1419 1514
rect 1471 1510 1475 1514
rect 1487 1510 1491 1514
rect 1527 1510 1531 1514
rect 1567 1510 1571 1514
rect 1583 1510 1587 1514
rect 1623 1510 1627 1514
rect 1663 1510 1667 1514
rect 111 1470 115 1474
rect 135 1470 139 1474
rect 167 1470 171 1474
rect 223 1470 227 1474
rect 295 1470 299 1474
rect 375 1470 379 1474
rect 455 1470 459 1474
rect 527 1470 531 1474
rect 599 1470 603 1474
rect 663 1470 667 1474
rect 671 1470 675 1474
rect 719 1470 723 1474
rect 743 1470 747 1474
rect 783 1470 787 1474
rect 815 1470 819 1474
rect 847 1470 851 1474
rect 879 1470 883 1474
rect 903 1470 907 1474
rect 943 1470 947 1474
rect 959 1470 963 1474
rect 1007 1470 1011 1474
rect 1015 1470 1019 1474
rect 1063 1470 1067 1474
rect 1071 1470 1075 1474
rect 1111 1470 1115 1474
rect 1119 1470 1123 1474
rect 1151 1470 1155 1474
rect 1159 1470 1163 1474
rect 1183 1470 1187 1474
rect 1207 1470 1211 1474
rect 1215 1470 1219 1474
rect 1255 1470 1259 1474
rect 1263 1470 1267 1474
rect 1295 1470 1299 1474
rect 1327 1470 1331 1474
rect 1351 1470 1355 1474
rect 1399 1470 1403 1474
rect 1415 1470 1419 1474
rect 1479 1470 1483 1474
rect 1487 1470 1491 1474
rect 1559 1470 1563 1474
rect 1567 1470 1571 1474
rect 1623 1470 1627 1474
rect 1663 1470 1667 1474
rect 111 1426 115 1430
rect 135 1426 139 1430
rect 167 1426 171 1430
rect 215 1426 219 1430
rect 223 1426 227 1430
rect 287 1426 291 1430
rect 295 1426 299 1430
rect 359 1426 363 1430
rect 375 1426 379 1430
rect 439 1426 443 1430
rect 455 1426 459 1430
rect 519 1426 523 1430
rect 527 1426 531 1430
rect 599 1426 603 1430
rect 663 1426 667 1430
rect 679 1426 683 1430
rect 719 1426 723 1430
rect 759 1426 763 1430
rect 783 1426 787 1430
rect 831 1426 835 1430
rect 847 1426 851 1430
rect 903 1426 907 1430
rect 959 1426 963 1430
rect 967 1426 971 1430
rect 1015 1426 1019 1430
rect 1031 1426 1035 1430
rect 1071 1426 1075 1430
rect 1103 1426 1107 1430
rect 1119 1426 1123 1430
rect 1159 1426 1163 1430
rect 1167 1426 1171 1430
rect 1207 1426 1211 1430
rect 1231 1426 1235 1430
rect 1263 1426 1267 1430
rect 1295 1426 1299 1430
rect 1327 1426 1331 1430
rect 1359 1426 1363 1430
rect 1399 1426 1403 1430
rect 1415 1426 1419 1430
rect 1463 1426 1467 1430
rect 1479 1426 1483 1430
rect 1503 1426 1507 1430
rect 1551 1426 1555 1430
rect 1559 1426 1563 1430
rect 1591 1426 1595 1430
rect 1623 1426 1627 1430
rect 1663 1426 1667 1430
rect 111 1386 115 1390
rect 135 1386 139 1390
rect 167 1386 171 1390
rect 215 1386 219 1390
rect 223 1386 227 1390
rect 287 1386 291 1390
rect 359 1386 363 1390
rect 431 1386 435 1390
rect 439 1386 443 1390
rect 503 1386 507 1390
rect 519 1386 523 1390
rect 583 1386 587 1390
rect 599 1386 603 1390
rect 663 1386 667 1390
rect 679 1386 683 1390
rect 743 1386 747 1390
rect 759 1386 763 1390
rect 815 1386 819 1390
rect 831 1386 835 1390
rect 887 1386 891 1390
rect 903 1386 907 1390
rect 959 1386 963 1390
rect 967 1386 971 1390
rect 1031 1386 1035 1390
rect 1103 1386 1107 1390
rect 1167 1386 1171 1390
rect 1175 1386 1179 1390
rect 1231 1386 1235 1390
rect 1239 1386 1243 1390
rect 1295 1386 1299 1390
rect 1303 1386 1307 1390
rect 1359 1386 1363 1390
rect 1367 1386 1371 1390
rect 1415 1386 1419 1390
rect 1431 1386 1435 1390
rect 1463 1386 1467 1390
rect 1495 1386 1499 1390
rect 1503 1386 1507 1390
rect 1551 1386 1555 1390
rect 1567 1386 1571 1390
rect 1591 1386 1595 1390
rect 1623 1386 1627 1390
rect 1663 1386 1667 1390
rect 111 1346 115 1350
rect 135 1346 139 1350
rect 167 1346 171 1350
rect 183 1346 187 1350
rect 223 1346 227 1350
rect 239 1346 243 1350
rect 287 1346 291 1350
rect 295 1346 299 1350
rect 351 1346 355 1350
rect 359 1346 363 1350
rect 399 1346 403 1350
rect 431 1346 435 1350
rect 455 1346 459 1350
rect 503 1346 507 1350
rect 511 1346 515 1350
rect 567 1346 571 1350
rect 583 1346 587 1350
rect 631 1346 635 1350
rect 663 1346 667 1350
rect 695 1346 699 1350
rect 743 1346 747 1350
rect 759 1346 763 1350
rect 815 1346 819 1350
rect 823 1346 827 1350
rect 887 1346 891 1350
rect 959 1346 963 1350
rect 1023 1346 1027 1350
rect 1031 1346 1035 1350
rect 1087 1346 1091 1350
rect 1103 1346 1107 1350
rect 1151 1346 1155 1350
rect 1175 1346 1179 1350
rect 1215 1346 1219 1350
rect 1239 1346 1243 1350
rect 1279 1346 1283 1350
rect 1303 1346 1307 1350
rect 1343 1346 1347 1350
rect 1367 1346 1371 1350
rect 1407 1346 1411 1350
rect 1431 1346 1435 1350
rect 1479 1346 1483 1350
rect 1495 1346 1499 1350
rect 1559 1346 1563 1350
rect 1567 1346 1571 1350
rect 1623 1346 1627 1350
rect 1663 1346 1667 1350
rect 111 1302 115 1306
rect 135 1302 139 1306
rect 183 1302 187 1306
rect 231 1302 235 1306
rect 239 1302 243 1306
rect 279 1302 283 1306
rect 295 1302 299 1306
rect 327 1302 331 1306
rect 351 1302 355 1306
rect 375 1302 379 1306
rect 399 1302 403 1306
rect 431 1302 435 1306
rect 455 1302 459 1306
rect 487 1302 491 1306
rect 511 1302 515 1306
rect 543 1302 547 1306
rect 567 1302 571 1306
rect 607 1302 611 1306
rect 631 1302 635 1306
rect 663 1302 667 1306
rect 695 1302 699 1306
rect 719 1302 723 1306
rect 759 1302 763 1306
rect 775 1302 779 1306
rect 823 1302 827 1306
rect 831 1302 835 1306
rect 887 1302 891 1306
rect 895 1302 899 1306
rect 959 1302 963 1306
rect 1023 1302 1027 1306
rect 1079 1302 1083 1306
rect 1087 1302 1091 1306
rect 1143 1302 1147 1306
rect 1151 1302 1155 1306
rect 1207 1302 1211 1306
rect 1215 1302 1219 1306
rect 1279 1302 1283 1306
rect 1343 1302 1347 1306
rect 1359 1302 1363 1306
rect 1407 1302 1411 1306
rect 1447 1302 1451 1306
rect 1479 1302 1483 1306
rect 1543 1302 1547 1306
rect 1559 1302 1563 1306
rect 1623 1302 1627 1306
rect 1663 1302 1667 1306
rect 111 1262 115 1266
rect 135 1262 139 1266
rect 167 1262 171 1266
rect 183 1262 187 1266
rect 223 1262 227 1266
rect 231 1262 235 1266
rect 279 1262 283 1266
rect 327 1262 331 1266
rect 375 1262 379 1266
rect 383 1262 387 1266
rect 431 1262 435 1266
rect 439 1262 443 1266
rect 487 1262 491 1266
rect 495 1262 499 1266
rect 543 1262 547 1266
rect 551 1262 555 1266
rect 607 1262 611 1266
rect 663 1262 667 1266
rect 719 1262 723 1266
rect 767 1262 771 1266
rect 775 1262 779 1266
rect 815 1262 819 1266
rect 831 1262 835 1266
rect 871 1262 875 1266
rect 895 1262 899 1266
rect 927 1262 931 1266
rect 959 1262 963 1266
rect 983 1262 987 1266
rect 1023 1262 1027 1266
rect 1039 1262 1043 1266
rect 1079 1262 1083 1266
rect 1095 1262 1099 1266
rect 1143 1262 1147 1266
rect 1159 1262 1163 1266
rect 1207 1262 1211 1266
rect 1231 1262 1235 1266
rect 1279 1262 1283 1266
rect 1319 1262 1323 1266
rect 1359 1262 1363 1266
rect 1423 1262 1427 1266
rect 1447 1262 1451 1266
rect 1535 1262 1539 1266
rect 1543 1262 1547 1266
rect 1623 1262 1627 1266
rect 1663 1262 1667 1266
rect 111 1218 115 1222
rect 135 1218 139 1222
rect 167 1218 171 1222
rect 223 1218 227 1222
rect 279 1218 283 1222
rect 327 1218 331 1222
rect 335 1218 339 1222
rect 383 1218 387 1222
rect 431 1218 435 1222
rect 439 1218 443 1222
rect 487 1218 491 1222
rect 495 1218 499 1222
rect 543 1218 547 1222
rect 551 1218 555 1222
rect 599 1218 603 1222
rect 607 1218 611 1222
rect 655 1218 659 1222
rect 663 1218 667 1222
rect 711 1218 715 1222
rect 719 1218 723 1222
rect 767 1218 771 1222
rect 815 1218 819 1222
rect 823 1218 827 1222
rect 871 1218 875 1222
rect 887 1218 891 1222
rect 927 1218 931 1222
rect 951 1218 955 1222
rect 983 1218 987 1222
rect 1015 1218 1019 1222
rect 1039 1218 1043 1222
rect 1079 1218 1083 1222
rect 1095 1218 1099 1222
rect 1143 1218 1147 1222
rect 1159 1218 1163 1222
rect 1207 1218 1211 1222
rect 1231 1218 1235 1222
rect 1279 1218 1283 1222
rect 1319 1218 1323 1222
rect 1359 1218 1363 1222
rect 1423 1218 1427 1222
rect 1447 1218 1451 1222
rect 1535 1218 1539 1222
rect 1543 1218 1547 1222
rect 1623 1218 1627 1222
rect 1663 1218 1667 1222
rect 111 1174 115 1178
rect 135 1174 139 1178
rect 167 1174 171 1178
rect 223 1174 227 1178
rect 279 1174 283 1178
rect 287 1174 291 1178
rect 335 1174 339 1178
rect 351 1174 355 1178
rect 383 1174 387 1178
rect 415 1174 419 1178
rect 431 1174 435 1178
rect 471 1174 475 1178
rect 487 1174 491 1178
rect 535 1174 539 1178
rect 543 1174 547 1178
rect 599 1174 603 1178
rect 655 1174 659 1178
rect 663 1174 667 1178
rect 711 1174 715 1178
rect 727 1174 731 1178
rect 767 1174 771 1178
rect 783 1174 787 1178
rect 823 1174 827 1178
rect 839 1174 843 1178
rect 887 1174 891 1178
rect 903 1174 907 1178
rect 951 1174 955 1178
rect 967 1174 971 1178
rect 1015 1174 1019 1178
rect 1031 1174 1035 1178
rect 1079 1174 1083 1178
rect 1095 1174 1099 1178
rect 1143 1174 1147 1178
rect 1159 1174 1163 1178
rect 1207 1174 1211 1178
rect 1215 1174 1219 1178
rect 1279 1174 1283 1178
rect 1343 1174 1347 1178
rect 1359 1174 1363 1178
rect 1407 1174 1411 1178
rect 1447 1174 1451 1178
rect 1479 1174 1483 1178
rect 1543 1174 1547 1178
rect 1559 1174 1563 1178
rect 1623 1174 1627 1178
rect 1663 1174 1667 1178
rect 111 1130 115 1134
rect 135 1130 139 1134
rect 143 1130 147 1134
rect 167 1130 171 1134
rect 175 1130 179 1134
rect 215 1130 219 1134
rect 223 1130 227 1134
rect 271 1130 275 1134
rect 287 1130 291 1134
rect 335 1130 339 1134
rect 351 1130 355 1134
rect 399 1130 403 1134
rect 415 1130 419 1134
rect 463 1130 467 1134
rect 471 1130 475 1134
rect 527 1130 531 1134
rect 535 1130 539 1134
rect 599 1130 603 1134
rect 663 1130 667 1134
rect 727 1130 731 1134
rect 783 1130 787 1134
rect 791 1130 795 1134
rect 839 1130 843 1134
rect 855 1130 859 1134
rect 903 1130 907 1134
rect 911 1130 915 1134
rect 967 1130 971 1134
rect 1023 1130 1027 1134
rect 1031 1130 1035 1134
rect 1087 1130 1091 1134
rect 1095 1130 1099 1134
rect 1151 1130 1155 1134
rect 1159 1130 1163 1134
rect 1215 1130 1219 1134
rect 1279 1130 1283 1134
rect 1335 1130 1339 1134
rect 1343 1130 1347 1134
rect 1391 1130 1395 1134
rect 1407 1130 1411 1134
rect 1447 1130 1451 1134
rect 1479 1130 1483 1134
rect 1495 1130 1499 1134
rect 1543 1130 1547 1134
rect 1559 1130 1563 1134
rect 1591 1130 1595 1134
rect 1623 1130 1627 1134
rect 1663 1130 1667 1134
rect 111 1086 115 1090
rect 143 1086 147 1090
rect 175 1086 179 1090
rect 215 1086 219 1090
rect 247 1086 251 1090
rect 271 1086 275 1090
rect 279 1086 283 1090
rect 311 1086 315 1090
rect 335 1086 339 1090
rect 351 1086 355 1090
rect 391 1086 395 1090
rect 399 1086 403 1090
rect 439 1086 443 1090
rect 463 1086 467 1090
rect 503 1086 507 1090
rect 527 1086 531 1090
rect 575 1086 579 1090
rect 599 1086 603 1090
rect 655 1086 659 1090
rect 663 1086 667 1090
rect 727 1086 731 1090
rect 735 1086 739 1090
rect 791 1086 795 1090
rect 815 1086 819 1090
rect 855 1086 859 1090
rect 895 1086 899 1090
rect 911 1086 915 1090
rect 967 1086 971 1090
rect 1023 1086 1027 1090
rect 1039 1086 1043 1090
rect 1087 1086 1091 1090
rect 1111 1086 1115 1090
rect 1151 1086 1155 1090
rect 1175 1086 1179 1090
rect 1215 1086 1219 1090
rect 1239 1086 1243 1090
rect 1279 1086 1283 1090
rect 1303 1086 1307 1090
rect 1335 1086 1339 1090
rect 1359 1086 1363 1090
rect 1391 1086 1395 1090
rect 1415 1086 1419 1090
rect 1447 1086 1451 1090
rect 1463 1086 1467 1090
rect 1495 1086 1499 1090
rect 1503 1086 1507 1090
rect 1543 1086 1547 1090
rect 1551 1086 1555 1090
rect 1591 1086 1595 1090
rect 1623 1086 1627 1090
rect 1663 1086 1667 1090
rect 111 1042 115 1046
rect 215 1042 219 1046
rect 247 1042 251 1046
rect 279 1042 283 1046
rect 295 1042 299 1046
rect 311 1042 315 1046
rect 327 1042 331 1046
rect 351 1042 355 1046
rect 359 1042 363 1046
rect 391 1042 395 1046
rect 423 1042 427 1046
rect 439 1042 443 1046
rect 455 1042 459 1046
rect 503 1042 507 1046
rect 559 1042 563 1046
rect 575 1042 579 1046
rect 631 1042 635 1046
rect 655 1042 659 1046
rect 711 1042 715 1046
rect 735 1042 739 1046
rect 799 1042 803 1046
rect 815 1042 819 1046
rect 879 1042 883 1046
rect 895 1042 899 1046
rect 959 1042 963 1046
rect 967 1042 971 1046
rect 1031 1042 1035 1046
rect 1039 1042 1043 1046
rect 1095 1042 1099 1046
rect 1111 1042 1115 1046
rect 1159 1042 1163 1046
rect 1175 1042 1179 1046
rect 1223 1042 1227 1046
rect 1239 1042 1243 1046
rect 1279 1042 1283 1046
rect 1303 1042 1307 1046
rect 1335 1042 1339 1046
rect 1359 1042 1363 1046
rect 1383 1042 1387 1046
rect 1415 1042 1419 1046
rect 1431 1042 1435 1046
rect 1463 1042 1467 1046
rect 1479 1042 1483 1046
rect 1503 1042 1507 1046
rect 1535 1042 1539 1046
rect 1551 1042 1555 1046
rect 1591 1042 1595 1046
rect 1623 1042 1627 1046
rect 1663 1042 1667 1046
rect 111 1002 115 1006
rect 247 1002 251 1006
rect 279 1002 283 1006
rect 295 1002 299 1006
rect 311 1002 315 1006
rect 327 1002 331 1006
rect 343 1002 347 1006
rect 359 1002 363 1006
rect 383 1002 387 1006
rect 391 1002 395 1006
rect 423 1002 427 1006
rect 455 1002 459 1006
rect 479 1002 483 1006
rect 503 1002 507 1006
rect 543 1002 547 1006
rect 559 1002 563 1006
rect 615 1002 619 1006
rect 631 1002 635 1006
rect 687 1002 691 1006
rect 711 1002 715 1006
rect 759 1002 763 1006
rect 799 1002 803 1006
rect 831 1002 835 1006
rect 879 1002 883 1006
rect 903 1002 907 1006
rect 959 1002 963 1006
rect 967 1002 971 1006
rect 1031 1002 1035 1006
rect 1095 1002 1099 1006
rect 1159 1002 1163 1006
rect 1223 1002 1227 1006
rect 1279 1002 1283 1006
rect 1287 1002 1291 1006
rect 1335 1002 1339 1006
rect 1343 1002 1347 1006
rect 1383 1002 1387 1006
rect 1399 1002 1403 1006
rect 1431 1002 1435 1006
rect 1447 1002 1451 1006
rect 1479 1002 1483 1006
rect 1495 1002 1499 1006
rect 1535 1002 1539 1006
rect 1543 1002 1547 1006
rect 1591 1002 1595 1006
rect 1623 1002 1627 1006
rect 1663 1002 1667 1006
rect 111 962 115 966
rect 167 962 171 966
rect 199 962 203 966
rect 239 962 243 966
rect 247 962 251 966
rect 279 962 283 966
rect 287 962 291 966
rect 311 962 315 966
rect 343 962 347 966
rect 383 962 387 966
rect 407 962 411 966
rect 423 962 427 966
rect 471 962 475 966
rect 479 962 483 966
rect 535 962 539 966
rect 543 962 547 966
rect 599 962 603 966
rect 615 962 619 966
rect 663 962 667 966
rect 687 962 691 966
rect 727 962 731 966
rect 759 962 763 966
rect 791 962 795 966
rect 831 962 835 966
rect 847 962 851 966
rect 903 962 907 966
rect 911 962 915 966
rect 967 962 971 966
rect 975 962 979 966
rect 1031 962 1035 966
rect 1039 962 1043 966
rect 1095 962 1099 966
rect 1103 962 1107 966
rect 1159 962 1163 966
rect 1167 962 1171 966
rect 1223 962 1227 966
rect 1231 962 1235 966
rect 1287 962 1291 966
rect 1343 962 1347 966
rect 1391 962 1395 966
rect 1399 962 1403 966
rect 1431 962 1435 966
rect 1447 962 1451 966
rect 1471 962 1475 966
rect 1495 962 1499 966
rect 1511 962 1515 966
rect 1543 962 1547 966
rect 1551 962 1555 966
rect 1591 962 1595 966
rect 1623 962 1627 966
rect 1663 962 1667 966
rect 111 918 115 922
rect 135 918 139 922
rect 167 918 171 922
rect 199 918 203 922
rect 207 918 211 922
rect 239 918 243 922
rect 271 918 275 922
rect 287 918 291 922
rect 335 918 339 922
rect 343 918 347 922
rect 407 918 411 922
rect 471 918 475 922
rect 535 918 539 922
rect 591 918 595 922
rect 599 918 603 922
rect 647 918 651 922
rect 663 918 667 922
rect 703 918 707 922
rect 727 918 731 922
rect 751 918 755 922
rect 791 918 795 922
rect 799 918 803 922
rect 847 918 851 922
rect 903 918 907 922
rect 911 918 915 922
rect 959 918 963 922
rect 975 918 979 922
rect 1023 918 1027 922
rect 1039 918 1043 922
rect 1087 918 1091 922
rect 1103 918 1107 922
rect 1143 918 1147 922
rect 1167 918 1171 922
rect 1199 918 1203 922
rect 1231 918 1235 922
rect 1255 918 1259 922
rect 1287 918 1291 922
rect 1319 918 1323 922
rect 1343 918 1347 922
rect 1383 918 1387 922
rect 1391 918 1395 922
rect 1431 918 1435 922
rect 1471 918 1475 922
rect 1511 918 1515 922
rect 1551 918 1555 922
rect 1591 918 1595 922
rect 1623 918 1627 922
rect 1663 918 1667 922
rect 111 874 115 878
rect 135 874 139 878
rect 167 874 171 878
rect 207 874 211 878
rect 271 874 275 878
rect 335 874 339 878
rect 407 874 411 878
rect 471 874 475 878
rect 535 874 539 878
rect 591 874 595 878
rect 599 874 603 878
rect 647 874 651 878
rect 655 874 659 878
rect 703 874 707 878
rect 751 874 755 878
rect 799 874 803 878
rect 847 874 851 878
rect 903 874 907 878
rect 959 874 963 878
rect 967 874 971 878
rect 1023 874 1027 878
rect 1039 874 1043 878
rect 1087 874 1091 878
rect 1103 874 1107 878
rect 1143 874 1147 878
rect 1167 874 1171 878
rect 1199 874 1203 878
rect 1231 874 1235 878
rect 1255 874 1259 878
rect 1287 874 1291 878
rect 1319 874 1323 878
rect 1343 874 1347 878
rect 1383 874 1387 878
rect 1399 874 1403 878
rect 1463 874 1467 878
rect 1663 874 1667 878
rect 111 834 115 838
rect 135 834 139 838
rect 167 834 171 838
rect 207 834 211 838
rect 215 834 219 838
rect 271 834 275 838
rect 279 834 283 838
rect 335 834 339 838
rect 343 834 347 838
rect 407 834 411 838
rect 415 834 419 838
rect 471 834 475 838
rect 479 834 483 838
rect 535 834 539 838
rect 543 834 547 838
rect 599 834 603 838
rect 607 834 611 838
rect 655 834 659 838
rect 671 834 675 838
rect 703 834 707 838
rect 735 834 739 838
rect 751 834 755 838
rect 791 834 795 838
rect 799 834 803 838
rect 847 834 851 838
rect 903 834 907 838
rect 911 834 915 838
rect 967 834 971 838
rect 975 834 979 838
rect 1039 834 1043 838
rect 1103 834 1107 838
rect 1111 834 1115 838
rect 1167 834 1171 838
rect 1183 834 1187 838
rect 1231 834 1235 838
rect 1247 834 1251 838
rect 1287 834 1291 838
rect 1311 834 1315 838
rect 1343 834 1347 838
rect 1367 834 1371 838
rect 1399 834 1403 838
rect 1423 834 1427 838
rect 1463 834 1467 838
rect 1479 834 1483 838
rect 1535 834 1539 838
rect 1591 834 1595 838
rect 1663 834 1667 838
rect 111 790 115 794
rect 135 790 139 794
rect 167 790 171 794
rect 175 790 179 794
rect 215 790 219 794
rect 231 790 235 794
rect 279 790 283 794
rect 295 790 299 794
rect 343 790 347 794
rect 367 790 371 794
rect 415 790 419 794
rect 447 790 451 794
rect 479 790 483 794
rect 527 790 531 794
rect 543 790 547 794
rect 607 790 611 794
rect 615 790 619 794
rect 671 790 675 794
rect 703 790 707 794
rect 735 790 739 794
rect 791 790 795 794
rect 847 790 851 794
rect 871 790 875 794
rect 911 790 915 794
rect 951 790 955 794
rect 975 790 979 794
rect 1023 790 1027 794
rect 1039 790 1043 794
rect 1095 790 1099 794
rect 1111 790 1115 794
rect 1167 790 1171 794
rect 1183 790 1187 794
rect 1231 790 1235 794
rect 1247 790 1251 794
rect 1295 790 1299 794
rect 1311 790 1315 794
rect 1359 790 1363 794
rect 1367 790 1371 794
rect 1415 790 1419 794
rect 1423 790 1427 794
rect 1471 790 1475 794
rect 1479 790 1483 794
rect 1527 790 1531 794
rect 1535 790 1539 794
rect 1591 790 1595 794
rect 1663 790 1667 794
rect 111 750 115 754
rect 135 750 139 754
rect 175 750 179 754
rect 215 750 219 754
rect 231 750 235 754
rect 247 750 251 754
rect 279 750 283 754
rect 295 750 299 754
rect 319 750 323 754
rect 359 750 363 754
rect 367 750 371 754
rect 399 750 403 754
rect 439 750 443 754
rect 447 750 451 754
rect 487 750 491 754
rect 527 750 531 754
rect 543 750 547 754
rect 607 750 611 754
rect 615 750 619 754
rect 671 750 675 754
rect 703 750 707 754
rect 735 750 739 754
rect 791 750 795 754
rect 799 750 803 754
rect 863 750 867 754
rect 871 750 875 754
rect 927 750 931 754
rect 951 750 955 754
rect 991 750 995 754
rect 1023 750 1027 754
rect 1055 750 1059 754
rect 1095 750 1099 754
rect 1119 750 1123 754
rect 1167 750 1171 754
rect 1183 750 1187 754
rect 1231 750 1235 754
rect 1239 750 1243 754
rect 1295 750 1299 754
rect 1351 750 1355 754
rect 1359 750 1363 754
rect 1407 750 1411 754
rect 1415 750 1419 754
rect 1463 750 1467 754
rect 1471 750 1475 754
rect 1519 750 1523 754
rect 1527 750 1531 754
rect 1583 750 1587 754
rect 1591 750 1595 754
rect 1623 750 1627 754
rect 1663 750 1667 754
rect 111 706 115 710
rect 215 706 219 710
rect 247 706 251 710
rect 279 706 283 710
rect 311 706 315 710
rect 319 706 323 710
rect 343 706 347 710
rect 359 706 363 710
rect 375 706 379 710
rect 399 706 403 710
rect 407 706 411 710
rect 439 706 443 710
rect 471 706 475 710
rect 487 706 491 710
rect 503 706 507 710
rect 543 706 547 710
rect 591 706 595 710
rect 607 706 611 710
rect 647 706 651 710
rect 671 706 675 710
rect 703 706 707 710
rect 735 706 739 710
rect 759 706 763 710
rect 799 706 803 710
rect 823 706 827 710
rect 863 706 867 710
rect 887 706 891 710
rect 927 706 931 710
rect 959 706 963 710
rect 991 706 995 710
rect 1023 706 1027 710
rect 1055 706 1059 710
rect 1087 706 1091 710
rect 1119 706 1123 710
rect 1159 706 1163 710
rect 1183 706 1187 710
rect 1223 706 1227 710
rect 1239 706 1243 710
rect 1287 706 1291 710
rect 1295 706 1299 710
rect 1351 706 1355 710
rect 1407 706 1411 710
rect 1415 706 1419 710
rect 1463 706 1467 710
rect 1471 706 1475 710
rect 1519 706 1523 710
rect 1527 706 1531 710
rect 1583 706 1587 710
rect 1623 706 1627 710
rect 1663 706 1667 710
rect 111 666 115 670
rect 279 666 283 670
rect 295 666 299 670
rect 311 666 315 670
rect 327 666 331 670
rect 343 666 347 670
rect 359 666 363 670
rect 375 666 379 670
rect 391 666 395 670
rect 407 666 411 670
rect 423 666 427 670
rect 439 666 443 670
rect 455 666 459 670
rect 471 666 475 670
rect 487 666 491 670
rect 503 666 507 670
rect 519 666 523 670
rect 543 666 547 670
rect 551 666 555 670
rect 591 666 595 670
rect 639 666 643 670
rect 647 666 651 670
rect 687 666 691 670
rect 703 666 707 670
rect 735 666 739 670
rect 759 666 763 670
rect 791 666 795 670
rect 823 666 827 670
rect 847 666 851 670
rect 887 666 891 670
rect 911 666 915 670
rect 959 666 963 670
rect 975 666 979 670
rect 1023 666 1027 670
rect 1047 666 1051 670
rect 1087 666 1091 670
rect 1127 666 1131 670
rect 1159 666 1163 670
rect 1215 666 1219 670
rect 1223 666 1227 670
rect 1287 666 1291 670
rect 1295 666 1299 670
rect 1351 666 1355 670
rect 1383 666 1387 670
rect 1415 666 1419 670
rect 1471 666 1475 670
rect 1527 666 1531 670
rect 1559 666 1563 670
rect 1583 666 1587 670
rect 1623 666 1627 670
rect 1663 666 1667 670
rect 111 626 115 630
rect 247 626 251 630
rect 279 626 283 630
rect 295 626 299 630
rect 319 626 323 630
rect 327 626 331 630
rect 359 626 363 630
rect 367 626 371 630
rect 391 626 395 630
rect 423 626 427 630
rect 455 626 459 630
rect 471 626 475 630
rect 487 626 491 630
rect 519 626 523 630
rect 551 626 555 630
rect 567 626 571 630
rect 591 626 595 630
rect 615 626 619 630
rect 639 626 643 630
rect 663 626 667 630
rect 687 626 691 630
rect 719 626 723 630
rect 735 626 739 630
rect 775 626 779 630
rect 791 626 795 630
rect 831 626 835 630
rect 847 626 851 630
rect 895 626 899 630
rect 911 626 915 630
rect 967 626 971 630
rect 975 626 979 630
rect 1047 626 1051 630
rect 1127 626 1131 630
rect 1207 626 1211 630
rect 1215 626 1219 630
rect 1287 626 1291 630
rect 1295 626 1299 630
rect 1359 626 1363 630
rect 1383 626 1387 630
rect 1431 626 1435 630
rect 1471 626 1475 630
rect 1503 626 1507 630
rect 1559 626 1563 630
rect 1575 626 1579 630
rect 1623 626 1627 630
rect 1663 626 1667 630
rect 111 586 115 590
rect 167 586 171 590
rect 215 586 219 590
rect 247 586 251 590
rect 271 586 275 590
rect 279 586 283 590
rect 319 586 323 590
rect 335 586 339 590
rect 367 586 371 590
rect 407 586 411 590
rect 423 586 427 590
rect 471 586 475 590
rect 487 586 491 590
rect 519 586 523 590
rect 559 586 563 590
rect 567 586 571 590
rect 615 586 619 590
rect 631 586 635 590
rect 663 586 667 590
rect 703 586 707 590
rect 719 586 723 590
rect 767 586 771 590
rect 775 586 779 590
rect 823 586 827 590
rect 831 586 835 590
rect 879 586 883 590
rect 895 586 899 590
rect 935 586 939 590
rect 967 586 971 590
rect 991 586 995 590
rect 1047 586 1051 590
rect 1103 586 1107 590
rect 1127 586 1131 590
rect 1159 586 1163 590
rect 1207 586 1211 590
rect 1215 586 1219 590
rect 1271 586 1275 590
rect 1287 586 1291 590
rect 1327 586 1331 590
rect 1359 586 1363 590
rect 1383 586 1387 590
rect 1431 586 1435 590
rect 1447 586 1451 590
rect 1503 586 1507 590
rect 1511 586 1515 590
rect 1575 586 1579 590
rect 1623 586 1627 590
rect 1663 586 1667 590
rect 111 542 115 546
rect 135 542 139 546
rect 167 542 171 546
rect 199 542 203 546
rect 215 542 219 546
rect 231 542 235 546
rect 271 542 275 546
rect 279 542 283 546
rect 327 542 331 546
rect 335 542 339 546
rect 375 542 379 546
rect 407 542 411 546
rect 431 542 435 546
rect 487 542 491 546
rect 495 542 499 546
rect 559 542 563 546
rect 623 542 627 546
rect 631 542 635 546
rect 687 542 691 546
rect 703 542 707 546
rect 751 542 755 546
rect 767 542 771 546
rect 815 542 819 546
rect 823 542 827 546
rect 879 542 883 546
rect 935 542 939 546
rect 943 542 947 546
rect 991 542 995 546
rect 1007 542 1011 546
rect 1047 542 1051 546
rect 1071 542 1075 546
rect 1103 542 1107 546
rect 1127 542 1131 546
rect 1159 542 1163 546
rect 1183 542 1187 546
rect 1215 542 1219 546
rect 1231 542 1235 546
rect 1271 542 1275 546
rect 1279 542 1283 546
rect 1327 542 1331 546
rect 1335 542 1339 546
rect 1383 542 1387 546
rect 1391 542 1395 546
rect 1447 542 1451 546
rect 1511 542 1515 546
rect 1575 542 1579 546
rect 1623 542 1627 546
rect 1663 542 1667 546
rect 111 502 115 506
rect 135 502 139 506
rect 167 502 171 506
rect 199 502 203 506
rect 231 502 235 506
rect 239 502 243 506
rect 279 502 283 506
rect 287 502 291 506
rect 327 502 331 506
rect 375 502 379 506
rect 423 502 427 506
rect 431 502 435 506
rect 479 502 483 506
rect 495 502 499 506
rect 543 502 547 506
rect 559 502 563 506
rect 615 502 619 506
rect 623 502 627 506
rect 687 502 691 506
rect 695 502 699 506
rect 751 502 755 506
rect 775 502 779 506
rect 815 502 819 506
rect 847 502 851 506
rect 879 502 883 506
rect 919 502 923 506
rect 943 502 947 506
rect 983 502 987 506
rect 1007 502 1011 506
rect 1039 502 1043 506
rect 1071 502 1075 506
rect 1095 502 1099 506
rect 1127 502 1131 506
rect 1143 502 1147 506
rect 1183 502 1187 506
rect 1191 502 1195 506
rect 1231 502 1235 506
rect 1239 502 1243 506
rect 1279 502 1283 506
rect 1287 502 1291 506
rect 1335 502 1339 506
rect 1383 502 1387 506
rect 1391 502 1395 506
rect 1431 502 1435 506
rect 1447 502 1451 506
rect 1479 502 1483 506
rect 1511 502 1515 506
rect 1535 502 1539 506
rect 1575 502 1579 506
rect 1591 502 1595 506
rect 1623 502 1627 506
rect 1663 502 1667 506
rect 111 462 115 466
rect 135 462 139 466
rect 151 462 155 466
rect 167 462 171 466
rect 199 462 203 466
rect 207 462 211 466
rect 239 462 243 466
rect 255 462 259 466
rect 287 462 291 466
rect 311 462 315 466
rect 327 462 331 466
rect 367 462 371 466
rect 375 462 379 466
rect 423 462 427 466
rect 439 462 443 466
rect 479 462 483 466
rect 519 462 523 466
rect 543 462 547 466
rect 599 462 603 466
rect 615 462 619 466
rect 679 462 683 466
rect 695 462 699 466
rect 759 462 763 466
rect 775 462 779 466
rect 839 462 843 466
rect 847 462 851 466
rect 911 462 915 466
rect 919 462 923 466
rect 983 462 987 466
rect 1039 462 1043 466
rect 1055 462 1059 466
rect 1095 462 1099 466
rect 1127 462 1131 466
rect 1143 462 1147 466
rect 1191 462 1195 466
rect 1199 462 1203 466
rect 1239 462 1243 466
rect 1263 462 1267 466
rect 1287 462 1291 466
rect 1319 462 1323 466
rect 1335 462 1339 466
rect 1375 462 1379 466
rect 1383 462 1387 466
rect 1431 462 1435 466
rect 1479 462 1483 466
rect 1495 462 1499 466
rect 1535 462 1539 466
rect 1591 462 1595 466
rect 1623 462 1627 466
rect 1663 462 1667 466
rect 111 422 115 426
rect 151 422 155 426
rect 175 422 179 426
rect 207 422 211 426
rect 223 422 227 426
rect 255 422 259 426
rect 271 422 275 426
rect 311 422 315 426
rect 319 422 323 426
rect 367 422 371 426
rect 415 422 419 426
rect 439 422 443 426
rect 471 422 475 426
rect 519 422 523 426
rect 527 422 531 426
rect 591 422 595 426
rect 599 422 603 426
rect 663 422 667 426
rect 679 422 683 426
rect 735 422 739 426
rect 759 422 763 426
rect 807 422 811 426
rect 839 422 843 426
rect 871 422 875 426
rect 911 422 915 426
rect 935 422 939 426
rect 983 422 987 426
rect 991 422 995 426
rect 1039 422 1043 426
rect 1055 422 1059 426
rect 1087 422 1091 426
rect 1127 422 1131 426
rect 1167 422 1171 426
rect 1199 422 1203 426
rect 1207 422 1211 426
rect 1247 422 1251 426
rect 1263 422 1267 426
rect 1287 422 1291 426
rect 1319 422 1323 426
rect 1335 422 1339 426
rect 1375 422 1379 426
rect 1383 422 1387 426
rect 1431 422 1435 426
rect 1495 422 1499 426
rect 1663 422 1667 426
rect 111 378 115 382
rect 135 378 139 382
rect 167 378 171 382
rect 175 378 179 382
rect 199 378 203 382
rect 223 378 227 382
rect 239 378 243 382
rect 271 378 275 382
rect 295 378 299 382
rect 319 378 323 382
rect 351 378 355 382
rect 367 378 371 382
rect 407 378 411 382
rect 415 378 419 382
rect 463 378 467 382
rect 471 378 475 382
rect 519 378 523 382
rect 527 378 531 382
rect 575 378 579 382
rect 591 378 595 382
rect 631 378 635 382
rect 663 378 667 382
rect 687 378 691 382
rect 735 378 739 382
rect 743 378 747 382
rect 799 378 803 382
rect 807 378 811 382
rect 855 378 859 382
rect 871 378 875 382
rect 919 378 923 382
rect 935 378 939 382
rect 983 378 987 382
rect 991 378 995 382
rect 1039 378 1043 382
rect 1087 378 1091 382
rect 1095 378 1099 382
rect 1127 378 1131 382
rect 1151 378 1155 382
rect 1167 378 1171 382
rect 1207 378 1211 382
rect 1247 378 1251 382
rect 1255 378 1259 382
rect 1287 378 1291 382
rect 1303 378 1307 382
rect 1335 378 1339 382
rect 1351 378 1355 382
rect 1383 378 1387 382
rect 1399 378 1403 382
rect 1447 378 1451 382
rect 1495 378 1499 382
rect 1543 378 1547 382
rect 1591 378 1595 382
rect 1623 378 1627 382
rect 1663 378 1667 382
rect 111 338 115 342
rect 135 338 139 342
rect 167 338 171 342
rect 199 338 203 342
rect 207 338 211 342
rect 239 338 243 342
rect 263 338 267 342
rect 295 338 299 342
rect 327 338 331 342
rect 351 338 355 342
rect 391 338 395 342
rect 407 338 411 342
rect 455 338 459 342
rect 463 338 467 342
rect 519 338 523 342
rect 575 338 579 342
rect 631 338 635 342
rect 687 338 691 342
rect 743 338 747 342
rect 751 338 755 342
rect 799 338 803 342
rect 815 338 819 342
rect 855 338 859 342
rect 879 338 883 342
rect 919 338 923 342
rect 951 338 955 342
rect 983 338 987 342
rect 1031 338 1035 342
rect 1039 338 1043 342
rect 1095 338 1099 342
rect 1111 338 1115 342
rect 1151 338 1155 342
rect 1191 338 1195 342
rect 1207 338 1211 342
rect 1255 338 1259 342
rect 1271 338 1275 342
rect 1303 338 1307 342
rect 1343 338 1347 342
rect 1351 338 1355 342
rect 1399 338 1403 342
rect 1407 338 1411 342
rect 1447 338 1451 342
rect 1463 338 1467 342
rect 1495 338 1499 342
rect 1519 338 1523 342
rect 1543 338 1547 342
rect 1583 338 1587 342
rect 1591 338 1595 342
rect 1623 338 1627 342
rect 1663 338 1667 342
rect 111 298 115 302
rect 135 298 139 302
rect 167 298 171 302
rect 207 298 211 302
rect 231 298 235 302
rect 263 298 267 302
rect 295 298 299 302
rect 327 298 331 302
rect 367 298 371 302
rect 391 298 395 302
rect 439 298 443 302
rect 455 298 459 302
rect 503 298 507 302
rect 519 298 523 302
rect 567 298 571 302
rect 575 298 579 302
rect 631 298 635 302
rect 687 298 691 302
rect 743 298 747 302
rect 751 298 755 302
rect 807 298 811 302
rect 815 298 819 302
rect 879 298 883 302
rect 951 298 955 302
rect 1031 298 1035 302
rect 1111 298 1115 302
rect 1191 298 1195 302
rect 1263 298 1267 302
rect 1271 298 1275 302
rect 1327 298 1331 302
rect 1343 298 1347 302
rect 1391 298 1395 302
rect 1407 298 1411 302
rect 1447 298 1451 302
rect 1463 298 1467 302
rect 1495 298 1499 302
rect 1519 298 1523 302
rect 1543 298 1547 302
rect 1583 298 1587 302
rect 1591 298 1595 302
rect 1623 298 1627 302
rect 1663 298 1667 302
rect 111 254 115 258
rect 135 254 139 258
rect 167 254 171 258
rect 175 254 179 258
rect 231 254 235 258
rect 247 254 251 258
rect 295 254 299 258
rect 319 254 323 258
rect 367 254 371 258
rect 383 254 387 258
rect 439 254 443 258
rect 447 254 451 258
rect 503 254 507 258
rect 519 254 523 258
rect 567 254 571 258
rect 591 254 595 258
rect 631 254 635 258
rect 663 254 667 258
rect 687 254 691 258
rect 743 254 747 258
rect 807 254 811 258
rect 823 254 827 258
rect 879 254 883 258
rect 895 254 899 258
rect 951 254 955 258
rect 967 254 971 258
rect 1031 254 1035 258
rect 1087 254 1091 258
rect 1111 254 1115 258
rect 1143 254 1147 258
rect 1191 254 1195 258
rect 1199 254 1203 258
rect 1255 254 1259 258
rect 1263 254 1267 258
rect 1311 254 1315 258
rect 1327 254 1331 258
rect 1367 254 1371 258
rect 1391 254 1395 258
rect 1415 254 1419 258
rect 1447 254 1451 258
rect 1463 254 1467 258
rect 1495 254 1499 258
rect 1519 254 1523 258
rect 1543 254 1547 258
rect 1575 254 1579 258
rect 1591 254 1595 258
rect 1623 254 1627 258
rect 1663 254 1667 258
rect 111 214 115 218
rect 135 214 139 218
rect 167 214 171 218
rect 175 214 179 218
rect 207 214 211 218
rect 247 214 251 218
rect 255 214 259 218
rect 303 214 307 218
rect 319 214 323 218
rect 343 214 347 218
rect 375 214 379 218
rect 383 214 387 218
rect 415 214 419 218
rect 447 214 451 218
rect 471 214 475 218
rect 519 214 523 218
rect 535 214 539 218
rect 591 214 595 218
rect 615 214 619 218
rect 663 214 667 218
rect 695 214 699 218
rect 743 214 747 218
rect 775 214 779 218
rect 823 214 827 218
rect 855 214 859 218
rect 895 214 899 218
rect 927 214 931 218
rect 967 214 971 218
rect 999 214 1003 218
rect 1031 214 1035 218
rect 1071 214 1075 218
rect 1087 214 1091 218
rect 1143 214 1147 218
rect 1199 214 1203 218
rect 1215 214 1219 218
rect 1255 214 1259 218
rect 1287 214 1291 218
rect 1311 214 1315 218
rect 1351 214 1355 218
rect 1367 214 1371 218
rect 1415 214 1419 218
rect 1463 214 1467 218
rect 1471 214 1475 218
rect 1519 214 1523 218
rect 1527 214 1531 218
rect 1575 214 1579 218
rect 1583 214 1587 218
rect 1623 214 1627 218
rect 1663 214 1667 218
rect 111 174 115 178
rect 135 174 139 178
rect 167 174 171 178
rect 175 174 179 178
rect 207 174 211 178
rect 231 174 235 178
rect 255 174 259 178
rect 287 174 291 178
rect 303 174 307 178
rect 343 174 347 178
rect 375 174 379 178
rect 399 174 403 178
rect 415 174 419 178
rect 455 174 459 178
rect 471 174 475 178
rect 511 174 515 178
rect 535 174 539 178
rect 575 174 579 178
rect 615 174 619 178
rect 639 174 643 178
rect 695 174 699 178
rect 703 174 707 178
rect 767 174 771 178
rect 775 174 779 178
rect 831 174 835 178
rect 855 174 859 178
rect 895 174 899 178
rect 927 174 931 178
rect 951 174 955 178
rect 999 174 1003 178
rect 1015 174 1019 178
rect 1071 174 1075 178
rect 1079 174 1083 178
rect 1143 174 1147 178
rect 1207 174 1211 178
rect 1215 174 1219 178
rect 1279 174 1283 178
rect 1287 174 1291 178
rect 1351 174 1355 178
rect 1415 174 1419 178
rect 1423 174 1427 178
rect 1471 174 1475 178
rect 1495 174 1499 178
rect 1527 174 1531 178
rect 1567 174 1571 178
rect 1583 174 1587 178
rect 1623 174 1627 178
rect 1663 174 1667 178
rect 111 118 115 122
rect 135 118 139 122
rect 167 118 171 122
rect 175 118 179 122
rect 199 118 203 122
rect 231 118 235 122
rect 263 118 267 122
rect 287 118 291 122
rect 295 118 299 122
rect 327 118 331 122
rect 343 118 347 122
rect 359 118 363 122
rect 391 118 395 122
rect 399 118 403 122
rect 423 118 427 122
rect 455 118 459 122
rect 463 118 467 122
rect 503 118 507 122
rect 511 118 515 122
rect 543 118 547 122
rect 575 118 579 122
rect 607 118 611 122
rect 639 118 643 122
rect 671 118 675 122
rect 703 118 707 122
rect 735 118 739 122
rect 767 118 771 122
rect 799 118 803 122
rect 831 118 835 122
rect 863 118 867 122
rect 895 118 899 122
rect 935 118 939 122
rect 951 118 955 122
rect 975 118 979 122
rect 1015 118 1019 122
rect 1063 118 1067 122
rect 1079 118 1083 122
rect 1103 118 1107 122
rect 1143 118 1147 122
rect 1183 118 1187 122
rect 1207 118 1211 122
rect 1223 118 1227 122
rect 1263 118 1267 122
rect 1279 118 1283 122
rect 1295 118 1299 122
rect 1335 118 1339 122
rect 1351 118 1355 122
rect 1375 118 1379 122
rect 1415 118 1419 122
rect 1423 118 1427 122
rect 1455 118 1459 122
rect 1495 118 1499 122
rect 1503 118 1507 122
rect 1551 118 1555 122
rect 1567 118 1571 122
rect 1591 118 1595 122
rect 1623 118 1627 122
rect 1663 118 1667 122
rect 111 78 115 82
rect 135 78 139 82
rect 167 78 171 82
rect 199 78 203 82
rect 231 78 235 82
rect 263 78 267 82
rect 295 78 299 82
rect 327 78 331 82
rect 359 78 363 82
rect 391 78 395 82
rect 423 78 427 82
rect 463 78 467 82
rect 503 78 507 82
rect 543 78 547 82
rect 575 78 579 82
rect 607 78 611 82
rect 639 78 643 82
rect 671 78 675 82
rect 703 78 707 82
rect 735 78 739 82
rect 767 78 771 82
rect 799 78 803 82
rect 831 78 835 82
rect 863 78 867 82
rect 895 78 899 82
rect 935 78 939 82
rect 975 78 979 82
rect 1015 78 1019 82
rect 1063 78 1067 82
rect 1103 78 1107 82
rect 1143 78 1147 82
rect 1183 78 1187 82
rect 1223 78 1227 82
rect 1263 78 1267 82
rect 1295 78 1299 82
rect 1335 78 1339 82
rect 1375 78 1379 82
rect 1415 78 1419 82
rect 1455 78 1459 82
rect 1503 78 1507 82
rect 1551 78 1555 82
rect 1591 78 1595 82
rect 1623 78 1627 82
rect 1663 78 1667 82
<< m4 >>
rect 96 1713 97 1719
rect 103 1718 1699 1719
rect 103 1714 111 1718
rect 115 1714 255 1718
rect 259 1714 287 1718
rect 291 1714 319 1718
rect 323 1714 359 1718
rect 363 1714 407 1718
rect 411 1714 455 1718
rect 459 1714 503 1718
rect 507 1714 551 1718
rect 555 1714 607 1718
rect 611 1714 663 1718
rect 667 1714 727 1718
rect 731 1714 783 1718
rect 787 1714 839 1718
rect 843 1714 895 1718
rect 899 1714 951 1718
rect 955 1714 1007 1718
rect 1011 1714 1063 1718
rect 1067 1714 1119 1718
rect 1123 1714 1175 1718
rect 1179 1714 1231 1718
rect 1235 1714 1287 1718
rect 1291 1714 1335 1718
rect 1339 1714 1375 1718
rect 1379 1714 1423 1718
rect 1427 1714 1471 1718
rect 1475 1714 1519 1718
rect 1523 1714 1663 1718
rect 1667 1714 1699 1718
rect 103 1713 1699 1714
rect 1705 1713 1706 1719
rect 84 1673 85 1679
rect 91 1678 1687 1679
rect 91 1674 111 1678
rect 115 1674 135 1678
rect 139 1674 167 1678
rect 171 1674 215 1678
rect 219 1674 255 1678
rect 259 1674 279 1678
rect 283 1674 287 1678
rect 291 1674 319 1678
rect 323 1674 343 1678
rect 347 1674 359 1678
rect 363 1674 407 1678
rect 411 1674 415 1678
rect 419 1674 455 1678
rect 459 1674 487 1678
rect 491 1674 503 1678
rect 507 1674 551 1678
rect 555 1674 559 1678
rect 563 1674 607 1678
rect 611 1674 631 1678
rect 635 1674 663 1678
rect 667 1674 711 1678
rect 715 1674 727 1678
rect 731 1674 783 1678
rect 787 1674 791 1678
rect 795 1674 839 1678
rect 843 1674 871 1678
rect 875 1674 895 1678
rect 899 1674 951 1678
rect 955 1674 1007 1678
rect 1011 1674 1031 1678
rect 1035 1674 1063 1678
rect 1067 1674 1103 1678
rect 1107 1674 1119 1678
rect 1123 1674 1175 1678
rect 1179 1674 1231 1678
rect 1235 1674 1247 1678
rect 1251 1674 1287 1678
rect 1291 1674 1319 1678
rect 1323 1674 1335 1678
rect 1339 1674 1375 1678
rect 1379 1674 1391 1678
rect 1395 1674 1423 1678
rect 1427 1674 1455 1678
rect 1459 1674 1471 1678
rect 1475 1674 1519 1678
rect 1523 1674 1583 1678
rect 1587 1674 1623 1678
rect 1627 1674 1663 1678
rect 1667 1674 1687 1678
rect 91 1673 1687 1674
rect 1693 1673 1694 1679
rect 96 1633 97 1639
rect 103 1638 1699 1639
rect 103 1634 111 1638
rect 115 1634 135 1638
rect 139 1634 167 1638
rect 171 1634 183 1638
rect 187 1634 215 1638
rect 219 1634 247 1638
rect 251 1634 279 1638
rect 283 1634 303 1638
rect 307 1634 343 1638
rect 347 1634 359 1638
rect 363 1634 415 1638
rect 419 1634 471 1638
rect 475 1634 487 1638
rect 491 1634 535 1638
rect 539 1634 559 1638
rect 563 1634 599 1638
rect 603 1634 631 1638
rect 635 1634 663 1638
rect 667 1634 711 1638
rect 715 1634 727 1638
rect 731 1634 791 1638
rect 795 1634 799 1638
rect 803 1634 871 1638
rect 875 1634 943 1638
rect 947 1634 951 1638
rect 955 1634 1023 1638
rect 1027 1634 1031 1638
rect 1035 1634 1103 1638
rect 1107 1634 1175 1638
rect 1179 1634 1247 1638
rect 1251 1634 1319 1638
rect 1323 1634 1391 1638
rect 1395 1634 1399 1638
rect 1403 1634 1455 1638
rect 1459 1634 1479 1638
rect 1483 1634 1519 1638
rect 1523 1634 1559 1638
rect 1563 1634 1583 1638
rect 1587 1634 1623 1638
rect 1627 1634 1663 1638
rect 1667 1634 1699 1638
rect 103 1633 1699 1634
rect 1705 1633 1706 1639
rect 84 1593 85 1599
rect 91 1598 1687 1599
rect 91 1594 111 1598
rect 115 1594 135 1598
rect 139 1594 167 1598
rect 171 1594 183 1598
rect 187 1594 223 1598
rect 227 1594 247 1598
rect 251 1594 279 1598
rect 283 1594 303 1598
rect 307 1594 335 1598
rect 339 1594 359 1598
rect 363 1594 383 1598
rect 387 1594 415 1598
rect 419 1594 431 1598
rect 435 1594 471 1598
rect 475 1594 479 1598
rect 483 1594 535 1598
rect 539 1594 599 1598
rect 603 1594 663 1598
rect 667 1594 727 1598
rect 731 1594 799 1598
rect 803 1594 871 1598
rect 875 1594 943 1598
rect 947 1594 951 1598
rect 955 1594 1023 1598
rect 1027 1594 1039 1598
rect 1043 1594 1103 1598
rect 1107 1594 1119 1598
rect 1123 1594 1175 1598
rect 1179 1594 1199 1598
rect 1203 1594 1247 1598
rect 1251 1594 1279 1598
rect 1283 1594 1319 1598
rect 1323 1594 1351 1598
rect 1355 1594 1399 1598
rect 1403 1594 1415 1598
rect 1419 1594 1471 1598
rect 1475 1594 1479 1598
rect 1483 1594 1527 1598
rect 1531 1594 1559 1598
rect 1563 1594 1583 1598
rect 1587 1594 1623 1598
rect 1627 1594 1663 1598
rect 1667 1594 1687 1598
rect 91 1593 1687 1594
rect 1693 1593 1694 1599
rect 96 1553 97 1559
rect 103 1558 1699 1559
rect 103 1554 111 1558
rect 115 1554 135 1558
rect 139 1554 167 1558
rect 171 1554 215 1558
rect 219 1554 223 1558
rect 227 1554 263 1558
rect 267 1554 279 1558
rect 283 1554 311 1558
rect 315 1554 335 1558
rect 339 1554 359 1558
rect 363 1554 383 1558
rect 387 1554 407 1558
rect 411 1554 431 1558
rect 435 1554 455 1558
rect 459 1554 479 1558
rect 483 1554 511 1558
rect 515 1554 535 1558
rect 539 1554 567 1558
rect 571 1554 599 1558
rect 603 1554 631 1558
rect 635 1554 663 1558
rect 667 1554 695 1558
rect 699 1554 727 1558
rect 731 1554 759 1558
rect 763 1554 799 1558
rect 803 1554 831 1558
rect 835 1554 871 1558
rect 875 1554 919 1558
rect 923 1554 951 1558
rect 955 1554 1007 1558
rect 1011 1554 1039 1558
rect 1043 1554 1095 1558
rect 1099 1554 1119 1558
rect 1123 1554 1183 1558
rect 1187 1554 1199 1558
rect 1203 1554 1263 1558
rect 1267 1554 1279 1558
rect 1283 1554 1335 1558
rect 1339 1554 1351 1558
rect 1355 1554 1407 1558
rect 1411 1554 1415 1558
rect 1419 1554 1471 1558
rect 1475 1554 1527 1558
rect 1531 1554 1583 1558
rect 1587 1554 1623 1558
rect 1627 1554 1663 1558
rect 1667 1554 1699 1558
rect 103 1553 1699 1554
rect 1705 1553 1706 1559
rect 84 1509 85 1515
rect 91 1514 1687 1515
rect 91 1510 111 1514
rect 115 1510 135 1514
rect 139 1510 167 1514
rect 171 1510 215 1514
rect 219 1510 223 1514
rect 227 1510 263 1514
rect 267 1510 295 1514
rect 299 1510 311 1514
rect 315 1510 359 1514
rect 363 1510 375 1514
rect 379 1510 407 1514
rect 411 1510 455 1514
rect 459 1510 511 1514
rect 515 1510 527 1514
rect 531 1510 567 1514
rect 571 1510 599 1514
rect 603 1510 631 1514
rect 635 1510 671 1514
rect 675 1510 695 1514
rect 699 1510 743 1514
rect 747 1510 759 1514
rect 763 1510 815 1514
rect 819 1510 831 1514
rect 835 1510 879 1514
rect 883 1510 919 1514
rect 923 1510 943 1514
rect 947 1510 1007 1514
rect 1011 1510 1063 1514
rect 1067 1510 1095 1514
rect 1099 1510 1111 1514
rect 1115 1510 1151 1514
rect 1155 1510 1183 1514
rect 1187 1510 1215 1514
rect 1219 1510 1255 1514
rect 1259 1510 1263 1514
rect 1267 1510 1295 1514
rect 1299 1510 1335 1514
rect 1339 1510 1351 1514
rect 1355 1510 1407 1514
rect 1411 1510 1415 1514
rect 1419 1510 1471 1514
rect 1475 1510 1487 1514
rect 1491 1510 1527 1514
rect 1531 1510 1567 1514
rect 1571 1510 1583 1514
rect 1587 1510 1623 1514
rect 1627 1510 1663 1514
rect 1667 1510 1687 1514
rect 91 1509 1687 1510
rect 1693 1509 1694 1515
rect 96 1469 97 1475
rect 103 1474 1699 1475
rect 103 1470 111 1474
rect 115 1470 135 1474
rect 139 1470 167 1474
rect 171 1470 223 1474
rect 227 1470 295 1474
rect 299 1470 375 1474
rect 379 1470 455 1474
rect 459 1470 527 1474
rect 531 1470 599 1474
rect 603 1470 663 1474
rect 667 1470 671 1474
rect 675 1470 719 1474
rect 723 1470 743 1474
rect 747 1470 783 1474
rect 787 1470 815 1474
rect 819 1470 847 1474
rect 851 1470 879 1474
rect 883 1470 903 1474
rect 907 1470 943 1474
rect 947 1470 959 1474
rect 963 1470 1007 1474
rect 1011 1470 1015 1474
rect 1019 1470 1063 1474
rect 1067 1470 1071 1474
rect 1075 1470 1111 1474
rect 1115 1470 1119 1474
rect 1123 1470 1151 1474
rect 1155 1470 1159 1474
rect 1163 1470 1183 1474
rect 1187 1470 1207 1474
rect 1211 1470 1215 1474
rect 1219 1470 1255 1474
rect 1259 1470 1263 1474
rect 1267 1470 1295 1474
rect 1299 1470 1327 1474
rect 1331 1470 1351 1474
rect 1355 1470 1399 1474
rect 1403 1470 1415 1474
rect 1419 1470 1479 1474
rect 1483 1470 1487 1474
rect 1491 1470 1559 1474
rect 1563 1470 1567 1474
rect 1571 1470 1623 1474
rect 1627 1470 1663 1474
rect 1667 1470 1699 1474
rect 103 1469 1699 1470
rect 1705 1469 1706 1475
rect 84 1425 85 1431
rect 91 1430 1687 1431
rect 91 1426 111 1430
rect 115 1426 135 1430
rect 139 1426 167 1430
rect 171 1426 215 1430
rect 219 1426 223 1430
rect 227 1426 287 1430
rect 291 1426 295 1430
rect 299 1426 359 1430
rect 363 1426 375 1430
rect 379 1426 439 1430
rect 443 1426 455 1430
rect 459 1426 519 1430
rect 523 1426 527 1430
rect 531 1426 599 1430
rect 603 1426 663 1430
rect 667 1426 679 1430
rect 683 1426 719 1430
rect 723 1426 759 1430
rect 763 1426 783 1430
rect 787 1426 831 1430
rect 835 1426 847 1430
rect 851 1426 903 1430
rect 907 1426 959 1430
rect 963 1426 967 1430
rect 971 1426 1015 1430
rect 1019 1426 1031 1430
rect 1035 1426 1071 1430
rect 1075 1426 1103 1430
rect 1107 1426 1119 1430
rect 1123 1426 1159 1430
rect 1163 1426 1167 1430
rect 1171 1426 1207 1430
rect 1211 1426 1231 1430
rect 1235 1426 1263 1430
rect 1267 1426 1295 1430
rect 1299 1426 1327 1430
rect 1331 1426 1359 1430
rect 1363 1426 1399 1430
rect 1403 1426 1415 1430
rect 1419 1426 1463 1430
rect 1467 1426 1479 1430
rect 1483 1426 1503 1430
rect 1507 1426 1551 1430
rect 1555 1426 1559 1430
rect 1563 1426 1591 1430
rect 1595 1426 1623 1430
rect 1627 1426 1663 1430
rect 1667 1426 1687 1430
rect 91 1425 1687 1426
rect 1693 1425 1694 1431
rect 96 1385 97 1391
rect 103 1390 1699 1391
rect 103 1386 111 1390
rect 115 1386 135 1390
rect 139 1386 167 1390
rect 171 1386 215 1390
rect 219 1386 223 1390
rect 227 1386 287 1390
rect 291 1386 359 1390
rect 363 1386 431 1390
rect 435 1386 439 1390
rect 443 1386 503 1390
rect 507 1386 519 1390
rect 523 1386 583 1390
rect 587 1386 599 1390
rect 603 1386 663 1390
rect 667 1386 679 1390
rect 683 1386 743 1390
rect 747 1386 759 1390
rect 763 1386 815 1390
rect 819 1386 831 1390
rect 835 1386 887 1390
rect 891 1386 903 1390
rect 907 1386 959 1390
rect 963 1386 967 1390
rect 971 1386 1031 1390
rect 1035 1386 1103 1390
rect 1107 1386 1167 1390
rect 1171 1386 1175 1390
rect 1179 1386 1231 1390
rect 1235 1386 1239 1390
rect 1243 1386 1295 1390
rect 1299 1386 1303 1390
rect 1307 1386 1359 1390
rect 1363 1386 1367 1390
rect 1371 1386 1415 1390
rect 1419 1386 1431 1390
rect 1435 1386 1463 1390
rect 1467 1386 1495 1390
rect 1499 1386 1503 1390
rect 1507 1386 1551 1390
rect 1555 1386 1567 1390
rect 1571 1386 1591 1390
rect 1595 1386 1623 1390
rect 1627 1386 1663 1390
rect 1667 1386 1699 1390
rect 103 1385 1699 1386
rect 1705 1385 1706 1391
rect 84 1345 85 1351
rect 91 1350 1687 1351
rect 91 1346 111 1350
rect 115 1346 135 1350
rect 139 1346 167 1350
rect 171 1346 183 1350
rect 187 1346 223 1350
rect 227 1346 239 1350
rect 243 1346 287 1350
rect 291 1346 295 1350
rect 299 1346 351 1350
rect 355 1346 359 1350
rect 363 1346 399 1350
rect 403 1346 431 1350
rect 435 1346 455 1350
rect 459 1346 503 1350
rect 507 1346 511 1350
rect 515 1346 567 1350
rect 571 1346 583 1350
rect 587 1346 631 1350
rect 635 1346 663 1350
rect 667 1346 695 1350
rect 699 1346 743 1350
rect 747 1346 759 1350
rect 763 1346 815 1350
rect 819 1346 823 1350
rect 827 1346 887 1350
rect 891 1346 959 1350
rect 963 1346 1023 1350
rect 1027 1346 1031 1350
rect 1035 1346 1087 1350
rect 1091 1346 1103 1350
rect 1107 1346 1151 1350
rect 1155 1346 1175 1350
rect 1179 1346 1215 1350
rect 1219 1346 1239 1350
rect 1243 1346 1279 1350
rect 1283 1346 1303 1350
rect 1307 1346 1343 1350
rect 1347 1346 1367 1350
rect 1371 1346 1407 1350
rect 1411 1346 1431 1350
rect 1435 1346 1479 1350
rect 1483 1346 1495 1350
rect 1499 1346 1559 1350
rect 1563 1346 1567 1350
rect 1571 1346 1623 1350
rect 1627 1346 1663 1350
rect 1667 1346 1687 1350
rect 91 1345 1687 1346
rect 1693 1345 1694 1351
rect 96 1301 97 1307
rect 103 1306 1699 1307
rect 103 1302 111 1306
rect 115 1302 135 1306
rect 139 1302 183 1306
rect 187 1302 231 1306
rect 235 1302 239 1306
rect 243 1302 279 1306
rect 283 1302 295 1306
rect 299 1302 327 1306
rect 331 1302 351 1306
rect 355 1302 375 1306
rect 379 1302 399 1306
rect 403 1302 431 1306
rect 435 1302 455 1306
rect 459 1302 487 1306
rect 491 1302 511 1306
rect 515 1302 543 1306
rect 547 1302 567 1306
rect 571 1302 607 1306
rect 611 1302 631 1306
rect 635 1302 663 1306
rect 667 1302 695 1306
rect 699 1302 719 1306
rect 723 1302 759 1306
rect 763 1302 775 1306
rect 779 1302 823 1306
rect 827 1302 831 1306
rect 835 1302 887 1306
rect 891 1302 895 1306
rect 899 1302 959 1306
rect 963 1302 1023 1306
rect 1027 1302 1079 1306
rect 1083 1302 1087 1306
rect 1091 1302 1143 1306
rect 1147 1302 1151 1306
rect 1155 1302 1207 1306
rect 1211 1302 1215 1306
rect 1219 1302 1279 1306
rect 1283 1302 1343 1306
rect 1347 1302 1359 1306
rect 1363 1302 1407 1306
rect 1411 1302 1447 1306
rect 1451 1302 1479 1306
rect 1483 1302 1543 1306
rect 1547 1302 1559 1306
rect 1563 1302 1623 1306
rect 1627 1302 1663 1306
rect 1667 1302 1699 1306
rect 103 1301 1699 1302
rect 1705 1301 1706 1307
rect 84 1261 85 1267
rect 91 1266 1687 1267
rect 91 1262 111 1266
rect 115 1262 135 1266
rect 139 1262 167 1266
rect 171 1262 183 1266
rect 187 1262 223 1266
rect 227 1262 231 1266
rect 235 1262 279 1266
rect 283 1262 327 1266
rect 331 1262 375 1266
rect 379 1262 383 1266
rect 387 1262 431 1266
rect 435 1262 439 1266
rect 443 1262 487 1266
rect 491 1262 495 1266
rect 499 1262 543 1266
rect 547 1262 551 1266
rect 555 1262 607 1266
rect 611 1262 663 1266
rect 667 1262 719 1266
rect 723 1262 767 1266
rect 771 1262 775 1266
rect 779 1262 815 1266
rect 819 1262 831 1266
rect 835 1262 871 1266
rect 875 1262 895 1266
rect 899 1262 927 1266
rect 931 1262 959 1266
rect 963 1262 983 1266
rect 987 1262 1023 1266
rect 1027 1262 1039 1266
rect 1043 1262 1079 1266
rect 1083 1262 1095 1266
rect 1099 1262 1143 1266
rect 1147 1262 1159 1266
rect 1163 1262 1207 1266
rect 1211 1262 1231 1266
rect 1235 1262 1279 1266
rect 1283 1262 1319 1266
rect 1323 1262 1359 1266
rect 1363 1262 1423 1266
rect 1427 1262 1447 1266
rect 1451 1262 1535 1266
rect 1539 1262 1543 1266
rect 1547 1262 1623 1266
rect 1627 1262 1663 1266
rect 1667 1262 1687 1266
rect 91 1261 1687 1262
rect 1693 1261 1694 1267
rect 96 1217 97 1223
rect 103 1222 1699 1223
rect 103 1218 111 1222
rect 115 1218 135 1222
rect 139 1218 167 1222
rect 171 1218 223 1222
rect 227 1218 279 1222
rect 283 1218 327 1222
rect 331 1218 335 1222
rect 339 1218 383 1222
rect 387 1218 431 1222
rect 435 1218 439 1222
rect 443 1218 487 1222
rect 491 1218 495 1222
rect 499 1218 543 1222
rect 547 1218 551 1222
rect 555 1218 599 1222
rect 603 1218 607 1222
rect 611 1218 655 1222
rect 659 1218 663 1222
rect 667 1218 711 1222
rect 715 1218 719 1222
rect 723 1218 767 1222
rect 771 1218 815 1222
rect 819 1218 823 1222
rect 827 1218 871 1222
rect 875 1218 887 1222
rect 891 1218 927 1222
rect 931 1218 951 1222
rect 955 1218 983 1222
rect 987 1218 1015 1222
rect 1019 1218 1039 1222
rect 1043 1218 1079 1222
rect 1083 1218 1095 1222
rect 1099 1218 1143 1222
rect 1147 1218 1159 1222
rect 1163 1218 1207 1222
rect 1211 1218 1231 1222
rect 1235 1218 1279 1222
rect 1283 1218 1319 1222
rect 1323 1218 1359 1222
rect 1363 1218 1423 1222
rect 1427 1218 1447 1222
rect 1451 1218 1535 1222
rect 1539 1218 1543 1222
rect 1547 1218 1623 1222
rect 1627 1218 1663 1222
rect 1667 1218 1699 1222
rect 103 1217 1699 1218
rect 1705 1217 1706 1223
rect 84 1173 85 1179
rect 91 1178 1687 1179
rect 91 1174 111 1178
rect 115 1174 135 1178
rect 139 1174 167 1178
rect 171 1174 223 1178
rect 227 1174 279 1178
rect 283 1174 287 1178
rect 291 1174 335 1178
rect 339 1174 351 1178
rect 355 1174 383 1178
rect 387 1174 415 1178
rect 419 1174 431 1178
rect 435 1174 471 1178
rect 475 1174 487 1178
rect 491 1174 535 1178
rect 539 1174 543 1178
rect 547 1174 599 1178
rect 603 1174 655 1178
rect 659 1174 663 1178
rect 667 1174 711 1178
rect 715 1174 727 1178
rect 731 1174 767 1178
rect 771 1174 783 1178
rect 787 1174 823 1178
rect 827 1174 839 1178
rect 843 1174 887 1178
rect 891 1174 903 1178
rect 907 1174 951 1178
rect 955 1174 967 1178
rect 971 1174 1015 1178
rect 1019 1174 1031 1178
rect 1035 1174 1079 1178
rect 1083 1174 1095 1178
rect 1099 1174 1143 1178
rect 1147 1174 1159 1178
rect 1163 1174 1207 1178
rect 1211 1174 1215 1178
rect 1219 1174 1279 1178
rect 1283 1174 1343 1178
rect 1347 1174 1359 1178
rect 1363 1174 1407 1178
rect 1411 1174 1447 1178
rect 1451 1174 1479 1178
rect 1483 1174 1543 1178
rect 1547 1174 1559 1178
rect 1563 1174 1623 1178
rect 1627 1174 1663 1178
rect 1667 1174 1687 1178
rect 91 1173 1687 1174
rect 1693 1173 1694 1179
rect 96 1129 97 1135
rect 103 1134 1699 1135
rect 103 1130 111 1134
rect 115 1130 135 1134
rect 139 1130 143 1134
rect 147 1130 167 1134
rect 171 1130 175 1134
rect 179 1130 215 1134
rect 219 1130 223 1134
rect 227 1130 271 1134
rect 275 1130 287 1134
rect 291 1130 335 1134
rect 339 1130 351 1134
rect 355 1130 399 1134
rect 403 1130 415 1134
rect 419 1130 463 1134
rect 467 1130 471 1134
rect 475 1130 527 1134
rect 531 1130 535 1134
rect 539 1130 599 1134
rect 603 1130 663 1134
rect 667 1130 727 1134
rect 731 1130 783 1134
rect 787 1130 791 1134
rect 795 1130 839 1134
rect 843 1130 855 1134
rect 859 1130 903 1134
rect 907 1130 911 1134
rect 915 1130 967 1134
rect 971 1130 1023 1134
rect 1027 1130 1031 1134
rect 1035 1130 1087 1134
rect 1091 1130 1095 1134
rect 1099 1130 1151 1134
rect 1155 1130 1159 1134
rect 1163 1130 1215 1134
rect 1219 1130 1279 1134
rect 1283 1130 1335 1134
rect 1339 1130 1343 1134
rect 1347 1130 1391 1134
rect 1395 1130 1407 1134
rect 1411 1130 1447 1134
rect 1451 1130 1479 1134
rect 1483 1130 1495 1134
rect 1499 1130 1543 1134
rect 1547 1130 1559 1134
rect 1563 1130 1591 1134
rect 1595 1130 1623 1134
rect 1627 1130 1663 1134
rect 1667 1130 1699 1134
rect 103 1129 1699 1130
rect 1705 1129 1706 1135
rect 84 1085 85 1091
rect 91 1090 1687 1091
rect 91 1086 111 1090
rect 115 1086 143 1090
rect 147 1086 175 1090
rect 179 1086 215 1090
rect 219 1086 247 1090
rect 251 1086 271 1090
rect 275 1086 279 1090
rect 283 1086 311 1090
rect 315 1086 335 1090
rect 339 1086 351 1090
rect 355 1086 391 1090
rect 395 1086 399 1090
rect 403 1086 439 1090
rect 443 1086 463 1090
rect 467 1086 503 1090
rect 507 1086 527 1090
rect 531 1086 575 1090
rect 579 1086 599 1090
rect 603 1086 655 1090
rect 659 1086 663 1090
rect 667 1086 727 1090
rect 731 1086 735 1090
rect 739 1086 791 1090
rect 795 1086 815 1090
rect 819 1086 855 1090
rect 859 1086 895 1090
rect 899 1086 911 1090
rect 915 1086 967 1090
rect 971 1086 1023 1090
rect 1027 1086 1039 1090
rect 1043 1086 1087 1090
rect 1091 1086 1111 1090
rect 1115 1086 1151 1090
rect 1155 1086 1175 1090
rect 1179 1086 1215 1090
rect 1219 1086 1239 1090
rect 1243 1086 1279 1090
rect 1283 1086 1303 1090
rect 1307 1086 1335 1090
rect 1339 1086 1359 1090
rect 1363 1086 1391 1090
rect 1395 1086 1415 1090
rect 1419 1086 1447 1090
rect 1451 1086 1463 1090
rect 1467 1086 1495 1090
rect 1499 1086 1503 1090
rect 1507 1086 1543 1090
rect 1547 1086 1551 1090
rect 1555 1086 1591 1090
rect 1595 1086 1623 1090
rect 1627 1086 1663 1090
rect 1667 1086 1687 1090
rect 91 1085 1687 1086
rect 1693 1085 1694 1091
rect 96 1041 97 1047
rect 103 1046 1699 1047
rect 103 1042 111 1046
rect 115 1042 215 1046
rect 219 1042 247 1046
rect 251 1042 279 1046
rect 283 1042 295 1046
rect 299 1042 311 1046
rect 315 1042 327 1046
rect 331 1042 351 1046
rect 355 1042 359 1046
rect 363 1042 391 1046
rect 395 1042 423 1046
rect 427 1042 439 1046
rect 443 1042 455 1046
rect 459 1042 503 1046
rect 507 1042 559 1046
rect 563 1042 575 1046
rect 579 1042 631 1046
rect 635 1042 655 1046
rect 659 1042 711 1046
rect 715 1042 735 1046
rect 739 1042 799 1046
rect 803 1042 815 1046
rect 819 1042 879 1046
rect 883 1042 895 1046
rect 899 1042 959 1046
rect 963 1042 967 1046
rect 971 1042 1031 1046
rect 1035 1042 1039 1046
rect 1043 1042 1095 1046
rect 1099 1042 1111 1046
rect 1115 1042 1159 1046
rect 1163 1042 1175 1046
rect 1179 1042 1223 1046
rect 1227 1042 1239 1046
rect 1243 1042 1279 1046
rect 1283 1042 1303 1046
rect 1307 1042 1335 1046
rect 1339 1042 1359 1046
rect 1363 1042 1383 1046
rect 1387 1042 1415 1046
rect 1419 1042 1431 1046
rect 1435 1042 1463 1046
rect 1467 1042 1479 1046
rect 1483 1042 1503 1046
rect 1507 1042 1535 1046
rect 1539 1042 1551 1046
rect 1555 1042 1591 1046
rect 1595 1042 1623 1046
rect 1627 1042 1663 1046
rect 1667 1042 1699 1046
rect 103 1041 1699 1042
rect 1705 1041 1706 1047
rect 84 1001 85 1007
rect 91 1006 1687 1007
rect 91 1002 111 1006
rect 115 1002 247 1006
rect 251 1002 279 1006
rect 283 1002 295 1006
rect 299 1002 311 1006
rect 315 1002 327 1006
rect 331 1002 343 1006
rect 347 1002 359 1006
rect 363 1002 383 1006
rect 387 1002 391 1006
rect 395 1002 423 1006
rect 427 1002 455 1006
rect 459 1002 479 1006
rect 483 1002 503 1006
rect 507 1002 543 1006
rect 547 1002 559 1006
rect 563 1002 615 1006
rect 619 1002 631 1006
rect 635 1002 687 1006
rect 691 1002 711 1006
rect 715 1002 759 1006
rect 763 1002 799 1006
rect 803 1002 831 1006
rect 835 1002 879 1006
rect 883 1002 903 1006
rect 907 1002 959 1006
rect 963 1002 967 1006
rect 971 1002 1031 1006
rect 1035 1002 1095 1006
rect 1099 1002 1159 1006
rect 1163 1002 1223 1006
rect 1227 1002 1279 1006
rect 1283 1002 1287 1006
rect 1291 1002 1335 1006
rect 1339 1002 1343 1006
rect 1347 1002 1383 1006
rect 1387 1002 1399 1006
rect 1403 1002 1431 1006
rect 1435 1002 1447 1006
rect 1451 1002 1479 1006
rect 1483 1002 1495 1006
rect 1499 1002 1535 1006
rect 1539 1002 1543 1006
rect 1547 1002 1591 1006
rect 1595 1002 1623 1006
rect 1627 1002 1663 1006
rect 1667 1002 1687 1006
rect 91 1001 1687 1002
rect 1693 1001 1694 1007
rect 96 961 97 967
rect 103 966 1699 967
rect 103 962 111 966
rect 115 962 167 966
rect 171 962 199 966
rect 203 962 239 966
rect 243 962 247 966
rect 251 962 279 966
rect 283 962 287 966
rect 291 962 311 966
rect 315 962 343 966
rect 347 962 383 966
rect 387 962 407 966
rect 411 962 423 966
rect 427 962 471 966
rect 475 962 479 966
rect 483 962 535 966
rect 539 962 543 966
rect 547 962 599 966
rect 603 962 615 966
rect 619 962 663 966
rect 667 962 687 966
rect 691 962 727 966
rect 731 962 759 966
rect 763 962 791 966
rect 795 962 831 966
rect 835 962 847 966
rect 851 962 903 966
rect 907 962 911 966
rect 915 962 967 966
rect 971 962 975 966
rect 979 962 1031 966
rect 1035 962 1039 966
rect 1043 962 1095 966
rect 1099 962 1103 966
rect 1107 962 1159 966
rect 1163 962 1167 966
rect 1171 962 1223 966
rect 1227 962 1231 966
rect 1235 962 1287 966
rect 1291 962 1343 966
rect 1347 962 1391 966
rect 1395 962 1399 966
rect 1403 962 1431 966
rect 1435 962 1447 966
rect 1451 962 1471 966
rect 1475 962 1495 966
rect 1499 962 1511 966
rect 1515 962 1543 966
rect 1547 962 1551 966
rect 1555 962 1591 966
rect 1595 962 1623 966
rect 1627 962 1663 966
rect 1667 962 1699 966
rect 103 961 1699 962
rect 1705 961 1706 967
rect 84 917 85 923
rect 91 922 1687 923
rect 91 918 111 922
rect 115 918 135 922
rect 139 918 167 922
rect 171 918 199 922
rect 203 918 207 922
rect 211 918 239 922
rect 243 918 271 922
rect 275 918 287 922
rect 291 918 335 922
rect 339 918 343 922
rect 347 918 407 922
rect 411 918 471 922
rect 475 918 535 922
rect 539 918 591 922
rect 595 918 599 922
rect 603 918 647 922
rect 651 918 663 922
rect 667 918 703 922
rect 707 918 727 922
rect 731 918 751 922
rect 755 918 791 922
rect 795 918 799 922
rect 803 918 847 922
rect 851 918 903 922
rect 907 918 911 922
rect 915 918 959 922
rect 963 918 975 922
rect 979 918 1023 922
rect 1027 918 1039 922
rect 1043 918 1087 922
rect 1091 918 1103 922
rect 1107 918 1143 922
rect 1147 918 1167 922
rect 1171 918 1199 922
rect 1203 918 1231 922
rect 1235 918 1255 922
rect 1259 918 1287 922
rect 1291 918 1319 922
rect 1323 918 1343 922
rect 1347 918 1383 922
rect 1387 918 1391 922
rect 1395 918 1431 922
rect 1435 918 1471 922
rect 1475 918 1511 922
rect 1515 918 1551 922
rect 1555 918 1591 922
rect 1595 918 1623 922
rect 1627 918 1663 922
rect 1667 918 1687 922
rect 91 917 1687 918
rect 1693 917 1694 923
rect 96 873 97 879
rect 103 878 1699 879
rect 103 874 111 878
rect 115 874 135 878
rect 139 874 167 878
rect 171 874 207 878
rect 211 874 271 878
rect 275 874 335 878
rect 339 874 407 878
rect 411 874 471 878
rect 475 874 535 878
rect 539 874 591 878
rect 595 874 599 878
rect 603 874 647 878
rect 651 874 655 878
rect 659 874 703 878
rect 707 874 751 878
rect 755 874 799 878
rect 803 874 847 878
rect 851 874 903 878
rect 907 874 959 878
rect 963 874 967 878
rect 971 874 1023 878
rect 1027 874 1039 878
rect 1043 874 1087 878
rect 1091 874 1103 878
rect 1107 874 1143 878
rect 1147 874 1167 878
rect 1171 874 1199 878
rect 1203 874 1231 878
rect 1235 874 1255 878
rect 1259 874 1287 878
rect 1291 874 1319 878
rect 1323 874 1343 878
rect 1347 874 1383 878
rect 1387 874 1399 878
rect 1403 874 1463 878
rect 1467 874 1663 878
rect 1667 874 1699 878
rect 103 873 1699 874
rect 1705 873 1706 879
rect 84 833 85 839
rect 91 838 1687 839
rect 91 834 111 838
rect 115 834 135 838
rect 139 834 167 838
rect 171 834 207 838
rect 211 834 215 838
rect 219 834 271 838
rect 275 834 279 838
rect 283 834 335 838
rect 339 834 343 838
rect 347 834 407 838
rect 411 834 415 838
rect 419 834 471 838
rect 475 834 479 838
rect 483 834 535 838
rect 539 834 543 838
rect 547 834 599 838
rect 603 834 607 838
rect 611 834 655 838
rect 659 834 671 838
rect 675 834 703 838
rect 707 834 735 838
rect 739 834 751 838
rect 755 834 791 838
rect 795 834 799 838
rect 803 834 847 838
rect 851 834 903 838
rect 907 834 911 838
rect 915 834 967 838
rect 971 834 975 838
rect 979 834 1039 838
rect 1043 834 1103 838
rect 1107 834 1111 838
rect 1115 834 1167 838
rect 1171 834 1183 838
rect 1187 834 1231 838
rect 1235 834 1247 838
rect 1251 834 1287 838
rect 1291 834 1311 838
rect 1315 834 1343 838
rect 1347 834 1367 838
rect 1371 834 1399 838
rect 1403 834 1423 838
rect 1427 834 1463 838
rect 1467 834 1479 838
rect 1483 834 1535 838
rect 1539 834 1591 838
rect 1595 834 1663 838
rect 1667 834 1687 838
rect 91 833 1687 834
rect 1693 833 1694 839
rect 96 789 97 795
rect 103 794 1699 795
rect 103 790 111 794
rect 115 790 135 794
rect 139 790 167 794
rect 171 790 175 794
rect 179 790 215 794
rect 219 790 231 794
rect 235 790 279 794
rect 283 790 295 794
rect 299 790 343 794
rect 347 790 367 794
rect 371 790 415 794
rect 419 790 447 794
rect 451 790 479 794
rect 483 790 527 794
rect 531 790 543 794
rect 547 790 607 794
rect 611 790 615 794
rect 619 790 671 794
rect 675 790 703 794
rect 707 790 735 794
rect 739 790 791 794
rect 795 790 847 794
rect 851 790 871 794
rect 875 790 911 794
rect 915 790 951 794
rect 955 790 975 794
rect 979 790 1023 794
rect 1027 790 1039 794
rect 1043 790 1095 794
rect 1099 790 1111 794
rect 1115 790 1167 794
rect 1171 790 1183 794
rect 1187 790 1231 794
rect 1235 790 1247 794
rect 1251 790 1295 794
rect 1299 790 1311 794
rect 1315 790 1359 794
rect 1363 790 1367 794
rect 1371 790 1415 794
rect 1419 790 1423 794
rect 1427 790 1471 794
rect 1475 790 1479 794
rect 1483 790 1527 794
rect 1531 790 1535 794
rect 1539 790 1591 794
rect 1595 790 1663 794
rect 1667 790 1699 794
rect 103 789 1699 790
rect 1705 789 1706 795
rect 84 749 85 755
rect 91 754 1687 755
rect 91 750 111 754
rect 115 750 135 754
rect 139 750 175 754
rect 179 750 215 754
rect 219 750 231 754
rect 235 750 247 754
rect 251 750 279 754
rect 283 750 295 754
rect 299 750 319 754
rect 323 750 359 754
rect 363 750 367 754
rect 371 750 399 754
rect 403 750 439 754
rect 443 750 447 754
rect 451 750 487 754
rect 491 750 527 754
rect 531 750 543 754
rect 547 750 607 754
rect 611 750 615 754
rect 619 750 671 754
rect 675 750 703 754
rect 707 750 735 754
rect 739 750 791 754
rect 795 750 799 754
rect 803 750 863 754
rect 867 750 871 754
rect 875 750 927 754
rect 931 750 951 754
rect 955 750 991 754
rect 995 750 1023 754
rect 1027 750 1055 754
rect 1059 750 1095 754
rect 1099 750 1119 754
rect 1123 750 1167 754
rect 1171 750 1183 754
rect 1187 750 1231 754
rect 1235 750 1239 754
rect 1243 750 1295 754
rect 1299 750 1351 754
rect 1355 750 1359 754
rect 1363 750 1407 754
rect 1411 750 1415 754
rect 1419 750 1463 754
rect 1467 750 1471 754
rect 1475 750 1519 754
rect 1523 750 1527 754
rect 1531 750 1583 754
rect 1587 750 1591 754
rect 1595 750 1623 754
rect 1627 750 1663 754
rect 1667 750 1687 754
rect 91 749 1687 750
rect 1693 749 1694 755
rect 96 705 97 711
rect 103 710 1699 711
rect 103 706 111 710
rect 115 706 215 710
rect 219 706 247 710
rect 251 706 279 710
rect 283 706 311 710
rect 315 706 319 710
rect 323 706 343 710
rect 347 706 359 710
rect 363 706 375 710
rect 379 706 399 710
rect 403 706 407 710
rect 411 706 439 710
rect 443 706 471 710
rect 475 706 487 710
rect 491 706 503 710
rect 507 706 543 710
rect 547 706 591 710
rect 595 706 607 710
rect 611 706 647 710
rect 651 706 671 710
rect 675 706 703 710
rect 707 706 735 710
rect 739 706 759 710
rect 763 706 799 710
rect 803 706 823 710
rect 827 706 863 710
rect 867 706 887 710
rect 891 706 927 710
rect 931 706 959 710
rect 963 706 991 710
rect 995 706 1023 710
rect 1027 706 1055 710
rect 1059 706 1087 710
rect 1091 706 1119 710
rect 1123 706 1159 710
rect 1163 706 1183 710
rect 1187 706 1223 710
rect 1227 706 1239 710
rect 1243 706 1287 710
rect 1291 706 1295 710
rect 1299 706 1351 710
rect 1355 706 1407 710
rect 1411 706 1415 710
rect 1419 706 1463 710
rect 1467 706 1471 710
rect 1475 706 1519 710
rect 1523 706 1527 710
rect 1531 706 1583 710
rect 1587 706 1623 710
rect 1627 706 1663 710
rect 1667 706 1699 710
rect 103 705 1699 706
rect 1705 705 1706 711
rect 84 665 85 671
rect 91 670 1687 671
rect 91 666 111 670
rect 115 666 279 670
rect 283 666 295 670
rect 299 666 311 670
rect 315 666 327 670
rect 331 666 343 670
rect 347 666 359 670
rect 363 666 375 670
rect 379 666 391 670
rect 395 666 407 670
rect 411 666 423 670
rect 427 666 439 670
rect 443 666 455 670
rect 459 666 471 670
rect 475 666 487 670
rect 491 666 503 670
rect 507 666 519 670
rect 523 666 543 670
rect 547 666 551 670
rect 555 666 591 670
rect 595 666 639 670
rect 643 666 647 670
rect 651 666 687 670
rect 691 666 703 670
rect 707 666 735 670
rect 739 666 759 670
rect 763 666 791 670
rect 795 666 823 670
rect 827 666 847 670
rect 851 666 887 670
rect 891 666 911 670
rect 915 666 959 670
rect 963 666 975 670
rect 979 666 1023 670
rect 1027 666 1047 670
rect 1051 666 1087 670
rect 1091 666 1127 670
rect 1131 666 1159 670
rect 1163 666 1215 670
rect 1219 666 1223 670
rect 1227 666 1287 670
rect 1291 666 1295 670
rect 1299 666 1351 670
rect 1355 666 1383 670
rect 1387 666 1415 670
rect 1419 666 1471 670
rect 1475 666 1527 670
rect 1531 666 1559 670
rect 1563 666 1583 670
rect 1587 666 1623 670
rect 1627 666 1663 670
rect 1667 666 1687 670
rect 91 665 1687 666
rect 1693 665 1694 671
rect 96 625 97 631
rect 103 630 1699 631
rect 103 626 111 630
rect 115 626 247 630
rect 251 626 279 630
rect 283 626 295 630
rect 299 626 319 630
rect 323 626 327 630
rect 331 626 359 630
rect 363 626 367 630
rect 371 626 391 630
rect 395 626 423 630
rect 427 626 455 630
rect 459 626 471 630
rect 475 626 487 630
rect 491 626 519 630
rect 523 626 551 630
rect 555 626 567 630
rect 571 626 591 630
rect 595 626 615 630
rect 619 626 639 630
rect 643 626 663 630
rect 667 626 687 630
rect 691 626 719 630
rect 723 626 735 630
rect 739 626 775 630
rect 779 626 791 630
rect 795 626 831 630
rect 835 626 847 630
rect 851 626 895 630
rect 899 626 911 630
rect 915 626 967 630
rect 971 626 975 630
rect 979 626 1047 630
rect 1051 626 1127 630
rect 1131 626 1207 630
rect 1211 626 1215 630
rect 1219 626 1287 630
rect 1291 626 1295 630
rect 1299 626 1359 630
rect 1363 626 1383 630
rect 1387 626 1431 630
rect 1435 626 1471 630
rect 1475 626 1503 630
rect 1507 626 1559 630
rect 1563 626 1575 630
rect 1579 626 1623 630
rect 1627 626 1663 630
rect 1667 626 1699 630
rect 103 625 1699 626
rect 1705 625 1706 631
rect 84 585 85 591
rect 91 590 1687 591
rect 91 586 111 590
rect 115 586 167 590
rect 171 586 215 590
rect 219 586 247 590
rect 251 586 271 590
rect 275 586 279 590
rect 283 586 319 590
rect 323 586 335 590
rect 339 586 367 590
rect 371 586 407 590
rect 411 586 423 590
rect 427 586 471 590
rect 475 586 487 590
rect 491 586 519 590
rect 523 586 559 590
rect 563 586 567 590
rect 571 586 615 590
rect 619 586 631 590
rect 635 586 663 590
rect 667 586 703 590
rect 707 586 719 590
rect 723 586 767 590
rect 771 586 775 590
rect 779 586 823 590
rect 827 586 831 590
rect 835 586 879 590
rect 883 586 895 590
rect 899 586 935 590
rect 939 586 967 590
rect 971 586 991 590
rect 995 586 1047 590
rect 1051 586 1103 590
rect 1107 586 1127 590
rect 1131 586 1159 590
rect 1163 586 1207 590
rect 1211 586 1215 590
rect 1219 586 1271 590
rect 1275 586 1287 590
rect 1291 586 1327 590
rect 1331 586 1359 590
rect 1363 586 1383 590
rect 1387 586 1431 590
rect 1435 586 1447 590
rect 1451 586 1503 590
rect 1507 586 1511 590
rect 1515 586 1575 590
rect 1579 586 1623 590
rect 1627 586 1663 590
rect 1667 586 1687 590
rect 91 585 1687 586
rect 1693 585 1694 591
rect 96 541 97 547
rect 103 546 1699 547
rect 103 542 111 546
rect 115 542 135 546
rect 139 542 167 546
rect 171 542 199 546
rect 203 542 215 546
rect 219 542 231 546
rect 235 542 271 546
rect 275 542 279 546
rect 283 542 327 546
rect 331 542 335 546
rect 339 542 375 546
rect 379 542 407 546
rect 411 542 431 546
rect 435 542 487 546
rect 491 542 495 546
rect 499 542 559 546
rect 563 542 623 546
rect 627 542 631 546
rect 635 542 687 546
rect 691 542 703 546
rect 707 542 751 546
rect 755 542 767 546
rect 771 542 815 546
rect 819 542 823 546
rect 827 542 879 546
rect 883 542 935 546
rect 939 542 943 546
rect 947 542 991 546
rect 995 542 1007 546
rect 1011 542 1047 546
rect 1051 542 1071 546
rect 1075 542 1103 546
rect 1107 542 1127 546
rect 1131 542 1159 546
rect 1163 542 1183 546
rect 1187 542 1215 546
rect 1219 542 1231 546
rect 1235 542 1271 546
rect 1275 542 1279 546
rect 1283 542 1327 546
rect 1331 542 1335 546
rect 1339 542 1383 546
rect 1387 542 1391 546
rect 1395 542 1447 546
rect 1451 542 1511 546
rect 1515 542 1575 546
rect 1579 542 1623 546
rect 1627 542 1663 546
rect 1667 542 1699 546
rect 103 541 1699 542
rect 1705 541 1706 547
rect 84 501 85 507
rect 91 506 1687 507
rect 91 502 111 506
rect 115 502 135 506
rect 139 502 167 506
rect 171 502 199 506
rect 203 502 231 506
rect 235 502 239 506
rect 243 502 279 506
rect 283 502 287 506
rect 291 502 327 506
rect 331 502 375 506
rect 379 502 423 506
rect 427 502 431 506
rect 435 502 479 506
rect 483 502 495 506
rect 499 502 543 506
rect 547 502 559 506
rect 563 502 615 506
rect 619 502 623 506
rect 627 502 687 506
rect 691 502 695 506
rect 699 502 751 506
rect 755 502 775 506
rect 779 502 815 506
rect 819 502 847 506
rect 851 502 879 506
rect 883 502 919 506
rect 923 502 943 506
rect 947 502 983 506
rect 987 502 1007 506
rect 1011 502 1039 506
rect 1043 502 1071 506
rect 1075 502 1095 506
rect 1099 502 1127 506
rect 1131 502 1143 506
rect 1147 502 1183 506
rect 1187 502 1191 506
rect 1195 502 1231 506
rect 1235 502 1239 506
rect 1243 502 1279 506
rect 1283 502 1287 506
rect 1291 502 1335 506
rect 1339 502 1383 506
rect 1387 502 1391 506
rect 1395 502 1431 506
rect 1435 502 1447 506
rect 1451 502 1479 506
rect 1483 502 1511 506
rect 1515 502 1535 506
rect 1539 502 1575 506
rect 1579 502 1591 506
rect 1595 502 1623 506
rect 1627 502 1663 506
rect 1667 502 1687 506
rect 91 501 1687 502
rect 1693 501 1694 507
rect 96 461 97 467
rect 103 466 1699 467
rect 103 462 111 466
rect 115 462 135 466
rect 139 462 151 466
rect 155 462 167 466
rect 171 462 199 466
rect 203 462 207 466
rect 211 462 239 466
rect 243 462 255 466
rect 259 462 287 466
rect 291 462 311 466
rect 315 462 327 466
rect 331 462 367 466
rect 371 462 375 466
rect 379 462 423 466
rect 427 462 439 466
rect 443 462 479 466
rect 483 462 519 466
rect 523 462 543 466
rect 547 462 599 466
rect 603 462 615 466
rect 619 462 679 466
rect 683 462 695 466
rect 699 462 759 466
rect 763 462 775 466
rect 779 462 839 466
rect 843 462 847 466
rect 851 462 911 466
rect 915 462 919 466
rect 923 462 983 466
rect 987 462 1039 466
rect 1043 462 1055 466
rect 1059 462 1095 466
rect 1099 462 1127 466
rect 1131 462 1143 466
rect 1147 462 1191 466
rect 1195 462 1199 466
rect 1203 462 1239 466
rect 1243 462 1263 466
rect 1267 462 1287 466
rect 1291 462 1319 466
rect 1323 462 1335 466
rect 1339 462 1375 466
rect 1379 462 1383 466
rect 1387 462 1431 466
rect 1435 462 1479 466
rect 1483 462 1495 466
rect 1499 462 1535 466
rect 1539 462 1591 466
rect 1595 462 1623 466
rect 1627 462 1663 466
rect 1667 462 1699 466
rect 103 461 1699 462
rect 1705 461 1706 467
rect 84 421 85 427
rect 91 426 1687 427
rect 91 422 111 426
rect 115 422 151 426
rect 155 422 175 426
rect 179 422 207 426
rect 211 422 223 426
rect 227 422 255 426
rect 259 422 271 426
rect 275 422 311 426
rect 315 422 319 426
rect 323 422 367 426
rect 371 422 415 426
rect 419 422 439 426
rect 443 422 471 426
rect 475 422 519 426
rect 523 422 527 426
rect 531 422 591 426
rect 595 422 599 426
rect 603 422 663 426
rect 667 422 679 426
rect 683 422 735 426
rect 739 422 759 426
rect 763 422 807 426
rect 811 422 839 426
rect 843 422 871 426
rect 875 422 911 426
rect 915 422 935 426
rect 939 422 983 426
rect 987 422 991 426
rect 995 422 1039 426
rect 1043 422 1055 426
rect 1059 422 1087 426
rect 1091 422 1127 426
rect 1131 422 1167 426
rect 1171 422 1199 426
rect 1203 422 1207 426
rect 1211 422 1247 426
rect 1251 422 1263 426
rect 1267 422 1287 426
rect 1291 422 1319 426
rect 1323 422 1335 426
rect 1339 422 1375 426
rect 1379 422 1383 426
rect 1387 422 1431 426
rect 1435 422 1495 426
rect 1499 422 1663 426
rect 1667 422 1687 426
rect 91 421 1687 422
rect 1693 421 1694 427
rect 96 377 97 383
rect 103 382 1699 383
rect 103 378 111 382
rect 115 378 135 382
rect 139 378 167 382
rect 171 378 175 382
rect 179 378 199 382
rect 203 378 223 382
rect 227 378 239 382
rect 243 378 271 382
rect 275 378 295 382
rect 299 378 319 382
rect 323 378 351 382
rect 355 378 367 382
rect 371 378 407 382
rect 411 378 415 382
rect 419 378 463 382
rect 467 378 471 382
rect 475 378 519 382
rect 523 378 527 382
rect 531 378 575 382
rect 579 378 591 382
rect 595 378 631 382
rect 635 378 663 382
rect 667 378 687 382
rect 691 378 735 382
rect 739 378 743 382
rect 747 378 799 382
rect 803 378 807 382
rect 811 378 855 382
rect 859 378 871 382
rect 875 378 919 382
rect 923 378 935 382
rect 939 378 983 382
rect 987 378 991 382
rect 995 378 1039 382
rect 1043 378 1087 382
rect 1091 378 1095 382
rect 1099 378 1127 382
rect 1131 378 1151 382
rect 1155 378 1167 382
rect 1171 378 1207 382
rect 1211 378 1247 382
rect 1251 378 1255 382
rect 1259 378 1287 382
rect 1291 378 1303 382
rect 1307 378 1335 382
rect 1339 378 1351 382
rect 1355 378 1383 382
rect 1387 378 1399 382
rect 1403 378 1447 382
rect 1451 378 1495 382
rect 1499 378 1543 382
rect 1547 378 1591 382
rect 1595 378 1623 382
rect 1627 378 1663 382
rect 1667 378 1699 382
rect 103 377 1699 378
rect 1705 377 1706 383
rect 84 337 85 343
rect 91 342 1687 343
rect 91 338 111 342
rect 115 338 135 342
rect 139 338 167 342
rect 171 338 199 342
rect 203 338 207 342
rect 211 338 239 342
rect 243 338 263 342
rect 267 338 295 342
rect 299 338 327 342
rect 331 338 351 342
rect 355 338 391 342
rect 395 338 407 342
rect 411 338 455 342
rect 459 338 463 342
rect 467 338 519 342
rect 523 338 575 342
rect 579 338 631 342
rect 635 338 687 342
rect 691 338 743 342
rect 747 338 751 342
rect 755 338 799 342
rect 803 338 815 342
rect 819 338 855 342
rect 859 338 879 342
rect 883 338 919 342
rect 923 338 951 342
rect 955 338 983 342
rect 987 338 1031 342
rect 1035 338 1039 342
rect 1043 338 1095 342
rect 1099 338 1111 342
rect 1115 338 1151 342
rect 1155 338 1191 342
rect 1195 338 1207 342
rect 1211 338 1255 342
rect 1259 338 1271 342
rect 1275 338 1303 342
rect 1307 338 1343 342
rect 1347 338 1351 342
rect 1355 338 1399 342
rect 1403 338 1407 342
rect 1411 338 1447 342
rect 1451 338 1463 342
rect 1467 338 1495 342
rect 1499 338 1519 342
rect 1523 338 1543 342
rect 1547 338 1583 342
rect 1587 338 1591 342
rect 1595 338 1623 342
rect 1627 338 1663 342
rect 1667 338 1687 342
rect 91 337 1687 338
rect 1693 337 1694 343
rect 96 297 97 303
rect 103 302 1699 303
rect 103 298 111 302
rect 115 298 135 302
rect 139 298 167 302
rect 171 298 207 302
rect 211 298 231 302
rect 235 298 263 302
rect 267 298 295 302
rect 299 298 327 302
rect 331 298 367 302
rect 371 298 391 302
rect 395 298 439 302
rect 443 298 455 302
rect 459 298 503 302
rect 507 298 519 302
rect 523 298 567 302
rect 571 298 575 302
rect 579 298 631 302
rect 635 298 687 302
rect 691 298 743 302
rect 747 298 751 302
rect 755 298 807 302
rect 811 298 815 302
rect 819 298 879 302
rect 883 298 951 302
rect 955 298 1031 302
rect 1035 298 1111 302
rect 1115 298 1191 302
rect 1195 298 1263 302
rect 1267 298 1271 302
rect 1275 298 1327 302
rect 1331 298 1343 302
rect 1347 298 1391 302
rect 1395 298 1407 302
rect 1411 298 1447 302
rect 1451 298 1463 302
rect 1467 298 1495 302
rect 1499 298 1519 302
rect 1523 298 1543 302
rect 1547 298 1583 302
rect 1587 298 1591 302
rect 1595 298 1623 302
rect 1627 298 1663 302
rect 1667 298 1699 302
rect 103 297 1699 298
rect 1705 297 1706 303
rect 84 253 85 259
rect 91 258 1687 259
rect 91 254 111 258
rect 115 254 135 258
rect 139 254 167 258
rect 171 254 175 258
rect 179 254 231 258
rect 235 254 247 258
rect 251 254 295 258
rect 299 254 319 258
rect 323 254 367 258
rect 371 254 383 258
rect 387 254 439 258
rect 443 254 447 258
rect 451 254 503 258
rect 507 254 519 258
rect 523 254 567 258
rect 571 254 591 258
rect 595 254 631 258
rect 635 254 663 258
rect 667 254 687 258
rect 691 254 743 258
rect 747 254 807 258
rect 811 254 823 258
rect 827 254 879 258
rect 883 254 895 258
rect 899 254 951 258
rect 955 254 967 258
rect 971 254 1031 258
rect 1035 254 1087 258
rect 1091 254 1111 258
rect 1115 254 1143 258
rect 1147 254 1191 258
rect 1195 254 1199 258
rect 1203 254 1255 258
rect 1259 254 1263 258
rect 1267 254 1311 258
rect 1315 254 1327 258
rect 1331 254 1367 258
rect 1371 254 1391 258
rect 1395 254 1415 258
rect 1419 254 1447 258
rect 1451 254 1463 258
rect 1467 254 1495 258
rect 1499 254 1519 258
rect 1523 254 1543 258
rect 1547 254 1575 258
rect 1579 254 1591 258
rect 1595 254 1623 258
rect 1627 254 1663 258
rect 1667 254 1687 258
rect 91 253 1687 254
rect 1693 253 1694 259
rect 96 213 97 219
rect 103 218 1699 219
rect 103 214 111 218
rect 115 214 135 218
rect 139 214 167 218
rect 171 214 175 218
rect 179 214 207 218
rect 211 214 247 218
rect 251 214 255 218
rect 259 214 303 218
rect 307 214 319 218
rect 323 214 343 218
rect 347 214 375 218
rect 379 214 383 218
rect 387 214 415 218
rect 419 214 447 218
rect 451 214 471 218
rect 475 214 519 218
rect 523 214 535 218
rect 539 214 591 218
rect 595 214 615 218
rect 619 214 663 218
rect 667 214 695 218
rect 699 214 743 218
rect 747 214 775 218
rect 779 214 823 218
rect 827 214 855 218
rect 859 214 895 218
rect 899 214 927 218
rect 931 214 967 218
rect 971 214 999 218
rect 1003 214 1031 218
rect 1035 214 1071 218
rect 1075 214 1087 218
rect 1091 214 1143 218
rect 1147 214 1199 218
rect 1203 214 1215 218
rect 1219 214 1255 218
rect 1259 214 1287 218
rect 1291 214 1311 218
rect 1315 214 1351 218
rect 1355 214 1367 218
rect 1371 214 1415 218
rect 1419 214 1463 218
rect 1467 214 1471 218
rect 1475 214 1519 218
rect 1523 214 1527 218
rect 1531 214 1575 218
rect 1579 214 1583 218
rect 1587 214 1623 218
rect 1627 214 1663 218
rect 1667 214 1699 218
rect 103 213 1699 214
rect 1705 213 1706 219
rect 84 173 85 179
rect 91 178 1687 179
rect 91 174 111 178
rect 115 174 135 178
rect 139 174 167 178
rect 171 174 175 178
rect 179 174 207 178
rect 211 174 231 178
rect 235 174 255 178
rect 259 174 287 178
rect 291 174 303 178
rect 307 174 343 178
rect 347 174 375 178
rect 379 174 399 178
rect 403 174 415 178
rect 419 174 455 178
rect 459 174 471 178
rect 475 174 511 178
rect 515 174 535 178
rect 539 174 575 178
rect 579 174 615 178
rect 619 174 639 178
rect 643 174 695 178
rect 699 174 703 178
rect 707 174 767 178
rect 771 174 775 178
rect 779 174 831 178
rect 835 174 855 178
rect 859 174 895 178
rect 899 174 927 178
rect 931 174 951 178
rect 955 174 999 178
rect 1003 174 1015 178
rect 1019 174 1071 178
rect 1075 174 1079 178
rect 1083 174 1143 178
rect 1147 174 1207 178
rect 1211 174 1215 178
rect 1219 174 1279 178
rect 1283 174 1287 178
rect 1291 174 1351 178
rect 1355 174 1415 178
rect 1419 174 1423 178
rect 1427 174 1471 178
rect 1475 174 1495 178
rect 1499 174 1527 178
rect 1531 174 1567 178
rect 1571 174 1583 178
rect 1587 174 1623 178
rect 1627 174 1663 178
rect 1667 174 1687 178
rect 91 173 1687 174
rect 1693 173 1694 179
rect 96 117 97 123
rect 103 122 1699 123
rect 103 118 111 122
rect 115 118 135 122
rect 139 118 167 122
rect 171 118 175 122
rect 179 118 199 122
rect 203 118 231 122
rect 235 118 263 122
rect 267 118 287 122
rect 291 118 295 122
rect 299 118 327 122
rect 331 118 343 122
rect 347 118 359 122
rect 363 118 391 122
rect 395 118 399 122
rect 403 118 423 122
rect 427 118 455 122
rect 459 118 463 122
rect 467 118 503 122
rect 507 118 511 122
rect 515 118 543 122
rect 547 118 575 122
rect 579 118 607 122
rect 611 118 639 122
rect 643 118 671 122
rect 675 118 703 122
rect 707 118 735 122
rect 739 118 767 122
rect 771 118 799 122
rect 803 118 831 122
rect 835 118 863 122
rect 867 118 895 122
rect 899 118 935 122
rect 939 118 951 122
rect 955 118 975 122
rect 979 118 1015 122
rect 1019 118 1063 122
rect 1067 118 1079 122
rect 1083 118 1103 122
rect 1107 118 1143 122
rect 1147 118 1183 122
rect 1187 118 1207 122
rect 1211 118 1223 122
rect 1227 118 1263 122
rect 1267 118 1279 122
rect 1283 118 1295 122
rect 1299 118 1335 122
rect 1339 118 1351 122
rect 1355 118 1375 122
rect 1379 118 1415 122
rect 1419 118 1423 122
rect 1427 118 1455 122
rect 1459 118 1495 122
rect 1499 118 1503 122
rect 1507 118 1551 122
rect 1555 118 1567 122
rect 1571 118 1591 122
rect 1595 118 1623 122
rect 1627 118 1663 122
rect 1667 118 1699 122
rect 103 117 1699 118
rect 1705 117 1706 123
rect 84 77 85 83
rect 91 82 1687 83
rect 91 78 111 82
rect 115 78 135 82
rect 139 78 167 82
rect 171 78 199 82
rect 203 78 231 82
rect 235 78 263 82
rect 267 78 295 82
rect 299 78 327 82
rect 331 78 359 82
rect 363 78 391 82
rect 395 78 423 82
rect 427 78 463 82
rect 467 78 503 82
rect 507 78 543 82
rect 547 78 575 82
rect 579 78 607 82
rect 611 78 639 82
rect 643 78 671 82
rect 675 78 703 82
rect 707 78 735 82
rect 739 78 767 82
rect 771 78 799 82
rect 803 78 831 82
rect 835 78 863 82
rect 867 78 895 82
rect 899 78 935 82
rect 939 78 975 82
rect 979 78 1015 82
rect 1019 78 1063 82
rect 1067 78 1103 82
rect 1107 78 1143 82
rect 1147 78 1183 82
rect 1187 78 1223 82
rect 1227 78 1263 82
rect 1267 78 1295 82
rect 1299 78 1335 82
rect 1339 78 1375 82
rect 1379 78 1415 82
rect 1419 78 1455 82
rect 1459 78 1503 82
rect 1507 78 1551 82
rect 1555 78 1591 82
rect 1595 78 1623 82
rect 1627 78 1663 82
rect 1667 78 1687 82
rect 91 77 1687 78
rect 1693 77 1694 83
<< m5c >>
rect 97 1713 103 1719
rect 1699 1713 1705 1719
rect 85 1673 91 1679
rect 1687 1673 1693 1679
rect 97 1633 103 1639
rect 1699 1633 1705 1639
rect 85 1593 91 1599
rect 1687 1593 1693 1599
rect 97 1553 103 1559
rect 1699 1553 1705 1559
rect 85 1509 91 1515
rect 1687 1509 1693 1515
rect 97 1469 103 1475
rect 1699 1469 1705 1475
rect 85 1425 91 1431
rect 1687 1425 1693 1431
rect 97 1385 103 1391
rect 1699 1385 1705 1391
rect 85 1345 91 1351
rect 1687 1345 1693 1351
rect 97 1301 103 1307
rect 1699 1301 1705 1307
rect 85 1261 91 1267
rect 1687 1261 1693 1267
rect 97 1217 103 1223
rect 1699 1217 1705 1223
rect 85 1173 91 1179
rect 1687 1173 1693 1179
rect 97 1129 103 1135
rect 1699 1129 1705 1135
rect 85 1085 91 1091
rect 1687 1085 1693 1091
rect 97 1041 103 1047
rect 1699 1041 1705 1047
rect 85 1001 91 1007
rect 1687 1001 1693 1007
rect 97 961 103 967
rect 1699 961 1705 967
rect 85 917 91 923
rect 1687 917 1693 923
rect 97 873 103 879
rect 1699 873 1705 879
rect 85 833 91 839
rect 1687 833 1693 839
rect 97 789 103 795
rect 1699 789 1705 795
rect 85 749 91 755
rect 1687 749 1693 755
rect 97 705 103 711
rect 1699 705 1705 711
rect 85 665 91 671
rect 1687 665 1693 671
rect 97 625 103 631
rect 1699 625 1705 631
rect 85 585 91 591
rect 1687 585 1693 591
rect 97 541 103 547
rect 1699 541 1705 547
rect 85 501 91 507
rect 1687 501 1693 507
rect 97 461 103 467
rect 1699 461 1705 467
rect 85 421 91 427
rect 1687 421 1693 427
rect 97 377 103 383
rect 1699 377 1705 383
rect 85 337 91 343
rect 1687 337 1693 343
rect 97 297 103 303
rect 1699 297 1705 303
rect 85 253 91 259
rect 1687 253 1693 259
rect 97 213 103 219
rect 1699 213 1705 219
rect 85 173 91 179
rect 1687 173 1693 179
rect 97 117 103 123
rect 1699 117 1705 123
rect 85 77 91 83
rect 1687 77 1693 83
<< m5 >>
rect 84 1679 92 1728
rect 84 1673 85 1679
rect 91 1673 92 1679
rect 84 1599 92 1673
rect 84 1593 85 1599
rect 91 1593 92 1599
rect 84 1515 92 1593
rect 84 1509 85 1515
rect 91 1509 92 1515
rect 84 1431 92 1509
rect 84 1425 85 1431
rect 91 1425 92 1431
rect 84 1351 92 1425
rect 84 1345 85 1351
rect 91 1345 92 1351
rect 84 1267 92 1345
rect 84 1261 85 1267
rect 91 1261 92 1267
rect 84 1179 92 1261
rect 84 1173 85 1179
rect 91 1173 92 1179
rect 84 1091 92 1173
rect 84 1085 85 1091
rect 91 1085 92 1091
rect 84 1007 92 1085
rect 84 1001 85 1007
rect 91 1001 92 1007
rect 84 923 92 1001
rect 84 917 85 923
rect 91 917 92 923
rect 84 839 92 917
rect 84 833 85 839
rect 91 833 92 839
rect 84 755 92 833
rect 84 749 85 755
rect 91 749 92 755
rect 84 671 92 749
rect 84 665 85 671
rect 91 665 92 671
rect 84 591 92 665
rect 84 585 85 591
rect 91 585 92 591
rect 84 507 92 585
rect 84 501 85 507
rect 91 501 92 507
rect 84 427 92 501
rect 84 421 85 427
rect 91 421 92 427
rect 84 343 92 421
rect 84 337 85 343
rect 91 337 92 343
rect 84 259 92 337
rect 84 253 85 259
rect 91 253 92 259
rect 84 179 92 253
rect 84 173 85 179
rect 91 173 92 179
rect 84 83 92 173
rect 84 77 85 83
rect 91 77 92 83
rect 84 72 92 77
rect 96 1719 104 1728
rect 96 1713 97 1719
rect 103 1713 104 1719
rect 96 1639 104 1713
rect 96 1633 97 1639
rect 103 1633 104 1639
rect 96 1559 104 1633
rect 96 1553 97 1559
rect 103 1553 104 1559
rect 96 1475 104 1553
rect 96 1469 97 1475
rect 103 1469 104 1475
rect 96 1391 104 1469
rect 96 1385 97 1391
rect 103 1385 104 1391
rect 96 1307 104 1385
rect 96 1301 97 1307
rect 103 1301 104 1307
rect 96 1223 104 1301
rect 96 1217 97 1223
rect 103 1217 104 1223
rect 96 1135 104 1217
rect 96 1129 97 1135
rect 103 1129 104 1135
rect 96 1047 104 1129
rect 96 1041 97 1047
rect 103 1041 104 1047
rect 96 967 104 1041
rect 96 961 97 967
rect 103 961 104 967
rect 96 879 104 961
rect 96 873 97 879
rect 103 873 104 879
rect 96 795 104 873
rect 96 789 97 795
rect 103 789 104 795
rect 96 711 104 789
rect 96 705 97 711
rect 103 705 104 711
rect 96 631 104 705
rect 96 625 97 631
rect 103 625 104 631
rect 96 547 104 625
rect 96 541 97 547
rect 103 541 104 547
rect 96 467 104 541
rect 96 461 97 467
rect 103 461 104 467
rect 96 383 104 461
rect 96 377 97 383
rect 103 377 104 383
rect 96 303 104 377
rect 96 297 97 303
rect 103 297 104 303
rect 96 219 104 297
rect 96 213 97 219
rect 103 213 104 219
rect 96 123 104 213
rect 96 117 97 123
rect 103 117 104 123
rect 96 72 104 117
rect 1686 1679 1694 1728
rect 1686 1673 1687 1679
rect 1693 1673 1694 1679
rect 1686 1599 1694 1673
rect 1686 1593 1687 1599
rect 1693 1593 1694 1599
rect 1686 1515 1694 1593
rect 1686 1509 1687 1515
rect 1693 1509 1694 1515
rect 1686 1431 1694 1509
rect 1686 1425 1687 1431
rect 1693 1425 1694 1431
rect 1686 1351 1694 1425
rect 1686 1345 1687 1351
rect 1693 1345 1694 1351
rect 1686 1267 1694 1345
rect 1686 1261 1687 1267
rect 1693 1261 1694 1267
rect 1686 1179 1694 1261
rect 1686 1173 1687 1179
rect 1693 1173 1694 1179
rect 1686 1091 1694 1173
rect 1686 1085 1687 1091
rect 1693 1085 1694 1091
rect 1686 1007 1694 1085
rect 1686 1001 1687 1007
rect 1693 1001 1694 1007
rect 1686 923 1694 1001
rect 1686 917 1687 923
rect 1693 917 1694 923
rect 1686 839 1694 917
rect 1686 833 1687 839
rect 1693 833 1694 839
rect 1686 755 1694 833
rect 1686 749 1687 755
rect 1693 749 1694 755
rect 1686 671 1694 749
rect 1686 665 1687 671
rect 1693 665 1694 671
rect 1686 591 1694 665
rect 1686 585 1687 591
rect 1693 585 1694 591
rect 1686 507 1694 585
rect 1686 501 1687 507
rect 1693 501 1694 507
rect 1686 427 1694 501
rect 1686 421 1687 427
rect 1693 421 1694 427
rect 1686 343 1694 421
rect 1686 337 1687 343
rect 1693 337 1694 343
rect 1686 259 1694 337
rect 1686 253 1687 259
rect 1693 253 1694 259
rect 1686 179 1694 253
rect 1686 173 1687 179
rect 1693 173 1694 179
rect 1686 83 1694 173
rect 1686 77 1687 83
rect 1693 77 1694 83
rect 1686 72 1694 77
rect 1698 1719 1706 1728
rect 1698 1713 1699 1719
rect 1705 1713 1706 1719
rect 1698 1639 1706 1713
rect 1698 1633 1699 1639
rect 1705 1633 1706 1639
rect 1698 1559 1706 1633
rect 1698 1553 1699 1559
rect 1705 1553 1706 1559
rect 1698 1475 1706 1553
rect 1698 1469 1699 1475
rect 1705 1469 1706 1475
rect 1698 1391 1706 1469
rect 1698 1385 1699 1391
rect 1705 1385 1706 1391
rect 1698 1307 1706 1385
rect 1698 1301 1699 1307
rect 1705 1301 1706 1307
rect 1698 1223 1706 1301
rect 1698 1217 1699 1223
rect 1705 1217 1706 1223
rect 1698 1135 1706 1217
rect 1698 1129 1699 1135
rect 1705 1129 1706 1135
rect 1698 1047 1706 1129
rect 1698 1041 1699 1047
rect 1705 1041 1706 1047
rect 1698 967 1706 1041
rect 1698 961 1699 967
rect 1705 961 1706 967
rect 1698 879 1706 961
rect 1698 873 1699 879
rect 1705 873 1706 879
rect 1698 795 1706 873
rect 1698 789 1699 795
rect 1705 789 1706 795
rect 1698 711 1706 789
rect 1698 705 1699 711
rect 1705 705 1706 711
rect 1698 631 1706 705
rect 1698 625 1699 631
rect 1705 625 1706 631
rect 1698 547 1706 625
rect 1698 541 1699 547
rect 1705 541 1706 547
rect 1698 467 1706 541
rect 1698 461 1699 467
rect 1705 461 1706 467
rect 1698 383 1706 461
rect 1698 377 1699 383
rect 1705 377 1706 383
rect 1698 303 1706 377
rect 1698 297 1699 303
rect 1705 297 1706 303
rect 1698 219 1706 297
rect 1698 213 1699 219
rect 1705 213 1706 219
rect 1698 123 1706 213
rect 1698 117 1699 123
rect 1705 117 1706 123
rect 1698 72 1706 117
use circuitwell  npwells
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use circuitppnp  ppnps
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use welltap_svt  __well_tap__77
timestamp 1731220528
transform 1 0 1656 0 1 1680
box 7 3 12 24
use welltap_svt  __well_tap__76
timestamp 1731220528
transform 1 0 104 0 1 1680
box 7 3 12 24
use welltap_svt  __well_tap__75
timestamp 1731220528
transform 1 0 1656 0 -1 1672
box 7 3 12 24
use welltap_svt  __well_tap__74
timestamp 1731220528
transform 1 0 104 0 -1 1672
box 7 3 12 24
use welltap_svt  __well_tap__73
timestamp 1731220528
transform 1 0 1656 0 1 1600
box 7 3 12 24
use welltap_svt  __well_tap__72
timestamp 1731220528
transform 1 0 104 0 1 1600
box 7 3 12 24
use welltap_svt  __well_tap__71
timestamp 1731220528
transform 1 0 1656 0 -1 1592
box 7 3 12 24
use welltap_svt  __well_tap__70
timestamp 1731220528
transform 1 0 104 0 -1 1592
box 7 3 12 24
use welltap_svt  __well_tap__69
timestamp 1731220528
transform 1 0 1656 0 1 1520
box 7 3 12 24
use welltap_svt  __well_tap__68
timestamp 1731220528
transform 1 0 104 0 1 1520
box 7 3 12 24
use welltap_svt  __well_tap__67
timestamp 1731220528
transform 1 0 1656 0 -1 1508
box 7 3 12 24
use welltap_svt  __well_tap__66
timestamp 1731220528
transform 1 0 104 0 -1 1508
box 7 3 12 24
use welltap_svt  __well_tap__65
timestamp 1731220528
transform 1 0 1656 0 1 1436
box 7 3 12 24
use welltap_svt  __well_tap__64
timestamp 1731220528
transform 1 0 104 0 1 1436
box 7 3 12 24
use welltap_svt  __well_tap__63
timestamp 1731220528
transform 1 0 1656 0 -1 1424
box 7 3 12 24
use welltap_svt  __well_tap__62
timestamp 1731220528
transform 1 0 104 0 -1 1424
box 7 3 12 24
use welltap_svt  __well_tap__61
timestamp 1731220528
transform 1 0 1656 0 1 1352
box 7 3 12 24
use welltap_svt  __well_tap__60
timestamp 1731220528
transform 1 0 104 0 1 1352
box 7 3 12 24
use welltap_svt  __well_tap__59
timestamp 1731220528
transform 1 0 1656 0 -1 1344
box 7 3 12 24
use welltap_svt  __well_tap__58
timestamp 1731220528
transform 1 0 104 0 -1 1344
box 7 3 12 24
use welltap_svt  __well_tap__57
timestamp 1731220528
transform 1 0 1656 0 1 1268
box 7 3 12 24
use welltap_svt  __well_tap__56
timestamp 1731220528
transform 1 0 104 0 1 1268
box 7 3 12 24
use welltap_svt  __well_tap__55
timestamp 1731220528
transform 1 0 1656 0 -1 1260
box 7 3 12 24
use welltap_svt  __well_tap__54
timestamp 1731220528
transform 1 0 104 0 -1 1260
box 7 3 12 24
use welltap_svt  __well_tap__53
timestamp 1731220528
transform 1 0 1656 0 1 1184
box 7 3 12 24
use welltap_svt  __well_tap__52
timestamp 1731220528
transform 1 0 104 0 1 1184
box 7 3 12 24
use welltap_svt  __well_tap__51
timestamp 1731220528
transform 1 0 1656 0 -1 1172
box 7 3 12 24
use welltap_svt  __well_tap__50
timestamp 1731220528
transform 1 0 104 0 -1 1172
box 7 3 12 24
use welltap_svt  __well_tap__49
timestamp 1731220528
transform 1 0 1656 0 1 1096
box 7 3 12 24
use welltap_svt  __well_tap__48
timestamp 1731220528
transform 1 0 104 0 1 1096
box 7 3 12 24
use welltap_svt  __well_tap__47
timestamp 1731220528
transform 1 0 1656 0 -1 1084
box 7 3 12 24
use welltap_svt  __well_tap__46
timestamp 1731220528
transform 1 0 104 0 -1 1084
box 7 3 12 24
use welltap_svt  __well_tap__45
timestamp 1731220528
transform 1 0 1656 0 1 1008
box 7 3 12 24
use welltap_svt  __well_tap__44
timestamp 1731220528
transform 1 0 104 0 1 1008
box 7 3 12 24
use welltap_svt  __well_tap__43
timestamp 1731220528
transform 1 0 1656 0 -1 1000
box 7 3 12 24
use welltap_svt  __well_tap__42
timestamp 1731220528
transform 1 0 104 0 -1 1000
box 7 3 12 24
use welltap_svt  __well_tap__41
timestamp 1731220528
transform 1 0 1656 0 1 928
box 7 3 12 24
use welltap_svt  __well_tap__40
timestamp 1731220528
transform 1 0 104 0 1 928
box 7 3 12 24
use welltap_svt  __well_tap__39
timestamp 1731220528
transform 1 0 1656 0 -1 916
box 7 3 12 24
use welltap_svt  __well_tap__38
timestamp 1731220528
transform 1 0 104 0 -1 916
box 7 3 12 24
use welltap_svt  __well_tap__37
timestamp 1731220528
transform 1 0 1656 0 1 840
box 7 3 12 24
use welltap_svt  __well_tap__36
timestamp 1731220528
transform 1 0 104 0 1 840
box 7 3 12 24
use welltap_svt  __well_tap__35
timestamp 1731220528
transform 1 0 1656 0 -1 832
box 7 3 12 24
use welltap_svt  __well_tap__34
timestamp 1731220528
transform 1 0 104 0 -1 832
box 7 3 12 24
use welltap_svt  __well_tap__33
timestamp 1731220528
transform 1 0 1656 0 1 756
box 7 3 12 24
use welltap_svt  __well_tap__32
timestamp 1731220528
transform 1 0 104 0 1 756
box 7 3 12 24
use welltap_svt  __well_tap__31
timestamp 1731220528
transform 1 0 1656 0 -1 748
box 7 3 12 24
use welltap_svt  __well_tap__30
timestamp 1731220528
transform 1 0 104 0 -1 748
box 7 3 12 24
use welltap_svt  __well_tap__29
timestamp 1731220528
transform 1 0 1656 0 1 672
box 7 3 12 24
use welltap_svt  __well_tap__28
timestamp 1731220528
transform 1 0 104 0 1 672
box 7 3 12 24
use welltap_svt  __well_tap__27
timestamp 1731220528
transform 1 0 1656 0 -1 664
box 7 3 12 24
use welltap_svt  __well_tap__26
timestamp 1731220528
transform 1 0 104 0 -1 664
box 7 3 12 24
use welltap_svt  __well_tap__25
timestamp 1731220528
transform 1 0 1656 0 1 592
box 7 3 12 24
use welltap_svt  __well_tap__24
timestamp 1731220528
transform 1 0 104 0 1 592
box 7 3 12 24
use welltap_svt  __well_tap__23
timestamp 1731220528
transform 1 0 1656 0 -1 584
box 7 3 12 24
use welltap_svt  __well_tap__22
timestamp 1731220528
transform 1 0 104 0 -1 584
box 7 3 12 24
use welltap_svt  __well_tap__21
timestamp 1731220528
transform 1 0 1656 0 1 508
box 7 3 12 24
use welltap_svt  __well_tap__20
timestamp 1731220528
transform 1 0 104 0 1 508
box 7 3 12 24
use welltap_svt  __well_tap__19
timestamp 1731220528
transform 1 0 1656 0 -1 500
box 7 3 12 24
use welltap_svt  __well_tap__18
timestamp 1731220528
transform 1 0 104 0 -1 500
box 7 3 12 24
use welltap_svt  __well_tap__17
timestamp 1731220528
transform 1 0 1656 0 1 428
box 7 3 12 24
use welltap_svt  __well_tap__16
timestamp 1731220528
transform 1 0 104 0 1 428
box 7 3 12 24
use welltap_svt  __well_tap__15
timestamp 1731220528
transform 1 0 1656 0 -1 420
box 7 3 12 24
use welltap_svt  __well_tap__14
timestamp 1731220528
transform 1 0 104 0 -1 420
box 7 3 12 24
use welltap_svt  __well_tap__13
timestamp 1731220528
transform 1 0 1656 0 1 344
box 7 3 12 24
use welltap_svt  __well_tap__12
timestamp 1731220528
transform 1 0 104 0 1 344
box 7 3 12 24
use welltap_svt  __well_tap__11
timestamp 1731220528
transform 1 0 1656 0 -1 336
box 7 3 12 24
use welltap_svt  __well_tap__10
timestamp 1731220528
transform 1 0 104 0 -1 336
box 7 3 12 24
use welltap_svt  __well_tap__9
timestamp 1731220528
transform 1 0 1656 0 1 264
box 7 3 12 24
use welltap_svt  __well_tap__8
timestamp 1731220528
transform 1 0 104 0 1 264
box 7 3 12 24
use welltap_svt  __well_tap__7
timestamp 1731220528
transform 1 0 1656 0 -1 252
box 7 3 12 24
use welltap_svt  __well_tap__6
timestamp 1731220528
transform 1 0 104 0 -1 252
box 7 3 12 24
use welltap_svt  __well_tap__5
timestamp 1731220528
transform 1 0 1656 0 1 180
box 7 3 12 24
use welltap_svt  __well_tap__4
timestamp 1731220528
transform 1 0 104 0 1 180
box 7 3 12 24
use welltap_svt  __well_tap__3
timestamp 1731220528
transform 1 0 1656 0 -1 172
box 7 3 12 24
use welltap_svt  __well_tap__2
timestamp 1731220528
transform 1 0 104 0 -1 172
box 7 3 12 24
use welltap_svt  __well_tap__1
timestamp 1731220528
transform 1 0 1656 0 1 84
box 7 3 12 24
use welltap_svt  __well_tap__0
timestamp 1731220528
transform 1 0 104 0 1 84
box 7 3 12 24
use _0_0std_0_0cells_0_0INVX1  tst_5999_6
timestamp 1731220528
transform 1 0 1584 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5998_6
timestamp 1731220528
transform 1 0 1616 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5997_6
timestamp 1731220528
transform 1 0 1616 0 -1 176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5996_6
timestamp 1731220528
transform 1 0 1616 0 1 176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5995_6
timestamp 1731220528
transform 1 0 1576 0 1 176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5994_6
timestamp 1731220528
transform 1 0 1520 0 1 176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5993_6
timestamp 1731220528
transform 1 0 1616 0 -1 256
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5992_6
timestamp 1731220528
transform 1 0 1568 0 -1 256
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5991_6
timestamp 1731220528
transform 1 0 1512 0 -1 256
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5990_6
timestamp 1731220528
transform 1 0 1456 0 -1 256
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5989_6
timestamp 1731220528
transform 1 0 1464 0 1 176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5988_6
timestamp 1731220528
transform 1 0 1408 0 1 176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5987_6
timestamp 1731220528
transform 1 0 1416 0 -1 176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5986_6
timestamp 1731220528
transform 1 0 1488 0 -1 176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5985_6
timestamp 1731220528
transform 1 0 1560 0 -1 176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5984_6
timestamp 1731220528
transform 1 0 1544 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5983_6
timestamp 1731220528
transform 1 0 1496 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5982_6
timestamp 1731220528
transform 1 0 1448 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5981_6
timestamp 1731220528
transform 1 0 1408 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5980_6
timestamp 1731220528
transform 1 0 1368 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5979_6
timestamp 1731220528
transform 1 0 1328 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5978_6
timestamp 1731220528
transform 1 0 1288 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5977_6
timestamp 1731220528
transform 1 0 1256 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5976_6
timestamp 1731220528
transform 1 0 1216 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5975_6
timestamp 1731220528
transform 1 0 1176 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5974_6
timestamp 1731220528
transform 1 0 1200 0 -1 176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5973_6
timestamp 1731220528
transform 1 0 1272 0 -1 176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5972_6
timestamp 1731220528
transform 1 0 1344 0 -1 176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5971_6
timestamp 1731220528
transform 1 0 1344 0 1 176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5970_6
timestamp 1731220528
transform 1 0 1280 0 1 176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5969_6
timestamp 1731220528
transform 1 0 1304 0 -1 256
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5968_6
timestamp 1731220528
transform 1 0 1360 0 -1 256
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5967_6
timestamp 1731220528
transform 1 0 1408 0 -1 256
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5966_6
timestamp 1731220528
transform 1 0 1384 0 1 260
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5965_6
timestamp 1731220528
transform 1 0 1320 0 1 260
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5964_6
timestamp 1731220528
transform 1 0 1440 0 1 260
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5963_6
timestamp 1731220528
transform 1 0 1488 0 1 260
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5962_6
timestamp 1731220528
transform 1 0 1536 0 1 260
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5961_6
timestamp 1731220528
transform 1 0 1584 0 1 260
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5960_6
timestamp 1731220528
transform 1 0 1616 0 1 260
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5959_6
timestamp 1731220528
transform 1 0 1616 0 -1 340
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5958_6
timestamp 1731220528
transform 1 0 1616 0 1 340
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5957_6
timestamp 1731220528
transform 1 0 1584 0 1 340
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5956_6
timestamp 1731220528
transform 1 0 1536 0 1 340
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5955_6
timestamp 1731220528
transform 1 0 1488 0 1 340
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5954_6
timestamp 1731220528
transform 1 0 1576 0 -1 340
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5953_6
timestamp 1731220528
transform 1 0 1512 0 -1 340
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5952_6
timestamp 1731220528
transform 1 0 1456 0 -1 340
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5951_6
timestamp 1731220528
transform 1 0 1400 0 -1 340
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5950_6
timestamp 1731220528
transform 1 0 1336 0 -1 340
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5949_6
timestamp 1731220528
transform 1 0 1440 0 1 340
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5948_6
timestamp 1731220528
transform 1 0 1392 0 1 340
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5947_6
timestamp 1731220528
transform 1 0 1344 0 1 340
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5946_6
timestamp 1731220528
transform 1 0 1296 0 1 340
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5945_6
timestamp 1731220528
transform 1 0 1248 0 1 340
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5944_6
timestamp 1731220528
transform 1 0 1200 0 1 340
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5943_6
timestamp 1731220528
transform 1 0 1160 0 -1 424
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5942_6
timestamp 1731220528
transform 1 0 1200 0 -1 424
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5941_6
timestamp 1731220528
transform 1 0 1240 0 -1 424
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5940_6
timestamp 1731220528
transform 1 0 1280 0 -1 424
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5939_6
timestamp 1731220528
transform 1 0 1376 0 -1 424
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5938_6
timestamp 1731220528
transform 1 0 1328 0 -1 424
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5937_6
timestamp 1731220528
transform 1 0 1312 0 1 424
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5936_6
timestamp 1731220528
transform 1 0 1256 0 1 424
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5935_6
timestamp 1731220528
transform 1 0 1368 0 1 424
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5934_6
timestamp 1731220528
transform 1 0 1424 0 1 424
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5933_6
timestamp 1731220528
transform 1 0 1488 0 1 424
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5932_6
timestamp 1731220528
transform 1 0 1472 0 -1 504
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5931_6
timestamp 1731220528
transform 1 0 1424 0 -1 504
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5930_6
timestamp 1731220528
transform 1 0 1528 0 -1 504
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5929_6
timestamp 1731220528
transform 1 0 1616 0 -1 504
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5928_6
timestamp 1731220528
transform 1 0 1584 0 -1 504
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5927_6
timestamp 1731220528
transform 1 0 1568 0 1 504
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5926_6
timestamp 1731220528
transform 1 0 1616 0 1 504
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5925_6
timestamp 1731220528
transform 1 0 1616 0 -1 588
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5924_6
timestamp 1731220528
transform 1 0 1616 0 1 588
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5923_6
timestamp 1731220528
transform 1 0 1616 0 -1 668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5922_6
timestamp 1731220528
transform 1 0 1616 0 1 668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5921_6
timestamp 1731220528
transform 1 0 1576 0 1 668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5920_6
timestamp 1731220528
transform 1 0 1616 0 -1 752
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5919_6
timestamp 1731220528
transform 1 0 1576 0 -1 752
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5918_6
timestamp 1731220528
transform 1 0 1520 0 1 668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5917_6
timestamp 1731220528
transform 1 0 1464 0 1 668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5916_6
timestamp 1731220528
transform 1 0 1464 0 -1 668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5915_6
timestamp 1731220528
transform 1 0 1552 0 -1 668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5914_6
timestamp 1731220528
transform 1 0 1568 0 1 588
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5913_6
timestamp 1731220528
transform 1 0 1496 0 1 588
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5912_6
timestamp 1731220528
transform 1 0 1424 0 1 588
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5911_6
timestamp 1731220528
transform 1 0 1352 0 1 588
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5910_6
timestamp 1731220528
transform 1 0 1568 0 -1 588
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5909_6
timestamp 1731220528
transform 1 0 1504 0 -1 588
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5908_6
timestamp 1731220528
transform 1 0 1440 0 -1 588
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5907_6
timestamp 1731220528
transform 1 0 1376 0 -1 588
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5906_6
timestamp 1731220528
transform 1 0 1320 0 -1 588
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5905_6
timestamp 1731220528
transform 1 0 1504 0 1 504
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5904_6
timestamp 1731220528
transform 1 0 1440 0 1 504
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5903_6
timestamp 1731220528
transform 1 0 1384 0 1 504
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5902_6
timestamp 1731220528
transform 1 0 1328 0 1 504
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5901_6
timestamp 1731220528
transform 1 0 1272 0 1 504
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5900_6
timestamp 1731220528
transform 1 0 1224 0 1 504
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5899_6
timestamp 1731220528
transform 1 0 1376 0 -1 504
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5898_6
timestamp 1731220528
transform 1 0 1328 0 -1 504
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5897_6
timestamp 1731220528
transform 1 0 1280 0 -1 504
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5896_6
timestamp 1731220528
transform 1 0 1232 0 -1 504
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5895_6
timestamp 1731220528
transform 1 0 1184 0 -1 504
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5894_6
timestamp 1731220528
transform 1 0 1136 0 -1 504
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5893_6
timestamp 1731220528
transform 1 0 1088 0 -1 504
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5892_6
timestamp 1731220528
transform 1 0 1032 0 -1 504
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5891_6
timestamp 1731220528
transform 1 0 976 0 -1 504
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5890_6
timestamp 1731220528
transform 1 0 912 0 -1 504
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5889_6
timestamp 1731220528
transform 1 0 1064 0 1 504
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5888_6
timestamp 1731220528
transform 1 0 1120 0 1 504
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5887_6
timestamp 1731220528
transform 1 0 1176 0 1 504
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5886_6
timestamp 1731220528
transform 1 0 1152 0 -1 588
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5885_6
timestamp 1731220528
transform 1 0 1208 0 -1 588
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5884_6
timestamp 1731220528
transform 1 0 1264 0 -1 588
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5883_6
timestamp 1731220528
transform 1 0 1280 0 1 588
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5882_6
timestamp 1731220528
transform 1 0 1200 0 1 588
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5881_6
timestamp 1731220528
transform 1 0 1208 0 -1 668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5880_6
timestamp 1731220528
transform 1 0 1288 0 -1 668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5879_6
timestamp 1731220528
transform 1 0 1376 0 -1 668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5878_6
timestamp 1731220528
transform 1 0 1408 0 1 668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5877_6
timestamp 1731220528
transform 1 0 1344 0 1 668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5876_6
timestamp 1731220528
transform 1 0 1280 0 1 668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5875_6
timestamp 1731220528
transform 1 0 1216 0 1 668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5874_6
timestamp 1731220528
transform 1 0 1152 0 1 668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5873_6
timestamp 1731220528
transform 1 0 1232 0 -1 752
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5872_6
timestamp 1731220528
transform 1 0 1288 0 -1 752
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5871_6
timestamp 1731220528
transform 1 0 1344 0 -1 752
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5870_6
timestamp 1731220528
transform 1 0 1400 0 -1 752
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5869_6
timestamp 1731220528
transform 1 0 1456 0 -1 752
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5868_6
timestamp 1731220528
transform 1 0 1512 0 -1 752
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5867_6
timestamp 1731220528
transform 1 0 1464 0 1 752
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5866_6
timestamp 1731220528
transform 1 0 1408 0 1 752
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5865_6
timestamp 1731220528
transform 1 0 1352 0 1 752
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5864_6
timestamp 1731220528
transform 1 0 1520 0 1 752
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5863_6
timestamp 1731220528
transform 1 0 1584 0 1 752
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5862_6
timestamp 1731220528
transform 1 0 1584 0 -1 836
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5861_6
timestamp 1731220528
transform 1 0 1528 0 -1 836
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5860_6
timestamp 1731220528
transform 1 0 1472 0 -1 836
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5859_6
timestamp 1731220528
transform 1 0 1416 0 -1 836
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5858_6
timestamp 1731220528
transform 1 0 1360 0 -1 836
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5857_6
timestamp 1731220528
transform 1 0 1304 0 -1 836
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5856_6
timestamp 1731220528
transform 1 0 1456 0 1 836
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5855_6
timestamp 1731220528
transform 1 0 1392 0 1 836
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5854_6
timestamp 1731220528
transform 1 0 1336 0 1 836
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5853_6
timestamp 1731220528
transform 1 0 1280 0 1 836
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5852_6
timestamp 1731220528
transform 1 0 1224 0 1 836
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5851_6
timestamp 1731220528
transform 1 0 1160 0 1 836
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5850_6
timestamp 1731220528
transform 1 0 1376 0 -1 920
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5849_6
timestamp 1731220528
transform 1 0 1312 0 -1 920
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5848_6
timestamp 1731220528
transform 1 0 1248 0 -1 920
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5847_6
timestamp 1731220528
transform 1 0 1192 0 -1 920
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5846_6
timestamp 1731220528
transform 1 0 1136 0 -1 920
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5845_6
timestamp 1731220528
transform 1 0 1224 0 1 924
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5844_6
timestamp 1731220528
transform 1 0 1280 0 1 924
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5843_6
timestamp 1731220528
transform 1 0 1336 0 1 924
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5842_6
timestamp 1731220528
transform 1 0 1280 0 -1 1004
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5841_6
timestamp 1731220528
transform 1 0 1336 0 -1 1004
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5840_6
timestamp 1731220528
transform 1 0 1392 0 -1 1004
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5839_6
timestamp 1731220528
transform 1 0 1376 0 1 1004
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5838_6
timestamp 1731220528
transform 1 0 1328 0 1 1004
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5837_6
timestamp 1731220528
transform 1 0 1424 0 1 1004
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5836_6
timestamp 1731220528
transform 1 0 1472 0 1 1004
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5835_6
timestamp 1731220528
transform 1 0 1528 0 1 1004
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5834_6
timestamp 1731220528
transform 1 0 1536 0 -1 1004
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5833_6
timestamp 1731220528
transform 1 0 1488 0 -1 1004
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5832_6
timestamp 1731220528
transform 1 0 1440 0 -1 1004
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5831_6
timestamp 1731220528
transform 1 0 1424 0 1 924
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5830_6
timestamp 1731220528
transform 1 0 1384 0 1 924
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5829_6
timestamp 1731220528
transform 1 0 1464 0 1 924
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5828_6
timestamp 1731220528
transform 1 0 1504 0 1 924
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5827_6
timestamp 1731220528
transform 1 0 1544 0 1 924
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5826_6
timestamp 1731220528
transform 1 0 1616 0 1 924
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5825_6
timestamp 1731220528
transform 1 0 1584 0 1 924
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5824_6
timestamp 1731220528
transform 1 0 1584 0 -1 1004
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5823_6
timestamp 1731220528
transform 1 0 1616 0 -1 1004
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5822_6
timestamp 1731220528
transform 1 0 1616 0 1 1004
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5821_6
timestamp 1731220528
transform 1 0 1584 0 1 1004
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5820_6
timestamp 1731220528
transform 1 0 1616 0 -1 1088
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5819_6
timestamp 1731220528
transform 1 0 1616 0 1 1092
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5818_6
timestamp 1731220528
transform 1 0 1584 0 1 1092
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5817_6
timestamp 1731220528
transform 1 0 1536 0 1 1092
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5816_6
timestamp 1731220528
transform 1 0 1584 0 -1 1088
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5815_6
timestamp 1731220528
transform 1 0 1544 0 -1 1088
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5814_6
timestamp 1731220528
transform 1 0 1496 0 -1 1088
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5813_6
timestamp 1731220528
transform 1 0 1456 0 -1 1088
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5812_6
timestamp 1731220528
transform 1 0 1408 0 -1 1088
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5811_6
timestamp 1731220528
transform 1 0 1352 0 -1 1088
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5810_6
timestamp 1731220528
transform 1 0 1488 0 1 1092
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5809_6
timestamp 1731220528
transform 1 0 1440 0 1 1092
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5808_6
timestamp 1731220528
transform 1 0 1384 0 1 1092
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5807_6
timestamp 1731220528
transform 1 0 1328 0 1 1092
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5806_6
timestamp 1731220528
transform 1 0 1552 0 -1 1176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5805_6
timestamp 1731220528
transform 1 0 1472 0 -1 1176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5804_6
timestamp 1731220528
transform 1 0 1400 0 -1 1176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5803_6
timestamp 1731220528
transform 1 0 1336 0 -1 1176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5802_6
timestamp 1731220528
transform 1 0 1272 0 -1 1176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5801_6
timestamp 1731220528
transform 1 0 1208 0 -1 1176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5800_6
timestamp 1731220528
transform 1 0 1536 0 1 1180
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5799_6
timestamp 1731220528
transform 1 0 1440 0 1 1180
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5798_6
timestamp 1731220528
transform 1 0 1352 0 1 1180
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5797_6
timestamp 1731220528
transform 1 0 1272 0 1 1180
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5796_6
timestamp 1731220528
transform 1 0 1200 0 1 1180
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5795_6
timestamp 1731220528
transform 1 0 1136 0 1 1180
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5794_6
timestamp 1731220528
transform 1 0 1528 0 -1 1264
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5793_6
timestamp 1731220528
transform 1 0 1416 0 -1 1264
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5792_6
timestamp 1731220528
transform 1 0 1312 0 -1 1264
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5791_6
timestamp 1731220528
transform 1 0 1224 0 -1 1264
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5790_6
timestamp 1731220528
transform 1 0 1152 0 -1 1264
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5789_6
timestamp 1731220528
transform 1 0 1088 0 -1 1264
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5788_6
timestamp 1731220528
transform 1 0 1136 0 1 1264
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5787_6
timestamp 1731220528
transform 1 0 1200 0 1 1264
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5786_6
timestamp 1731220528
transform 1 0 1272 0 1 1264
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5785_6
timestamp 1731220528
transform 1 0 1536 0 1 1264
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5784_6
timestamp 1731220528
transform 1 0 1440 0 1 1264
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5783_6
timestamp 1731220528
transform 1 0 1352 0 1 1264
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5782_6
timestamp 1731220528
transform 1 0 1336 0 -1 1348
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5781_6
timestamp 1731220528
transform 1 0 1272 0 -1 1348
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5780_6
timestamp 1731220528
transform 1 0 1208 0 -1 1348
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5779_6
timestamp 1731220528
transform 1 0 1400 0 -1 1348
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5778_6
timestamp 1731220528
transform 1 0 1552 0 -1 1348
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5777_6
timestamp 1731220528
transform 1 0 1472 0 -1 1348
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5776_6
timestamp 1731220528
transform 1 0 1424 0 1 1348
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5775_6
timestamp 1731220528
transform 1 0 1360 0 1 1348
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5774_6
timestamp 1731220528
transform 1 0 1296 0 1 1348
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5773_6
timestamp 1731220528
transform 1 0 1560 0 1 1348
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5772_6
timestamp 1731220528
transform 1 0 1488 0 1 1348
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5771_6
timestamp 1731220528
transform 1 0 1456 0 -1 1428
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5770_6
timestamp 1731220528
transform 1 0 1408 0 -1 1428
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5769_6
timestamp 1731220528
transform 1 0 1352 0 -1 1428
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5768_6
timestamp 1731220528
transform 1 0 1496 0 -1 1428
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5767_6
timestamp 1731220528
transform 1 0 1552 0 1 1432
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5766_6
timestamp 1731220528
transform 1 0 1544 0 -1 1428
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5765_6
timestamp 1731220528
transform 1 0 1584 0 -1 1428
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5764_6
timestamp 1731220528
transform 1 0 1616 0 1 1348
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5763_6
timestamp 1731220528
transform 1 0 1616 0 1 1264
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5762_6
timestamp 1731220528
transform 1 0 1616 0 -1 1176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5761_6
timestamp 1731220528
transform 1 0 1616 0 1 1180
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5760_6
timestamp 1731220528
transform 1 0 1616 0 -1 1264
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5759_6
timestamp 1731220528
transform 1 0 1616 0 -1 1348
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5758_6
timestamp 1731220528
transform 1 0 1616 0 -1 1428
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5757_6
timestamp 1731220528
transform 1 0 1616 0 1 1432
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5756_6
timestamp 1731220528
transform 1 0 1616 0 -1 1512
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5755_6
timestamp 1731220528
transform 1 0 1616 0 1 1516
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5754_6
timestamp 1731220528
transform 1 0 1616 0 -1 1596
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5753_6
timestamp 1731220528
transform 1 0 1616 0 1 1596
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5752_6
timestamp 1731220528
transform 1 0 1616 0 -1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5751_6
timestamp 1731220528
transform 1 0 1576 0 -1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5750_6
timestamp 1731220528
transform 1 0 1520 0 -1 1596
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5749_6
timestamp 1731220528
transform 1 0 1576 0 -1 1596
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5748_6
timestamp 1731220528
transform 1 0 1576 0 1 1516
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5747_6
timestamp 1731220528
transform 1 0 1520 0 1 1516
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5746_6
timestamp 1731220528
transform 1 0 1464 0 1 1516
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5745_6
timestamp 1731220528
transform 1 0 1400 0 1 1516
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5744_6
timestamp 1731220528
transform 1 0 1328 0 1 1516
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5743_6
timestamp 1731220528
transform 1 0 1344 0 -1 1596
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5742_6
timestamp 1731220528
transform 1 0 1464 0 -1 1596
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5741_6
timestamp 1731220528
transform 1 0 1408 0 -1 1596
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5740_6
timestamp 1731220528
transform 1 0 1392 0 1 1596
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5739_6
timestamp 1731220528
transform 1 0 1472 0 1 1596
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5738_6
timestamp 1731220528
transform 1 0 1552 0 1 1596
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5737_6
timestamp 1731220528
transform 1 0 1512 0 -1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5736_6
timestamp 1731220528
transform 1 0 1448 0 -1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5735_6
timestamp 1731220528
transform 1 0 1384 0 -1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5734_6
timestamp 1731220528
transform 1 0 1512 0 1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5733_6
timestamp 1731220528
transform 1 0 1464 0 1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5732_6
timestamp 1731220528
transform 1 0 1416 0 1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5731_6
timestamp 1731220528
transform 1 0 1368 0 1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5730_6
timestamp 1731220528
transform 1 0 1328 0 1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5729_6
timestamp 1731220528
transform 1 0 1280 0 1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5728_6
timestamp 1731220528
transform 1 0 1224 0 1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5727_6
timestamp 1731220528
transform 1 0 1240 0 -1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5726_6
timestamp 1731220528
transform 1 0 1312 0 -1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5725_6
timestamp 1731220528
transform 1 0 1312 0 1 1596
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5724_6
timestamp 1731220528
transform 1 0 1240 0 1 1596
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5723_6
timestamp 1731220528
transform 1 0 1272 0 -1 1596
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5722_6
timestamp 1731220528
transform 1 0 1256 0 1 1516
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5721_6
timestamp 1731220528
transform 1 0 1560 0 -1 1512
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5720_6
timestamp 1731220528
transform 1 0 1480 0 -1 1512
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5719_6
timestamp 1731220528
transform 1 0 1408 0 -1 1512
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5718_6
timestamp 1731220528
transform 1 0 1344 0 -1 1512
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5717_6
timestamp 1731220528
transform 1 0 1288 0 -1 1512
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5716_6
timestamp 1731220528
transform 1 0 1248 0 -1 1512
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5715_6
timestamp 1731220528
transform 1 0 1472 0 1 1432
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5714_6
timestamp 1731220528
transform 1 0 1392 0 1 1432
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5713_6
timestamp 1731220528
transform 1 0 1320 0 1 1432
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5712_6
timestamp 1731220528
transform 1 0 1256 0 1 1432
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5711_6
timestamp 1731220528
transform 1 0 1200 0 1 1432
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5710_6
timestamp 1731220528
transform 1 0 1152 0 1 1432
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5709_6
timestamp 1731220528
transform 1 0 1208 0 -1 1512
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5708_6
timestamp 1731220528
transform 1 0 1176 0 -1 1512
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5707_6
timestamp 1731220528
transform 1 0 1144 0 -1 1512
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5706_6
timestamp 1731220528
transform 1 0 1104 0 -1 1512
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5705_6
timestamp 1731220528
transform 1 0 1056 0 -1 1512
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5704_6
timestamp 1731220528
transform 1 0 1000 0 -1 1512
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5703_6
timestamp 1731220528
transform 1 0 1008 0 1 1432
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5702_6
timestamp 1731220528
transform 1 0 1064 0 1 1432
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5701_6
timestamp 1731220528
transform 1 0 1112 0 1 1432
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5700_6
timestamp 1731220528
transform 1 0 1288 0 -1 1428
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5699_6
timestamp 1731220528
transform 1 0 1224 0 -1 1428
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5698_6
timestamp 1731220528
transform 1 0 1160 0 -1 1428
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5697_6
timestamp 1731220528
transform 1 0 1096 0 -1 1428
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5696_6
timestamp 1731220528
transform 1 0 1024 0 -1 1428
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5695_6
timestamp 1731220528
transform 1 0 960 0 -1 1428
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5694_6
timestamp 1731220528
transform 1 0 1232 0 1 1348
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5693_6
timestamp 1731220528
transform 1 0 1168 0 1 1348
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5692_6
timestamp 1731220528
transform 1 0 1096 0 1 1348
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5691_6
timestamp 1731220528
transform 1 0 1024 0 1 1348
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5690_6
timestamp 1731220528
transform 1 0 952 0 1 1348
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5689_6
timestamp 1731220528
transform 1 0 880 0 1 1348
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5688_6
timestamp 1731220528
transform 1 0 1144 0 -1 1348
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5687_6
timestamp 1731220528
transform 1 0 1080 0 -1 1348
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5686_6
timestamp 1731220528
transform 1 0 1016 0 -1 1348
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5685_6
timestamp 1731220528
transform 1 0 952 0 -1 1348
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5684_6
timestamp 1731220528
transform 1 0 880 0 -1 1348
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5683_6
timestamp 1731220528
transform 1 0 816 0 -1 1348
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5682_6
timestamp 1731220528
transform 1 0 1072 0 1 1264
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5681_6
timestamp 1731220528
transform 1 0 1016 0 1 1264
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5680_6
timestamp 1731220528
transform 1 0 952 0 1 1264
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5679_6
timestamp 1731220528
transform 1 0 888 0 1 1264
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5678_6
timestamp 1731220528
transform 1 0 824 0 1 1264
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5677_6
timestamp 1731220528
transform 1 0 768 0 1 1264
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5676_6
timestamp 1731220528
transform 1 0 760 0 -1 1264
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5675_6
timestamp 1731220528
transform 1 0 712 0 1 1264
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5674_6
timestamp 1731220528
transform 1 0 712 0 -1 1264
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5673_6
timestamp 1731220528
transform 1 0 656 0 -1 1264
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5672_6
timestamp 1731220528
transform 1 0 808 0 -1 1264
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5671_6
timestamp 1731220528
transform 1 0 864 0 -1 1264
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5670_6
timestamp 1731220528
transform 1 0 1032 0 -1 1264
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5669_6
timestamp 1731220528
transform 1 0 976 0 -1 1264
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5668_6
timestamp 1731220528
transform 1 0 920 0 -1 1264
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5667_6
timestamp 1731220528
transform 1 0 880 0 1 1180
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5666_6
timestamp 1731220528
transform 1 0 816 0 1 1180
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5665_6
timestamp 1731220528
transform 1 0 760 0 1 1180
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5664_6
timestamp 1731220528
transform 1 0 944 0 1 1180
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5663_6
timestamp 1731220528
transform 1 0 1072 0 1 1180
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5662_6
timestamp 1731220528
transform 1 0 1008 0 1 1180
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5661_6
timestamp 1731220528
transform 1 0 960 0 -1 1176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5660_6
timestamp 1731220528
transform 1 0 896 0 -1 1176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5659_6
timestamp 1731220528
transform 1 0 832 0 -1 1176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5658_6
timestamp 1731220528
transform 1 0 1152 0 -1 1176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5657_6
timestamp 1731220528
transform 1 0 1088 0 -1 1176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5656_6
timestamp 1731220528
transform 1 0 1024 0 -1 1176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5655_6
timestamp 1731220528
transform 1 0 1016 0 1 1092
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5654_6
timestamp 1731220528
transform 1 0 960 0 1 1092
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5653_6
timestamp 1731220528
transform 1 0 904 0 1 1092
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5652_6
timestamp 1731220528
transform 1 0 1080 0 1 1092
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5651_6
timestamp 1731220528
transform 1 0 1272 0 1 1092
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5650_6
timestamp 1731220528
transform 1 0 1208 0 1 1092
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5649_6
timestamp 1731220528
transform 1 0 1144 0 1 1092
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5648_6
timestamp 1731220528
transform 1 0 1104 0 -1 1088
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5647_6
timestamp 1731220528
transform 1 0 1032 0 -1 1088
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5646_6
timestamp 1731220528
transform 1 0 960 0 -1 1088
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5645_6
timestamp 1731220528
transform 1 0 1168 0 -1 1088
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5644_6
timestamp 1731220528
transform 1 0 1232 0 -1 1088
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5643_6
timestamp 1731220528
transform 1 0 1296 0 -1 1088
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5642_6
timestamp 1731220528
transform 1 0 1272 0 1 1004
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5641_6
timestamp 1731220528
transform 1 0 1216 0 1 1004
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5640_6
timestamp 1731220528
transform 1 0 1152 0 1 1004
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5639_6
timestamp 1731220528
transform 1 0 1088 0 1 1004
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5638_6
timestamp 1731220528
transform 1 0 1024 0 1 1004
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5637_6
timestamp 1731220528
transform 1 0 952 0 1 1004
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5636_6
timestamp 1731220528
transform 1 0 1216 0 -1 1004
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5635_6
timestamp 1731220528
transform 1 0 1152 0 -1 1004
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5634_6
timestamp 1731220528
transform 1 0 1088 0 -1 1004
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5633_6
timestamp 1731220528
transform 1 0 1024 0 -1 1004
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5632_6
timestamp 1731220528
transform 1 0 960 0 -1 1004
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5631_6
timestamp 1731220528
transform 1 0 896 0 -1 1004
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5630_6
timestamp 1731220528
transform 1 0 1160 0 1 924
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5629_6
timestamp 1731220528
transform 1 0 1096 0 1 924
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5628_6
timestamp 1731220528
transform 1 0 1032 0 1 924
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5627_6
timestamp 1731220528
transform 1 0 968 0 1 924
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5626_6
timestamp 1731220528
transform 1 0 904 0 1 924
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5625_6
timestamp 1731220528
transform 1 0 840 0 1 924
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5624_6
timestamp 1731220528
transform 1 0 1080 0 -1 920
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5623_6
timestamp 1731220528
transform 1 0 1016 0 -1 920
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5622_6
timestamp 1731220528
transform 1 0 952 0 -1 920
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5621_6
timestamp 1731220528
transform 1 0 896 0 -1 920
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5620_6
timestamp 1731220528
transform 1 0 840 0 -1 920
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5619_6
timestamp 1731220528
transform 1 0 792 0 -1 920
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5618_6
timestamp 1731220528
transform 1 0 792 0 1 836
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5617_6
timestamp 1731220528
transform 1 0 840 0 1 836
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5616_6
timestamp 1731220528
transform 1 0 896 0 1 836
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5615_6
timestamp 1731220528
transform 1 0 960 0 1 836
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5614_6
timestamp 1731220528
transform 1 0 1096 0 1 836
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5613_6
timestamp 1731220528
transform 1 0 1032 0 1 836
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5612_6
timestamp 1731220528
transform 1 0 1032 0 -1 836
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5611_6
timestamp 1731220528
transform 1 0 968 0 -1 836
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5610_6
timestamp 1731220528
transform 1 0 904 0 -1 836
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5609_6
timestamp 1731220528
transform 1 0 1104 0 -1 836
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5608_6
timestamp 1731220528
transform 1 0 1176 0 -1 836
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5607_6
timestamp 1731220528
transform 1 0 1240 0 -1 836
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5606_6
timestamp 1731220528
transform 1 0 1288 0 1 752
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5605_6
timestamp 1731220528
transform 1 0 1224 0 1 752
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5604_6
timestamp 1731220528
transform 1 0 1160 0 1 752
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5603_6
timestamp 1731220528
transform 1 0 1088 0 1 752
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5602_6
timestamp 1731220528
transform 1 0 1016 0 1 752
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5601_6
timestamp 1731220528
transform 1 0 944 0 1 752
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5600_6
timestamp 1731220528
transform 1 0 1176 0 -1 752
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5599_6
timestamp 1731220528
transform 1 0 1112 0 -1 752
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5598_6
timestamp 1731220528
transform 1 0 1048 0 -1 752
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5597_6
timestamp 1731220528
transform 1 0 984 0 -1 752
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5596_6
timestamp 1731220528
transform 1 0 920 0 -1 752
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5595_6
timestamp 1731220528
transform 1 0 952 0 1 668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5594_6
timestamp 1731220528
transform 1 0 1080 0 1 668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5593_6
timestamp 1731220528
transform 1 0 1016 0 1 668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5592_6
timestamp 1731220528
transform 1 0 968 0 -1 668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5591_6
timestamp 1731220528
transform 1 0 1040 0 -1 668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5590_6
timestamp 1731220528
transform 1 0 1120 0 -1 668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5589_6
timestamp 1731220528
transform 1 0 1120 0 1 588
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5588_6
timestamp 1731220528
transform 1 0 1040 0 1 588
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5587_6
timestamp 1731220528
transform 1 0 1096 0 -1 588
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5586_6
timestamp 1731220528
transform 1 0 1040 0 -1 588
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5585_6
timestamp 1731220528
transform 1 0 984 0 -1 588
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5584_6
timestamp 1731220528
transform 1 0 1000 0 1 504
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5583_6
timestamp 1731220528
transform 1 0 936 0 1 504
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5582_6
timestamp 1731220528
transform 1 0 872 0 1 504
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5581_6
timestamp 1731220528
transform 1 0 872 0 -1 588
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5580_6
timestamp 1731220528
transform 1 0 816 0 -1 588
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5579_6
timestamp 1731220528
transform 1 0 928 0 -1 588
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5578_6
timestamp 1731220528
transform 1 0 960 0 1 588
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5577_6
timestamp 1731220528
transform 1 0 888 0 1 588
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5576_6
timestamp 1731220528
transform 1 0 824 0 1 588
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5575_6
timestamp 1731220528
transform 1 0 784 0 -1 668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5574_6
timestamp 1731220528
transform 1 0 840 0 -1 668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5573_6
timestamp 1731220528
transform 1 0 904 0 -1 668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5572_6
timestamp 1731220528
transform 1 0 880 0 1 668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5571_6
timestamp 1731220528
transform 1 0 816 0 1 668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5570_6
timestamp 1731220528
transform 1 0 752 0 1 668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5569_6
timestamp 1731220528
transform 1 0 728 0 -1 752
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5568_6
timestamp 1731220528
transform 1 0 792 0 -1 752
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5567_6
timestamp 1731220528
transform 1 0 856 0 -1 752
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5566_6
timestamp 1731220528
transform 1 0 864 0 1 752
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5565_6
timestamp 1731220528
transform 1 0 784 0 1 752
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5564_6
timestamp 1731220528
transform 1 0 696 0 1 752
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5563_6
timestamp 1731220528
transform 1 0 840 0 -1 836
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5562_6
timestamp 1731220528
transform 1 0 784 0 -1 836
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5561_6
timestamp 1731220528
transform 1 0 728 0 -1 836
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5560_6
timestamp 1731220528
transform 1 0 664 0 -1 836
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5559_6
timestamp 1731220528
transform 1 0 744 0 1 836
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5558_6
timestamp 1731220528
transform 1 0 696 0 1 836
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5557_6
timestamp 1731220528
transform 1 0 528 0 1 836
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5556_6
timestamp 1731220528
transform 1 0 464 0 1 836
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5555_6
timestamp 1731220528
transform 1 0 464 0 -1 920
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5554_6
timestamp 1731220528
transform 1 0 528 0 -1 920
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5553_6
timestamp 1731220528
transform 1 0 584 0 -1 920
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5552_6
timestamp 1731220528
transform 1 0 656 0 1 924
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5551_6
timestamp 1731220528
transform 1 0 592 0 1 924
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5550_6
timestamp 1731220528
transform 1 0 528 0 1 924
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5549_6
timestamp 1731220528
transform 1 0 464 0 1 924
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5548_6
timestamp 1731220528
transform 1 0 680 0 -1 1004
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5547_6
timestamp 1731220528
transform 1 0 608 0 -1 1004
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5546_6
timestamp 1731220528
transform 1 0 536 0 -1 1004
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5545_6
timestamp 1731220528
transform 1 0 472 0 -1 1004
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5544_6
timestamp 1731220528
transform 1 0 704 0 1 1004
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5543_6
timestamp 1731220528
transform 1 0 624 0 1 1004
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5542_6
timestamp 1731220528
transform 1 0 552 0 1 1004
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5541_6
timestamp 1731220528
transform 1 0 496 0 1 1004
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5540_6
timestamp 1731220528
transform 1 0 648 0 -1 1088
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5539_6
timestamp 1731220528
transform 1 0 568 0 -1 1088
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5538_6
timestamp 1731220528
transform 1 0 496 0 -1 1088
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5537_6
timestamp 1731220528
transform 1 0 432 0 -1 1088
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5536_6
timestamp 1731220528
transform 1 0 384 0 -1 1088
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5535_6
timestamp 1731220528
transform 1 0 344 0 -1 1088
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5534_6
timestamp 1731220528
transform 1 0 304 0 -1 1088
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5533_6
timestamp 1731220528
transform 1 0 448 0 1 1004
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5532_6
timestamp 1731220528
transform 1 0 416 0 1 1004
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5531_6
timestamp 1731220528
transform 1 0 384 0 1 1004
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5530_6
timestamp 1731220528
transform 1 0 352 0 1 1004
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5529_6
timestamp 1731220528
transform 1 0 320 0 1 1004
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5528_6
timestamp 1731220528
transform 1 0 288 0 1 1004
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5527_6
timestamp 1731220528
transform 1 0 416 0 -1 1004
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5526_6
timestamp 1731220528
transform 1 0 376 0 -1 1004
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5525_6
timestamp 1731220528
transform 1 0 336 0 -1 1004
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5524_6
timestamp 1731220528
transform 1 0 304 0 -1 1004
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5523_6
timestamp 1731220528
transform 1 0 272 0 -1 1004
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5522_6
timestamp 1731220528
transform 1 0 240 0 -1 1004
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5521_6
timestamp 1731220528
transform 1 0 400 0 1 924
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5520_6
timestamp 1731220528
transform 1 0 336 0 1 924
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5519_6
timestamp 1731220528
transform 1 0 280 0 1 924
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5518_6
timestamp 1731220528
transform 1 0 232 0 1 924
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5517_6
timestamp 1731220528
transform 1 0 192 0 1 924
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5516_6
timestamp 1731220528
transform 1 0 160 0 1 924
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5515_6
timestamp 1731220528
transform 1 0 400 0 -1 920
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5514_6
timestamp 1731220528
transform 1 0 328 0 -1 920
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5513_6
timestamp 1731220528
transform 1 0 264 0 -1 920
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5512_6
timestamp 1731220528
transform 1 0 200 0 -1 920
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5511_6
timestamp 1731220528
transform 1 0 160 0 -1 920
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5510_6
timestamp 1731220528
transform 1 0 128 0 -1 920
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5509_6
timestamp 1731220528
transform 1 0 400 0 1 836
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5508_6
timestamp 1731220528
transform 1 0 328 0 1 836
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5507_6
timestamp 1731220528
transform 1 0 264 0 1 836
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5506_6
timestamp 1731220528
transform 1 0 200 0 1 836
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5505_6
timestamp 1731220528
transform 1 0 160 0 1 836
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5504_6
timestamp 1731220528
transform 1 0 128 0 1 836
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5503_6
timestamp 1731220528
transform 1 0 128 0 -1 836
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5502_6
timestamp 1731220528
transform 1 0 160 0 -1 836
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5501_6
timestamp 1731220528
transform 1 0 208 0 -1 836
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5500_6
timestamp 1731220528
transform 1 0 408 0 -1 836
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5499_6
timestamp 1731220528
transform 1 0 336 0 -1 836
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5498_6
timestamp 1731220528
transform 1 0 272 0 -1 836
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5497_6
timestamp 1731220528
transform 1 0 224 0 1 752
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5496_6
timestamp 1731220528
transform 1 0 168 0 1 752
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5495_6
timestamp 1731220528
transform 1 0 128 0 1 752
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5494_6
timestamp 1731220528
transform 1 0 440 0 1 752
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5493_6
timestamp 1731220528
transform 1 0 360 0 1 752
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5492_6
timestamp 1731220528
transform 1 0 288 0 1 752
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5491_6
timestamp 1731220528
transform 1 0 272 0 -1 752
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5490_6
timestamp 1731220528
transform 1 0 240 0 -1 752
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5489_6
timestamp 1731220528
transform 1 0 208 0 -1 752
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5488_6
timestamp 1731220528
transform 1 0 312 0 -1 752
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5487_6
timestamp 1731220528
transform 1 0 392 0 -1 752
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5486_6
timestamp 1731220528
transform 1 0 352 0 -1 752
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5485_6
timestamp 1731220528
transform 1 0 336 0 1 668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5484_6
timestamp 1731220528
transform 1 0 304 0 1 668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5483_6
timestamp 1731220528
transform 1 0 272 0 1 668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5482_6
timestamp 1731220528
transform 1 0 368 0 1 668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5481_6
timestamp 1731220528
transform 1 0 400 0 1 668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5480_6
timestamp 1731220528
transform 1 0 432 0 1 668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5479_6
timestamp 1731220528
transform 1 0 480 0 -1 668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5478_6
timestamp 1731220528
transform 1 0 448 0 -1 668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5477_6
timestamp 1731220528
transform 1 0 416 0 -1 668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5476_6
timestamp 1731220528
transform 1 0 384 0 -1 668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5475_6
timestamp 1731220528
transform 1 0 352 0 -1 668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5474_6
timestamp 1731220528
transform 1 0 320 0 -1 668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5473_6
timestamp 1731220528
transform 1 0 288 0 -1 668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5472_6
timestamp 1731220528
transform 1 0 464 0 1 588
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5471_6
timestamp 1731220528
transform 1 0 416 0 1 588
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5470_6
timestamp 1731220528
transform 1 0 360 0 1 588
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5469_6
timestamp 1731220528
transform 1 0 312 0 1 588
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5468_6
timestamp 1731220528
transform 1 0 272 0 1 588
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5467_6
timestamp 1731220528
transform 1 0 240 0 1 588
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5466_6
timestamp 1731220528
transform 1 0 480 0 -1 588
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5465_6
timestamp 1731220528
transform 1 0 400 0 -1 588
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5464_6
timestamp 1731220528
transform 1 0 328 0 -1 588
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5463_6
timestamp 1731220528
transform 1 0 264 0 -1 588
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5462_6
timestamp 1731220528
transform 1 0 208 0 -1 588
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5461_6
timestamp 1731220528
transform 1 0 160 0 -1 588
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5460_6
timestamp 1731220528
transform 1 0 320 0 1 504
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5459_6
timestamp 1731220528
transform 1 0 272 0 1 504
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5458_6
timestamp 1731220528
transform 1 0 224 0 1 504
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5457_6
timestamp 1731220528
transform 1 0 192 0 1 504
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5456_6
timestamp 1731220528
transform 1 0 160 0 1 504
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5455_6
timestamp 1731220528
transform 1 0 128 0 1 504
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5454_6
timestamp 1731220528
transform 1 0 232 0 -1 504
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5453_6
timestamp 1731220528
transform 1 0 192 0 -1 504
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5452_6
timestamp 1731220528
transform 1 0 160 0 -1 504
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5451_6
timestamp 1731220528
transform 1 0 128 0 -1 504
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5450_6
timestamp 1731220528
transform 1 0 280 0 -1 504
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5449_6
timestamp 1731220528
transform 1 0 248 0 1 424
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5448_6
timestamp 1731220528
transform 1 0 200 0 1 424
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5447_6
timestamp 1731220528
transform 1 0 144 0 1 424
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5446_6
timestamp 1731220528
transform 1 0 168 0 -1 424
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5445_6
timestamp 1731220528
transform 1 0 216 0 -1 424
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5444_6
timestamp 1731220528
transform 1 0 192 0 1 340
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5443_6
timestamp 1731220528
transform 1 0 160 0 1 340
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5442_6
timestamp 1731220528
transform 1 0 128 0 1 340
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5441_6
timestamp 1731220528
transform 1 0 160 0 -1 340
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5440_6
timestamp 1731220528
transform 1 0 128 0 -1 340
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5439_6
timestamp 1731220528
transform 1 0 128 0 1 260
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5438_6
timestamp 1731220528
transform 1 0 160 0 1 260
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5437_6
timestamp 1731220528
transform 1 0 224 0 1 260
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5436_6
timestamp 1731220528
transform 1 0 168 0 -1 256
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5435_6
timestamp 1731220528
transform 1 0 128 0 -1 256
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5434_6
timestamp 1731220528
transform 1 0 128 0 1 176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5433_6
timestamp 1731220528
transform 1 0 160 0 1 176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5432_6
timestamp 1731220528
transform 1 0 200 0 1 176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5431_6
timestamp 1731220528
transform 1 0 224 0 -1 176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5430_6
timestamp 1731220528
transform 1 0 168 0 -1 176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5429_6
timestamp 1731220528
transform 1 0 128 0 -1 176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5428_6
timestamp 1731220528
transform 1 0 128 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5427_6
timestamp 1731220528
transform 1 0 160 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5426_6
timestamp 1731220528
transform 1 0 192 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5425_6
timestamp 1731220528
transform 1 0 224 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5424_6
timestamp 1731220528
transform 1 0 256 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5423_6
timestamp 1731220528
transform 1 0 288 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5422_6
timestamp 1731220528
transform 1 0 320 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5421_6
timestamp 1731220528
transform 1 0 352 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5420_6
timestamp 1731220528
transform 1 0 384 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5419_6
timestamp 1731220528
transform 1 0 416 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5418_6
timestamp 1731220528
transform 1 0 392 0 -1 176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5417_6
timestamp 1731220528
transform 1 0 336 0 -1 176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5416_6
timestamp 1731220528
transform 1 0 280 0 -1 176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5415_6
timestamp 1731220528
transform 1 0 248 0 1 176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5414_6
timestamp 1731220528
transform 1 0 296 0 1 176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5413_6
timestamp 1731220528
transform 1 0 336 0 1 176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5412_6
timestamp 1731220528
transform 1 0 440 0 -1 256
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5411_6
timestamp 1731220528
transform 1 0 376 0 -1 256
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5410_6
timestamp 1731220528
transform 1 0 312 0 -1 256
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5409_6
timestamp 1731220528
transform 1 0 240 0 -1 256
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5408_6
timestamp 1731220528
transform 1 0 288 0 1 260
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5407_6
timestamp 1731220528
transform 1 0 360 0 1 260
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5406_6
timestamp 1731220528
transform 1 0 432 0 1 260
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5405_6
timestamp 1731220528
transform 1 0 384 0 -1 340
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5404_6
timestamp 1731220528
transform 1 0 320 0 -1 340
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5403_6
timestamp 1731220528
transform 1 0 256 0 -1 340
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5402_6
timestamp 1731220528
transform 1 0 200 0 -1 340
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5401_6
timestamp 1731220528
transform 1 0 232 0 1 340
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5400_6
timestamp 1731220528
transform 1 0 288 0 1 340
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5399_6
timestamp 1731220528
transform 1 0 344 0 1 340
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5398_6
timestamp 1731220528
transform 1 0 400 0 1 340
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5397_6
timestamp 1731220528
transform 1 0 408 0 -1 424
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5396_6
timestamp 1731220528
transform 1 0 360 0 -1 424
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5395_6
timestamp 1731220528
transform 1 0 312 0 -1 424
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5394_6
timestamp 1731220528
transform 1 0 264 0 -1 424
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5393_6
timestamp 1731220528
transform 1 0 304 0 1 424
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5392_6
timestamp 1731220528
transform 1 0 432 0 1 424
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5391_6
timestamp 1731220528
transform 1 0 360 0 1 424
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5390_6
timestamp 1731220528
transform 1 0 320 0 -1 504
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5389_6
timestamp 1731220528
transform 1 0 368 0 -1 504
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5388_6
timestamp 1731220528
transform 1 0 416 0 -1 504
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5387_6
timestamp 1731220528
transform 1 0 472 0 -1 504
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5386_6
timestamp 1731220528
transform 1 0 424 0 1 504
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5385_6
timestamp 1731220528
transform 1 0 368 0 1 504
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5384_6
timestamp 1731220528
transform 1 0 488 0 1 504
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5383_6
timestamp 1731220528
transform 1 0 552 0 1 504
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5382_6
timestamp 1731220528
transform 1 0 616 0 1 504
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5381_6
timestamp 1731220528
transform 1 0 608 0 -1 504
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5380_6
timestamp 1731220528
transform 1 0 536 0 -1 504
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5379_6
timestamp 1731220528
transform 1 0 688 0 -1 504
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5378_6
timestamp 1731220528
transform 1 0 672 0 1 424
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5377_6
timestamp 1731220528
transform 1 0 592 0 1 424
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5376_6
timestamp 1731220528
transform 1 0 512 0 1 424
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5375_6
timestamp 1731220528
transform 1 0 464 0 -1 424
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5374_6
timestamp 1731220528
transform 1 0 520 0 -1 424
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5373_6
timestamp 1731220528
transform 1 0 584 0 -1 424
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5372_6
timestamp 1731220528
transform 1 0 656 0 -1 424
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5371_6
timestamp 1731220528
transform 1 0 624 0 1 340
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5370_6
timestamp 1731220528
transform 1 0 568 0 1 340
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5369_6
timestamp 1731220528
transform 1 0 512 0 1 340
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5368_6
timestamp 1731220528
transform 1 0 456 0 1 340
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5367_6
timestamp 1731220528
transform 1 0 448 0 -1 340
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5366_6
timestamp 1731220528
transform 1 0 512 0 -1 340
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5365_6
timestamp 1731220528
transform 1 0 680 0 -1 340
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5364_6
timestamp 1731220528
transform 1 0 744 0 -1 340
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5363_6
timestamp 1731220528
transform 1 0 680 0 1 260
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5362_6
timestamp 1731220528
transform 1 0 624 0 1 260
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5361_6
timestamp 1731220528
transform 1 0 656 0 -1 256
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5360_6
timestamp 1731220528
transform 1 0 736 0 -1 256
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5359_6
timestamp 1731220528
transform 1 0 816 0 -1 256
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5358_6
timestamp 1731220528
transform 1 0 888 0 -1 256
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5357_6
timestamp 1731220528
transform 1 0 1024 0 1 260
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5356_6
timestamp 1731220528
transform 1 0 944 0 1 260
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5355_6
timestamp 1731220528
transform 1 0 872 0 1 260
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5354_6
timestamp 1731220528
transform 1 0 800 0 1 260
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5353_6
timestamp 1731220528
transform 1 0 736 0 1 260
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5352_6
timestamp 1731220528
transform 1 0 808 0 -1 340
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5351_6
timestamp 1731220528
transform 1 0 872 0 -1 340
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5350_6
timestamp 1731220528
transform 1 0 944 0 -1 340
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5349_6
timestamp 1731220528
transform 1 0 1024 0 -1 340
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5348_6
timestamp 1731220528
transform 1 0 1032 0 1 340
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5347_6
timestamp 1731220528
transform 1 0 976 0 1 340
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5346_6
timestamp 1731220528
transform 1 0 912 0 1 340
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5345_6
timestamp 1731220528
transform 1 0 848 0 1 340
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5344_6
timestamp 1731220528
transform 1 0 864 0 -1 424
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5343_6
timestamp 1731220528
transform 1 0 984 0 -1 424
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5342_6
timestamp 1731220528
transform 1 0 928 0 -1 424
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5341_6
timestamp 1731220528
transform 1 0 904 0 1 424
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5340_6
timestamp 1731220528
transform 1 0 832 0 1 424
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5339_6
timestamp 1731220528
transform 1 0 976 0 1 424
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5338_6
timestamp 1731220528
transform 1 0 1048 0 1 424
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5337_6
timestamp 1731220528
transform 1 0 1120 0 1 424
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5336_6
timestamp 1731220528
transform 1 0 1192 0 1 424
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5335_6
timestamp 1731220528
transform 1 0 1120 0 -1 424
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5334_6
timestamp 1731220528
transform 1 0 1080 0 -1 424
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5333_6
timestamp 1731220528
transform 1 0 1032 0 -1 424
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5332_6
timestamp 1731220528
transform 1 0 1088 0 1 340
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5331_6
timestamp 1731220528
transform 1 0 1144 0 1 340
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5330_6
timestamp 1731220528
transform 1 0 1104 0 -1 340
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5329_6
timestamp 1731220528
transform 1 0 1184 0 -1 340
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5328_6
timestamp 1731220528
transform 1 0 1264 0 -1 340
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5327_6
timestamp 1731220528
transform 1 0 1256 0 1 260
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5326_6
timestamp 1731220528
transform 1 0 1184 0 1 260
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5325_6
timestamp 1731220528
transform 1 0 1104 0 1 260
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5324_6
timestamp 1731220528
transform 1 0 1248 0 -1 256
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5323_6
timestamp 1731220528
transform 1 0 1192 0 -1 256
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5322_6
timestamp 1731220528
transform 1 0 1136 0 -1 256
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5321_6
timestamp 1731220528
transform 1 0 1080 0 -1 256
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5320_6
timestamp 1731220528
transform 1 0 1024 0 -1 256
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5319_6
timestamp 1731220528
transform 1 0 960 0 -1 256
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5318_6
timestamp 1731220528
transform 1 0 1208 0 1 176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5317_6
timestamp 1731220528
transform 1 0 1136 0 1 176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5316_6
timestamp 1731220528
transform 1 0 1064 0 1 176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5315_6
timestamp 1731220528
transform 1 0 992 0 1 176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5314_6
timestamp 1731220528
transform 1 0 920 0 1 176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5313_6
timestamp 1731220528
transform 1 0 848 0 1 176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5312_6
timestamp 1731220528
transform 1 0 1136 0 -1 176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5311_6
timestamp 1731220528
transform 1 0 1072 0 -1 176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5310_6
timestamp 1731220528
transform 1 0 1008 0 -1 176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5309_6
timestamp 1731220528
transform 1 0 944 0 -1 176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5308_6
timestamp 1731220528
transform 1 0 888 0 -1 176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5307_6
timestamp 1731220528
transform 1 0 824 0 -1 176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5306_6
timestamp 1731220528
transform 1 0 1136 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5305_6
timestamp 1731220528
transform 1 0 1096 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5304_6
timestamp 1731220528
transform 1 0 1056 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5303_6
timestamp 1731220528
transform 1 0 1008 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5302_6
timestamp 1731220528
transform 1 0 968 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5301_6
timestamp 1731220528
transform 1 0 928 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5300_6
timestamp 1731220528
transform 1 0 888 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5299_6
timestamp 1731220528
transform 1 0 856 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5298_6
timestamp 1731220528
transform 1 0 824 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5297_6
timestamp 1731220528
transform 1 0 792 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5296_6
timestamp 1731220528
transform 1 0 760 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5295_6
timestamp 1731220528
transform 1 0 728 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5294_6
timestamp 1731220528
transform 1 0 696 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5293_6
timestamp 1731220528
transform 1 0 664 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5292_6
timestamp 1731220528
transform 1 0 632 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5291_6
timestamp 1731220528
transform 1 0 600 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5290_6
timestamp 1731220528
transform 1 0 568 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5289_6
timestamp 1731220528
transform 1 0 536 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5288_6
timestamp 1731220528
transform 1 0 496 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5287_6
timestamp 1731220528
transform 1 0 456 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5286_6
timestamp 1731220528
transform 1 0 760 0 -1 176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5285_6
timestamp 1731220528
transform 1 0 696 0 -1 176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5284_6
timestamp 1731220528
transform 1 0 632 0 -1 176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5283_6
timestamp 1731220528
transform 1 0 568 0 -1 176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5282_6
timestamp 1731220528
transform 1 0 504 0 -1 176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5281_6
timestamp 1731220528
transform 1 0 448 0 -1 176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5280_6
timestamp 1731220528
transform 1 0 768 0 1 176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5279_6
timestamp 1731220528
transform 1 0 688 0 1 176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5278_6
timestamp 1731220528
transform 1 0 608 0 1 176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5277_6
timestamp 1731220528
transform 1 0 464 0 1 176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5276_6
timestamp 1731220528
transform 1 0 408 0 1 176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5275_6
timestamp 1731220528
transform 1 0 368 0 1 176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5274_6
timestamp 1731220528
transform 1 0 528 0 1 176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5273_6
timestamp 1731220528
transform 1 0 584 0 -1 256
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5272_6
timestamp 1731220528
transform 1 0 512 0 -1 256
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5271_6
timestamp 1731220528
transform 1 0 496 0 1 260
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5270_6
timestamp 1731220528
transform 1 0 560 0 1 260
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5269_6
timestamp 1731220528
transform 1 0 568 0 -1 340
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5268_6
timestamp 1731220528
transform 1 0 624 0 -1 340
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5267_6
timestamp 1731220528
transform 1 0 680 0 1 340
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5266_6
timestamp 1731220528
transform 1 0 792 0 1 340
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5265_6
timestamp 1731220528
transform 1 0 736 0 1 340
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5264_6
timestamp 1731220528
transform 1 0 728 0 -1 424
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5263_6
timestamp 1731220528
transform 1 0 800 0 -1 424
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5262_6
timestamp 1731220528
transform 1 0 752 0 1 424
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5261_6
timestamp 1731220528
transform 1 0 840 0 -1 504
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5260_6
timestamp 1731220528
transform 1 0 768 0 -1 504
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5259_6
timestamp 1731220528
transform 1 0 744 0 1 504
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5258_6
timestamp 1731220528
transform 1 0 680 0 1 504
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5257_6
timestamp 1731220528
transform 1 0 808 0 1 504
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5256_6
timestamp 1731220528
transform 1 0 760 0 -1 588
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5255_6
timestamp 1731220528
transform 1 0 696 0 -1 588
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5254_6
timestamp 1731220528
transform 1 0 624 0 -1 588
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5253_6
timestamp 1731220528
transform 1 0 552 0 -1 588
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5252_6
timestamp 1731220528
transform 1 0 768 0 1 588
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5251_6
timestamp 1731220528
transform 1 0 712 0 1 588
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5250_6
timestamp 1731220528
transform 1 0 656 0 1 588
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5249_6
timestamp 1731220528
transform 1 0 608 0 1 588
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5248_6
timestamp 1731220528
transform 1 0 560 0 1 588
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5247_6
timestamp 1731220528
transform 1 0 512 0 1 588
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5246_6
timestamp 1731220528
transform 1 0 728 0 -1 668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5245_6
timestamp 1731220528
transform 1 0 680 0 -1 668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5244_6
timestamp 1731220528
transform 1 0 632 0 -1 668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5243_6
timestamp 1731220528
transform 1 0 584 0 -1 668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5242_6
timestamp 1731220528
transform 1 0 544 0 -1 668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5241_6
timestamp 1731220528
transform 1 0 512 0 -1 668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5240_6
timestamp 1731220528
transform 1 0 696 0 1 668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5239_6
timestamp 1731220528
transform 1 0 640 0 1 668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5238_6
timestamp 1731220528
transform 1 0 584 0 1 668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5237_6
timestamp 1731220528
transform 1 0 536 0 1 668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5236_6
timestamp 1731220528
transform 1 0 496 0 1 668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5235_6
timestamp 1731220528
transform 1 0 464 0 1 668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5234_6
timestamp 1731220528
transform 1 0 432 0 -1 752
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5233_6
timestamp 1731220528
transform 1 0 480 0 -1 752
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5232_6
timestamp 1731220528
transform 1 0 536 0 -1 752
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5231_6
timestamp 1731220528
transform 1 0 600 0 -1 752
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5230_6
timestamp 1731220528
transform 1 0 664 0 -1 752
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5229_6
timestamp 1731220528
transform 1 0 608 0 1 752
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5228_6
timestamp 1731220528
transform 1 0 520 0 1 752
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5227_6
timestamp 1731220528
transform 1 0 472 0 -1 836
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5226_6
timestamp 1731220528
transform 1 0 536 0 -1 836
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5225_6
timestamp 1731220528
transform 1 0 600 0 -1 836
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5224_6
timestamp 1731220528
transform 1 0 592 0 1 836
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5223_6
timestamp 1731220528
transform 1 0 648 0 1 836
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5222_6
timestamp 1731220528
transform 1 0 640 0 -1 920
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5221_6
timestamp 1731220528
transform 1 0 696 0 -1 920
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5220_6
timestamp 1731220528
transform 1 0 744 0 -1 920
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5219_6
timestamp 1731220528
transform 1 0 720 0 1 924
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5218_6
timestamp 1731220528
transform 1 0 784 0 1 924
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5217_6
timestamp 1731220528
transform 1 0 752 0 -1 1004
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5216_6
timestamp 1731220528
transform 1 0 824 0 -1 1004
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5215_6
timestamp 1731220528
transform 1 0 872 0 1 1004
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5214_6
timestamp 1731220528
transform 1 0 792 0 1 1004
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5213_6
timestamp 1731220528
transform 1 0 728 0 -1 1088
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5212_6
timestamp 1731220528
transform 1 0 808 0 -1 1088
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5211_6
timestamp 1731220528
transform 1 0 888 0 -1 1088
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5210_6
timestamp 1731220528
transform 1 0 848 0 1 1092
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5209_6
timestamp 1731220528
transform 1 0 784 0 1 1092
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5208_6
timestamp 1731220528
transform 1 0 720 0 1 1092
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5207_6
timestamp 1731220528
transform 1 0 656 0 1 1092
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5206_6
timestamp 1731220528
transform 1 0 592 0 1 1092
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5205_6
timestamp 1731220528
transform 1 0 520 0 1 1092
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5204_6
timestamp 1731220528
transform 1 0 776 0 -1 1176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5203_6
timestamp 1731220528
transform 1 0 720 0 -1 1176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5202_6
timestamp 1731220528
transform 1 0 656 0 -1 1176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5201_6
timestamp 1731220528
transform 1 0 592 0 -1 1176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5200_6
timestamp 1731220528
transform 1 0 528 0 -1 1176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5199_6
timestamp 1731220528
transform 1 0 464 0 -1 1176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5198_6
timestamp 1731220528
transform 1 0 704 0 1 1180
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5197_6
timestamp 1731220528
transform 1 0 648 0 1 1180
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5196_6
timestamp 1731220528
transform 1 0 592 0 1 1180
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5195_6
timestamp 1731220528
transform 1 0 536 0 1 1180
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5194_6
timestamp 1731220528
transform 1 0 480 0 1 1180
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5193_6
timestamp 1731220528
transform 1 0 424 0 1 1180
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5192_6
timestamp 1731220528
transform 1 0 600 0 -1 1264
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5191_6
timestamp 1731220528
transform 1 0 544 0 -1 1264
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5190_6
timestamp 1731220528
transform 1 0 488 0 -1 1264
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5189_6
timestamp 1731220528
transform 1 0 432 0 -1 1264
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5188_6
timestamp 1731220528
transform 1 0 424 0 1 1264
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5187_6
timestamp 1731220528
transform 1 0 480 0 1 1264
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5186_6
timestamp 1731220528
transform 1 0 536 0 1 1264
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5185_6
timestamp 1731220528
transform 1 0 656 0 1 1264
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5184_6
timestamp 1731220528
transform 1 0 600 0 1 1264
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5183_6
timestamp 1731220528
transform 1 0 560 0 -1 1348
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5182_6
timestamp 1731220528
transform 1 0 504 0 -1 1348
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5181_6
timestamp 1731220528
transform 1 0 448 0 -1 1348
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5180_6
timestamp 1731220528
transform 1 0 624 0 -1 1348
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5179_6
timestamp 1731220528
transform 1 0 752 0 -1 1348
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5178_6
timestamp 1731220528
transform 1 0 688 0 -1 1348
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5177_6
timestamp 1731220528
transform 1 0 656 0 1 1348
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5176_6
timestamp 1731220528
transform 1 0 576 0 1 1348
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5175_6
timestamp 1731220528
transform 1 0 496 0 1 1348
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5174_6
timestamp 1731220528
transform 1 0 808 0 1 1348
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5173_6
timestamp 1731220528
transform 1 0 736 0 1 1348
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5172_6
timestamp 1731220528
transform 1 0 672 0 -1 1428
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5171_6
timestamp 1731220528
transform 1 0 592 0 -1 1428
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5170_6
timestamp 1731220528
transform 1 0 512 0 -1 1428
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5169_6
timestamp 1731220528
transform 1 0 752 0 -1 1428
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5168_6
timestamp 1731220528
transform 1 0 824 0 -1 1428
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5167_6
timestamp 1731220528
transform 1 0 896 0 -1 1428
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5166_6
timestamp 1731220528
transform 1 0 840 0 1 1432
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5165_6
timestamp 1731220528
transform 1 0 896 0 1 1432
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5164_6
timestamp 1731220528
transform 1 0 952 0 1 1432
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5163_6
timestamp 1731220528
transform 1 0 936 0 -1 1512
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5162_6
timestamp 1731220528
transform 1 0 912 0 1 1516
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5161_6
timestamp 1731220528
transform 1 0 1000 0 1 1516
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5160_6
timestamp 1731220528
transform 1 0 1088 0 1 1516
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5159_6
timestamp 1731220528
transform 1 0 1176 0 1 1516
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5158_6
timestamp 1731220528
transform 1 0 1192 0 -1 1596
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5157_6
timestamp 1731220528
transform 1 0 1112 0 -1 1596
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5156_6
timestamp 1731220528
transform 1 0 1032 0 -1 1596
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5155_6
timestamp 1731220528
transform 1 0 944 0 -1 1596
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5154_6
timestamp 1731220528
transform 1 0 1016 0 1 1596
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5153_6
timestamp 1731220528
transform 1 0 1096 0 1 1596
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5152_6
timestamp 1731220528
transform 1 0 1168 0 1 1596
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5151_6
timestamp 1731220528
transform 1 0 1096 0 -1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5150_6
timestamp 1731220528
transform 1 0 1024 0 -1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5149_6
timestamp 1731220528
transform 1 0 1168 0 -1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5148_6
timestamp 1731220528
transform 1 0 1168 0 1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5147_6
timestamp 1731220528
transform 1 0 1112 0 1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5146_6
timestamp 1731220528
transform 1 0 1056 0 1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5145_6
timestamp 1731220528
transform 1 0 1000 0 1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5144_6
timestamp 1731220528
transform 1 0 944 0 1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5143_6
timestamp 1731220528
transform 1 0 888 0 1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5142_6
timestamp 1731220528
transform 1 0 832 0 1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5141_6
timestamp 1731220528
transform 1 0 864 0 -1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5140_6
timestamp 1731220528
transform 1 0 944 0 -1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5139_6
timestamp 1731220528
transform 1 0 936 0 1 1596
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5138_6
timestamp 1731220528
transform 1 0 864 0 1 1596
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5137_6
timestamp 1731220528
transform 1 0 792 0 1 1596
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5136_6
timestamp 1731220528
transform 1 0 792 0 -1 1596
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5135_6
timestamp 1731220528
transform 1 0 864 0 -1 1596
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5134_6
timestamp 1731220528
transform 1 0 824 0 1 1516
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5133_6
timestamp 1731220528
transform 1 0 872 0 -1 1512
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5132_6
timestamp 1731220528
transform 1 0 808 0 -1 1512
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5131_6
timestamp 1731220528
transform 1 0 736 0 -1 1512
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5130_6
timestamp 1731220528
transform 1 0 776 0 1 1432
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5129_6
timestamp 1731220528
transform 1 0 712 0 1 1432
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5128_6
timestamp 1731220528
transform 1 0 656 0 1 1432
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5127_6
timestamp 1731220528
transform 1 0 592 0 1 1432
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5126_6
timestamp 1731220528
transform 1 0 520 0 1 1432
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5125_6
timestamp 1731220528
transform 1 0 520 0 -1 1512
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5124_6
timestamp 1731220528
transform 1 0 592 0 -1 1512
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5123_6
timestamp 1731220528
transform 1 0 664 0 -1 1512
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5122_6
timestamp 1731220528
transform 1 0 752 0 1 1516
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5121_6
timestamp 1731220528
transform 1 0 688 0 1 1516
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5120_6
timestamp 1731220528
transform 1 0 624 0 1 1516
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5119_6
timestamp 1731220528
transform 1 0 656 0 -1 1596
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5118_6
timestamp 1731220528
transform 1 0 720 0 -1 1596
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5117_6
timestamp 1731220528
transform 1 0 720 0 1 1596
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5116_6
timestamp 1731220528
transform 1 0 656 0 1 1596
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5115_6
timestamp 1731220528
transform 1 0 624 0 -1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5114_6
timestamp 1731220528
transform 1 0 704 0 -1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5113_6
timestamp 1731220528
transform 1 0 784 0 -1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5112_6
timestamp 1731220528
transform 1 0 776 0 1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5111_6
timestamp 1731220528
transform 1 0 720 0 1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5110_6
timestamp 1731220528
transform 1 0 656 0 1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5109_6
timestamp 1731220528
transform 1 0 600 0 1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5108_6
timestamp 1731220528
transform 1 0 544 0 1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5107_6
timestamp 1731220528
transform 1 0 496 0 1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5106_6
timestamp 1731220528
transform 1 0 480 0 -1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5105_6
timestamp 1731220528
transform 1 0 408 0 -1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5104_6
timestamp 1731220528
transform 1 0 552 0 -1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5103_6
timestamp 1731220528
transform 1 0 592 0 1 1596
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5102_6
timestamp 1731220528
transform 1 0 528 0 1 1596
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5101_6
timestamp 1731220528
transform 1 0 464 0 1 1596
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5100_6
timestamp 1731220528
transform 1 0 472 0 -1 1596
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_599_6
timestamp 1731220528
transform 1 0 528 0 -1 1596
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_598_6
timestamp 1731220528
transform 1 0 592 0 -1 1596
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_597_6
timestamp 1731220528
transform 1 0 560 0 1 1516
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_596_6
timestamp 1731220528
transform 1 0 504 0 1 1516
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_595_6
timestamp 1731220528
transform 1 0 448 0 1 1516
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_594_6
timestamp 1731220528
transform 1 0 400 0 1 1516
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_593_6
timestamp 1731220528
transform 1 0 352 0 1 1516
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_592_6
timestamp 1731220528
transform 1 0 328 0 -1 1596
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_591_6
timestamp 1731220528
transform 1 0 376 0 -1 1596
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_590_6
timestamp 1731220528
transform 1 0 424 0 -1 1596
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_589_6
timestamp 1731220528
transform 1 0 408 0 1 1596
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_588_6
timestamp 1731220528
transform 1 0 352 0 1 1596
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_587_6
timestamp 1731220528
transform 1 0 296 0 1 1596
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_586_6
timestamp 1731220528
transform 1 0 240 0 1 1596
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_585_6
timestamp 1731220528
transform 1 0 176 0 1 1596
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_584_6
timestamp 1731220528
transform 1 0 272 0 -1 1596
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_583_6
timestamp 1731220528
transform 1 0 216 0 -1 1596
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_582_6
timestamp 1731220528
transform 1 0 208 0 1 1516
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_581_6
timestamp 1731220528
transform 1 0 256 0 1 1516
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_580_6
timestamp 1731220528
transform 1 0 304 0 1 1516
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_579_6
timestamp 1731220528
transform 1 0 448 0 -1 1512
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_578_6
timestamp 1731220528
transform 1 0 368 0 -1 1512
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_577_6
timestamp 1731220528
transform 1 0 288 0 -1 1512
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_576_6
timestamp 1731220528
transform 1 0 216 0 -1 1512
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_575_6
timestamp 1731220528
transform 1 0 160 0 -1 1512
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_574_6
timestamp 1731220528
transform 1 0 216 0 1 1432
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_573_6
timestamp 1731220528
transform 1 0 288 0 1 1432
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_572_6
timestamp 1731220528
transform 1 0 368 0 1 1432
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_571_6
timestamp 1731220528
transform 1 0 448 0 1 1432
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_570_6
timestamp 1731220528
transform 1 0 432 0 -1 1428
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_569_6
timestamp 1731220528
transform 1 0 352 0 -1 1428
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_568_6
timestamp 1731220528
transform 1 0 280 0 -1 1428
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_567_6
timestamp 1731220528
transform 1 0 216 0 1 1348
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_566_6
timestamp 1731220528
transform 1 0 280 0 1 1348
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_565_6
timestamp 1731220528
transform 1 0 352 0 1 1348
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_564_6
timestamp 1731220528
transform 1 0 424 0 1 1348
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_563_6
timestamp 1731220528
transform 1 0 392 0 -1 1348
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_562_6
timestamp 1731220528
transform 1 0 344 0 -1 1348
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_561_6
timestamp 1731220528
transform 1 0 288 0 -1 1348
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_560_6
timestamp 1731220528
transform 1 0 232 0 -1 1348
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_559_6
timestamp 1731220528
transform 1 0 368 0 1 1264
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_558_6
timestamp 1731220528
transform 1 0 320 0 1 1264
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_557_6
timestamp 1731220528
transform 1 0 272 0 1 1264
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_556_6
timestamp 1731220528
transform 1 0 272 0 -1 1264
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_555_6
timestamp 1731220528
transform 1 0 320 0 -1 1264
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_554_6
timestamp 1731220528
transform 1 0 376 0 -1 1264
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_553_6
timestamp 1731220528
transform 1 0 376 0 1 1180
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_552_6
timestamp 1731220528
transform 1 0 328 0 1 1180
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_551_6
timestamp 1731220528
transform 1 0 272 0 1 1180
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_550_6
timestamp 1731220528
transform 1 0 280 0 -1 1176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_549_6
timestamp 1731220528
transform 1 0 344 0 -1 1176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_548_6
timestamp 1731220528
transform 1 0 408 0 -1 1176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_547_6
timestamp 1731220528
transform 1 0 456 0 1 1092
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_546_6
timestamp 1731220528
transform 1 0 392 0 1 1092
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_545_6
timestamp 1731220528
transform 1 0 328 0 1 1092
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_544_6
timestamp 1731220528
transform 1 0 272 0 -1 1088
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_543_6
timestamp 1731220528
transform 1 0 240 0 -1 1088
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_542_6
timestamp 1731220528
transform 1 0 208 0 -1 1088
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_541_6
timestamp 1731220528
transform 1 0 264 0 1 1092
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_540_6
timestamp 1731220528
transform 1 0 208 0 1 1092
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_539_6
timestamp 1731220528
transform 1 0 168 0 1 1092
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_538_6
timestamp 1731220528
transform 1 0 136 0 1 1092
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_537_6
timestamp 1731220528
transform 1 0 128 0 -1 1176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_536_6
timestamp 1731220528
transform 1 0 160 0 -1 1176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_535_6
timestamp 1731220528
transform 1 0 216 0 -1 1176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_534_6
timestamp 1731220528
transform 1 0 216 0 1 1180
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_533_6
timestamp 1731220528
transform 1 0 160 0 1 1180
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_532_6
timestamp 1731220528
transform 1 0 128 0 1 1180
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_531_6
timestamp 1731220528
transform 1 0 128 0 -1 1264
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_530_6
timestamp 1731220528
transform 1 0 160 0 -1 1264
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_529_6
timestamp 1731220528
transform 1 0 216 0 -1 1264
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_528_6
timestamp 1731220528
transform 1 0 224 0 1 1264
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_527_6
timestamp 1731220528
transform 1 0 176 0 1 1264
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_526_6
timestamp 1731220528
transform 1 0 128 0 1 1264
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_525_6
timestamp 1731220528
transform 1 0 128 0 -1 1348
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_524_6
timestamp 1731220528
transform 1 0 176 0 -1 1348
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_523_6
timestamp 1731220528
transform 1 0 160 0 1 1348
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_522_6
timestamp 1731220528
transform 1 0 128 0 1 1348
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_521_6
timestamp 1731220528
transform 1 0 208 0 -1 1428
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_520_6
timestamp 1731220528
transform 1 0 160 0 -1 1428
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_519_6
timestamp 1731220528
transform 1 0 128 0 -1 1428
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_518_6
timestamp 1731220528
transform 1 0 128 0 1 1432
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_517_6
timestamp 1731220528
transform 1 0 160 0 1 1432
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_516_6
timestamp 1731220528
transform 1 0 128 0 -1 1512
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_515_6
timestamp 1731220528
transform 1 0 128 0 1 1516
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_514_6
timestamp 1731220528
transform 1 0 160 0 1 1516
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_513_6
timestamp 1731220528
transform 1 0 160 0 -1 1596
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_512_6
timestamp 1731220528
transform 1 0 128 0 -1 1596
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_511_6
timestamp 1731220528
transform 1 0 128 0 1 1596
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_510_6
timestamp 1731220528
transform 1 0 128 0 -1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_59_6
timestamp 1731220528
transform 1 0 160 0 -1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_58_6
timestamp 1731220528
transform 1 0 208 0 -1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_57_6
timestamp 1731220528
transform 1 0 272 0 -1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_56_6
timestamp 1731220528
transform 1 0 336 0 -1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_55_6
timestamp 1731220528
transform 1 0 312 0 1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_54_6
timestamp 1731220528
transform 1 0 280 0 1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_53_6
timestamp 1731220528
transform 1 0 248 0 1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_52_6
timestamp 1731220528
transform 1 0 352 0 1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_51_6
timestamp 1731220528
transform 1 0 400 0 1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_50_6
timestamp 1731220528
transform 1 0 448 0 1 1676
box 8 7 28 34
<< end >>
