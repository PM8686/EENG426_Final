magic
tech sky130l
timestamp 1731220653
<< m2 >>
rect 134 2576 140 2577
rect 110 2573 116 2574
rect 110 2569 111 2573
rect 115 2569 116 2573
rect 134 2572 135 2576
rect 139 2572 140 2576
rect 134 2571 140 2572
rect 190 2576 196 2577
rect 190 2572 191 2576
rect 195 2572 196 2576
rect 190 2571 196 2572
rect 246 2576 252 2577
rect 246 2572 247 2576
rect 251 2572 252 2576
rect 246 2571 252 2572
rect 302 2576 308 2577
rect 302 2572 303 2576
rect 307 2572 308 2576
rect 302 2571 308 2572
rect 358 2576 364 2577
rect 358 2572 359 2576
rect 363 2572 364 2576
rect 358 2571 364 2572
rect 1286 2573 1292 2574
rect 110 2568 116 2569
rect 1286 2569 1287 2573
rect 1291 2569 1292 2573
rect 1286 2568 1292 2569
rect 110 2556 116 2557
rect 1286 2556 1292 2557
rect 110 2552 111 2556
rect 115 2552 116 2556
rect 110 2551 116 2552
rect 150 2555 156 2556
rect 150 2551 151 2555
rect 155 2551 156 2555
rect 150 2550 156 2551
rect 206 2555 212 2556
rect 206 2551 207 2555
rect 211 2551 212 2555
rect 206 2550 212 2551
rect 262 2555 268 2556
rect 262 2551 263 2555
rect 267 2551 268 2555
rect 262 2550 268 2551
rect 318 2555 324 2556
rect 318 2551 319 2555
rect 323 2551 324 2555
rect 318 2550 324 2551
rect 374 2555 380 2556
rect 374 2551 375 2555
rect 379 2551 380 2555
rect 1286 2552 1287 2556
rect 1291 2552 1292 2556
rect 1494 2556 1500 2557
rect 1286 2551 1292 2552
rect 1326 2553 1332 2554
rect 374 2550 380 2551
rect 1326 2549 1327 2553
rect 1331 2549 1332 2553
rect 1494 2552 1495 2556
rect 1499 2552 1500 2556
rect 1494 2551 1500 2552
rect 1550 2556 1556 2557
rect 1550 2552 1551 2556
rect 1555 2552 1556 2556
rect 1550 2551 1556 2552
rect 1606 2556 1612 2557
rect 1606 2552 1607 2556
rect 1611 2552 1612 2556
rect 1606 2551 1612 2552
rect 1662 2556 1668 2557
rect 1662 2552 1663 2556
rect 1667 2552 1668 2556
rect 1662 2551 1668 2552
rect 1718 2556 1724 2557
rect 1718 2552 1719 2556
rect 1723 2552 1724 2556
rect 1718 2551 1724 2552
rect 1774 2556 1780 2557
rect 1774 2552 1775 2556
rect 1779 2552 1780 2556
rect 1774 2551 1780 2552
rect 1830 2556 1836 2557
rect 1830 2552 1831 2556
rect 1835 2552 1836 2556
rect 1830 2551 1836 2552
rect 1886 2556 1892 2557
rect 1886 2552 1887 2556
rect 1891 2552 1892 2556
rect 1886 2551 1892 2552
rect 1942 2556 1948 2557
rect 1942 2552 1943 2556
rect 1947 2552 1948 2556
rect 1942 2551 1948 2552
rect 1998 2556 2004 2557
rect 1998 2552 1999 2556
rect 2003 2552 2004 2556
rect 1998 2551 2004 2552
rect 2054 2556 2060 2557
rect 2054 2552 2055 2556
rect 2059 2552 2060 2556
rect 2054 2551 2060 2552
rect 2110 2556 2116 2557
rect 2110 2552 2111 2556
rect 2115 2552 2116 2556
rect 2110 2551 2116 2552
rect 2166 2556 2172 2557
rect 2166 2552 2167 2556
rect 2171 2552 2172 2556
rect 2166 2551 2172 2552
rect 2502 2553 2508 2554
rect 1326 2548 1332 2549
rect 2502 2549 2503 2553
rect 2507 2549 2508 2553
rect 2502 2548 2508 2549
rect 1326 2536 1332 2537
rect 2502 2536 2508 2537
rect 1326 2532 1327 2536
rect 1331 2532 1332 2536
rect 1326 2531 1332 2532
rect 1510 2535 1516 2536
rect 1510 2531 1511 2535
rect 1515 2531 1516 2535
rect 1510 2530 1516 2531
rect 1566 2535 1572 2536
rect 1566 2531 1567 2535
rect 1571 2531 1572 2535
rect 1566 2530 1572 2531
rect 1622 2535 1628 2536
rect 1622 2531 1623 2535
rect 1627 2531 1628 2535
rect 1622 2530 1628 2531
rect 1678 2535 1684 2536
rect 1678 2531 1679 2535
rect 1683 2531 1684 2535
rect 1678 2530 1684 2531
rect 1734 2535 1740 2536
rect 1734 2531 1735 2535
rect 1739 2531 1740 2535
rect 1734 2530 1740 2531
rect 1790 2535 1796 2536
rect 1790 2531 1791 2535
rect 1795 2531 1796 2535
rect 1790 2530 1796 2531
rect 1846 2535 1852 2536
rect 1846 2531 1847 2535
rect 1851 2531 1852 2535
rect 1846 2530 1852 2531
rect 1902 2535 1908 2536
rect 1902 2531 1903 2535
rect 1907 2531 1908 2535
rect 1902 2530 1908 2531
rect 1958 2535 1964 2536
rect 1958 2531 1959 2535
rect 1963 2531 1964 2535
rect 1958 2530 1964 2531
rect 2014 2535 2020 2536
rect 2014 2531 2015 2535
rect 2019 2531 2020 2535
rect 2014 2530 2020 2531
rect 2070 2535 2076 2536
rect 2070 2531 2071 2535
rect 2075 2531 2076 2535
rect 2070 2530 2076 2531
rect 2126 2535 2132 2536
rect 2126 2531 2127 2535
rect 2131 2531 2132 2535
rect 2126 2530 2132 2531
rect 2182 2535 2188 2536
rect 2182 2531 2183 2535
rect 2187 2531 2188 2535
rect 2502 2532 2503 2536
rect 2507 2532 2508 2536
rect 2502 2531 2508 2532
rect 2182 2530 2188 2531
rect 222 2505 228 2506
rect 110 2504 116 2505
rect 110 2500 111 2504
rect 115 2500 116 2504
rect 222 2501 223 2505
rect 227 2501 228 2505
rect 222 2500 228 2501
rect 278 2505 284 2506
rect 278 2501 279 2505
rect 283 2501 284 2505
rect 278 2500 284 2501
rect 342 2505 348 2506
rect 342 2501 343 2505
rect 347 2501 348 2505
rect 342 2500 348 2501
rect 414 2505 420 2506
rect 414 2501 415 2505
rect 419 2501 420 2505
rect 414 2500 420 2501
rect 486 2505 492 2506
rect 486 2501 487 2505
rect 491 2501 492 2505
rect 486 2500 492 2501
rect 550 2505 556 2506
rect 550 2501 551 2505
rect 555 2501 556 2505
rect 550 2500 556 2501
rect 614 2505 620 2506
rect 614 2501 615 2505
rect 619 2501 620 2505
rect 614 2500 620 2501
rect 678 2505 684 2506
rect 678 2501 679 2505
rect 683 2501 684 2505
rect 678 2500 684 2501
rect 742 2505 748 2506
rect 742 2501 743 2505
rect 747 2501 748 2505
rect 742 2500 748 2501
rect 806 2505 812 2506
rect 806 2501 807 2505
rect 811 2501 812 2505
rect 806 2500 812 2501
rect 870 2505 876 2506
rect 870 2501 871 2505
rect 875 2501 876 2505
rect 870 2500 876 2501
rect 934 2505 940 2506
rect 934 2501 935 2505
rect 939 2501 940 2505
rect 934 2500 940 2501
rect 998 2505 1004 2506
rect 998 2501 999 2505
rect 1003 2501 1004 2505
rect 998 2500 1004 2501
rect 1062 2505 1068 2506
rect 1062 2501 1063 2505
rect 1067 2501 1068 2505
rect 1062 2500 1068 2501
rect 1286 2504 1292 2505
rect 1286 2500 1287 2504
rect 1291 2500 1292 2504
rect 110 2499 116 2500
rect 1286 2499 1292 2500
rect 110 2487 116 2488
rect 110 2483 111 2487
rect 115 2483 116 2487
rect 1286 2487 1292 2488
rect 110 2482 116 2483
rect 206 2484 212 2485
rect 206 2480 207 2484
rect 211 2480 212 2484
rect 206 2479 212 2480
rect 262 2484 268 2485
rect 262 2480 263 2484
rect 267 2480 268 2484
rect 262 2479 268 2480
rect 326 2484 332 2485
rect 326 2480 327 2484
rect 331 2480 332 2484
rect 326 2479 332 2480
rect 398 2484 404 2485
rect 398 2480 399 2484
rect 403 2480 404 2484
rect 398 2479 404 2480
rect 470 2484 476 2485
rect 470 2480 471 2484
rect 475 2480 476 2484
rect 470 2479 476 2480
rect 534 2484 540 2485
rect 534 2480 535 2484
rect 539 2480 540 2484
rect 534 2479 540 2480
rect 598 2484 604 2485
rect 598 2480 599 2484
rect 603 2480 604 2484
rect 598 2479 604 2480
rect 662 2484 668 2485
rect 662 2480 663 2484
rect 667 2480 668 2484
rect 662 2479 668 2480
rect 726 2484 732 2485
rect 726 2480 727 2484
rect 731 2480 732 2484
rect 726 2479 732 2480
rect 790 2484 796 2485
rect 790 2480 791 2484
rect 795 2480 796 2484
rect 790 2479 796 2480
rect 854 2484 860 2485
rect 854 2480 855 2484
rect 859 2480 860 2484
rect 854 2479 860 2480
rect 918 2484 924 2485
rect 918 2480 919 2484
rect 923 2480 924 2484
rect 918 2479 924 2480
rect 982 2484 988 2485
rect 982 2480 983 2484
rect 987 2480 988 2484
rect 982 2479 988 2480
rect 1046 2484 1052 2485
rect 1046 2480 1047 2484
rect 1051 2480 1052 2484
rect 1286 2483 1287 2487
rect 1291 2483 1292 2487
rect 1542 2485 1548 2486
rect 1286 2482 1292 2483
rect 1326 2484 1332 2485
rect 1046 2479 1052 2480
rect 1326 2480 1327 2484
rect 1331 2480 1332 2484
rect 1542 2481 1543 2485
rect 1547 2481 1548 2485
rect 1542 2480 1548 2481
rect 1606 2485 1612 2486
rect 1606 2481 1607 2485
rect 1611 2481 1612 2485
rect 1606 2480 1612 2481
rect 1678 2485 1684 2486
rect 1678 2481 1679 2485
rect 1683 2481 1684 2485
rect 1678 2480 1684 2481
rect 1750 2485 1756 2486
rect 1750 2481 1751 2485
rect 1755 2481 1756 2485
rect 1750 2480 1756 2481
rect 1822 2485 1828 2486
rect 1822 2481 1823 2485
rect 1827 2481 1828 2485
rect 1822 2480 1828 2481
rect 1894 2485 1900 2486
rect 1894 2481 1895 2485
rect 1899 2481 1900 2485
rect 1894 2480 1900 2481
rect 1966 2485 1972 2486
rect 1966 2481 1967 2485
rect 1971 2481 1972 2485
rect 1966 2480 1972 2481
rect 2038 2485 2044 2486
rect 2038 2481 2039 2485
rect 2043 2481 2044 2485
rect 2038 2480 2044 2481
rect 2110 2485 2116 2486
rect 2110 2481 2111 2485
rect 2115 2481 2116 2485
rect 2110 2480 2116 2481
rect 2182 2485 2188 2486
rect 2182 2481 2183 2485
rect 2187 2481 2188 2485
rect 2182 2480 2188 2481
rect 2502 2484 2508 2485
rect 2502 2480 2503 2484
rect 2507 2480 2508 2484
rect 1326 2479 1332 2480
rect 2502 2479 2508 2480
rect 1326 2467 1332 2468
rect 166 2464 172 2465
rect 110 2461 116 2462
rect 110 2457 111 2461
rect 115 2457 116 2461
rect 166 2460 167 2464
rect 171 2460 172 2464
rect 166 2459 172 2460
rect 222 2464 228 2465
rect 222 2460 223 2464
rect 227 2460 228 2464
rect 222 2459 228 2460
rect 278 2464 284 2465
rect 278 2460 279 2464
rect 283 2460 284 2464
rect 278 2459 284 2460
rect 334 2464 340 2465
rect 334 2460 335 2464
rect 339 2460 340 2464
rect 334 2459 340 2460
rect 390 2464 396 2465
rect 390 2460 391 2464
rect 395 2460 396 2464
rect 390 2459 396 2460
rect 446 2464 452 2465
rect 446 2460 447 2464
rect 451 2460 452 2464
rect 446 2459 452 2460
rect 502 2464 508 2465
rect 502 2460 503 2464
rect 507 2460 508 2464
rect 502 2459 508 2460
rect 558 2464 564 2465
rect 558 2460 559 2464
rect 563 2460 564 2464
rect 558 2459 564 2460
rect 614 2464 620 2465
rect 614 2460 615 2464
rect 619 2460 620 2464
rect 614 2459 620 2460
rect 670 2464 676 2465
rect 670 2460 671 2464
rect 675 2460 676 2464
rect 670 2459 676 2460
rect 726 2464 732 2465
rect 726 2460 727 2464
rect 731 2460 732 2464
rect 726 2459 732 2460
rect 782 2464 788 2465
rect 782 2460 783 2464
rect 787 2460 788 2464
rect 782 2459 788 2460
rect 838 2464 844 2465
rect 838 2460 839 2464
rect 843 2460 844 2464
rect 838 2459 844 2460
rect 894 2464 900 2465
rect 894 2460 895 2464
rect 899 2460 900 2464
rect 894 2459 900 2460
rect 950 2464 956 2465
rect 950 2460 951 2464
rect 955 2460 956 2464
rect 950 2459 956 2460
rect 1006 2464 1012 2465
rect 1006 2460 1007 2464
rect 1011 2460 1012 2464
rect 1006 2459 1012 2460
rect 1062 2464 1068 2465
rect 1062 2460 1063 2464
rect 1067 2460 1068 2464
rect 1326 2463 1327 2467
rect 1331 2463 1332 2467
rect 2502 2467 2508 2468
rect 1326 2462 1332 2463
rect 1526 2464 1532 2465
rect 1062 2459 1068 2460
rect 1286 2461 1292 2462
rect 110 2456 116 2457
rect 1286 2457 1287 2461
rect 1291 2457 1292 2461
rect 1526 2460 1527 2464
rect 1531 2460 1532 2464
rect 1526 2459 1532 2460
rect 1590 2464 1596 2465
rect 1590 2460 1591 2464
rect 1595 2460 1596 2464
rect 1590 2459 1596 2460
rect 1662 2464 1668 2465
rect 1662 2460 1663 2464
rect 1667 2460 1668 2464
rect 1662 2459 1668 2460
rect 1734 2464 1740 2465
rect 1734 2460 1735 2464
rect 1739 2460 1740 2464
rect 1734 2459 1740 2460
rect 1806 2464 1812 2465
rect 1806 2460 1807 2464
rect 1811 2460 1812 2464
rect 1806 2459 1812 2460
rect 1878 2464 1884 2465
rect 1878 2460 1879 2464
rect 1883 2460 1884 2464
rect 1878 2459 1884 2460
rect 1950 2464 1956 2465
rect 1950 2460 1951 2464
rect 1955 2460 1956 2464
rect 1950 2459 1956 2460
rect 2022 2464 2028 2465
rect 2022 2460 2023 2464
rect 2027 2460 2028 2464
rect 2022 2459 2028 2460
rect 2094 2464 2100 2465
rect 2094 2460 2095 2464
rect 2099 2460 2100 2464
rect 2094 2459 2100 2460
rect 2166 2464 2172 2465
rect 2166 2460 2167 2464
rect 2171 2460 2172 2464
rect 2502 2463 2503 2467
rect 2507 2463 2508 2467
rect 2502 2462 2508 2463
rect 2166 2459 2172 2460
rect 1286 2456 1292 2457
rect 1542 2448 1548 2449
rect 1326 2445 1332 2446
rect 110 2444 116 2445
rect 1286 2444 1292 2445
rect 110 2440 111 2444
rect 115 2440 116 2444
rect 110 2439 116 2440
rect 182 2443 188 2444
rect 182 2439 183 2443
rect 187 2439 188 2443
rect 182 2438 188 2439
rect 238 2443 244 2444
rect 238 2439 239 2443
rect 243 2439 244 2443
rect 238 2438 244 2439
rect 294 2443 300 2444
rect 294 2439 295 2443
rect 299 2439 300 2443
rect 294 2438 300 2439
rect 350 2443 356 2444
rect 350 2439 351 2443
rect 355 2439 356 2443
rect 350 2438 356 2439
rect 406 2443 412 2444
rect 406 2439 407 2443
rect 411 2439 412 2443
rect 406 2438 412 2439
rect 462 2443 468 2444
rect 462 2439 463 2443
rect 467 2439 468 2443
rect 462 2438 468 2439
rect 518 2443 524 2444
rect 518 2439 519 2443
rect 523 2439 524 2443
rect 518 2438 524 2439
rect 574 2443 580 2444
rect 574 2439 575 2443
rect 579 2439 580 2443
rect 574 2438 580 2439
rect 630 2443 636 2444
rect 630 2439 631 2443
rect 635 2439 636 2443
rect 630 2438 636 2439
rect 686 2443 692 2444
rect 686 2439 687 2443
rect 691 2439 692 2443
rect 686 2438 692 2439
rect 742 2443 748 2444
rect 742 2439 743 2443
rect 747 2439 748 2443
rect 742 2438 748 2439
rect 798 2443 804 2444
rect 798 2439 799 2443
rect 803 2439 804 2443
rect 798 2438 804 2439
rect 854 2443 860 2444
rect 854 2439 855 2443
rect 859 2439 860 2443
rect 854 2438 860 2439
rect 910 2443 916 2444
rect 910 2439 911 2443
rect 915 2439 916 2443
rect 910 2438 916 2439
rect 966 2443 972 2444
rect 966 2439 967 2443
rect 971 2439 972 2443
rect 966 2438 972 2439
rect 1022 2443 1028 2444
rect 1022 2439 1023 2443
rect 1027 2439 1028 2443
rect 1022 2438 1028 2439
rect 1078 2443 1084 2444
rect 1078 2439 1079 2443
rect 1083 2439 1084 2443
rect 1286 2440 1287 2444
rect 1291 2440 1292 2444
rect 1326 2441 1327 2445
rect 1331 2441 1332 2445
rect 1542 2444 1543 2448
rect 1547 2444 1548 2448
rect 1542 2443 1548 2444
rect 1606 2448 1612 2449
rect 1606 2444 1607 2448
rect 1611 2444 1612 2448
rect 1606 2443 1612 2444
rect 1670 2448 1676 2449
rect 1670 2444 1671 2448
rect 1675 2444 1676 2448
rect 1670 2443 1676 2444
rect 1742 2448 1748 2449
rect 1742 2444 1743 2448
rect 1747 2444 1748 2448
rect 1742 2443 1748 2444
rect 1814 2448 1820 2449
rect 1814 2444 1815 2448
rect 1819 2444 1820 2448
rect 1814 2443 1820 2444
rect 1878 2448 1884 2449
rect 1878 2444 1879 2448
rect 1883 2444 1884 2448
rect 1878 2443 1884 2444
rect 1950 2448 1956 2449
rect 1950 2444 1951 2448
rect 1955 2444 1956 2448
rect 1950 2443 1956 2444
rect 2022 2448 2028 2449
rect 2022 2444 2023 2448
rect 2027 2444 2028 2448
rect 2022 2443 2028 2444
rect 2094 2448 2100 2449
rect 2094 2444 2095 2448
rect 2099 2444 2100 2448
rect 2094 2443 2100 2444
rect 2166 2448 2172 2449
rect 2166 2444 2167 2448
rect 2171 2444 2172 2448
rect 2166 2443 2172 2444
rect 2502 2445 2508 2446
rect 1326 2440 1332 2441
rect 2502 2441 2503 2445
rect 2507 2441 2508 2445
rect 2502 2440 2508 2441
rect 1286 2439 1292 2440
rect 1078 2438 1084 2439
rect 1326 2428 1332 2429
rect 2502 2428 2508 2429
rect 1326 2424 1327 2428
rect 1331 2424 1332 2428
rect 1326 2423 1332 2424
rect 1558 2427 1564 2428
rect 1558 2423 1559 2427
rect 1563 2423 1564 2427
rect 1558 2422 1564 2423
rect 1622 2427 1628 2428
rect 1622 2423 1623 2427
rect 1627 2423 1628 2427
rect 1622 2422 1628 2423
rect 1686 2427 1692 2428
rect 1686 2423 1687 2427
rect 1691 2423 1692 2427
rect 1686 2422 1692 2423
rect 1758 2427 1764 2428
rect 1758 2423 1759 2427
rect 1763 2423 1764 2427
rect 1758 2422 1764 2423
rect 1830 2427 1836 2428
rect 1830 2423 1831 2427
rect 1835 2423 1836 2427
rect 1830 2422 1836 2423
rect 1894 2427 1900 2428
rect 1894 2423 1895 2427
rect 1899 2423 1900 2427
rect 1894 2422 1900 2423
rect 1966 2427 1972 2428
rect 1966 2423 1967 2427
rect 1971 2423 1972 2427
rect 1966 2422 1972 2423
rect 2038 2427 2044 2428
rect 2038 2423 2039 2427
rect 2043 2423 2044 2427
rect 2038 2422 2044 2423
rect 2110 2427 2116 2428
rect 2110 2423 2111 2427
rect 2115 2423 2116 2427
rect 2110 2422 2116 2423
rect 2182 2427 2188 2428
rect 2182 2423 2183 2427
rect 2187 2423 2188 2427
rect 2502 2424 2503 2428
rect 2507 2424 2508 2428
rect 2502 2423 2508 2424
rect 2182 2422 2188 2423
rect 518 2381 524 2382
rect 110 2380 116 2381
rect 110 2376 111 2380
rect 115 2376 116 2380
rect 518 2377 519 2381
rect 523 2377 524 2381
rect 518 2376 524 2377
rect 574 2381 580 2382
rect 574 2377 575 2381
rect 579 2377 580 2381
rect 574 2376 580 2377
rect 630 2381 636 2382
rect 630 2377 631 2381
rect 635 2377 636 2381
rect 630 2376 636 2377
rect 686 2381 692 2382
rect 686 2377 687 2381
rect 691 2377 692 2381
rect 686 2376 692 2377
rect 1286 2380 1292 2381
rect 1286 2376 1287 2380
rect 1291 2376 1292 2380
rect 110 2375 116 2376
rect 1286 2375 1292 2376
rect 1566 2373 1572 2374
rect 1326 2372 1332 2373
rect 1326 2368 1327 2372
rect 1331 2368 1332 2372
rect 1566 2369 1567 2373
rect 1571 2369 1572 2373
rect 1566 2368 1572 2369
rect 1622 2373 1628 2374
rect 1622 2369 1623 2373
rect 1627 2369 1628 2373
rect 1622 2368 1628 2369
rect 1678 2373 1684 2374
rect 1678 2369 1679 2373
rect 1683 2369 1684 2373
rect 1678 2368 1684 2369
rect 1734 2373 1740 2374
rect 1734 2369 1735 2373
rect 1739 2369 1740 2373
rect 1734 2368 1740 2369
rect 1790 2373 1796 2374
rect 1790 2369 1791 2373
rect 1795 2369 1796 2373
rect 1790 2368 1796 2369
rect 1854 2373 1860 2374
rect 1854 2369 1855 2373
rect 1859 2369 1860 2373
rect 1854 2368 1860 2369
rect 1918 2373 1924 2374
rect 1918 2369 1919 2373
rect 1923 2369 1924 2373
rect 1918 2368 1924 2369
rect 1982 2373 1988 2374
rect 1982 2369 1983 2373
rect 1987 2369 1988 2373
rect 1982 2368 1988 2369
rect 2046 2373 2052 2374
rect 2046 2369 2047 2373
rect 2051 2369 2052 2373
rect 2046 2368 2052 2369
rect 2110 2373 2116 2374
rect 2110 2369 2111 2373
rect 2115 2369 2116 2373
rect 2110 2368 2116 2369
rect 2502 2372 2508 2373
rect 2502 2368 2503 2372
rect 2507 2368 2508 2372
rect 1326 2367 1332 2368
rect 2502 2367 2508 2368
rect 110 2363 116 2364
rect 110 2359 111 2363
rect 115 2359 116 2363
rect 1286 2363 1292 2364
rect 110 2358 116 2359
rect 502 2360 508 2361
rect 502 2356 503 2360
rect 507 2356 508 2360
rect 502 2355 508 2356
rect 558 2360 564 2361
rect 558 2356 559 2360
rect 563 2356 564 2360
rect 558 2355 564 2356
rect 614 2360 620 2361
rect 614 2356 615 2360
rect 619 2356 620 2360
rect 614 2355 620 2356
rect 670 2360 676 2361
rect 670 2356 671 2360
rect 675 2356 676 2360
rect 1286 2359 1287 2363
rect 1291 2359 1292 2363
rect 1286 2358 1292 2359
rect 670 2355 676 2356
rect 1326 2355 1332 2356
rect 1326 2351 1327 2355
rect 1331 2351 1332 2355
rect 2502 2355 2508 2356
rect 1326 2350 1332 2351
rect 1550 2352 1556 2353
rect 1550 2348 1551 2352
rect 1555 2348 1556 2352
rect 1550 2347 1556 2348
rect 1606 2352 1612 2353
rect 1606 2348 1607 2352
rect 1611 2348 1612 2352
rect 1606 2347 1612 2348
rect 1662 2352 1668 2353
rect 1662 2348 1663 2352
rect 1667 2348 1668 2352
rect 1662 2347 1668 2348
rect 1718 2352 1724 2353
rect 1718 2348 1719 2352
rect 1723 2348 1724 2352
rect 1718 2347 1724 2348
rect 1774 2352 1780 2353
rect 1774 2348 1775 2352
rect 1779 2348 1780 2352
rect 1774 2347 1780 2348
rect 1838 2352 1844 2353
rect 1838 2348 1839 2352
rect 1843 2348 1844 2352
rect 1838 2347 1844 2348
rect 1902 2352 1908 2353
rect 1902 2348 1903 2352
rect 1907 2348 1908 2352
rect 1902 2347 1908 2348
rect 1966 2352 1972 2353
rect 1966 2348 1967 2352
rect 1971 2348 1972 2352
rect 1966 2347 1972 2348
rect 2030 2352 2036 2353
rect 2030 2348 2031 2352
rect 2035 2348 2036 2352
rect 2030 2347 2036 2348
rect 2094 2352 2100 2353
rect 2094 2348 2095 2352
rect 2099 2348 2100 2352
rect 2502 2351 2503 2355
rect 2507 2351 2508 2355
rect 2502 2350 2508 2351
rect 2094 2347 2100 2348
rect 318 2340 324 2341
rect 110 2337 116 2338
rect 110 2333 111 2337
rect 115 2333 116 2337
rect 318 2336 319 2340
rect 323 2336 324 2340
rect 318 2335 324 2336
rect 390 2340 396 2341
rect 390 2336 391 2340
rect 395 2336 396 2340
rect 390 2335 396 2336
rect 462 2340 468 2341
rect 462 2336 463 2340
rect 467 2336 468 2340
rect 462 2335 468 2336
rect 534 2340 540 2341
rect 534 2336 535 2340
rect 539 2336 540 2340
rect 534 2335 540 2336
rect 606 2340 612 2341
rect 606 2336 607 2340
rect 611 2336 612 2340
rect 606 2335 612 2336
rect 678 2340 684 2341
rect 678 2336 679 2340
rect 683 2336 684 2340
rect 678 2335 684 2336
rect 742 2340 748 2341
rect 742 2336 743 2340
rect 747 2336 748 2340
rect 742 2335 748 2336
rect 806 2340 812 2341
rect 806 2336 807 2340
rect 811 2336 812 2340
rect 806 2335 812 2336
rect 862 2340 868 2341
rect 862 2336 863 2340
rect 867 2336 868 2340
rect 862 2335 868 2336
rect 926 2340 932 2341
rect 926 2336 927 2340
rect 931 2336 932 2340
rect 926 2335 932 2336
rect 990 2340 996 2341
rect 990 2336 991 2340
rect 995 2336 996 2340
rect 990 2335 996 2336
rect 1054 2340 1060 2341
rect 1054 2336 1055 2340
rect 1059 2336 1060 2340
rect 1054 2335 1060 2336
rect 1110 2340 1116 2341
rect 1110 2336 1111 2340
rect 1115 2336 1116 2340
rect 1110 2335 1116 2336
rect 1166 2340 1172 2341
rect 1166 2336 1167 2340
rect 1171 2336 1172 2340
rect 1166 2335 1172 2336
rect 1222 2340 1228 2341
rect 1222 2336 1223 2340
rect 1227 2336 1228 2340
rect 1222 2335 1228 2336
rect 1286 2337 1292 2338
rect 110 2332 116 2333
rect 1286 2333 1287 2337
rect 1291 2333 1292 2337
rect 1286 2332 1292 2333
rect 1470 2332 1476 2333
rect 1326 2329 1332 2330
rect 1326 2325 1327 2329
rect 1331 2325 1332 2329
rect 1470 2328 1471 2332
rect 1475 2328 1476 2332
rect 1470 2327 1476 2328
rect 1534 2332 1540 2333
rect 1534 2328 1535 2332
rect 1539 2328 1540 2332
rect 1534 2327 1540 2328
rect 1606 2332 1612 2333
rect 1606 2328 1607 2332
rect 1611 2328 1612 2332
rect 1606 2327 1612 2328
rect 1686 2332 1692 2333
rect 1686 2328 1687 2332
rect 1691 2328 1692 2332
rect 1686 2327 1692 2328
rect 1758 2332 1764 2333
rect 1758 2328 1759 2332
rect 1763 2328 1764 2332
rect 1758 2327 1764 2328
rect 1830 2332 1836 2333
rect 1830 2328 1831 2332
rect 1835 2328 1836 2332
rect 1830 2327 1836 2328
rect 1902 2332 1908 2333
rect 1902 2328 1903 2332
rect 1907 2328 1908 2332
rect 1902 2327 1908 2328
rect 1982 2332 1988 2333
rect 1982 2328 1983 2332
rect 1987 2328 1988 2332
rect 1982 2327 1988 2328
rect 2062 2332 2068 2333
rect 2062 2328 2063 2332
rect 2067 2328 2068 2332
rect 2062 2327 2068 2328
rect 2142 2332 2148 2333
rect 2142 2328 2143 2332
rect 2147 2328 2148 2332
rect 2142 2327 2148 2328
rect 2502 2329 2508 2330
rect 1326 2324 1332 2325
rect 2502 2325 2503 2329
rect 2507 2325 2508 2329
rect 2502 2324 2508 2325
rect 110 2320 116 2321
rect 1286 2320 1292 2321
rect 110 2316 111 2320
rect 115 2316 116 2320
rect 110 2315 116 2316
rect 334 2319 340 2320
rect 334 2315 335 2319
rect 339 2315 340 2319
rect 334 2314 340 2315
rect 406 2319 412 2320
rect 406 2315 407 2319
rect 411 2315 412 2319
rect 406 2314 412 2315
rect 478 2319 484 2320
rect 478 2315 479 2319
rect 483 2315 484 2319
rect 478 2314 484 2315
rect 550 2319 556 2320
rect 550 2315 551 2319
rect 555 2315 556 2319
rect 550 2314 556 2315
rect 622 2319 628 2320
rect 622 2315 623 2319
rect 627 2315 628 2319
rect 622 2314 628 2315
rect 694 2319 700 2320
rect 694 2315 695 2319
rect 699 2315 700 2319
rect 694 2314 700 2315
rect 758 2319 764 2320
rect 758 2315 759 2319
rect 763 2315 764 2319
rect 758 2314 764 2315
rect 822 2319 828 2320
rect 822 2315 823 2319
rect 827 2315 828 2319
rect 822 2314 828 2315
rect 878 2319 884 2320
rect 878 2315 879 2319
rect 883 2315 884 2319
rect 878 2314 884 2315
rect 942 2319 948 2320
rect 942 2315 943 2319
rect 947 2315 948 2319
rect 942 2314 948 2315
rect 1006 2319 1012 2320
rect 1006 2315 1007 2319
rect 1011 2315 1012 2319
rect 1006 2314 1012 2315
rect 1070 2319 1076 2320
rect 1070 2315 1071 2319
rect 1075 2315 1076 2319
rect 1070 2314 1076 2315
rect 1126 2319 1132 2320
rect 1126 2315 1127 2319
rect 1131 2315 1132 2319
rect 1126 2314 1132 2315
rect 1182 2319 1188 2320
rect 1182 2315 1183 2319
rect 1187 2315 1188 2319
rect 1182 2314 1188 2315
rect 1238 2319 1244 2320
rect 1238 2315 1239 2319
rect 1243 2315 1244 2319
rect 1286 2316 1287 2320
rect 1291 2316 1292 2320
rect 1286 2315 1292 2316
rect 1238 2314 1244 2315
rect 1326 2312 1332 2313
rect 2502 2312 2508 2313
rect 1326 2308 1327 2312
rect 1331 2308 1332 2312
rect 1326 2307 1332 2308
rect 1486 2311 1492 2312
rect 1486 2307 1487 2311
rect 1491 2307 1492 2311
rect 1486 2306 1492 2307
rect 1550 2311 1556 2312
rect 1550 2307 1551 2311
rect 1555 2307 1556 2311
rect 1550 2306 1556 2307
rect 1622 2311 1628 2312
rect 1622 2307 1623 2311
rect 1627 2307 1628 2311
rect 1622 2306 1628 2307
rect 1702 2311 1708 2312
rect 1702 2307 1703 2311
rect 1707 2307 1708 2311
rect 1702 2306 1708 2307
rect 1774 2311 1780 2312
rect 1774 2307 1775 2311
rect 1779 2307 1780 2311
rect 1774 2306 1780 2307
rect 1846 2311 1852 2312
rect 1846 2307 1847 2311
rect 1851 2307 1852 2311
rect 1846 2306 1852 2307
rect 1918 2311 1924 2312
rect 1918 2307 1919 2311
rect 1923 2307 1924 2311
rect 1918 2306 1924 2307
rect 1998 2311 2004 2312
rect 1998 2307 1999 2311
rect 2003 2307 2004 2311
rect 1998 2306 2004 2307
rect 2078 2311 2084 2312
rect 2078 2307 2079 2311
rect 2083 2307 2084 2311
rect 2078 2306 2084 2307
rect 2158 2311 2164 2312
rect 2158 2307 2159 2311
rect 2163 2307 2164 2311
rect 2502 2308 2503 2312
rect 2507 2308 2508 2312
rect 2502 2307 2508 2308
rect 2158 2306 2164 2307
rect 174 2261 180 2262
rect 110 2260 116 2261
rect 110 2256 111 2260
rect 115 2256 116 2260
rect 174 2257 175 2261
rect 179 2257 180 2261
rect 174 2256 180 2257
rect 270 2261 276 2262
rect 270 2257 271 2261
rect 275 2257 276 2261
rect 270 2256 276 2257
rect 374 2261 380 2262
rect 374 2257 375 2261
rect 379 2257 380 2261
rect 374 2256 380 2257
rect 478 2261 484 2262
rect 478 2257 479 2261
rect 483 2257 484 2261
rect 478 2256 484 2257
rect 590 2261 596 2262
rect 590 2257 591 2261
rect 595 2257 596 2261
rect 590 2256 596 2257
rect 702 2261 708 2262
rect 702 2257 703 2261
rect 707 2257 708 2261
rect 702 2256 708 2257
rect 806 2261 812 2262
rect 806 2257 807 2261
rect 811 2257 812 2261
rect 806 2256 812 2257
rect 910 2261 916 2262
rect 910 2257 911 2261
rect 915 2257 916 2261
rect 910 2256 916 2257
rect 1014 2261 1020 2262
rect 1014 2257 1015 2261
rect 1019 2257 1020 2261
rect 1014 2256 1020 2257
rect 1126 2261 1132 2262
rect 1126 2257 1127 2261
rect 1131 2257 1132 2261
rect 1126 2256 1132 2257
rect 1238 2261 1244 2262
rect 1382 2261 1388 2262
rect 1238 2257 1239 2261
rect 1243 2257 1244 2261
rect 1238 2256 1244 2257
rect 1286 2260 1292 2261
rect 1286 2256 1287 2260
rect 1291 2256 1292 2260
rect 110 2255 116 2256
rect 1286 2255 1292 2256
rect 1326 2260 1332 2261
rect 1326 2256 1327 2260
rect 1331 2256 1332 2260
rect 1382 2257 1383 2261
rect 1387 2257 1388 2261
rect 1382 2256 1388 2257
rect 1478 2261 1484 2262
rect 1478 2257 1479 2261
rect 1483 2257 1484 2261
rect 1478 2256 1484 2257
rect 1582 2261 1588 2262
rect 1582 2257 1583 2261
rect 1587 2257 1588 2261
rect 1582 2256 1588 2257
rect 1686 2261 1692 2262
rect 1686 2257 1687 2261
rect 1691 2257 1692 2261
rect 1686 2256 1692 2257
rect 1790 2261 1796 2262
rect 1790 2257 1791 2261
rect 1795 2257 1796 2261
rect 1790 2256 1796 2257
rect 1902 2261 1908 2262
rect 1902 2257 1903 2261
rect 1907 2257 1908 2261
rect 1902 2256 1908 2257
rect 2014 2261 2020 2262
rect 2014 2257 2015 2261
rect 2019 2257 2020 2261
rect 2014 2256 2020 2257
rect 2126 2261 2132 2262
rect 2126 2257 2127 2261
rect 2131 2257 2132 2261
rect 2126 2256 2132 2257
rect 2238 2261 2244 2262
rect 2238 2257 2239 2261
rect 2243 2257 2244 2261
rect 2238 2256 2244 2257
rect 2502 2260 2508 2261
rect 2502 2256 2503 2260
rect 2507 2256 2508 2260
rect 1326 2255 1332 2256
rect 2502 2255 2508 2256
rect 110 2243 116 2244
rect 110 2239 111 2243
rect 115 2239 116 2243
rect 1286 2243 1292 2244
rect 110 2238 116 2239
rect 158 2240 164 2241
rect 158 2236 159 2240
rect 163 2236 164 2240
rect 158 2235 164 2236
rect 254 2240 260 2241
rect 254 2236 255 2240
rect 259 2236 260 2240
rect 254 2235 260 2236
rect 358 2240 364 2241
rect 358 2236 359 2240
rect 363 2236 364 2240
rect 358 2235 364 2236
rect 462 2240 468 2241
rect 462 2236 463 2240
rect 467 2236 468 2240
rect 462 2235 468 2236
rect 574 2240 580 2241
rect 574 2236 575 2240
rect 579 2236 580 2240
rect 574 2235 580 2236
rect 686 2240 692 2241
rect 686 2236 687 2240
rect 691 2236 692 2240
rect 686 2235 692 2236
rect 790 2240 796 2241
rect 790 2236 791 2240
rect 795 2236 796 2240
rect 790 2235 796 2236
rect 894 2240 900 2241
rect 894 2236 895 2240
rect 899 2236 900 2240
rect 894 2235 900 2236
rect 998 2240 1004 2241
rect 998 2236 999 2240
rect 1003 2236 1004 2240
rect 998 2235 1004 2236
rect 1110 2240 1116 2241
rect 1110 2236 1111 2240
rect 1115 2236 1116 2240
rect 1110 2235 1116 2236
rect 1222 2240 1228 2241
rect 1222 2236 1223 2240
rect 1227 2236 1228 2240
rect 1286 2239 1287 2243
rect 1291 2239 1292 2243
rect 1286 2238 1292 2239
rect 1326 2243 1332 2244
rect 1326 2239 1327 2243
rect 1331 2239 1332 2243
rect 2502 2243 2508 2244
rect 1326 2238 1332 2239
rect 1366 2240 1372 2241
rect 1222 2235 1228 2236
rect 1366 2236 1367 2240
rect 1371 2236 1372 2240
rect 1366 2235 1372 2236
rect 1462 2240 1468 2241
rect 1462 2236 1463 2240
rect 1467 2236 1468 2240
rect 1462 2235 1468 2236
rect 1566 2240 1572 2241
rect 1566 2236 1567 2240
rect 1571 2236 1572 2240
rect 1566 2235 1572 2236
rect 1670 2240 1676 2241
rect 1670 2236 1671 2240
rect 1675 2236 1676 2240
rect 1670 2235 1676 2236
rect 1774 2240 1780 2241
rect 1774 2236 1775 2240
rect 1779 2236 1780 2240
rect 1774 2235 1780 2236
rect 1886 2240 1892 2241
rect 1886 2236 1887 2240
rect 1891 2236 1892 2240
rect 1886 2235 1892 2236
rect 1998 2240 2004 2241
rect 1998 2236 1999 2240
rect 2003 2236 2004 2240
rect 1998 2235 2004 2236
rect 2110 2240 2116 2241
rect 2110 2236 2111 2240
rect 2115 2236 2116 2240
rect 2110 2235 2116 2236
rect 2222 2240 2228 2241
rect 2222 2236 2223 2240
rect 2227 2236 2228 2240
rect 2502 2239 2503 2243
rect 2507 2239 2508 2243
rect 2502 2238 2508 2239
rect 2222 2235 2228 2236
rect 142 2228 148 2229
rect 110 2225 116 2226
rect 110 2221 111 2225
rect 115 2221 116 2225
rect 142 2224 143 2228
rect 147 2224 148 2228
rect 142 2223 148 2224
rect 230 2228 236 2229
rect 230 2224 231 2228
rect 235 2224 236 2228
rect 230 2223 236 2224
rect 318 2228 324 2229
rect 318 2224 319 2228
rect 323 2224 324 2228
rect 318 2223 324 2224
rect 414 2228 420 2229
rect 414 2224 415 2228
rect 419 2224 420 2228
rect 414 2223 420 2224
rect 518 2228 524 2229
rect 518 2224 519 2228
rect 523 2224 524 2228
rect 518 2223 524 2224
rect 622 2228 628 2229
rect 622 2224 623 2228
rect 627 2224 628 2228
rect 622 2223 628 2224
rect 726 2228 732 2229
rect 726 2224 727 2228
rect 731 2224 732 2228
rect 726 2223 732 2224
rect 830 2228 836 2229
rect 830 2224 831 2228
rect 835 2224 836 2228
rect 830 2223 836 2224
rect 934 2228 940 2229
rect 934 2224 935 2228
rect 939 2224 940 2228
rect 934 2223 940 2224
rect 1038 2228 1044 2229
rect 1038 2224 1039 2228
rect 1043 2224 1044 2228
rect 1038 2223 1044 2224
rect 1142 2228 1148 2229
rect 1142 2224 1143 2228
rect 1147 2224 1148 2228
rect 1142 2223 1148 2224
rect 1222 2228 1228 2229
rect 1222 2224 1223 2228
rect 1227 2224 1228 2228
rect 1366 2228 1372 2229
rect 1222 2223 1228 2224
rect 1286 2225 1292 2226
rect 110 2220 116 2221
rect 1286 2221 1287 2225
rect 1291 2221 1292 2225
rect 1286 2220 1292 2221
rect 1326 2225 1332 2226
rect 1326 2221 1327 2225
rect 1331 2221 1332 2225
rect 1366 2224 1367 2228
rect 1371 2224 1372 2228
rect 1366 2223 1372 2224
rect 1486 2228 1492 2229
rect 1486 2224 1487 2228
rect 1491 2224 1492 2228
rect 1486 2223 1492 2224
rect 1606 2228 1612 2229
rect 1606 2224 1607 2228
rect 1611 2224 1612 2228
rect 1606 2223 1612 2224
rect 1718 2228 1724 2229
rect 1718 2224 1719 2228
rect 1723 2224 1724 2228
rect 1718 2223 1724 2224
rect 1814 2228 1820 2229
rect 1814 2224 1815 2228
rect 1819 2224 1820 2228
rect 1814 2223 1820 2224
rect 1902 2228 1908 2229
rect 1902 2224 1903 2228
rect 1907 2224 1908 2228
rect 1902 2223 1908 2224
rect 1982 2228 1988 2229
rect 1982 2224 1983 2228
rect 1987 2224 1988 2228
rect 1982 2223 1988 2224
rect 2054 2228 2060 2229
rect 2054 2224 2055 2228
rect 2059 2224 2060 2228
rect 2054 2223 2060 2224
rect 2126 2228 2132 2229
rect 2126 2224 2127 2228
rect 2131 2224 2132 2228
rect 2126 2223 2132 2224
rect 2190 2228 2196 2229
rect 2190 2224 2191 2228
rect 2195 2224 2196 2228
rect 2190 2223 2196 2224
rect 2254 2228 2260 2229
rect 2254 2224 2255 2228
rect 2259 2224 2260 2228
rect 2254 2223 2260 2224
rect 2318 2228 2324 2229
rect 2318 2224 2319 2228
rect 2323 2224 2324 2228
rect 2318 2223 2324 2224
rect 2382 2228 2388 2229
rect 2382 2224 2383 2228
rect 2387 2224 2388 2228
rect 2382 2223 2388 2224
rect 2438 2228 2444 2229
rect 2438 2224 2439 2228
rect 2443 2224 2444 2228
rect 2438 2223 2444 2224
rect 2502 2225 2508 2226
rect 1326 2220 1332 2221
rect 2502 2221 2503 2225
rect 2507 2221 2508 2225
rect 2502 2220 2508 2221
rect 110 2208 116 2209
rect 1286 2208 1292 2209
rect 110 2204 111 2208
rect 115 2204 116 2208
rect 110 2203 116 2204
rect 158 2207 164 2208
rect 158 2203 159 2207
rect 163 2203 164 2207
rect 158 2202 164 2203
rect 246 2207 252 2208
rect 246 2203 247 2207
rect 251 2203 252 2207
rect 246 2202 252 2203
rect 334 2207 340 2208
rect 334 2203 335 2207
rect 339 2203 340 2207
rect 334 2202 340 2203
rect 430 2207 436 2208
rect 430 2203 431 2207
rect 435 2203 436 2207
rect 430 2202 436 2203
rect 534 2207 540 2208
rect 534 2203 535 2207
rect 539 2203 540 2207
rect 534 2202 540 2203
rect 638 2207 644 2208
rect 638 2203 639 2207
rect 643 2203 644 2207
rect 638 2202 644 2203
rect 742 2207 748 2208
rect 742 2203 743 2207
rect 747 2203 748 2207
rect 742 2202 748 2203
rect 846 2207 852 2208
rect 846 2203 847 2207
rect 851 2203 852 2207
rect 846 2202 852 2203
rect 950 2207 956 2208
rect 950 2203 951 2207
rect 955 2203 956 2207
rect 950 2202 956 2203
rect 1054 2207 1060 2208
rect 1054 2203 1055 2207
rect 1059 2203 1060 2207
rect 1054 2202 1060 2203
rect 1158 2207 1164 2208
rect 1158 2203 1159 2207
rect 1163 2203 1164 2207
rect 1158 2202 1164 2203
rect 1238 2207 1244 2208
rect 1238 2203 1239 2207
rect 1243 2203 1244 2207
rect 1286 2204 1287 2208
rect 1291 2204 1292 2208
rect 1286 2203 1292 2204
rect 1326 2208 1332 2209
rect 2502 2208 2508 2209
rect 1326 2204 1327 2208
rect 1331 2204 1332 2208
rect 1326 2203 1332 2204
rect 1382 2207 1388 2208
rect 1382 2203 1383 2207
rect 1387 2203 1388 2207
rect 1238 2202 1244 2203
rect 1382 2202 1388 2203
rect 1502 2207 1508 2208
rect 1502 2203 1503 2207
rect 1507 2203 1508 2207
rect 1502 2202 1508 2203
rect 1622 2207 1628 2208
rect 1622 2203 1623 2207
rect 1627 2203 1628 2207
rect 1622 2202 1628 2203
rect 1734 2207 1740 2208
rect 1734 2203 1735 2207
rect 1739 2203 1740 2207
rect 1734 2202 1740 2203
rect 1830 2207 1836 2208
rect 1830 2203 1831 2207
rect 1835 2203 1836 2207
rect 1830 2202 1836 2203
rect 1918 2207 1924 2208
rect 1918 2203 1919 2207
rect 1923 2203 1924 2207
rect 1918 2202 1924 2203
rect 1998 2207 2004 2208
rect 1998 2203 1999 2207
rect 2003 2203 2004 2207
rect 1998 2202 2004 2203
rect 2070 2207 2076 2208
rect 2070 2203 2071 2207
rect 2075 2203 2076 2207
rect 2070 2202 2076 2203
rect 2142 2207 2148 2208
rect 2142 2203 2143 2207
rect 2147 2203 2148 2207
rect 2142 2202 2148 2203
rect 2206 2207 2212 2208
rect 2206 2203 2207 2207
rect 2211 2203 2212 2207
rect 2206 2202 2212 2203
rect 2270 2207 2276 2208
rect 2270 2203 2271 2207
rect 2275 2203 2276 2207
rect 2270 2202 2276 2203
rect 2334 2207 2340 2208
rect 2334 2203 2335 2207
rect 2339 2203 2340 2207
rect 2334 2202 2340 2203
rect 2398 2207 2404 2208
rect 2398 2203 2399 2207
rect 2403 2203 2404 2207
rect 2398 2202 2404 2203
rect 2454 2207 2460 2208
rect 2454 2203 2455 2207
rect 2459 2203 2460 2207
rect 2502 2204 2503 2208
rect 2507 2204 2508 2208
rect 2502 2203 2508 2204
rect 2454 2202 2460 2203
rect 254 2157 260 2158
rect 110 2156 116 2157
rect 110 2152 111 2156
rect 115 2152 116 2156
rect 254 2153 255 2157
rect 259 2153 260 2157
rect 254 2152 260 2153
rect 350 2157 356 2158
rect 350 2153 351 2157
rect 355 2153 356 2157
rect 350 2152 356 2153
rect 454 2157 460 2158
rect 454 2153 455 2157
rect 459 2153 460 2157
rect 454 2152 460 2153
rect 558 2157 564 2158
rect 558 2153 559 2157
rect 563 2153 564 2157
rect 558 2152 564 2153
rect 662 2157 668 2158
rect 662 2153 663 2157
rect 667 2153 668 2157
rect 662 2152 668 2153
rect 766 2157 772 2158
rect 766 2153 767 2157
rect 771 2153 772 2157
rect 766 2152 772 2153
rect 862 2157 868 2158
rect 862 2153 863 2157
rect 867 2153 868 2157
rect 862 2152 868 2153
rect 958 2157 964 2158
rect 958 2153 959 2157
rect 963 2153 964 2157
rect 958 2152 964 2153
rect 1054 2157 1060 2158
rect 1054 2153 1055 2157
rect 1059 2153 1060 2157
rect 1054 2152 1060 2153
rect 1158 2157 1164 2158
rect 1158 2153 1159 2157
rect 1163 2153 1164 2157
rect 1158 2152 1164 2153
rect 1238 2157 1244 2158
rect 1238 2153 1239 2157
rect 1243 2153 1244 2157
rect 1238 2152 1244 2153
rect 1286 2156 1292 2157
rect 1286 2152 1287 2156
rect 1291 2152 1292 2156
rect 110 2151 116 2152
rect 1286 2151 1292 2152
rect 110 2139 116 2140
rect 110 2135 111 2139
rect 115 2135 116 2139
rect 1286 2139 1292 2140
rect 110 2134 116 2135
rect 238 2136 244 2137
rect 238 2132 239 2136
rect 243 2132 244 2136
rect 238 2131 244 2132
rect 334 2136 340 2137
rect 334 2132 335 2136
rect 339 2132 340 2136
rect 334 2131 340 2132
rect 438 2136 444 2137
rect 438 2132 439 2136
rect 443 2132 444 2136
rect 438 2131 444 2132
rect 542 2136 548 2137
rect 542 2132 543 2136
rect 547 2132 548 2136
rect 542 2131 548 2132
rect 646 2136 652 2137
rect 646 2132 647 2136
rect 651 2132 652 2136
rect 646 2131 652 2132
rect 750 2136 756 2137
rect 750 2132 751 2136
rect 755 2132 756 2136
rect 750 2131 756 2132
rect 846 2136 852 2137
rect 846 2132 847 2136
rect 851 2132 852 2136
rect 846 2131 852 2132
rect 942 2136 948 2137
rect 942 2132 943 2136
rect 947 2132 948 2136
rect 942 2131 948 2132
rect 1038 2136 1044 2137
rect 1038 2132 1039 2136
rect 1043 2132 1044 2136
rect 1038 2131 1044 2132
rect 1142 2136 1148 2137
rect 1142 2132 1143 2136
rect 1147 2132 1148 2136
rect 1142 2131 1148 2132
rect 1222 2136 1228 2137
rect 1222 2132 1223 2136
rect 1227 2132 1228 2136
rect 1286 2135 1287 2139
rect 1291 2135 1292 2139
rect 1406 2137 1412 2138
rect 1286 2134 1292 2135
rect 1326 2136 1332 2137
rect 1222 2131 1228 2132
rect 1326 2132 1327 2136
rect 1331 2132 1332 2136
rect 1406 2133 1407 2137
rect 1411 2133 1412 2137
rect 1406 2132 1412 2133
rect 1622 2137 1628 2138
rect 1622 2133 1623 2137
rect 1627 2133 1628 2137
rect 1622 2132 1628 2133
rect 1814 2137 1820 2138
rect 1814 2133 1815 2137
rect 1819 2133 1820 2137
rect 1814 2132 1820 2133
rect 1990 2137 1996 2138
rect 1990 2133 1991 2137
rect 1995 2133 1996 2137
rect 1990 2132 1996 2133
rect 2158 2137 2164 2138
rect 2158 2133 2159 2137
rect 2163 2133 2164 2137
rect 2158 2132 2164 2133
rect 2318 2137 2324 2138
rect 2318 2133 2319 2137
rect 2323 2133 2324 2137
rect 2318 2132 2324 2133
rect 2454 2137 2460 2138
rect 2454 2133 2455 2137
rect 2459 2133 2460 2137
rect 2454 2132 2460 2133
rect 2502 2136 2508 2137
rect 2502 2132 2503 2136
rect 2507 2132 2508 2136
rect 1326 2131 1332 2132
rect 2502 2131 2508 2132
rect 302 2124 308 2125
rect 110 2121 116 2122
rect 110 2117 111 2121
rect 115 2117 116 2121
rect 302 2120 303 2124
rect 307 2120 308 2124
rect 302 2119 308 2120
rect 358 2124 364 2125
rect 358 2120 359 2124
rect 363 2120 364 2124
rect 358 2119 364 2120
rect 422 2124 428 2125
rect 422 2120 423 2124
rect 427 2120 428 2124
rect 422 2119 428 2120
rect 486 2124 492 2125
rect 486 2120 487 2124
rect 491 2120 492 2124
rect 486 2119 492 2120
rect 558 2124 564 2125
rect 558 2120 559 2124
rect 563 2120 564 2124
rect 558 2119 564 2120
rect 630 2124 636 2125
rect 630 2120 631 2124
rect 635 2120 636 2124
rect 630 2119 636 2120
rect 710 2124 716 2125
rect 710 2120 711 2124
rect 715 2120 716 2124
rect 710 2119 716 2120
rect 798 2124 804 2125
rect 798 2120 799 2124
rect 803 2120 804 2124
rect 798 2119 804 2120
rect 886 2124 892 2125
rect 886 2120 887 2124
rect 891 2120 892 2124
rect 886 2119 892 2120
rect 974 2124 980 2125
rect 974 2120 975 2124
rect 979 2120 980 2124
rect 974 2119 980 2120
rect 1062 2124 1068 2125
rect 1062 2120 1063 2124
rect 1067 2120 1068 2124
rect 1062 2119 1068 2120
rect 1150 2124 1156 2125
rect 1150 2120 1151 2124
rect 1155 2120 1156 2124
rect 1150 2119 1156 2120
rect 1222 2124 1228 2125
rect 1222 2120 1223 2124
rect 1227 2120 1228 2124
rect 1222 2119 1228 2120
rect 1286 2121 1292 2122
rect 110 2116 116 2117
rect 1286 2117 1287 2121
rect 1291 2117 1292 2121
rect 1286 2116 1292 2117
rect 1326 2119 1332 2120
rect 1326 2115 1327 2119
rect 1331 2115 1332 2119
rect 2502 2119 2508 2120
rect 1326 2114 1332 2115
rect 1390 2116 1396 2117
rect 1390 2112 1391 2116
rect 1395 2112 1396 2116
rect 1390 2111 1396 2112
rect 1606 2116 1612 2117
rect 1606 2112 1607 2116
rect 1611 2112 1612 2116
rect 1606 2111 1612 2112
rect 1798 2116 1804 2117
rect 1798 2112 1799 2116
rect 1803 2112 1804 2116
rect 1798 2111 1804 2112
rect 1974 2116 1980 2117
rect 1974 2112 1975 2116
rect 1979 2112 1980 2116
rect 1974 2111 1980 2112
rect 2142 2116 2148 2117
rect 2142 2112 2143 2116
rect 2147 2112 2148 2116
rect 2142 2111 2148 2112
rect 2302 2116 2308 2117
rect 2302 2112 2303 2116
rect 2307 2112 2308 2116
rect 2302 2111 2308 2112
rect 2438 2116 2444 2117
rect 2438 2112 2439 2116
rect 2443 2112 2444 2116
rect 2502 2115 2503 2119
rect 2507 2115 2508 2119
rect 2502 2114 2508 2115
rect 2438 2111 2444 2112
rect 110 2104 116 2105
rect 1286 2104 1292 2105
rect 110 2100 111 2104
rect 115 2100 116 2104
rect 110 2099 116 2100
rect 318 2103 324 2104
rect 318 2099 319 2103
rect 323 2099 324 2103
rect 318 2098 324 2099
rect 374 2103 380 2104
rect 374 2099 375 2103
rect 379 2099 380 2103
rect 374 2098 380 2099
rect 438 2103 444 2104
rect 438 2099 439 2103
rect 443 2099 444 2103
rect 438 2098 444 2099
rect 502 2103 508 2104
rect 502 2099 503 2103
rect 507 2099 508 2103
rect 502 2098 508 2099
rect 574 2103 580 2104
rect 574 2099 575 2103
rect 579 2099 580 2103
rect 574 2098 580 2099
rect 646 2103 652 2104
rect 646 2099 647 2103
rect 651 2099 652 2103
rect 646 2098 652 2099
rect 726 2103 732 2104
rect 726 2099 727 2103
rect 731 2099 732 2103
rect 726 2098 732 2099
rect 814 2103 820 2104
rect 814 2099 815 2103
rect 819 2099 820 2103
rect 814 2098 820 2099
rect 902 2103 908 2104
rect 902 2099 903 2103
rect 907 2099 908 2103
rect 902 2098 908 2099
rect 990 2103 996 2104
rect 990 2099 991 2103
rect 995 2099 996 2103
rect 990 2098 996 2099
rect 1078 2103 1084 2104
rect 1078 2099 1079 2103
rect 1083 2099 1084 2103
rect 1078 2098 1084 2099
rect 1166 2103 1172 2104
rect 1166 2099 1167 2103
rect 1171 2099 1172 2103
rect 1166 2098 1172 2099
rect 1238 2103 1244 2104
rect 1238 2099 1239 2103
rect 1243 2099 1244 2103
rect 1286 2100 1287 2104
rect 1291 2100 1292 2104
rect 1382 2104 1388 2105
rect 1286 2099 1292 2100
rect 1326 2101 1332 2102
rect 1238 2098 1244 2099
rect 1326 2097 1327 2101
rect 1331 2097 1332 2101
rect 1382 2100 1383 2104
rect 1387 2100 1388 2104
rect 1382 2099 1388 2100
rect 1550 2104 1556 2105
rect 1550 2100 1551 2104
rect 1555 2100 1556 2104
rect 1550 2099 1556 2100
rect 1710 2104 1716 2105
rect 1710 2100 1711 2104
rect 1715 2100 1716 2104
rect 1710 2099 1716 2100
rect 1854 2104 1860 2105
rect 1854 2100 1855 2104
rect 1859 2100 1860 2104
rect 1854 2099 1860 2100
rect 1990 2104 1996 2105
rect 1990 2100 1991 2104
rect 1995 2100 1996 2104
rect 1990 2099 1996 2100
rect 2118 2104 2124 2105
rect 2118 2100 2119 2104
rect 2123 2100 2124 2104
rect 2118 2099 2124 2100
rect 2238 2104 2244 2105
rect 2238 2100 2239 2104
rect 2243 2100 2244 2104
rect 2238 2099 2244 2100
rect 2366 2104 2372 2105
rect 2366 2100 2367 2104
rect 2371 2100 2372 2104
rect 2366 2099 2372 2100
rect 2502 2101 2508 2102
rect 1326 2096 1332 2097
rect 2502 2097 2503 2101
rect 2507 2097 2508 2101
rect 2502 2096 2508 2097
rect 1326 2084 1332 2085
rect 2502 2084 2508 2085
rect 1326 2080 1327 2084
rect 1331 2080 1332 2084
rect 1326 2079 1332 2080
rect 1398 2083 1404 2084
rect 1398 2079 1399 2083
rect 1403 2079 1404 2083
rect 1398 2078 1404 2079
rect 1566 2083 1572 2084
rect 1566 2079 1567 2083
rect 1571 2079 1572 2083
rect 1566 2078 1572 2079
rect 1726 2083 1732 2084
rect 1726 2079 1727 2083
rect 1731 2079 1732 2083
rect 1726 2078 1732 2079
rect 1870 2083 1876 2084
rect 1870 2079 1871 2083
rect 1875 2079 1876 2083
rect 1870 2078 1876 2079
rect 2006 2083 2012 2084
rect 2006 2079 2007 2083
rect 2011 2079 2012 2083
rect 2006 2078 2012 2079
rect 2134 2083 2140 2084
rect 2134 2079 2135 2083
rect 2139 2079 2140 2083
rect 2134 2078 2140 2079
rect 2254 2083 2260 2084
rect 2254 2079 2255 2083
rect 2259 2079 2260 2083
rect 2254 2078 2260 2079
rect 2382 2083 2388 2084
rect 2382 2079 2383 2083
rect 2387 2079 2388 2083
rect 2502 2080 2503 2084
rect 2507 2080 2508 2084
rect 2502 2079 2508 2080
rect 2382 2078 2388 2079
rect 398 2049 404 2050
rect 110 2048 116 2049
rect 110 2044 111 2048
rect 115 2044 116 2048
rect 398 2045 399 2049
rect 403 2045 404 2049
rect 398 2044 404 2045
rect 454 2049 460 2050
rect 454 2045 455 2049
rect 459 2045 460 2049
rect 454 2044 460 2045
rect 510 2049 516 2050
rect 510 2045 511 2049
rect 515 2045 516 2049
rect 510 2044 516 2045
rect 574 2049 580 2050
rect 574 2045 575 2049
rect 579 2045 580 2049
rect 574 2044 580 2045
rect 638 2049 644 2050
rect 638 2045 639 2049
rect 643 2045 644 2049
rect 638 2044 644 2045
rect 710 2049 716 2050
rect 710 2045 711 2049
rect 715 2045 716 2049
rect 710 2044 716 2045
rect 790 2049 796 2050
rect 790 2045 791 2049
rect 795 2045 796 2049
rect 790 2044 796 2045
rect 862 2049 868 2050
rect 862 2045 863 2049
rect 867 2045 868 2049
rect 862 2044 868 2045
rect 942 2049 948 2050
rect 942 2045 943 2049
rect 947 2045 948 2049
rect 942 2044 948 2045
rect 1022 2049 1028 2050
rect 1022 2045 1023 2049
rect 1027 2045 1028 2049
rect 1022 2044 1028 2045
rect 1102 2049 1108 2050
rect 1102 2045 1103 2049
rect 1107 2045 1108 2049
rect 1102 2044 1108 2045
rect 1182 2049 1188 2050
rect 1182 2045 1183 2049
rect 1187 2045 1188 2049
rect 1182 2044 1188 2045
rect 1238 2049 1244 2050
rect 1238 2045 1239 2049
rect 1243 2045 1244 2049
rect 1238 2044 1244 2045
rect 1286 2048 1292 2049
rect 1286 2044 1287 2048
rect 1291 2044 1292 2048
rect 110 2043 116 2044
rect 1286 2043 1292 2044
rect 110 2031 116 2032
rect 110 2027 111 2031
rect 115 2027 116 2031
rect 1286 2031 1292 2032
rect 110 2026 116 2027
rect 382 2028 388 2029
rect 382 2024 383 2028
rect 387 2024 388 2028
rect 382 2023 388 2024
rect 438 2028 444 2029
rect 438 2024 439 2028
rect 443 2024 444 2028
rect 438 2023 444 2024
rect 494 2028 500 2029
rect 494 2024 495 2028
rect 499 2024 500 2028
rect 494 2023 500 2024
rect 558 2028 564 2029
rect 558 2024 559 2028
rect 563 2024 564 2028
rect 558 2023 564 2024
rect 622 2028 628 2029
rect 622 2024 623 2028
rect 627 2024 628 2028
rect 622 2023 628 2024
rect 694 2028 700 2029
rect 694 2024 695 2028
rect 699 2024 700 2028
rect 694 2023 700 2024
rect 774 2028 780 2029
rect 774 2024 775 2028
rect 779 2024 780 2028
rect 774 2023 780 2024
rect 846 2028 852 2029
rect 846 2024 847 2028
rect 851 2024 852 2028
rect 846 2023 852 2024
rect 926 2028 932 2029
rect 926 2024 927 2028
rect 931 2024 932 2028
rect 926 2023 932 2024
rect 1006 2028 1012 2029
rect 1006 2024 1007 2028
rect 1011 2024 1012 2028
rect 1006 2023 1012 2024
rect 1086 2028 1092 2029
rect 1086 2024 1087 2028
rect 1091 2024 1092 2028
rect 1086 2023 1092 2024
rect 1166 2028 1172 2029
rect 1166 2024 1167 2028
rect 1171 2024 1172 2028
rect 1166 2023 1172 2024
rect 1222 2028 1228 2029
rect 1222 2024 1223 2028
rect 1227 2024 1228 2028
rect 1286 2027 1287 2031
rect 1291 2027 1292 2031
rect 1446 2029 1452 2030
rect 1286 2026 1292 2027
rect 1326 2028 1332 2029
rect 1222 2023 1228 2024
rect 1326 2024 1327 2028
rect 1331 2024 1332 2028
rect 1446 2025 1447 2029
rect 1451 2025 1452 2029
rect 1446 2024 1452 2025
rect 1550 2029 1556 2030
rect 1550 2025 1551 2029
rect 1555 2025 1556 2029
rect 1550 2024 1556 2025
rect 1654 2029 1660 2030
rect 1654 2025 1655 2029
rect 1659 2025 1660 2029
rect 1654 2024 1660 2025
rect 1750 2029 1756 2030
rect 1750 2025 1751 2029
rect 1755 2025 1756 2029
rect 1750 2024 1756 2025
rect 1838 2029 1844 2030
rect 1838 2025 1839 2029
rect 1843 2025 1844 2029
rect 1838 2024 1844 2025
rect 1926 2029 1932 2030
rect 1926 2025 1927 2029
rect 1931 2025 1932 2029
rect 1926 2024 1932 2025
rect 2022 2029 2028 2030
rect 2022 2025 2023 2029
rect 2027 2025 2028 2029
rect 2022 2024 2028 2025
rect 2118 2029 2124 2030
rect 2118 2025 2119 2029
rect 2123 2025 2124 2029
rect 2118 2024 2124 2025
rect 2502 2028 2508 2029
rect 2502 2024 2503 2028
rect 2507 2024 2508 2028
rect 1326 2023 1332 2024
rect 2502 2023 2508 2024
rect 230 2012 236 2013
rect 110 2009 116 2010
rect 110 2005 111 2009
rect 115 2005 116 2009
rect 230 2008 231 2012
rect 235 2008 236 2012
rect 230 2007 236 2008
rect 286 2012 292 2013
rect 286 2008 287 2012
rect 291 2008 292 2012
rect 286 2007 292 2008
rect 358 2012 364 2013
rect 358 2008 359 2012
rect 363 2008 364 2012
rect 358 2007 364 2008
rect 438 2012 444 2013
rect 438 2008 439 2012
rect 443 2008 444 2012
rect 438 2007 444 2008
rect 534 2012 540 2013
rect 534 2008 535 2012
rect 539 2008 540 2012
rect 534 2007 540 2008
rect 630 2012 636 2013
rect 630 2008 631 2012
rect 635 2008 636 2012
rect 630 2007 636 2008
rect 734 2012 740 2013
rect 734 2008 735 2012
rect 739 2008 740 2012
rect 734 2007 740 2008
rect 846 2012 852 2013
rect 846 2008 847 2012
rect 851 2008 852 2012
rect 846 2007 852 2008
rect 958 2012 964 2013
rect 958 2008 959 2012
rect 963 2008 964 2012
rect 958 2007 964 2008
rect 1078 2012 1084 2013
rect 1078 2008 1079 2012
rect 1083 2008 1084 2012
rect 1078 2007 1084 2008
rect 1198 2012 1204 2013
rect 1198 2008 1199 2012
rect 1203 2008 1204 2012
rect 1326 2011 1332 2012
rect 1198 2007 1204 2008
rect 1286 2009 1292 2010
rect 110 2004 116 2005
rect 1286 2005 1287 2009
rect 1291 2005 1292 2009
rect 1326 2007 1327 2011
rect 1331 2007 1332 2011
rect 2502 2011 2508 2012
rect 1326 2006 1332 2007
rect 1430 2008 1436 2009
rect 1286 2004 1292 2005
rect 1430 2004 1431 2008
rect 1435 2004 1436 2008
rect 1430 2003 1436 2004
rect 1534 2008 1540 2009
rect 1534 2004 1535 2008
rect 1539 2004 1540 2008
rect 1534 2003 1540 2004
rect 1638 2008 1644 2009
rect 1638 2004 1639 2008
rect 1643 2004 1644 2008
rect 1638 2003 1644 2004
rect 1734 2008 1740 2009
rect 1734 2004 1735 2008
rect 1739 2004 1740 2008
rect 1734 2003 1740 2004
rect 1822 2008 1828 2009
rect 1822 2004 1823 2008
rect 1827 2004 1828 2008
rect 1822 2003 1828 2004
rect 1910 2008 1916 2009
rect 1910 2004 1911 2008
rect 1915 2004 1916 2008
rect 1910 2003 1916 2004
rect 2006 2008 2012 2009
rect 2006 2004 2007 2008
rect 2011 2004 2012 2008
rect 2006 2003 2012 2004
rect 2102 2008 2108 2009
rect 2102 2004 2103 2008
rect 2107 2004 2108 2008
rect 2502 2007 2503 2011
rect 2507 2007 2508 2011
rect 2502 2006 2508 2007
rect 2102 2003 2108 2004
rect 110 1992 116 1993
rect 1286 1992 1292 1993
rect 110 1988 111 1992
rect 115 1988 116 1992
rect 110 1987 116 1988
rect 246 1991 252 1992
rect 246 1987 247 1991
rect 251 1987 252 1991
rect 246 1986 252 1987
rect 302 1991 308 1992
rect 302 1987 303 1991
rect 307 1987 308 1991
rect 302 1986 308 1987
rect 374 1991 380 1992
rect 374 1987 375 1991
rect 379 1987 380 1991
rect 374 1986 380 1987
rect 454 1991 460 1992
rect 454 1987 455 1991
rect 459 1987 460 1991
rect 454 1986 460 1987
rect 550 1991 556 1992
rect 550 1987 551 1991
rect 555 1987 556 1991
rect 550 1986 556 1987
rect 646 1991 652 1992
rect 646 1987 647 1991
rect 651 1987 652 1991
rect 646 1986 652 1987
rect 750 1991 756 1992
rect 750 1987 751 1991
rect 755 1987 756 1991
rect 750 1986 756 1987
rect 862 1991 868 1992
rect 862 1987 863 1991
rect 867 1987 868 1991
rect 862 1986 868 1987
rect 974 1991 980 1992
rect 974 1987 975 1991
rect 979 1987 980 1991
rect 974 1986 980 1987
rect 1094 1991 1100 1992
rect 1094 1987 1095 1991
rect 1099 1987 1100 1991
rect 1094 1986 1100 1987
rect 1214 1991 1220 1992
rect 1214 1987 1215 1991
rect 1219 1987 1220 1991
rect 1286 1988 1287 1992
rect 1291 1988 1292 1992
rect 1454 1992 1460 1993
rect 1286 1987 1292 1988
rect 1326 1989 1332 1990
rect 1214 1986 1220 1987
rect 1326 1985 1327 1989
rect 1331 1985 1332 1989
rect 1454 1988 1455 1992
rect 1459 1988 1460 1992
rect 1454 1987 1460 1988
rect 1510 1992 1516 1993
rect 1510 1988 1511 1992
rect 1515 1988 1516 1992
rect 1510 1987 1516 1988
rect 1574 1992 1580 1993
rect 1574 1988 1575 1992
rect 1579 1988 1580 1992
rect 1574 1987 1580 1988
rect 1638 1992 1644 1993
rect 1638 1988 1639 1992
rect 1643 1988 1644 1992
rect 1638 1987 1644 1988
rect 1702 1992 1708 1993
rect 1702 1988 1703 1992
rect 1707 1988 1708 1992
rect 1702 1987 1708 1988
rect 1766 1992 1772 1993
rect 1766 1988 1767 1992
rect 1771 1988 1772 1992
rect 1766 1987 1772 1988
rect 1830 1992 1836 1993
rect 1830 1988 1831 1992
rect 1835 1988 1836 1992
rect 1830 1987 1836 1988
rect 1894 1992 1900 1993
rect 1894 1988 1895 1992
rect 1899 1988 1900 1992
rect 1894 1987 1900 1988
rect 1958 1992 1964 1993
rect 1958 1988 1959 1992
rect 1963 1988 1964 1992
rect 1958 1987 1964 1988
rect 2030 1992 2036 1993
rect 2030 1988 2031 1992
rect 2035 1988 2036 1992
rect 2030 1987 2036 1988
rect 2502 1989 2508 1990
rect 1326 1984 1332 1985
rect 2502 1985 2503 1989
rect 2507 1985 2508 1989
rect 2502 1984 2508 1985
rect 1326 1972 1332 1973
rect 2502 1972 2508 1973
rect 1326 1968 1327 1972
rect 1331 1968 1332 1972
rect 1326 1967 1332 1968
rect 1470 1971 1476 1972
rect 1470 1967 1471 1971
rect 1475 1967 1476 1971
rect 1470 1966 1476 1967
rect 1526 1971 1532 1972
rect 1526 1967 1527 1971
rect 1531 1967 1532 1971
rect 1526 1966 1532 1967
rect 1590 1971 1596 1972
rect 1590 1967 1591 1971
rect 1595 1967 1596 1971
rect 1590 1966 1596 1967
rect 1654 1971 1660 1972
rect 1654 1967 1655 1971
rect 1659 1967 1660 1971
rect 1654 1966 1660 1967
rect 1718 1971 1724 1972
rect 1718 1967 1719 1971
rect 1723 1967 1724 1971
rect 1718 1966 1724 1967
rect 1782 1971 1788 1972
rect 1782 1967 1783 1971
rect 1787 1967 1788 1971
rect 1782 1966 1788 1967
rect 1846 1971 1852 1972
rect 1846 1967 1847 1971
rect 1851 1967 1852 1971
rect 1846 1966 1852 1967
rect 1910 1971 1916 1972
rect 1910 1967 1911 1971
rect 1915 1967 1916 1971
rect 1910 1966 1916 1967
rect 1974 1971 1980 1972
rect 1974 1967 1975 1971
rect 1979 1967 1980 1971
rect 1974 1966 1980 1967
rect 2046 1971 2052 1972
rect 2046 1967 2047 1971
rect 2051 1967 2052 1971
rect 2502 1968 2503 1972
rect 2507 1968 2508 1972
rect 2502 1967 2508 1968
rect 2046 1966 2052 1967
rect 150 1937 156 1938
rect 110 1936 116 1937
rect 110 1932 111 1936
rect 115 1932 116 1936
rect 150 1933 151 1937
rect 155 1933 156 1937
rect 150 1932 156 1933
rect 214 1937 220 1938
rect 214 1933 215 1937
rect 219 1933 220 1937
rect 214 1932 220 1933
rect 318 1937 324 1938
rect 318 1933 319 1937
rect 323 1933 324 1937
rect 318 1932 324 1933
rect 438 1937 444 1938
rect 438 1933 439 1937
rect 443 1933 444 1937
rect 438 1932 444 1933
rect 582 1937 588 1938
rect 582 1933 583 1937
rect 587 1933 588 1937
rect 582 1932 588 1933
rect 742 1937 748 1938
rect 742 1933 743 1937
rect 747 1933 748 1937
rect 742 1932 748 1933
rect 918 1937 924 1938
rect 918 1933 919 1937
rect 923 1933 924 1937
rect 918 1932 924 1933
rect 1094 1937 1100 1938
rect 1094 1933 1095 1937
rect 1099 1933 1100 1937
rect 1094 1932 1100 1933
rect 1286 1936 1292 1937
rect 1286 1932 1287 1936
rect 1291 1932 1292 1936
rect 110 1931 116 1932
rect 1286 1931 1292 1932
rect 110 1919 116 1920
rect 110 1915 111 1919
rect 115 1915 116 1919
rect 1286 1919 1292 1920
rect 110 1914 116 1915
rect 134 1916 140 1917
rect 134 1912 135 1916
rect 139 1912 140 1916
rect 134 1911 140 1912
rect 198 1916 204 1917
rect 198 1912 199 1916
rect 203 1912 204 1916
rect 198 1911 204 1912
rect 302 1916 308 1917
rect 302 1912 303 1916
rect 307 1912 308 1916
rect 302 1911 308 1912
rect 422 1916 428 1917
rect 422 1912 423 1916
rect 427 1912 428 1916
rect 422 1911 428 1912
rect 566 1916 572 1917
rect 566 1912 567 1916
rect 571 1912 572 1916
rect 566 1911 572 1912
rect 726 1916 732 1917
rect 726 1912 727 1916
rect 731 1912 732 1916
rect 726 1911 732 1912
rect 902 1916 908 1917
rect 902 1912 903 1916
rect 907 1912 908 1916
rect 902 1911 908 1912
rect 1078 1916 1084 1917
rect 1078 1912 1079 1916
rect 1083 1912 1084 1916
rect 1286 1915 1287 1919
rect 1291 1915 1292 1919
rect 1566 1917 1572 1918
rect 1286 1914 1292 1915
rect 1326 1916 1332 1917
rect 1078 1911 1084 1912
rect 1326 1912 1327 1916
rect 1331 1912 1332 1916
rect 1566 1913 1567 1917
rect 1571 1913 1572 1917
rect 1566 1912 1572 1913
rect 1630 1917 1636 1918
rect 1630 1913 1631 1917
rect 1635 1913 1636 1917
rect 1630 1912 1636 1913
rect 1702 1917 1708 1918
rect 1702 1913 1703 1917
rect 1707 1913 1708 1917
rect 1702 1912 1708 1913
rect 1774 1917 1780 1918
rect 1774 1913 1775 1917
rect 1779 1913 1780 1917
rect 1774 1912 1780 1913
rect 1846 1917 1852 1918
rect 1846 1913 1847 1917
rect 1851 1913 1852 1917
rect 1846 1912 1852 1913
rect 1918 1917 1924 1918
rect 1918 1913 1919 1917
rect 1923 1913 1924 1917
rect 1918 1912 1924 1913
rect 1998 1917 2004 1918
rect 1998 1913 1999 1917
rect 2003 1913 2004 1917
rect 1998 1912 2004 1913
rect 2086 1917 2092 1918
rect 2086 1913 2087 1917
rect 2091 1913 2092 1917
rect 2086 1912 2092 1913
rect 2182 1917 2188 1918
rect 2182 1913 2183 1917
rect 2187 1913 2188 1917
rect 2182 1912 2188 1913
rect 2278 1917 2284 1918
rect 2278 1913 2279 1917
rect 2283 1913 2284 1917
rect 2278 1912 2284 1913
rect 2374 1917 2380 1918
rect 2374 1913 2375 1917
rect 2379 1913 2380 1917
rect 2374 1912 2380 1913
rect 2454 1917 2460 1918
rect 2454 1913 2455 1917
rect 2459 1913 2460 1917
rect 2454 1912 2460 1913
rect 2502 1916 2508 1917
rect 2502 1912 2503 1916
rect 2507 1912 2508 1916
rect 1326 1911 1332 1912
rect 2502 1911 2508 1912
rect 1326 1899 1332 1900
rect 134 1896 140 1897
rect 110 1893 116 1894
rect 110 1889 111 1893
rect 115 1889 116 1893
rect 134 1892 135 1896
rect 139 1892 140 1896
rect 134 1891 140 1892
rect 190 1896 196 1897
rect 190 1892 191 1896
rect 195 1892 196 1896
rect 190 1891 196 1892
rect 270 1896 276 1897
rect 270 1892 271 1896
rect 275 1892 276 1896
rect 270 1891 276 1892
rect 358 1896 364 1897
rect 358 1892 359 1896
rect 363 1892 364 1896
rect 358 1891 364 1892
rect 454 1896 460 1897
rect 454 1892 455 1896
rect 459 1892 460 1896
rect 454 1891 460 1892
rect 542 1896 548 1897
rect 542 1892 543 1896
rect 547 1892 548 1896
rect 542 1891 548 1892
rect 630 1896 636 1897
rect 630 1892 631 1896
rect 635 1892 636 1896
rect 630 1891 636 1892
rect 718 1896 724 1897
rect 718 1892 719 1896
rect 723 1892 724 1896
rect 718 1891 724 1892
rect 798 1896 804 1897
rect 798 1892 799 1896
rect 803 1892 804 1896
rect 798 1891 804 1892
rect 870 1896 876 1897
rect 870 1892 871 1896
rect 875 1892 876 1896
rect 870 1891 876 1892
rect 942 1896 948 1897
rect 942 1892 943 1896
rect 947 1892 948 1896
rect 942 1891 948 1892
rect 1014 1896 1020 1897
rect 1014 1892 1015 1896
rect 1019 1892 1020 1896
rect 1014 1891 1020 1892
rect 1086 1896 1092 1897
rect 1086 1892 1087 1896
rect 1091 1892 1092 1896
rect 1086 1891 1092 1892
rect 1158 1896 1164 1897
rect 1158 1892 1159 1896
rect 1163 1892 1164 1896
rect 1326 1895 1327 1899
rect 1331 1895 1332 1899
rect 2502 1899 2508 1900
rect 1326 1894 1332 1895
rect 1550 1896 1556 1897
rect 1158 1891 1164 1892
rect 1286 1893 1292 1894
rect 110 1888 116 1889
rect 1286 1889 1287 1893
rect 1291 1889 1292 1893
rect 1550 1892 1551 1896
rect 1555 1892 1556 1896
rect 1550 1891 1556 1892
rect 1614 1896 1620 1897
rect 1614 1892 1615 1896
rect 1619 1892 1620 1896
rect 1614 1891 1620 1892
rect 1686 1896 1692 1897
rect 1686 1892 1687 1896
rect 1691 1892 1692 1896
rect 1686 1891 1692 1892
rect 1758 1896 1764 1897
rect 1758 1892 1759 1896
rect 1763 1892 1764 1896
rect 1758 1891 1764 1892
rect 1830 1896 1836 1897
rect 1830 1892 1831 1896
rect 1835 1892 1836 1896
rect 1830 1891 1836 1892
rect 1902 1896 1908 1897
rect 1902 1892 1903 1896
rect 1907 1892 1908 1896
rect 1902 1891 1908 1892
rect 1982 1896 1988 1897
rect 1982 1892 1983 1896
rect 1987 1892 1988 1896
rect 1982 1891 1988 1892
rect 2070 1896 2076 1897
rect 2070 1892 2071 1896
rect 2075 1892 2076 1896
rect 2070 1891 2076 1892
rect 2166 1896 2172 1897
rect 2166 1892 2167 1896
rect 2171 1892 2172 1896
rect 2166 1891 2172 1892
rect 2262 1896 2268 1897
rect 2262 1892 2263 1896
rect 2267 1892 2268 1896
rect 2262 1891 2268 1892
rect 2358 1896 2364 1897
rect 2358 1892 2359 1896
rect 2363 1892 2364 1896
rect 2358 1891 2364 1892
rect 2438 1896 2444 1897
rect 2438 1892 2439 1896
rect 2443 1892 2444 1896
rect 2502 1895 2503 1899
rect 2507 1895 2508 1899
rect 2502 1894 2508 1895
rect 2438 1891 2444 1892
rect 1286 1888 1292 1889
rect 1606 1880 1612 1881
rect 1326 1877 1332 1878
rect 110 1876 116 1877
rect 1286 1876 1292 1877
rect 110 1872 111 1876
rect 115 1872 116 1876
rect 110 1871 116 1872
rect 150 1875 156 1876
rect 150 1871 151 1875
rect 155 1871 156 1875
rect 150 1870 156 1871
rect 206 1875 212 1876
rect 206 1871 207 1875
rect 211 1871 212 1875
rect 206 1870 212 1871
rect 286 1875 292 1876
rect 286 1871 287 1875
rect 291 1871 292 1875
rect 286 1870 292 1871
rect 374 1875 380 1876
rect 374 1871 375 1875
rect 379 1871 380 1875
rect 374 1870 380 1871
rect 470 1875 476 1876
rect 470 1871 471 1875
rect 475 1871 476 1875
rect 470 1870 476 1871
rect 558 1875 564 1876
rect 558 1871 559 1875
rect 563 1871 564 1875
rect 558 1870 564 1871
rect 646 1875 652 1876
rect 646 1871 647 1875
rect 651 1871 652 1875
rect 646 1870 652 1871
rect 734 1875 740 1876
rect 734 1871 735 1875
rect 739 1871 740 1875
rect 734 1870 740 1871
rect 814 1875 820 1876
rect 814 1871 815 1875
rect 819 1871 820 1875
rect 814 1870 820 1871
rect 886 1875 892 1876
rect 886 1871 887 1875
rect 891 1871 892 1875
rect 886 1870 892 1871
rect 958 1875 964 1876
rect 958 1871 959 1875
rect 963 1871 964 1875
rect 958 1870 964 1871
rect 1030 1875 1036 1876
rect 1030 1871 1031 1875
rect 1035 1871 1036 1875
rect 1030 1870 1036 1871
rect 1102 1875 1108 1876
rect 1102 1871 1103 1875
rect 1107 1871 1108 1875
rect 1102 1870 1108 1871
rect 1174 1875 1180 1876
rect 1174 1871 1175 1875
rect 1179 1871 1180 1875
rect 1286 1872 1287 1876
rect 1291 1872 1292 1876
rect 1326 1873 1327 1877
rect 1331 1873 1332 1877
rect 1606 1876 1607 1880
rect 1611 1876 1612 1880
rect 1606 1875 1612 1876
rect 1662 1880 1668 1881
rect 1662 1876 1663 1880
rect 1667 1876 1668 1880
rect 1662 1875 1668 1876
rect 1726 1880 1732 1881
rect 1726 1876 1727 1880
rect 1731 1876 1732 1880
rect 1726 1875 1732 1876
rect 1798 1880 1804 1881
rect 1798 1876 1799 1880
rect 1803 1876 1804 1880
rect 1798 1875 1804 1876
rect 1870 1880 1876 1881
rect 1870 1876 1871 1880
rect 1875 1876 1876 1880
rect 1870 1875 1876 1876
rect 1942 1880 1948 1881
rect 1942 1876 1943 1880
rect 1947 1876 1948 1880
rect 1942 1875 1948 1876
rect 2006 1880 2012 1881
rect 2006 1876 2007 1880
rect 2011 1876 2012 1880
rect 2006 1875 2012 1876
rect 2070 1880 2076 1881
rect 2070 1876 2071 1880
rect 2075 1876 2076 1880
rect 2070 1875 2076 1876
rect 2134 1880 2140 1881
rect 2134 1876 2135 1880
rect 2139 1876 2140 1880
rect 2134 1875 2140 1876
rect 2198 1880 2204 1881
rect 2198 1876 2199 1880
rect 2203 1876 2204 1880
rect 2198 1875 2204 1876
rect 2262 1880 2268 1881
rect 2262 1876 2263 1880
rect 2267 1876 2268 1880
rect 2262 1875 2268 1876
rect 2326 1880 2332 1881
rect 2326 1876 2327 1880
rect 2331 1876 2332 1880
rect 2326 1875 2332 1876
rect 2382 1880 2388 1881
rect 2382 1876 2383 1880
rect 2387 1876 2388 1880
rect 2382 1875 2388 1876
rect 2438 1880 2444 1881
rect 2438 1876 2439 1880
rect 2443 1876 2444 1880
rect 2438 1875 2444 1876
rect 2502 1877 2508 1878
rect 1326 1872 1332 1873
rect 2502 1873 2503 1877
rect 2507 1873 2508 1877
rect 2502 1872 2508 1873
rect 1286 1871 1292 1872
rect 1174 1870 1180 1871
rect 1326 1860 1332 1861
rect 2502 1860 2508 1861
rect 1326 1856 1327 1860
rect 1331 1856 1332 1860
rect 1326 1855 1332 1856
rect 1622 1859 1628 1860
rect 1622 1855 1623 1859
rect 1627 1855 1628 1859
rect 1622 1854 1628 1855
rect 1678 1859 1684 1860
rect 1678 1855 1679 1859
rect 1683 1855 1684 1859
rect 1678 1854 1684 1855
rect 1742 1859 1748 1860
rect 1742 1855 1743 1859
rect 1747 1855 1748 1859
rect 1742 1854 1748 1855
rect 1814 1859 1820 1860
rect 1814 1855 1815 1859
rect 1819 1855 1820 1859
rect 1814 1854 1820 1855
rect 1886 1859 1892 1860
rect 1886 1855 1887 1859
rect 1891 1855 1892 1859
rect 1886 1854 1892 1855
rect 1958 1859 1964 1860
rect 1958 1855 1959 1859
rect 1963 1855 1964 1859
rect 1958 1854 1964 1855
rect 2022 1859 2028 1860
rect 2022 1855 2023 1859
rect 2027 1855 2028 1859
rect 2022 1854 2028 1855
rect 2086 1859 2092 1860
rect 2086 1855 2087 1859
rect 2091 1855 2092 1859
rect 2086 1854 2092 1855
rect 2150 1859 2156 1860
rect 2150 1855 2151 1859
rect 2155 1855 2156 1859
rect 2150 1854 2156 1855
rect 2214 1859 2220 1860
rect 2214 1855 2215 1859
rect 2219 1855 2220 1859
rect 2214 1854 2220 1855
rect 2278 1859 2284 1860
rect 2278 1855 2279 1859
rect 2283 1855 2284 1859
rect 2278 1854 2284 1855
rect 2342 1859 2348 1860
rect 2342 1855 2343 1859
rect 2347 1855 2348 1859
rect 2342 1854 2348 1855
rect 2398 1859 2404 1860
rect 2398 1855 2399 1859
rect 2403 1855 2404 1859
rect 2398 1854 2404 1855
rect 2454 1859 2460 1860
rect 2454 1855 2455 1859
rect 2459 1855 2460 1859
rect 2502 1856 2503 1860
rect 2507 1856 2508 1860
rect 2502 1855 2508 1856
rect 2454 1854 2460 1855
rect 150 1825 156 1826
rect 110 1824 116 1825
rect 110 1820 111 1824
rect 115 1820 116 1824
rect 150 1821 151 1825
rect 155 1821 156 1825
rect 150 1820 156 1821
rect 206 1825 212 1826
rect 206 1821 207 1825
rect 211 1821 212 1825
rect 206 1820 212 1821
rect 294 1825 300 1826
rect 294 1821 295 1825
rect 299 1821 300 1825
rect 294 1820 300 1821
rect 390 1825 396 1826
rect 390 1821 391 1825
rect 395 1821 396 1825
rect 390 1820 396 1821
rect 494 1825 500 1826
rect 494 1821 495 1825
rect 499 1821 500 1825
rect 494 1820 500 1821
rect 590 1825 596 1826
rect 590 1821 591 1825
rect 595 1821 596 1825
rect 590 1820 596 1821
rect 686 1825 692 1826
rect 686 1821 687 1825
rect 691 1821 692 1825
rect 686 1820 692 1821
rect 774 1825 780 1826
rect 774 1821 775 1825
rect 779 1821 780 1825
rect 774 1820 780 1821
rect 854 1825 860 1826
rect 854 1821 855 1825
rect 859 1821 860 1825
rect 854 1820 860 1821
rect 926 1825 932 1826
rect 926 1821 927 1825
rect 931 1821 932 1825
rect 926 1820 932 1821
rect 998 1825 1004 1826
rect 998 1821 999 1825
rect 1003 1821 1004 1825
rect 998 1820 1004 1821
rect 1078 1825 1084 1826
rect 1078 1821 1079 1825
rect 1083 1821 1084 1825
rect 1078 1820 1084 1821
rect 1158 1825 1164 1826
rect 1158 1821 1159 1825
rect 1163 1821 1164 1825
rect 1158 1820 1164 1821
rect 1286 1824 1292 1825
rect 1286 1820 1287 1824
rect 1291 1820 1292 1824
rect 110 1819 116 1820
rect 1286 1819 1292 1820
rect 110 1807 116 1808
rect 110 1803 111 1807
rect 115 1803 116 1807
rect 1286 1807 1292 1808
rect 110 1802 116 1803
rect 134 1804 140 1805
rect 134 1800 135 1804
rect 139 1800 140 1804
rect 134 1799 140 1800
rect 190 1804 196 1805
rect 190 1800 191 1804
rect 195 1800 196 1804
rect 190 1799 196 1800
rect 278 1804 284 1805
rect 278 1800 279 1804
rect 283 1800 284 1804
rect 278 1799 284 1800
rect 374 1804 380 1805
rect 374 1800 375 1804
rect 379 1800 380 1804
rect 374 1799 380 1800
rect 478 1804 484 1805
rect 478 1800 479 1804
rect 483 1800 484 1804
rect 478 1799 484 1800
rect 574 1804 580 1805
rect 574 1800 575 1804
rect 579 1800 580 1804
rect 574 1799 580 1800
rect 670 1804 676 1805
rect 670 1800 671 1804
rect 675 1800 676 1804
rect 670 1799 676 1800
rect 758 1804 764 1805
rect 758 1800 759 1804
rect 763 1800 764 1804
rect 758 1799 764 1800
rect 838 1804 844 1805
rect 838 1800 839 1804
rect 843 1800 844 1804
rect 838 1799 844 1800
rect 910 1804 916 1805
rect 910 1800 911 1804
rect 915 1800 916 1804
rect 910 1799 916 1800
rect 982 1804 988 1805
rect 982 1800 983 1804
rect 987 1800 988 1804
rect 982 1799 988 1800
rect 1062 1804 1068 1805
rect 1062 1800 1063 1804
rect 1067 1800 1068 1804
rect 1062 1799 1068 1800
rect 1142 1804 1148 1805
rect 1142 1800 1143 1804
rect 1147 1800 1148 1804
rect 1286 1803 1287 1807
rect 1291 1803 1292 1807
rect 1630 1805 1636 1806
rect 1286 1802 1292 1803
rect 1326 1804 1332 1805
rect 1142 1799 1148 1800
rect 1326 1800 1327 1804
rect 1331 1800 1332 1804
rect 1630 1801 1631 1805
rect 1635 1801 1636 1805
rect 1630 1800 1636 1801
rect 1718 1805 1724 1806
rect 1718 1801 1719 1805
rect 1723 1801 1724 1805
rect 1718 1800 1724 1801
rect 1814 1805 1820 1806
rect 1814 1801 1815 1805
rect 1819 1801 1820 1805
rect 1814 1800 1820 1801
rect 1926 1805 1932 1806
rect 1926 1801 1927 1805
rect 1931 1801 1932 1805
rect 1926 1800 1932 1801
rect 2054 1805 2060 1806
rect 2054 1801 2055 1805
rect 2059 1801 2060 1805
rect 2054 1800 2060 1801
rect 2190 1805 2196 1806
rect 2190 1801 2191 1805
rect 2195 1801 2196 1805
rect 2190 1800 2196 1801
rect 2334 1805 2340 1806
rect 2334 1801 2335 1805
rect 2339 1801 2340 1805
rect 2334 1800 2340 1801
rect 2454 1805 2460 1806
rect 2454 1801 2455 1805
rect 2459 1801 2460 1805
rect 2454 1800 2460 1801
rect 2502 1804 2508 1805
rect 2502 1800 2503 1804
rect 2507 1800 2508 1804
rect 1326 1799 1332 1800
rect 2502 1799 2508 1800
rect 1326 1787 1332 1788
rect 1326 1783 1327 1787
rect 1331 1783 1332 1787
rect 2502 1787 2508 1788
rect 1326 1782 1332 1783
rect 1614 1784 1620 1785
rect 134 1780 140 1781
rect 110 1777 116 1778
rect 110 1773 111 1777
rect 115 1773 116 1777
rect 134 1776 135 1780
rect 139 1776 140 1780
rect 134 1775 140 1776
rect 198 1780 204 1781
rect 198 1776 199 1780
rect 203 1776 204 1780
rect 198 1775 204 1776
rect 294 1780 300 1781
rect 294 1776 295 1780
rect 299 1776 300 1780
rect 294 1775 300 1776
rect 398 1780 404 1781
rect 398 1776 399 1780
rect 403 1776 404 1780
rect 398 1775 404 1776
rect 502 1780 508 1781
rect 502 1776 503 1780
rect 507 1776 508 1780
rect 502 1775 508 1776
rect 606 1780 612 1781
rect 606 1776 607 1780
rect 611 1776 612 1780
rect 606 1775 612 1776
rect 702 1780 708 1781
rect 702 1776 703 1780
rect 707 1776 708 1780
rect 702 1775 708 1776
rect 798 1780 804 1781
rect 798 1776 799 1780
rect 803 1776 804 1780
rect 798 1775 804 1776
rect 886 1780 892 1781
rect 886 1776 887 1780
rect 891 1776 892 1780
rect 886 1775 892 1776
rect 974 1780 980 1781
rect 974 1776 975 1780
rect 979 1776 980 1780
rect 974 1775 980 1776
rect 1062 1780 1068 1781
rect 1062 1776 1063 1780
rect 1067 1776 1068 1780
rect 1062 1775 1068 1776
rect 1150 1780 1156 1781
rect 1150 1776 1151 1780
rect 1155 1776 1156 1780
rect 1614 1780 1615 1784
rect 1619 1780 1620 1784
rect 1614 1779 1620 1780
rect 1702 1784 1708 1785
rect 1702 1780 1703 1784
rect 1707 1780 1708 1784
rect 1702 1779 1708 1780
rect 1798 1784 1804 1785
rect 1798 1780 1799 1784
rect 1803 1780 1804 1784
rect 1798 1779 1804 1780
rect 1910 1784 1916 1785
rect 1910 1780 1911 1784
rect 1915 1780 1916 1784
rect 1910 1779 1916 1780
rect 2038 1784 2044 1785
rect 2038 1780 2039 1784
rect 2043 1780 2044 1784
rect 2038 1779 2044 1780
rect 2174 1784 2180 1785
rect 2174 1780 2175 1784
rect 2179 1780 2180 1784
rect 2174 1779 2180 1780
rect 2318 1784 2324 1785
rect 2318 1780 2319 1784
rect 2323 1780 2324 1784
rect 2318 1779 2324 1780
rect 2438 1784 2444 1785
rect 2438 1780 2439 1784
rect 2443 1780 2444 1784
rect 2502 1783 2503 1787
rect 2507 1783 2508 1787
rect 2502 1782 2508 1783
rect 2438 1779 2444 1780
rect 1150 1775 1156 1776
rect 1286 1777 1292 1778
rect 110 1772 116 1773
rect 1286 1773 1287 1777
rect 1291 1773 1292 1777
rect 1286 1772 1292 1773
rect 1526 1772 1532 1773
rect 1326 1769 1332 1770
rect 1326 1765 1327 1769
rect 1331 1765 1332 1769
rect 1526 1768 1527 1772
rect 1531 1768 1532 1772
rect 1526 1767 1532 1768
rect 1606 1772 1612 1773
rect 1606 1768 1607 1772
rect 1611 1768 1612 1772
rect 1606 1767 1612 1768
rect 1694 1772 1700 1773
rect 1694 1768 1695 1772
rect 1699 1768 1700 1772
rect 1694 1767 1700 1768
rect 1790 1772 1796 1773
rect 1790 1768 1791 1772
rect 1795 1768 1796 1772
rect 1790 1767 1796 1768
rect 1878 1772 1884 1773
rect 1878 1768 1879 1772
rect 1883 1768 1884 1772
rect 1878 1767 1884 1768
rect 1966 1772 1972 1773
rect 1966 1768 1967 1772
rect 1971 1768 1972 1772
rect 1966 1767 1972 1768
rect 2054 1772 2060 1773
rect 2054 1768 2055 1772
rect 2059 1768 2060 1772
rect 2054 1767 2060 1768
rect 2134 1772 2140 1773
rect 2134 1768 2135 1772
rect 2139 1768 2140 1772
rect 2134 1767 2140 1768
rect 2214 1772 2220 1773
rect 2214 1768 2215 1772
rect 2219 1768 2220 1772
rect 2214 1767 2220 1768
rect 2294 1772 2300 1773
rect 2294 1768 2295 1772
rect 2299 1768 2300 1772
rect 2294 1767 2300 1768
rect 2374 1772 2380 1773
rect 2374 1768 2375 1772
rect 2379 1768 2380 1772
rect 2374 1767 2380 1768
rect 2438 1772 2444 1773
rect 2438 1768 2439 1772
rect 2443 1768 2444 1772
rect 2438 1767 2444 1768
rect 2502 1769 2508 1770
rect 1326 1764 1332 1765
rect 2502 1765 2503 1769
rect 2507 1765 2508 1769
rect 2502 1764 2508 1765
rect 110 1760 116 1761
rect 1286 1760 1292 1761
rect 110 1756 111 1760
rect 115 1756 116 1760
rect 110 1755 116 1756
rect 150 1759 156 1760
rect 150 1755 151 1759
rect 155 1755 156 1759
rect 150 1754 156 1755
rect 214 1759 220 1760
rect 214 1755 215 1759
rect 219 1755 220 1759
rect 214 1754 220 1755
rect 310 1759 316 1760
rect 310 1755 311 1759
rect 315 1755 316 1759
rect 310 1754 316 1755
rect 414 1759 420 1760
rect 414 1755 415 1759
rect 419 1755 420 1759
rect 414 1754 420 1755
rect 518 1759 524 1760
rect 518 1755 519 1759
rect 523 1755 524 1759
rect 518 1754 524 1755
rect 622 1759 628 1760
rect 622 1755 623 1759
rect 627 1755 628 1759
rect 622 1754 628 1755
rect 718 1759 724 1760
rect 718 1755 719 1759
rect 723 1755 724 1759
rect 718 1754 724 1755
rect 814 1759 820 1760
rect 814 1755 815 1759
rect 819 1755 820 1759
rect 814 1754 820 1755
rect 902 1759 908 1760
rect 902 1755 903 1759
rect 907 1755 908 1759
rect 902 1754 908 1755
rect 990 1759 996 1760
rect 990 1755 991 1759
rect 995 1755 996 1759
rect 990 1754 996 1755
rect 1078 1759 1084 1760
rect 1078 1755 1079 1759
rect 1083 1755 1084 1759
rect 1078 1754 1084 1755
rect 1166 1759 1172 1760
rect 1166 1755 1167 1759
rect 1171 1755 1172 1759
rect 1286 1756 1287 1760
rect 1291 1756 1292 1760
rect 1286 1755 1292 1756
rect 1166 1754 1172 1755
rect 1326 1752 1332 1753
rect 2502 1752 2508 1753
rect 1326 1748 1327 1752
rect 1331 1748 1332 1752
rect 1326 1747 1332 1748
rect 1542 1751 1548 1752
rect 1542 1747 1543 1751
rect 1547 1747 1548 1751
rect 1542 1746 1548 1747
rect 1622 1751 1628 1752
rect 1622 1747 1623 1751
rect 1627 1747 1628 1751
rect 1622 1746 1628 1747
rect 1710 1751 1716 1752
rect 1710 1747 1711 1751
rect 1715 1747 1716 1751
rect 1710 1746 1716 1747
rect 1806 1751 1812 1752
rect 1806 1747 1807 1751
rect 1811 1747 1812 1751
rect 1806 1746 1812 1747
rect 1894 1751 1900 1752
rect 1894 1747 1895 1751
rect 1899 1747 1900 1751
rect 1894 1746 1900 1747
rect 1982 1751 1988 1752
rect 1982 1747 1983 1751
rect 1987 1747 1988 1751
rect 1982 1746 1988 1747
rect 2070 1751 2076 1752
rect 2070 1747 2071 1751
rect 2075 1747 2076 1751
rect 2070 1746 2076 1747
rect 2150 1751 2156 1752
rect 2150 1747 2151 1751
rect 2155 1747 2156 1751
rect 2150 1746 2156 1747
rect 2230 1751 2236 1752
rect 2230 1747 2231 1751
rect 2235 1747 2236 1751
rect 2230 1746 2236 1747
rect 2310 1751 2316 1752
rect 2310 1747 2311 1751
rect 2315 1747 2316 1751
rect 2310 1746 2316 1747
rect 2390 1751 2396 1752
rect 2390 1747 2391 1751
rect 2395 1747 2396 1751
rect 2390 1746 2396 1747
rect 2454 1751 2460 1752
rect 2454 1747 2455 1751
rect 2459 1747 2460 1751
rect 2502 1748 2503 1752
rect 2507 1748 2508 1752
rect 2502 1747 2508 1748
rect 2454 1746 2460 1747
rect 166 1705 172 1706
rect 110 1704 116 1705
rect 110 1700 111 1704
rect 115 1700 116 1704
rect 166 1701 167 1705
rect 171 1701 172 1705
rect 166 1700 172 1701
rect 238 1705 244 1706
rect 238 1701 239 1705
rect 243 1701 244 1705
rect 238 1700 244 1701
rect 318 1705 324 1706
rect 318 1701 319 1705
rect 323 1701 324 1705
rect 318 1700 324 1701
rect 406 1705 412 1706
rect 406 1701 407 1705
rect 411 1701 412 1705
rect 406 1700 412 1701
rect 502 1705 508 1706
rect 502 1701 503 1705
rect 507 1701 508 1705
rect 502 1700 508 1701
rect 606 1705 612 1706
rect 606 1701 607 1705
rect 611 1701 612 1705
rect 606 1700 612 1701
rect 710 1705 716 1706
rect 710 1701 711 1705
rect 715 1701 716 1705
rect 710 1700 716 1701
rect 822 1705 828 1706
rect 822 1701 823 1705
rect 827 1701 828 1705
rect 822 1700 828 1701
rect 934 1705 940 1706
rect 934 1701 935 1705
rect 939 1701 940 1705
rect 934 1700 940 1701
rect 1046 1705 1052 1706
rect 1046 1701 1047 1705
rect 1051 1701 1052 1705
rect 1046 1700 1052 1701
rect 1158 1705 1164 1706
rect 1158 1701 1159 1705
rect 1163 1701 1164 1705
rect 1158 1700 1164 1701
rect 1286 1704 1292 1705
rect 1286 1700 1287 1704
rect 1291 1700 1292 1704
rect 110 1699 116 1700
rect 1286 1699 1292 1700
rect 1398 1697 1404 1698
rect 1326 1696 1332 1697
rect 1326 1692 1327 1696
rect 1331 1692 1332 1696
rect 1398 1693 1399 1697
rect 1403 1693 1404 1697
rect 1398 1692 1404 1693
rect 1462 1697 1468 1698
rect 1462 1693 1463 1697
rect 1467 1693 1468 1697
rect 1462 1692 1468 1693
rect 1542 1697 1548 1698
rect 1542 1693 1543 1697
rect 1547 1693 1548 1697
rect 1542 1692 1548 1693
rect 1630 1697 1636 1698
rect 1630 1693 1631 1697
rect 1635 1693 1636 1697
rect 1630 1692 1636 1693
rect 1726 1697 1732 1698
rect 1726 1693 1727 1697
rect 1731 1693 1732 1697
rect 1726 1692 1732 1693
rect 1822 1697 1828 1698
rect 1822 1693 1823 1697
rect 1827 1693 1828 1697
rect 1822 1692 1828 1693
rect 1918 1697 1924 1698
rect 1918 1693 1919 1697
rect 1923 1693 1924 1697
rect 1918 1692 1924 1693
rect 2014 1697 2020 1698
rect 2014 1693 2015 1697
rect 2019 1693 2020 1697
rect 2014 1692 2020 1693
rect 2110 1697 2116 1698
rect 2110 1693 2111 1697
rect 2115 1693 2116 1697
rect 2110 1692 2116 1693
rect 2198 1697 2204 1698
rect 2198 1693 2199 1697
rect 2203 1693 2204 1697
rect 2198 1692 2204 1693
rect 2286 1697 2292 1698
rect 2286 1693 2287 1697
rect 2291 1693 2292 1697
rect 2286 1692 2292 1693
rect 2382 1697 2388 1698
rect 2382 1693 2383 1697
rect 2387 1693 2388 1697
rect 2382 1692 2388 1693
rect 2454 1697 2460 1698
rect 2454 1693 2455 1697
rect 2459 1693 2460 1697
rect 2454 1692 2460 1693
rect 2502 1696 2508 1697
rect 2502 1692 2503 1696
rect 2507 1692 2508 1696
rect 1326 1691 1332 1692
rect 2502 1691 2508 1692
rect 110 1687 116 1688
rect 110 1683 111 1687
rect 115 1683 116 1687
rect 1286 1687 1292 1688
rect 110 1682 116 1683
rect 150 1684 156 1685
rect 150 1680 151 1684
rect 155 1680 156 1684
rect 150 1679 156 1680
rect 222 1684 228 1685
rect 222 1680 223 1684
rect 227 1680 228 1684
rect 222 1679 228 1680
rect 302 1684 308 1685
rect 302 1680 303 1684
rect 307 1680 308 1684
rect 302 1679 308 1680
rect 390 1684 396 1685
rect 390 1680 391 1684
rect 395 1680 396 1684
rect 390 1679 396 1680
rect 486 1684 492 1685
rect 486 1680 487 1684
rect 491 1680 492 1684
rect 486 1679 492 1680
rect 590 1684 596 1685
rect 590 1680 591 1684
rect 595 1680 596 1684
rect 590 1679 596 1680
rect 694 1684 700 1685
rect 694 1680 695 1684
rect 699 1680 700 1684
rect 694 1679 700 1680
rect 806 1684 812 1685
rect 806 1680 807 1684
rect 811 1680 812 1684
rect 806 1679 812 1680
rect 918 1684 924 1685
rect 918 1680 919 1684
rect 923 1680 924 1684
rect 918 1679 924 1680
rect 1030 1684 1036 1685
rect 1030 1680 1031 1684
rect 1035 1680 1036 1684
rect 1030 1679 1036 1680
rect 1142 1684 1148 1685
rect 1142 1680 1143 1684
rect 1147 1680 1148 1684
rect 1286 1683 1287 1687
rect 1291 1683 1292 1687
rect 1286 1682 1292 1683
rect 1142 1679 1148 1680
rect 1326 1679 1332 1680
rect 1326 1675 1327 1679
rect 1331 1675 1332 1679
rect 2502 1679 2508 1680
rect 1326 1674 1332 1675
rect 1382 1676 1388 1677
rect 1382 1672 1383 1676
rect 1387 1672 1388 1676
rect 1382 1671 1388 1672
rect 1446 1676 1452 1677
rect 1446 1672 1447 1676
rect 1451 1672 1452 1676
rect 1446 1671 1452 1672
rect 1526 1676 1532 1677
rect 1526 1672 1527 1676
rect 1531 1672 1532 1676
rect 1526 1671 1532 1672
rect 1614 1676 1620 1677
rect 1614 1672 1615 1676
rect 1619 1672 1620 1676
rect 1614 1671 1620 1672
rect 1710 1676 1716 1677
rect 1710 1672 1711 1676
rect 1715 1672 1716 1676
rect 1710 1671 1716 1672
rect 1806 1676 1812 1677
rect 1806 1672 1807 1676
rect 1811 1672 1812 1676
rect 1806 1671 1812 1672
rect 1902 1676 1908 1677
rect 1902 1672 1903 1676
rect 1907 1672 1908 1676
rect 1902 1671 1908 1672
rect 1998 1676 2004 1677
rect 1998 1672 1999 1676
rect 2003 1672 2004 1676
rect 1998 1671 2004 1672
rect 2094 1676 2100 1677
rect 2094 1672 2095 1676
rect 2099 1672 2100 1676
rect 2094 1671 2100 1672
rect 2182 1676 2188 1677
rect 2182 1672 2183 1676
rect 2187 1672 2188 1676
rect 2182 1671 2188 1672
rect 2270 1676 2276 1677
rect 2270 1672 2271 1676
rect 2275 1672 2276 1676
rect 2270 1671 2276 1672
rect 2366 1676 2372 1677
rect 2366 1672 2367 1676
rect 2371 1672 2372 1676
rect 2366 1671 2372 1672
rect 2438 1676 2444 1677
rect 2438 1672 2439 1676
rect 2443 1672 2444 1676
rect 2502 1675 2503 1679
rect 2507 1675 2508 1679
rect 2502 1674 2508 1675
rect 2438 1671 2444 1672
rect 254 1668 260 1669
rect 110 1665 116 1666
rect 110 1661 111 1665
rect 115 1661 116 1665
rect 254 1664 255 1668
rect 259 1664 260 1668
rect 254 1663 260 1664
rect 318 1668 324 1669
rect 318 1664 319 1668
rect 323 1664 324 1668
rect 318 1663 324 1664
rect 398 1668 404 1669
rect 398 1664 399 1668
rect 403 1664 404 1668
rect 398 1663 404 1664
rect 486 1668 492 1669
rect 486 1664 487 1668
rect 491 1664 492 1668
rect 486 1663 492 1664
rect 574 1668 580 1669
rect 574 1664 575 1668
rect 579 1664 580 1668
rect 574 1663 580 1664
rect 670 1668 676 1669
rect 670 1664 671 1668
rect 675 1664 676 1668
rect 670 1663 676 1664
rect 766 1668 772 1669
rect 766 1664 767 1668
rect 771 1664 772 1668
rect 766 1663 772 1664
rect 862 1668 868 1669
rect 862 1664 863 1668
rect 867 1664 868 1668
rect 862 1663 868 1664
rect 958 1668 964 1669
rect 958 1664 959 1668
rect 963 1664 964 1668
rect 958 1663 964 1664
rect 1062 1668 1068 1669
rect 1062 1664 1063 1668
rect 1067 1664 1068 1668
rect 1062 1663 1068 1664
rect 1166 1668 1172 1669
rect 1166 1664 1167 1668
rect 1171 1664 1172 1668
rect 1166 1663 1172 1664
rect 1286 1665 1292 1666
rect 110 1660 116 1661
rect 1286 1661 1287 1665
rect 1291 1661 1292 1665
rect 1286 1660 1292 1661
rect 1350 1660 1356 1661
rect 1326 1657 1332 1658
rect 1326 1653 1327 1657
rect 1331 1653 1332 1657
rect 1350 1656 1351 1660
rect 1355 1656 1356 1660
rect 1350 1655 1356 1656
rect 1406 1660 1412 1661
rect 1406 1656 1407 1660
rect 1411 1656 1412 1660
rect 1406 1655 1412 1656
rect 1494 1660 1500 1661
rect 1494 1656 1495 1660
rect 1499 1656 1500 1660
rect 1494 1655 1500 1656
rect 1582 1660 1588 1661
rect 1582 1656 1583 1660
rect 1587 1656 1588 1660
rect 1582 1655 1588 1656
rect 1678 1660 1684 1661
rect 1678 1656 1679 1660
rect 1683 1656 1684 1660
rect 1678 1655 1684 1656
rect 1782 1660 1788 1661
rect 1782 1656 1783 1660
rect 1787 1656 1788 1660
rect 1782 1655 1788 1656
rect 1894 1660 1900 1661
rect 1894 1656 1895 1660
rect 1899 1656 1900 1660
rect 1894 1655 1900 1656
rect 2022 1660 2028 1661
rect 2022 1656 2023 1660
rect 2027 1656 2028 1660
rect 2022 1655 2028 1656
rect 2158 1660 2164 1661
rect 2158 1656 2159 1660
rect 2163 1656 2164 1660
rect 2158 1655 2164 1656
rect 2302 1660 2308 1661
rect 2302 1656 2303 1660
rect 2307 1656 2308 1660
rect 2302 1655 2308 1656
rect 2438 1660 2444 1661
rect 2438 1656 2439 1660
rect 2443 1656 2444 1660
rect 2438 1655 2444 1656
rect 2502 1657 2508 1658
rect 1326 1652 1332 1653
rect 2502 1653 2503 1657
rect 2507 1653 2508 1657
rect 2502 1652 2508 1653
rect 110 1648 116 1649
rect 1286 1648 1292 1649
rect 110 1644 111 1648
rect 115 1644 116 1648
rect 110 1643 116 1644
rect 270 1647 276 1648
rect 270 1643 271 1647
rect 275 1643 276 1647
rect 270 1642 276 1643
rect 334 1647 340 1648
rect 334 1643 335 1647
rect 339 1643 340 1647
rect 334 1642 340 1643
rect 414 1647 420 1648
rect 414 1643 415 1647
rect 419 1643 420 1647
rect 414 1642 420 1643
rect 502 1647 508 1648
rect 502 1643 503 1647
rect 507 1643 508 1647
rect 502 1642 508 1643
rect 590 1647 596 1648
rect 590 1643 591 1647
rect 595 1643 596 1647
rect 590 1642 596 1643
rect 686 1647 692 1648
rect 686 1643 687 1647
rect 691 1643 692 1647
rect 686 1642 692 1643
rect 782 1647 788 1648
rect 782 1643 783 1647
rect 787 1643 788 1647
rect 782 1642 788 1643
rect 878 1647 884 1648
rect 878 1643 879 1647
rect 883 1643 884 1647
rect 878 1642 884 1643
rect 974 1647 980 1648
rect 974 1643 975 1647
rect 979 1643 980 1647
rect 974 1642 980 1643
rect 1078 1647 1084 1648
rect 1078 1643 1079 1647
rect 1083 1643 1084 1647
rect 1078 1642 1084 1643
rect 1182 1647 1188 1648
rect 1182 1643 1183 1647
rect 1187 1643 1188 1647
rect 1286 1644 1287 1648
rect 1291 1644 1292 1648
rect 1286 1643 1292 1644
rect 1182 1642 1188 1643
rect 1326 1640 1332 1641
rect 2502 1640 2508 1641
rect 1326 1636 1327 1640
rect 1331 1636 1332 1640
rect 1326 1635 1332 1636
rect 1366 1639 1372 1640
rect 1366 1635 1367 1639
rect 1371 1635 1372 1639
rect 1366 1634 1372 1635
rect 1422 1639 1428 1640
rect 1422 1635 1423 1639
rect 1427 1635 1428 1639
rect 1422 1634 1428 1635
rect 1510 1639 1516 1640
rect 1510 1635 1511 1639
rect 1515 1635 1516 1639
rect 1510 1634 1516 1635
rect 1598 1639 1604 1640
rect 1598 1635 1599 1639
rect 1603 1635 1604 1639
rect 1598 1634 1604 1635
rect 1694 1639 1700 1640
rect 1694 1635 1695 1639
rect 1699 1635 1700 1639
rect 1694 1634 1700 1635
rect 1798 1639 1804 1640
rect 1798 1635 1799 1639
rect 1803 1635 1804 1639
rect 1798 1634 1804 1635
rect 1910 1639 1916 1640
rect 1910 1635 1911 1639
rect 1915 1635 1916 1639
rect 1910 1634 1916 1635
rect 2038 1639 2044 1640
rect 2038 1635 2039 1639
rect 2043 1635 2044 1639
rect 2038 1634 2044 1635
rect 2174 1639 2180 1640
rect 2174 1635 2175 1639
rect 2179 1635 2180 1639
rect 2174 1634 2180 1635
rect 2318 1639 2324 1640
rect 2318 1635 2319 1639
rect 2323 1635 2324 1639
rect 2318 1634 2324 1635
rect 2454 1639 2460 1640
rect 2454 1635 2455 1639
rect 2459 1635 2460 1639
rect 2502 1636 2503 1640
rect 2507 1636 2508 1640
rect 2502 1635 2508 1636
rect 2454 1634 2460 1635
rect 302 1593 308 1594
rect 110 1592 116 1593
rect 110 1588 111 1592
rect 115 1588 116 1592
rect 302 1589 303 1593
rect 307 1589 308 1593
rect 302 1588 308 1589
rect 358 1593 364 1594
rect 358 1589 359 1593
rect 363 1589 364 1593
rect 358 1588 364 1589
rect 430 1593 436 1594
rect 430 1589 431 1593
rect 435 1589 436 1593
rect 430 1588 436 1589
rect 510 1593 516 1594
rect 510 1589 511 1593
rect 515 1589 516 1593
rect 510 1588 516 1589
rect 598 1593 604 1594
rect 598 1589 599 1593
rect 603 1589 604 1593
rect 598 1588 604 1589
rect 694 1593 700 1594
rect 694 1589 695 1593
rect 699 1589 700 1593
rect 694 1588 700 1589
rect 790 1593 796 1594
rect 790 1589 791 1593
rect 795 1589 796 1593
rect 790 1588 796 1589
rect 894 1593 900 1594
rect 894 1589 895 1593
rect 899 1589 900 1593
rect 894 1588 900 1589
rect 1006 1593 1012 1594
rect 1006 1589 1007 1593
rect 1011 1589 1012 1593
rect 1006 1588 1012 1589
rect 1118 1593 1124 1594
rect 1118 1589 1119 1593
rect 1123 1589 1124 1593
rect 1118 1588 1124 1589
rect 1286 1592 1292 1593
rect 1286 1588 1287 1592
rect 1291 1588 1292 1592
rect 1366 1589 1372 1590
rect 110 1587 116 1588
rect 1286 1587 1292 1588
rect 1326 1588 1332 1589
rect 1326 1584 1327 1588
rect 1331 1584 1332 1588
rect 1366 1585 1367 1589
rect 1371 1585 1372 1589
rect 1366 1584 1372 1585
rect 1422 1589 1428 1590
rect 1422 1585 1423 1589
rect 1427 1585 1428 1589
rect 1422 1584 1428 1585
rect 1478 1589 1484 1590
rect 1478 1585 1479 1589
rect 1483 1585 1484 1589
rect 1478 1584 1484 1585
rect 1558 1589 1564 1590
rect 1558 1585 1559 1589
rect 1563 1585 1564 1589
rect 1558 1584 1564 1585
rect 1638 1589 1644 1590
rect 1638 1585 1639 1589
rect 1643 1585 1644 1589
rect 1638 1584 1644 1585
rect 1718 1589 1724 1590
rect 1718 1585 1719 1589
rect 1723 1585 1724 1589
rect 1718 1584 1724 1585
rect 1790 1589 1796 1590
rect 1790 1585 1791 1589
rect 1795 1585 1796 1589
rect 1790 1584 1796 1585
rect 1870 1589 1876 1590
rect 1870 1585 1871 1589
rect 1875 1585 1876 1589
rect 1870 1584 1876 1585
rect 1950 1589 1956 1590
rect 1950 1585 1951 1589
rect 1955 1585 1956 1589
rect 1950 1584 1956 1585
rect 2030 1589 2036 1590
rect 2030 1585 2031 1589
rect 2035 1585 2036 1589
rect 2030 1584 2036 1585
rect 2502 1588 2508 1589
rect 2502 1584 2503 1588
rect 2507 1584 2508 1588
rect 1326 1583 1332 1584
rect 2502 1583 2508 1584
rect 110 1575 116 1576
rect 110 1571 111 1575
rect 115 1571 116 1575
rect 1286 1575 1292 1576
rect 110 1570 116 1571
rect 286 1572 292 1573
rect 286 1568 287 1572
rect 291 1568 292 1572
rect 286 1567 292 1568
rect 342 1572 348 1573
rect 342 1568 343 1572
rect 347 1568 348 1572
rect 342 1567 348 1568
rect 414 1572 420 1573
rect 414 1568 415 1572
rect 419 1568 420 1572
rect 414 1567 420 1568
rect 494 1572 500 1573
rect 494 1568 495 1572
rect 499 1568 500 1572
rect 494 1567 500 1568
rect 582 1572 588 1573
rect 582 1568 583 1572
rect 587 1568 588 1572
rect 582 1567 588 1568
rect 678 1572 684 1573
rect 678 1568 679 1572
rect 683 1568 684 1572
rect 678 1567 684 1568
rect 774 1572 780 1573
rect 774 1568 775 1572
rect 779 1568 780 1572
rect 774 1567 780 1568
rect 878 1572 884 1573
rect 878 1568 879 1572
rect 883 1568 884 1572
rect 878 1567 884 1568
rect 990 1572 996 1573
rect 990 1568 991 1572
rect 995 1568 996 1572
rect 990 1567 996 1568
rect 1102 1572 1108 1573
rect 1102 1568 1103 1572
rect 1107 1568 1108 1572
rect 1286 1571 1287 1575
rect 1291 1571 1292 1575
rect 1286 1570 1292 1571
rect 1326 1571 1332 1572
rect 1102 1567 1108 1568
rect 1326 1567 1327 1571
rect 1331 1567 1332 1571
rect 2502 1571 2508 1572
rect 1326 1566 1332 1567
rect 1350 1568 1356 1569
rect 1350 1564 1351 1568
rect 1355 1564 1356 1568
rect 1350 1563 1356 1564
rect 1406 1568 1412 1569
rect 1406 1564 1407 1568
rect 1411 1564 1412 1568
rect 1406 1563 1412 1564
rect 1462 1568 1468 1569
rect 1462 1564 1463 1568
rect 1467 1564 1468 1568
rect 1462 1563 1468 1564
rect 1542 1568 1548 1569
rect 1542 1564 1543 1568
rect 1547 1564 1548 1568
rect 1542 1563 1548 1564
rect 1622 1568 1628 1569
rect 1622 1564 1623 1568
rect 1627 1564 1628 1568
rect 1622 1563 1628 1564
rect 1702 1568 1708 1569
rect 1702 1564 1703 1568
rect 1707 1564 1708 1568
rect 1702 1563 1708 1564
rect 1774 1568 1780 1569
rect 1774 1564 1775 1568
rect 1779 1564 1780 1568
rect 1774 1563 1780 1564
rect 1854 1568 1860 1569
rect 1854 1564 1855 1568
rect 1859 1564 1860 1568
rect 1854 1563 1860 1564
rect 1934 1568 1940 1569
rect 1934 1564 1935 1568
rect 1939 1564 1940 1568
rect 1934 1563 1940 1564
rect 2014 1568 2020 1569
rect 2014 1564 2015 1568
rect 2019 1564 2020 1568
rect 2502 1567 2503 1571
rect 2507 1567 2508 1571
rect 2502 1566 2508 1567
rect 2014 1563 2020 1564
rect 246 1560 252 1561
rect 110 1557 116 1558
rect 110 1553 111 1557
rect 115 1553 116 1557
rect 246 1556 247 1560
rect 251 1556 252 1560
rect 246 1555 252 1556
rect 318 1560 324 1561
rect 318 1556 319 1560
rect 323 1556 324 1560
rect 318 1555 324 1556
rect 398 1560 404 1561
rect 398 1556 399 1560
rect 403 1556 404 1560
rect 398 1555 404 1556
rect 486 1560 492 1561
rect 486 1556 487 1560
rect 491 1556 492 1560
rect 486 1555 492 1556
rect 582 1560 588 1561
rect 582 1556 583 1560
rect 587 1556 588 1560
rect 582 1555 588 1556
rect 670 1560 676 1561
rect 670 1556 671 1560
rect 675 1556 676 1560
rect 670 1555 676 1556
rect 758 1560 764 1561
rect 758 1556 759 1560
rect 763 1556 764 1560
rect 758 1555 764 1556
rect 846 1560 852 1561
rect 846 1556 847 1560
rect 851 1556 852 1560
rect 846 1555 852 1556
rect 926 1560 932 1561
rect 926 1556 927 1560
rect 931 1556 932 1560
rect 926 1555 932 1556
rect 1006 1560 1012 1561
rect 1006 1556 1007 1560
rect 1011 1556 1012 1560
rect 1006 1555 1012 1556
rect 1086 1560 1092 1561
rect 1086 1556 1087 1560
rect 1091 1556 1092 1560
rect 1086 1555 1092 1556
rect 1166 1560 1172 1561
rect 1166 1556 1167 1560
rect 1171 1556 1172 1560
rect 1166 1555 1172 1556
rect 1222 1560 1228 1561
rect 1222 1556 1223 1560
rect 1227 1556 1228 1560
rect 1222 1555 1228 1556
rect 1286 1557 1292 1558
rect 110 1552 116 1553
rect 1286 1553 1287 1557
rect 1291 1553 1292 1557
rect 1350 1556 1356 1557
rect 1286 1552 1292 1553
rect 1326 1553 1332 1554
rect 1326 1549 1327 1553
rect 1331 1549 1332 1553
rect 1350 1552 1351 1556
rect 1355 1552 1356 1556
rect 1350 1551 1356 1552
rect 1470 1556 1476 1557
rect 1470 1552 1471 1556
rect 1475 1552 1476 1556
rect 1470 1551 1476 1552
rect 1606 1556 1612 1557
rect 1606 1552 1607 1556
rect 1611 1552 1612 1556
rect 1606 1551 1612 1552
rect 1734 1556 1740 1557
rect 1734 1552 1735 1556
rect 1739 1552 1740 1556
rect 1734 1551 1740 1552
rect 1870 1556 1876 1557
rect 1870 1552 1871 1556
rect 1875 1552 1876 1556
rect 1870 1551 1876 1552
rect 2006 1556 2012 1557
rect 2006 1552 2007 1556
rect 2011 1552 2012 1556
rect 2006 1551 2012 1552
rect 2502 1553 2508 1554
rect 1326 1548 1332 1549
rect 2502 1549 2503 1553
rect 2507 1549 2508 1553
rect 2502 1548 2508 1549
rect 110 1540 116 1541
rect 1286 1540 1292 1541
rect 110 1536 111 1540
rect 115 1536 116 1540
rect 110 1535 116 1536
rect 262 1539 268 1540
rect 262 1535 263 1539
rect 267 1535 268 1539
rect 262 1534 268 1535
rect 334 1539 340 1540
rect 334 1535 335 1539
rect 339 1535 340 1539
rect 334 1534 340 1535
rect 414 1539 420 1540
rect 414 1535 415 1539
rect 419 1535 420 1539
rect 414 1534 420 1535
rect 502 1539 508 1540
rect 502 1535 503 1539
rect 507 1535 508 1539
rect 502 1534 508 1535
rect 598 1539 604 1540
rect 598 1535 599 1539
rect 603 1535 604 1539
rect 598 1534 604 1535
rect 686 1539 692 1540
rect 686 1535 687 1539
rect 691 1535 692 1539
rect 686 1534 692 1535
rect 774 1539 780 1540
rect 774 1535 775 1539
rect 779 1535 780 1539
rect 774 1534 780 1535
rect 862 1539 868 1540
rect 862 1535 863 1539
rect 867 1535 868 1539
rect 862 1534 868 1535
rect 942 1539 948 1540
rect 942 1535 943 1539
rect 947 1535 948 1539
rect 942 1534 948 1535
rect 1022 1539 1028 1540
rect 1022 1535 1023 1539
rect 1027 1535 1028 1539
rect 1022 1534 1028 1535
rect 1102 1539 1108 1540
rect 1102 1535 1103 1539
rect 1107 1535 1108 1539
rect 1102 1534 1108 1535
rect 1182 1539 1188 1540
rect 1182 1535 1183 1539
rect 1187 1535 1188 1539
rect 1182 1534 1188 1535
rect 1238 1539 1244 1540
rect 1238 1535 1239 1539
rect 1243 1535 1244 1539
rect 1286 1536 1287 1540
rect 1291 1536 1292 1540
rect 1286 1535 1292 1536
rect 1326 1536 1332 1537
rect 2502 1536 2508 1537
rect 1238 1534 1244 1535
rect 1326 1532 1327 1536
rect 1331 1532 1332 1536
rect 1326 1531 1332 1532
rect 1366 1535 1372 1536
rect 1366 1531 1367 1535
rect 1371 1531 1372 1535
rect 1366 1530 1372 1531
rect 1486 1535 1492 1536
rect 1486 1531 1487 1535
rect 1491 1531 1492 1535
rect 1486 1530 1492 1531
rect 1622 1535 1628 1536
rect 1622 1531 1623 1535
rect 1627 1531 1628 1535
rect 1622 1530 1628 1531
rect 1750 1535 1756 1536
rect 1750 1531 1751 1535
rect 1755 1531 1756 1535
rect 1750 1530 1756 1531
rect 1886 1535 1892 1536
rect 1886 1531 1887 1535
rect 1891 1531 1892 1535
rect 1886 1530 1892 1531
rect 2022 1535 2028 1536
rect 2022 1531 2023 1535
rect 2027 1531 2028 1535
rect 2502 1532 2503 1536
rect 2507 1532 2508 1536
rect 2502 1531 2508 1532
rect 2022 1530 2028 1531
rect 1366 1485 1372 1486
rect 1326 1484 1332 1485
rect 278 1481 284 1482
rect 110 1480 116 1481
rect 110 1476 111 1480
rect 115 1476 116 1480
rect 278 1477 279 1481
rect 283 1477 284 1481
rect 278 1476 284 1477
rect 342 1481 348 1482
rect 342 1477 343 1481
rect 347 1477 348 1481
rect 342 1476 348 1477
rect 414 1481 420 1482
rect 414 1477 415 1481
rect 419 1477 420 1481
rect 414 1476 420 1477
rect 494 1481 500 1482
rect 494 1477 495 1481
rect 499 1477 500 1481
rect 494 1476 500 1477
rect 574 1481 580 1482
rect 574 1477 575 1481
rect 579 1477 580 1481
rect 574 1476 580 1477
rect 654 1481 660 1482
rect 654 1477 655 1481
rect 659 1477 660 1481
rect 654 1476 660 1477
rect 734 1481 740 1482
rect 734 1477 735 1481
rect 739 1477 740 1481
rect 734 1476 740 1477
rect 814 1481 820 1482
rect 814 1477 815 1481
rect 819 1477 820 1481
rect 814 1476 820 1477
rect 894 1481 900 1482
rect 894 1477 895 1481
rect 899 1477 900 1481
rect 894 1476 900 1477
rect 974 1481 980 1482
rect 974 1477 975 1481
rect 979 1477 980 1481
rect 974 1476 980 1477
rect 1054 1481 1060 1482
rect 1054 1477 1055 1481
rect 1059 1477 1060 1481
rect 1054 1476 1060 1477
rect 1142 1481 1148 1482
rect 1142 1477 1143 1481
rect 1147 1477 1148 1481
rect 1142 1476 1148 1477
rect 1286 1480 1292 1481
rect 1286 1476 1287 1480
rect 1291 1476 1292 1480
rect 1326 1480 1327 1484
rect 1331 1480 1332 1484
rect 1366 1481 1367 1485
rect 1371 1481 1372 1485
rect 1366 1480 1372 1481
rect 1422 1485 1428 1486
rect 1422 1481 1423 1485
rect 1427 1481 1428 1485
rect 1422 1480 1428 1481
rect 1478 1485 1484 1486
rect 1478 1481 1479 1485
rect 1483 1481 1484 1485
rect 1478 1480 1484 1481
rect 1550 1485 1556 1486
rect 1550 1481 1551 1485
rect 1555 1481 1556 1485
rect 1550 1480 1556 1481
rect 1630 1485 1636 1486
rect 1630 1481 1631 1485
rect 1635 1481 1636 1485
rect 1630 1480 1636 1481
rect 1710 1485 1716 1486
rect 1710 1481 1711 1485
rect 1715 1481 1716 1485
rect 1710 1480 1716 1481
rect 1790 1485 1796 1486
rect 1790 1481 1791 1485
rect 1795 1481 1796 1485
rect 1790 1480 1796 1481
rect 1870 1485 1876 1486
rect 1870 1481 1871 1485
rect 1875 1481 1876 1485
rect 1870 1480 1876 1481
rect 1950 1485 1956 1486
rect 1950 1481 1951 1485
rect 1955 1481 1956 1485
rect 1950 1480 1956 1481
rect 2030 1485 2036 1486
rect 2030 1481 2031 1485
rect 2035 1481 2036 1485
rect 2030 1480 2036 1481
rect 2118 1485 2124 1486
rect 2118 1481 2119 1485
rect 2123 1481 2124 1485
rect 2118 1480 2124 1481
rect 2502 1484 2508 1485
rect 2502 1480 2503 1484
rect 2507 1480 2508 1484
rect 1326 1479 1332 1480
rect 2502 1479 2508 1480
rect 110 1475 116 1476
rect 1286 1475 1292 1476
rect 1326 1467 1332 1468
rect 110 1463 116 1464
rect 110 1459 111 1463
rect 115 1459 116 1463
rect 1286 1463 1292 1464
rect 110 1458 116 1459
rect 262 1460 268 1461
rect 262 1456 263 1460
rect 267 1456 268 1460
rect 262 1455 268 1456
rect 326 1460 332 1461
rect 326 1456 327 1460
rect 331 1456 332 1460
rect 326 1455 332 1456
rect 398 1460 404 1461
rect 398 1456 399 1460
rect 403 1456 404 1460
rect 398 1455 404 1456
rect 478 1460 484 1461
rect 478 1456 479 1460
rect 483 1456 484 1460
rect 478 1455 484 1456
rect 558 1460 564 1461
rect 558 1456 559 1460
rect 563 1456 564 1460
rect 558 1455 564 1456
rect 638 1460 644 1461
rect 638 1456 639 1460
rect 643 1456 644 1460
rect 638 1455 644 1456
rect 718 1460 724 1461
rect 718 1456 719 1460
rect 723 1456 724 1460
rect 718 1455 724 1456
rect 798 1460 804 1461
rect 798 1456 799 1460
rect 803 1456 804 1460
rect 798 1455 804 1456
rect 878 1460 884 1461
rect 878 1456 879 1460
rect 883 1456 884 1460
rect 878 1455 884 1456
rect 958 1460 964 1461
rect 958 1456 959 1460
rect 963 1456 964 1460
rect 958 1455 964 1456
rect 1038 1460 1044 1461
rect 1038 1456 1039 1460
rect 1043 1456 1044 1460
rect 1038 1455 1044 1456
rect 1126 1460 1132 1461
rect 1126 1456 1127 1460
rect 1131 1456 1132 1460
rect 1286 1459 1287 1463
rect 1291 1459 1292 1463
rect 1326 1463 1327 1467
rect 1331 1463 1332 1467
rect 2502 1467 2508 1468
rect 1326 1462 1332 1463
rect 1350 1464 1356 1465
rect 1350 1460 1351 1464
rect 1355 1460 1356 1464
rect 1350 1459 1356 1460
rect 1406 1464 1412 1465
rect 1406 1460 1407 1464
rect 1411 1460 1412 1464
rect 1406 1459 1412 1460
rect 1462 1464 1468 1465
rect 1462 1460 1463 1464
rect 1467 1460 1468 1464
rect 1462 1459 1468 1460
rect 1534 1464 1540 1465
rect 1534 1460 1535 1464
rect 1539 1460 1540 1464
rect 1534 1459 1540 1460
rect 1614 1464 1620 1465
rect 1614 1460 1615 1464
rect 1619 1460 1620 1464
rect 1614 1459 1620 1460
rect 1694 1464 1700 1465
rect 1694 1460 1695 1464
rect 1699 1460 1700 1464
rect 1694 1459 1700 1460
rect 1774 1464 1780 1465
rect 1774 1460 1775 1464
rect 1779 1460 1780 1464
rect 1774 1459 1780 1460
rect 1854 1464 1860 1465
rect 1854 1460 1855 1464
rect 1859 1460 1860 1464
rect 1854 1459 1860 1460
rect 1934 1464 1940 1465
rect 1934 1460 1935 1464
rect 1939 1460 1940 1464
rect 1934 1459 1940 1460
rect 2014 1464 2020 1465
rect 2014 1460 2015 1464
rect 2019 1460 2020 1464
rect 2014 1459 2020 1460
rect 2102 1464 2108 1465
rect 2102 1460 2103 1464
rect 2107 1460 2108 1464
rect 2502 1463 2503 1467
rect 2507 1463 2508 1467
rect 2502 1462 2508 1463
rect 2102 1459 2108 1460
rect 1286 1458 1292 1459
rect 1126 1455 1132 1456
rect 190 1444 196 1445
rect 110 1441 116 1442
rect 110 1437 111 1441
rect 115 1437 116 1441
rect 190 1440 191 1444
rect 195 1440 196 1444
rect 190 1439 196 1440
rect 254 1444 260 1445
rect 254 1440 255 1444
rect 259 1440 260 1444
rect 254 1439 260 1440
rect 326 1444 332 1445
rect 326 1440 327 1444
rect 331 1440 332 1444
rect 326 1439 332 1440
rect 406 1444 412 1445
rect 406 1440 407 1444
rect 411 1440 412 1444
rect 406 1439 412 1440
rect 502 1444 508 1445
rect 502 1440 503 1444
rect 507 1440 508 1444
rect 502 1439 508 1440
rect 606 1444 612 1445
rect 606 1440 607 1444
rect 611 1440 612 1444
rect 606 1439 612 1440
rect 710 1444 716 1445
rect 710 1440 711 1444
rect 715 1440 716 1444
rect 710 1439 716 1440
rect 814 1444 820 1445
rect 814 1440 815 1444
rect 819 1440 820 1444
rect 814 1439 820 1440
rect 918 1444 924 1445
rect 918 1440 919 1444
rect 923 1440 924 1444
rect 918 1439 924 1440
rect 1022 1444 1028 1445
rect 1022 1440 1023 1444
rect 1027 1440 1028 1444
rect 1022 1439 1028 1440
rect 1126 1444 1132 1445
rect 1126 1440 1127 1444
rect 1131 1440 1132 1444
rect 1126 1439 1132 1440
rect 1222 1444 1228 1445
rect 1222 1440 1223 1444
rect 1227 1440 1228 1444
rect 1358 1444 1364 1445
rect 1222 1439 1228 1440
rect 1286 1441 1292 1442
rect 110 1436 116 1437
rect 1286 1437 1287 1441
rect 1291 1437 1292 1441
rect 1286 1436 1292 1437
rect 1326 1441 1332 1442
rect 1326 1437 1327 1441
rect 1331 1437 1332 1441
rect 1358 1440 1359 1444
rect 1363 1440 1364 1444
rect 1358 1439 1364 1440
rect 1446 1444 1452 1445
rect 1446 1440 1447 1444
rect 1451 1440 1452 1444
rect 1446 1439 1452 1440
rect 1534 1444 1540 1445
rect 1534 1440 1535 1444
rect 1539 1440 1540 1444
rect 1534 1439 1540 1440
rect 1630 1444 1636 1445
rect 1630 1440 1631 1444
rect 1635 1440 1636 1444
rect 1630 1439 1636 1440
rect 1726 1444 1732 1445
rect 1726 1440 1727 1444
rect 1731 1440 1732 1444
rect 1726 1439 1732 1440
rect 1814 1444 1820 1445
rect 1814 1440 1815 1444
rect 1819 1440 1820 1444
rect 1814 1439 1820 1440
rect 1902 1444 1908 1445
rect 1902 1440 1903 1444
rect 1907 1440 1908 1444
rect 1902 1439 1908 1440
rect 1990 1444 1996 1445
rect 1990 1440 1991 1444
rect 1995 1440 1996 1444
rect 1990 1439 1996 1440
rect 2070 1444 2076 1445
rect 2070 1440 2071 1444
rect 2075 1440 2076 1444
rect 2070 1439 2076 1440
rect 2158 1444 2164 1445
rect 2158 1440 2159 1444
rect 2163 1440 2164 1444
rect 2158 1439 2164 1440
rect 2246 1444 2252 1445
rect 2246 1440 2247 1444
rect 2251 1440 2252 1444
rect 2246 1439 2252 1440
rect 2502 1441 2508 1442
rect 1326 1436 1332 1437
rect 2502 1437 2503 1441
rect 2507 1437 2508 1441
rect 2502 1436 2508 1437
rect 110 1424 116 1425
rect 1286 1424 1292 1425
rect 110 1420 111 1424
rect 115 1420 116 1424
rect 110 1419 116 1420
rect 206 1423 212 1424
rect 206 1419 207 1423
rect 211 1419 212 1423
rect 206 1418 212 1419
rect 270 1423 276 1424
rect 270 1419 271 1423
rect 275 1419 276 1423
rect 270 1418 276 1419
rect 342 1423 348 1424
rect 342 1419 343 1423
rect 347 1419 348 1423
rect 342 1418 348 1419
rect 422 1423 428 1424
rect 422 1419 423 1423
rect 427 1419 428 1423
rect 422 1418 428 1419
rect 518 1423 524 1424
rect 518 1419 519 1423
rect 523 1419 524 1423
rect 518 1418 524 1419
rect 622 1423 628 1424
rect 622 1419 623 1423
rect 627 1419 628 1423
rect 622 1418 628 1419
rect 726 1423 732 1424
rect 726 1419 727 1423
rect 731 1419 732 1423
rect 726 1418 732 1419
rect 830 1423 836 1424
rect 830 1419 831 1423
rect 835 1419 836 1423
rect 830 1418 836 1419
rect 934 1423 940 1424
rect 934 1419 935 1423
rect 939 1419 940 1423
rect 934 1418 940 1419
rect 1038 1423 1044 1424
rect 1038 1419 1039 1423
rect 1043 1419 1044 1423
rect 1038 1418 1044 1419
rect 1142 1423 1148 1424
rect 1142 1419 1143 1423
rect 1147 1419 1148 1423
rect 1142 1418 1148 1419
rect 1238 1423 1244 1424
rect 1238 1419 1239 1423
rect 1243 1419 1244 1423
rect 1286 1420 1287 1424
rect 1291 1420 1292 1424
rect 1286 1419 1292 1420
rect 1326 1424 1332 1425
rect 2502 1424 2508 1425
rect 1326 1420 1327 1424
rect 1331 1420 1332 1424
rect 1326 1419 1332 1420
rect 1374 1423 1380 1424
rect 1374 1419 1375 1423
rect 1379 1419 1380 1423
rect 1238 1418 1244 1419
rect 1374 1418 1380 1419
rect 1462 1423 1468 1424
rect 1462 1419 1463 1423
rect 1467 1419 1468 1423
rect 1462 1418 1468 1419
rect 1550 1423 1556 1424
rect 1550 1419 1551 1423
rect 1555 1419 1556 1423
rect 1550 1418 1556 1419
rect 1646 1423 1652 1424
rect 1646 1419 1647 1423
rect 1651 1419 1652 1423
rect 1646 1418 1652 1419
rect 1742 1423 1748 1424
rect 1742 1419 1743 1423
rect 1747 1419 1748 1423
rect 1742 1418 1748 1419
rect 1830 1423 1836 1424
rect 1830 1419 1831 1423
rect 1835 1419 1836 1423
rect 1830 1418 1836 1419
rect 1918 1423 1924 1424
rect 1918 1419 1919 1423
rect 1923 1419 1924 1423
rect 1918 1418 1924 1419
rect 2006 1423 2012 1424
rect 2006 1419 2007 1423
rect 2011 1419 2012 1423
rect 2006 1418 2012 1419
rect 2086 1423 2092 1424
rect 2086 1419 2087 1423
rect 2091 1419 2092 1423
rect 2086 1418 2092 1419
rect 2174 1423 2180 1424
rect 2174 1419 2175 1423
rect 2179 1419 2180 1423
rect 2174 1418 2180 1419
rect 2262 1423 2268 1424
rect 2262 1419 2263 1423
rect 2267 1419 2268 1423
rect 2502 1420 2503 1424
rect 2507 1420 2508 1424
rect 2502 1419 2508 1420
rect 2262 1418 2268 1419
rect 1566 1373 1572 1374
rect 1326 1372 1332 1373
rect 150 1369 156 1370
rect 110 1368 116 1369
rect 110 1364 111 1368
rect 115 1364 116 1368
rect 150 1365 151 1369
rect 155 1365 156 1369
rect 150 1364 156 1365
rect 222 1369 228 1370
rect 222 1365 223 1369
rect 227 1365 228 1369
rect 222 1364 228 1365
rect 294 1369 300 1370
rect 294 1365 295 1369
rect 299 1365 300 1369
rect 294 1364 300 1365
rect 358 1369 364 1370
rect 358 1365 359 1369
rect 363 1365 364 1369
rect 358 1364 364 1365
rect 430 1369 436 1370
rect 430 1365 431 1369
rect 435 1365 436 1369
rect 430 1364 436 1365
rect 502 1369 508 1370
rect 502 1365 503 1369
rect 507 1365 508 1369
rect 502 1364 508 1365
rect 582 1369 588 1370
rect 582 1365 583 1369
rect 587 1365 588 1369
rect 582 1364 588 1365
rect 662 1369 668 1370
rect 662 1365 663 1369
rect 667 1365 668 1369
rect 662 1364 668 1365
rect 750 1369 756 1370
rect 750 1365 751 1369
rect 755 1365 756 1369
rect 750 1364 756 1365
rect 838 1369 844 1370
rect 838 1365 839 1369
rect 843 1365 844 1369
rect 838 1364 844 1365
rect 926 1369 932 1370
rect 926 1365 927 1369
rect 931 1365 932 1369
rect 926 1364 932 1365
rect 1014 1369 1020 1370
rect 1014 1365 1015 1369
rect 1019 1365 1020 1369
rect 1014 1364 1020 1365
rect 1102 1369 1108 1370
rect 1102 1365 1103 1369
rect 1107 1365 1108 1369
rect 1102 1364 1108 1365
rect 1198 1369 1204 1370
rect 1198 1365 1199 1369
rect 1203 1365 1204 1369
rect 1198 1364 1204 1365
rect 1286 1368 1292 1369
rect 1286 1364 1287 1368
rect 1291 1364 1292 1368
rect 1326 1368 1327 1372
rect 1331 1368 1332 1372
rect 1566 1369 1567 1373
rect 1571 1369 1572 1373
rect 1566 1368 1572 1369
rect 1646 1373 1652 1374
rect 1646 1369 1647 1373
rect 1651 1369 1652 1373
rect 1646 1368 1652 1369
rect 1734 1373 1740 1374
rect 1734 1369 1735 1373
rect 1739 1369 1740 1373
rect 1734 1368 1740 1369
rect 1830 1373 1836 1374
rect 1830 1369 1831 1373
rect 1835 1369 1836 1373
rect 1830 1368 1836 1369
rect 1918 1373 1924 1374
rect 1918 1369 1919 1373
rect 1923 1369 1924 1373
rect 1918 1368 1924 1369
rect 2006 1373 2012 1374
rect 2006 1369 2007 1373
rect 2011 1369 2012 1373
rect 2006 1368 2012 1369
rect 2094 1373 2100 1374
rect 2094 1369 2095 1373
rect 2099 1369 2100 1373
rect 2094 1368 2100 1369
rect 2174 1373 2180 1374
rect 2174 1369 2175 1373
rect 2179 1369 2180 1373
rect 2174 1368 2180 1369
rect 2246 1373 2252 1374
rect 2246 1369 2247 1373
rect 2251 1369 2252 1373
rect 2246 1368 2252 1369
rect 2318 1373 2324 1374
rect 2318 1369 2319 1373
rect 2323 1369 2324 1373
rect 2318 1368 2324 1369
rect 2398 1373 2404 1374
rect 2398 1369 2399 1373
rect 2403 1369 2404 1373
rect 2398 1368 2404 1369
rect 2454 1373 2460 1374
rect 2454 1369 2455 1373
rect 2459 1369 2460 1373
rect 2454 1368 2460 1369
rect 2502 1372 2508 1373
rect 2502 1368 2503 1372
rect 2507 1368 2508 1372
rect 1326 1367 1332 1368
rect 2502 1367 2508 1368
rect 110 1363 116 1364
rect 1286 1363 1292 1364
rect 1326 1355 1332 1356
rect 110 1351 116 1352
rect 110 1347 111 1351
rect 115 1347 116 1351
rect 1286 1351 1292 1352
rect 110 1346 116 1347
rect 134 1348 140 1349
rect 134 1344 135 1348
rect 139 1344 140 1348
rect 134 1343 140 1344
rect 206 1348 212 1349
rect 206 1344 207 1348
rect 211 1344 212 1348
rect 206 1343 212 1344
rect 278 1348 284 1349
rect 278 1344 279 1348
rect 283 1344 284 1348
rect 278 1343 284 1344
rect 342 1348 348 1349
rect 342 1344 343 1348
rect 347 1344 348 1348
rect 342 1343 348 1344
rect 414 1348 420 1349
rect 414 1344 415 1348
rect 419 1344 420 1348
rect 414 1343 420 1344
rect 486 1348 492 1349
rect 486 1344 487 1348
rect 491 1344 492 1348
rect 486 1343 492 1344
rect 566 1348 572 1349
rect 566 1344 567 1348
rect 571 1344 572 1348
rect 566 1343 572 1344
rect 646 1348 652 1349
rect 646 1344 647 1348
rect 651 1344 652 1348
rect 646 1343 652 1344
rect 734 1348 740 1349
rect 734 1344 735 1348
rect 739 1344 740 1348
rect 734 1343 740 1344
rect 822 1348 828 1349
rect 822 1344 823 1348
rect 827 1344 828 1348
rect 822 1343 828 1344
rect 910 1348 916 1349
rect 910 1344 911 1348
rect 915 1344 916 1348
rect 910 1343 916 1344
rect 998 1348 1004 1349
rect 998 1344 999 1348
rect 1003 1344 1004 1348
rect 998 1343 1004 1344
rect 1086 1348 1092 1349
rect 1086 1344 1087 1348
rect 1091 1344 1092 1348
rect 1086 1343 1092 1344
rect 1182 1348 1188 1349
rect 1182 1344 1183 1348
rect 1187 1344 1188 1348
rect 1286 1347 1287 1351
rect 1291 1347 1292 1351
rect 1326 1351 1327 1355
rect 1331 1351 1332 1355
rect 2502 1355 2508 1356
rect 1326 1350 1332 1351
rect 1550 1352 1556 1353
rect 1550 1348 1551 1352
rect 1555 1348 1556 1352
rect 1550 1347 1556 1348
rect 1630 1352 1636 1353
rect 1630 1348 1631 1352
rect 1635 1348 1636 1352
rect 1630 1347 1636 1348
rect 1718 1352 1724 1353
rect 1718 1348 1719 1352
rect 1723 1348 1724 1352
rect 1718 1347 1724 1348
rect 1814 1352 1820 1353
rect 1814 1348 1815 1352
rect 1819 1348 1820 1352
rect 1814 1347 1820 1348
rect 1902 1352 1908 1353
rect 1902 1348 1903 1352
rect 1907 1348 1908 1352
rect 1902 1347 1908 1348
rect 1990 1352 1996 1353
rect 1990 1348 1991 1352
rect 1995 1348 1996 1352
rect 1990 1347 1996 1348
rect 2078 1352 2084 1353
rect 2078 1348 2079 1352
rect 2083 1348 2084 1352
rect 2078 1347 2084 1348
rect 2158 1352 2164 1353
rect 2158 1348 2159 1352
rect 2163 1348 2164 1352
rect 2158 1347 2164 1348
rect 2230 1352 2236 1353
rect 2230 1348 2231 1352
rect 2235 1348 2236 1352
rect 2230 1347 2236 1348
rect 2302 1352 2308 1353
rect 2302 1348 2303 1352
rect 2307 1348 2308 1352
rect 2302 1347 2308 1348
rect 2382 1352 2388 1353
rect 2382 1348 2383 1352
rect 2387 1348 2388 1352
rect 2382 1347 2388 1348
rect 2438 1352 2444 1353
rect 2438 1348 2439 1352
rect 2443 1348 2444 1352
rect 2502 1351 2503 1355
rect 2507 1351 2508 1355
rect 2502 1350 2508 1351
rect 2438 1347 2444 1348
rect 1286 1346 1292 1347
rect 1182 1343 1188 1344
rect 1582 1340 1588 1341
rect 1326 1337 1332 1338
rect 1326 1333 1327 1337
rect 1331 1333 1332 1337
rect 1582 1336 1583 1340
rect 1587 1336 1588 1340
rect 1582 1335 1588 1336
rect 1646 1340 1652 1341
rect 1646 1336 1647 1340
rect 1651 1336 1652 1340
rect 1646 1335 1652 1336
rect 1726 1340 1732 1341
rect 1726 1336 1727 1340
rect 1731 1336 1732 1340
rect 1726 1335 1732 1336
rect 1806 1340 1812 1341
rect 1806 1336 1807 1340
rect 1811 1336 1812 1340
rect 1806 1335 1812 1336
rect 1894 1340 1900 1341
rect 1894 1336 1895 1340
rect 1899 1336 1900 1340
rect 1894 1335 1900 1336
rect 1982 1340 1988 1341
rect 1982 1336 1983 1340
rect 1987 1336 1988 1340
rect 1982 1335 1988 1336
rect 2062 1340 2068 1341
rect 2062 1336 2063 1340
rect 2067 1336 2068 1340
rect 2062 1335 2068 1336
rect 2142 1340 2148 1341
rect 2142 1336 2143 1340
rect 2147 1336 2148 1340
rect 2142 1335 2148 1336
rect 2222 1340 2228 1341
rect 2222 1336 2223 1340
rect 2227 1336 2228 1340
rect 2222 1335 2228 1336
rect 2302 1340 2308 1341
rect 2302 1336 2303 1340
rect 2307 1336 2308 1340
rect 2302 1335 2308 1336
rect 2382 1340 2388 1341
rect 2382 1336 2383 1340
rect 2387 1336 2388 1340
rect 2382 1335 2388 1336
rect 2438 1340 2444 1341
rect 2438 1336 2439 1340
rect 2443 1336 2444 1340
rect 2438 1335 2444 1336
rect 2502 1337 2508 1338
rect 1326 1332 1332 1333
rect 2502 1333 2503 1337
rect 2507 1333 2508 1337
rect 2502 1332 2508 1333
rect 134 1320 140 1321
rect 110 1317 116 1318
rect 110 1313 111 1317
rect 115 1313 116 1317
rect 134 1316 135 1320
rect 139 1316 140 1320
rect 134 1315 140 1316
rect 238 1320 244 1321
rect 238 1316 239 1320
rect 243 1316 244 1320
rect 238 1315 244 1316
rect 366 1320 372 1321
rect 366 1316 367 1320
rect 371 1316 372 1320
rect 366 1315 372 1316
rect 478 1320 484 1321
rect 478 1316 479 1320
rect 483 1316 484 1320
rect 478 1315 484 1316
rect 582 1320 588 1321
rect 582 1316 583 1320
rect 587 1316 588 1320
rect 582 1315 588 1316
rect 686 1320 692 1321
rect 686 1316 687 1320
rect 691 1316 692 1320
rect 686 1315 692 1316
rect 782 1320 788 1321
rect 782 1316 783 1320
rect 787 1316 788 1320
rect 782 1315 788 1316
rect 878 1320 884 1321
rect 878 1316 879 1320
rect 883 1316 884 1320
rect 878 1315 884 1316
rect 974 1320 980 1321
rect 974 1316 975 1320
rect 979 1316 980 1320
rect 1326 1320 1332 1321
rect 2502 1320 2508 1321
rect 974 1315 980 1316
rect 1286 1317 1292 1318
rect 110 1312 116 1313
rect 1286 1313 1287 1317
rect 1291 1313 1292 1317
rect 1326 1316 1327 1320
rect 1331 1316 1332 1320
rect 1326 1315 1332 1316
rect 1598 1319 1604 1320
rect 1598 1315 1599 1319
rect 1603 1315 1604 1319
rect 1598 1314 1604 1315
rect 1662 1319 1668 1320
rect 1662 1315 1663 1319
rect 1667 1315 1668 1319
rect 1662 1314 1668 1315
rect 1742 1319 1748 1320
rect 1742 1315 1743 1319
rect 1747 1315 1748 1319
rect 1742 1314 1748 1315
rect 1822 1319 1828 1320
rect 1822 1315 1823 1319
rect 1827 1315 1828 1319
rect 1822 1314 1828 1315
rect 1910 1319 1916 1320
rect 1910 1315 1911 1319
rect 1915 1315 1916 1319
rect 1910 1314 1916 1315
rect 1998 1319 2004 1320
rect 1998 1315 1999 1319
rect 2003 1315 2004 1319
rect 1998 1314 2004 1315
rect 2078 1319 2084 1320
rect 2078 1315 2079 1319
rect 2083 1315 2084 1319
rect 2078 1314 2084 1315
rect 2158 1319 2164 1320
rect 2158 1315 2159 1319
rect 2163 1315 2164 1319
rect 2158 1314 2164 1315
rect 2238 1319 2244 1320
rect 2238 1315 2239 1319
rect 2243 1315 2244 1319
rect 2238 1314 2244 1315
rect 2318 1319 2324 1320
rect 2318 1315 2319 1319
rect 2323 1315 2324 1319
rect 2318 1314 2324 1315
rect 2398 1319 2404 1320
rect 2398 1315 2399 1319
rect 2403 1315 2404 1319
rect 2398 1314 2404 1315
rect 2454 1319 2460 1320
rect 2454 1315 2455 1319
rect 2459 1315 2460 1319
rect 2502 1316 2503 1320
rect 2507 1316 2508 1320
rect 2502 1315 2508 1316
rect 2454 1314 2460 1315
rect 1286 1312 1292 1313
rect 110 1300 116 1301
rect 1286 1300 1292 1301
rect 110 1296 111 1300
rect 115 1296 116 1300
rect 110 1295 116 1296
rect 150 1299 156 1300
rect 150 1295 151 1299
rect 155 1295 156 1299
rect 150 1294 156 1295
rect 254 1299 260 1300
rect 254 1295 255 1299
rect 259 1295 260 1299
rect 254 1294 260 1295
rect 382 1299 388 1300
rect 382 1295 383 1299
rect 387 1295 388 1299
rect 382 1294 388 1295
rect 494 1299 500 1300
rect 494 1295 495 1299
rect 499 1295 500 1299
rect 494 1294 500 1295
rect 598 1299 604 1300
rect 598 1295 599 1299
rect 603 1295 604 1299
rect 598 1294 604 1295
rect 702 1299 708 1300
rect 702 1295 703 1299
rect 707 1295 708 1299
rect 702 1294 708 1295
rect 798 1299 804 1300
rect 798 1295 799 1299
rect 803 1295 804 1299
rect 798 1294 804 1295
rect 894 1299 900 1300
rect 894 1295 895 1299
rect 899 1295 900 1299
rect 894 1294 900 1295
rect 990 1299 996 1300
rect 990 1295 991 1299
rect 995 1295 996 1299
rect 1286 1296 1287 1300
rect 1291 1296 1292 1300
rect 1286 1295 1292 1296
rect 990 1294 996 1295
rect 1566 1269 1572 1270
rect 1326 1268 1332 1269
rect 1326 1264 1327 1268
rect 1331 1264 1332 1268
rect 1566 1265 1567 1269
rect 1571 1265 1572 1269
rect 1566 1264 1572 1265
rect 1630 1269 1636 1270
rect 1630 1265 1631 1269
rect 1635 1265 1636 1269
rect 1630 1264 1636 1265
rect 1710 1269 1716 1270
rect 1710 1265 1711 1269
rect 1715 1265 1716 1269
rect 1710 1264 1716 1265
rect 1798 1269 1804 1270
rect 1798 1265 1799 1269
rect 1803 1265 1804 1269
rect 1798 1264 1804 1265
rect 1894 1269 1900 1270
rect 1894 1265 1895 1269
rect 1899 1265 1900 1269
rect 1894 1264 1900 1265
rect 1990 1269 1996 1270
rect 1990 1265 1991 1269
rect 1995 1265 1996 1269
rect 1990 1264 1996 1265
rect 2094 1269 2100 1270
rect 2094 1265 2095 1269
rect 2099 1265 2100 1269
rect 2094 1264 2100 1265
rect 2206 1269 2212 1270
rect 2206 1265 2207 1269
rect 2211 1265 2212 1269
rect 2206 1264 2212 1265
rect 2318 1269 2324 1270
rect 2318 1265 2319 1269
rect 2323 1265 2324 1269
rect 2318 1264 2324 1265
rect 2502 1268 2508 1269
rect 2502 1264 2503 1268
rect 2507 1264 2508 1268
rect 1326 1263 1332 1264
rect 2502 1263 2508 1264
rect 1326 1251 1332 1252
rect 1326 1247 1327 1251
rect 1331 1247 1332 1251
rect 2502 1251 2508 1252
rect 1326 1246 1332 1247
rect 1550 1248 1556 1249
rect 1550 1244 1551 1248
rect 1555 1244 1556 1248
rect 1550 1243 1556 1244
rect 1614 1248 1620 1249
rect 1614 1244 1615 1248
rect 1619 1244 1620 1248
rect 1614 1243 1620 1244
rect 1694 1248 1700 1249
rect 1694 1244 1695 1248
rect 1699 1244 1700 1248
rect 1694 1243 1700 1244
rect 1782 1248 1788 1249
rect 1782 1244 1783 1248
rect 1787 1244 1788 1248
rect 1782 1243 1788 1244
rect 1878 1248 1884 1249
rect 1878 1244 1879 1248
rect 1883 1244 1884 1248
rect 1878 1243 1884 1244
rect 1974 1248 1980 1249
rect 1974 1244 1975 1248
rect 1979 1244 1980 1248
rect 1974 1243 1980 1244
rect 2078 1248 2084 1249
rect 2078 1244 2079 1248
rect 2083 1244 2084 1248
rect 2078 1243 2084 1244
rect 2190 1248 2196 1249
rect 2190 1244 2191 1248
rect 2195 1244 2196 1248
rect 2190 1243 2196 1244
rect 2302 1248 2308 1249
rect 2302 1244 2303 1248
rect 2307 1244 2308 1248
rect 2502 1247 2503 1251
rect 2507 1247 2508 1251
rect 2502 1246 2508 1247
rect 2302 1243 2308 1244
rect 150 1241 156 1242
rect 110 1240 116 1241
rect 110 1236 111 1240
rect 115 1236 116 1240
rect 150 1237 151 1241
rect 155 1237 156 1241
rect 150 1236 156 1237
rect 214 1241 220 1242
rect 214 1237 215 1241
rect 219 1237 220 1241
rect 214 1236 220 1237
rect 302 1241 308 1242
rect 302 1237 303 1241
rect 307 1237 308 1241
rect 302 1236 308 1237
rect 390 1241 396 1242
rect 390 1237 391 1241
rect 395 1237 396 1241
rect 390 1236 396 1237
rect 470 1241 476 1242
rect 470 1237 471 1241
rect 475 1237 476 1241
rect 470 1236 476 1237
rect 550 1241 556 1242
rect 550 1237 551 1241
rect 555 1237 556 1241
rect 550 1236 556 1237
rect 622 1241 628 1242
rect 622 1237 623 1241
rect 627 1237 628 1241
rect 622 1236 628 1237
rect 694 1241 700 1242
rect 694 1237 695 1241
rect 699 1237 700 1241
rect 694 1236 700 1237
rect 766 1241 772 1242
rect 766 1237 767 1241
rect 771 1237 772 1241
rect 766 1236 772 1237
rect 838 1241 844 1242
rect 838 1237 839 1241
rect 843 1237 844 1241
rect 838 1236 844 1237
rect 918 1241 924 1242
rect 918 1237 919 1241
rect 923 1237 924 1241
rect 918 1236 924 1237
rect 1286 1240 1292 1241
rect 1286 1236 1287 1240
rect 1291 1236 1292 1240
rect 110 1235 116 1236
rect 1286 1235 1292 1236
rect 1518 1232 1524 1233
rect 1326 1229 1332 1230
rect 1326 1225 1327 1229
rect 1331 1225 1332 1229
rect 1518 1228 1519 1232
rect 1523 1228 1524 1232
rect 1518 1227 1524 1228
rect 1574 1232 1580 1233
rect 1574 1228 1575 1232
rect 1579 1228 1580 1232
rect 1574 1227 1580 1228
rect 1630 1232 1636 1233
rect 1630 1228 1631 1232
rect 1635 1228 1636 1232
rect 1630 1227 1636 1228
rect 1686 1232 1692 1233
rect 1686 1228 1687 1232
rect 1691 1228 1692 1232
rect 1686 1227 1692 1228
rect 1742 1232 1748 1233
rect 1742 1228 1743 1232
rect 1747 1228 1748 1232
rect 1742 1227 1748 1228
rect 1798 1232 1804 1233
rect 1798 1228 1799 1232
rect 1803 1228 1804 1232
rect 1798 1227 1804 1228
rect 1854 1232 1860 1233
rect 1854 1228 1855 1232
rect 1859 1228 1860 1232
rect 1854 1227 1860 1228
rect 1910 1232 1916 1233
rect 1910 1228 1911 1232
rect 1915 1228 1916 1232
rect 1910 1227 1916 1228
rect 1966 1232 1972 1233
rect 1966 1228 1967 1232
rect 1971 1228 1972 1232
rect 1966 1227 1972 1228
rect 2030 1232 2036 1233
rect 2030 1228 2031 1232
rect 2035 1228 2036 1232
rect 2030 1227 2036 1228
rect 2102 1232 2108 1233
rect 2102 1228 2103 1232
rect 2107 1228 2108 1232
rect 2102 1227 2108 1228
rect 2182 1232 2188 1233
rect 2182 1228 2183 1232
rect 2187 1228 2188 1232
rect 2182 1227 2188 1228
rect 2270 1232 2276 1233
rect 2270 1228 2271 1232
rect 2275 1228 2276 1232
rect 2270 1227 2276 1228
rect 2366 1232 2372 1233
rect 2366 1228 2367 1232
rect 2371 1228 2372 1232
rect 2366 1227 2372 1228
rect 2438 1232 2444 1233
rect 2438 1228 2439 1232
rect 2443 1228 2444 1232
rect 2438 1227 2444 1228
rect 2502 1229 2508 1230
rect 1326 1224 1332 1225
rect 2502 1225 2503 1229
rect 2507 1225 2508 1229
rect 2502 1224 2508 1225
rect 110 1223 116 1224
rect 110 1219 111 1223
rect 115 1219 116 1223
rect 1286 1223 1292 1224
rect 110 1218 116 1219
rect 134 1220 140 1221
rect 134 1216 135 1220
rect 139 1216 140 1220
rect 134 1215 140 1216
rect 198 1220 204 1221
rect 198 1216 199 1220
rect 203 1216 204 1220
rect 198 1215 204 1216
rect 286 1220 292 1221
rect 286 1216 287 1220
rect 291 1216 292 1220
rect 286 1215 292 1216
rect 374 1220 380 1221
rect 374 1216 375 1220
rect 379 1216 380 1220
rect 374 1215 380 1216
rect 454 1220 460 1221
rect 454 1216 455 1220
rect 459 1216 460 1220
rect 454 1215 460 1216
rect 534 1220 540 1221
rect 534 1216 535 1220
rect 539 1216 540 1220
rect 534 1215 540 1216
rect 606 1220 612 1221
rect 606 1216 607 1220
rect 611 1216 612 1220
rect 606 1215 612 1216
rect 678 1220 684 1221
rect 678 1216 679 1220
rect 683 1216 684 1220
rect 678 1215 684 1216
rect 750 1220 756 1221
rect 750 1216 751 1220
rect 755 1216 756 1220
rect 750 1215 756 1216
rect 822 1220 828 1221
rect 822 1216 823 1220
rect 827 1216 828 1220
rect 822 1215 828 1216
rect 902 1220 908 1221
rect 902 1216 903 1220
rect 907 1216 908 1220
rect 1286 1219 1287 1223
rect 1291 1219 1292 1223
rect 1286 1218 1292 1219
rect 902 1215 908 1216
rect 1326 1212 1332 1213
rect 2502 1212 2508 1213
rect 1326 1208 1327 1212
rect 1331 1208 1332 1212
rect 1326 1207 1332 1208
rect 1534 1211 1540 1212
rect 1534 1207 1535 1211
rect 1539 1207 1540 1211
rect 1534 1206 1540 1207
rect 1590 1211 1596 1212
rect 1590 1207 1591 1211
rect 1595 1207 1596 1211
rect 1590 1206 1596 1207
rect 1646 1211 1652 1212
rect 1646 1207 1647 1211
rect 1651 1207 1652 1211
rect 1646 1206 1652 1207
rect 1702 1211 1708 1212
rect 1702 1207 1703 1211
rect 1707 1207 1708 1211
rect 1702 1206 1708 1207
rect 1758 1211 1764 1212
rect 1758 1207 1759 1211
rect 1763 1207 1764 1211
rect 1758 1206 1764 1207
rect 1814 1211 1820 1212
rect 1814 1207 1815 1211
rect 1819 1207 1820 1211
rect 1814 1206 1820 1207
rect 1870 1211 1876 1212
rect 1870 1207 1871 1211
rect 1875 1207 1876 1211
rect 1870 1206 1876 1207
rect 1926 1211 1932 1212
rect 1926 1207 1927 1211
rect 1931 1207 1932 1211
rect 1926 1206 1932 1207
rect 1982 1211 1988 1212
rect 1982 1207 1983 1211
rect 1987 1207 1988 1211
rect 1982 1206 1988 1207
rect 2046 1211 2052 1212
rect 2046 1207 2047 1211
rect 2051 1207 2052 1211
rect 2046 1206 2052 1207
rect 2118 1211 2124 1212
rect 2118 1207 2119 1211
rect 2123 1207 2124 1211
rect 2118 1206 2124 1207
rect 2198 1211 2204 1212
rect 2198 1207 2199 1211
rect 2203 1207 2204 1211
rect 2198 1206 2204 1207
rect 2286 1211 2292 1212
rect 2286 1207 2287 1211
rect 2291 1207 2292 1211
rect 2286 1206 2292 1207
rect 2382 1211 2388 1212
rect 2382 1207 2383 1211
rect 2387 1207 2388 1211
rect 2382 1206 2388 1207
rect 2454 1211 2460 1212
rect 2454 1207 2455 1211
rect 2459 1207 2460 1211
rect 2502 1208 2503 1212
rect 2507 1208 2508 1212
rect 2502 1207 2508 1208
rect 2454 1206 2460 1207
rect 134 1204 140 1205
rect 110 1201 116 1202
rect 110 1197 111 1201
rect 115 1197 116 1201
rect 134 1200 135 1204
rect 139 1200 140 1204
rect 134 1199 140 1200
rect 190 1204 196 1205
rect 190 1200 191 1204
rect 195 1200 196 1204
rect 190 1199 196 1200
rect 270 1204 276 1205
rect 270 1200 271 1204
rect 275 1200 276 1204
rect 270 1199 276 1200
rect 350 1204 356 1205
rect 350 1200 351 1204
rect 355 1200 356 1204
rect 350 1199 356 1200
rect 430 1204 436 1205
rect 430 1200 431 1204
rect 435 1200 436 1204
rect 430 1199 436 1200
rect 510 1204 516 1205
rect 510 1200 511 1204
rect 515 1200 516 1204
rect 510 1199 516 1200
rect 582 1204 588 1205
rect 582 1200 583 1204
rect 587 1200 588 1204
rect 582 1199 588 1200
rect 646 1204 652 1205
rect 646 1200 647 1204
rect 651 1200 652 1204
rect 646 1199 652 1200
rect 718 1204 724 1205
rect 718 1200 719 1204
rect 723 1200 724 1204
rect 718 1199 724 1200
rect 790 1204 796 1205
rect 790 1200 791 1204
rect 795 1200 796 1204
rect 790 1199 796 1200
rect 862 1204 868 1205
rect 862 1200 863 1204
rect 867 1200 868 1204
rect 862 1199 868 1200
rect 1286 1201 1292 1202
rect 110 1196 116 1197
rect 1286 1197 1287 1201
rect 1291 1197 1292 1201
rect 1286 1196 1292 1197
rect 110 1184 116 1185
rect 1286 1184 1292 1185
rect 110 1180 111 1184
rect 115 1180 116 1184
rect 110 1179 116 1180
rect 150 1183 156 1184
rect 150 1179 151 1183
rect 155 1179 156 1183
rect 150 1178 156 1179
rect 206 1183 212 1184
rect 206 1179 207 1183
rect 211 1179 212 1183
rect 206 1178 212 1179
rect 286 1183 292 1184
rect 286 1179 287 1183
rect 291 1179 292 1183
rect 286 1178 292 1179
rect 366 1183 372 1184
rect 366 1179 367 1183
rect 371 1179 372 1183
rect 366 1178 372 1179
rect 446 1183 452 1184
rect 446 1179 447 1183
rect 451 1179 452 1183
rect 446 1178 452 1179
rect 526 1183 532 1184
rect 526 1179 527 1183
rect 531 1179 532 1183
rect 526 1178 532 1179
rect 598 1183 604 1184
rect 598 1179 599 1183
rect 603 1179 604 1183
rect 598 1178 604 1179
rect 662 1183 668 1184
rect 662 1179 663 1183
rect 667 1179 668 1183
rect 662 1178 668 1179
rect 734 1183 740 1184
rect 734 1179 735 1183
rect 739 1179 740 1183
rect 734 1178 740 1179
rect 806 1183 812 1184
rect 806 1179 807 1183
rect 811 1179 812 1183
rect 806 1178 812 1179
rect 878 1183 884 1184
rect 878 1179 879 1183
rect 883 1179 884 1183
rect 1286 1180 1287 1184
rect 1291 1180 1292 1184
rect 1286 1179 1292 1180
rect 878 1178 884 1179
rect 1566 1157 1572 1158
rect 1326 1156 1332 1157
rect 1326 1152 1327 1156
rect 1331 1152 1332 1156
rect 1566 1153 1567 1157
rect 1571 1153 1572 1157
rect 1566 1152 1572 1153
rect 1630 1157 1636 1158
rect 1630 1153 1631 1157
rect 1635 1153 1636 1157
rect 1630 1152 1636 1153
rect 1702 1157 1708 1158
rect 1702 1153 1703 1157
rect 1707 1153 1708 1157
rect 1702 1152 1708 1153
rect 1790 1157 1796 1158
rect 1790 1153 1791 1157
rect 1795 1153 1796 1157
rect 1790 1152 1796 1153
rect 1902 1157 1908 1158
rect 1902 1153 1903 1157
rect 1907 1153 1908 1157
rect 1902 1152 1908 1153
rect 2030 1157 2036 1158
rect 2030 1153 2031 1157
rect 2035 1153 2036 1157
rect 2030 1152 2036 1153
rect 2174 1157 2180 1158
rect 2174 1153 2175 1157
rect 2179 1153 2180 1157
rect 2174 1152 2180 1153
rect 2326 1157 2332 1158
rect 2326 1153 2327 1157
rect 2331 1153 2332 1157
rect 2326 1152 2332 1153
rect 2454 1157 2460 1158
rect 2454 1153 2455 1157
rect 2459 1153 2460 1157
rect 2454 1152 2460 1153
rect 2502 1156 2508 1157
rect 2502 1152 2503 1156
rect 2507 1152 2508 1156
rect 1326 1151 1332 1152
rect 2502 1151 2508 1152
rect 1326 1139 1332 1140
rect 1326 1135 1327 1139
rect 1331 1135 1332 1139
rect 2502 1139 2508 1140
rect 1326 1134 1332 1135
rect 1550 1136 1556 1137
rect 1550 1132 1551 1136
rect 1555 1132 1556 1136
rect 1550 1131 1556 1132
rect 1614 1136 1620 1137
rect 1614 1132 1615 1136
rect 1619 1132 1620 1136
rect 1614 1131 1620 1132
rect 1686 1136 1692 1137
rect 1686 1132 1687 1136
rect 1691 1132 1692 1136
rect 1686 1131 1692 1132
rect 1774 1136 1780 1137
rect 1774 1132 1775 1136
rect 1779 1132 1780 1136
rect 1774 1131 1780 1132
rect 1886 1136 1892 1137
rect 1886 1132 1887 1136
rect 1891 1132 1892 1136
rect 1886 1131 1892 1132
rect 2014 1136 2020 1137
rect 2014 1132 2015 1136
rect 2019 1132 2020 1136
rect 2014 1131 2020 1132
rect 2158 1136 2164 1137
rect 2158 1132 2159 1136
rect 2163 1132 2164 1136
rect 2158 1131 2164 1132
rect 2310 1136 2316 1137
rect 2310 1132 2311 1136
rect 2315 1132 2316 1136
rect 2310 1131 2316 1132
rect 2438 1136 2444 1137
rect 2438 1132 2439 1136
rect 2443 1132 2444 1136
rect 2502 1135 2503 1139
rect 2507 1135 2508 1139
rect 2502 1134 2508 1135
rect 2438 1131 2444 1132
rect 182 1129 188 1130
rect 110 1128 116 1129
rect 110 1124 111 1128
rect 115 1124 116 1128
rect 182 1125 183 1129
rect 187 1125 188 1129
rect 182 1124 188 1125
rect 278 1129 284 1130
rect 278 1125 279 1129
rect 283 1125 284 1129
rect 278 1124 284 1125
rect 374 1129 380 1130
rect 374 1125 375 1129
rect 379 1125 380 1129
rect 374 1124 380 1125
rect 470 1129 476 1130
rect 470 1125 471 1129
rect 475 1125 476 1129
rect 470 1124 476 1125
rect 566 1129 572 1130
rect 566 1125 567 1129
rect 571 1125 572 1129
rect 566 1124 572 1125
rect 654 1129 660 1130
rect 654 1125 655 1129
rect 659 1125 660 1129
rect 654 1124 660 1125
rect 734 1129 740 1130
rect 734 1125 735 1129
rect 739 1125 740 1129
rect 734 1124 740 1125
rect 806 1129 812 1130
rect 806 1125 807 1129
rect 811 1125 812 1129
rect 806 1124 812 1125
rect 878 1129 884 1130
rect 878 1125 879 1129
rect 883 1125 884 1129
rect 878 1124 884 1125
rect 958 1129 964 1130
rect 958 1125 959 1129
rect 963 1125 964 1129
rect 958 1124 964 1125
rect 1038 1129 1044 1130
rect 1038 1125 1039 1129
rect 1043 1125 1044 1129
rect 1038 1124 1044 1125
rect 1286 1128 1292 1129
rect 1286 1124 1287 1128
rect 1291 1124 1292 1128
rect 110 1123 116 1124
rect 1286 1123 1292 1124
rect 1382 1124 1388 1125
rect 1326 1121 1332 1122
rect 1326 1117 1327 1121
rect 1331 1117 1332 1121
rect 1382 1120 1383 1124
rect 1387 1120 1388 1124
rect 1382 1119 1388 1120
rect 1446 1124 1452 1125
rect 1446 1120 1447 1124
rect 1451 1120 1452 1124
rect 1446 1119 1452 1120
rect 1518 1124 1524 1125
rect 1518 1120 1519 1124
rect 1523 1120 1524 1124
rect 1518 1119 1524 1120
rect 1590 1124 1596 1125
rect 1590 1120 1591 1124
rect 1595 1120 1596 1124
rect 1590 1119 1596 1120
rect 1670 1124 1676 1125
rect 1670 1120 1671 1124
rect 1675 1120 1676 1124
rect 1670 1119 1676 1120
rect 1750 1124 1756 1125
rect 1750 1120 1751 1124
rect 1755 1120 1756 1124
rect 1750 1119 1756 1120
rect 1830 1124 1836 1125
rect 1830 1120 1831 1124
rect 1835 1120 1836 1124
rect 1830 1119 1836 1120
rect 1910 1124 1916 1125
rect 1910 1120 1911 1124
rect 1915 1120 1916 1124
rect 1910 1119 1916 1120
rect 1982 1124 1988 1125
rect 1982 1120 1983 1124
rect 1987 1120 1988 1124
rect 1982 1119 1988 1120
rect 2054 1124 2060 1125
rect 2054 1120 2055 1124
rect 2059 1120 2060 1124
rect 2054 1119 2060 1120
rect 2134 1124 2140 1125
rect 2134 1120 2135 1124
rect 2139 1120 2140 1124
rect 2134 1119 2140 1120
rect 2214 1124 2220 1125
rect 2214 1120 2215 1124
rect 2219 1120 2220 1124
rect 2214 1119 2220 1120
rect 2502 1121 2508 1122
rect 1326 1116 1332 1117
rect 2502 1117 2503 1121
rect 2507 1117 2508 1121
rect 2502 1116 2508 1117
rect 110 1111 116 1112
rect 110 1107 111 1111
rect 115 1107 116 1111
rect 1286 1111 1292 1112
rect 110 1106 116 1107
rect 166 1108 172 1109
rect 166 1104 167 1108
rect 171 1104 172 1108
rect 166 1103 172 1104
rect 262 1108 268 1109
rect 262 1104 263 1108
rect 267 1104 268 1108
rect 262 1103 268 1104
rect 358 1108 364 1109
rect 358 1104 359 1108
rect 363 1104 364 1108
rect 358 1103 364 1104
rect 454 1108 460 1109
rect 454 1104 455 1108
rect 459 1104 460 1108
rect 454 1103 460 1104
rect 550 1108 556 1109
rect 550 1104 551 1108
rect 555 1104 556 1108
rect 550 1103 556 1104
rect 638 1108 644 1109
rect 638 1104 639 1108
rect 643 1104 644 1108
rect 638 1103 644 1104
rect 718 1108 724 1109
rect 718 1104 719 1108
rect 723 1104 724 1108
rect 718 1103 724 1104
rect 790 1108 796 1109
rect 790 1104 791 1108
rect 795 1104 796 1108
rect 790 1103 796 1104
rect 862 1108 868 1109
rect 862 1104 863 1108
rect 867 1104 868 1108
rect 862 1103 868 1104
rect 942 1108 948 1109
rect 942 1104 943 1108
rect 947 1104 948 1108
rect 942 1103 948 1104
rect 1022 1108 1028 1109
rect 1022 1104 1023 1108
rect 1027 1104 1028 1108
rect 1286 1107 1287 1111
rect 1291 1107 1292 1111
rect 1286 1106 1292 1107
rect 1022 1103 1028 1104
rect 1326 1104 1332 1105
rect 2502 1104 2508 1105
rect 1326 1100 1327 1104
rect 1331 1100 1332 1104
rect 1326 1099 1332 1100
rect 1398 1103 1404 1104
rect 1398 1099 1399 1103
rect 1403 1099 1404 1103
rect 1398 1098 1404 1099
rect 1462 1103 1468 1104
rect 1462 1099 1463 1103
rect 1467 1099 1468 1103
rect 1462 1098 1468 1099
rect 1534 1103 1540 1104
rect 1534 1099 1535 1103
rect 1539 1099 1540 1103
rect 1534 1098 1540 1099
rect 1606 1103 1612 1104
rect 1606 1099 1607 1103
rect 1611 1099 1612 1103
rect 1606 1098 1612 1099
rect 1686 1103 1692 1104
rect 1686 1099 1687 1103
rect 1691 1099 1692 1103
rect 1686 1098 1692 1099
rect 1766 1103 1772 1104
rect 1766 1099 1767 1103
rect 1771 1099 1772 1103
rect 1766 1098 1772 1099
rect 1846 1103 1852 1104
rect 1846 1099 1847 1103
rect 1851 1099 1852 1103
rect 1846 1098 1852 1099
rect 1926 1103 1932 1104
rect 1926 1099 1927 1103
rect 1931 1099 1932 1103
rect 1926 1098 1932 1099
rect 1998 1103 2004 1104
rect 1998 1099 1999 1103
rect 2003 1099 2004 1103
rect 1998 1098 2004 1099
rect 2070 1103 2076 1104
rect 2070 1099 2071 1103
rect 2075 1099 2076 1103
rect 2070 1098 2076 1099
rect 2150 1103 2156 1104
rect 2150 1099 2151 1103
rect 2155 1099 2156 1103
rect 2150 1098 2156 1099
rect 2230 1103 2236 1104
rect 2230 1099 2231 1103
rect 2235 1099 2236 1103
rect 2502 1100 2503 1104
rect 2507 1100 2508 1104
rect 2502 1099 2508 1100
rect 2230 1098 2236 1099
rect 206 1088 212 1089
rect 110 1085 116 1086
rect 110 1081 111 1085
rect 115 1081 116 1085
rect 206 1084 207 1088
rect 211 1084 212 1088
rect 206 1083 212 1084
rect 278 1088 284 1089
rect 278 1084 279 1088
rect 283 1084 284 1088
rect 278 1083 284 1084
rect 358 1088 364 1089
rect 358 1084 359 1088
rect 363 1084 364 1088
rect 358 1083 364 1084
rect 446 1088 452 1089
rect 446 1084 447 1088
rect 451 1084 452 1088
rect 446 1083 452 1084
rect 542 1088 548 1089
rect 542 1084 543 1088
rect 547 1084 548 1088
rect 542 1083 548 1084
rect 638 1088 644 1089
rect 638 1084 639 1088
rect 643 1084 644 1088
rect 638 1083 644 1084
rect 726 1088 732 1089
rect 726 1084 727 1088
rect 731 1084 732 1088
rect 726 1083 732 1084
rect 814 1088 820 1089
rect 814 1084 815 1088
rect 819 1084 820 1088
rect 814 1083 820 1084
rect 894 1088 900 1089
rect 894 1084 895 1088
rect 899 1084 900 1088
rect 894 1083 900 1084
rect 974 1088 980 1089
rect 974 1084 975 1088
rect 979 1084 980 1088
rect 974 1083 980 1084
rect 1054 1088 1060 1089
rect 1054 1084 1055 1088
rect 1059 1084 1060 1088
rect 1054 1083 1060 1084
rect 1142 1088 1148 1089
rect 1142 1084 1143 1088
rect 1147 1084 1148 1088
rect 1142 1083 1148 1084
rect 1286 1085 1292 1086
rect 110 1080 116 1081
rect 1286 1081 1287 1085
rect 1291 1081 1292 1085
rect 1286 1080 1292 1081
rect 110 1068 116 1069
rect 1286 1068 1292 1069
rect 110 1064 111 1068
rect 115 1064 116 1068
rect 110 1063 116 1064
rect 222 1067 228 1068
rect 222 1063 223 1067
rect 227 1063 228 1067
rect 222 1062 228 1063
rect 294 1067 300 1068
rect 294 1063 295 1067
rect 299 1063 300 1067
rect 294 1062 300 1063
rect 374 1067 380 1068
rect 374 1063 375 1067
rect 379 1063 380 1067
rect 374 1062 380 1063
rect 462 1067 468 1068
rect 462 1063 463 1067
rect 467 1063 468 1067
rect 462 1062 468 1063
rect 558 1067 564 1068
rect 558 1063 559 1067
rect 563 1063 564 1067
rect 558 1062 564 1063
rect 654 1067 660 1068
rect 654 1063 655 1067
rect 659 1063 660 1067
rect 654 1062 660 1063
rect 742 1067 748 1068
rect 742 1063 743 1067
rect 747 1063 748 1067
rect 742 1062 748 1063
rect 830 1067 836 1068
rect 830 1063 831 1067
rect 835 1063 836 1067
rect 830 1062 836 1063
rect 910 1067 916 1068
rect 910 1063 911 1067
rect 915 1063 916 1067
rect 910 1062 916 1063
rect 990 1067 996 1068
rect 990 1063 991 1067
rect 995 1063 996 1067
rect 990 1062 996 1063
rect 1070 1067 1076 1068
rect 1070 1063 1071 1067
rect 1075 1063 1076 1067
rect 1070 1062 1076 1063
rect 1158 1067 1164 1068
rect 1158 1063 1159 1067
rect 1163 1063 1164 1067
rect 1286 1064 1287 1068
rect 1291 1064 1292 1068
rect 1286 1063 1292 1064
rect 1158 1062 1164 1063
rect 1366 1045 1372 1046
rect 1326 1044 1332 1045
rect 1326 1040 1327 1044
rect 1331 1040 1332 1044
rect 1366 1041 1367 1045
rect 1371 1041 1372 1045
rect 1366 1040 1372 1041
rect 1454 1045 1460 1046
rect 1454 1041 1455 1045
rect 1459 1041 1460 1045
rect 1454 1040 1460 1041
rect 1574 1045 1580 1046
rect 1574 1041 1575 1045
rect 1579 1041 1580 1045
rect 1574 1040 1580 1041
rect 1694 1045 1700 1046
rect 1694 1041 1695 1045
rect 1699 1041 1700 1045
rect 1694 1040 1700 1041
rect 1814 1045 1820 1046
rect 1814 1041 1815 1045
rect 1819 1041 1820 1045
rect 1814 1040 1820 1041
rect 1926 1045 1932 1046
rect 1926 1041 1927 1045
rect 1931 1041 1932 1045
rect 1926 1040 1932 1041
rect 2038 1045 2044 1046
rect 2038 1041 2039 1045
rect 2043 1041 2044 1045
rect 2038 1040 2044 1041
rect 2150 1045 2156 1046
rect 2150 1041 2151 1045
rect 2155 1041 2156 1045
rect 2150 1040 2156 1041
rect 2254 1045 2260 1046
rect 2254 1041 2255 1045
rect 2259 1041 2260 1045
rect 2254 1040 2260 1041
rect 2366 1045 2372 1046
rect 2366 1041 2367 1045
rect 2371 1041 2372 1045
rect 2366 1040 2372 1041
rect 2454 1045 2460 1046
rect 2454 1041 2455 1045
rect 2459 1041 2460 1045
rect 2454 1040 2460 1041
rect 2502 1044 2508 1045
rect 2502 1040 2503 1044
rect 2507 1040 2508 1044
rect 1326 1039 1332 1040
rect 2502 1039 2508 1040
rect 1326 1027 1332 1028
rect 1326 1023 1327 1027
rect 1331 1023 1332 1027
rect 2502 1027 2508 1028
rect 1326 1022 1332 1023
rect 1350 1024 1356 1025
rect 1350 1020 1351 1024
rect 1355 1020 1356 1024
rect 1350 1019 1356 1020
rect 1438 1024 1444 1025
rect 1438 1020 1439 1024
rect 1443 1020 1444 1024
rect 1438 1019 1444 1020
rect 1558 1024 1564 1025
rect 1558 1020 1559 1024
rect 1563 1020 1564 1024
rect 1558 1019 1564 1020
rect 1678 1024 1684 1025
rect 1678 1020 1679 1024
rect 1683 1020 1684 1024
rect 1678 1019 1684 1020
rect 1798 1024 1804 1025
rect 1798 1020 1799 1024
rect 1803 1020 1804 1024
rect 1798 1019 1804 1020
rect 1910 1024 1916 1025
rect 1910 1020 1911 1024
rect 1915 1020 1916 1024
rect 1910 1019 1916 1020
rect 2022 1024 2028 1025
rect 2022 1020 2023 1024
rect 2027 1020 2028 1024
rect 2022 1019 2028 1020
rect 2134 1024 2140 1025
rect 2134 1020 2135 1024
rect 2139 1020 2140 1024
rect 2134 1019 2140 1020
rect 2238 1024 2244 1025
rect 2238 1020 2239 1024
rect 2243 1020 2244 1024
rect 2238 1019 2244 1020
rect 2350 1024 2356 1025
rect 2350 1020 2351 1024
rect 2355 1020 2356 1024
rect 2350 1019 2356 1020
rect 2438 1024 2444 1025
rect 2438 1020 2439 1024
rect 2443 1020 2444 1024
rect 2502 1023 2503 1027
rect 2507 1023 2508 1027
rect 2502 1022 2508 1023
rect 2438 1019 2444 1020
rect 294 1009 300 1010
rect 110 1008 116 1009
rect 110 1004 111 1008
rect 115 1004 116 1008
rect 294 1005 295 1009
rect 299 1005 300 1009
rect 294 1004 300 1005
rect 382 1009 388 1010
rect 382 1005 383 1009
rect 387 1005 388 1009
rect 382 1004 388 1005
rect 478 1009 484 1010
rect 478 1005 479 1009
rect 483 1005 484 1009
rect 478 1004 484 1005
rect 574 1009 580 1010
rect 574 1005 575 1009
rect 579 1005 580 1009
rect 574 1004 580 1005
rect 670 1009 676 1010
rect 670 1005 671 1009
rect 675 1005 676 1009
rect 670 1004 676 1005
rect 766 1009 772 1010
rect 766 1005 767 1009
rect 771 1005 772 1009
rect 766 1004 772 1005
rect 854 1009 860 1010
rect 854 1005 855 1009
rect 859 1005 860 1009
rect 854 1004 860 1005
rect 942 1009 948 1010
rect 942 1005 943 1009
rect 947 1005 948 1009
rect 942 1004 948 1005
rect 1022 1009 1028 1010
rect 1022 1005 1023 1009
rect 1027 1005 1028 1009
rect 1022 1004 1028 1005
rect 1102 1009 1108 1010
rect 1102 1005 1103 1009
rect 1107 1005 1108 1009
rect 1102 1004 1108 1005
rect 1182 1009 1188 1010
rect 1182 1005 1183 1009
rect 1187 1005 1188 1009
rect 1182 1004 1188 1005
rect 1238 1009 1244 1010
rect 1238 1005 1239 1009
rect 1243 1005 1244 1009
rect 1238 1004 1244 1005
rect 1286 1008 1292 1009
rect 1286 1004 1287 1008
rect 1291 1004 1292 1008
rect 1350 1008 1356 1009
rect 110 1003 116 1004
rect 1286 1003 1292 1004
rect 1326 1005 1332 1006
rect 1326 1001 1327 1005
rect 1331 1001 1332 1005
rect 1350 1004 1351 1008
rect 1355 1004 1356 1008
rect 1350 1003 1356 1004
rect 1510 1008 1516 1009
rect 1510 1004 1511 1008
rect 1515 1004 1516 1008
rect 1510 1003 1516 1004
rect 1678 1008 1684 1009
rect 1678 1004 1679 1008
rect 1683 1004 1684 1008
rect 1678 1003 1684 1004
rect 1822 1008 1828 1009
rect 1822 1004 1823 1008
rect 1827 1004 1828 1008
rect 1822 1003 1828 1004
rect 1950 1008 1956 1009
rect 1950 1004 1951 1008
rect 1955 1004 1956 1008
rect 1950 1003 1956 1004
rect 2070 1008 2076 1009
rect 2070 1004 2071 1008
rect 2075 1004 2076 1008
rect 2070 1003 2076 1004
rect 2174 1008 2180 1009
rect 2174 1004 2175 1008
rect 2179 1004 2180 1008
rect 2174 1003 2180 1004
rect 2270 1008 2276 1009
rect 2270 1004 2271 1008
rect 2275 1004 2276 1008
rect 2270 1003 2276 1004
rect 2366 1008 2372 1009
rect 2366 1004 2367 1008
rect 2371 1004 2372 1008
rect 2366 1003 2372 1004
rect 2438 1008 2444 1009
rect 2438 1004 2439 1008
rect 2443 1004 2444 1008
rect 2438 1003 2444 1004
rect 2502 1005 2508 1006
rect 1326 1000 1332 1001
rect 2502 1001 2503 1005
rect 2507 1001 2508 1005
rect 2502 1000 2508 1001
rect 110 991 116 992
rect 110 987 111 991
rect 115 987 116 991
rect 1286 991 1292 992
rect 110 986 116 987
rect 278 988 284 989
rect 278 984 279 988
rect 283 984 284 988
rect 278 983 284 984
rect 366 988 372 989
rect 366 984 367 988
rect 371 984 372 988
rect 366 983 372 984
rect 462 988 468 989
rect 462 984 463 988
rect 467 984 468 988
rect 462 983 468 984
rect 558 988 564 989
rect 558 984 559 988
rect 563 984 564 988
rect 558 983 564 984
rect 654 988 660 989
rect 654 984 655 988
rect 659 984 660 988
rect 654 983 660 984
rect 750 988 756 989
rect 750 984 751 988
rect 755 984 756 988
rect 750 983 756 984
rect 838 988 844 989
rect 838 984 839 988
rect 843 984 844 988
rect 838 983 844 984
rect 926 988 932 989
rect 926 984 927 988
rect 931 984 932 988
rect 926 983 932 984
rect 1006 988 1012 989
rect 1006 984 1007 988
rect 1011 984 1012 988
rect 1006 983 1012 984
rect 1086 988 1092 989
rect 1086 984 1087 988
rect 1091 984 1092 988
rect 1086 983 1092 984
rect 1166 988 1172 989
rect 1166 984 1167 988
rect 1171 984 1172 988
rect 1166 983 1172 984
rect 1222 988 1228 989
rect 1222 984 1223 988
rect 1227 984 1228 988
rect 1286 987 1287 991
rect 1291 987 1292 991
rect 1286 986 1292 987
rect 1326 988 1332 989
rect 2502 988 2508 989
rect 1222 983 1228 984
rect 1326 984 1327 988
rect 1331 984 1332 988
rect 1326 983 1332 984
rect 1366 987 1372 988
rect 1366 983 1367 987
rect 1371 983 1372 987
rect 1366 982 1372 983
rect 1526 987 1532 988
rect 1526 983 1527 987
rect 1531 983 1532 987
rect 1526 982 1532 983
rect 1694 987 1700 988
rect 1694 983 1695 987
rect 1699 983 1700 987
rect 1694 982 1700 983
rect 1838 987 1844 988
rect 1838 983 1839 987
rect 1843 983 1844 987
rect 1838 982 1844 983
rect 1966 987 1972 988
rect 1966 983 1967 987
rect 1971 983 1972 987
rect 1966 982 1972 983
rect 2086 987 2092 988
rect 2086 983 2087 987
rect 2091 983 2092 987
rect 2086 982 2092 983
rect 2190 987 2196 988
rect 2190 983 2191 987
rect 2195 983 2196 987
rect 2190 982 2196 983
rect 2286 987 2292 988
rect 2286 983 2287 987
rect 2291 983 2292 987
rect 2286 982 2292 983
rect 2382 987 2388 988
rect 2382 983 2383 987
rect 2387 983 2388 987
rect 2382 982 2388 983
rect 2454 987 2460 988
rect 2454 983 2455 987
rect 2459 983 2460 987
rect 2502 984 2503 988
rect 2507 984 2508 988
rect 2502 983 2508 984
rect 2454 982 2460 983
rect 270 976 276 977
rect 110 973 116 974
rect 110 969 111 973
rect 115 969 116 973
rect 270 972 271 976
rect 275 972 276 976
rect 270 971 276 972
rect 358 976 364 977
rect 358 972 359 976
rect 363 972 364 976
rect 358 971 364 972
rect 454 976 460 977
rect 454 972 455 976
rect 459 972 460 976
rect 454 971 460 972
rect 550 976 556 977
rect 550 972 551 976
rect 555 972 556 976
rect 550 971 556 972
rect 654 976 660 977
rect 654 972 655 976
rect 659 972 660 976
rect 654 971 660 972
rect 750 976 756 977
rect 750 972 751 976
rect 755 972 756 976
rect 750 971 756 972
rect 838 976 844 977
rect 838 972 839 976
rect 843 972 844 976
rect 838 971 844 972
rect 926 976 932 977
rect 926 972 927 976
rect 931 972 932 976
rect 926 971 932 972
rect 1006 976 1012 977
rect 1006 972 1007 976
rect 1011 972 1012 976
rect 1006 971 1012 972
rect 1086 976 1092 977
rect 1086 972 1087 976
rect 1091 972 1092 976
rect 1086 971 1092 972
rect 1166 976 1172 977
rect 1166 972 1167 976
rect 1171 972 1172 976
rect 1166 971 1172 972
rect 1222 976 1228 977
rect 1222 972 1223 976
rect 1227 972 1228 976
rect 1222 971 1228 972
rect 1286 973 1292 974
rect 110 968 116 969
rect 1286 969 1287 973
rect 1291 969 1292 973
rect 1286 968 1292 969
rect 110 956 116 957
rect 1286 956 1292 957
rect 110 952 111 956
rect 115 952 116 956
rect 110 951 116 952
rect 286 955 292 956
rect 286 951 287 955
rect 291 951 292 955
rect 286 950 292 951
rect 374 955 380 956
rect 374 951 375 955
rect 379 951 380 955
rect 374 950 380 951
rect 470 955 476 956
rect 470 951 471 955
rect 475 951 476 955
rect 470 950 476 951
rect 566 955 572 956
rect 566 951 567 955
rect 571 951 572 955
rect 566 950 572 951
rect 670 955 676 956
rect 670 951 671 955
rect 675 951 676 955
rect 670 950 676 951
rect 766 955 772 956
rect 766 951 767 955
rect 771 951 772 955
rect 766 950 772 951
rect 854 955 860 956
rect 854 951 855 955
rect 859 951 860 955
rect 854 950 860 951
rect 942 955 948 956
rect 942 951 943 955
rect 947 951 948 955
rect 942 950 948 951
rect 1022 955 1028 956
rect 1022 951 1023 955
rect 1027 951 1028 955
rect 1022 950 1028 951
rect 1102 955 1108 956
rect 1102 951 1103 955
rect 1107 951 1108 955
rect 1102 950 1108 951
rect 1182 955 1188 956
rect 1182 951 1183 955
rect 1187 951 1188 955
rect 1182 950 1188 951
rect 1238 955 1244 956
rect 1238 951 1239 955
rect 1243 951 1244 955
rect 1286 952 1287 956
rect 1291 952 1292 956
rect 1286 951 1292 952
rect 1238 950 1244 951
rect 1366 925 1372 926
rect 1326 924 1332 925
rect 1326 920 1327 924
rect 1331 920 1332 924
rect 1366 921 1367 925
rect 1371 921 1372 925
rect 1366 920 1372 921
rect 1422 925 1428 926
rect 1422 921 1423 925
rect 1427 921 1428 925
rect 1422 920 1428 921
rect 1502 925 1508 926
rect 1502 921 1503 925
rect 1507 921 1508 925
rect 1502 920 1508 921
rect 1606 925 1612 926
rect 1606 921 1607 925
rect 1611 921 1612 925
rect 1606 920 1612 921
rect 1718 925 1724 926
rect 1718 921 1719 925
rect 1723 921 1724 925
rect 1718 920 1724 921
rect 1830 925 1836 926
rect 1830 921 1831 925
rect 1835 921 1836 925
rect 1830 920 1836 921
rect 1934 925 1940 926
rect 1934 921 1935 925
rect 1939 921 1940 925
rect 1934 920 1940 921
rect 2030 925 2036 926
rect 2030 921 2031 925
rect 2035 921 2036 925
rect 2030 920 2036 921
rect 2126 925 2132 926
rect 2126 921 2127 925
rect 2131 921 2132 925
rect 2126 920 2132 921
rect 2214 925 2220 926
rect 2214 921 2215 925
rect 2219 921 2220 925
rect 2214 920 2220 921
rect 2294 925 2300 926
rect 2294 921 2295 925
rect 2299 921 2300 925
rect 2294 920 2300 921
rect 2374 925 2380 926
rect 2374 921 2375 925
rect 2379 921 2380 925
rect 2374 920 2380 921
rect 2454 925 2460 926
rect 2454 921 2455 925
rect 2459 921 2460 925
rect 2454 920 2460 921
rect 2502 924 2508 925
rect 2502 920 2503 924
rect 2507 920 2508 924
rect 1326 919 1332 920
rect 2502 919 2508 920
rect 1326 907 1332 908
rect 1326 903 1327 907
rect 1331 903 1332 907
rect 2502 907 2508 908
rect 1326 902 1332 903
rect 1350 904 1356 905
rect 1350 900 1351 904
rect 1355 900 1356 904
rect 1350 899 1356 900
rect 1406 904 1412 905
rect 1406 900 1407 904
rect 1411 900 1412 904
rect 1406 899 1412 900
rect 1486 904 1492 905
rect 1486 900 1487 904
rect 1491 900 1492 904
rect 1486 899 1492 900
rect 1590 904 1596 905
rect 1590 900 1591 904
rect 1595 900 1596 904
rect 1590 899 1596 900
rect 1702 904 1708 905
rect 1702 900 1703 904
rect 1707 900 1708 904
rect 1702 899 1708 900
rect 1814 904 1820 905
rect 1814 900 1815 904
rect 1819 900 1820 904
rect 1814 899 1820 900
rect 1918 904 1924 905
rect 1918 900 1919 904
rect 1923 900 1924 904
rect 1918 899 1924 900
rect 2014 904 2020 905
rect 2014 900 2015 904
rect 2019 900 2020 904
rect 2014 899 2020 900
rect 2110 904 2116 905
rect 2110 900 2111 904
rect 2115 900 2116 904
rect 2110 899 2116 900
rect 2198 904 2204 905
rect 2198 900 2199 904
rect 2203 900 2204 904
rect 2198 899 2204 900
rect 2278 904 2284 905
rect 2278 900 2279 904
rect 2283 900 2284 904
rect 2278 899 2284 900
rect 2358 904 2364 905
rect 2358 900 2359 904
rect 2363 900 2364 904
rect 2358 899 2364 900
rect 2438 904 2444 905
rect 2438 900 2439 904
rect 2443 900 2444 904
rect 2502 903 2503 907
rect 2507 903 2508 907
rect 2502 902 2508 903
rect 2438 899 2444 900
rect 270 897 276 898
rect 110 896 116 897
rect 110 892 111 896
rect 115 892 116 896
rect 270 893 271 897
rect 275 893 276 897
rect 270 892 276 893
rect 342 897 348 898
rect 342 893 343 897
rect 347 893 348 897
rect 342 892 348 893
rect 422 897 428 898
rect 422 893 423 897
rect 427 893 428 897
rect 422 892 428 893
rect 518 897 524 898
rect 518 893 519 897
rect 523 893 524 897
rect 518 892 524 893
rect 614 897 620 898
rect 614 893 615 897
rect 619 893 620 897
rect 614 892 620 893
rect 710 897 716 898
rect 710 893 711 897
rect 715 893 716 897
rect 710 892 716 893
rect 806 897 812 898
rect 806 893 807 897
rect 811 893 812 897
rect 806 892 812 893
rect 902 897 908 898
rect 902 893 903 897
rect 907 893 908 897
rect 902 892 908 893
rect 990 897 996 898
rect 990 893 991 897
rect 995 893 996 897
rect 990 892 996 893
rect 1086 897 1092 898
rect 1086 893 1087 897
rect 1091 893 1092 897
rect 1086 892 1092 893
rect 1182 897 1188 898
rect 1182 893 1183 897
rect 1187 893 1188 897
rect 1182 892 1188 893
rect 1286 896 1292 897
rect 1286 892 1287 896
rect 1291 892 1292 896
rect 110 891 116 892
rect 1286 891 1292 892
rect 1430 888 1436 889
rect 1326 885 1332 886
rect 1326 881 1327 885
rect 1331 881 1332 885
rect 1430 884 1431 888
rect 1435 884 1436 888
rect 1430 883 1436 884
rect 1486 888 1492 889
rect 1486 884 1487 888
rect 1491 884 1492 888
rect 1486 883 1492 884
rect 1550 888 1556 889
rect 1550 884 1551 888
rect 1555 884 1556 888
rect 1550 883 1556 884
rect 1622 888 1628 889
rect 1622 884 1623 888
rect 1627 884 1628 888
rect 1622 883 1628 884
rect 1702 888 1708 889
rect 1702 884 1703 888
rect 1707 884 1708 888
rect 1702 883 1708 884
rect 1790 888 1796 889
rect 1790 884 1791 888
rect 1795 884 1796 888
rect 1790 883 1796 884
rect 1894 888 1900 889
rect 1894 884 1895 888
rect 1899 884 1900 888
rect 1894 883 1900 884
rect 2014 888 2020 889
rect 2014 884 2015 888
rect 2019 884 2020 888
rect 2014 883 2020 884
rect 2142 888 2148 889
rect 2142 884 2143 888
rect 2147 884 2148 888
rect 2142 883 2148 884
rect 2278 888 2284 889
rect 2278 884 2279 888
rect 2283 884 2284 888
rect 2278 883 2284 884
rect 2422 888 2428 889
rect 2422 884 2423 888
rect 2427 884 2428 888
rect 2422 883 2428 884
rect 2502 885 2508 886
rect 1326 880 1332 881
rect 2502 881 2503 885
rect 2507 881 2508 885
rect 2502 880 2508 881
rect 110 879 116 880
rect 110 875 111 879
rect 115 875 116 879
rect 1286 879 1292 880
rect 110 874 116 875
rect 254 876 260 877
rect 254 872 255 876
rect 259 872 260 876
rect 254 871 260 872
rect 326 876 332 877
rect 326 872 327 876
rect 331 872 332 876
rect 326 871 332 872
rect 406 876 412 877
rect 406 872 407 876
rect 411 872 412 876
rect 406 871 412 872
rect 502 876 508 877
rect 502 872 503 876
rect 507 872 508 876
rect 502 871 508 872
rect 598 876 604 877
rect 598 872 599 876
rect 603 872 604 876
rect 598 871 604 872
rect 694 876 700 877
rect 694 872 695 876
rect 699 872 700 876
rect 694 871 700 872
rect 790 876 796 877
rect 790 872 791 876
rect 795 872 796 876
rect 790 871 796 872
rect 886 876 892 877
rect 886 872 887 876
rect 891 872 892 876
rect 886 871 892 872
rect 974 876 980 877
rect 974 872 975 876
rect 979 872 980 876
rect 974 871 980 872
rect 1070 876 1076 877
rect 1070 872 1071 876
rect 1075 872 1076 876
rect 1070 871 1076 872
rect 1166 876 1172 877
rect 1166 872 1167 876
rect 1171 872 1172 876
rect 1286 875 1287 879
rect 1291 875 1292 879
rect 1286 874 1292 875
rect 1166 871 1172 872
rect 1326 868 1332 869
rect 2502 868 2508 869
rect 1326 864 1327 868
rect 1331 864 1332 868
rect 1326 863 1332 864
rect 1446 867 1452 868
rect 1446 863 1447 867
rect 1451 863 1452 867
rect 1446 862 1452 863
rect 1502 867 1508 868
rect 1502 863 1503 867
rect 1507 863 1508 867
rect 1502 862 1508 863
rect 1566 867 1572 868
rect 1566 863 1567 867
rect 1571 863 1572 867
rect 1566 862 1572 863
rect 1638 867 1644 868
rect 1638 863 1639 867
rect 1643 863 1644 867
rect 1638 862 1644 863
rect 1718 867 1724 868
rect 1718 863 1719 867
rect 1723 863 1724 867
rect 1718 862 1724 863
rect 1806 867 1812 868
rect 1806 863 1807 867
rect 1811 863 1812 867
rect 1806 862 1812 863
rect 1910 867 1916 868
rect 1910 863 1911 867
rect 1915 863 1916 867
rect 1910 862 1916 863
rect 2030 867 2036 868
rect 2030 863 2031 867
rect 2035 863 2036 867
rect 2030 862 2036 863
rect 2158 867 2164 868
rect 2158 863 2159 867
rect 2163 863 2164 867
rect 2158 862 2164 863
rect 2294 867 2300 868
rect 2294 863 2295 867
rect 2299 863 2300 867
rect 2294 862 2300 863
rect 2438 867 2444 868
rect 2438 863 2439 867
rect 2443 863 2444 867
rect 2502 864 2503 868
rect 2507 864 2508 868
rect 2502 863 2508 864
rect 2438 862 2444 863
rect 246 860 252 861
rect 110 857 116 858
rect 110 853 111 857
rect 115 853 116 857
rect 246 856 247 860
rect 251 856 252 860
rect 246 855 252 856
rect 310 860 316 861
rect 310 856 311 860
rect 315 856 316 860
rect 310 855 316 856
rect 374 860 380 861
rect 374 856 375 860
rect 379 856 380 860
rect 374 855 380 856
rect 438 860 444 861
rect 438 856 439 860
rect 443 856 444 860
rect 438 855 444 856
rect 502 860 508 861
rect 502 856 503 860
rect 507 856 508 860
rect 502 855 508 856
rect 566 860 572 861
rect 566 856 567 860
rect 571 856 572 860
rect 566 855 572 856
rect 630 860 636 861
rect 630 856 631 860
rect 635 856 636 860
rect 630 855 636 856
rect 694 860 700 861
rect 694 856 695 860
rect 699 856 700 860
rect 694 855 700 856
rect 758 860 764 861
rect 758 856 759 860
rect 763 856 764 860
rect 758 855 764 856
rect 830 860 836 861
rect 830 856 831 860
rect 835 856 836 860
rect 830 855 836 856
rect 902 860 908 861
rect 902 856 903 860
rect 907 856 908 860
rect 902 855 908 856
rect 1286 857 1292 858
rect 110 852 116 853
rect 1286 853 1287 857
rect 1291 853 1292 857
rect 1286 852 1292 853
rect 110 840 116 841
rect 1286 840 1292 841
rect 110 836 111 840
rect 115 836 116 840
rect 110 835 116 836
rect 262 839 268 840
rect 262 835 263 839
rect 267 835 268 839
rect 262 834 268 835
rect 326 839 332 840
rect 326 835 327 839
rect 331 835 332 839
rect 326 834 332 835
rect 390 839 396 840
rect 390 835 391 839
rect 395 835 396 839
rect 390 834 396 835
rect 454 839 460 840
rect 454 835 455 839
rect 459 835 460 839
rect 454 834 460 835
rect 518 839 524 840
rect 518 835 519 839
rect 523 835 524 839
rect 518 834 524 835
rect 582 839 588 840
rect 582 835 583 839
rect 587 835 588 839
rect 582 834 588 835
rect 646 839 652 840
rect 646 835 647 839
rect 651 835 652 839
rect 646 834 652 835
rect 710 839 716 840
rect 710 835 711 839
rect 715 835 716 839
rect 710 834 716 835
rect 774 839 780 840
rect 774 835 775 839
rect 779 835 780 839
rect 774 834 780 835
rect 846 839 852 840
rect 846 835 847 839
rect 851 835 852 839
rect 846 834 852 835
rect 918 839 924 840
rect 918 835 919 839
rect 923 835 924 839
rect 1286 836 1287 840
rect 1291 836 1292 840
rect 1286 835 1292 836
rect 918 834 924 835
rect 1590 813 1596 814
rect 1326 812 1332 813
rect 1326 808 1327 812
rect 1331 808 1332 812
rect 1590 809 1591 813
rect 1595 809 1596 813
rect 1590 808 1596 809
rect 1646 813 1652 814
rect 1646 809 1647 813
rect 1651 809 1652 813
rect 1646 808 1652 809
rect 1702 813 1708 814
rect 1702 809 1703 813
rect 1707 809 1708 813
rect 1702 808 1708 809
rect 1766 813 1772 814
rect 1766 809 1767 813
rect 1771 809 1772 813
rect 1766 808 1772 809
rect 1846 813 1852 814
rect 1846 809 1847 813
rect 1851 809 1852 813
rect 1846 808 1852 809
rect 1926 813 1932 814
rect 1926 809 1927 813
rect 1931 809 1932 813
rect 1926 808 1932 809
rect 2014 813 2020 814
rect 2014 809 2015 813
rect 2019 809 2020 813
rect 2014 808 2020 809
rect 2102 813 2108 814
rect 2102 809 2103 813
rect 2107 809 2108 813
rect 2102 808 2108 809
rect 2190 813 2196 814
rect 2190 809 2191 813
rect 2195 809 2196 813
rect 2190 808 2196 809
rect 2286 813 2292 814
rect 2286 809 2287 813
rect 2291 809 2292 813
rect 2286 808 2292 809
rect 2382 813 2388 814
rect 2382 809 2383 813
rect 2387 809 2388 813
rect 2382 808 2388 809
rect 2454 813 2460 814
rect 2454 809 2455 813
rect 2459 809 2460 813
rect 2454 808 2460 809
rect 2502 812 2508 813
rect 2502 808 2503 812
rect 2507 808 2508 812
rect 1326 807 1332 808
rect 2502 807 2508 808
rect 1326 795 1332 796
rect 1326 791 1327 795
rect 1331 791 1332 795
rect 2502 795 2508 796
rect 1326 790 1332 791
rect 1574 792 1580 793
rect 1574 788 1575 792
rect 1579 788 1580 792
rect 1574 787 1580 788
rect 1630 792 1636 793
rect 1630 788 1631 792
rect 1635 788 1636 792
rect 1630 787 1636 788
rect 1686 792 1692 793
rect 1686 788 1687 792
rect 1691 788 1692 792
rect 1686 787 1692 788
rect 1750 792 1756 793
rect 1750 788 1751 792
rect 1755 788 1756 792
rect 1750 787 1756 788
rect 1830 792 1836 793
rect 1830 788 1831 792
rect 1835 788 1836 792
rect 1830 787 1836 788
rect 1910 792 1916 793
rect 1910 788 1911 792
rect 1915 788 1916 792
rect 1910 787 1916 788
rect 1998 792 2004 793
rect 1998 788 1999 792
rect 2003 788 2004 792
rect 1998 787 2004 788
rect 2086 792 2092 793
rect 2086 788 2087 792
rect 2091 788 2092 792
rect 2086 787 2092 788
rect 2174 792 2180 793
rect 2174 788 2175 792
rect 2179 788 2180 792
rect 2174 787 2180 788
rect 2270 792 2276 793
rect 2270 788 2271 792
rect 2275 788 2276 792
rect 2270 787 2276 788
rect 2366 792 2372 793
rect 2366 788 2367 792
rect 2371 788 2372 792
rect 2366 787 2372 788
rect 2438 792 2444 793
rect 2438 788 2439 792
rect 2443 788 2444 792
rect 2502 791 2503 795
rect 2507 791 2508 795
rect 2502 790 2508 791
rect 2438 787 2444 788
rect 214 785 220 786
rect 110 784 116 785
rect 110 780 111 784
rect 115 780 116 784
rect 214 781 215 785
rect 219 781 220 785
rect 214 780 220 781
rect 302 785 308 786
rect 302 781 303 785
rect 307 781 308 785
rect 302 780 308 781
rect 390 785 396 786
rect 390 781 391 785
rect 395 781 396 785
rect 390 780 396 781
rect 478 785 484 786
rect 478 781 479 785
rect 483 781 484 785
rect 478 780 484 781
rect 558 785 564 786
rect 558 781 559 785
rect 563 781 564 785
rect 558 780 564 781
rect 630 785 636 786
rect 630 781 631 785
rect 635 781 636 785
rect 630 780 636 781
rect 702 785 708 786
rect 702 781 703 785
rect 707 781 708 785
rect 702 780 708 781
rect 766 785 772 786
rect 766 781 767 785
rect 771 781 772 785
rect 766 780 772 781
rect 830 785 836 786
rect 830 781 831 785
rect 835 781 836 785
rect 830 780 836 781
rect 894 785 900 786
rect 894 781 895 785
rect 899 781 900 785
rect 894 780 900 781
rect 966 785 972 786
rect 966 781 967 785
rect 971 781 972 785
rect 966 780 972 781
rect 1038 785 1044 786
rect 1038 781 1039 785
rect 1043 781 1044 785
rect 1038 780 1044 781
rect 1286 784 1292 785
rect 1286 780 1287 784
rect 1291 780 1292 784
rect 110 779 116 780
rect 1286 779 1292 780
rect 1566 776 1572 777
rect 1326 773 1332 774
rect 1326 769 1327 773
rect 1331 769 1332 773
rect 1566 772 1567 776
rect 1571 772 1572 776
rect 1566 771 1572 772
rect 1622 776 1628 777
rect 1622 772 1623 776
rect 1627 772 1628 776
rect 1622 771 1628 772
rect 1686 776 1692 777
rect 1686 772 1687 776
rect 1691 772 1692 776
rect 1686 771 1692 772
rect 1758 776 1764 777
rect 1758 772 1759 776
rect 1763 772 1764 776
rect 1758 771 1764 772
rect 1830 776 1836 777
rect 1830 772 1831 776
rect 1835 772 1836 776
rect 1830 771 1836 772
rect 1918 776 1924 777
rect 1918 772 1919 776
rect 1923 772 1924 776
rect 1918 771 1924 772
rect 2014 776 2020 777
rect 2014 772 2015 776
rect 2019 772 2020 776
rect 2014 771 2020 772
rect 2118 776 2124 777
rect 2118 772 2119 776
rect 2123 772 2124 776
rect 2118 771 2124 772
rect 2230 776 2236 777
rect 2230 772 2231 776
rect 2235 772 2236 776
rect 2230 771 2236 772
rect 2342 776 2348 777
rect 2342 772 2343 776
rect 2347 772 2348 776
rect 2342 771 2348 772
rect 2438 776 2444 777
rect 2438 772 2439 776
rect 2443 772 2444 776
rect 2438 771 2444 772
rect 2502 773 2508 774
rect 1326 768 1332 769
rect 2502 769 2503 773
rect 2507 769 2508 773
rect 2502 768 2508 769
rect 110 767 116 768
rect 110 763 111 767
rect 115 763 116 767
rect 1286 767 1292 768
rect 110 762 116 763
rect 198 764 204 765
rect 198 760 199 764
rect 203 760 204 764
rect 198 759 204 760
rect 286 764 292 765
rect 286 760 287 764
rect 291 760 292 764
rect 286 759 292 760
rect 374 764 380 765
rect 374 760 375 764
rect 379 760 380 764
rect 374 759 380 760
rect 462 764 468 765
rect 462 760 463 764
rect 467 760 468 764
rect 462 759 468 760
rect 542 764 548 765
rect 542 760 543 764
rect 547 760 548 764
rect 542 759 548 760
rect 614 764 620 765
rect 614 760 615 764
rect 619 760 620 764
rect 614 759 620 760
rect 686 764 692 765
rect 686 760 687 764
rect 691 760 692 764
rect 686 759 692 760
rect 750 764 756 765
rect 750 760 751 764
rect 755 760 756 764
rect 750 759 756 760
rect 814 764 820 765
rect 814 760 815 764
rect 819 760 820 764
rect 814 759 820 760
rect 878 764 884 765
rect 878 760 879 764
rect 883 760 884 764
rect 878 759 884 760
rect 950 764 956 765
rect 950 760 951 764
rect 955 760 956 764
rect 950 759 956 760
rect 1022 764 1028 765
rect 1022 760 1023 764
rect 1027 760 1028 764
rect 1286 763 1287 767
rect 1291 763 1292 767
rect 1286 762 1292 763
rect 1022 759 1028 760
rect 1326 756 1332 757
rect 2502 756 2508 757
rect 134 752 140 753
rect 110 749 116 750
rect 110 745 111 749
rect 115 745 116 749
rect 134 748 135 752
rect 139 748 140 752
rect 134 747 140 748
rect 254 752 260 753
rect 254 748 255 752
rect 259 748 260 752
rect 254 747 260 748
rect 390 752 396 753
rect 390 748 391 752
rect 395 748 396 752
rect 390 747 396 748
rect 518 752 524 753
rect 518 748 519 752
rect 523 748 524 752
rect 518 747 524 748
rect 646 752 652 753
rect 646 748 647 752
rect 651 748 652 752
rect 646 747 652 748
rect 774 752 780 753
rect 774 748 775 752
rect 779 748 780 752
rect 774 747 780 748
rect 902 752 908 753
rect 902 748 903 752
rect 907 748 908 752
rect 902 747 908 748
rect 1038 752 1044 753
rect 1038 748 1039 752
rect 1043 748 1044 752
rect 1326 752 1327 756
rect 1331 752 1332 756
rect 1326 751 1332 752
rect 1582 755 1588 756
rect 1582 751 1583 755
rect 1587 751 1588 755
rect 1582 750 1588 751
rect 1638 755 1644 756
rect 1638 751 1639 755
rect 1643 751 1644 755
rect 1638 750 1644 751
rect 1702 755 1708 756
rect 1702 751 1703 755
rect 1707 751 1708 755
rect 1702 750 1708 751
rect 1774 755 1780 756
rect 1774 751 1775 755
rect 1779 751 1780 755
rect 1774 750 1780 751
rect 1846 755 1852 756
rect 1846 751 1847 755
rect 1851 751 1852 755
rect 1846 750 1852 751
rect 1934 755 1940 756
rect 1934 751 1935 755
rect 1939 751 1940 755
rect 1934 750 1940 751
rect 2030 755 2036 756
rect 2030 751 2031 755
rect 2035 751 2036 755
rect 2030 750 2036 751
rect 2134 755 2140 756
rect 2134 751 2135 755
rect 2139 751 2140 755
rect 2134 750 2140 751
rect 2246 755 2252 756
rect 2246 751 2247 755
rect 2251 751 2252 755
rect 2246 750 2252 751
rect 2358 755 2364 756
rect 2358 751 2359 755
rect 2363 751 2364 755
rect 2358 750 2364 751
rect 2454 755 2460 756
rect 2454 751 2455 755
rect 2459 751 2460 755
rect 2502 752 2503 756
rect 2507 752 2508 756
rect 2502 751 2508 752
rect 2454 750 2460 751
rect 1038 747 1044 748
rect 1286 749 1292 750
rect 110 744 116 745
rect 1286 745 1287 749
rect 1291 745 1292 749
rect 1286 744 1292 745
rect 110 732 116 733
rect 1286 732 1292 733
rect 110 728 111 732
rect 115 728 116 732
rect 110 727 116 728
rect 150 731 156 732
rect 150 727 151 731
rect 155 727 156 731
rect 150 726 156 727
rect 270 731 276 732
rect 270 727 271 731
rect 275 727 276 731
rect 270 726 276 727
rect 406 731 412 732
rect 406 727 407 731
rect 411 727 412 731
rect 406 726 412 727
rect 534 731 540 732
rect 534 727 535 731
rect 539 727 540 731
rect 534 726 540 727
rect 662 731 668 732
rect 662 727 663 731
rect 667 727 668 731
rect 662 726 668 727
rect 790 731 796 732
rect 790 727 791 731
rect 795 727 796 731
rect 790 726 796 727
rect 918 731 924 732
rect 918 727 919 731
rect 923 727 924 731
rect 918 726 924 727
rect 1054 731 1060 732
rect 1054 727 1055 731
rect 1059 727 1060 731
rect 1286 728 1287 732
rect 1291 728 1292 732
rect 1286 727 1292 728
rect 1054 726 1060 727
rect 1366 705 1372 706
rect 1326 704 1332 705
rect 1326 700 1327 704
rect 1331 700 1332 704
rect 1366 701 1367 705
rect 1371 701 1372 705
rect 1366 700 1372 701
rect 1430 705 1436 706
rect 1430 701 1431 705
rect 1435 701 1436 705
rect 1430 700 1436 701
rect 1526 705 1532 706
rect 1526 701 1527 705
rect 1531 701 1532 705
rect 1526 700 1532 701
rect 1630 705 1636 706
rect 1630 701 1631 705
rect 1635 701 1636 705
rect 1630 700 1636 701
rect 1734 705 1740 706
rect 1734 701 1735 705
rect 1739 701 1740 705
rect 1734 700 1740 701
rect 1838 705 1844 706
rect 1838 701 1839 705
rect 1843 701 1844 705
rect 1838 700 1844 701
rect 1942 705 1948 706
rect 1942 701 1943 705
rect 1947 701 1948 705
rect 1942 700 1948 701
rect 2046 705 2052 706
rect 2046 701 2047 705
rect 2051 701 2052 705
rect 2046 700 2052 701
rect 2150 705 2156 706
rect 2150 701 2151 705
rect 2155 701 2156 705
rect 2150 700 2156 701
rect 2254 705 2260 706
rect 2254 701 2255 705
rect 2259 701 2260 705
rect 2254 700 2260 701
rect 2366 705 2372 706
rect 2366 701 2367 705
rect 2371 701 2372 705
rect 2366 700 2372 701
rect 2454 705 2460 706
rect 2454 701 2455 705
rect 2459 701 2460 705
rect 2454 700 2460 701
rect 2502 704 2508 705
rect 2502 700 2503 704
rect 2507 700 2508 704
rect 1326 699 1332 700
rect 2502 699 2508 700
rect 1326 687 1332 688
rect 1326 683 1327 687
rect 1331 683 1332 687
rect 2502 687 2508 688
rect 1326 682 1332 683
rect 1350 684 1356 685
rect 150 681 156 682
rect 110 680 116 681
rect 110 676 111 680
rect 115 676 116 680
rect 150 677 151 681
rect 155 677 156 681
rect 150 676 156 677
rect 206 681 212 682
rect 206 677 207 681
rect 211 677 212 681
rect 206 676 212 677
rect 294 681 300 682
rect 294 677 295 681
rect 299 677 300 681
rect 294 676 300 677
rect 390 681 396 682
rect 390 677 391 681
rect 395 677 396 681
rect 390 676 396 677
rect 502 681 508 682
rect 502 677 503 681
rect 507 677 508 681
rect 502 676 508 677
rect 622 681 628 682
rect 622 677 623 681
rect 627 677 628 681
rect 622 676 628 677
rect 742 681 748 682
rect 742 677 743 681
rect 747 677 748 681
rect 742 676 748 677
rect 870 681 876 682
rect 870 677 871 681
rect 875 677 876 681
rect 870 676 876 677
rect 998 681 1004 682
rect 998 677 999 681
rect 1003 677 1004 681
rect 998 676 1004 677
rect 1126 681 1132 682
rect 1126 677 1127 681
rect 1131 677 1132 681
rect 1126 676 1132 677
rect 1238 681 1244 682
rect 1238 677 1239 681
rect 1243 677 1244 681
rect 1238 676 1244 677
rect 1286 680 1292 681
rect 1286 676 1287 680
rect 1291 676 1292 680
rect 1350 680 1351 684
rect 1355 680 1356 684
rect 1350 679 1356 680
rect 1414 684 1420 685
rect 1414 680 1415 684
rect 1419 680 1420 684
rect 1414 679 1420 680
rect 1510 684 1516 685
rect 1510 680 1511 684
rect 1515 680 1516 684
rect 1510 679 1516 680
rect 1614 684 1620 685
rect 1614 680 1615 684
rect 1619 680 1620 684
rect 1614 679 1620 680
rect 1718 684 1724 685
rect 1718 680 1719 684
rect 1723 680 1724 684
rect 1718 679 1724 680
rect 1822 684 1828 685
rect 1822 680 1823 684
rect 1827 680 1828 684
rect 1822 679 1828 680
rect 1926 684 1932 685
rect 1926 680 1927 684
rect 1931 680 1932 684
rect 1926 679 1932 680
rect 2030 684 2036 685
rect 2030 680 2031 684
rect 2035 680 2036 684
rect 2030 679 2036 680
rect 2134 684 2140 685
rect 2134 680 2135 684
rect 2139 680 2140 684
rect 2134 679 2140 680
rect 2238 684 2244 685
rect 2238 680 2239 684
rect 2243 680 2244 684
rect 2238 679 2244 680
rect 2350 684 2356 685
rect 2350 680 2351 684
rect 2355 680 2356 684
rect 2350 679 2356 680
rect 2438 684 2444 685
rect 2438 680 2439 684
rect 2443 680 2444 684
rect 2502 683 2503 687
rect 2507 683 2508 687
rect 2502 682 2508 683
rect 2438 679 2444 680
rect 110 675 116 676
rect 1286 675 1292 676
rect 110 663 116 664
rect 110 659 111 663
rect 115 659 116 663
rect 1286 663 1292 664
rect 110 658 116 659
rect 134 660 140 661
rect 134 656 135 660
rect 139 656 140 660
rect 134 655 140 656
rect 190 660 196 661
rect 190 656 191 660
rect 195 656 196 660
rect 190 655 196 656
rect 278 660 284 661
rect 278 656 279 660
rect 283 656 284 660
rect 278 655 284 656
rect 374 660 380 661
rect 374 656 375 660
rect 379 656 380 660
rect 374 655 380 656
rect 486 660 492 661
rect 486 656 487 660
rect 491 656 492 660
rect 486 655 492 656
rect 606 660 612 661
rect 606 656 607 660
rect 611 656 612 660
rect 606 655 612 656
rect 726 660 732 661
rect 726 656 727 660
rect 731 656 732 660
rect 726 655 732 656
rect 854 660 860 661
rect 854 656 855 660
rect 859 656 860 660
rect 854 655 860 656
rect 982 660 988 661
rect 982 656 983 660
rect 987 656 988 660
rect 982 655 988 656
rect 1110 660 1116 661
rect 1110 656 1111 660
rect 1115 656 1116 660
rect 1110 655 1116 656
rect 1222 660 1228 661
rect 1222 656 1223 660
rect 1227 656 1228 660
rect 1286 659 1287 663
rect 1291 659 1292 663
rect 1286 658 1292 659
rect 1350 660 1356 661
rect 1222 655 1228 656
rect 1326 657 1332 658
rect 1326 653 1327 657
rect 1331 653 1332 657
rect 1350 656 1351 660
rect 1355 656 1356 660
rect 1350 655 1356 656
rect 1414 660 1420 661
rect 1414 656 1415 660
rect 1419 656 1420 660
rect 1414 655 1420 656
rect 1510 660 1516 661
rect 1510 656 1511 660
rect 1515 656 1516 660
rect 1510 655 1516 656
rect 1606 660 1612 661
rect 1606 656 1607 660
rect 1611 656 1612 660
rect 1606 655 1612 656
rect 1710 660 1716 661
rect 1710 656 1711 660
rect 1715 656 1716 660
rect 1710 655 1716 656
rect 1822 660 1828 661
rect 1822 656 1823 660
rect 1827 656 1828 660
rect 1822 655 1828 656
rect 1934 660 1940 661
rect 1934 656 1935 660
rect 1939 656 1940 660
rect 1934 655 1940 656
rect 2054 660 2060 661
rect 2054 656 2055 660
rect 2059 656 2060 660
rect 2054 655 2060 656
rect 2182 660 2188 661
rect 2182 656 2183 660
rect 2187 656 2188 660
rect 2182 655 2188 656
rect 2318 660 2324 661
rect 2318 656 2319 660
rect 2323 656 2324 660
rect 2318 655 2324 656
rect 2438 660 2444 661
rect 2438 656 2439 660
rect 2443 656 2444 660
rect 2438 655 2444 656
rect 2502 657 2508 658
rect 1326 652 1332 653
rect 2502 653 2503 657
rect 2507 653 2508 657
rect 2502 652 2508 653
rect 150 644 156 645
rect 110 641 116 642
rect 110 637 111 641
rect 115 637 116 641
rect 150 640 151 644
rect 155 640 156 644
rect 150 639 156 640
rect 262 644 268 645
rect 262 640 263 644
rect 267 640 268 644
rect 262 639 268 640
rect 366 644 372 645
rect 366 640 367 644
rect 371 640 372 644
rect 366 639 372 640
rect 462 644 468 645
rect 462 640 463 644
rect 467 640 468 644
rect 462 639 468 640
rect 558 644 564 645
rect 558 640 559 644
rect 563 640 564 644
rect 558 639 564 640
rect 654 644 660 645
rect 654 640 655 644
rect 659 640 660 644
rect 654 639 660 640
rect 750 644 756 645
rect 750 640 751 644
rect 755 640 756 644
rect 750 639 756 640
rect 846 644 852 645
rect 846 640 847 644
rect 851 640 852 644
rect 846 639 852 640
rect 942 644 948 645
rect 942 640 943 644
rect 947 640 948 644
rect 942 639 948 640
rect 1038 644 1044 645
rect 1038 640 1039 644
rect 1043 640 1044 644
rect 1038 639 1044 640
rect 1142 644 1148 645
rect 1142 640 1143 644
rect 1147 640 1148 644
rect 1142 639 1148 640
rect 1222 644 1228 645
rect 1222 640 1223 644
rect 1227 640 1228 644
rect 1222 639 1228 640
rect 1286 641 1292 642
rect 110 636 116 637
rect 1286 637 1287 641
rect 1291 637 1292 641
rect 1286 636 1292 637
rect 1326 640 1332 641
rect 2502 640 2508 641
rect 1326 636 1327 640
rect 1331 636 1332 640
rect 1326 635 1332 636
rect 1366 639 1372 640
rect 1366 635 1367 639
rect 1371 635 1372 639
rect 1366 634 1372 635
rect 1430 639 1436 640
rect 1430 635 1431 639
rect 1435 635 1436 639
rect 1430 634 1436 635
rect 1526 639 1532 640
rect 1526 635 1527 639
rect 1531 635 1532 639
rect 1526 634 1532 635
rect 1622 639 1628 640
rect 1622 635 1623 639
rect 1627 635 1628 639
rect 1622 634 1628 635
rect 1726 639 1732 640
rect 1726 635 1727 639
rect 1731 635 1732 639
rect 1726 634 1732 635
rect 1838 639 1844 640
rect 1838 635 1839 639
rect 1843 635 1844 639
rect 1838 634 1844 635
rect 1950 639 1956 640
rect 1950 635 1951 639
rect 1955 635 1956 639
rect 1950 634 1956 635
rect 2070 639 2076 640
rect 2070 635 2071 639
rect 2075 635 2076 639
rect 2070 634 2076 635
rect 2198 639 2204 640
rect 2198 635 2199 639
rect 2203 635 2204 639
rect 2198 634 2204 635
rect 2334 639 2340 640
rect 2334 635 2335 639
rect 2339 635 2340 639
rect 2334 634 2340 635
rect 2454 639 2460 640
rect 2454 635 2455 639
rect 2459 635 2460 639
rect 2502 636 2503 640
rect 2507 636 2508 640
rect 2502 635 2508 636
rect 2454 634 2460 635
rect 110 624 116 625
rect 1286 624 1292 625
rect 110 620 111 624
rect 115 620 116 624
rect 110 619 116 620
rect 166 623 172 624
rect 166 619 167 623
rect 171 619 172 623
rect 166 618 172 619
rect 278 623 284 624
rect 278 619 279 623
rect 283 619 284 623
rect 278 618 284 619
rect 382 623 388 624
rect 382 619 383 623
rect 387 619 388 623
rect 382 618 388 619
rect 478 623 484 624
rect 478 619 479 623
rect 483 619 484 623
rect 478 618 484 619
rect 574 623 580 624
rect 574 619 575 623
rect 579 619 580 623
rect 574 618 580 619
rect 670 623 676 624
rect 670 619 671 623
rect 675 619 676 623
rect 670 618 676 619
rect 766 623 772 624
rect 766 619 767 623
rect 771 619 772 623
rect 766 618 772 619
rect 862 623 868 624
rect 862 619 863 623
rect 867 619 868 623
rect 862 618 868 619
rect 958 623 964 624
rect 958 619 959 623
rect 963 619 964 623
rect 958 618 964 619
rect 1054 623 1060 624
rect 1054 619 1055 623
rect 1059 619 1060 623
rect 1054 618 1060 619
rect 1158 623 1164 624
rect 1158 619 1159 623
rect 1163 619 1164 623
rect 1158 618 1164 619
rect 1238 623 1244 624
rect 1238 619 1239 623
rect 1243 619 1244 623
rect 1286 620 1287 624
rect 1291 620 1292 624
rect 1286 619 1292 620
rect 1238 618 1244 619
rect 1382 589 1388 590
rect 1326 588 1332 589
rect 1326 584 1327 588
rect 1331 584 1332 588
rect 1382 585 1383 589
rect 1387 585 1388 589
rect 1382 584 1388 585
rect 1462 589 1468 590
rect 1462 585 1463 589
rect 1467 585 1468 589
rect 1462 584 1468 585
rect 1550 589 1556 590
rect 1550 585 1551 589
rect 1555 585 1556 589
rect 1550 584 1556 585
rect 1646 589 1652 590
rect 1646 585 1647 589
rect 1651 585 1652 589
rect 1646 584 1652 585
rect 1742 589 1748 590
rect 1742 585 1743 589
rect 1747 585 1748 589
rect 1742 584 1748 585
rect 1846 589 1852 590
rect 1846 585 1847 589
rect 1851 585 1852 589
rect 1846 584 1852 585
rect 1958 589 1964 590
rect 1958 585 1959 589
rect 1963 585 1964 589
rect 1958 584 1964 585
rect 2078 589 2084 590
rect 2078 585 2079 589
rect 2083 585 2084 589
rect 2078 584 2084 585
rect 2206 589 2212 590
rect 2206 585 2207 589
rect 2211 585 2212 589
rect 2206 584 2212 585
rect 2342 589 2348 590
rect 2342 585 2343 589
rect 2347 585 2348 589
rect 2342 584 2348 585
rect 2454 589 2460 590
rect 2454 585 2455 589
rect 2459 585 2460 589
rect 2454 584 2460 585
rect 2502 588 2508 589
rect 2502 584 2503 588
rect 2507 584 2508 588
rect 1326 583 1332 584
rect 2502 583 2508 584
rect 150 573 156 574
rect 110 572 116 573
rect 110 568 111 572
rect 115 568 116 572
rect 150 569 151 573
rect 155 569 156 573
rect 150 568 156 569
rect 238 573 244 574
rect 238 569 239 573
rect 243 569 244 573
rect 238 568 244 569
rect 334 573 340 574
rect 334 569 335 573
rect 339 569 340 573
rect 334 568 340 569
rect 430 573 436 574
rect 430 569 431 573
rect 435 569 436 573
rect 430 568 436 569
rect 534 573 540 574
rect 534 569 535 573
rect 539 569 540 573
rect 534 568 540 569
rect 630 573 636 574
rect 630 569 631 573
rect 635 569 636 573
rect 630 568 636 569
rect 726 573 732 574
rect 726 569 727 573
rect 731 569 732 573
rect 726 568 732 569
rect 822 573 828 574
rect 822 569 823 573
rect 827 569 828 573
rect 822 568 828 569
rect 910 573 916 574
rect 910 569 911 573
rect 915 569 916 573
rect 910 568 916 569
rect 998 573 1004 574
rect 998 569 999 573
rect 1003 569 1004 573
rect 998 568 1004 569
rect 1086 573 1092 574
rect 1086 569 1087 573
rect 1091 569 1092 573
rect 1086 568 1092 569
rect 1182 573 1188 574
rect 1182 569 1183 573
rect 1187 569 1188 573
rect 1182 568 1188 569
rect 1286 572 1292 573
rect 1286 568 1287 572
rect 1291 568 1292 572
rect 110 567 116 568
rect 1286 567 1292 568
rect 1326 571 1332 572
rect 1326 567 1327 571
rect 1331 567 1332 571
rect 2502 571 2508 572
rect 1326 566 1332 567
rect 1366 568 1372 569
rect 1366 564 1367 568
rect 1371 564 1372 568
rect 1366 563 1372 564
rect 1446 568 1452 569
rect 1446 564 1447 568
rect 1451 564 1452 568
rect 1446 563 1452 564
rect 1534 568 1540 569
rect 1534 564 1535 568
rect 1539 564 1540 568
rect 1534 563 1540 564
rect 1630 568 1636 569
rect 1630 564 1631 568
rect 1635 564 1636 568
rect 1630 563 1636 564
rect 1726 568 1732 569
rect 1726 564 1727 568
rect 1731 564 1732 568
rect 1726 563 1732 564
rect 1830 568 1836 569
rect 1830 564 1831 568
rect 1835 564 1836 568
rect 1830 563 1836 564
rect 1942 568 1948 569
rect 1942 564 1943 568
rect 1947 564 1948 568
rect 1942 563 1948 564
rect 2062 568 2068 569
rect 2062 564 2063 568
rect 2067 564 2068 568
rect 2062 563 2068 564
rect 2190 568 2196 569
rect 2190 564 2191 568
rect 2195 564 2196 568
rect 2190 563 2196 564
rect 2326 568 2332 569
rect 2326 564 2327 568
rect 2331 564 2332 568
rect 2326 563 2332 564
rect 2438 568 2444 569
rect 2438 564 2439 568
rect 2443 564 2444 568
rect 2502 567 2503 571
rect 2507 567 2508 571
rect 2502 566 2508 567
rect 2438 563 2444 564
rect 1374 556 1380 557
rect 110 555 116 556
rect 110 551 111 555
rect 115 551 116 555
rect 1286 555 1292 556
rect 110 550 116 551
rect 134 552 140 553
rect 134 548 135 552
rect 139 548 140 552
rect 134 547 140 548
rect 222 552 228 553
rect 222 548 223 552
rect 227 548 228 552
rect 222 547 228 548
rect 318 552 324 553
rect 318 548 319 552
rect 323 548 324 552
rect 318 547 324 548
rect 414 552 420 553
rect 414 548 415 552
rect 419 548 420 552
rect 414 547 420 548
rect 518 552 524 553
rect 518 548 519 552
rect 523 548 524 552
rect 518 547 524 548
rect 614 552 620 553
rect 614 548 615 552
rect 619 548 620 552
rect 614 547 620 548
rect 710 552 716 553
rect 710 548 711 552
rect 715 548 716 552
rect 710 547 716 548
rect 806 552 812 553
rect 806 548 807 552
rect 811 548 812 552
rect 806 547 812 548
rect 894 552 900 553
rect 894 548 895 552
rect 899 548 900 552
rect 894 547 900 548
rect 982 552 988 553
rect 982 548 983 552
rect 987 548 988 552
rect 982 547 988 548
rect 1070 552 1076 553
rect 1070 548 1071 552
rect 1075 548 1076 552
rect 1070 547 1076 548
rect 1166 552 1172 553
rect 1166 548 1167 552
rect 1171 548 1172 552
rect 1286 551 1287 555
rect 1291 551 1292 555
rect 1286 550 1292 551
rect 1326 553 1332 554
rect 1326 549 1327 553
rect 1331 549 1332 553
rect 1374 552 1375 556
rect 1379 552 1380 556
rect 1374 551 1380 552
rect 1454 556 1460 557
rect 1454 552 1455 556
rect 1459 552 1460 556
rect 1454 551 1460 552
rect 1550 556 1556 557
rect 1550 552 1551 556
rect 1555 552 1556 556
rect 1550 551 1556 552
rect 1646 556 1652 557
rect 1646 552 1647 556
rect 1651 552 1652 556
rect 1646 551 1652 552
rect 1750 556 1756 557
rect 1750 552 1751 556
rect 1755 552 1756 556
rect 1750 551 1756 552
rect 1854 556 1860 557
rect 1854 552 1855 556
rect 1859 552 1860 556
rect 1854 551 1860 552
rect 1958 556 1964 557
rect 1958 552 1959 556
rect 1963 552 1964 556
rect 1958 551 1964 552
rect 2054 556 2060 557
rect 2054 552 2055 556
rect 2059 552 2060 556
rect 2054 551 2060 552
rect 2150 556 2156 557
rect 2150 552 2151 556
rect 2155 552 2156 556
rect 2150 551 2156 552
rect 2254 556 2260 557
rect 2254 552 2255 556
rect 2259 552 2260 556
rect 2254 551 2260 552
rect 2358 556 2364 557
rect 2358 552 2359 556
rect 2363 552 2364 556
rect 2358 551 2364 552
rect 2438 556 2444 557
rect 2438 552 2439 556
rect 2443 552 2444 556
rect 2438 551 2444 552
rect 2502 553 2508 554
rect 1326 548 1332 549
rect 2502 549 2503 553
rect 2507 549 2508 553
rect 2502 548 2508 549
rect 1166 547 1172 548
rect 1326 536 1332 537
rect 2502 536 2508 537
rect 142 532 148 533
rect 110 529 116 530
rect 110 525 111 529
rect 115 525 116 529
rect 142 528 143 532
rect 147 528 148 532
rect 142 527 148 528
rect 238 532 244 533
rect 238 528 239 532
rect 243 528 244 532
rect 238 527 244 528
rect 334 532 340 533
rect 334 528 335 532
rect 339 528 340 532
rect 334 527 340 528
rect 430 532 436 533
rect 430 528 431 532
rect 435 528 436 532
rect 430 527 436 528
rect 526 532 532 533
rect 526 528 527 532
rect 531 528 532 532
rect 526 527 532 528
rect 622 532 628 533
rect 622 528 623 532
rect 627 528 628 532
rect 622 527 628 528
rect 710 532 716 533
rect 710 528 711 532
rect 715 528 716 532
rect 710 527 716 528
rect 790 532 796 533
rect 790 528 791 532
rect 795 528 796 532
rect 790 527 796 528
rect 870 532 876 533
rect 870 528 871 532
rect 875 528 876 532
rect 870 527 876 528
rect 950 532 956 533
rect 950 528 951 532
rect 955 528 956 532
rect 950 527 956 528
rect 1030 532 1036 533
rect 1030 528 1031 532
rect 1035 528 1036 532
rect 1326 532 1327 536
rect 1331 532 1332 536
rect 1326 531 1332 532
rect 1390 535 1396 536
rect 1390 531 1391 535
rect 1395 531 1396 535
rect 1390 530 1396 531
rect 1470 535 1476 536
rect 1470 531 1471 535
rect 1475 531 1476 535
rect 1470 530 1476 531
rect 1566 535 1572 536
rect 1566 531 1567 535
rect 1571 531 1572 535
rect 1566 530 1572 531
rect 1662 535 1668 536
rect 1662 531 1663 535
rect 1667 531 1668 535
rect 1662 530 1668 531
rect 1766 535 1772 536
rect 1766 531 1767 535
rect 1771 531 1772 535
rect 1766 530 1772 531
rect 1870 535 1876 536
rect 1870 531 1871 535
rect 1875 531 1876 535
rect 1870 530 1876 531
rect 1974 535 1980 536
rect 1974 531 1975 535
rect 1979 531 1980 535
rect 1974 530 1980 531
rect 2070 535 2076 536
rect 2070 531 2071 535
rect 2075 531 2076 535
rect 2070 530 2076 531
rect 2166 535 2172 536
rect 2166 531 2167 535
rect 2171 531 2172 535
rect 2166 530 2172 531
rect 2270 535 2276 536
rect 2270 531 2271 535
rect 2275 531 2276 535
rect 2270 530 2276 531
rect 2374 535 2380 536
rect 2374 531 2375 535
rect 2379 531 2380 535
rect 2374 530 2380 531
rect 2454 535 2460 536
rect 2454 531 2455 535
rect 2459 531 2460 535
rect 2502 532 2503 536
rect 2507 532 2508 536
rect 2502 531 2508 532
rect 2454 530 2460 531
rect 1030 527 1036 528
rect 1286 529 1292 530
rect 110 524 116 525
rect 1286 525 1287 529
rect 1291 525 1292 529
rect 1286 524 1292 525
rect 110 512 116 513
rect 1286 512 1292 513
rect 110 508 111 512
rect 115 508 116 512
rect 110 507 116 508
rect 158 511 164 512
rect 158 507 159 511
rect 163 507 164 511
rect 158 506 164 507
rect 254 511 260 512
rect 254 507 255 511
rect 259 507 260 511
rect 254 506 260 507
rect 350 511 356 512
rect 350 507 351 511
rect 355 507 356 511
rect 350 506 356 507
rect 446 511 452 512
rect 446 507 447 511
rect 451 507 452 511
rect 446 506 452 507
rect 542 511 548 512
rect 542 507 543 511
rect 547 507 548 511
rect 542 506 548 507
rect 638 511 644 512
rect 638 507 639 511
rect 643 507 644 511
rect 638 506 644 507
rect 726 511 732 512
rect 726 507 727 511
rect 731 507 732 511
rect 726 506 732 507
rect 806 511 812 512
rect 806 507 807 511
rect 811 507 812 511
rect 806 506 812 507
rect 886 511 892 512
rect 886 507 887 511
rect 891 507 892 511
rect 886 506 892 507
rect 966 511 972 512
rect 966 507 967 511
rect 971 507 972 511
rect 966 506 972 507
rect 1046 511 1052 512
rect 1046 507 1047 511
rect 1051 507 1052 511
rect 1286 508 1287 512
rect 1291 508 1292 512
rect 1286 507 1292 508
rect 1046 506 1052 507
rect 1366 481 1372 482
rect 1326 480 1332 481
rect 1326 476 1327 480
rect 1331 476 1332 480
rect 1366 477 1367 481
rect 1371 477 1372 481
rect 1366 476 1372 477
rect 1454 481 1460 482
rect 1454 477 1455 481
rect 1459 477 1460 481
rect 1454 476 1460 477
rect 1574 481 1580 482
rect 1574 477 1575 481
rect 1579 477 1580 481
rect 1574 476 1580 477
rect 1694 481 1700 482
rect 1694 477 1695 481
rect 1699 477 1700 481
rect 1694 476 1700 477
rect 1806 481 1812 482
rect 1806 477 1807 481
rect 1811 477 1812 481
rect 1806 476 1812 477
rect 1918 481 1924 482
rect 1918 477 1919 481
rect 1923 477 1924 481
rect 1918 476 1924 477
rect 2022 481 2028 482
rect 2022 477 2023 481
rect 2027 477 2028 481
rect 2022 476 2028 477
rect 2118 481 2124 482
rect 2118 477 2119 481
rect 2123 477 2124 481
rect 2118 476 2124 477
rect 2206 481 2212 482
rect 2206 477 2207 481
rect 2211 477 2212 481
rect 2206 476 2212 477
rect 2294 481 2300 482
rect 2294 477 2295 481
rect 2299 477 2300 481
rect 2294 476 2300 477
rect 2382 481 2388 482
rect 2382 477 2383 481
rect 2387 477 2388 481
rect 2382 476 2388 477
rect 2454 481 2460 482
rect 2454 477 2455 481
rect 2459 477 2460 481
rect 2454 476 2460 477
rect 2502 480 2508 481
rect 2502 476 2503 480
rect 2507 476 2508 480
rect 1326 475 1332 476
rect 2502 475 2508 476
rect 1326 463 1332 464
rect 1326 459 1327 463
rect 1331 459 1332 463
rect 2502 463 2508 464
rect 1326 458 1332 459
rect 1350 460 1356 461
rect 150 457 156 458
rect 110 456 116 457
rect 110 452 111 456
rect 115 452 116 456
rect 150 453 151 457
rect 155 453 156 457
rect 150 452 156 453
rect 206 457 212 458
rect 206 453 207 457
rect 211 453 212 457
rect 206 452 212 453
rect 286 457 292 458
rect 286 453 287 457
rect 291 453 292 457
rect 286 452 292 453
rect 374 457 380 458
rect 374 453 375 457
rect 379 453 380 457
rect 374 452 380 453
rect 462 457 468 458
rect 462 453 463 457
rect 467 453 468 457
rect 462 452 468 453
rect 558 457 564 458
rect 558 453 559 457
rect 563 453 564 457
rect 558 452 564 453
rect 654 457 660 458
rect 654 453 655 457
rect 659 453 660 457
rect 654 452 660 453
rect 750 457 756 458
rect 750 453 751 457
rect 755 453 756 457
rect 750 452 756 453
rect 846 457 852 458
rect 846 453 847 457
rect 851 453 852 457
rect 846 452 852 453
rect 950 457 956 458
rect 950 453 951 457
rect 955 453 956 457
rect 950 452 956 453
rect 1054 457 1060 458
rect 1054 453 1055 457
rect 1059 453 1060 457
rect 1054 452 1060 453
rect 1158 457 1164 458
rect 1158 453 1159 457
rect 1163 453 1164 457
rect 1158 452 1164 453
rect 1238 457 1244 458
rect 1238 453 1239 457
rect 1243 453 1244 457
rect 1238 452 1244 453
rect 1286 456 1292 457
rect 1286 452 1287 456
rect 1291 452 1292 456
rect 1350 456 1351 460
rect 1355 456 1356 460
rect 1350 455 1356 456
rect 1438 460 1444 461
rect 1438 456 1439 460
rect 1443 456 1444 460
rect 1438 455 1444 456
rect 1558 460 1564 461
rect 1558 456 1559 460
rect 1563 456 1564 460
rect 1558 455 1564 456
rect 1678 460 1684 461
rect 1678 456 1679 460
rect 1683 456 1684 460
rect 1678 455 1684 456
rect 1790 460 1796 461
rect 1790 456 1791 460
rect 1795 456 1796 460
rect 1790 455 1796 456
rect 1902 460 1908 461
rect 1902 456 1903 460
rect 1907 456 1908 460
rect 1902 455 1908 456
rect 2006 460 2012 461
rect 2006 456 2007 460
rect 2011 456 2012 460
rect 2006 455 2012 456
rect 2102 460 2108 461
rect 2102 456 2103 460
rect 2107 456 2108 460
rect 2102 455 2108 456
rect 2190 460 2196 461
rect 2190 456 2191 460
rect 2195 456 2196 460
rect 2190 455 2196 456
rect 2278 460 2284 461
rect 2278 456 2279 460
rect 2283 456 2284 460
rect 2278 455 2284 456
rect 2366 460 2372 461
rect 2366 456 2367 460
rect 2371 456 2372 460
rect 2366 455 2372 456
rect 2438 460 2444 461
rect 2438 456 2439 460
rect 2443 456 2444 460
rect 2502 459 2503 463
rect 2507 459 2508 463
rect 2502 458 2508 459
rect 2438 455 2444 456
rect 110 451 116 452
rect 1286 451 1292 452
rect 110 439 116 440
rect 110 435 111 439
rect 115 435 116 439
rect 1286 439 1292 440
rect 110 434 116 435
rect 134 436 140 437
rect 134 432 135 436
rect 139 432 140 436
rect 134 431 140 432
rect 190 436 196 437
rect 190 432 191 436
rect 195 432 196 436
rect 190 431 196 432
rect 270 436 276 437
rect 270 432 271 436
rect 275 432 276 436
rect 270 431 276 432
rect 358 436 364 437
rect 358 432 359 436
rect 363 432 364 436
rect 358 431 364 432
rect 446 436 452 437
rect 446 432 447 436
rect 451 432 452 436
rect 446 431 452 432
rect 542 436 548 437
rect 542 432 543 436
rect 547 432 548 436
rect 542 431 548 432
rect 638 436 644 437
rect 638 432 639 436
rect 643 432 644 436
rect 638 431 644 432
rect 734 436 740 437
rect 734 432 735 436
rect 739 432 740 436
rect 734 431 740 432
rect 830 436 836 437
rect 830 432 831 436
rect 835 432 836 436
rect 830 431 836 432
rect 934 436 940 437
rect 934 432 935 436
rect 939 432 940 436
rect 934 431 940 432
rect 1038 436 1044 437
rect 1038 432 1039 436
rect 1043 432 1044 436
rect 1038 431 1044 432
rect 1142 436 1148 437
rect 1142 432 1143 436
rect 1147 432 1148 436
rect 1142 431 1148 432
rect 1222 436 1228 437
rect 1222 432 1223 436
rect 1227 432 1228 436
rect 1286 435 1287 439
rect 1291 435 1292 439
rect 1286 434 1292 435
rect 1582 436 1588 437
rect 1222 431 1228 432
rect 1326 433 1332 434
rect 1326 429 1327 433
rect 1331 429 1332 433
rect 1582 432 1583 436
rect 1587 432 1588 436
rect 1582 431 1588 432
rect 1638 436 1644 437
rect 1638 432 1639 436
rect 1643 432 1644 436
rect 1638 431 1644 432
rect 1694 436 1700 437
rect 1694 432 1695 436
rect 1699 432 1700 436
rect 1694 431 1700 432
rect 1758 436 1764 437
rect 1758 432 1759 436
rect 1763 432 1764 436
rect 1758 431 1764 432
rect 1830 436 1836 437
rect 1830 432 1831 436
rect 1835 432 1836 436
rect 1830 431 1836 432
rect 1910 436 1916 437
rect 1910 432 1911 436
rect 1915 432 1916 436
rect 1910 431 1916 432
rect 1990 436 1996 437
rect 1990 432 1991 436
rect 1995 432 1996 436
rect 1990 431 1996 432
rect 2078 436 2084 437
rect 2078 432 2079 436
rect 2083 432 2084 436
rect 2078 431 2084 432
rect 2174 436 2180 437
rect 2174 432 2175 436
rect 2179 432 2180 436
rect 2174 431 2180 432
rect 2270 436 2276 437
rect 2270 432 2271 436
rect 2275 432 2276 436
rect 2270 431 2276 432
rect 2366 436 2372 437
rect 2366 432 2367 436
rect 2371 432 2372 436
rect 2366 431 2372 432
rect 2438 436 2444 437
rect 2438 432 2439 436
rect 2443 432 2444 436
rect 2438 431 2444 432
rect 2502 433 2508 434
rect 1326 428 1332 429
rect 2502 429 2503 433
rect 2507 429 2508 433
rect 2502 428 2508 429
rect 134 424 140 425
rect 110 421 116 422
rect 110 417 111 421
rect 115 417 116 421
rect 134 420 135 424
rect 139 420 140 424
rect 134 419 140 420
rect 190 424 196 425
rect 190 420 191 424
rect 195 420 196 424
rect 190 419 196 420
rect 278 424 284 425
rect 278 420 279 424
rect 283 420 284 424
rect 278 419 284 420
rect 382 424 388 425
rect 382 420 383 424
rect 387 420 388 424
rect 382 419 388 420
rect 494 424 500 425
rect 494 420 495 424
rect 499 420 500 424
rect 494 419 500 420
rect 606 424 612 425
rect 606 420 607 424
rect 611 420 612 424
rect 606 419 612 420
rect 718 424 724 425
rect 718 420 719 424
rect 723 420 724 424
rect 718 419 724 420
rect 830 424 836 425
rect 830 420 831 424
rect 835 420 836 424
rect 830 419 836 420
rect 934 424 940 425
rect 934 420 935 424
rect 939 420 940 424
rect 934 419 940 420
rect 1038 424 1044 425
rect 1038 420 1039 424
rect 1043 420 1044 424
rect 1038 419 1044 420
rect 1142 424 1148 425
rect 1142 420 1143 424
rect 1147 420 1148 424
rect 1142 419 1148 420
rect 1222 424 1228 425
rect 1222 420 1223 424
rect 1227 420 1228 424
rect 1222 419 1228 420
rect 1286 421 1292 422
rect 110 416 116 417
rect 1286 417 1287 421
rect 1291 417 1292 421
rect 1286 416 1292 417
rect 1326 416 1332 417
rect 2502 416 2508 417
rect 1326 412 1327 416
rect 1331 412 1332 416
rect 1326 411 1332 412
rect 1598 415 1604 416
rect 1598 411 1599 415
rect 1603 411 1604 415
rect 1598 410 1604 411
rect 1654 415 1660 416
rect 1654 411 1655 415
rect 1659 411 1660 415
rect 1654 410 1660 411
rect 1710 415 1716 416
rect 1710 411 1711 415
rect 1715 411 1716 415
rect 1710 410 1716 411
rect 1774 415 1780 416
rect 1774 411 1775 415
rect 1779 411 1780 415
rect 1774 410 1780 411
rect 1846 415 1852 416
rect 1846 411 1847 415
rect 1851 411 1852 415
rect 1846 410 1852 411
rect 1926 415 1932 416
rect 1926 411 1927 415
rect 1931 411 1932 415
rect 1926 410 1932 411
rect 2006 415 2012 416
rect 2006 411 2007 415
rect 2011 411 2012 415
rect 2006 410 2012 411
rect 2094 415 2100 416
rect 2094 411 2095 415
rect 2099 411 2100 415
rect 2094 410 2100 411
rect 2190 415 2196 416
rect 2190 411 2191 415
rect 2195 411 2196 415
rect 2190 410 2196 411
rect 2286 415 2292 416
rect 2286 411 2287 415
rect 2291 411 2292 415
rect 2286 410 2292 411
rect 2382 415 2388 416
rect 2382 411 2383 415
rect 2387 411 2388 415
rect 2382 410 2388 411
rect 2454 415 2460 416
rect 2454 411 2455 415
rect 2459 411 2460 415
rect 2502 412 2503 416
rect 2507 412 2508 416
rect 2502 411 2508 412
rect 2454 410 2460 411
rect 110 404 116 405
rect 1286 404 1292 405
rect 110 400 111 404
rect 115 400 116 404
rect 110 399 116 400
rect 150 403 156 404
rect 150 399 151 403
rect 155 399 156 403
rect 150 398 156 399
rect 206 403 212 404
rect 206 399 207 403
rect 211 399 212 403
rect 206 398 212 399
rect 294 403 300 404
rect 294 399 295 403
rect 299 399 300 403
rect 294 398 300 399
rect 398 403 404 404
rect 398 399 399 403
rect 403 399 404 403
rect 398 398 404 399
rect 510 403 516 404
rect 510 399 511 403
rect 515 399 516 403
rect 510 398 516 399
rect 622 403 628 404
rect 622 399 623 403
rect 627 399 628 403
rect 622 398 628 399
rect 734 403 740 404
rect 734 399 735 403
rect 739 399 740 403
rect 734 398 740 399
rect 846 403 852 404
rect 846 399 847 403
rect 851 399 852 403
rect 846 398 852 399
rect 950 403 956 404
rect 950 399 951 403
rect 955 399 956 403
rect 950 398 956 399
rect 1054 403 1060 404
rect 1054 399 1055 403
rect 1059 399 1060 403
rect 1054 398 1060 399
rect 1158 403 1164 404
rect 1158 399 1159 403
rect 1163 399 1164 403
rect 1158 398 1164 399
rect 1238 403 1244 404
rect 1238 399 1239 403
rect 1243 399 1244 403
rect 1286 400 1287 404
rect 1291 400 1292 404
rect 1286 399 1292 400
rect 1238 398 1244 399
rect 1678 361 1684 362
rect 1326 360 1332 361
rect 1326 356 1327 360
rect 1331 356 1332 360
rect 1678 357 1679 361
rect 1683 357 1684 361
rect 1678 356 1684 357
rect 1734 361 1740 362
rect 1734 357 1735 361
rect 1739 357 1740 361
rect 1734 356 1740 357
rect 1798 361 1804 362
rect 1798 357 1799 361
rect 1803 357 1804 361
rect 1798 356 1804 357
rect 1870 361 1876 362
rect 1870 357 1871 361
rect 1875 357 1876 361
rect 1870 356 1876 357
rect 1942 361 1948 362
rect 1942 357 1943 361
rect 1947 357 1948 361
rect 1942 356 1948 357
rect 2022 361 2028 362
rect 2022 357 2023 361
rect 2027 357 2028 361
rect 2022 356 2028 357
rect 2110 361 2116 362
rect 2110 357 2111 361
rect 2115 357 2116 361
rect 2110 356 2116 357
rect 2198 361 2204 362
rect 2198 357 2199 361
rect 2203 357 2204 361
rect 2198 356 2204 357
rect 2286 361 2292 362
rect 2286 357 2287 361
rect 2291 357 2292 361
rect 2286 356 2292 357
rect 2374 361 2380 362
rect 2374 357 2375 361
rect 2379 357 2380 361
rect 2374 356 2380 357
rect 2454 361 2460 362
rect 2454 357 2455 361
rect 2459 357 2460 361
rect 2454 356 2460 357
rect 2502 360 2508 361
rect 2502 356 2503 360
rect 2507 356 2508 360
rect 1326 355 1332 356
rect 2502 355 2508 356
rect 150 349 156 350
rect 110 348 116 349
rect 110 344 111 348
rect 115 344 116 348
rect 150 345 151 349
rect 155 345 156 349
rect 150 344 156 345
rect 230 349 236 350
rect 230 345 231 349
rect 235 345 236 349
rect 230 344 236 345
rect 334 349 340 350
rect 334 345 335 349
rect 339 345 340 349
rect 334 344 340 345
rect 438 349 444 350
rect 438 345 439 349
rect 443 345 444 349
rect 438 344 444 345
rect 542 349 548 350
rect 542 345 543 349
rect 547 345 548 349
rect 542 344 548 345
rect 646 349 652 350
rect 646 345 647 349
rect 651 345 652 349
rect 646 344 652 345
rect 750 349 756 350
rect 750 345 751 349
rect 755 345 756 349
rect 750 344 756 345
rect 846 349 852 350
rect 846 345 847 349
rect 851 345 852 349
rect 846 344 852 345
rect 934 349 940 350
rect 934 345 935 349
rect 939 345 940 349
rect 934 344 940 345
rect 1014 349 1020 350
rect 1014 345 1015 349
rect 1019 345 1020 349
rect 1014 344 1020 345
rect 1094 349 1100 350
rect 1094 345 1095 349
rect 1099 345 1100 349
rect 1094 344 1100 345
rect 1174 349 1180 350
rect 1174 345 1175 349
rect 1179 345 1180 349
rect 1174 344 1180 345
rect 1238 349 1244 350
rect 1238 345 1239 349
rect 1243 345 1244 349
rect 1238 344 1244 345
rect 1286 348 1292 349
rect 1286 344 1287 348
rect 1291 344 1292 348
rect 110 343 116 344
rect 1286 343 1292 344
rect 1326 343 1332 344
rect 1326 339 1327 343
rect 1331 339 1332 343
rect 2502 343 2508 344
rect 1326 338 1332 339
rect 1662 340 1668 341
rect 1662 336 1663 340
rect 1667 336 1668 340
rect 1662 335 1668 336
rect 1718 340 1724 341
rect 1718 336 1719 340
rect 1723 336 1724 340
rect 1718 335 1724 336
rect 1782 340 1788 341
rect 1782 336 1783 340
rect 1787 336 1788 340
rect 1782 335 1788 336
rect 1854 340 1860 341
rect 1854 336 1855 340
rect 1859 336 1860 340
rect 1854 335 1860 336
rect 1926 340 1932 341
rect 1926 336 1927 340
rect 1931 336 1932 340
rect 1926 335 1932 336
rect 2006 340 2012 341
rect 2006 336 2007 340
rect 2011 336 2012 340
rect 2006 335 2012 336
rect 2094 340 2100 341
rect 2094 336 2095 340
rect 2099 336 2100 340
rect 2094 335 2100 336
rect 2182 340 2188 341
rect 2182 336 2183 340
rect 2187 336 2188 340
rect 2182 335 2188 336
rect 2270 340 2276 341
rect 2270 336 2271 340
rect 2275 336 2276 340
rect 2270 335 2276 336
rect 2358 340 2364 341
rect 2358 336 2359 340
rect 2363 336 2364 340
rect 2358 335 2364 336
rect 2438 340 2444 341
rect 2438 336 2439 340
rect 2443 336 2444 340
rect 2502 339 2503 343
rect 2507 339 2508 343
rect 2502 338 2508 339
rect 2438 335 2444 336
rect 110 331 116 332
rect 110 327 111 331
rect 115 327 116 331
rect 1286 331 1292 332
rect 110 326 116 327
rect 134 328 140 329
rect 134 324 135 328
rect 139 324 140 328
rect 134 323 140 324
rect 214 328 220 329
rect 214 324 215 328
rect 219 324 220 328
rect 214 323 220 324
rect 318 328 324 329
rect 318 324 319 328
rect 323 324 324 328
rect 318 323 324 324
rect 422 328 428 329
rect 422 324 423 328
rect 427 324 428 328
rect 422 323 428 324
rect 526 328 532 329
rect 526 324 527 328
rect 531 324 532 328
rect 526 323 532 324
rect 630 328 636 329
rect 630 324 631 328
rect 635 324 636 328
rect 630 323 636 324
rect 734 328 740 329
rect 734 324 735 328
rect 739 324 740 328
rect 734 323 740 324
rect 830 328 836 329
rect 830 324 831 328
rect 835 324 836 328
rect 830 323 836 324
rect 918 328 924 329
rect 918 324 919 328
rect 923 324 924 328
rect 918 323 924 324
rect 998 328 1004 329
rect 998 324 999 328
rect 1003 324 1004 328
rect 998 323 1004 324
rect 1078 328 1084 329
rect 1078 324 1079 328
rect 1083 324 1084 328
rect 1078 323 1084 324
rect 1158 328 1164 329
rect 1158 324 1159 328
rect 1163 324 1164 328
rect 1158 323 1164 324
rect 1222 328 1228 329
rect 1222 324 1223 328
rect 1227 324 1228 328
rect 1286 327 1287 331
rect 1291 327 1292 331
rect 1286 326 1292 327
rect 1222 323 1228 324
rect 1350 320 1356 321
rect 1326 317 1332 318
rect 1326 313 1327 317
rect 1331 313 1332 317
rect 1350 316 1351 320
rect 1355 316 1356 320
rect 1350 315 1356 316
rect 1454 320 1460 321
rect 1454 316 1455 320
rect 1459 316 1460 320
rect 1454 315 1460 316
rect 1582 320 1588 321
rect 1582 316 1583 320
rect 1587 316 1588 320
rect 1582 315 1588 316
rect 1710 320 1716 321
rect 1710 316 1711 320
rect 1715 316 1716 320
rect 1710 315 1716 316
rect 1838 320 1844 321
rect 1838 316 1839 320
rect 1843 316 1844 320
rect 1838 315 1844 316
rect 1950 320 1956 321
rect 1950 316 1951 320
rect 1955 316 1956 320
rect 1950 315 1956 316
rect 2062 320 2068 321
rect 2062 316 2063 320
rect 2067 316 2068 320
rect 2062 315 2068 316
rect 2166 320 2172 321
rect 2166 316 2167 320
rect 2171 316 2172 320
rect 2166 315 2172 316
rect 2262 320 2268 321
rect 2262 316 2263 320
rect 2267 316 2268 320
rect 2262 315 2268 316
rect 2358 320 2364 321
rect 2358 316 2359 320
rect 2363 316 2364 320
rect 2358 315 2364 316
rect 2438 320 2444 321
rect 2438 316 2439 320
rect 2443 316 2444 320
rect 2438 315 2444 316
rect 2502 317 2508 318
rect 134 312 140 313
rect 110 309 116 310
rect 110 305 111 309
rect 115 305 116 309
rect 134 308 135 312
rect 139 308 140 312
rect 134 307 140 308
rect 214 312 220 313
rect 214 308 215 312
rect 219 308 220 312
rect 214 307 220 308
rect 318 312 324 313
rect 318 308 319 312
rect 323 308 324 312
rect 318 307 324 308
rect 422 312 428 313
rect 422 308 423 312
rect 427 308 428 312
rect 422 307 428 308
rect 534 312 540 313
rect 534 308 535 312
rect 539 308 540 312
rect 534 307 540 308
rect 638 312 644 313
rect 638 308 639 312
rect 643 308 644 312
rect 638 307 644 308
rect 742 312 748 313
rect 742 308 743 312
rect 747 308 748 312
rect 742 307 748 308
rect 846 312 852 313
rect 846 308 847 312
rect 851 308 852 312
rect 846 307 852 308
rect 942 312 948 313
rect 942 308 943 312
rect 947 308 948 312
rect 942 307 948 308
rect 1038 312 1044 313
rect 1038 308 1039 312
rect 1043 308 1044 312
rect 1038 307 1044 308
rect 1142 312 1148 313
rect 1142 308 1143 312
rect 1147 308 1148 312
rect 1142 307 1148 308
rect 1222 312 1228 313
rect 1326 312 1332 313
rect 2502 313 2503 317
rect 2507 313 2508 317
rect 2502 312 2508 313
rect 1222 308 1223 312
rect 1227 308 1228 312
rect 1222 307 1228 308
rect 1286 309 1292 310
rect 110 304 116 305
rect 1286 305 1287 309
rect 1291 305 1292 309
rect 1286 304 1292 305
rect 1326 300 1332 301
rect 2502 300 2508 301
rect 1326 296 1327 300
rect 1331 296 1332 300
rect 1326 295 1332 296
rect 1366 299 1372 300
rect 1366 295 1367 299
rect 1371 295 1372 299
rect 1366 294 1372 295
rect 1470 299 1476 300
rect 1470 295 1471 299
rect 1475 295 1476 299
rect 1470 294 1476 295
rect 1598 299 1604 300
rect 1598 295 1599 299
rect 1603 295 1604 299
rect 1598 294 1604 295
rect 1726 299 1732 300
rect 1726 295 1727 299
rect 1731 295 1732 299
rect 1726 294 1732 295
rect 1854 299 1860 300
rect 1854 295 1855 299
rect 1859 295 1860 299
rect 1854 294 1860 295
rect 1966 299 1972 300
rect 1966 295 1967 299
rect 1971 295 1972 299
rect 1966 294 1972 295
rect 2078 299 2084 300
rect 2078 295 2079 299
rect 2083 295 2084 299
rect 2078 294 2084 295
rect 2182 299 2188 300
rect 2182 295 2183 299
rect 2187 295 2188 299
rect 2182 294 2188 295
rect 2278 299 2284 300
rect 2278 295 2279 299
rect 2283 295 2284 299
rect 2278 294 2284 295
rect 2374 299 2380 300
rect 2374 295 2375 299
rect 2379 295 2380 299
rect 2374 294 2380 295
rect 2454 299 2460 300
rect 2454 295 2455 299
rect 2459 295 2460 299
rect 2502 296 2503 300
rect 2507 296 2508 300
rect 2502 295 2508 296
rect 2454 294 2460 295
rect 110 292 116 293
rect 1286 292 1292 293
rect 110 288 111 292
rect 115 288 116 292
rect 110 287 116 288
rect 150 291 156 292
rect 150 287 151 291
rect 155 287 156 291
rect 150 286 156 287
rect 230 291 236 292
rect 230 287 231 291
rect 235 287 236 291
rect 230 286 236 287
rect 334 291 340 292
rect 334 287 335 291
rect 339 287 340 291
rect 334 286 340 287
rect 438 291 444 292
rect 438 287 439 291
rect 443 287 444 291
rect 438 286 444 287
rect 550 291 556 292
rect 550 287 551 291
rect 555 287 556 291
rect 550 286 556 287
rect 654 291 660 292
rect 654 287 655 291
rect 659 287 660 291
rect 654 286 660 287
rect 758 291 764 292
rect 758 287 759 291
rect 763 287 764 291
rect 758 286 764 287
rect 862 291 868 292
rect 862 287 863 291
rect 867 287 868 291
rect 862 286 868 287
rect 958 291 964 292
rect 958 287 959 291
rect 963 287 964 291
rect 958 286 964 287
rect 1054 291 1060 292
rect 1054 287 1055 291
rect 1059 287 1060 291
rect 1054 286 1060 287
rect 1158 291 1164 292
rect 1158 287 1159 291
rect 1163 287 1164 291
rect 1158 286 1164 287
rect 1238 291 1244 292
rect 1238 287 1239 291
rect 1243 287 1244 291
rect 1286 288 1287 292
rect 1291 288 1292 292
rect 1286 287 1292 288
rect 1238 286 1244 287
rect 150 241 156 242
rect 110 240 116 241
rect 110 236 111 240
rect 115 236 116 240
rect 150 237 151 241
rect 155 237 156 241
rect 150 236 156 237
rect 222 241 228 242
rect 222 237 223 241
rect 227 237 228 241
rect 222 236 228 237
rect 318 241 324 242
rect 318 237 319 241
rect 323 237 324 241
rect 318 236 324 237
rect 422 241 428 242
rect 422 237 423 241
rect 427 237 428 241
rect 422 236 428 237
rect 534 241 540 242
rect 534 237 535 241
rect 539 237 540 241
rect 534 236 540 237
rect 646 241 652 242
rect 646 237 647 241
rect 651 237 652 241
rect 646 236 652 237
rect 758 241 764 242
rect 758 237 759 241
rect 763 237 764 241
rect 758 236 764 237
rect 870 241 876 242
rect 870 237 871 241
rect 875 237 876 241
rect 870 236 876 237
rect 982 241 988 242
rect 982 237 983 241
rect 987 237 988 241
rect 982 236 988 237
rect 1102 241 1108 242
rect 1102 237 1103 241
rect 1107 237 1108 241
rect 1102 236 1108 237
rect 1222 241 1228 242
rect 1366 241 1372 242
rect 1222 237 1223 241
rect 1227 237 1228 241
rect 1222 236 1228 237
rect 1286 240 1292 241
rect 1286 236 1287 240
rect 1291 236 1292 240
rect 110 235 116 236
rect 1286 235 1292 236
rect 1326 240 1332 241
rect 1326 236 1327 240
rect 1331 236 1332 240
rect 1366 237 1367 241
rect 1371 237 1372 241
rect 1366 236 1372 237
rect 1446 241 1452 242
rect 1446 237 1447 241
rect 1451 237 1452 241
rect 1446 236 1452 237
rect 1550 241 1556 242
rect 1550 237 1551 241
rect 1555 237 1556 241
rect 1550 236 1556 237
rect 1654 241 1660 242
rect 1654 237 1655 241
rect 1659 237 1660 241
rect 1654 236 1660 237
rect 1758 241 1764 242
rect 1758 237 1759 241
rect 1763 237 1764 241
rect 1758 236 1764 237
rect 1862 241 1868 242
rect 1862 237 1863 241
rect 1867 237 1868 241
rect 1862 236 1868 237
rect 1966 241 1972 242
rect 1966 237 1967 241
rect 1971 237 1972 241
rect 1966 236 1972 237
rect 2070 241 2076 242
rect 2070 237 2071 241
rect 2075 237 2076 241
rect 2070 236 2076 237
rect 2174 241 2180 242
rect 2174 237 2175 241
rect 2179 237 2180 241
rect 2174 236 2180 237
rect 2270 241 2276 242
rect 2270 237 2271 241
rect 2275 237 2276 241
rect 2270 236 2276 237
rect 2374 241 2380 242
rect 2374 237 2375 241
rect 2379 237 2380 241
rect 2374 236 2380 237
rect 2454 241 2460 242
rect 2454 237 2455 241
rect 2459 237 2460 241
rect 2454 236 2460 237
rect 2502 240 2508 241
rect 2502 236 2503 240
rect 2507 236 2508 240
rect 1326 235 1332 236
rect 2502 235 2508 236
rect 110 223 116 224
rect 110 219 111 223
rect 115 219 116 223
rect 1286 223 1292 224
rect 110 218 116 219
rect 134 220 140 221
rect 134 216 135 220
rect 139 216 140 220
rect 134 215 140 216
rect 206 220 212 221
rect 206 216 207 220
rect 211 216 212 220
rect 206 215 212 216
rect 302 220 308 221
rect 302 216 303 220
rect 307 216 308 220
rect 302 215 308 216
rect 406 220 412 221
rect 406 216 407 220
rect 411 216 412 220
rect 406 215 412 216
rect 518 220 524 221
rect 518 216 519 220
rect 523 216 524 220
rect 518 215 524 216
rect 630 220 636 221
rect 630 216 631 220
rect 635 216 636 220
rect 630 215 636 216
rect 742 220 748 221
rect 742 216 743 220
rect 747 216 748 220
rect 742 215 748 216
rect 854 220 860 221
rect 854 216 855 220
rect 859 216 860 220
rect 854 215 860 216
rect 966 220 972 221
rect 966 216 967 220
rect 971 216 972 220
rect 966 215 972 216
rect 1086 220 1092 221
rect 1086 216 1087 220
rect 1091 216 1092 220
rect 1086 215 1092 216
rect 1206 220 1212 221
rect 1206 216 1207 220
rect 1211 216 1212 220
rect 1286 219 1287 223
rect 1291 219 1292 223
rect 1286 218 1292 219
rect 1326 223 1332 224
rect 1326 219 1327 223
rect 1331 219 1332 223
rect 2502 223 2508 224
rect 1326 218 1332 219
rect 1350 220 1356 221
rect 1206 215 1212 216
rect 1350 216 1351 220
rect 1355 216 1356 220
rect 1350 215 1356 216
rect 1430 220 1436 221
rect 1430 216 1431 220
rect 1435 216 1436 220
rect 1430 215 1436 216
rect 1534 220 1540 221
rect 1534 216 1535 220
rect 1539 216 1540 220
rect 1534 215 1540 216
rect 1638 220 1644 221
rect 1638 216 1639 220
rect 1643 216 1644 220
rect 1638 215 1644 216
rect 1742 220 1748 221
rect 1742 216 1743 220
rect 1747 216 1748 220
rect 1742 215 1748 216
rect 1846 220 1852 221
rect 1846 216 1847 220
rect 1851 216 1852 220
rect 1846 215 1852 216
rect 1950 220 1956 221
rect 1950 216 1951 220
rect 1955 216 1956 220
rect 1950 215 1956 216
rect 2054 220 2060 221
rect 2054 216 2055 220
rect 2059 216 2060 220
rect 2054 215 2060 216
rect 2158 220 2164 221
rect 2158 216 2159 220
rect 2163 216 2164 220
rect 2158 215 2164 216
rect 2254 220 2260 221
rect 2254 216 2255 220
rect 2259 216 2260 220
rect 2254 215 2260 216
rect 2358 220 2364 221
rect 2358 216 2359 220
rect 2363 216 2364 220
rect 2358 215 2364 216
rect 2438 220 2444 221
rect 2438 216 2439 220
rect 2443 216 2444 220
rect 2502 219 2503 223
rect 2507 219 2508 223
rect 2502 218 2508 219
rect 2438 215 2444 216
rect 182 204 188 205
rect 110 201 116 202
rect 110 197 111 201
rect 115 197 116 201
rect 182 200 183 204
rect 187 200 188 204
rect 182 199 188 200
rect 278 204 284 205
rect 278 200 279 204
rect 283 200 284 204
rect 278 199 284 200
rect 382 204 388 205
rect 382 200 383 204
rect 387 200 388 204
rect 382 199 388 200
rect 486 204 492 205
rect 486 200 487 204
rect 491 200 492 204
rect 486 199 492 200
rect 590 204 596 205
rect 590 200 591 204
rect 595 200 596 204
rect 590 199 596 200
rect 694 204 700 205
rect 694 200 695 204
rect 699 200 700 204
rect 694 199 700 200
rect 798 204 804 205
rect 798 200 799 204
rect 803 200 804 204
rect 798 199 804 200
rect 894 204 900 205
rect 894 200 895 204
rect 899 200 900 204
rect 894 199 900 200
rect 998 204 1004 205
rect 998 200 999 204
rect 1003 200 1004 204
rect 998 199 1004 200
rect 1102 204 1108 205
rect 1102 200 1103 204
rect 1107 200 1108 204
rect 1350 204 1356 205
rect 1102 199 1108 200
rect 1286 201 1292 202
rect 110 196 116 197
rect 1286 197 1287 201
rect 1291 197 1292 201
rect 1286 196 1292 197
rect 1326 201 1332 202
rect 1326 197 1327 201
rect 1331 197 1332 201
rect 1350 200 1351 204
rect 1355 200 1356 204
rect 1350 199 1356 200
rect 1406 204 1412 205
rect 1406 200 1407 204
rect 1411 200 1412 204
rect 1406 199 1412 200
rect 1470 204 1476 205
rect 1470 200 1471 204
rect 1475 200 1476 204
rect 1470 199 1476 200
rect 1550 204 1556 205
rect 1550 200 1551 204
rect 1555 200 1556 204
rect 1550 199 1556 200
rect 1638 204 1644 205
rect 1638 200 1639 204
rect 1643 200 1644 204
rect 1638 199 1644 200
rect 1718 204 1724 205
rect 1718 200 1719 204
rect 1723 200 1724 204
rect 1718 199 1724 200
rect 1806 204 1812 205
rect 1806 200 1807 204
rect 1811 200 1812 204
rect 1806 199 1812 200
rect 1894 204 1900 205
rect 1894 200 1895 204
rect 1899 200 1900 204
rect 1894 199 1900 200
rect 1990 204 1996 205
rect 1990 200 1991 204
rect 1995 200 1996 204
rect 1990 199 1996 200
rect 2102 204 2108 205
rect 2102 200 2103 204
rect 2107 200 2108 204
rect 2102 199 2108 200
rect 2214 204 2220 205
rect 2214 200 2215 204
rect 2219 200 2220 204
rect 2214 199 2220 200
rect 2334 204 2340 205
rect 2334 200 2335 204
rect 2339 200 2340 204
rect 2334 199 2340 200
rect 2438 204 2444 205
rect 2438 200 2439 204
rect 2443 200 2444 204
rect 2438 199 2444 200
rect 2502 201 2508 202
rect 1326 196 1332 197
rect 2502 197 2503 201
rect 2507 197 2508 201
rect 2502 196 2508 197
rect 110 184 116 185
rect 1286 184 1292 185
rect 110 180 111 184
rect 115 180 116 184
rect 110 179 116 180
rect 198 183 204 184
rect 198 179 199 183
rect 203 179 204 183
rect 198 178 204 179
rect 294 183 300 184
rect 294 179 295 183
rect 299 179 300 183
rect 294 178 300 179
rect 398 183 404 184
rect 398 179 399 183
rect 403 179 404 183
rect 398 178 404 179
rect 502 183 508 184
rect 502 179 503 183
rect 507 179 508 183
rect 502 178 508 179
rect 606 183 612 184
rect 606 179 607 183
rect 611 179 612 183
rect 606 178 612 179
rect 710 183 716 184
rect 710 179 711 183
rect 715 179 716 183
rect 710 178 716 179
rect 814 183 820 184
rect 814 179 815 183
rect 819 179 820 183
rect 814 178 820 179
rect 910 183 916 184
rect 910 179 911 183
rect 915 179 916 183
rect 910 178 916 179
rect 1014 183 1020 184
rect 1014 179 1015 183
rect 1019 179 1020 183
rect 1014 178 1020 179
rect 1118 183 1124 184
rect 1118 179 1119 183
rect 1123 179 1124 183
rect 1286 180 1287 184
rect 1291 180 1292 184
rect 1286 179 1292 180
rect 1326 184 1332 185
rect 2502 184 2508 185
rect 1326 180 1327 184
rect 1331 180 1332 184
rect 1326 179 1332 180
rect 1366 183 1372 184
rect 1366 179 1367 183
rect 1371 179 1372 183
rect 1118 178 1124 179
rect 1366 178 1372 179
rect 1422 183 1428 184
rect 1422 179 1423 183
rect 1427 179 1428 183
rect 1422 178 1428 179
rect 1486 183 1492 184
rect 1486 179 1487 183
rect 1491 179 1492 183
rect 1486 178 1492 179
rect 1566 183 1572 184
rect 1566 179 1567 183
rect 1571 179 1572 183
rect 1566 178 1572 179
rect 1654 183 1660 184
rect 1654 179 1655 183
rect 1659 179 1660 183
rect 1654 178 1660 179
rect 1734 183 1740 184
rect 1734 179 1735 183
rect 1739 179 1740 183
rect 1734 178 1740 179
rect 1822 183 1828 184
rect 1822 179 1823 183
rect 1827 179 1828 183
rect 1822 178 1828 179
rect 1910 183 1916 184
rect 1910 179 1911 183
rect 1915 179 1916 183
rect 1910 178 1916 179
rect 2006 183 2012 184
rect 2006 179 2007 183
rect 2011 179 2012 183
rect 2006 178 2012 179
rect 2118 183 2124 184
rect 2118 179 2119 183
rect 2123 179 2124 183
rect 2118 178 2124 179
rect 2230 183 2236 184
rect 2230 179 2231 183
rect 2235 179 2236 183
rect 2230 178 2236 179
rect 2350 183 2356 184
rect 2350 179 2351 183
rect 2355 179 2356 183
rect 2350 178 2356 179
rect 2454 183 2460 184
rect 2454 179 2455 183
rect 2459 179 2460 183
rect 2502 180 2503 184
rect 2507 180 2508 184
rect 2502 179 2508 180
rect 2454 178 2460 179
rect 150 125 156 126
rect 110 124 116 125
rect 110 120 111 124
rect 115 120 116 124
rect 150 121 151 125
rect 155 121 156 125
rect 150 120 156 121
rect 206 125 212 126
rect 206 121 207 125
rect 211 121 212 125
rect 206 120 212 121
rect 262 125 268 126
rect 262 121 263 125
rect 267 121 268 125
rect 262 120 268 121
rect 318 125 324 126
rect 318 121 319 125
rect 323 121 324 125
rect 318 120 324 121
rect 374 125 380 126
rect 374 121 375 125
rect 379 121 380 125
rect 374 120 380 121
rect 430 125 436 126
rect 430 121 431 125
rect 435 121 436 125
rect 430 120 436 121
rect 486 125 492 126
rect 486 121 487 125
rect 491 121 492 125
rect 486 120 492 121
rect 542 125 548 126
rect 542 121 543 125
rect 547 121 548 125
rect 542 120 548 121
rect 598 125 604 126
rect 598 121 599 125
rect 603 121 604 125
rect 598 120 604 121
rect 654 125 660 126
rect 654 121 655 125
rect 659 121 660 125
rect 654 120 660 121
rect 710 125 716 126
rect 710 121 711 125
rect 715 121 716 125
rect 710 120 716 121
rect 766 125 772 126
rect 766 121 767 125
rect 771 121 772 125
rect 766 120 772 121
rect 830 125 836 126
rect 830 121 831 125
rect 835 121 836 125
rect 830 120 836 121
rect 894 125 900 126
rect 894 121 895 125
rect 899 121 900 125
rect 894 120 900 121
rect 958 125 964 126
rect 958 121 959 125
rect 963 121 964 125
rect 958 120 964 121
rect 1022 125 1028 126
rect 1022 121 1023 125
rect 1027 121 1028 125
rect 1022 120 1028 121
rect 1086 125 1092 126
rect 1086 121 1087 125
rect 1091 121 1092 125
rect 1086 120 1092 121
rect 1150 125 1156 126
rect 1150 121 1151 125
rect 1155 121 1156 125
rect 1150 120 1156 121
rect 1286 124 1292 125
rect 1286 120 1287 124
rect 1291 120 1292 124
rect 110 119 116 120
rect 1286 119 1292 120
rect 1366 113 1372 114
rect 1326 112 1332 113
rect 1326 108 1327 112
rect 1331 108 1332 112
rect 1366 109 1367 113
rect 1371 109 1372 113
rect 1366 108 1372 109
rect 1422 113 1428 114
rect 1422 109 1423 113
rect 1427 109 1428 113
rect 1422 108 1428 109
rect 1478 113 1484 114
rect 1478 109 1479 113
rect 1483 109 1484 113
rect 1478 108 1484 109
rect 1534 113 1540 114
rect 1534 109 1535 113
rect 1539 109 1540 113
rect 1534 108 1540 109
rect 1590 113 1596 114
rect 1590 109 1591 113
rect 1595 109 1596 113
rect 1590 108 1596 109
rect 1646 113 1652 114
rect 1646 109 1647 113
rect 1651 109 1652 113
rect 1646 108 1652 109
rect 1702 113 1708 114
rect 1702 109 1703 113
rect 1707 109 1708 113
rect 1702 108 1708 109
rect 1758 113 1764 114
rect 1758 109 1759 113
rect 1763 109 1764 113
rect 1758 108 1764 109
rect 1822 113 1828 114
rect 1822 109 1823 113
rect 1827 109 1828 113
rect 1822 108 1828 109
rect 1878 113 1884 114
rect 1878 109 1879 113
rect 1883 109 1884 113
rect 1878 108 1884 109
rect 1942 113 1948 114
rect 1942 109 1943 113
rect 1947 109 1948 113
rect 1942 108 1948 109
rect 2006 113 2012 114
rect 2006 109 2007 113
rect 2011 109 2012 113
rect 2006 108 2012 109
rect 2070 113 2076 114
rect 2070 109 2071 113
rect 2075 109 2076 113
rect 2070 108 2076 109
rect 2142 113 2148 114
rect 2142 109 2143 113
rect 2147 109 2148 113
rect 2142 108 2148 109
rect 2222 113 2228 114
rect 2222 109 2223 113
rect 2227 109 2228 113
rect 2222 108 2228 109
rect 2302 113 2308 114
rect 2302 109 2303 113
rect 2307 109 2308 113
rect 2302 108 2308 109
rect 2390 113 2396 114
rect 2390 109 2391 113
rect 2395 109 2396 113
rect 2390 108 2396 109
rect 2454 113 2460 114
rect 2454 109 2455 113
rect 2459 109 2460 113
rect 2454 108 2460 109
rect 2502 112 2508 113
rect 2502 108 2503 112
rect 2507 108 2508 112
rect 110 107 116 108
rect 110 103 111 107
rect 115 103 116 107
rect 1286 107 1292 108
rect 1326 107 1332 108
rect 2502 107 2508 108
rect 110 102 116 103
rect 134 104 140 105
rect 134 100 135 104
rect 139 100 140 104
rect 134 99 140 100
rect 190 104 196 105
rect 190 100 191 104
rect 195 100 196 104
rect 190 99 196 100
rect 246 104 252 105
rect 246 100 247 104
rect 251 100 252 104
rect 246 99 252 100
rect 302 104 308 105
rect 302 100 303 104
rect 307 100 308 104
rect 302 99 308 100
rect 358 104 364 105
rect 358 100 359 104
rect 363 100 364 104
rect 358 99 364 100
rect 414 104 420 105
rect 414 100 415 104
rect 419 100 420 104
rect 414 99 420 100
rect 470 104 476 105
rect 470 100 471 104
rect 475 100 476 104
rect 470 99 476 100
rect 526 104 532 105
rect 526 100 527 104
rect 531 100 532 104
rect 526 99 532 100
rect 582 104 588 105
rect 582 100 583 104
rect 587 100 588 104
rect 582 99 588 100
rect 638 104 644 105
rect 638 100 639 104
rect 643 100 644 104
rect 638 99 644 100
rect 694 104 700 105
rect 694 100 695 104
rect 699 100 700 104
rect 694 99 700 100
rect 750 104 756 105
rect 750 100 751 104
rect 755 100 756 104
rect 750 99 756 100
rect 814 104 820 105
rect 814 100 815 104
rect 819 100 820 104
rect 814 99 820 100
rect 878 104 884 105
rect 878 100 879 104
rect 883 100 884 104
rect 878 99 884 100
rect 942 104 948 105
rect 942 100 943 104
rect 947 100 948 104
rect 942 99 948 100
rect 1006 104 1012 105
rect 1006 100 1007 104
rect 1011 100 1012 104
rect 1006 99 1012 100
rect 1070 104 1076 105
rect 1070 100 1071 104
rect 1075 100 1076 104
rect 1070 99 1076 100
rect 1134 104 1140 105
rect 1134 100 1135 104
rect 1139 100 1140 104
rect 1286 103 1287 107
rect 1291 103 1292 107
rect 1286 102 1292 103
rect 1134 99 1140 100
rect 1326 95 1332 96
rect 1326 91 1327 95
rect 1331 91 1332 95
rect 2502 95 2508 96
rect 1326 90 1332 91
rect 1350 92 1356 93
rect 1350 88 1351 92
rect 1355 88 1356 92
rect 1350 87 1356 88
rect 1406 92 1412 93
rect 1406 88 1407 92
rect 1411 88 1412 92
rect 1406 87 1412 88
rect 1462 92 1468 93
rect 1462 88 1463 92
rect 1467 88 1468 92
rect 1462 87 1468 88
rect 1518 92 1524 93
rect 1518 88 1519 92
rect 1523 88 1524 92
rect 1518 87 1524 88
rect 1574 92 1580 93
rect 1574 88 1575 92
rect 1579 88 1580 92
rect 1574 87 1580 88
rect 1630 92 1636 93
rect 1630 88 1631 92
rect 1635 88 1636 92
rect 1630 87 1636 88
rect 1686 92 1692 93
rect 1686 88 1687 92
rect 1691 88 1692 92
rect 1686 87 1692 88
rect 1742 92 1748 93
rect 1742 88 1743 92
rect 1747 88 1748 92
rect 1742 87 1748 88
rect 1806 92 1812 93
rect 1806 88 1807 92
rect 1811 88 1812 92
rect 1806 87 1812 88
rect 1862 92 1868 93
rect 1862 88 1863 92
rect 1867 88 1868 92
rect 1862 87 1868 88
rect 1926 92 1932 93
rect 1926 88 1927 92
rect 1931 88 1932 92
rect 1926 87 1932 88
rect 1990 92 1996 93
rect 1990 88 1991 92
rect 1995 88 1996 92
rect 1990 87 1996 88
rect 2054 92 2060 93
rect 2054 88 2055 92
rect 2059 88 2060 92
rect 2054 87 2060 88
rect 2126 92 2132 93
rect 2126 88 2127 92
rect 2131 88 2132 92
rect 2126 87 2132 88
rect 2206 92 2212 93
rect 2206 88 2207 92
rect 2211 88 2212 92
rect 2206 87 2212 88
rect 2286 92 2292 93
rect 2286 88 2287 92
rect 2291 88 2292 92
rect 2286 87 2292 88
rect 2374 92 2380 93
rect 2374 88 2375 92
rect 2379 88 2380 92
rect 2374 87 2380 88
rect 2438 92 2444 93
rect 2438 88 2439 92
rect 2443 88 2444 92
rect 2502 91 2503 95
rect 2507 91 2508 95
rect 2502 90 2508 91
rect 2438 87 2444 88
<< m3c >>
rect 111 2569 115 2573
rect 135 2572 139 2576
rect 191 2572 195 2576
rect 247 2572 251 2576
rect 303 2572 307 2576
rect 359 2572 363 2576
rect 1287 2569 1291 2573
rect 111 2552 115 2556
rect 151 2551 155 2555
rect 207 2551 211 2555
rect 263 2551 267 2555
rect 319 2551 323 2555
rect 375 2551 379 2555
rect 1287 2552 1291 2556
rect 1327 2549 1331 2553
rect 1495 2552 1499 2556
rect 1551 2552 1555 2556
rect 1607 2552 1611 2556
rect 1663 2552 1667 2556
rect 1719 2552 1723 2556
rect 1775 2552 1779 2556
rect 1831 2552 1835 2556
rect 1887 2552 1891 2556
rect 1943 2552 1947 2556
rect 1999 2552 2003 2556
rect 2055 2552 2059 2556
rect 2111 2552 2115 2556
rect 2167 2552 2171 2556
rect 2503 2549 2507 2553
rect 1327 2532 1331 2536
rect 1511 2531 1515 2535
rect 1567 2531 1571 2535
rect 1623 2531 1627 2535
rect 1679 2531 1683 2535
rect 1735 2531 1739 2535
rect 1791 2531 1795 2535
rect 1847 2531 1851 2535
rect 1903 2531 1907 2535
rect 1959 2531 1963 2535
rect 2015 2531 2019 2535
rect 2071 2531 2075 2535
rect 2127 2531 2131 2535
rect 2183 2531 2187 2535
rect 2503 2532 2507 2536
rect 111 2500 115 2504
rect 223 2501 227 2505
rect 279 2501 283 2505
rect 343 2501 347 2505
rect 415 2501 419 2505
rect 487 2501 491 2505
rect 551 2501 555 2505
rect 615 2501 619 2505
rect 679 2501 683 2505
rect 743 2501 747 2505
rect 807 2501 811 2505
rect 871 2501 875 2505
rect 935 2501 939 2505
rect 999 2501 1003 2505
rect 1063 2501 1067 2505
rect 1287 2500 1291 2504
rect 111 2483 115 2487
rect 207 2480 211 2484
rect 263 2480 267 2484
rect 327 2480 331 2484
rect 399 2480 403 2484
rect 471 2480 475 2484
rect 535 2480 539 2484
rect 599 2480 603 2484
rect 663 2480 667 2484
rect 727 2480 731 2484
rect 791 2480 795 2484
rect 855 2480 859 2484
rect 919 2480 923 2484
rect 983 2480 987 2484
rect 1047 2480 1051 2484
rect 1287 2483 1291 2487
rect 1327 2480 1331 2484
rect 1543 2481 1547 2485
rect 1607 2481 1611 2485
rect 1679 2481 1683 2485
rect 1751 2481 1755 2485
rect 1823 2481 1827 2485
rect 1895 2481 1899 2485
rect 1967 2481 1971 2485
rect 2039 2481 2043 2485
rect 2111 2481 2115 2485
rect 2183 2481 2187 2485
rect 2503 2480 2507 2484
rect 111 2457 115 2461
rect 167 2460 171 2464
rect 223 2460 227 2464
rect 279 2460 283 2464
rect 335 2460 339 2464
rect 391 2460 395 2464
rect 447 2460 451 2464
rect 503 2460 507 2464
rect 559 2460 563 2464
rect 615 2460 619 2464
rect 671 2460 675 2464
rect 727 2460 731 2464
rect 783 2460 787 2464
rect 839 2460 843 2464
rect 895 2460 899 2464
rect 951 2460 955 2464
rect 1007 2460 1011 2464
rect 1063 2460 1067 2464
rect 1327 2463 1331 2467
rect 1287 2457 1291 2461
rect 1527 2460 1531 2464
rect 1591 2460 1595 2464
rect 1663 2460 1667 2464
rect 1735 2460 1739 2464
rect 1807 2460 1811 2464
rect 1879 2460 1883 2464
rect 1951 2460 1955 2464
rect 2023 2460 2027 2464
rect 2095 2460 2099 2464
rect 2167 2460 2171 2464
rect 2503 2463 2507 2467
rect 111 2440 115 2444
rect 183 2439 187 2443
rect 239 2439 243 2443
rect 295 2439 299 2443
rect 351 2439 355 2443
rect 407 2439 411 2443
rect 463 2439 467 2443
rect 519 2439 523 2443
rect 575 2439 579 2443
rect 631 2439 635 2443
rect 687 2439 691 2443
rect 743 2439 747 2443
rect 799 2439 803 2443
rect 855 2439 859 2443
rect 911 2439 915 2443
rect 967 2439 971 2443
rect 1023 2439 1027 2443
rect 1079 2439 1083 2443
rect 1287 2440 1291 2444
rect 1327 2441 1331 2445
rect 1543 2444 1547 2448
rect 1607 2444 1611 2448
rect 1671 2444 1675 2448
rect 1743 2444 1747 2448
rect 1815 2444 1819 2448
rect 1879 2444 1883 2448
rect 1951 2444 1955 2448
rect 2023 2444 2027 2448
rect 2095 2444 2099 2448
rect 2167 2444 2171 2448
rect 2503 2441 2507 2445
rect 1327 2424 1331 2428
rect 1559 2423 1563 2427
rect 1623 2423 1627 2427
rect 1687 2423 1691 2427
rect 1759 2423 1763 2427
rect 1831 2423 1835 2427
rect 1895 2423 1899 2427
rect 1967 2423 1971 2427
rect 2039 2423 2043 2427
rect 2111 2423 2115 2427
rect 2183 2423 2187 2427
rect 2503 2424 2507 2428
rect 111 2376 115 2380
rect 519 2377 523 2381
rect 575 2377 579 2381
rect 631 2377 635 2381
rect 687 2377 691 2381
rect 1287 2376 1291 2380
rect 1327 2368 1331 2372
rect 1567 2369 1571 2373
rect 1623 2369 1627 2373
rect 1679 2369 1683 2373
rect 1735 2369 1739 2373
rect 1791 2369 1795 2373
rect 1855 2369 1859 2373
rect 1919 2369 1923 2373
rect 1983 2369 1987 2373
rect 2047 2369 2051 2373
rect 2111 2369 2115 2373
rect 2503 2368 2507 2372
rect 111 2359 115 2363
rect 503 2356 507 2360
rect 559 2356 563 2360
rect 615 2356 619 2360
rect 671 2356 675 2360
rect 1287 2359 1291 2363
rect 1327 2351 1331 2355
rect 1551 2348 1555 2352
rect 1607 2348 1611 2352
rect 1663 2348 1667 2352
rect 1719 2348 1723 2352
rect 1775 2348 1779 2352
rect 1839 2348 1843 2352
rect 1903 2348 1907 2352
rect 1967 2348 1971 2352
rect 2031 2348 2035 2352
rect 2095 2348 2099 2352
rect 2503 2351 2507 2355
rect 111 2333 115 2337
rect 319 2336 323 2340
rect 391 2336 395 2340
rect 463 2336 467 2340
rect 535 2336 539 2340
rect 607 2336 611 2340
rect 679 2336 683 2340
rect 743 2336 747 2340
rect 807 2336 811 2340
rect 863 2336 867 2340
rect 927 2336 931 2340
rect 991 2336 995 2340
rect 1055 2336 1059 2340
rect 1111 2336 1115 2340
rect 1167 2336 1171 2340
rect 1223 2336 1227 2340
rect 1287 2333 1291 2337
rect 1327 2325 1331 2329
rect 1471 2328 1475 2332
rect 1535 2328 1539 2332
rect 1607 2328 1611 2332
rect 1687 2328 1691 2332
rect 1759 2328 1763 2332
rect 1831 2328 1835 2332
rect 1903 2328 1907 2332
rect 1983 2328 1987 2332
rect 2063 2328 2067 2332
rect 2143 2328 2147 2332
rect 2503 2325 2507 2329
rect 111 2316 115 2320
rect 335 2315 339 2319
rect 407 2315 411 2319
rect 479 2315 483 2319
rect 551 2315 555 2319
rect 623 2315 627 2319
rect 695 2315 699 2319
rect 759 2315 763 2319
rect 823 2315 827 2319
rect 879 2315 883 2319
rect 943 2315 947 2319
rect 1007 2315 1011 2319
rect 1071 2315 1075 2319
rect 1127 2315 1131 2319
rect 1183 2315 1187 2319
rect 1239 2315 1243 2319
rect 1287 2316 1291 2320
rect 1327 2308 1331 2312
rect 1487 2307 1491 2311
rect 1551 2307 1555 2311
rect 1623 2307 1627 2311
rect 1703 2307 1707 2311
rect 1775 2307 1779 2311
rect 1847 2307 1851 2311
rect 1919 2307 1923 2311
rect 1999 2307 2003 2311
rect 2079 2307 2083 2311
rect 2159 2307 2163 2311
rect 2503 2308 2507 2312
rect 111 2256 115 2260
rect 175 2257 179 2261
rect 271 2257 275 2261
rect 375 2257 379 2261
rect 479 2257 483 2261
rect 591 2257 595 2261
rect 703 2257 707 2261
rect 807 2257 811 2261
rect 911 2257 915 2261
rect 1015 2257 1019 2261
rect 1127 2257 1131 2261
rect 1239 2257 1243 2261
rect 1287 2256 1291 2260
rect 1327 2256 1331 2260
rect 1383 2257 1387 2261
rect 1479 2257 1483 2261
rect 1583 2257 1587 2261
rect 1687 2257 1691 2261
rect 1791 2257 1795 2261
rect 1903 2257 1907 2261
rect 2015 2257 2019 2261
rect 2127 2257 2131 2261
rect 2239 2257 2243 2261
rect 2503 2256 2507 2260
rect 111 2239 115 2243
rect 159 2236 163 2240
rect 255 2236 259 2240
rect 359 2236 363 2240
rect 463 2236 467 2240
rect 575 2236 579 2240
rect 687 2236 691 2240
rect 791 2236 795 2240
rect 895 2236 899 2240
rect 999 2236 1003 2240
rect 1111 2236 1115 2240
rect 1223 2236 1227 2240
rect 1287 2239 1291 2243
rect 1327 2239 1331 2243
rect 1367 2236 1371 2240
rect 1463 2236 1467 2240
rect 1567 2236 1571 2240
rect 1671 2236 1675 2240
rect 1775 2236 1779 2240
rect 1887 2236 1891 2240
rect 1999 2236 2003 2240
rect 2111 2236 2115 2240
rect 2223 2236 2227 2240
rect 2503 2239 2507 2243
rect 111 2221 115 2225
rect 143 2224 147 2228
rect 231 2224 235 2228
rect 319 2224 323 2228
rect 415 2224 419 2228
rect 519 2224 523 2228
rect 623 2224 627 2228
rect 727 2224 731 2228
rect 831 2224 835 2228
rect 935 2224 939 2228
rect 1039 2224 1043 2228
rect 1143 2224 1147 2228
rect 1223 2224 1227 2228
rect 1287 2221 1291 2225
rect 1327 2221 1331 2225
rect 1367 2224 1371 2228
rect 1487 2224 1491 2228
rect 1607 2224 1611 2228
rect 1719 2224 1723 2228
rect 1815 2224 1819 2228
rect 1903 2224 1907 2228
rect 1983 2224 1987 2228
rect 2055 2224 2059 2228
rect 2127 2224 2131 2228
rect 2191 2224 2195 2228
rect 2255 2224 2259 2228
rect 2319 2224 2323 2228
rect 2383 2224 2387 2228
rect 2439 2224 2443 2228
rect 2503 2221 2507 2225
rect 111 2204 115 2208
rect 159 2203 163 2207
rect 247 2203 251 2207
rect 335 2203 339 2207
rect 431 2203 435 2207
rect 535 2203 539 2207
rect 639 2203 643 2207
rect 743 2203 747 2207
rect 847 2203 851 2207
rect 951 2203 955 2207
rect 1055 2203 1059 2207
rect 1159 2203 1163 2207
rect 1239 2203 1243 2207
rect 1287 2204 1291 2208
rect 1327 2204 1331 2208
rect 1383 2203 1387 2207
rect 1503 2203 1507 2207
rect 1623 2203 1627 2207
rect 1735 2203 1739 2207
rect 1831 2203 1835 2207
rect 1919 2203 1923 2207
rect 1999 2203 2003 2207
rect 2071 2203 2075 2207
rect 2143 2203 2147 2207
rect 2207 2203 2211 2207
rect 2271 2203 2275 2207
rect 2335 2203 2339 2207
rect 2399 2203 2403 2207
rect 2455 2203 2459 2207
rect 2503 2204 2507 2208
rect 111 2152 115 2156
rect 255 2153 259 2157
rect 351 2153 355 2157
rect 455 2153 459 2157
rect 559 2153 563 2157
rect 663 2153 667 2157
rect 767 2153 771 2157
rect 863 2153 867 2157
rect 959 2153 963 2157
rect 1055 2153 1059 2157
rect 1159 2153 1163 2157
rect 1239 2153 1243 2157
rect 1287 2152 1291 2156
rect 111 2135 115 2139
rect 239 2132 243 2136
rect 335 2132 339 2136
rect 439 2132 443 2136
rect 543 2132 547 2136
rect 647 2132 651 2136
rect 751 2132 755 2136
rect 847 2132 851 2136
rect 943 2132 947 2136
rect 1039 2132 1043 2136
rect 1143 2132 1147 2136
rect 1223 2132 1227 2136
rect 1287 2135 1291 2139
rect 1327 2132 1331 2136
rect 1407 2133 1411 2137
rect 1623 2133 1627 2137
rect 1815 2133 1819 2137
rect 1991 2133 1995 2137
rect 2159 2133 2163 2137
rect 2319 2133 2323 2137
rect 2455 2133 2459 2137
rect 2503 2132 2507 2136
rect 111 2117 115 2121
rect 303 2120 307 2124
rect 359 2120 363 2124
rect 423 2120 427 2124
rect 487 2120 491 2124
rect 559 2120 563 2124
rect 631 2120 635 2124
rect 711 2120 715 2124
rect 799 2120 803 2124
rect 887 2120 891 2124
rect 975 2120 979 2124
rect 1063 2120 1067 2124
rect 1151 2120 1155 2124
rect 1223 2120 1227 2124
rect 1287 2117 1291 2121
rect 1327 2115 1331 2119
rect 1391 2112 1395 2116
rect 1607 2112 1611 2116
rect 1799 2112 1803 2116
rect 1975 2112 1979 2116
rect 2143 2112 2147 2116
rect 2303 2112 2307 2116
rect 2439 2112 2443 2116
rect 2503 2115 2507 2119
rect 111 2100 115 2104
rect 319 2099 323 2103
rect 375 2099 379 2103
rect 439 2099 443 2103
rect 503 2099 507 2103
rect 575 2099 579 2103
rect 647 2099 651 2103
rect 727 2099 731 2103
rect 815 2099 819 2103
rect 903 2099 907 2103
rect 991 2099 995 2103
rect 1079 2099 1083 2103
rect 1167 2099 1171 2103
rect 1239 2099 1243 2103
rect 1287 2100 1291 2104
rect 1327 2097 1331 2101
rect 1383 2100 1387 2104
rect 1551 2100 1555 2104
rect 1711 2100 1715 2104
rect 1855 2100 1859 2104
rect 1991 2100 1995 2104
rect 2119 2100 2123 2104
rect 2239 2100 2243 2104
rect 2367 2100 2371 2104
rect 2503 2097 2507 2101
rect 1327 2080 1331 2084
rect 1399 2079 1403 2083
rect 1567 2079 1571 2083
rect 1727 2079 1731 2083
rect 1871 2079 1875 2083
rect 2007 2079 2011 2083
rect 2135 2079 2139 2083
rect 2255 2079 2259 2083
rect 2383 2079 2387 2083
rect 2503 2080 2507 2084
rect 111 2044 115 2048
rect 399 2045 403 2049
rect 455 2045 459 2049
rect 511 2045 515 2049
rect 575 2045 579 2049
rect 639 2045 643 2049
rect 711 2045 715 2049
rect 791 2045 795 2049
rect 863 2045 867 2049
rect 943 2045 947 2049
rect 1023 2045 1027 2049
rect 1103 2045 1107 2049
rect 1183 2045 1187 2049
rect 1239 2045 1243 2049
rect 1287 2044 1291 2048
rect 111 2027 115 2031
rect 383 2024 387 2028
rect 439 2024 443 2028
rect 495 2024 499 2028
rect 559 2024 563 2028
rect 623 2024 627 2028
rect 695 2024 699 2028
rect 775 2024 779 2028
rect 847 2024 851 2028
rect 927 2024 931 2028
rect 1007 2024 1011 2028
rect 1087 2024 1091 2028
rect 1167 2024 1171 2028
rect 1223 2024 1227 2028
rect 1287 2027 1291 2031
rect 1327 2024 1331 2028
rect 1447 2025 1451 2029
rect 1551 2025 1555 2029
rect 1655 2025 1659 2029
rect 1751 2025 1755 2029
rect 1839 2025 1843 2029
rect 1927 2025 1931 2029
rect 2023 2025 2027 2029
rect 2119 2025 2123 2029
rect 2503 2024 2507 2028
rect 111 2005 115 2009
rect 231 2008 235 2012
rect 287 2008 291 2012
rect 359 2008 363 2012
rect 439 2008 443 2012
rect 535 2008 539 2012
rect 631 2008 635 2012
rect 735 2008 739 2012
rect 847 2008 851 2012
rect 959 2008 963 2012
rect 1079 2008 1083 2012
rect 1199 2008 1203 2012
rect 1287 2005 1291 2009
rect 1327 2007 1331 2011
rect 1431 2004 1435 2008
rect 1535 2004 1539 2008
rect 1639 2004 1643 2008
rect 1735 2004 1739 2008
rect 1823 2004 1827 2008
rect 1911 2004 1915 2008
rect 2007 2004 2011 2008
rect 2103 2004 2107 2008
rect 2503 2007 2507 2011
rect 111 1988 115 1992
rect 247 1987 251 1991
rect 303 1987 307 1991
rect 375 1987 379 1991
rect 455 1987 459 1991
rect 551 1987 555 1991
rect 647 1987 651 1991
rect 751 1987 755 1991
rect 863 1987 867 1991
rect 975 1987 979 1991
rect 1095 1987 1099 1991
rect 1215 1987 1219 1991
rect 1287 1988 1291 1992
rect 1327 1985 1331 1989
rect 1455 1988 1459 1992
rect 1511 1988 1515 1992
rect 1575 1988 1579 1992
rect 1639 1988 1643 1992
rect 1703 1988 1707 1992
rect 1767 1988 1771 1992
rect 1831 1988 1835 1992
rect 1895 1988 1899 1992
rect 1959 1988 1963 1992
rect 2031 1988 2035 1992
rect 2503 1985 2507 1989
rect 1327 1968 1331 1972
rect 1471 1967 1475 1971
rect 1527 1967 1531 1971
rect 1591 1967 1595 1971
rect 1655 1967 1659 1971
rect 1719 1967 1723 1971
rect 1783 1967 1787 1971
rect 1847 1967 1851 1971
rect 1911 1967 1915 1971
rect 1975 1967 1979 1971
rect 2047 1967 2051 1971
rect 2503 1968 2507 1972
rect 111 1932 115 1936
rect 151 1933 155 1937
rect 215 1933 219 1937
rect 319 1933 323 1937
rect 439 1933 443 1937
rect 583 1933 587 1937
rect 743 1933 747 1937
rect 919 1933 923 1937
rect 1095 1933 1099 1937
rect 1287 1932 1291 1936
rect 111 1915 115 1919
rect 135 1912 139 1916
rect 199 1912 203 1916
rect 303 1912 307 1916
rect 423 1912 427 1916
rect 567 1912 571 1916
rect 727 1912 731 1916
rect 903 1912 907 1916
rect 1079 1912 1083 1916
rect 1287 1915 1291 1919
rect 1327 1912 1331 1916
rect 1567 1913 1571 1917
rect 1631 1913 1635 1917
rect 1703 1913 1707 1917
rect 1775 1913 1779 1917
rect 1847 1913 1851 1917
rect 1919 1913 1923 1917
rect 1999 1913 2003 1917
rect 2087 1913 2091 1917
rect 2183 1913 2187 1917
rect 2279 1913 2283 1917
rect 2375 1913 2379 1917
rect 2455 1913 2459 1917
rect 2503 1912 2507 1916
rect 111 1889 115 1893
rect 135 1892 139 1896
rect 191 1892 195 1896
rect 271 1892 275 1896
rect 359 1892 363 1896
rect 455 1892 459 1896
rect 543 1892 547 1896
rect 631 1892 635 1896
rect 719 1892 723 1896
rect 799 1892 803 1896
rect 871 1892 875 1896
rect 943 1892 947 1896
rect 1015 1892 1019 1896
rect 1087 1892 1091 1896
rect 1159 1892 1163 1896
rect 1327 1895 1331 1899
rect 1287 1889 1291 1893
rect 1551 1892 1555 1896
rect 1615 1892 1619 1896
rect 1687 1892 1691 1896
rect 1759 1892 1763 1896
rect 1831 1892 1835 1896
rect 1903 1892 1907 1896
rect 1983 1892 1987 1896
rect 2071 1892 2075 1896
rect 2167 1892 2171 1896
rect 2263 1892 2267 1896
rect 2359 1892 2363 1896
rect 2439 1892 2443 1896
rect 2503 1895 2507 1899
rect 111 1872 115 1876
rect 151 1871 155 1875
rect 207 1871 211 1875
rect 287 1871 291 1875
rect 375 1871 379 1875
rect 471 1871 475 1875
rect 559 1871 563 1875
rect 647 1871 651 1875
rect 735 1871 739 1875
rect 815 1871 819 1875
rect 887 1871 891 1875
rect 959 1871 963 1875
rect 1031 1871 1035 1875
rect 1103 1871 1107 1875
rect 1175 1871 1179 1875
rect 1287 1872 1291 1876
rect 1327 1873 1331 1877
rect 1607 1876 1611 1880
rect 1663 1876 1667 1880
rect 1727 1876 1731 1880
rect 1799 1876 1803 1880
rect 1871 1876 1875 1880
rect 1943 1876 1947 1880
rect 2007 1876 2011 1880
rect 2071 1876 2075 1880
rect 2135 1876 2139 1880
rect 2199 1876 2203 1880
rect 2263 1876 2267 1880
rect 2327 1876 2331 1880
rect 2383 1876 2387 1880
rect 2439 1876 2443 1880
rect 2503 1873 2507 1877
rect 1327 1856 1331 1860
rect 1623 1855 1627 1859
rect 1679 1855 1683 1859
rect 1743 1855 1747 1859
rect 1815 1855 1819 1859
rect 1887 1855 1891 1859
rect 1959 1855 1963 1859
rect 2023 1855 2027 1859
rect 2087 1855 2091 1859
rect 2151 1855 2155 1859
rect 2215 1855 2219 1859
rect 2279 1855 2283 1859
rect 2343 1855 2347 1859
rect 2399 1855 2403 1859
rect 2455 1855 2459 1859
rect 2503 1856 2507 1860
rect 111 1820 115 1824
rect 151 1821 155 1825
rect 207 1821 211 1825
rect 295 1821 299 1825
rect 391 1821 395 1825
rect 495 1821 499 1825
rect 591 1821 595 1825
rect 687 1821 691 1825
rect 775 1821 779 1825
rect 855 1821 859 1825
rect 927 1821 931 1825
rect 999 1821 1003 1825
rect 1079 1821 1083 1825
rect 1159 1821 1163 1825
rect 1287 1820 1291 1824
rect 111 1803 115 1807
rect 135 1800 139 1804
rect 191 1800 195 1804
rect 279 1800 283 1804
rect 375 1800 379 1804
rect 479 1800 483 1804
rect 575 1800 579 1804
rect 671 1800 675 1804
rect 759 1800 763 1804
rect 839 1800 843 1804
rect 911 1800 915 1804
rect 983 1800 987 1804
rect 1063 1800 1067 1804
rect 1143 1800 1147 1804
rect 1287 1803 1291 1807
rect 1327 1800 1331 1804
rect 1631 1801 1635 1805
rect 1719 1801 1723 1805
rect 1815 1801 1819 1805
rect 1927 1801 1931 1805
rect 2055 1801 2059 1805
rect 2191 1801 2195 1805
rect 2335 1801 2339 1805
rect 2455 1801 2459 1805
rect 2503 1800 2507 1804
rect 1327 1783 1331 1787
rect 111 1773 115 1777
rect 135 1776 139 1780
rect 199 1776 203 1780
rect 295 1776 299 1780
rect 399 1776 403 1780
rect 503 1776 507 1780
rect 607 1776 611 1780
rect 703 1776 707 1780
rect 799 1776 803 1780
rect 887 1776 891 1780
rect 975 1776 979 1780
rect 1063 1776 1067 1780
rect 1151 1776 1155 1780
rect 1615 1780 1619 1784
rect 1703 1780 1707 1784
rect 1799 1780 1803 1784
rect 1911 1780 1915 1784
rect 2039 1780 2043 1784
rect 2175 1780 2179 1784
rect 2319 1780 2323 1784
rect 2439 1780 2443 1784
rect 2503 1783 2507 1787
rect 1287 1773 1291 1777
rect 1327 1765 1331 1769
rect 1527 1768 1531 1772
rect 1607 1768 1611 1772
rect 1695 1768 1699 1772
rect 1791 1768 1795 1772
rect 1879 1768 1883 1772
rect 1967 1768 1971 1772
rect 2055 1768 2059 1772
rect 2135 1768 2139 1772
rect 2215 1768 2219 1772
rect 2295 1768 2299 1772
rect 2375 1768 2379 1772
rect 2439 1768 2443 1772
rect 2503 1765 2507 1769
rect 111 1756 115 1760
rect 151 1755 155 1759
rect 215 1755 219 1759
rect 311 1755 315 1759
rect 415 1755 419 1759
rect 519 1755 523 1759
rect 623 1755 627 1759
rect 719 1755 723 1759
rect 815 1755 819 1759
rect 903 1755 907 1759
rect 991 1755 995 1759
rect 1079 1755 1083 1759
rect 1167 1755 1171 1759
rect 1287 1756 1291 1760
rect 1327 1748 1331 1752
rect 1543 1747 1547 1751
rect 1623 1747 1627 1751
rect 1711 1747 1715 1751
rect 1807 1747 1811 1751
rect 1895 1747 1899 1751
rect 1983 1747 1987 1751
rect 2071 1747 2075 1751
rect 2151 1747 2155 1751
rect 2231 1747 2235 1751
rect 2311 1747 2315 1751
rect 2391 1747 2395 1751
rect 2455 1747 2459 1751
rect 2503 1748 2507 1752
rect 111 1700 115 1704
rect 167 1701 171 1705
rect 239 1701 243 1705
rect 319 1701 323 1705
rect 407 1701 411 1705
rect 503 1701 507 1705
rect 607 1701 611 1705
rect 711 1701 715 1705
rect 823 1701 827 1705
rect 935 1701 939 1705
rect 1047 1701 1051 1705
rect 1159 1701 1163 1705
rect 1287 1700 1291 1704
rect 1327 1692 1331 1696
rect 1399 1693 1403 1697
rect 1463 1693 1467 1697
rect 1543 1693 1547 1697
rect 1631 1693 1635 1697
rect 1727 1693 1731 1697
rect 1823 1693 1827 1697
rect 1919 1693 1923 1697
rect 2015 1693 2019 1697
rect 2111 1693 2115 1697
rect 2199 1693 2203 1697
rect 2287 1693 2291 1697
rect 2383 1693 2387 1697
rect 2455 1693 2459 1697
rect 2503 1692 2507 1696
rect 111 1683 115 1687
rect 151 1680 155 1684
rect 223 1680 227 1684
rect 303 1680 307 1684
rect 391 1680 395 1684
rect 487 1680 491 1684
rect 591 1680 595 1684
rect 695 1680 699 1684
rect 807 1680 811 1684
rect 919 1680 923 1684
rect 1031 1680 1035 1684
rect 1143 1680 1147 1684
rect 1287 1683 1291 1687
rect 1327 1675 1331 1679
rect 1383 1672 1387 1676
rect 1447 1672 1451 1676
rect 1527 1672 1531 1676
rect 1615 1672 1619 1676
rect 1711 1672 1715 1676
rect 1807 1672 1811 1676
rect 1903 1672 1907 1676
rect 1999 1672 2003 1676
rect 2095 1672 2099 1676
rect 2183 1672 2187 1676
rect 2271 1672 2275 1676
rect 2367 1672 2371 1676
rect 2439 1672 2443 1676
rect 2503 1675 2507 1679
rect 111 1661 115 1665
rect 255 1664 259 1668
rect 319 1664 323 1668
rect 399 1664 403 1668
rect 487 1664 491 1668
rect 575 1664 579 1668
rect 671 1664 675 1668
rect 767 1664 771 1668
rect 863 1664 867 1668
rect 959 1664 963 1668
rect 1063 1664 1067 1668
rect 1167 1664 1171 1668
rect 1287 1661 1291 1665
rect 1327 1653 1331 1657
rect 1351 1656 1355 1660
rect 1407 1656 1411 1660
rect 1495 1656 1499 1660
rect 1583 1656 1587 1660
rect 1679 1656 1683 1660
rect 1783 1656 1787 1660
rect 1895 1656 1899 1660
rect 2023 1656 2027 1660
rect 2159 1656 2163 1660
rect 2303 1656 2307 1660
rect 2439 1656 2443 1660
rect 2503 1653 2507 1657
rect 111 1644 115 1648
rect 271 1643 275 1647
rect 335 1643 339 1647
rect 415 1643 419 1647
rect 503 1643 507 1647
rect 591 1643 595 1647
rect 687 1643 691 1647
rect 783 1643 787 1647
rect 879 1643 883 1647
rect 975 1643 979 1647
rect 1079 1643 1083 1647
rect 1183 1643 1187 1647
rect 1287 1644 1291 1648
rect 1327 1636 1331 1640
rect 1367 1635 1371 1639
rect 1423 1635 1427 1639
rect 1511 1635 1515 1639
rect 1599 1635 1603 1639
rect 1695 1635 1699 1639
rect 1799 1635 1803 1639
rect 1911 1635 1915 1639
rect 2039 1635 2043 1639
rect 2175 1635 2179 1639
rect 2319 1635 2323 1639
rect 2455 1635 2459 1639
rect 2503 1636 2507 1640
rect 111 1588 115 1592
rect 303 1589 307 1593
rect 359 1589 363 1593
rect 431 1589 435 1593
rect 511 1589 515 1593
rect 599 1589 603 1593
rect 695 1589 699 1593
rect 791 1589 795 1593
rect 895 1589 899 1593
rect 1007 1589 1011 1593
rect 1119 1589 1123 1593
rect 1287 1588 1291 1592
rect 1327 1584 1331 1588
rect 1367 1585 1371 1589
rect 1423 1585 1427 1589
rect 1479 1585 1483 1589
rect 1559 1585 1563 1589
rect 1639 1585 1643 1589
rect 1719 1585 1723 1589
rect 1791 1585 1795 1589
rect 1871 1585 1875 1589
rect 1951 1585 1955 1589
rect 2031 1585 2035 1589
rect 2503 1584 2507 1588
rect 111 1571 115 1575
rect 287 1568 291 1572
rect 343 1568 347 1572
rect 415 1568 419 1572
rect 495 1568 499 1572
rect 583 1568 587 1572
rect 679 1568 683 1572
rect 775 1568 779 1572
rect 879 1568 883 1572
rect 991 1568 995 1572
rect 1103 1568 1107 1572
rect 1287 1571 1291 1575
rect 1327 1567 1331 1571
rect 1351 1564 1355 1568
rect 1407 1564 1411 1568
rect 1463 1564 1467 1568
rect 1543 1564 1547 1568
rect 1623 1564 1627 1568
rect 1703 1564 1707 1568
rect 1775 1564 1779 1568
rect 1855 1564 1859 1568
rect 1935 1564 1939 1568
rect 2015 1564 2019 1568
rect 2503 1567 2507 1571
rect 111 1553 115 1557
rect 247 1556 251 1560
rect 319 1556 323 1560
rect 399 1556 403 1560
rect 487 1556 491 1560
rect 583 1556 587 1560
rect 671 1556 675 1560
rect 759 1556 763 1560
rect 847 1556 851 1560
rect 927 1556 931 1560
rect 1007 1556 1011 1560
rect 1087 1556 1091 1560
rect 1167 1556 1171 1560
rect 1223 1556 1227 1560
rect 1287 1553 1291 1557
rect 1327 1549 1331 1553
rect 1351 1552 1355 1556
rect 1471 1552 1475 1556
rect 1607 1552 1611 1556
rect 1735 1552 1739 1556
rect 1871 1552 1875 1556
rect 2007 1552 2011 1556
rect 2503 1549 2507 1553
rect 111 1536 115 1540
rect 263 1535 267 1539
rect 335 1535 339 1539
rect 415 1535 419 1539
rect 503 1535 507 1539
rect 599 1535 603 1539
rect 687 1535 691 1539
rect 775 1535 779 1539
rect 863 1535 867 1539
rect 943 1535 947 1539
rect 1023 1535 1027 1539
rect 1103 1535 1107 1539
rect 1183 1535 1187 1539
rect 1239 1535 1243 1539
rect 1287 1536 1291 1540
rect 1327 1532 1331 1536
rect 1367 1531 1371 1535
rect 1487 1531 1491 1535
rect 1623 1531 1627 1535
rect 1751 1531 1755 1535
rect 1887 1531 1891 1535
rect 2023 1531 2027 1535
rect 2503 1532 2507 1536
rect 111 1476 115 1480
rect 279 1477 283 1481
rect 343 1477 347 1481
rect 415 1477 419 1481
rect 495 1477 499 1481
rect 575 1477 579 1481
rect 655 1477 659 1481
rect 735 1477 739 1481
rect 815 1477 819 1481
rect 895 1477 899 1481
rect 975 1477 979 1481
rect 1055 1477 1059 1481
rect 1143 1477 1147 1481
rect 1287 1476 1291 1480
rect 1327 1480 1331 1484
rect 1367 1481 1371 1485
rect 1423 1481 1427 1485
rect 1479 1481 1483 1485
rect 1551 1481 1555 1485
rect 1631 1481 1635 1485
rect 1711 1481 1715 1485
rect 1791 1481 1795 1485
rect 1871 1481 1875 1485
rect 1951 1481 1955 1485
rect 2031 1481 2035 1485
rect 2119 1481 2123 1485
rect 2503 1480 2507 1484
rect 111 1459 115 1463
rect 263 1456 267 1460
rect 327 1456 331 1460
rect 399 1456 403 1460
rect 479 1456 483 1460
rect 559 1456 563 1460
rect 639 1456 643 1460
rect 719 1456 723 1460
rect 799 1456 803 1460
rect 879 1456 883 1460
rect 959 1456 963 1460
rect 1039 1456 1043 1460
rect 1127 1456 1131 1460
rect 1287 1459 1291 1463
rect 1327 1463 1331 1467
rect 1351 1460 1355 1464
rect 1407 1460 1411 1464
rect 1463 1460 1467 1464
rect 1535 1460 1539 1464
rect 1615 1460 1619 1464
rect 1695 1460 1699 1464
rect 1775 1460 1779 1464
rect 1855 1460 1859 1464
rect 1935 1460 1939 1464
rect 2015 1460 2019 1464
rect 2103 1460 2107 1464
rect 2503 1463 2507 1467
rect 111 1437 115 1441
rect 191 1440 195 1444
rect 255 1440 259 1444
rect 327 1440 331 1444
rect 407 1440 411 1444
rect 503 1440 507 1444
rect 607 1440 611 1444
rect 711 1440 715 1444
rect 815 1440 819 1444
rect 919 1440 923 1444
rect 1023 1440 1027 1444
rect 1127 1440 1131 1444
rect 1223 1440 1227 1444
rect 1287 1437 1291 1441
rect 1327 1437 1331 1441
rect 1359 1440 1363 1444
rect 1447 1440 1451 1444
rect 1535 1440 1539 1444
rect 1631 1440 1635 1444
rect 1727 1440 1731 1444
rect 1815 1440 1819 1444
rect 1903 1440 1907 1444
rect 1991 1440 1995 1444
rect 2071 1440 2075 1444
rect 2159 1440 2163 1444
rect 2247 1440 2251 1444
rect 2503 1437 2507 1441
rect 111 1420 115 1424
rect 207 1419 211 1423
rect 271 1419 275 1423
rect 343 1419 347 1423
rect 423 1419 427 1423
rect 519 1419 523 1423
rect 623 1419 627 1423
rect 727 1419 731 1423
rect 831 1419 835 1423
rect 935 1419 939 1423
rect 1039 1419 1043 1423
rect 1143 1419 1147 1423
rect 1239 1419 1243 1423
rect 1287 1420 1291 1424
rect 1327 1420 1331 1424
rect 1375 1419 1379 1423
rect 1463 1419 1467 1423
rect 1551 1419 1555 1423
rect 1647 1419 1651 1423
rect 1743 1419 1747 1423
rect 1831 1419 1835 1423
rect 1919 1419 1923 1423
rect 2007 1419 2011 1423
rect 2087 1419 2091 1423
rect 2175 1419 2179 1423
rect 2263 1419 2267 1423
rect 2503 1420 2507 1424
rect 111 1364 115 1368
rect 151 1365 155 1369
rect 223 1365 227 1369
rect 295 1365 299 1369
rect 359 1365 363 1369
rect 431 1365 435 1369
rect 503 1365 507 1369
rect 583 1365 587 1369
rect 663 1365 667 1369
rect 751 1365 755 1369
rect 839 1365 843 1369
rect 927 1365 931 1369
rect 1015 1365 1019 1369
rect 1103 1365 1107 1369
rect 1199 1365 1203 1369
rect 1287 1364 1291 1368
rect 1327 1368 1331 1372
rect 1567 1369 1571 1373
rect 1647 1369 1651 1373
rect 1735 1369 1739 1373
rect 1831 1369 1835 1373
rect 1919 1369 1923 1373
rect 2007 1369 2011 1373
rect 2095 1369 2099 1373
rect 2175 1369 2179 1373
rect 2247 1369 2251 1373
rect 2319 1369 2323 1373
rect 2399 1369 2403 1373
rect 2455 1369 2459 1373
rect 2503 1368 2507 1372
rect 111 1347 115 1351
rect 135 1344 139 1348
rect 207 1344 211 1348
rect 279 1344 283 1348
rect 343 1344 347 1348
rect 415 1344 419 1348
rect 487 1344 491 1348
rect 567 1344 571 1348
rect 647 1344 651 1348
rect 735 1344 739 1348
rect 823 1344 827 1348
rect 911 1344 915 1348
rect 999 1344 1003 1348
rect 1087 1344 1091 1348
rect 1183 1344 1187 1348
rect 1287 1347 1291 1351
rect 1327 1351 1331 1355
rect 1551 1348 1555 1352
rect 1631 1348 1635 1352
rect 1719 1348 1723 1352
rect 1815 1348 1819 1352
rect 1903 1348 1907 1352
rect 1991 1348 1995 1352
rect 2079 1348 2083 1352
rect 2159 1348 2163 1352
rect 2231 1348 2235 1352
rect 2303 1348 2307 1352
rect 2383 1348 2387 1352
rect 2439 1348 2443 1352
rect 2503 1351 2507 1355
rect 1327 1333 1331 1337
rect 1583 1336 1587 1340
rect 1647 1336 1651 1340
rect 1727 1336 1731 1340
rect 1807 1336 1811 1340
rect 1895 1336 1899 1340
rect 1983 1336 1987 1340
rect 2063 1336 2067 1340
rect 2143 1336 2147 1340
rect 2223 1336 2227 1340
rect 2303 1336 2307 1340
rect 2383 1336 2387 1340
rect 2439 1336 2443 1340
rect 2503 1333 2507 1337
rect 111 1313 115 1317
rect 135 1316 139 1320
rect 239 1316 243 1320
rect 367 1316 371 1320
rect 479 1316 483 1320
rect 583 1316 587 1320
rect 687 1316 691 1320
rect 783 1316 787 1320
rect 879 1316 883 1320
rect 975 1316 979 1320
rect 1287 1313 1291 1317
rect 1327 1316 1331 1320
rect 1599 1315 1603 1319
rect 1663 1315 1667 1319
rect 1743 1315 1747 1319
rect 1823 1315 1827 1319
rect 1911 1315 1915 1319
rect 1999 1315 2003 1319
rect 2079 1315 2083 1319
rect 2159 1315 2163 1319
rect 2239 1315 2243 1319
rect 2319 1315 2323 1319
rect 2399 1315 2403 1319
rect 2455 1315 2459 1319
rect 2503 1316 2507 1320
rect 111 1296 115 1300
rect 151 1295 155 1299
rect 255 1295 259 1299
rect 383 1295 387 1299
rect 495 1295 499 1299
rect 599 1295 603 1299
rect 703 1295 707 1299
rect 799 1295 803 1299
rect 895 1295 899 1299
rect 991 1295 995 1299
rect 1287 1296 1291 1300
rect 1327 1264 1331 1268
rect 1567 1265 1571 1269
rect 1631 1265 1635 1269
rect 1711 1265 1715 1269
rect 1799 1265 1803 1269
rect 1895 1265 1899 1269
rect 1991 1265 1995 1269
rect 2095 1265 2099 1269
rect 2207 1265 2211 1269
rect 2319 1265 2323 1269
rect 2503 1264 2507 1268
rect 1327 1247 1331 1251
rect 1551 1244 1555 1248
rect 1615 1244 1619 1248
rect 1695 1244 1699 1248
rect 1783 1244 1787 1248
rect 1879 1244 1883 1248
rect 1975 1244 1979 1248
rect 2079 1244 2083 1248
rect 2191 1244 2195 1248
rect 2303 1244 2307 1248
rect 2503 1247 2507 1251
rect 111 1236 115 1240
rect 151 1237 155 1241
rect 215 1237 219 1241
rect 303 1237 307 1241
rect 391 1237 395 1241
rect 471 1237 475 1241
rect 551 1237 555 1241
rect 623 1237 627 1241
rect 695 1237 699 1241
rect 767 1237 771 1241
rect 839 1237 843 1241
rect 919 1237 923 1241
rect 1287 1236 1291 1240
rect 1327 1225 1331 1229
rect 1519 1228 1523 1232
rect 1575 1228 1579 1232
rect 1631 1228 1635 1232
rect 1687 1228 1691 1232
rect 1743 1228 1747 1232
rect 1799 1228 1803 1232
rect 1855 1228 1859 1232
rect 1911 1228 1915 1232
rect 1967 1228 1971 1232
rect 2031 1228 2035 1232
rect 2103 1228 2107 1232
rect 2183 1228 2187 1232
rect 2271 1228 2275 1232
rect 2367 1228 2371 1232
rect 2439 1228 2443 1232
rect 2503 1225 2507 1229
rect 111 1219 115 1223
rect 135 1216 139 1220
rect 199 1216 203 1220
rect 287 1216 291 1220
rect 375 1216 379 1220
rect 455 1216 459 1220
rect 535 1216 539 1220
rect 607 1216 611 1220
rect 679 1216 683 1220
rect 751 1216 755 1220
rect 823 1216 827 1220
rect 903 1216 907 1220
rect 1287 1219 1291 1223
rect 1327 1208 1331 1212
rect 1535 1207 1539 1211
rect 1591 1207 1595 1211
rect 1647 1207 1651 1211
rect 1703 1207 1707 1211
rect 1759 1207 1763 1211
rect 1815 1207 1819 1211
rect 1871 1207 1875 1211
rect 1927 1207 1931 1211
rect 1983 1207 1987 1211
rect 2047 1207 2051 1211
rect 2119 1207 2123 1211
rect 2199 1207 2203 1211
rect 2287 1207 2291 1211
rect 2383 1207 2387 1211
rect 2455 1207 2459 1211
rect 2503 1208 2507 1212
rect 111 1197 115 1201
rect 135 1200 139 1204
rect 191 1200 195 1204
rect 271 1200 275 1204
rect 351 1200 355 1204
rect 431 1200 435 1204
rect 511 1200 515 1204
rect 583 1200 587 1204
rect 647 1200 651 1204
rect 719 1200 723 1204
rect 791 1200 795 1204
rect 863 1200 867 1204
rect 1287 1197 1291 1201
rect 111 1180 115 1184
rect 151 1179 155 1183
rect 207 1179 211 1183
rect 287 1179 291 1183
rect 367 1179 371 1183
rect 447 1179 451 1183
rect 527 1179 531 1183
rect 599 1179 603 1183
rect 663 1179 667 1183
rect 735 1179 739 1183
rect 807 1179 811 1183
rect 879 1179 883 1183
rect 1287 1180 1291 1184
rect 1327 1152 1331 1156
rect 1567 1153 1571 1157
rect 1631 1153 1635 1157
rect 1703 1153 1707 1157
rect 1791 1153 1795 1157
rect 1903 1153 1907 1157
rect 2031 1153 2035 1157
rect 2175 1153 2179 1157
rect 2327 1153 2331 1157
rect 2455 1153 2459 1157
rect 2503 1152 2507 1156
rect 1327 1135 1331 1139
rect 1551 1132 1555 1136
rect 1615 1132 1619 1136
rect 1687 1132 1691 1136
rect 1775 1132 1779 1136
rect 1887 1132 1891 1136
rect 2015 1132 2019 1136
rect 2159 1132 2163 1136
rect 2311 1132 2315 1136
rect 2439 1132 2443 1136
rect 2503 1135 2507 1139
rect 111 1124 115 1128
rect 183 1125 187 1129
rect 279 1125 283 1129
rect 375 1125 379 1129
rect 471 1125 475 1129
rect 567 1125 571 1129
rect 655 1125 659 1129
rect 735 1125 739 1129
rect 807 1125 811 1129
rect 879 1125 883 1129
rect 959 1125 963 1129
rect 1039 1125 1043 1129
rect 1287 1124 1291 1128
rect 1327 1117 1331 1121
rect 1383 1120 1387 1124
rect 1447 1120 1451 1124
rect 1519 1120 1523 1124
rect 1591 1120 1595 1124
rect 1671 1120 1675 1124
rect 1751 1120 1755 1124
rect 1831 1120 1835 1124
rect 1911 1120 1915 1124
rect 1983 1120 1987 1124
rect 2055 1120 2059 1124
rect 2135 1120 2139 1124
rect 2215 1120 2219 1124
rect 2503 1117 2507 1121
rect 111 1107 115 1111
rect 167 1104 171 1108
rect 263 1104 267 1108
rect 359 1104 363 1108
rect 455 1104 459 1108
rect 551 1104 555 1108
rect 639 1104 643 1108
rect 719 1104 723 1108
rect 791 1104 795 1108
rect 863 1104 867 1108
rect 943 1104 947 1108
rect 1023 1104 1027 1108
rect 1287 1107 1291 1111
rect 1327 1100 1331 1104
rect 1399 1099 1403 1103
rect 1463 1099 1467 1103
rect 1535 1099 1539 1103
rect 1607 1099 1611 1103
rect 1687 1099 1691 1103
rect 1767 1099 1771 1103
rect 1847 1099 1851 1103
rect 1927 1099 1931 1103
rect 1999 1099 2003 1103
rect 2071 1099 2075 1103
rect 2151 1099 2155 1103
rect 2231 1099 2235 1103
rect 2503 1100 2507 1104
rect 111 1081 115 1085
rect 207 1084 211 1088
rect 279 1084 283 1088
rect 359 1084 363 1088
rect 447 1084 451 1088
rect 543 1084 547 1088
rect 639 1084 643 1088
rect 727 1084 731 1088
rect 815 1084 819 1088
rect 895 1084 899 1088
rect 975 1084 979 1088
rect 1055 1084 1059 1088
rect 1143 1084 1147 1088
rect 1287 1081 1291 1085
rect 111 1064 115 1068
rect 223 1063 227 1067
rect 295 1063 299 1067
rect 375 1063 379 1067
rect 463 1063 467 1067
rect 559 1063 563 1067
rect 655 1063 659 1067
rect 743 1063 747 1067
rect 831 1063 835 1067
rect 911 1063 915 1067
rect 991 1063 995 1067
rect 1071 1063 1075 1067
rect 1159 1063 1163 1067
rect 1287 1064 1291 1068
rect 1327 1040 1331 1044
rect 1367 1041 1371 1045
rect 1455 1041 1459 1045
rect 1575 1041 1579 1045
rect 1695 1041 1699 1045
rect 1815 1041 1819 1045
rect 1927 1041 1931 1045
rect 2039 1041 2043 1045
rect 2151 1041 2155 1045
rect 2255 1041 2259 1045
rect 2367 1041 2371 1045
rect 2455 1041 2459 1045
rect 2503 1040 2507 1044
rect 1327 1023 1331 1027
rect 1351 1020 1355 1024
rect 1439 1020 1443 1024
rect 1559 1020 1563 1024
rect 1679 1020 1683 1024
rect 1799 1020 1803 1024
rect 1911 1020 1915 1024
rect 2023 1020 2027 1024
rect 2135 1020 2139 1024
rect 2239 1020 2243 1024
rect 2351 1020 2355 1024
rect 2439 1020 2443 1024
rect 2503 1023 2507 1027
rect 111 1004 115 1008
rect 295 1005 299 1009
rect 383 1005 387 1009
rect 479 1005 483 1009
rect 575 1005 579 1009
rect 671 1005 675 1009
rect 767 1005 771 1009
rect 855 1005 859 1009
rect 943 1005 947 1009
rect 1023 1005 1027 1009
rect 1103 1005 1107 1009
rect 1183 1005 1187 1009
rect 1239 1005 1243 1009
rect 1287 1004 1291 1008
rect 1327 1001 1331 1005
rect 1351 1004 1355 1008
rect 1511 1004 1515 1008
rect 1679 1004 1683 1008
rect 1823 1004 1827 1008
rect 1951 1004 1955 1008
rect 2071 1004 2075 1008
rect 2175 1004 2179 1008
rect 2271 1004 2275 1008
rect 2367 1004 2371 1008
rect 2439 1004 2443 1008
rect 2503 1001 2507 1005
rect 111 987 115 991
rect 279 984 283 988
rect 367 984 371 988
rect 463 984 467 988
rect 559 984 563 988
rect 655 984 659 988
rect 751 984 755 988
rect 839 984 843 988
rect 927 984 931 988
rect 1007 984 1011 988
rect 1087 984 1091 988
rect 1167 984 1171 988
rect 1223 984 1227 988
rect 1287 987 1291 991
rect 1327 984 1331 988
rect 1367 983 1371 987
rect 1527 983 1531 987
rect 1695 983 1699 987
rect 1839 983 1843 987
rect 1967 983 1971 987
rect 2087 983 2091 987
rect 2191 983 2195 987
rect 2287 983 2291 987
rect 2383 983 2387 987
rect 2455 983 2459 987
rect 2503 984 2507 988
rect 111 969 115 973
rect 271 972 275 976
rect 359 972 363 976
rect 455 972 459 976
rect 551 972 555 976
rect 655 972 659 976
rect 751 972 755 976
rect 839 972 843 976
rect 927 972 931 976
rect 1007 972 1011 976
rect 1087 972 1091 976
rect 1167 972 1171 976
rect 1223 972 1227 976
rect 1287 969 1291 973
rect 111 952 115 956
rect 287 951 291 955
rect 375 951 379 955
rect 471 951 475 955
rect 567 951 571 955
rect 671 951 675 955
rect 767 951 771 955
rect 855 951 859 955
rect 943 951 947 955
rect 1023 951 1027 955
rect 1103 951 1107 955
rect 1183 951 1187 955
rect 1239 951 1243 955
rect 1287 952 1291 956
rect 1327 920 1331 924
rect 1367 921 1371 925
rect 1423 921 1427 925
rect 1503 921 1507 925
rect 1607 921 1611 925
rect 1719 921 1723 925
rect 1831 921 1835 925
rect 1935 921 1939 925
rect 2031 921 2035 925
rect 2127 921 2131 925
rect 2215 921 2219 925
rect 2295 921 2299 925
rect 2375 921 2379 925
rect 2455 921 2459 925
rect 2503 920 2507 924
rect 1327 903 1331 907
rect 1351 900 1355 904
rect 1407 900 1411 904
rect 1487 900 1491 904
rect 1591 900 1595 904
rect 1703 900 1707 904
rect 1815 900 1819 904
rect 1919 900 1923 904
rect 2015 900 2019 904
rect 2111 900 2115 904
rect 2199 900 2203 904
rect 2279 900 2283 904
rect 2359 900 2363 904
rect 2439 900 2443 904
rect 2503 903 2507 907
rect 111 892 115 896
rect 271 893 275 897
rect 343 893 347 897
rect 423 893 427 897
rect 519 893 523 897
rect 615 893 619 897
rect 711 893 715 897
rect 807 893 811 897
rect 903 893 907 897
rect 991 893 995 897
rect 1087 893 1091 897
rect 1183 893 1187 897
rect 1287 892 1291 896
rect 1327 881 1331 885
rect 1431 884 1435 888
rect 1487 884 1491 888
rect 1551 884 1555 888
rect 1623 884 1627 888
rect 1703 884 1707 888
rect 1791 884 1795 888
rect 1895 884 1899 888
rect 2015 884 2019 888
rect 2143 884 2147 888
rect 2279 884 2283 888
rect 2423 884 2427 888
rect 2503 881 2507 885
rect 111 875 115 879
rect 255 872 259 876
rect 327 872 331 876
rect 407 872 411 876
rect 503 872 507 876
rect 599 872 603 876
rect 695 872 699 876
rect 791 872 795 876
rect 887 872 891 876
rect 975 872 979 876
rect 1071 872 1075 876
rect 1167 872 1171 876
rect 1287 875 1291 879
rect 1327 864 1331 868
rect 1447 863 1451 867
rect 1503 863 1507 867
rect 1567 863 1571 867
rect 1639 863 1643 867
rect 1719 863 1723 867
rect 1807 863 1811 867
rect 1911 863 1915 867
rect 2031 863 2035 867
rect 2159 863 2163 867
rect 2295 863 2299 867
rect 2439 863 2443 867
rect 2503 864 2507 868
rect 111 853 115 857
rect 247 856 251 860
rect 311 856 315 860
rect 375 856 379 860
rect 439 856 443 860
rect 503 856 507 860
rect 567 856 571 860
rect 631 856 635 860
rect 695 856 699 860
rect 759 856 763 860
rect 831 856 835 860
rect 903 856 907 860
rect 1287 853 1291 857
rect 111 836 115 840
rect 263 835 267 839
rect 327 835 331 839
rect 391 835 395 839
rect 455 835 459 839
rect 519 835 523 839
rect 583 835 587 839
rect 647 835 651 839
rect 711 835 715 839
rect 775 835 779 839
rect 847 835 851 839
rect 919 835 923 839
rect 1287 836 1291 840
rect 1327 808 1331 812
rect 1591 809 1595 813
rect 1647 809 1651 813
rect 1703 809 1707 813
rect 1767 809 1771 813
rect 1847 809 1851 813
rect 1927 809 1931 813
rect 2015 809 2019 813
rect 2103 809 2107 813
rect 2191 809 2195 813
rect 2287 809 2291 813
rect 2383 809 2387 813
rect 2455 809 2459 813
rect 2503 808 2507 812
rect 1327 791 1331 795
rect 1575 788 1579 792
rect 1631 788 1635 792
rect 1687 788 1691 792
rect 1751 788 1755 792
rect 1831 788 1835 792
rect 1911 788 1915 792
rect 1999 788 2003 792
rect 2087 788 2091 792
rect 2175 788 2179 792
rect 2271 788 2275 792
rect 2367 788 2371 792
rect 2439 788 2443 792
rect 2503 791 2507 795
rect 111 780 115 784
rect 215 781 219 785
rect 303 781 307 785
rect 391 781 395 785
rect 479 781 483 785
rect 559 781 563 785
rect 631 781 635 785
rect 703 781 707 785
rect 767 781 771 785
rect 831 781 835 785
rect 895 781 899 785
rect 967 781 971 785
rect 1039 781 1043 785
rect 1287 780 1291 784
rect 1327 769 1331 773
rect 1567 772 1571 776
rect 1623 772 1627 776
rect 1687 772 1691 776
rect 1759 772 1763 776
rect 1831 772 1835 776
rect 1919 772 1923 776
rect 2015 772 2019 776
rect 2119 772 2123 776
rect 2231 772 2235 776
rect 2343 772 2347 776
rect 2439 772 2443 776
rect 2503 769 2507 773
rect 111 763 115 767
rect 199 760 203 764
rect 287 760 291 764
rect 375 760 379 764
rect 463 760 467 764
rect 543 760 547 764
rect 615 760 619 764
rect 687 760 691 764
rect 751 760 755 764
rect 815 760 819 764
rect 879 760 883 764
rect 951 760 955 764
rect 1023 760 1027 764
rect 1287 763 1291 767
rect 111 745 115 749
rect 135 748 139 752
rect 255 748 259 752
rect 391 748 395 752
rect 519 748 523 752
rect 647 748 651 752
rect 775 748 779 752
rect 903 748 907 752
rect 1039 748 1043 752
rect 1327 752 1331 756
rect 1583 751 1587 755
rect 1639 751 1643 755
rect 1703 751 1707 755
rect 1775 751 1779 755
rect 1847 751 1851 755
rect 1935 751 1939 755
rect 2031 751 2035 755
rect 2135 751 2139 755
rect 2247 751 2251 755
rect 2359 751 2363 755
rect 2455 751 2459 755
rect 2503 752 2507 756
rect 1287 745 1291 749
rect 111 728 115 732
rect 151 727 155 731
rect 271 727 275 731
rect 407 727 411 731
rect 535 727 539 731
rect 663 727 667 731
rect 791 727 795 731
rect 919 727 923 731
rect 1055 727 1059 731
rect 1287 728 1291 732
rect 1327 700 1331 704
rect 1367 701 1371 705
rect 1431 701 1435 705
rect 1527 701 1531 705
rect 1631 701 1635 705
rect 1735 701 1739 705
rect 1839 701 1843 705
rect 1943 701 1947 705
rect 2047 701 2051 705
rect 2151 701 2155 705
rect 2255 701 2259 705
rect 2367 701 2371 705
rect 2455 701 2459 705
rect 2503 700 2507 704
rect 1327 683 1331 687
rect 111 676 115 680
rect 151 677 155 681
rect 207 677 211 681
rect 295 677 299 681
rect 391 677 395 681
rect 503 677 507 681
rect 623 677 627 681
rect 743 677 747 681
rect 871 677 875 681
rect 999 677 1003 681
rect 1127 677 1131 681
rect 1239 677 1243 681
rect 1287 676 1291 680
rect 1351 680 1355 684
rect 1415 680 1419 684
rect 1511 680 1515 684
rect 1615 680 1619 684
rect 1719 680 1723 684
rect 1823 680 1827 684
rect 1927 680 1931 684
rect 2031 680 2035 684
rect 2135 680 2139 684
rect 2239 680 2243 684
rect 2351 680 2355 684
rect 2439 680 2443 684
rect 2503 683 2507 687
rect 111 659 115 663
rect 135 656 139 660
rect 191 656 195 660
rect 279 656 283 660
rect 375 656 379 660
rect 487 656 491 660
rect 607 656 611 660
rect 727 656 731 660
rect 855 656 859 660
rect 983 656 987 660
rect 1111 656 1115 660
rect 1223 656 1227 660
rect 1287 659 1291 663
rect 1327 653 1331 657
rect 1351 656 1355 660
rect 1415 656 1419 660
rect 1511 656 1515 660
rect 1607 656 1611 660
rect 1711 656 1715 660
rect 1823 656 1827 660
rect 1935 656 1939 660
rect 2055 656 2059 660
rect 2183 656 2187 660
rect 2319 656 2323 660
rect 2439 656 2443 660
rect 2503 653 2507 657
rect 111 637 115 641
rect 151 640 155 644
rect 263 640 267 644
rect 367 640 371 644
rect 463 640 467 644
rect 559 640 563 644
rect 655 640 659 644
rect 751 640 755 644
rect 847 640 851 644
rect 943 640 947 644
rect 1039 640 1043 644
rect 1143 640 1147 644
rect 1223 640 1227 644
rect 1287 637 1291 641
rect 1327 636 1331 640
rect 1367 635 1371 639
rect 1431 635 1435 639
rect 1527 635 1531 639
rect 1623 635 1627 639
rect 1727 635 1731 639
rect 1839 635 1843 639
rect 1951 635 1955 639
rect 2071 635 2075 639
rect 2199 635 2203 639
rect 2335 635 2339 639
rect 2455 635 2459 639
rect 2503 636 2507 640
rect 111 620 115 624
rect 167 619 171 623
rect 279 619 283 623
rect 383 619 387 623
rect 479 619 483 623
rect 575 619 579 623
rect 671 619 675 623
rect 767 619 771 623
rect 863 619 867 623
rect 959 619 963 623
rect 1055 619 1059 623
rect 1159 619 1163 623
rect 1239 619 1243 623
rect 1287 620 1291 624
rect 1327 584 1331 588
rect 1383 585 1387 589
rect 1463 585 1467 589
rect 1551 585 1555 589
rect 1647 585 1651 589
rect 1743 585 1747 589
rect 1847 585 1851 589
rect 1959 585 1963 589
rect 2079 585 2083 589
rect 2207 585 2211 589
rect 2343 585 2347 589
rect 2455 585 2459 589
rect 2503 584 2507 588
rect 111 568 115 572
rect 151 569 155 573
rect 239 569 243 573
rect 335 569 339 573
rect 431 569 435 573
rect 535 569 539 573
rect 631 569 635 573
rect 727 569 731 573
rect 823 569 827 573
rect 911 569 915 573
rect 999 569 1003 573
rect 1087 569 1091 573
rect 1183 569 1187 573
rect 1287 568 1291 572
rect 1327 567 1331 571
rect 1367 564 1371 568
rect 1447 564 1451 568
rect 1535 564 1539 568
rect 1631 564 1635 568
rect 1727 564 1731 568
rect 1831 564 1835 568
rect 1943 564 1947 568
rect 2063 564 2067 568
rect 2191 564 2195 568
rect 2327 564 2331 568
rect 2439 564 2443 568
rect 2503 567 2507 571
rect 111 551 115 555
rect 135 548 139 552
rect 223 548 227 552
rect 319 548 323 552
rect 415 548 419 552
rect 519 548 523 552
rect 615 548 619 552
rect 711 548 715 552
rect 807 548 811 552
rect 895 548 899 552
rect 983 548 987 552
rect 1071 548 1075 552
rect 1167 548 1171 552
rect 1287 551 1291 555
rect 1327 549 1331 553
rect 1375 552 1379 556
rect 1455 552 1459 556
rect 1551 552 1555 556
rect 1647 552 1651 556
rect 1751 552 1755 556
rect 1855 552 1859 556
rect 1959 552 1963 556
rect 2055 552 2059 556
rect 2151 552 2155 556
rect 2255 552 2259 556
rect 2359 552 2363 556
rect 2439 552 2443 556
rect 2503 549 2507 553
rect 111 525 115 529
rect 143 528 147 532
rect 239 528 243 532
rect 335 528 339 532
rect 431 528 435 532
rect 527 528 531 532
rect 623 528 627 532
rect 711 528 715 532
rect 791 528 795 532
rect 871 528 875 532
rect 951 528 955 532
rect 1031 528 1035 532
rect 1327 532 1331 536
rect 1391 531 1395 535
rect 1471 531 1475 535
rect 1567 531 1571 535
rect 1663 531 1667 535
rect 1767 531 1771 535
rect 1871 531 1875 535
rect 1975 531 1979 535
rect 2071 531 2075 535
rect 2167 531 2171 535
rect 2271 531 2275 535
rect 2375 531 2379 535
rect 2455 531 2459 535
rect 2503 532 2507 536
rect 1287 525 1291 529
rect 111 508 115 512
rect 159 507 163 511
rect 255 507 259 511
rect 351 507 355 511
rect 447 507 451 511
rect 543 507 547 511
rect 639 507 643 511
rect 727 507 731 511
rect 807 507 811 511
rect 887 507 891 511
rect 967 507 971 511
rect 1047 507 1051 511
rect 1287 508 1291 512
rect 1327 476 1331 480
rect 1367 477 1371 481
rect 1455 477 1459 481
rect 1575 477 1579 481
rect 1695 477 1699 481
rect 1807 477 1811 481
rect 1919 477 1923 481
rect 2023 477 2027 481
rect 2119 477 2123 481
rect 2207 477 2211 481
rect 2295 477 2299 481
rect 2383 477 2387 481
rect 2455 477 2459 481
rect 2503 476 2507 480
rect 1327 459 1331 463
rect 111 452 115 456
rect 151 453 155 457
rect 207 453 211 457
rect 287 453 291 457
rect 375 453 379 457
rect 463 453 467 457
rect 559 453 563 457
rect 655 453 659 457
rect 751 453 755 457
rect 847 453 851 457
rect 951 453 955 457
rect 1055 453 1059 457
rect 1159 453 1163 457
rect 1239 453 1243 457
rect 1287 452 1291 456
rect 1351 456 1355 460
rect 1439 456 1443 460
rect 1559 456 1563 460
rect 1679 456 1683 460
rect 1791 456 1795 460
rect 1903 456 1907 460
rect 2007 456 2011 460
rect 2103 456 2107 460
rect 2191 456 2195 460
rect 2279 456 2283 460
rect 2367 456 2371 460
rect 2439 456 2443 460
rect 2503 459 2507 463
rect 111 435 115 439
rect 135 432 139 436
rect 191 432 195 436
rect 271 432 275 436
rect 359 432 363 436
rect 447 432 451 436
rect 543 432 547 436
rect 639 432 643 436
rect 735 432 739 436
rect 831 432 835 436
rect 935 432 939 436
rect 1039 432 1043 436
rect 1143 432 1147 436
rect 1223 432 1227 436
rect 1287 435 1291 439
rect 1327 429 1331 433
rect 1583 432 1587 436
rect 1639 432 1643 436
rect 1695 432 1699 436
rect 1759 432 1763 436
rect 1831 432 1835 436
rect 1911 432 1915 436
rect 1991 432 1995 436
rect 2079 432 2083 436
rect 2175 432 2179 436
rect 2271 432 2275 436
rect 2367 432 2371 436
rect 2439 432 2443 436
rect 2503 429 2507 433
rect 111 417 115 421
rect 135 420 139 424
rect 191 420 195 424
rect 279 420 283 424
rect 383 420 387 424
rect 495 420 499 424
rect 607 420 611 424
rect 719 420 723 424
rect 831 420 835 424
rect 935 420 939 424
rect 1039 420 1043 424
rect 1143 420 1147 424
rect 1223 420 1227 424
rect 1287 417 1291 421
rect 1327 412 1331 416
rect 1599 411 1603 415
rect 1655 411 1659 415
rect 1711 411 1715 415
rect 1775 411 1779 415
rect 1847 411 1851 415
rect 1927 411 1931 415
rect 2007 411 2011 415
rect 2095 411 2099 415
rect 2191 411 2195 415
rect 2287 411 2291 415
rect 2383 411 2387 415
rect 2455 411 2459 415
rect 2503 412 2507 416
rect 111 400 115 404
rect 151 399 155 403
rect 207 399 211 403
rect 295 399 299 403
rect 399 399 403 403
rect 511 399 515 403
rect 623 399 627 403
rect 735 399 739 403
rect 847 399 851 403
rect 951 399 955 403
rect 1055 399 1059 403
rect 1159 399 1163 403
rect 1239 399 1243 403
rect 1287 400 1291 404
rect 1327 356 1331 360
rect 1679 357 1683 361
rect 1735 357 1739 361
rect 1799 357 1803 361
rect 1871 357 1875 361
rect 1943 357 1947 361
rect 2023 357 2027 361
rect 2111 357 2115 361
rect 2199 357 2203 361
rect 2287 357 2291 361
rect 2375 357 2379 361
rect 2455 357 2459 361
rect 2503 356 2507 360
rect 111 344 115 348
rect 151 345 155 349
rect 231 345 235 349
rect 335 345 339 349
rect 439 345 443 349
rect 543 345 547 349
rect 647 345 651 349
rect 751 345 755 349
rect 847 345 851 349
rect 935 345 939 349
rect 1015 345 1019 349
rect 1095 345 1099 349
rect 1175 345 1179 349
rect 1239 345 1243 349
rect 1287 344 1291 348
rect 1327 339 1331 343
rect 1663 336 1667 340
rect 1719 336 1723 340
rect 1783 336 1787 340
rect 1855 336 1859 340
rect 1927 336 1931 340
rect 2007 336 2011 340
rect 2095 336 2099 340
rect 2183 336 2187 340
rect 2271 336 2275 340
rect 2359 336 2363 340
rect 2439 336 2443 340
rect 2503 339 2507 343
rect 111 327 115 331
rect 135 324 139 328
rect 215 324 219 328
rect 319 324 323 328
rect 423 324 427 328
rect 527 324 531 328
rect 631 324 635 328
rect 735 324 739 328
rect 831 324 835 328
rect 919 324 923 328
rect 999 324 1003 328
rect 1079 324 1083 328
rect 1159 324 1163 328
rect 1223 324 1227 328
rect 1287 327 1291 331
rect 1327 313 1331 317
rect 1351 316 1355 320
rect 1455 316 1459 320
rect 1583 316 1587 320
rect 1711 316 1715 320
rect 1839 316 1843 320
rect 1951 316 1955 320
rect 2063 316 2067 320
rect 2167 316 2171 320
rect 2263 316 2267 320
rect 2359 316 2363 320
rect 2439 316 2443 320
rect 111 305 115 309
rect 135 308 139 312
rect 215 308 219 312
rect 319 308 323 312
rect 423 308 427 312
rect 535 308 539 312
rect 639 308 643 312
rect 743 308 747 312
rect 847 308 851 312
rect 943 308 947 312
rect 1039 308 1043 312
rect 1143 308 1147 312
rect 2503 313 2507 317
rect 1223 308 1227 312
rect 1287 305 1291 309
rect 1327 296 1331 300
rect 1367 295 1371 299
rect 1471 295 1475 299
rect 1599 295 1603 299
rect 1727 295 1731 299
rect 1855 295 1859 299
rect 1967 295 1971 299
rect 2079 295 2083 299
rect 2183 295 2187 299
rect 2279 295 2283 299
rect 2375 295 2379 299
rect 2455 295 2459 299
rect 2503 296 2507 300
rect 111 288 115 292
rect 151 287 155 291
rect 231 287 235 291
rect 335 287 339 291
rect 439 287 443 291
rect 551 287 555 291
rect 655 287 659 291
rect 759 287 763 291
rect 863 287 867 291
rect 959 287 963 291
rect 1055 287 1059 291
rect 1159 287 1163 291
rect 1239 287 1243 291
rect 1287 288 1291 292
rect 111 236 115 240
rect 151 237 155 241
rect 223 237 227 241
rect 319 237 323 241
rect 423 237 427 241
rect 535 237 539 241
rect 647 237 651 241
rect 759 237 763 241
rect 871 237 875 241
rect 983 237 987 241
rect 1103 237 1107 241
rect 1223 237 1227 241
rect 1287 236 1291 240
rect 1327 236 1331 240
rect 1367 237 1371 241
rect 1447 237 1451 241
rect 1551 237 1555 241
rect 1655 237 1659 241
rect 1759 237 1763 241
rect 1863 237 1867 241
rect 1967 237 1971 241
rect 2071 237 2075 241
rect 2175 237 2179 241
rect 2271 237 2275 241
rect 2375 237 2379 241
rect 2455 237 2459 241
rect 2503 236 2507 240
rect 111 219 115 223
rect 135 216 139 220
rect 207 216 211 220
rect 303 216 307 220
rect 407 216 411 220
rect 519 216 523 220
rect 631 216 635 220
rect 743 216 747 220
rect 855 216 859 220
rect 967 216 971 220
rect 1087 216 1091 220
rect 1207 216 1211 220
rect 1287 219 1291 223
rect 1327 219 1331 223
rect 1351 216 1355 220
rect 1431 216 1435 220
rect 1535 216 1539 220
rect 1639 216 1643 220
rect 1743 216 1747 220
rect 1847 216 1851 220
rect 1951 216 1955 220
rect 2055 216 2059 220
rect 2159 216 2163 220
rect 2255 216 2259 220
rect 2359 216 2363 220
rect 2439 216 2443 220
rect 2503 219 2507 223
rect 111 197 115 201
rect 183 200 187 204
rect 279 200 283 204
rect 383 200 387 204
rect 487 200 491 204
rect 591 200 595 204
rect 695 200 699 204
rect 799 200 803 204
rect 895 200 899 204
rect 999 200 1003 204
rect 1103 200 1107 204
rect 1287 197 1291 201
rect 1327 197 1331 201
rect 1351 200 1355 204
rect 1407 200 1411 204
rect 1471 200 1475 204
rect 1551 200 1555 204
rect 1639 200 1643 204
rect 1719 200 1723 204
rect 1807 200 1811 204
rect 1895 200 1899 204
rect 1991 200 1995 204
rect 2103 200 2107 204
rect 2215 200 2219 204
rect 2335 200 2339 204
rect 2439 200 2443 204
rect 2503 197 2507 201
rect 111 180 115 184
rect 199 179 203 183
rect 295 179 299 183
rect 399 179 403 183
rect 503 179 507 183
rect 607 179 611 183
rect 711 179 715 183
rect 815 179 819 183
rect 911 179 915 183
rect 1015 179 1019 183
rect 1119 179 1123 183
rect 1287 180 1291 184
rect 1327 180 1331 184
rect 1367 179 1371 183
rect 1423 179 1427 183
rect 1487 179 1491 183
rect 1567 179 1571 183
rect 1655 179 1659 183
rect 1735 179 1739 183
rect 1823 179 1827 183
rect 1911 179 1915 183
rect 2007 179 2011 183
rect 2119 179 2123 183
rect 2231 179 2235 183
rect 2351 179 2355 183
rect 2455 179 2459 183
rect 2503 180 2507 184
rect 111 120 115 124
rect 151 121 155 125
rect 207 121 211 125
rect 263 121 267 125
rect 319 121 323 125
rect 375 121 379 125
rect 431 121 435 125
rect 487 121 491 125
rect 543 121 547 125
rect 599 121 603 125
rect 655 121 659 125
rect 711 121 715 125
rect 767 121 771 125
rect 831 121 835 125
rect 895 121 899 125
rect 959 121 963 125
rect 1023 121 1027 125
rect 1087 121 1091 125
rect 1151 121 1155 125
rect 1287 120 1291 124
rect 1327 108 1331 112
rect 1367 109 1371 113
rect 1423 109 1427 113
rect 1479 109 1483 113
rect 1535 109 1539 113
rect 1591 109 1595 113
rect 1647 109 1651 113
rect 1703 109 1707 113
rect 1759 109 1763 113
rect 1823 109 1827 113
rect 1879 109 1883 113
rect 1943 109 1947 113
rect 2007 109 2011 113
rect 2071 109 2075 113
rect 2143 109 2147 113
rect 2223 109 2227 113
rect 2303 109 2307 113
rect 2391 109 2395 113
rect 2455 109 2459 113
rect 2503 108 2507 112
rect 111 103 115 107
rect 135 100 139 104
rect 191 100 195 104
rect 247 100 251 104
rect 303 100 307 104
rect 359 100 363 104
rect 415 100 419 104
rect 471 100 475 104
rect 527 100 531 104
rect 583 100 587 104
rect 639 100 643 104
rect 695 100 699 104
rect 751 100 755 104
rect 815 100 819 104
rect 879 100 883 104
rect 943 100 947 104
rect 1007 100 1011 104
rect 1071 100 1075 104
rect 1135 100 1139 104
rect 1287 103 1291 107
rect 1327 91 1331 95
rect 1351 88 1355 92
rect 1407 88 1411 92
rect 1463 88 1467 92
rect 1519 88 1523 92
rect 1575 88 1579 92
rect 1631 88 1635 92
rect 1687 88 1691 92
rect 1743 88 1747 92
rect 1807 88 1811 92
rect 1863 88 1867 92
rect 1927 88 1931 92
rect 1991 88 1995 92
rect 2055 88 2059 92
rect 2127 88 2131 92
rect 2207 88 2211 92
rect 2287 88 2291 92
rect 2375 88 2379 92
rect 2439 88 2443 92
rect 2503 91 2507 95
<< m3 >>
rect 111 2582 115 2583
rect 111 2577 115 2578
rect 135 2582 139 2583
rect 135 2577 139 2578
rect 191 2582 195 2583
rect 191 2577 195 2578
rect 247 2582 251 2583
rect 247 2577 251 2578
rect 303 2582 307 2583
rect 303 2577 307 2578
rect 359 2582 363 2583
rect 359 2577 363 2578
rect 1287 2582 1291 2583
rect 1287 2577 1291 2578
rect 112 2574 114 2577
rect 134 2576 140 2577
rect 110 2573 116 2574
rect 110 2569 111 2573
rect 115 2569 116 2573
rect 134 2572 135 2576
rect 139 2572 140 2576
rect 134 2571 140 2572
rect 190 2576 196 2577
rect 190 2572 191 2576
rect 195 2572 196 2576
rect 190 2571 196 2572
rect 246 2576 252 2577
rect 246 2572 247 2576
rect 251 2572 252 2576
rect 246 2571 252 2572
rect 302 2576 308 2577
rect 302 2572 303 2576
rect 307 2572 308 2576
rect 302 2571 308 2572
rect 358 2576 364 2577
rect 358 2572 359 2576
rect 363 2572 364 2576
rect 1288 2574 1290 2577
rect 358 2571 364 2572
rect 1286 2573 1292 2574
rect 110 2568 116 2569
rect 1286 2569 1287 2573
rect 1291 2569 1292 2573
rect 1286 2568 1292 2569
rect 1327 2562 1331 2563
rect 1327 2557 1331 2558
rect 1495 2562 1499 2563
rect 1495 2557 1499 2558
rect 1551 2562 1555 2563
rect 1551 2557 1555 2558
rect 1607 2562 1611 2563
rect 1607 2557 1611 2558
rect 1663 2562 1667 2563
rect 1663 2557 1667 2558
rect 1719 2562 1723 2563
rect 1719 2557 1723 2558
rect 1775 2562 1779 2563
rect 1775 2557 1779 2558
rect 1831 2562 1835 2563
rect 1831 2557 1835 2558
rect 1887 2562 1891 2563
rect 1887 2557 1891 2558
rect 1943 2562 1947 2563
rect 1943 2557 1947 2558
rect 1999 2562 2003 2563
rect 1999 2557 2003 2558
rect 2055 2562 2059 2563
rect 2055 2557 2059 2558
rect 2111 2562 2115 2563
rect 2111 2557 2115 2558
rect 2167 2562 2171 2563
rect 2167 2557 2171 2558
rect 2503 2562 2507 2563
rect 2503 2557 2507 2558
rect 110 2556 116 2557
rect 1286 2556 1292 2557
rect 110 2552 111 2556
rect 115 2552 116 2556
rect 110 2551 116 2552
rect 150 2555 156 2556
rect 150 2551 151 2555
rect 155 2551 156 2555
rect 112 2531 114 2551
rect 150 2550 156 2551
rect 206 2555 212 2556
rect 206 2551 207 2555
rect 211 2551 212 2555
rect 206 2550 212 2551
rect 262 2555 268 2556
rect 262 2551 263 2555
rect 267 2551 268 2555
rect 262 2550 268 2551
rect 318 2555 324 2556
rect 318 2551 319 2555
rect 323 2551 324 2555
rect 318 2550 324 2551
rect 374 2555 380 2556
rect 374 2551 375 2555
rect 379 2551 380 2555
rect 1286 2552 1287 2556
rect 1291 2552 1292 2556
rect 1328 2554 1330 2557
rect 1494 2556 1500 2557
rect 1286 2551 1292 2552
rect 1326 2553 1332 2554
rect 374 2550 380 2551
rect 152 2531 154 2550
rect 208 2531 210 2550
rect 264 2531 266 2550
rect 320 2531 322 2550
rect 376 2531 378 2550
rect 1288 2531 1290 2551
rect 1326 2549 1327 2553
rect 1331 2549 1332 2553
rect 1494 2552 1495 2556
rect 1499 2552 1500 2556
rect 1494 2551 1500 2552
rect 1550 2556 1556 2557
rect 1550 2552 1551 2556
rect 1555 2552 1556 2556
rect 1550 2551 1556 2552
rect 1606 2556 1612 2557
rect 1606 2552 1607 2556
rect 1611 2552 1612 2556
rect 1606 2551 1612 2552
rect 1662 2556 1668 2557
rect 1662 2552 1663 2556
rect 1667 2552 1668 2556
rect 1662 2551 1668 2552
rect 1718 2556 1724 2557
rect 1718 2552 1719 2556
rect 1723 2552 1724 2556
rect 1718 2551 1724 2552
rect 1774 2556 1780 2557
rect 1774 2552 1775 2556
rect 1779 2552 1780 2556
rect 1774 2551 1780 2552
rect 1830 2556 1836 2557
rect 1830 2552 1831 2556
rect 1835 2552 1836 2556
rect 1830 2551 1836 2552
rect 1886 2556 1892 2557
rect 1886 2552 1887 2556
rect 1891 2552 1892 2556
rect 1886 2551 1892 2552
rect 1942 2556 1948 2557
rect 1942 2552 1943 2556
rect 1947 2552 1948 2556
rect 1942 2551 1948 2552
rect 1998 2556 2004 2557
rect 1998 2552 1999 2556
rect 2003 2552 2004 2556
rect 1998 2551 2004 2552
rect 2054 2556 2060 2557
rect 2054 2552 2055 2556
rect 2059 2552 2060 2556
rect 2054 2551 2060 2552
rect 2110 2556 2116 2557
rect 2110 2552 2111 2556
rect 2115 2552 2116 2556
rect 2110 2551 2116 2552
rect 2166 2556 2172 2557
rect 2166 2552 2167 2556
rect 2171 2552 2172 2556
rect 2504 2554 2506 2557
rect 2166 2551 2172 2552
rect 2502 2553 2508 2554
rect 1326 2548 1332 2549
rect 2502 2549 2503 2553
rect 2507 2549 2508 2553
rect 2502 2548 2508 2549
rect 1326 2536 1332 2537
rect 2502 2536 2508 2537
rect 1326 2532 1327 2536
rect 1331 2532 1332 2536
rect 1326 2531 1332 2532
rect 1510 2535 1516 2536
rect 1510 2531 1511 2535
rect 1515 2531 1516 2535
rect 111 2530 115 2531
rect 111 2525 115 2526
rect 151 2530 155 2531
rect 151 2525 155 2526
rect 207 2530 211 2531
rect 207 2525 211 2526
rect 223 2530 227 2531
rect 223 2525 227 2526
rect 263 2530 267 2531
rect 263 2525 267 2526
rect 279 2530 283 2531
rect 279 2525 283 2526
rect 319 2530 323 2531
rect 319 2525 323 2526
rect 343 2530 347 2531
rect 343 2525 347 2526
rect 375 2530 379 2531
rect 375 2525 379 2526
rect 415 2530 419 2531
rect 415 2525 419 2526
rect 487 2530 491 2531
rect 487 2525 491 2526
rect 551 2530 555 2531
rect 551 2525 555 2526
rect 615 2530 619 2531
rect 615 2525 619 2526
rect 679 2530 683 2531
rect 679 2525 683 2526
rect 743 2530 747 2531
rect 743 2525 747 2526
rect 807 2530 811 2531
rect 807 2525 811 2526
rect 871 2530 875 2531
rect 871 2525 875 2526
rect 935 2530 939 2531
rect 935 2525 939 2526
rect 999 2530 1003 2531
rect 999 2525 1003 2526
rect 1063 2530 1067 2531
rect 1063 2525 1067 2526
rect 1287 2530 1291 2531
rect 1287 2525 1291 2526
rect 112 2505 114 2525
rect 224 2506 226 2525
rect 280 2506 282 2525
rect 344 2506 346 2525
rect 416 2506 418 2525
rect 488 2506 490 2525
rect 552 2506 554 2525
rect 616 2506 618 2525
rect 680 2506 682 2525
rect 744 2506 746 2525
rect 808 2506 810 2525
rect 872 2506 874 2525
rect 936 2506 938 2525
rect 1000 2506 1002 2525
rect 1064 2506 1066 2525
rect 222 2505 228 2506
rect 110 2504 116 2505
rect 110 2500 111 2504
rect 115 2500 116 2504
rect 222 2501 223 2505
rect 227 2501 228 2505
rect 222 2500 228 2501
rect 278 2505 284 2506
rect 278 2501 279 2505
rect 283 2501 284 2505
rect 278 2500 284 2501
rect 342 2505 348 2506
rect 342 2501 343 2505
rect 347 2501 348 2505
rect 342 2500 348 2501
rect 414 2505 420 2506
rect 414 2501 415 2505
rect 419 2501 420 2505
rect 414 2500 420 2501
rect 486 2505 492 2506
rect 486 2501 487 2505
rect 491 2501 492 2505
rect 486 2500 492 2501
rect 550 2505 556 2506
rect 550 2501 551 2505
rect 555 2501 556 2505
rect 550 2500 556 2501
rect 614 2505 620 2506
rect 614 2501 615 2505
rect 619 2501 620 2505
rect 614 2500 620 2501
rect 678 2505 684 2506
rect 678 2501 679 2505
rect 683 2501 684 2505
rect 678 2500 684 2501
rect 742 2505 748 2506
rect 742 2501 743 2505
rect 747 2501 748 2505
rect 742 2500 748 2501
rect 806 2505 812 2506
rect 806 2501 807 2505
rect 811 2501 812 2505
rect 806 2500 812 2501
rect 870 2505 876 2506
rect 870 2501 871 2505
rect 875 2501 876 2505
rect 870 2500 876 2501
rect 934 2505 940 2506
rect 934 2501 935 2505
rect 939 2501 940 2505
rect 934 2500 940 2501
rect 998 2505 1004 2506
rect 998 2501 999 2505
rect 1003 2501 1004 2505
rect 998 2500 1004 2501
rect 1062 2505 1068 2506
rect 1288 2505 1290 2525
rect 1328 2511 1330 2531
rect 1510 2530 1516 2531
rect 1566 2535 1572 2536
rect 1566 2531 1567 2535
rect 1571 2531 1572 2535
rect 1566 2530 1572 2531
rect 1622 2535 1628 2536
rect 1622 2531 1623 2535
rect 1627 2531 1628 2535
rect 1622 2530 1628 2531
rect 1678 2535 1684 2536
rect 1678 2531 1679 2535
rect 1683 2531 1684 2535
rect 1678 2530 1684 2531
rect 1734 2535 1740 2536
rect 1734 2531 1735 2535
rect 1739 2531 1740 2535
rect 1734 2530 1740 2531
rect 1790 2535 1796 2536
rect 1790 2531 1791 2535
rect 1795 2531 1796 2535
rect 1790 2530 1796 2531
rect 1846 2535 1852 2536
rect 1846 2531 1847 2535
rect 1851 2531 1852 2535
rect 1846 2530 1852 2531
rect 1902 2535 1908 2536
rect 1902 2531 1903 2535
rect 1907 2531 1908 2535
rect 1902 2530 1908 2531
rect 1958 2535 1964 2536
rect 1958 2531 1959 2535
rect 1963 2531 1964 2535
rect 1958 2530 1964 2531
rect 2014 2535 2020 2536
rect 2014 2531 2015 2535
rect 2019 2531 2020 2535
rect 2014 2530 2020 2531
rect 2070 2535 2076 2536
rect 2070 2531 2071 2535
rect 2075 2531 2076 2535
rect 2070 2530 2076 2531
rect 2126 2535 2132 2536
rect 2126 2531 2127 2535
rect 2131 2531 2132 2535
rect 2126 2530 2132 2531
rect 2182 2535 2188 2536
rect 2182 2531 2183 2535
rect 2187 2531 2188 2535
rect 2502 2532 2503 2536
rect 2507 2532 2508 2536
rect 2502 2531 2508 2532
rect 2182 2530 2188 2531
rect 1512 2511 1514 2530
rect 1568 2511 1570 2530
rect 1624 2511 1626 2530
rect 1680 2511 1682 2530
rect 1736 2511 1738 2530
rect 1792 2511 1794 2530
rect 1848 2511 1850 2530
rect 1904 2511 1906 2530
rect 1960 2511 1962 2530
rect 2016 2511 2018 2530
rect 2072 2511 2074 2530
rect 2128 2511 2130 2530
rect 2184 2511 2186 2530
rect 2504 2511 2506 2531
rect 1327 2510 1331 2511
rect 1327 2505 1331 2506
rect 1511 2510 1515 2511
rect 1511 2505 1515 2506
rect 1543 2510 1547 2511
rect 1543 2505 1547 2506
rect 1567 2510 1571 2511
rect 1567 2505 1571 2506
rect 1607 2510 1611 2511
rect 1607 2505 1611 2506
rect 1623 2510 1627 2511
rect 1623 2505 1627 2506
rect 1679 2510 1683 2511
rect 1679 2505 1683 2506
rect 1735 2510 1739 2511
rect 1735 2505 1739 2506
rect 1751 2510 1755 2511
rect 1751 2505 1755 2506
rect 1791 2510 1795 2511
rect 1791 2505 1795 2506
rect 1823 2510 1827 2511
rect 1823 2505 1827 2506
rect 1847 2510 1851 2511
rect 1847 2505 1851 2506
rect 1895 2510 1899 2511
rect 1895 2505 1899 2506
rect 1903 2510 1907 2511
rect 1903 2505 1907 2506
rect 1959 2510 1963 2511
rect 1959 2505 1963 2506
rect 1967 2510 1971 2511
rect 1967 2505 1971 2506
rect 2015 2510 2019 2511
rect 2015 2505 2019 2506
rect 2039 2510 2043 2511
rect 2039 2505 2043 2506
rect 2071 2510 2075 2511
rect 2071 2505 2075 2506
rect 2111 2510 2115 2511
rect 2111 2505 2115 2506
rect 2127 2510 2131 2511
rect 2127 2505 2131 2506
rect 2183 2510 2187 2511
rect 2183 2505 2187 2506
rect 2503 2510 2507 2511
rect 2503 2505 2507 2506
rect 1062 2501 1063 2505
rect 1067 2501 1068 2505
rect 1062 2500 1068 2501
rect 1286 2504 1292 2505
rect 1286 2500 1287 2504
rect 1291 2500 1292 2504
rect 110 2499 116 2500
rect 1286 2499 1292 2500
rect 110 2487 116 2488
rect 110 2483 111 2487
rect 115 2483 116 2487
rect 1286 2487 1292 2488
rect 110 2482 116 2483
rect 206 2484 212 2485
rect 112 2471 114 2482
rect 206 2480 207 2484
rect 211 2480 212 2484
rect 206 2479 212 2480
rect 262 2484 268 2485
rect 262 2480 263 2484
rect 267 2480 268 2484
rect 262 2479 268 2480
rect 326 2484 332 2485
rect 326 2480 327 2484
rect 331 2480 332 2484
rect 326 2479 332 2480
rect 398 2484 404 2485
rect 398 2480 399 2484
rect 403 2480 404 2484
rect 398 2479 404 2480
rect 470 2484 476 2485
rect 470 2480 471 2484
rect 475 2480 476 2484
rect 470 2479 476 2480
rect 534 2484 540 2485
rect 534 2480 535 2484
rect 539 2480 540 2484
rect 534 2479 540 2480
rect 598 2484 604 2485
rect 598 2480 599 2484
rect 603 2480 604 2484
rect 598 2479 604 2480
rect 662 2484 668 2485
rect 662 2480 663 2484
rect 667 2480 668 2484
rect 662 2479 668 2480
rect 726 2484 732 2485
rect 726 2480 727 2484
rect 731 2480 732 2484
rect 726 2479 732 2480
rect 790 2484 796 2485
rect 790 2480 791 2484
rect 795 2480 796 2484
rect 790 2479 796 2480
rect 854 2484 860 2485
rect 854 2480 855 2484
rect 859 2480 860 2484
rect 854 2479 860 2480
rect 918 2484 924 2485
rect 918 2480 919 2484
rect 923 2480 924 2484
rect 918 2479 924 2480
rect 982 2484 988 2485
rect 982 2480 983 2484
rect 987 2480 988 2484
rect 982 2479 988 2480
rect 1046 2484 1052 2485
rect 1046 2480 1047 2484
rect 1051 2480 1052 2484
rect 1286 2483 1287 2487
rect 1291 2483 1292 2487
rect 1328 2485 1330 2505
rect 1544 2486 1546 2505
rect 1608 2486 1610 2505
rect 1680 2486 1682 2505
rect 1752 2486 1754 2505
rect 1824 2486 1826 2505
rect 1896 2486 1898 2505
rect 1968 2486 1970 2505
rect 2040 2486 2042 2505
rect 2112 2486 2114 2505
rect 2184 2486 2186 2505
rect 1542 2485 1548 2486
rect 1286 2482 1292 2483
rect 1326 2484 1332 2485
rect 1046 2479 1052 2480
rect 208 2471 210 2479
rect 264 2471 266 2479
rect 328 2471 330 2479
rect 400 2471 402 2479
rect 472 2471 474 2479
rect 536 2471 538 2479
rect 600 2471 602 2479
rect 664 2471 666 2479
rect 728 2471 730 2479
rect 792 2471 794 2479
rect 856 2471 858 2479
rect 920 2471 922 2479
rect 984 2471 986 2479
rect 1048 2471 1050 2479
rect 1288 2471 1290 2482
rect 1326 2480 1327 2484
rect 1331 2480 1332 2484
rect 1542 2481 1543 2485
rect 1547 2481 1548 2485
rect 1542 2480 1548 2481
rect 1606 2485 1612 2486
rect 1606 2481 1607 2485
rect 1611 2481 1612 2485
rect 1606 2480 1612 2481
rect 1678 2485 1684 2486
rect 1678 2481 1679 2485
rect 1683 2481 1684 2485
rect 1678 2480 1684 2481
rect 1750 2485 1756 2486
rect 1750 2481 1751 2485
rect 1755 2481 1756 2485
rect 1750 2480 1756 2481
rect 1822 2485 1828 2486
rect 1822 2481 1823 2485
rect 1827 2481 1828 2485
rect 1822 2480 1828 2481
rect 1894 2485 1900 2486
rect 1894 2481 1895 2485
rect 1899 2481 1900 2485
rect 1894 2480 1900 2481
rect 1966 2485 1972 2486
rect 1966 2481 1967 2485
rect 1971 2481 1972 2485
rect 1966 2480 1972 2481
rect 2038 2485 2044 2486
rect 2038 2481 2039 2485
rect 2043 2481 2044 2485
rect 2038 2480 2044 2481
rect 2110 2485 2116 2486
rect 2110 2481 2111 2485
rect 2115 2481 2116 2485
rect 2110 2480 2116 2481
rect 2182 2485 2188 2486
rect 2504 2485 2506 2505
rect 2182 2481 2183 2485
rect 2187 2481 2188 2485
rect 2182 2480 2188 2481
rect 2502 2484 2508 2485
rect 2502 2480 2503 2484
rect 2507 2480 2508 2484
rect 1326 2479 1332 2480
rect 2502 2479 2508 2480
rect 111 2470 115 2471
rect 111 2465 115 2466
rect 167 2470 171 2471
rect 167 2465 171 2466
rect 207 2470 211 2471
rect 207 2465 211 2466
rect 223 2470 227 2471
rect 223 2465 227 2466
rect 263 2470 267 2471
rect 263 2465 267 2466
rect 279 2470 283 2471
rect 279 2465 283 2466
rect 327 2470 331 2471
rect 327 2465 331 2466
rect 335 2470 339 2471
rect 335 2465 339 2466
rect 391 2470 395 2471
rect 391 2465 395 2466
rect 399 2470 403 2471
rect 399 2465 403 2466
rect 447 2470 451 2471
rect 447 2465 451 2466
rect 471 2470 475 2471
rect 471 2465 475 2466
rect 503 2470 507 2471
rect 503 2465 507 2466
rect 535 2470 539 2471
rect 535 2465 539 2466
rect 559 2470 563 2471
rect 559 2465 563 2466
rect 599 2470 603 2471
rect 599 2465 603 2466
rect 615 2470 619 2471
rect 615 2465 619 2466
rect 663 2470 667 2471
rect 663 2465 667 2466
rect 671 2470 675 2471
rect 671 2465 675 2466
rect 727 2470 731 2471
rect 727 2465 731 2466
rect 783 2470 787 2471
rect 783 2465 787 2466
rect 791 2470 795 2471
rect 791 2465 795 2466
rect 839 2470 843 2471
rect 839 2465 843 2466
rect 855 2470 859 2471
rect 855 2465 859 2466
rect 895 2470 899 2471
rect 895 2465 899 2466
rect 919 2470 923 2471
rect 919 2465 923 2466
rect 951 2470 955 2471
rect 951 2465 955 2466
rect 983 2470 987 2471
rect 983 2465 987 2466
rect 1007 2470 1011 2471
rect 1007 2465 1011 2466
rect 1047 2470 1051 2471
rect 1047 2465 1051 2466
rect 1063 2470 1067 2471
rect 1063 2465 1067 2466
rect 1287 2470 1291 2471
rect 1287 2465 1291 2466
rect 1326 2467 1332 2468
rect 112 2462 114 2465
rect 166 2464 172 2465
rect 110 2461 116 2462
rect 110 2457 111 2461
rect 115 2457 116 2461
rect 166 2460 167 2464
rect 171 2460 172 2464
rect 166 2459 172 2460
rect 222 2464 228 2465
rect 222 2460 223 2464
rect 227 2460 228 2464
rect 222 2459 228 2460
rect 278 2464 284 2465
rect 278 2460 279 2464
rect 283 2460 284 2464
rect 278 2459 284 2460
rect 334 2464 340 2465
rect 334 2460 335 2464
rect 339 2460 340 2464
rect 334 2459 340 2460
rect 390 2464 396 2465
rect 390 2460 391 2464
rect 395 2460 396 2464
rect 390 2459 396 2460
rect 446 2464 452 2465
rect 446 2460 447 2464
rect 451 2460 452 2464
rect 446 2459 452 2460
rect 502 2464 508 2465
rect 502 2460 503 2464
rect 507 2460 508 2464
rect 502 2459 508 2460
rect 558 2464 564 2465
rect 558 2460 559 2464
rect 563 2460 564 2464
rect 558 2459 564 2460
rect 614 2464 620 2465
rect 614 2460 615 2464
rect 619 2460 620 2464
rect 614 2459 620 2460
rect 670 2464 676 2465
rect 670 2460 671 2464
rect 675 2460 676 2464
rect 670 2459 676 2460
rect 726 2464 732 2465
rect 726 2460 727 2464
rect 731 2460 732 2464
rect 726 2459 732 2460
rect 782 2464 788 2465
rect 782 2460 783 2464
rect 787 2460 788 2464
rect 782 2459 788 2460
rect 838 2464 844 2465
rect 838 2460 839 2464
rect 843 2460 844 2464
rect 838 2459 844 2460
rect 894 2464 900 2465
rect 894 2460 895 2464
rect 899 2460 900 2464
rect 894 2459 900 2460
rect 950 2464 956 2465
rect 950 2460 951 2464
rect 955 2460 956 2464
rect 950 2459 956 2460
rect 1006 2464 1012 2465
rect 1006 2460 1007 2464
rect 1011 2460 1012 2464
rect 1006 2459 1012 2460
rect 1062 2464 1068 2465
rect 1062 2460 1063 2464
rect 1067 2460 1068 2464
rect 1288 2462 1290 2465
rect 1326 2463 1327 2467
rect 1331 2463 1332 2467
rect 2502 2467 2508 2468
rect 1326 2462 1332 2463
rect 1526 2464 1532 2465
rect 1062 2459 1068 2460
rect 1286 2461 1292 2462
rect 110 2456 116 2457
rect 1286 2457 1287 2461
rect 1291 2457 1292 2461
rect 1286 2456 1292 2457
rect 1328 2455 1330 2462
rect 1526 2460 1527 2464
rect 1531 2460 1532 2464
rect 1526 2459 1532 2460
rect 1590 2464 1596 2465
rect 1590 2460 1591 2464
rect 1595 2460 1596 2464
rect 1590 2459 1596 2460
rect 1662 2464 1668 2465
rect 1662 2460 1663 2464
rect 1667 2460 1668 2464
rect 1662 2459 1668 2460
rect 1734 2464 1740 2465
rect 1734 2460 1735 2464
rect 1739 2460 1740 2464
rect 1734 2459 1740 2460
rect 1806 2464 1812 2465
rect 1806 2460 1807 2464
rect 1811 2460 1812 2464
rect 1806 2459 1812 2460
rect 1878 2464 1884 2465
rect 1878 2460 1879 2464
rect 1883 2460 1884 2464
rect 1878 2459 1884 2460
rect 1950 2464 1956 2465
rect 1950 2460 1951 2464
rect 1955 2460 1956 2464
rect 1950 2459 1956 2460
rect 2022 2464 2028 2465
rect 2022 2460 2023 2464
rect 2027 2460 2028 2464
rect 2022 2459 2028 2460
rect 2094 2464 2100 2465
rect 2094 2460 2095 2464
rect 2099 2460 2100 2464
rect 2094 2459 2100 2460
rect 2166 2464 2172 2465
rect 2166 2460 2167 2464
rect 2171 2460 2172 2464
rect 2502 2463 2503 2467
rect 2507 2463 2508 2467
rect 2502 2462 2508 2463
rect 2166 2459 2172 2460
rect 1528 2455 1530 2459
rect 1592 2455 1594 2459
rect 1664 2455 1666 2459
rect 1736 2455 1738 2459
rect 1808 2455 1810 2459
rect 1880 2455 1882 2459
rect 1952 2455 1954 2459
rect 2024 2455 2026 2459
rect 2096 2455 2098 2459
rect 2168 2455 2170 2459
rect 2504 2455 2506 2462
rect 1327 2454 1331 2455
rect 1327 2449 1331 2450
rect 1527 2454 1531 2455
rect 1527 2449 1531 2450
rect 1543 2454 1547 2455
rect 1543 2449 1547 2450
rect 1591 2454 1595 2455
rect 1591 2449 1595 2450
rect 1607 2454 1611 2455
rect 1607 2449 1611 2450
rect 1663 2454 1667 2455
rect 1663 2449 1667 2450
rect 1671 2454 1675 2455
rect 1671 2449 1675 2450
rect 1735 2454 1739 2455
rect 1735 2449 1739 2450
rect 1743 2454 1747 2455
rect 1743 2449 1747 2450
rect 1807 2454 1811 2455
rect 1807 2449 1811 2450
rect 1815 2454 1819 2455
rect 1815 2449 1819 2450
rect 1879 2454 1883 2455
rect 1879 2449 1883 2450
rect 1951 2454 1955 2455
rect 1951 2449 1955 2450
rect 2023 2454 2027 2455
rect 2023 2449 2027 2450
rect 2095 2454 2099 2455
rect 2095 2449 2099 2450
rect 2167 2454 2171 2455
rect 2167 2449 2171 2450
rect 2503 2454 2507 2455
rect 2503 2449 2507 2450
rect 1328 2446 1330 2449
rect 1542 2448 1548 2449
rect 1326 2445 1332 2446
rect 110 2444 116 2445
rect 1286 2444 1292 2445
rect 110 2440 111 2444
rect 115 2440 116 2444
rect 110 2439 116 2440
rect 182 2443 188 2444
rect 182 2439 183 2443
rect 187 2439 188 2443
rect 112 2407 114 2439
rect 182 2438 188 2439
rect 238 2443 244 2444
rect 238 2439 239 2443
rect 243 2439 244 2443
rect 238 2438 244 2439
rect 294 2443 300 2444
rect 294 2439 295 2443
rect 299 2439 300 2443
rect 294 2438 300 2439
rect 350 2443 356 2444
rect 350 2439 351 2443
rect 355 2439 356 2443
rect 350 2438 356 2439
rect 406 2443 412 2444
rect 406 2439 407 2443
rect 411 2439 412 2443
rect 406 2438 412 2439
rect 462 2443 468 2444
rect 462 2439 463 2443
rect 467 2439 468 2443
rect 462 2438 468 2439
rect 518 2443 524 2444
rect 518 2439 519 2443
rect 523 2439 524 2443
rect 518 2438 524 2439
rect 574 2443 580 2444
rect 574 2439 575 2443
rect 579 2439 580 2443
rect 574 2438 580 2439
rect 630 2443 636 2444
rect 630 2439 631 2443
rect 635 2439 636 2443
rect 630 2438 636 2439
rect 686 2443 692 2444
rect 686 2439 687 2443
rect 691 2439 692 2443
rect 686 2438 692 2439
rect 742 2443 748 2444
rect 742 2439 743 2443
rect 747 2439 748 2443
rect 742 2438 748 2439
rect 798 2443 804 2444
rect 798 2439 799 2443
rect 803 2439 804 2443
rect 798 2438 804 2439
rect 854 2443 860 2444
rect 854 2439 855 2443
rect 859 2439 860 2443
rect 854 2438 860 2439
rect 910 2443 916 2444
rect 910 2439 911 2443
rect 915 2439 916 2443
rect 910 2438 916 2439
rect 966 2443 972 2444
rect 966 2439 967 2443
rect 971 2439 972 2443
rect 966 2438 972 2439
rect 1022 2443 1028 2444
rect 1022 2439 1023 2443
rect 1027 2439 1028 2443
rect 1022 2438 1028 2439
rect 1078 2443 1084 2444
rect 1078 2439 1079 2443
rect 1083 2439 1084 2443
rect 1286 2440 1287 2444
rect 1291 2440 1292 2444
rect 1326 2441 1327 2445
rect 1331 2441 1332 2445
rect 1542 2444 1543 2448
rect 1547 2444 1548 2448
rect 1542 2443 1548 2444
rect 1606 2448 1612 2449
rect 1606 2444 1607 2448
rect 1611 2444 1612 2448
rect 1606 2443 1612 2444
rect 1670 2448 1676 2449
rect 1670 2444 1671 2448
rect 1675 2444 1676 2448
rect 1670 2443 1676 2444
rect 1742 2448 1748 2449
rect 1742 2444 1743 2448
rect 1747 2444 1748 2448
rect 1742 2443 1748 2444
rect 1814 2448 1820 2449
rect 1814 2444 1815 2448
rect 1819 2444 1820 2448
rect 1814 2443 1820 2444
rect 1878 2448 1884 2449
rect 1878 2444 1879 2448
rect 1883 2444 1884 2448
rect 1878 2443 1884 2444
rect 1950 2448 1956 2449
rect 1950 2444 1951 2448
rect 1955 2444 1956 2448
rect 1950 2443 1956 2444
rect 2022 2448 2028 2449
rect 2022 2444 2023 2448
rect 2027 2444 2028 2448
rect 2022 2443 2028 2444
rect 2094 2448 2100 2449
rect 2094 2444 2095 2448
rect 2099 2444 2100 2448
rect 2094 2443 2100 2444
rect 2166 2448 2172 2449
rect 2166 2444 2167 2448
rect 2171 2444 2172 2448
rect 2504 2446 2506 2449
rect 2166 2443 2172 2444
rect 2502 2445 2508 2446
rect 1326 2440 1332 2441
rect 2502 2441 2503 2445
rect 2507 2441 2508 2445
rect 2502 2440 2508 2441
rect 1286 2439 1292 2440
rect 1078 2438 1084 2439
rect 184 2407 186 2438
rect 240 2407 242 2438
rect 296 2407 298 2438
rect 352 2407 354 2438
rect 408 2407 410 2438
rect 464 2407 466 2438
rect 520 2407 522 2438
rect 576 2407 578 2438
rect 632 2407 634 2438
rect 688 2407 690 2438
rect 744 2407 746 2438
rect 800 2407 802 2438
rect 856 2407 858 2438
rect 912 2407 914 2438
rect 968 2407 970 2438
rect 1024 2407 1026 2438
rect 1080 2407 1082 2438
rect 1288 2407 1290 2439
rect 1326 2428 1332 2429
rect 2502 2428 2508 2429
rect 1326 2424 1327 2428
rect 1331 2424 1332 2428
rect 1326 2423 1332 2424
rect 1558 2427 1564 2428
rect 1558 2423 1559 2427
rect 1563 2423 1564 2427
rect 111 2406 115 2407
rect 111 2401 115 2402
rect 183 2406 187 2407
rect 183 2401 187 2402
rect 239 2406 243 2407
rect 239 2401 243 2402
rect 295 2406 299 2407
rect 295 2401 299 2402
rect 351 2406 355 2407
rect 351 2401 355 2402
rect 407 2406 411 2407
rect 407 2401 411 2402
rect 463 2406 467 2407
rect 463 2401 467 2402
rect 519 2406 523 2407
rect 519 2401 523 2402
rect 575 2406 579 2407
rect 575 2401 579 2402
rect 631 2406 635 2407
rect 631 2401 635 2402
rect 687 2406 691 2407
rect 687 2401 691 2402
rect 743 2406 747 2407
rect 743 2401 747 2402
rect 799 2406 803 2407
rect 799 2401 803 2402
rect 855 2406 859 2407
rect 855 2401 859 2402
rect 911 2406 915 2407
rect 911 2401 915 2402
rect 967 2406 971 2407
rect 967 2401 971 2402
rect 1023 2406 1027 2407
rect 1023 2401 1027 2402
rect 1079 2406 1083 2407
rect 1079 2401 1083 2402
rect 1287 2406 1291 2407
rect 1287 2401 1291 2402
rect 112 2381 114 2401
rect 520 2382 522 2401
rect 576 2382 578 2401
rect 632 2382 634 2401
rect 688 2382 690 2401
rect 518 2381 524 2382
rect 110 2380 116 2381
rect 110 2376 111 2380
rect 115 2376 116 2380
rect 518 2377 519 2381
rect 523 2377 524 2381
rect 518 2376 524 2377
rect 574 2381 580 2382
rect 574 2377 575 2381
rect 579 2377 580 2381
rect 574 2376 580 2377
rect 630 2381 636 2382
rect 630 2377 631 2381
rect 635 2377 636 2381
rect 630 2376 636 2377
rect 686 2381 692 2382
rect 1288 2381 1290 2401
rect 1328 2399 1330 2423
rect 1558 2422 1564 2423
rect 1622 2427 1628 2428
rect 1622 2423 1623 2427
rect 1627 2423 1628 2427
rect 1622 2422 1628 2423
rect 1686 2427 1692 2428
rect 1686 2423 1687 2427
rect 1691 2423 1692 2427
rect 1686 2422 1692 2423
rect 1758 2427 1764 2428
rect 1758 2423 1759 2427
rect 1763 2423 1764 2427
rect 1758 2422 1764 2423
rect 1830 2427 1836 2428
rect 1830 2423 1831 2427
rect 1835 2423 1836 2427
rect 1830 2422 1836 2423
rect 1894 2427 1900 2428
rect 1894 2423 1895 2427
rect 1899 2423 1900 2427
rect 1894 2422 1900 2423
rect 1966 2427 1972 2428
rect 1966 2423 1967 2427
rect 1971 2423 1972 2427
rect 1966 2422 1972 2423
rect 2038 2427 2044 2428
rect 2038 2423 2039 2427
rect 2043 2423 2044 2427
rect 2038 2422 2044 2423
rect 2110 2427 2116 2428
rect 2110 2423 2111 2427
rect 2115 2423 2116 2427
rect 2110 2422 2116 2423
rect 2182 2427 2188 2428
rect 2182 2423 2183 2427
rect 2187 2423 2188 2427
rect 2502 2424 2503 2428
rect 2507 2424 2508 2428
rect 2502 2423 2508 2424
rect 2182 2422 2188 2423
rect 1560 2399 1562 2422
rect 1624 2399 1626 2422
rect 1688 2399 1690 2422
rect 1760 2399 1762 2422
rect 1832 2399 1834 2422
rect 1896 2399 1898 2422
rect 1968 2399 1970 2422
rect 2040 2399 2042 2422
rect 2112 2399 2114 2422
rect 2184 2399 2186 2422
rect 2504 2399 2506 2423
rect 1327 2398 1331 2399
rect 1327 2393 1331 2394
rect 1559 2398 1563 2399
rect 1559 2393 1563 2394
rect 1567 2398 1571 2399
rect 1567 2393 1571 2394
rect 1623 2398 1627 2399
rect 1623 2393 1627 2394
rect 1679 2398 1683 2399
rect 1679 2393 1683 2394
rect 1687 2398 1691 2399
rect 1687 2393 1691 2394
rect 1735 2398 1739 2399
rect 1735 2393 1739 2394
rect 1759 2398 1763 2399
rect 1759 2393 1763 2394
rect 1791 2398 1795 2399
rect 1791 2393 1795 2394
rect 1831 2398 1835 2399
rect 1831 2393 1835 2394
rect 1855 2398 1859 2399
rect 1855 2393 1859 2394
rect 1895 2398 1899 2399
rect 1895 2393 1899 2394
rect 1919 2398 1923 2399
rect 1919 2393 1923 2394
rect 1967 2398 1971 2399
rect 1967 2393 1971 2394
rect 1983 2398 1987 2399
rect 1983 2393 1987 2394
rect 2039 2398 2043 2399
rect 2039 2393 2043 2394
rect 2047 2398 2051 2399
rect 2047 2393 2051 2394
rect 2111 2398 2115 2399
rect 2111 2393 2115 2394
rect 2183 2398 2187 2399
rect 2183 2393 2187 2394
rect 2503 2398 2507 2399
rect 2503 2393 2507 2394
rect 686 2377 687 2381
rect 691 2377 692 2381
rect 686 2376 692 2377
rect 1286 2380 1292 2381
rect 1286 2376 1287 2380
rect 1291 2376 1292 2380
rect 110 2375 116 2376
rect 1286 2375 1292 2376
rect 1328 2373 1330 2393
rect 1568 2374 1570 2393
rect 1624 2374 1626 2393
rect 1680 2374 1682 2393
rect 1736 2374 1738 2393
rect 1792 2374 1794 2393
rect 1856 2374 1858 2393
rect 1920 2374 1922 2393
rect 1984 2374 1986 2393
rect 2048 2374 2050 2393
rect 2112 2374 2114 2393
rect 1566 2373 1572 2374
rect 1326 2372 1332 2373
rect 1326 2368 1327 2372
rect 1331 2368 1332 2372
rect 1566 2369 1567 2373
rect 1571 2369 1572 2373
rect 1566 2368 1572 2369
rect 1622 2373 1628 2374
rect 1622 2369 1623 2373
rect 1627 2369 1628 2373
rect 1622 2368 1628 2369
rect 1678 2373 1684 2374
rect 1678 2369 1679 2373
rect 1683 2369 1684 2373
rect 1678 2368 1684 2369
rect 1734 2373 1740 2374
rect 1734 2369 1735 2373
rect 1739 2369 1740 2373
rect 1734 2368 1740 2369
rect 1790 2373 1796 2374
rect 1790 2369 1791 2373
rect 1795 2369 1796 2373
rect 1790 2368 1796 2369
rect 1854 2373 1860 2374
rect 1854 2369 1855 2373
rect 1859 2369 1860 2373
rect 1854 2368 1860 2369
rect 1918 2373 1924 2374
rect 1918 2369 1919 2373
rect 1923 2369 1924 2373
rect 1918 2368 1924 2369
rect 1982 2373 1988 2374
rect 1982 2369 1983 2373
rect 1987 2369 1988 2373
rect 1982 2368 1988 2369
rect 2046 2373 2052 2374
rect 2046 2369 2047 2373
rect 2051 2369 2052 2373
rect 2046 2368 2052 2369
rect 2110 2373 2116 2374
rect 2504 2373 2506 2393
rect 2110 2369 2111 2373
rect 2115 2369 2116 2373
rect 2110 2368 2116 2369
rect 2502 2372 2508 2373
rect 2502 2368 2503 2372
rect 2507 2368 2508 2372
rect 1326 2367 1332 2368
rect 2502 2367 2508 2368
rect 110 2363 116 2364
rect 110 2359 111 2363
rect 115 2359 116 2363
rect 1286 2363 1292 2364
rect 110 2358 116 2359
rect 502 2360 508 2361
rect 112 2347 114 2358
rect 502 2356 503 2360
rect 507 2356 508 2360
rect 502 2355 508 2356
rect 558 2360 564 2361
rect 558 2356 559 2360
rect 563 2356 564 2360
rect 558 2355 564 2356
rect 614 2360 620 2361
rect 614 2356 615 2360
rect 619 2356 620 2360
rect 614 2355 620 2356
rect 670 2360 676 2361
rect 670 2356 671 2360
rect 675 2356 676 2360
rect 1286 2359 1287 2363
rect 1291 2359 1292 2363
rect 1286 2358 1292 2359
rect 670 2355 676 2356
rect 504 2347 506 2355
rect 560 2347 562 2355
rect 616 2347 618 2355
rect 672 2347 674 2355
rect 1288 2347 1290 2358
rect 1326 2355 1332 2356
rect 1326 2351 1327 2355
rect 1331 2351 1332 2355
rect 2502 2355 2508 2356
rect 1326 2350 1332 2351
rect 1550 2352 1556 2353
rect 111 2346 115 2347
rect 111 2341 115 2342
rect 319 2346 323 2347
rect 319 2341 323 2342
rect 391 2346 395 2347
rect 391 2341 395 2342
rect 463 2346 467 2347
rect 463 2341 467 2342
rect 503 2346 507 2347
rect 503 2341 507 2342
rect 535 2346 539 2347
rect 535 2341 539 2342
rect 559 2346 563 2347
rect 559 2341 563 2342
rect 607 2346 611 2347
rect 607 2341 611 2342
rect 615 2346 619 2347
rect 615 2341 619 2342
rect 671 2346 675 2347
rect 671 2341 675 2342
rect 679 2346 683 2347
rect 679 2341 683 2342
rect 743 2346 747 2347
rect 743 2341 747 2342
rect 807 2346 811 2347
rect 807 2341 811 2342
rect 863 2346 867 2347
rect 863 2341 867 2342
rect 927 2346 931 2347
rect 927 2341 931 2342
rect 991 2346 995 2347
rect 991 2341 995 2342
rect 1055 2346 1059 2347
rect 1055 2341 1059 2342
rect 1111 2346 1115 2347
rect 1111 2341 1115 2342
rect 1167 2346 1171 2347
rect 1167 2341 1171 2342
rect 1223 2346 1227 2347
rect 1223 2341 1227 2342
rect 1287 2346 1291 2347
rect 1287 2341 1291 2342
rect 112 2338 114 2341
rect 318 2340 324 2341
rect 110 2337 116 2338
rect 110 2333 111 2337
rect 115 2333 116 2337
rect 318 2336 319 2340
rect 323 2336 324 2340
rect 318 2335 324 2336
rect 390 2340 396 2341
rect 390 2336 391 2340
rect 395 2336 396 2340
rect 390 2335 396 2336
rect 462 2340 468 2341
rect 462 2336 463 2340
rect 467 2336 468 2340
rect 462 2335 468 2336
rect 534 2340 540 2341
rect 534 2336 535 2340
rect 539 2336 540 2340
rect 534 2335 540 2336
rect 606 2340 612 2341
rect 606 2336 607 2340
rect 611 2336 612 2340
rect 606 2335 612 2336
rect 678 2340 684 2341
rect 678 2336 679 2340
rect 683 2336 684 2340
rect 678 2335 684 2336
rect 742 2340 748 2341
rect 742 2336 743 2340
rect 747 2336 748 2340
rect 742 2335 748 2336
rect 806 2340 812 2341
rect 806 2336 807 2340
rect 811 2336 812 2340
rect 806 2335 812 2336
rect 862 2340 868 2341
rect 862 2336 863 2340
rect 867 2336 868 2340
rect 862 2335 868 2336
rect 926 2340 932 2341
rect 926 2336 927 2340
rect 931 2336 932 2340
rect 926 2335 932 2336
rect 990 2340 996 2341
rect 990 2336 991 2340
rect 995 2336 996 2340
rect 990 2335 996 2336
rect 1054 2340 1060 2341
rect 1054 2336 1055 2340
rect 1059 2336 1060 2340
rect 1054 2335 1060 2336
rect 1110 2340 1116 2341
rect 1110 2336 1111 2340
rect 1115 2336 1116 2340
rect 1110 2335 1116 2336
rect 1166 2340 1172 2341
rect 1166 2336 1167 2340
rect 1171 2336 1172 2340
rect 1166 2335 1172 2336
rect 1222 2340 1228 2341
rect 1222 2336 1223 2340
rect 1227 2336 1228 2340
rect 1288 2338 1290 2341
rect 1328 2339 1330 2350
rect 1550 2348 1551 2352
rect 1555 2348 1556 2352
rect 1550 2347 1556 2348
rect 1606 2352 1612 2353
rect 1606 2348 1607 2352
rect 1611 2348 1612 2352
rect 1606 2347 1612 2348
rect 1662 2352 1668 2353
rect 1662 2348 1663 2352
rect 1667 2348 1668 2352
rect 1662 2347 1668 2348
rect 1718 2352 1724 2353
rect 1718 2348 1719 2352
rect 1723 2348 1724 2352
rect 1718 2347 1724 2348
rect 1774 2352 1780 2353
rect 1774 2348 1775 2352
rect 1779 2348 1780 2352
rect 1774 2347 1780 2348
rect 1838 2352 1844 2353
rect 1838 2348 1839 2352
rect 1843 2348 1844 2352
rect 1838 2347 1844 2348
rect 1902 2352 1908 2353
rect 1902 2348 1903 2352
rect 1907 2348 1908 2352
rect 1902 2347 1908 2348
rect 1966 2352 1972 2353
rect 1966 2348 1967 2352
rect 1971 2348 1972 2352
rect 1966 2347 1972 2348
rect 2030 2352 2036 2353
rect 2030 2348 2031 2352
rect 2035 2348 2036 2352
rect 2030 2347 2036 2348
rect 2094 2352 2100 2353
rect 2094 2348 2095 2352
rect 2099 2348 2100 2352
rect 2502 2351 2503 2355
rect 2507 2351 2508 2355
rect 2502 2350 2508 2351
rect 2094 2347 2100 2348
rect 1552 2339 1554 2347
rect 1608 2339 1610 2347
rect 1664 2339 1666 2347
rect 1720 2339 1722 2347
rect 1776 2339 1778 2347
rect 1840 2339 1842 2347
rect 1904 2339 1906 2347
rect 1968 2339 1970 2347
rect 2032 2339 2034 2347
rect 2096 2339 2098 2347
rect 2504 2339 2506 2350
rect 1327 2338 1331 2339
rect 1222 2335 1228 2336
rect 1286 2337 1292 2338
rect 110 2332 116 2333
rect 1286 2333 1287 2337
rect 1291 2333 1292 2337
rect 1327 2333 1331 2334
rect 1471 2338 1475 2339
rect 1471 2333 1475 2334
rect 1535 2338 1539 2339
rect 1535 2333 1539 2334
rect 1551 2338 1555 2339
rect 1551 2333 1555 2334
rect 1607 2338 1611 2339
rect 1607 2333 1611 2334
rect 1663 2338 1667 2339
rect 1663 2333 1667 2334
rect 1687 2338 1691 2339
rect 1687 2333 1691 2334
rect 1719 2338 1723 2339
rect 1719 2333 1723 2334
rect 1759 2338 1763 2339
rect 1759 2333 1763 2334
rect 1775 2338 1779 2339
rect 1775 2333 1779 2334
rect 1831 2338 1835 2339
rect 1831 2333 1835 2334
rect 1839 2338 1843 2339
rect 1839 2333 1843 2334
rect 1903 2338 1907 2339
rect 1903 2333 1907 2334
rect 1967 2338 1971 2339
rect 1967 2333 1971 2334
rect 1983 2338 1987 2339
rect 1983 2333 1987 2334
rect 2031 2338 2035 2339
rect 2031 2333 2035 2334
rect 2063 2338 2067 2339
rect 2063 2333 2067 2334
rect 2095 2338 2099 2339
rect 2095 2333 2099 2334
rect 2143 2338 2147 2339
rect 2143 2333 2147 2334
rect 2503 2338 2507 2339
rect 2503 2333 2507 2334
rect 1286 2332 1292 2333
rect 1328 2330 1330 2333
rect 1470 2332 1476 2333
rect 1326 2329 1332 2330
rect 1326 2325 1327 2329
rect 1331 2325 1332 2329
rect 1470 2328 1471 2332
rect 1475 2328 1476 2332
rect 1470 2327 1476 2328
rect 1534 2332 1540 2333
rect 1534 2328 1535 2332
rect 1539 2328 1540 2332
rect 1534 2327 1540 2328
rect 1606 2332 1612 2333
rect 1606 2328 1607 2332
rect 1611 2328 1612 2332
rect 1606 2327 1612 2328
rect 1686 2332 1692 2333
rect 1686 2328 1687 2332
rect 1691 2328 1692 2332
rect 1686 2327 1692 2328
rect 1758 2332 1764 2333
rect 1758 2328 1759 2332
rect 1763 2328 1764 2332
rect 1758 2327 1764 2328
rect 1830 2332 1836 2333
rect 1830 2328 1831 2332
rect 1835 2328 1836 2332
rect 1830 2327 1836 2328
rect 1902 2332 1908 2333
rect 1902 2328 1903 2332
rect 1907 2328 1908 2332
rect 1902 2327 1908 2328
rect 1982 2332 1988 2333
rect 1982 2328 1983 2332
rect 1987 2328 1988 2332
rect 1982 2327 1988 2328
rect 2062 2332 2068 2333
rect 2062 2328 2063 2332
rect 2067 2328 2068 2332
rect 2062 2327 2068 2328
rect 2142 2332 2148 2333
rect 2142 2328 2143 2332
rect 2147 2328 2148 2332
rect 2504 2330 2506 2333
rect 2142 2327 2148 2328
rect 2502 2329 2508 2330
rect 1326 2324 1332 2325
rect 2502 2325 2503 2329
rect 2507 2325 2508 2329
rect 2502 2324 2508 2325
rect 110 2320 116 2321
rect 1286 2320 1292 2321
rect 110 2316 111 2320
rect 115 2316 116 2320
rect 110 2315 116 2316
rect 334 2319 340 2320
rect 334 2315 335 2319
rect 339 2315 340 2319
rect 112 2287 114 2315
rect 334 2314 340 2315
rect 406 2319 412 2320
rect 406 2315 407 2319
rect 411 2315 412 2319
rect 406 2314 412 2315
rect 478 2319 484 2320
rect 478 2315 479 2319
rect 483 2315 484 2319
rect 478 2314 484 2315
rect 550 2319 556 2320
rect 550 2315 551 2319
rect 555 2315 556 2319
rect 550 2314 556 2315
rect 622 2319 628 2320
rect 622 2315 623 2319
rect 627 2315 628 2319
rect 622 2314 628 2315
rect 694 2319 700 2320
rect 694 2315 695 2319
rect 699 2315 700 2319
rect 694 2314 700 2315
rect 758 2319 764 2320
rect 758 2315 759 2319
rect 763 2315 764 2319
rect 758 2314 764 2315
rect 822 2319 828 2320
rect 822 2315 823 2319
rect 827 2315 828 2319
rect 822 2314 828 2315
rect 878 2319 884 2320
rect 878 2315 879 2319
rect 883 2315 884 2319
rect 878 2314 884 2315
rect 942 2319 948 2320
rect 942 2315 943 2319
rect 947 2315 948 2319
rect 942 2314 948 2315
rect 1006 2319 1012 2320
rect 1006 2315 1007 2319
rect 1011 2315 1012 2319
rect 1006 2314 1012 2315
rect 1070 2319 1076 2320
rect 1070 2315 1071 2319
rect 1075 2315 1076 2319
rect 1070 2314 1076 2315
rect 1126 2319 1132 2320
rect 1126 2315 1127 2319
rect 1131 2315 1132 2319
rect 1126 2314 1132 2315
rect 1182 2319 1188 2320
rect 1182 2315 1183 2319
rect 1187 2315 1188 2319
rect 1182 2314 1188 2315
rect 1238 2319 1244 2320
rect 1238 2315 1239 2319
rect 1243 2315 1244 2319
rect 1286 2316 1287 2320
rect 1291 2316 1292 2320
rect 1286 2315 1292 2316
rect 1238 2314 1244 2315
rect 336 2287 338 2314
rect 408 2287 410 2314
rect 480 2287 482 2314
rect 552 2287 554 2314
rect 624 2287 626 2314
rect 696 2287 698 2314
rect 760 2287 762 2314
rect 824 2287 826 2314
rect 880 2287 882 2314
rect 944 2287 946 2314
rect 1008 2287 1010 2314
rect 1072 2287 1074 2314
rect 1128 2287 1130 2314
rect 1184 2287 1186 2314
rect 1240 2287 1242 2314
rect 1288 2287 1290 2315
rect 1326 2312 1332 2313
rect 2502 2312 2508 2313
rect 1326 2308 1327 2312
rect 1331 2308 1332 2312
rect 1326 2307 1332 2308
rect 1486 2311 1492 2312
rect 1486 2307 1487 2311
rect 1491 2307 1492 2311
rect 1328 2287 1330 2307
rect 1486 2306 1492 2307
rect 1550 2311 1556 2312
rect 1550 2307 1551 2311
rect 1555 2307 1556 2311
rect 1550 2306 1556 2307
rect 1622 2311 1628 2312
rect 1622 2307 1623 2311
rect 1627 2307 1628 2311
rect 1622 2306 1628 2307
rect 1702 2311 1708 2312
rect 1702 2307 1703 2311
rect 1707 2307 1708 2311
rect 1702 2306 1708 2307
rect 1774 2311 1780 2312
rect 1774 2307 1775 2311
rect 1779 2307 1780 2311
rect 1774 2306 1780 2307
rect 1846 2311 1852 2312
rect 1846 2307 1847 2311
rect 1851 2307 1852 2311
rect 1846 2306 1852 2307
rect 1918 2311 1924 2312
rect 1918 2307 1919 2311
rect 1923 2307 1924 2311
rect 1918 2306 1924 2307
rect 1998 2311 2004 2312
rect 1998 2307 1999 2311
rect 2003 2307 2004 2311
rect 1998 2306 2004 2307
rect 2078 2311 2084 2312
rect 2078 2307 2079 2311
rect 2083 2307 2084 2311
rect 2078 2306 2084 2307
rect 2158 2311 2164 2312
rect 2158 2307 2159 2311
rect 2163 2307 2164 2311
rect 2502 2308 2503 2312
rect 2507 2308 2508 2312
rect 2502 2307 2508 2308
rect 2158 2306 2164 2307
rect 1488 2287 1490 2306
rect 1552 2287 1554 2306
rect 1624 2287 1626 2306
rect 1704 2287 1706 2306
rect 1776 2287 1778 2306
rect 1848 2287 1850 2306
rect 1920 2287 1922 2306
rect 2000 2287 2002 2306
rect 2080 2287 2082 2306
rect 2160 2287 2162 2306
rect 2504 2287 2506 2307
rect 111 2286 115 2287
rect 111 2281 115 2282
rect 175 2286 179 2287
rect 175 2281 179 2282
rect 271 2286 275 2287
rect 271 2281 275 2282
rect 335 2286 339 2287
rect 335 2281 339 2282
rect 375 2286 379 2287
rect 375 2281 379 2282
rect 407 2286 411 2287
rect 407 2281 411 2282
rect 479 2286 483 2287
rect 479 2281 483 2282
rect 551 2286 555 2287
rect 551 2281 555 2282
rect 591 2286 595 2287
rect 591 2281 595 2282
rect 623 2286 627 2287
rect 623 2281 627 2282
rect 695 2286 699 2287
rect 695 2281 699 2282
rect 703 2286 707 2287
rect 703 2281 707 2282
rect 759 2286 763 2287
rect 759 2281 763 2282
rect 807 2286 811 2287
rect 807 2281 811 2282
rect 823 2286 827 2287
rect 823 2281 827 2282
rect 879 2286 883 2287
rect 879 2281 883 2282
rect 911 2286 915 2287
rect 911 2281 915 2282
rect 943 2286 947 2287
rect 943 2281 947 2282
rect 1007 2286 1011 2287
rect 1007 2281 1011 2282
rect 1015 2286 1019 2287
rect 1015 2281 1019 2282
rect 1071 2286 1075 2287
rect 1071 2281 1075 2282
rect 1127 2286 1131 2287
rect 1127 2281 1131 2282
rect 1183 2286 1187 2287
rect 1183 2281 1187 2282
rect 1239 2286 1243 2287
rect 1239 2281 1243 2282
rect 1287 2286 1291 2287
rect 1287 2281 1291 2282
rect 1327 2286 1331 2287
rect 1327 2281 1331 2282
rect 1383 2286 1387 2287
rect 1383 2281 1387 2282
rect 1479 2286 1483 2287
rect 1479 2281 1483 2282
rect 1487 2286 1491 2287
rect 1487 2281 1491 2282
rect 1551 2286 1555 2287
rect 1551 2281 1555 2282
rect 1583 2286 1587 2287
rect 1583 2281 1587 2282
rect 1623 2286 1627 2287
rect 1623 2281 1627 2282
rect 1687 2286 1691 2287
rect 1687 2281 1691 2282
rect 1703 2286 1707 2287
rect 1703 2281 1707 2282
rect 1775 2286 1779 2287
rect 1775 2281 1779 2282
rect 1791 2286 1795 2287
rect 1791 2281 1795 2282
rect 1847 2286 1851 2287
rect 1847 2281 1851 2282
rect 1903 2286 1907 2287
rect 1903 2281 1907 2282
rect 1919 2286 1923 2287
rect 1919 2281 1923 2282
rect 1999 2286 2003 2287
rect 1999 2281 2003 2282
rect 2015 2286 2019 2287
rect 2015 2281 2019 2282
rect 2079 2286 2083 2287
rect 2079 2281 2083 2282
rect 2127 2286 2131 2287
rect 2127 2281 2131 2282
rect 2159 2286 2163 2287
rect 2159 2281 2163 2282
rect 2239 2286 2243 2287
rect 2239 2281 2243 2282
rect 2503 2286 2507 2287
rect 2503 2281 2507 2282
rect 112 2261 114 2281
rect 176 2262 178 2281
rect 272 2262 274 2281
rect 376 2262 378 2281
rect 480 2262 482 2281
rect 592 2262 594 2281
rect 704 2262 706 2281
rect 808 2262 810 2281
rect 912 2262 914 2281
rect 1016 2262 1018 2281
rect 1128 2262 1130 2281
rect 1240 2262 1242 2281
rect 174 2261 180 2262
rect 110 2260 116 2261
rect 110 2256 111 2260
rect 115 2256 116 2260
rect 174 2257 175 2261
rect 179 2257 180 2261
rect 174 2256 180 2257
rect 270 2261 276 2262
rect 270 2257 271 2261
rect 275 2257 276 2261
rect 270 2256 276 2257
rect 374 2261 380 2262
rect 374 2257 375 2261
rect 379 2257 380 2261
rect 374 2256 380 2257
rect 478 2261 484 2262
rect 478 2257 479 2261
rect 483 2257 484 2261
rect 478 2256 484 2257
rect 590 2261 596 2262
rect 590 2257 591 2261
rect 595 2257 596 2261
rect 590 2256 596 2257
rect 702 2261 708 2262
rect 702 2257 703 2261
rect 707 2257 708 2261
rect 702 2256 708 2257
rect 806 2261 812 2262
rect 806 2257 807 2261
rect 811 2257 812 2261
rect 806 2256 812 2257
rect 910 2261 916 2262
rect 910 2257 911 2261
rect 915 2257 916 2261
rect 910 2256 916 2257
rect 1014 2261 1020 2262
rect 1014 2257 1015 2261
rect 1019 2257 1020 2261
rect 1014 2256 1020 2257
rect 1126 2261 1132 2262
rect 1126 2257 1127 2261
rect 1131 2257 1132 2261
rect 1126 2256 1132 2257
rect 1238 2261 1244 2262
rect 1288 2261 1290 2281
rect 1328 2261 1330 2281
rect 1384 2262 1386 2281
rect 1480 2262 1482 2281
rect 1584 2262 1586 2281
rect 1688 2262 1690 2281
rect 1792 2262 1794 2281
rect 1904 2262 1906 2281
rect 2016 2262 2018 2281
rect 2128 2262 2130 2281
rect 2240 2262 2242 2281
rect 1382 2261 1388 2262
rect 1238 2257 1239 2261
rect 1243 2257 1244 2261
rect 1238 2256 1244 2257
rect 1286 2260 1292 2261
rect 1286 2256 1287 2260
rect 1291 2256 1292 2260
rect 110 2255 116 2256
rect 1286 2255 1292 2256
rect 1326 2260 1332 2261
rect 1326 2256 1327 2260
rect 1331 2256 1332 2260
rect 1382 2257 1383 2261
rect 1387 2257 1388 2261
rect 1382 2256 1388 2257
rect 1478 2261 1484 2262
rect 1478 2257 1479 2261
rect 1483 2257 1484 2261
rect 1478 2256 1484 2257
rect 1582 2261 1588 2262
rect 1582 2257 1583 2261
rect 1587 2257 1588 2261
rect 1582 2256 1588 2257
rect 1686 2261 1692 2262
rect 1686 2257 1687 2261
rect 1691 2257 1692 2261
rect 1686 2256 1692 2257
rect 1790 2261 1796 2262
rect 1790 2257 1791 2261
rect 1795 2257 1796 2261
rect 1790 2256 1796 2257
rect 1902 2261 1908 2262
rect 1902 2257 1903 2261
rect 1907 2257 1908 2261
rect 1902 2256 1908 2257
rect 2014 2261 2020 2262
rect 2014 2257 2015 2261
rect 2019 2257 2020 2261
rect 2014 2256 2020 2257
rect 2126 2261 2132 2262
rect 2126 2257 2127 2261
rect 2131 2257 2132 2261
rect 2126 2256 2132 2257
rect 2238 2261 2244 2262
rect 2504 2261 2506 2281
rect 2238 2257 2239 2261
rect 2243 2257 2244 2261
rect 2238 2256 2244 2257
rect 2502 2260 2508 2261
rect 2502 2256 2503 2260
rect 2507 2256 2508 2260
rect 1326 2255 1332 2256
rect 2502 2255 2508 2256
rect 110 2243 116 2244
rect 110 2239 111 2243
rect 115 2239 116 2243
rect 1286 2243 1292 2244
rect 110 2238 116 2239
rect 158 2240 164 2241
rect 112 2235 114 2238
rect 158 2236 159 2240
rect 163 2236 164 2240
rect 158 2235 164 2236
rect 254 2240 260 2241
rect 254 2236 255 2240
rect 259 2236 260 2240
rect 254 2235 260 2236
rect 358 2240 364 2241
rect 358 2236 359 2240
rect 363 2236 364 2240
rect 358 2235 364 2236
rect 462 2240 468 2241
rect 462 2236 463 2240
rect 467 2236 468 2240
rect 462 2235 468 2236
rect 574 2240 580 2241
rect 574 2236 575 2240
rect 579 2236 580 2240
rect 574 2235 580 2236
rect 686 2240 692 2241
rect 686 2236 687 2240
rect 691 2236 692 2240
rect 686 2235 692 2236
rect 790 2240 796 2241
rect 790 2236 791 2240
rect 795 2236 796 2240
rect 790 2235 796 2236
rect 894 2240 900 2241
rect 894 2236 895 2240
rect 899 2236 900 2240
rect 894 2235 900 2236
rect 998 2240 1004 2241
rect 998 2236 999 2240
rect 1003 2236 1004 2240
rect 998 2235 1004 2236
rect 1110 2240 1116 2241
rect 1110 2236 1111 2240
rect 1115 2236 1116 2240
rect 1110 2235 1116 2236
rect 1222 2240 1228 2241
rect 1222 2236 1223 2240
rect 1227 2236 1228 2240
rect 1286 2239 1287 2243
rect 1291 2239 1292 2243
rect 1286 2238 1292 2239
rect 1326 2243 1332 2244
rect 1326 2239 1327 2243
rect 1331 2239 1332 2243
rect 2502 2243 2508 2244
rect 1326 2238 1332 2239
rect 1366 2240 1372 2241
rect 1222 2235 1228 2236
rect 1288 2235 1290 2238
rect 1328 2235 1330 2238
rect 1366 2236 1367 2240
rect 1371 2236 1372 2240
rect 1366 2235 1372 2236
rect 1462 2240 1468 2241
rect 1462 2236 1463 2240
rect 1467 2236 1468 2240
rect 1462 2235 1468 2236
rect 1566 2240 1572 2241
rect 1566 2236 1567 2240
rect 1571 2236 1572 2240
rect 1566 2235 1572 2236
rect 1670 2240 1676 2241
rect 1670 2236 1671 2240
rect 1675 2236 1676 2240
rect 1670 2235 1676 2236
rect 1774 2240 1780 2241
rect 1774 2236 1775 2240
rect 1779 2236 1780 2240
rect 1774 2235 1780 2236
rect 1886 2240 1892 2241
rect 1886 2236 1887 2240
rect 1891 2236 1892 2240
rect 1886 2235 1892 2236
rect 1998 2240 2004 2241
rect 1998 2236 1999 2240
rect 2003 2236 2004 2240
rect 1998 2235 2004 2236
rect 2110 2240 2116 2241
rect 2110 2236 2111 2240
rect 2115 2236 2116 2240
rect 2110 2235 2116 2236
rect 2222 2240 2228 2241
rect 2222 2236 2223 2240
rect 2227 2236 2228 2240
rect 2502 2239 2503 2243
rect 2507 2239 2508 2243
rect 2502 2238 2508 2239
rect 2222 2235 2228 2236
rect 2504 2235 2506 2238
rect 111 2234 115 2235
rect 111 2229 115 2230
rect 143 2234 147 2235
rect 143 2229 147 2230
rect 159 2234 163 2235
rect 159 2229 163 2230
rect 231 2234 235 2235
rect 231 2229 235 2230
rect 255 2234 259 2235
rect 255 2229 259 2230
rect 319 2234 323 2235
rect 319 2229 323 2230
rect 359 2234 363 2235
rect 359 2229 363 2230
rect 415 2234 419 2235
rect 415 2229 419 2230
rect 463 2234 467 2235
rect 463 2229 467 2230
rect 519 2234 523 2235
rect 519 2229 523 2230
rect 575 2234 579 2235
rect 575 2229 579 2230
rect 623 2234 627 2235
rect 623 2229 627 2230
rect 687 2234 691 2235
rect 687 2229 691 2230
rect 727 2234 731 2235
rect 727 2229 731 2230
rect 791 2234 795 2235
rect 791 2229 795 2230
rect 831 2234 835 2235
rect 831 2229 835 2230
rect 895 2234 899 2235
rect 895 2229 899 2230
rect 935 2234 939 2235
rect 935 2229 939 2230
rect 999 2234 1003 2235
rect 999 2229 1003 2230
rect 1039 2234 1043 2235
rect 1039 2229 1043 2230
rect 1111 2234 1115 2235
rect 1111 2229 1115 2230
rect 1143 2234 1147 2235
rect 1143 2229 1147 2230
rect 1223 2234 1227 2235
rect 1223 2229 1227 2230
rect 1287 2234 1291 2235
rect 1287 2229 1291 2230
rect 1327 2234 1331 2235
rect 1327 2229 1331 2230
rect 1367 2234 1371 2235
rect 1367 2229 1371 2230
rect 1463 2234 1467 2235
rect 1463 2229 1467 2230
rect 1487 2234 1491 2235
rect 1487 2229 1491 2230
rect 1567 2234 1571 2235
rect 1567 2229 1571 2230
rect 1607 2234 1611 2235
rect 1607 2229 1611 2230
rect 1671 2234 1675 2235
rect 1671 2229 1675 2230
rect 1719 2234 1723 2235
rect 1719 2229 1723 2230
rect 1775 2234 1779 2235
rect 1775 2229 1779 2230
rect 1815 2234 1819 2235
rect 1815 2229 1819 2230
rect 1887 2234 1891 2235
rect 1887 2229 1891 2230
rect 1903 2234 1907 2235
rect 1903 2229 1907 2230
rect 1983 2234 1987 2235
rect 1983 2229 1987 2230
rect 1999 2234 2003 2235
rect 1999 2229 2003 2230
rect 2055 2234 2059 2235
rect 2055 2229 2059 2230
rect 2111 2234 2115 2235
rect 2111 2229 2115 2230
rect 2127 2234 2131 2235
rect 2127 2229 2131 2230
rect 2191 2234 2195 2235
rect 2191 2229 2195 2230
rect 2223 2234 2227 2235
rect 2223 2229 2227 2230
rect 2255 2234 2259 2235
rect 2255 2229 2259 2230
rect 2319 2234 2323 2235
rect 2319 2229 2323 2230
rect 2383 2234 2387 2235
rect 2383 2229 2387 2230
rect 2439 2234 2443 2235
rect 2439 2229 2443 2230
rect 2503 2234 2507 2235
rect 2503 2229 2507 2230
rect 112 2226 114 2229
rect 142 2228 148 2229
rect 110 2225 116 2226
rect 110 2221 111 2225
rect 115 2221 116 2225
rect 142 2224 143 2228
rect 147 2224 148 2228
rect 142 2223 148 2224
rect 230 2228 236 2229
rect 230 2224 231 2228
rect 235 2224 236 2228
rect 230 2223 236 2224
rect 318 2228 324 2229
rect 318 2224 319 2228
rect 323 2224 324 2228
rect 318 2223 324 2224
rect 414 2228 420 2229
rect 414 2224 415 2228
rect 419 2224 420 2228
rect 414 2223 420 2224
rect 518 2228 524 2229
rect 518 2224 519 2228
rect 523 2224 524 2228
rect 518 2223 524 2224
rect 622 2228 628 2229
rect 622 2224 623 2228
rect 627 2224 628 2228
rect 622 2223 628 2224
rect 726 2228 732 2229
rect 726 2224 727 2228
rect 731 2224 732 2228
rect 726 2223 732 2224
rect 830 2228 836 2229
rect 830 2224 831 2228
rect 835 2224 836 2228
rect 830 2223 836 2224
rect 934 2228 940 2229
rect 934 2224 935 2228
rect 939 2224 940 2228
rect 934 2223 940 2224
rect 1038 2228 1044 2229
rect 1038 2224 1039 2228
rect 1043 2224 1044 2228
rect 1038 2223 1044 2224
rect 1142 2228 1148 2229
rect 1142 2224 1143 2228
rect 1147 2224 1148 2228
rect 1142 2223 1148 2224
rect 1222 2228 1228 2229
rect 1222 2224 1223 2228
rect 1227 2224 1228 2228
rect 1288 2226 1290 2229
rect 1328 2226 1330 2229
rect 1366 2228 1372 2229
rect 1222 2223 1228 2224
rect 1286 2225 1292 2226
rect 110 2220 116 2221
rect 1286 2221 1287 2225
rect 1291 2221 1292 2225
rect 1286 2220 1292 2221
rect 1326 2225 1332 2226
rect 1326 2221 1327 2225
rect 1331 2221 1332 2225
rect 1366 2224 1367 2228
rect 1371 2224 1372 2228
rect 1366 2223 1372 2224
rect 1486 2228 1492 2229
rect 1486 2224 1487 2228
rect 1491 2224 1492 2228
rect 1486 2223 1492 2224
rect 1606 2228 1612 2229
rect 1606 2224 1607 2228
rect 1611 2224 1612 2228
rect 1606 2223 1612 2224
rect 1718 2228 1724 2229
rect 1718 2224 1719 2228
rect 1723 2224 1724 2228
rect 1718 2223 1724 2224
rect 1814 2228 1820 2229
rect 1814 2224 1815 2228
rect 1819 2224 1820 2228
rect 1814 2223 1820 2224
rect 1902 2228 1908 2229
rect 1902 2224 1903 2228
rect 1907 2224 1908 2228
rect 1902 2223 1908 2224
rect 1982 2228 1988 2229
rect 1982 2224 1983 2228
rect 1987 2224 1988 2228
rect 1982 2223 1988 2224
rect 2054 2228 2060 2229
rect 2054 2224 2055 2228
rect 2059 2224 2060 2228
rect 2054 2223 2060 2224
rect 2126 2228 2132 2229
rect 2126 2224 2127 2228
rect 2131 2224 2132 2228
rect 2126 2223 2132 2224
rect 2190 2228 2196 2229
rect 2190 2224 2191 2228
rect 2195 2224 2196 2228
rect 2190 2223 2196 2224
rect 2254 2228 2260 2229
rect 2254 2224 2255 2228
rect 2259 2224 2260 2228
rect 2254 2223 2260 2224
rect 2318 2228 2324 2229
rect 2318 2224 2319 2228
rect 2323 2224 2324 2228
rect 2318 2223 2324 2224
rect 2382 2228 2388 2229
rect 2382 2224 2383 2228
rect 2387 2224 2388 2228
rect 2382 2223 2388 2224
rect 2438 2228 2444 2229
rect 2438 2224 2439 2228
rect 2443 2224 2444 2228
rect 2504 2226 2506 2229
rect 2438 2223 2444 2224
rect 2502 2225 2508 2226
rect 1326 2220 1332 2221
rect 2502 2221 2503 2225
rect 2507 2221 2508 2225
rect 2502 2220 2508 2221
rect 110 2208 116 2209
rect 1286 2208 1292 2209
rect 110 2204 111 2208
rect 115 2204 116 2208
rect 110 2203 116 2204
rect 158 2207 164 2208
rect 158 2203 159 2207
rect 163 2203 164 2207
rect 112 2183 114 2203
rect 158 2202 164 2203
rect 246 2207 252 2208
rect 246 2203 247 2207
rect 251 2203 252 2207
rect 246 2202 252 2203
rect 334 2207 340 2208
rect 334 2203 335 2207
rect 339 2203 340 2207
rect 334 2202 340 2203
rect 430 2207 436 2208
rect 430 2203 431 2207
rect 435 2203 436 2207
rect 430 2202 436 2203
rect 534 2207 540 2208
rect 534 2203 535 2207
rect 539 2203 540 2207
rect 534 2202 540 2203
rect 638 2207 644 2208
rect 638 2203 639 2207
rect 643 2203 644 2207
rect 638 2202 644 2203
rect 742 2207 748 2208
rect 742 2203 743 2207
rect 747 2203 748 2207
rect 742 2202 748 2203
rect 846 2207 852 2208
rect 846 2203 847 2207
rect 851 2203 852 2207
rect 846 2202 852 2203
rect 950 2207 956 2208
rect 950 2203 951 2207
rect 955 2203 956 2207
rect 950 2202 956 2203
rect 1054 2207 1060 2208
rect 1054 2203 1055 2207
rect 1059 2203 1060 2207
rect 1054 2202 1060 2203
rect 1158 2207 1164 2208
rect 1158 2203 1159 2207
rect 1163 2203 1164 2207
rect 1158 2202 1164 2203
rect 1238 2207 1244 2208
rect 1238 2203 1239 2207
rect 1243 2203 1244 2207
rect 1286 2204 1287 2208
rect 1291 2204 1292 2208
rect 1286 2203 1292 2204
rect 1326 2208 1332 2209
rect 2502 2208 2508 2209
rect 1326 2204 1327 2208
rect 1331 2204 1332 2208
rect 1326 2203 1332 2204
rect 1382 2207 1388 2208
rect 1382 2203 1383 2207
rect 1387 2203 1388 2207
rect 1238 2202 1244 2203
rect 160 2183 162 2202
rect 248 2183 250 2202
rect 336 2183 338 2202
rect 432 2183 434 2202
rect 536 2183 538 2202
rect 640 2183 642 2202
rect 744 2183 746 2202
rect 848 2183 850 2202
rect 952 2183 954 2202
rect 1056 2183 1058 2202
rect 1160 2183 1162 2202
rect 1240 2183 1242 2202
rect 1288 2183 1290 2203
rect 111 2182 115 2183
rect 111 2177 115 2178
rect 159 2182 163 2183
rect 159 2177 163 2178
rect 247 2182 251 2183
rect 247 2177 251 2178
rect 255 2182 259 2183
rect 255 2177 259 2178
rect 335 2182 339 2183
rect 335 2177 339 2178
rect 351 2182 355 2183
rect 351 2177 355 2178
rect 431 2182 435 2183
rect 431 2177 435 2178
rect 455 2182 459 2183
rect 455 2177 459 2178
rect 535 2182 539 2183
rect 535 2177 539 2178
rect 559 2182 563 2183
rect 559 2177 563 2178
rect 639 2182 643 2183
rect 639 2177 643 2178
rect 663 2182 667 2183
rect 663 2177 667 2178
rect 743 2182 747 2183
rect 743 2177 747 2178
rect 767 2182 771 2183
rect 767 2177 771 2178
rect 847 2182 851 2183
rect 847 2177 851 2178
rect 863 2182 867 2183
rect 863 2177 867 2178
rect 951 2182 955 2183
rect 951 2177 955 2178
rect 959 2182 963 2183
rect 959 2177 963 2178
rect 1055 2182 1059 2183
rect 1055 2177 1059 2178
rect 1159 2182 1163 2183
rect 1159 2177 1163 2178
rect 1239 2182 1243 2183
rect 1239 2177 1243 2178
rect 1287 2182 1291 2183
rect 1287 2177 1291 2178
rect 112 2157 114 2177
rect 256 2158 258 2177
rect 352 2158 354 2177
rect 456 2158 458 2177
rect 560 2158 562 2177
rect 664 2158 666 2177
rect 768 2158 770 2177
rect 864 2158 866 2177
rect 960 2158 962 2177
rect 1056 2158 1058 2177
rect 1160 2158 1162 2177
rect 1240 2158 1242 2177
rect 254 2157 260 2158
rect 110 2156 116 2157
rect 110 2152 111 2156
rect 115 2152 116 2156
rect 254 2153 255 2157
rect 259 2153 260 2157
rect 254 2152 260 2153
rect 350 2157 356 2158
rect 350 2153 351 2157
rect 355 2153 356 2157
rect 350 2152 356 2153
rect 454 2157 460 2158
rect 454 2153 455 2157
rect 459 2153 460 2157
rect 454 2152 460 2153
rect 558 2157 564 2158
rect 558 2153 559 2157
rect 563 2153 564 2157
rect 558 2152 564 2153
rect 662 2157 668 2158
rect 662 2153 663 2157
rect 667 2153 668 2157
rect 662 2152 668 2153
rect 766 2157 772 2158
rect 766 2153 767 2157
rect 771 2153 772 2157
rect 766 2152 772 2153
rect 862 2157 868 2158
rect 862 2153 863 2157
rect 867 2153 868 2157
rect 862 2152 868 2153
rect 958 2157 964 2158
rect 958 2153 959 2157
rect 963 2153 964 2157
rect 958 2152 964 2153
rect 1054 2157 1060 2158
rect 1054 2153 1055 2157
rect 1059 2153 1060 2157
rect 1054 2152 1060 2153
rect 1158 2157 1164 2158
rect 1158 2153 1159 2157
rect 1163 2153 1164 2157
rect 1158 2152 1164 2153
rect 1238 2157 1244 2158
rect 1288 2157 1290 2177
rect 1328 2163 1330 2203
rect 1382 2202 1388 2203
rect 1502 2207 1508 2208
rect 1502 2203 1503 2207
rect 1507 2203 1508 2207
rect 1502 2202 1508 2203
rect 1622 2207 1628 2208
rect 1622 2203 1623 2207
rect 1627 2203 1628 2207
rect 1622 2202 1628 2203
rect 1734 2207 1740 2208
rect 1734 2203 1735 2207
rect 1739 2203 1740 2207
rect 1734 2202 1740 2203
rect 1830 2207 1836 2208
rect 1830 2203 1831 2207
rect 1835 2203 1836 2207
rect 1830 2202 1836 2203
rect 1918 2207 1924 2208
rect 1918 2203 1919 2207
rect 1923 2203 1924 2207
rect 1918 2202 1924 2203
rect 1998 2207 2004 2208
rect 1998 2203 1999 2207
rect 2003 2203 2004 2207
rect 1998 2202 2004 2203
rect 2070 2207 2076 2208
rect 2070 2203 2071 2207
rect 2075 2203 2076 2207
rect 2070 2202 2076 2203
rect 2142 2207 2148 2208
rect 2142 2203 2143 2207
rect 2147 2203 2148 2207
rect 2142 2202 2148 2203
rect 2206 2207 2212 2208
rect 2206 2203 2207 2207
rect 2211 2203 2212 2207
rect 2206 2202 2212 2203
rect 2270 2207 2276 2208
rect 2270 2203 2271 2207
rect 2275 2203 2276 2207
rect 2270 2202 2276 2203
rect 2334 2207 2340 2208
rect 2334 2203 2335 2207
rect 2339 2203 2340 2207
rect 2334 2202 2340 2203
rect 2398 2207 2404 2208
rect 2398 2203 2399 2207
rect 2403 2203 2404 2207
rect 2398 2202 2404 2203
rect 2454 2207 2460 2208
rect 2454 2203 2455 2207
rect 2459 2203 2460 2207
rect 2502 2204 2503 2208
rect 2507 2204 2508 2208
rect 2502 2203 2508 2204
rect 2454 2202 2460 2203
rect 1384 2163 1386 2202
rect 1504 2163 1506 2202
rect 1624 2163 1626 2202
rect 1736 2163 1738 2202
rect 1832 2163 1834 2202
rect 1920 2163 1922 2202
rect 2000 2163 2002 2202
rect 2072 2163 2074 2202
rect 2144 2163 2146 2202
rect 2208 2163 2210 2202
rect 2272 2163 2274 2202
rect 2336 2163 2338 2202
rect 2400 2163 2402 2202
rect 2456 2163 2458 2202
rect 2504 2163 2506 2203
rect 1327 2162 1331 2163
rect 1327 2157 1331 2158
rect 1383 2162 1387 2163
rect 1383 2157 1387 2158
rect 1407 2162 1411 2163
rect 1407 2157 1411 2158
rect 1503 2162 1507 2163
rect 1503 2157 1507 2158
rect 1623 2162 1627 2163
rect 1623 2157 1627 2158
rect 1735 2162 1739 2163
rect 1735 2157 1739 2158
rect 1815 2162 1819 2163
rect 1815 2157 1819 2158
rect 1831 2162 1835 2163
rect 1831 2157 1835 2158
rect 1919 2162 1923 2163
rect 1919 2157 1923 2158
rect 1991 2162 1995 2163
rect 1991 2157 1995 2158
rect 1999 2162 2003 2163
rect 1999 2157 2003 2158
rect 2071 2162 2075 2163
rect 2071 2157 2075 2158
rect 2143 2162 2147 2163
rect 2143 2157 2147 2158
rect 2159 2162 2163 2163
rect 2159 2157 2163 2158
rect 2207 2162 2211 2163
rect 2207 2157 2211 2158
rect 2271 2162 2275 2163
rect 2271 2157 2275 2158
rect 2319 2162 2323 2163
rect 2319 2157 2323 2158
rect 2335 2162 2339 2163
rect 2335 2157 2339 2158
rect 2399 2162 2403 2163
rect 2399 2157 2403 2158
rect 2455 2162 2459 2163
rect 2455 2157 2459 2158
rect 2503 2162 2507 2163
rect 2503 2157 2507 2158
rect 1238 2153 1239 2157
rect 1243 2153 1244 2157
rect 1238 2152 1244 2153
rect 1286 2156 1292 2157
rect 1286 2152 1287 2156
rect 1291 2152 1292 2156
rect 110 2151 116 2152
rect 1286 2151 1292 2152
rect 110 2139 116 2140
rect 110 2135 111 2139
rect 115 2135 116 2139
rect 1286 2139 1292 2140
rect 110 2134 116 2135
rect 238 2136 244 2137
rect 112 2131 114 2134
rect 238 2132 239 2136
rect 243 2132 244 2136
rect 238 2131 244 2132
rect 334 2136 340 2137
rect 334 2132 335 2136
rect 339 2132 340 2136
rect 334 2131 340 2132
rect 438 2136 444 2137
rect 438 2132 439 2136
rect 443 2132 444 2136
rect 438 2131 444 2132
rect 542 2136 548 2137
rect 542 2132 543 2136
rect 547 2132 548 2136
rect 542 2131 548 2132
rect 646 2136 652 2137
rect 646 2132 647 2136
rect 651 2132 652 2136
rect 646 2131 652 2132
rect 750 2136 756 2137
rect 750 2132 751 2136
rect 755 2132 756 2136
rect 750 2131 756 2132
rect 846 2136 852 2137
rect 846 2132 847 2136
rect 851 2132 852 2136
rect 846 2131 852 2132
rect 942 2136 948 2137
rect 942 2132 943 2136
rect 947 2132 948 2136
rect 942 2131 948 2132
rect 1038 2136 1044 2137
rect 1038 2132 1039 2136
rect 1043 2132 1044 2136
rect 1038 2131 1044 2132
rect 1142 2136 1148 2137
rect 1142 2132 1143 2136
rect 1147 2132 1148 2136
rect 1142 2131 1148 2132
rect 1222 2136 1228 2137
rect 1222 2132 1223 2136
rect 1227 2132 1228 2136
rect 1286 2135 1287 2139
rect 1291 2135 1292 2139
rect 1328 2137 1330 2157
rect 1408 2138 1410 2157
rect 1624 2138 1626 2157
rect 1816 2138 1818 2157
rect 1992 2138 1994 2157
rect 2160 2138 2162 2157
rect 2320 2138 2322 2157
rect 2456 2138 2458 2157
rect 1406 2137 1412 2138
rect 1286 2134 1292 2135
rect 1326 2136 1332 2137
rect 1222 2131 1228 2132
rect 1288 2131 1290 2134
rect 1326 2132 1327 2136
rect 1331 2132 1332 2136
rect 1406 2133 1407 2137
rect 1411 2133 1412 2137
rect 1406 2132 1412 2133
rect 1622 2137 1628 2138
rect 1622 2133 1623 2137
rect 1627 2133 1628 2137
rect 1622 2132 1628 2133
rect 1814 2137 1820 2138
rect 1814 2133 1815 2137
rect 1819 2133 1820 2137
rect 1814 2132 1820 2133
rect 1990 2137 1996 2138
rect 1990 2133 1991 2137
rect 1995 2133 1996 2137
rect 1990 2132 1996 2133
rect 2158 2137 2164 2138
rect 2158 2133 2159 2137
rect 2163 2133 2164 2137
rect 2158 2132 2164 2133
rect 2318 2137 2324 2138
rect 2318 2133 2319 2137
rect 2323 2133 2324 2137
rect 2318 2132 2324 2133
rect 2454 2137 2460 2138
rect 2504 2137 2506 2157
rect 2454 2133 2455 2137
rect 2459 2133 2460 2137
rect 2454 2132 2460 2133
rect 2502 2136 2508 2137
rect 2502 2132 2503 2136
rect 2507 2132 2508 2136
rect 1326 2131 1332 2132
rect 2502 2131 2508 2132
rect 111 2130 115 2131
rect 111 2125 115 2126
rect 239 2130 243 2131
rect 239 2125 243 2126
rect 303 2130 307 2131
rect 303 2125 307 2126
rect 335 2130 339 2131
rect 335 2125 339 2126
rect 359 2130 363 2131
rect 359 2125 363 2126
rect 423 2130 427 2131
rect 423 2125 427 2126
rect 439 2130 443 2131
rect 439 2125 443 2126
rect 487 2130 491 2131
rect 487 2125 491 2126
rect 543 2130 547 2131
rect 543 2125 547 2126
rect 559 2130 563 2131
rect 559 2125 563 2126
rect 631 2130 635 2131
rect 631 2125 635 2126
rect 647 2130 651 2131
rect 647 2125 651 2126
rect 711 2130 715 2131
rect 711 2125 715 2126
rect 751 2130 755 2131
rect 751 2125 755 2126
rect 799 2130 803 2131
rect 799 2125 803 2126
rect 847 2130 851 2131
rect 847 2125 851 2126
rect 887 2130 891 2131
rect 887 2125 891 2126
rect 943 2130 947 2131
rect 943 2125 947 2126
rect 975 2130 979 2131
rect 975 2125 979 2126
rect 1039 2130 1043 2131
rect 1039 2125 1043 2126
rect 1063 2130 1067 2131
rect 1063 2125 1067 2126
rect 1143 2130 1147 2131
rect 1143 2125 1147 2126
rect 1151 2130 1155 2131
rect 1151 2125 1155 2126
rect 1223 2130 1227 2131
rect 1223 2125 1227 2126
rect 1287 2130 1291 2131
rect 1287 2125 1291 2126
rect 112 2122 114 2125
rect 302 2124 308 2125
rect 110 2121 116 2122
rect 110 2117 111 2121
rect 115 2117 116 2121
rect 302 2120 303 2124
rect 307 2120 308 2124
rect 302 2119 308 2120
rect 358 2124 364 2125
rect 358 2120 359 2124
rect 363 2120 364 2124
rect 358 2119 364 2120
rect 422 2124 428 2125
rect 422 2120 423 2124
rect 427 2120 428 2124
rect 422 2119 428 2120
rect 486 2124 492 2125
rect 486 2120 487 2124
rect 491 2120 492 2124
rect 486 2119 492 2120
rect 558 2124 564 2125
rect 558 2120 559 2124
rect 563 2120 564 2124
rect 558 2119 564 2120
rect 630 2124 636 2125
rect 630 2120 631 2124
rect 635 2120 636 2124
rect 630 2119 636 2120
rect 710 2124 716 2125
rect 710 2120 711 2124
rect 715 2120 716 2124
rect 710 2119 716 2120
rect 798 2124 804 2125
rect 798 2120 799 2124
rect 803 2120 804 2124
rect 798 2119 804 2120
rect 886 2124 892 2125
rect 886 2120 887 2124
rect 891 2120 892 2124
rect 886 2119 892 2120
rect 974 2124 980 2125
rect 974 2120 975 2124
rect 979 2120 980 2124
rect 974 2119 980 2120
rect 1062 2124 1068 2125
rect 1062 2120 1063 2124
rect 1067 2120 1068 2124
rect 1062 2119 1068 2120
rect 1150 2124 1156 2125
rect 1150 2120 1151 2124
rect 1155 2120 1156 2124
rect 1150 2119 1156 2120
rect 1222 2124 1228 2125
rect 1222 2120 1223 2124
rect 1227 2120 1228 2124
rect 1288 2122 1290 2125
rect 1222 2119 1228 2120
rect 1286 2121 1292 2122
rect 110 2116 116 2117
rect 1286 2117 1287 2121
rect 1291 2117 1292 2121
rect 1286 2116 1292 2117
rect 1326 2119 1332 2120
rect 1326 2115 1327 2119
rect 1331 2115 1332 2119
rect 2502 2119 2508 2120
rect 1326 2114 1332 2115
rect 1390 2116 1396 2117
rect 1328 2111 1330 2114
rect 1390 2112 1391 2116
rect 1395 2112 1396 2116
rect 1390 2111 1396 2112
rect 1606 2116 1612 2117
rect 1606 2112 1607 2116
rect 1611 2112 1612 2116
rect 1606 2111 1612 2112
rect 1798 2116 1804 2117
rect 1798 2112 1799 2116
rect 1803 2112 1804 2116
rect 1798 2111 1804 2112
rect 1974 2116 1980 2117
rect 1974 2112 1975 2116
rect 1979 2112 1980 2116
rect 1974 2111 1980 2112
rect 2142 2116 2148 2117
rect 2142 2112 2143 2116
rect 2147 2112 2148 2116
rect 2142 2111 2148 2112
rect 2302 2116 2308 2117
rect 2302 2112 2303 2116
rect 2307 2112 2308 2116
rect 2302 2111 2308 2112
rect 2438 2116 2444 2117
rect 2438 2112 2439 2116
rect 2443 2112 2444 2116
rect 2502 2115 2503 2119
rect 2507 2115 2508 2119
rect 2502 2114 2508 2115
rect 2438 2111 2444 2112
rect 2504 2111 2506 2114
rect 1327 2110 1331 2111
rect 1327 2105 1331 2106
rect 1383 2110 1387 2111
rect 1383 2105 1387 2106
rect 1391 2110 1395 2111
rect 1391 2105 1395 2106
rect 1551 2110 1555 2111
rect 1551 2105 1555 2106
rect 1607 2110 1611 2111
rect 1607 2105 1611 2106
rect 1711 2110 1715 2111
rect 1711 2105 1715 2106
rect 1799 2110 1803 2111
rect 1799 2105 1803 2106
rect 1855 2110 1859 2111
rect 1855 2105 1859 2106
rect 1975 2110 1979 2111
rect 1975 2105 1979 2106
rect 1991 2110 1995 2111
rect 1991 2105 1995 2106
rect 2119 2110 2123 2111
rect 2119 2105 2123 2106
rect 2143 2110 2147 2111
rect 2143 2105 2147 2106
rect 2239 2110 2243 2111
rect 2239 2105 2243 2106
rect 2303 2110 2307 2111
rect 2303 2105 2307 2106
rect 2367 2110 2371 2111
rect 2367 2105 2371 2106
rect 2439 2110 2443 2111
rect 2439 2105 2443 2106
rect 2503 2110 2507 2111
rect 2503 2105 2507 2106
rect 110 2104 116 2105
rect 1286 2104 1292 2105
rect 110 2100 111 2104
rect 115 2100 116 2104
rect 110 2099 116 2100
rect 318 2103 324 2104
rect 318 2099 319 2103
rect 323 2099 324 2103
rect 112 2075 114 2099
rect 318 2098 324 2099
rect 374 2103 380 2104
rect 374 2099 375 2103
rect 379 2099 380 2103
rect 374 2098 380 2099
rect 438 2103 444 2104
rect 438 2099 439 2103
rect 443 2099 444 2103
rect 438 2098 444 2099
rect 502 2103 508 2104
rect 502 2099 503 2103
rect 507 2099 508 2103
rect 502 2098 508 2099
rect 574 2103 580 2104
rect 574 2099 575 2103
rect 579 2099 580 2103
rect 574 2098 580 2099
rect 646 2103 652 2104
rect 646 2099 647 2103
rect 651 2099 652 2103
rect 646 2098 652 2099
rect 726 2103 732 2104
rect 726 2099 727 2103
rect 731 2099 732 2103
rect 726 2098 732 2099
rect 814 2103 820 2104
rect 814 2099 815 2103
rect 819 2099 820 2103
rect 814 2098 820 2099
rect 902 2103 908 2104
rect 902 2099 903 2103
rect 907 2099 908 2103
rect 902 2098 908 2099
rect 990 2103 996 2104
rect 990 2099 991 2103
rect 995 2099 996 2103
rect 990 2098 996 2099
rect 1078 2103 1084 2104
rect 1078 2099 1079 2103
rect 1083 2099 1084 2103
rect 1078 2098 1084 2099
rect 1166 2103 1172 2104
rect 1166 2099 1167 2103
rect 1171 2099 1172 2103
rect 1166 2098 1172 2099
rect 1238 2103 1244 2104
rect 1238 2099 1239 2103
rect 1243 2099 1244 2103
rect 1286 2100 1287 2104
rect 1291 2100 1292 2104
rect 1328 2102 1330 2105
rect 1382 2104 1388 2105
rect 1286 2099 1292 2100
rect 1326 2101 1332 2102
rect 1238 2098 1244 2099
rect 320 2075 322 2098
rect 376 2075 378 2098
rect 440 2075 442 2098
rect 504 2075 506 2098
rect 576 2075 578 2098
rect 648 2075 650 2098
rect 728 2075 730 2098
rect 816 2075 818 2098
rect 904 2075 906 2098
rect 992 2075 994 2098
rect 1080 2075 1082 2098
rect 1168 2075 1170 2098
rect 1240 2075 1242 2098
rect 1288 2075 1290 2099
rect 1326 2097 1327 2101
rect 1331 2097 1332 2101
rect 1382 2100 1383 2104
rect 1387 2100 1388 2104
rect 1382 2099 1388 2100
rect 1550 2104 1556 2105
rect 1550 2100 1551 2104
rect 1555 2100 1556 2104
rect 1550 2099 1556 2100
rect 1710 2104 1716 2105
rect 1710 2100 1711 2104
rect 1715 2100 1716 2104
rect 1710 2099 1716 2100
rect 1854 2104 1860 2105
rect 1854 2100 1855 2104
rect 1859 2100 1860 2104
rect 1854 2099 1860 2100
rect 1990 2104 1996 2105
rect 1990 2100 1991 2104
rect 1995 2100 1996 2104
rect 1990 2099 1996 2100
rect 2118 2104 2124 2105
rect 2118 2100 2119 2104
rect 2123 2100 2124 2104
rect 2118 2099 2124 2100
rect 2238 2104 2244 2105
rect 2238 2100 2239 2104
rect 2243 2100 2244 2104
rect 2238 2099 2244 2100
rect 2366 2104 2372 2105
rect 2366 2100 2367 2104
rect 2371 2100 2372 2104
rect 2504 2102 2506 2105
rect 2366 2099 2372 2100
rect 2502 2101 2508 2102
rect 1326 2096 1332 2097
rect 2502 2097 2503 2101
rect 2507 2097 2508 2101
rect 2502 2096 2508 2097
rect 1326 2084 1332 2085
rect 2502 2084 2508 2085
rect 1326 2080 1327 2084
rect 1331 2080 1332 2084
rect 1326 2079 1332 2080
rect 1398 2083 1404 2084
rect 1398 2079 1399 2083
rect 1403 2079 1404 2083
rect 111 2074 115 2075
rect 111 2069 115 2070
rect 319 2074 323 2075
rect 319 2069 323 2070
rect 375 2074 379 2075
rect 375 2069 379 2070
rect 399 2074 403 2075
rect 399 2069 403 2070
rect 439 2074 443 2075
rect 439 2069 443 2070
rect 455 2074 459 2075
rect 455 2069 459 2070
rect 503 2074 507 2075
rect 503 2069 507 2070
rect 511 2074 515 2075
rect 511 2069 515 2070
rect 575 2074 579 2075
rect 575 2069 579 2070
rect 639 2074 643 2075
rect 639 2069 643 2070
rect 647 2074 651 2075
rect 647 2069 651 2070
rect 711 2074 715 2075
rect 711 2069 715 2070
rect 727 2074 731 2075
rect 727 2069 731 2070
rect 791 2074 795 2075
rect 791 2069 795 2070
rect 815 2074 819 2075
rect 815 2069 819 2070
rect 863 2074 867 2075
rect 863 2069 867 2070
rect 903 2074 907 2075
rect 903 2069 907 2070
rect 943 2074 947 2075
rect 943 2069 947 2070
rect 991 2074 995 2075
rect 991 2069 995 2070
rect 1023 2074 1027 2075
rect 1023 2069 1027 2070
rect 1079 2074 1083 2075
rect 1079 2069 1083 2070
rect 1103 2074 1107 2075
rect 1103 2069 1107 2070
rect 1167 2074 1171 2075
rect 1167 2069 1171 2070
rect 1183 2074 1187 2075
rect 1183 2069 1187 2070
rect 1239 2074 1243 2075
rect 1239 2069 1243 2070
rect 1287 2074 1291 2075
rect 1287 2069 1291 2070
rect 112 2049 114 2069
rect 400 2050 402 2069
rect 456 2050 458 2069
rect 512 2050 514 2069
rect 576 2050 578 2069
rect 640 2050 642 2069
rect 712 2050 714 2069
rect 792 2050 794 2069
rect 864 2050 866 2069
rect 944 2050 946 2069
rect 1024 2050 1026 2069
rect 1104 2050 1106 2069
rect 1184 2050 1186 2069
rect 1240 2050 1242 2069
rect 398 2049 404 2050
rect 110 2048 116 2049
rect 110 2044 111 2048
rect 115 2044 116 2048
rect 398 2045 399 2049
rect 403 2045 404 2049
rect 398 2044 404 2045
rect 454 2049 460 2050
rect 454 2045 455 2049
rect 459 2045 460 2049
rect 454 2044 460 2045
rect 510 2049 516 2050
rect 510 2045 511 2049
rect 515 2045 516 2049
rect 510 2044 516 2045
rect 574 2049 580 2050
rect 574 2045 575 2049
rect 579 2045 580 2049
rect 574 2044 580 2045
rect 638 2049 644 2050
rect 638 2045 639 2049
rect 643 2045 644 2049
rect 638 2044 644 2045
rect 710 2049 716 2050
rect 710 2045 711 2049
rect 715 2045 716 2049
rect 710 2044 716 2045
rect 790 2049 796 2050
rect 790 2045 791 2049
rect 795 2045 796 2049
rect 790 2044 796 2045
rect 862 2049 868 2050
rect 862 2045 863 2049
rect 867 2045 868 2049
rect 862 2044 868 2045
rect 942 2049 948 2050
rect 942 2045 943 2049
rect 947 2045 948 2049
rect 942 2044 948 2045
rect 1022 2049 1028 2050
rect 1022 2045 1023 2049
rect 1027 2045 1028 2049
rect 1022 2044 1028 2045
rect 1102 2049 1108 2050
rect 1102 2045 1103 2049
rect 1107 2045 1108 2049
rect 1102 2044 1108 2045
rect 1182 2049 1188 2050
rect 1182 2045 1183 2049
rect 1187 2045 1188 2049
rect 1182 2044 1188 2045
rect 1238 2049 1244 2050
rect 1288 2049 1290 2069
rect 1328 2055 1330 2079
rect 1398 2078 1404 2079
rect 1566 2083 1572 2084
rect 1566 2079 1567 2083
rect 1571 2079 1572 2083
rect 1566 2078 1572 2079
rect 1726 2083 1732 2084
rect 1726 2079 1727 2083
rect 1731 2079 1732 2083
rect 1726 2078 1732 2079
rect 1870 2083 1876 2084
rect 1870 2079 1871 2083
rect 1875 2079 1876 2083
rect 1870 2078 1876 2079
rect 2006 2083 2012 2084
rect 2006 2079 2007 2083
rect 2011 2079 2012 2083
rect 2006 2078 2012 2079
rect 2134 2083 2140 2084
rect 2134 2079 2135 2083
rect 2139 2079 2140 2083
rect 2134 2078 2140 2079
rect 2254 2083 2260 2084
rect 2254 2079 2255 2083
rect 2259 2079 2260 2083
rect 2254 2078 2260 2079
rect 2382 2083 2388 2084
rect 2382 2079 2383 2083
rect 2387 2079 2388 2083
rect 2502 2080 2503 2084
rect 2507 2080 2508 2084
rect 2502 2079 2508 2080
rect 2382 2078 2388 2079
rect 1400 2055 1402 2078
rect 1568 2055 1570 2078
rect 1728 2055 1730 2078
rect 1872 2055 1874 2078
rect 2008 2055 2010 2078
rect 2136 2055 2138 2078
rect 2256 2055 2258 2078
rect 2384 2055 2386 2078
rect 2504 2055 2506 2079
rect 1327 2054 1331 2055
rect 1327 2049 1331 2050
rect 1399 2054 1403 2055
rect 1399 2049 1403 2050
rect 1447 2054 1451 2055
rect 1447 2049 1451 2050
rect 1551 2054 1555 2055
rect 1551 2049 1555 2050
rect 1567 2054 1571 2055
rect 1567 2049 1571 2050
rect 1655 2054 1659 2055
rect 1655 2049 1659 2050
rect 1727 2054 1731 2055
rect 1727 2049 1731 2050
rect 1751 2054 1755 2055
rect 1751 2049 1755 2050
rect 1839 2054 1843 2055
rect 1839 2049 1843 2050
rect 1871 2054 1875 2055
rect 1871 2049 1875 2050
rect 1927 2054 1931 2055
rect 1927 2049 1931 2050
rect 2007 2054 2011 2055
rect 2007 2049 2011 2050
rect 2023 2054 2027 2055
rect 2023 2049 2027 2050
rect 2119 2054 2123 2055
rect 2119 2049 2123 2050
rect 2135 2054 2139 2055
rect 2135 2049 2139 2050
rect 2255 2054 2259 2055
rect 2255 2049 2259 2050
rect 2383 2054 2387 2055
rect 2383 2049 2387 2050
rect 2503 2054 2507 2055
rect 2503 2049 2507 2050
rect 1238 2045 1239 2049
rect 1243 2045 1244 2049
rect 1238 2044 1244 2045
rect 1286 2048 1292 2049
rect 1286 2044 1287 2048
rect 1291 2044 1292 2048
rect 110 2043 116 2044
rect 1286 2043 1292 2044
rect 110 2031 116 2032
rect 110 2027 111 2031
rect 115 2027 116 2031
rect 1286 2031 1292 2032
rect 110 2026 116 2027
rect 382 2028 388 2029
rect 112 2019 114 2026
rect 382 2024 383 2028
rect 387 2024 388 2028
rect 382 2023 388 2024
rect 438 2028 444 2029
rect 438 2024 439 2028
rect 443 2024 444 2028
rect 438 2023 444 2024
rect 494 2028 500 2029
rect 494 2024 495 2028
rect 499 2024 500 2028
rect 494 2023 500 2024
rect 558 2028 564 2029
rect 558 2024 559 2028
rect 563 2024 564 2028
rect 558 2023 564 2024
rect 622 2028 628 2029
rect 622 2024 623 2028
rect 627 2024 628 2028
rect 622 2023 628 2024
rect 694 2028 700 2029
rect 694 2024 695 2028
rect 699 2024 700 2028
rect 694 2023 700 2024
rect 774 2028 780 2029
rect 774 2024 775 2028
rect 779 2024 780 2028
rect 774 2023 780 2024
rect 846 2028 852 2029
rect 846 2024 847 2028
rect 851 2024 852 2028
rect 846 2023 852 2024
rect 926 2028 932 2029
rect 926 2024 927 2028
rect 931 2024 932 2028
rect 926 2023 932 2024
rect 1006 2028 1012 2029
rect 1006 2024 1007 2028
rect 1011 2024 1012 2028
rect 1006 2023 1012 2024
rect 1086 2028 1092 2029
rect 1086 2024 1087 2028
rect 1091 2024 1092 2028
rect 1086 2023 1092 2024
rect 1166 2028 1172 2029
rect 1166 2024 1167 2028
rect 1171 2024 1172 2028
rect 1166 2023 1172 2024
rect 1222 2028 1228 2029
rect 1222 2024 1223 2028
rect 1227 2024 1228 2028
rect 1286 2027 1287 2031
rect 1291 2027 1292 2031
rect 1328 2029 1330 2049
rect 1448 2030 1450 2049
rect 1552 2030 1554 2049
rect 1656 2030 1658 2049
rect 1752 2030 1754 2049
rect 1840 2030 1842 2049
rect 1928 2030 1930 2049
rect 2024 2030 2026 2049
rect 2120 2030 2122 2049
rect 1446 2029 1452 2030
rect 1286 2026 1292 2027
rect 1326 2028 1332 2029
rect 1222 2023 1228 2024
rect 384 2019 386 2023
rect 440 2019 442 2023
rect 496 2019 498 2023
rect 560 2019 562 2023
rect 624 2019 626 2023
rect 696 2019 698 2023
rect 776 2019 778 2023
rect 848 2019 850 2023
rect 928 2019 930 2023
rect 1008 2019 1010 2023
rect 1088 2019 1090 2023
rect 1168 2019 1170 2023
rect 1224 2019 1226 2023
rect 1288 2019 1290 2026
rect 1326 2024 1327 2028
rect 1331 2024 1332 2028
rect 1446 2025 1447 2029
rect 1451 2025 1452 2029
rect 1446 2024 1452 2025
rect 1550 2029 1556 2030
rect 1550 2025 1551 2029
rect 1555 2025 1556 2029
rect 1550 2024 1556 2025
rect 1654 2029 1660 2030
rect 1654 2025 1655 2029
rect 1659 2025 1660 2029
rect 1654 2024 1660 2025
rect 1750 2029 1756 2030
rect 1750 2025 1751 2029
rect 1755 2025 1756 2029
rect 1750 2024 1756 2025
rect 1838 2029 1844 2030
rect 1838 2025 1839 2029
rect 1843 2025 1844 2029
rect 1838 2024 1844 2025
rect 1926 2029 1932 2030
rect 1926 2025 1927 2029
rect 1931 2025 1932 2029
rect 1926 2024 1932 2025
rect 2022 2029 2028 2030
rect 2022 2025 2023 2029
rect 2027 2025 2028 2029
rect 2022 2024 2028 2025
rect 2118 2029 2124 2030
rect 2504 2029 2506 2049
rect 2118 2025 2119 2029
rect 2123 2025 2124 2029
rect 2118 2024 2124 2025
rect 2502 2028 2508 2029
rect 2502 2024 2503 2028
rect 2507 2024 2508 2028
rect 1326 2023 1332 2024
rect 2502 2023 2508 2024
rect 111 2018 115 2019
rect 111 2013 115 2014
rect 231 2018 235 2019
rect 231 2013 235 2014
rect 287 2018 291 2019
rect 287 2013 291 2014
rect 359 2018 363 2019
rect 359 2013 363 2014
rect 383 2018 387 2019
rect 383 2013 387 2014
rect 439 2018 443 2019
rect 439 2013 443 2014
rect 495 2018 499 2019
rect 495 2013 499 2014
rect 535 2018 539 2019
rect 535 2013 539 2014
rect 559 2018 563 2019
rect 559 2013 563 2014
rect 623 2018 627 2019
rect 623 2013 627 2014
rect 631 2018 635 2019
rect 631 2013 635 2014
rect 695 2018 699 2019
rect 695 2013 699 2014
rect 735 2018 739 2019
rect 735 2013 739 2014
rect 775 2018 779 2019
rect 775 2013 779 2014
rect 847 2018 851 2019
rect 847 2013 851 2014
rect 927 2018 931 2019
rect 927 2013 931 2014
rect 959 2018 963 2019
rect 959 2013 963 2014
rect 1007 2018 1011 2019
rect 1007 2013 1011 2014
rect 1079 2018 1083 2019
rect 1079 2013 1083 2014
rect 1087 2018 1091 2019
rect 1087 2013 1091 2014
rect 1167 2018 1171 2019
rect 1167 2013 1171 2014
rect 1199 2018 1203 2019
rect 1199 2013 1203 2014
rect 1223 2018 1227 2019
rect 1223 2013 1227 2014
rect 1287 2018 1291 2019
rect 1287 2013 1291 2014
rect 112 2010 114 2013
rect 230 2012 236 2013
rect 110 2009 116 2010
rect 110 2005 111 2009
rect 115 2005 116 2009
rect 230 2008 231 2012
rect 235 2008 236 2012
rect 230 2007 236 2008
rect 286 2012 292 2013
rect 286 2008 287 2012
rect 291 2008 292 2012
rect 286 2007 292 2008
rect 358 2012 364 2013
rect 358 2008 359 2012
rect 363 2008 364 2012
rect 358 2007 364 2008
rect 438 2012 444 2013
rect 438 2008 439 2012
rect 443 2008 444 2012
rect 438 2007 444 2008
rect 534 2012 540 2013
rect 534 2008 535 2012
rect 539 2008 540 2012
rect 534 2007 540 2008
rect 630 2012 636 2013
rect 630 2008 631 2012
rect 635 2008 636 2012
rect 630 2007 636 2008
rect 734 2012 740 2013
rect 734 2008 735 2012
rect 739 2008 740 2012
rect 734 2007 740 2008
rect 846 2012 852 2013
rect 846 2008 847 2012
rect 851 2008 852 2012
rect 846 2007 852 2008
rect 958 2012 964 2013
rect 958 2008 959 2012
rect 963 2008 964 2012
rect 958 2007 964 2008
rect 1078 2012 1084 2013
rect 1078 2008 1079 2012
rect 1083 2008 1084 2012
rect 1078 2007 1084 2008
rect 1198 2012 1204 2013
rect 1198 2008 1199 2012
rect 1203 2008 1204 2012
rect 1288 2010 1290 2013
rect 1326 2011 1332 2012
rect 1198 2007 1204 2008
rect 1286 2009 1292 2010
rect 110 2004 116 2005
rect 1286 2005 1287 2009
rect 1291 2005 1292 2009
rect 1326 2007 1327 2011
rect 1331 2007 1332 2011
rect 2502 2011 2508 2012
rect 1326 2006 1332 2007
rect 1430 2008 1436 2009
rect 1286 2004 1292 2005
rect 1328 1999 1330 2006
rect 1430 2004 1431 2008
rect 1435 2004 1436 2008
rect 1430 2003 1436 2004
rect 1534 2008 1540 2009
rect 1534 2004 1535 2008
rect 1539 2004 1540 2008
rect 1534 2003 1540 2004
rect 1638 2008 1644 2009
rect 1638 2004 1639 2008
rect 1643 2004 1644 2008
rect 1638 2003 1644 2004
rect 1734 2008 1740 2009
rect 1734 2004 1735 2008
rect 1739 2004 1740 2008
rect 1734 2003 1740 2004
rect 1822 2008 1828 2009
rect 1822 2004 1823 2008
rect 1827 2004 1828 2008
rect 1822 2003 1828 2004
rect 1910 2008 1916 2009
rect 1910 2004 1911 2008
rect 1915 2004 1916 2008
rect 1910 2003 1916 2004
rect 2006 2008 2012 2009
rect 2006 2004 2007 2008
rect 2011 2004 2012 2008
rect 2006 2003 2012 2004
rect 2102 2008 2108 2009
rect 2102 2004 2103 2008
rect 2107 2004 2108 2008
rect 2502 2007 2503 2011
rect 2507 2007 2508 2011
rect 2502 2006 2508 2007
rect 2102 2003 2108 2004
rect 1432 1999 1434 2003
rect 1536 1999 1538 2003
rect 1640 1999 1642 2003
rect 1736 1999 1738 2003
rect 1824 1999 1826 2003
rect 1912 1999 1914 2003
rect 2008 1999 2010 2003
rect 2104 1999 2106 2003
rect 2504 1999 2506 2006
rect 1327 1998 1331 1999
rect 1327 1993 1331 1994
rect 1431 1998 1435 1999
rect 1431 1993 1435 1994
rect 1455 1998 1459 1999
rect 1455 1993 1459 1994
rect 1511 1998 1515 1999
rect 1511 1993 1515 1994
rect 1535 1998 1539 1999
rect 1535 1993 1539 1994
rect 1575 1998 1579 1999
rect 1575 1993 1579 1994
rect 1639 1998 1643 1999
rect 1639 1993 1643 1994
rect 1703 1998 1707 1999
rect 1703 1993 1707 1994
rect 1735 1998 1739 1999
rect 1735 1993 1739 1994
rect 1767 1998 1771 1999
rect 1767 1993 1771 1994
rect 1823 1998 1827 1999
rect 1823 1993 1827 1994
rect 1831 1998 1835 1999
rect 1831 1993 1835 1994
rect 1895 1998 1899 1999
rect 1895 1993 1899 1994
rect 1911 1998 1915 1999
rect 1911 1993 1915 1994
rect 1959 1998 1963 1999
rect 1959 1993 1963 1994
rect 2007 1998 2011 1999
rect 2007 1993 2011 1994
rect 2031 1998 2035 1999
rect 2031 1993 2035 1994
rect 2103 1998 2107 1999
rect 2103 1993 2107 1994
rect 2503 1998 2507 1999
rect 2503 1993 2507 1994
rect 110 1992 116 1993
rect 1286 1992 1292 1993
rect 110 1988 111 1992
rect 115 1988 116 1992
rect 110 1987 116 1988
rect 246 1991 252 1992
rect 246 1987 247 1991
rect 251 1987 252 1991
rect 112 1963 114 1987
rect 246 1986 252 1987
rect 302 1991 308 1992
rect 302 1987 303 1991
rect 307 1987 308 1991
rect 302 1986 308 1987
rect 374 1991 380 1992
rect 374 1987 375 1991
rect 379 1987 380 1991
rect 374 1986 380 1987
rect 454 1991 460 1992
rect 454 1987 455 1991
rect 459 1987 460 1991
rect 454 1986 460 1987
rect 550 1991 556 1992
rect 550 1987 551 1991
rect 555 1987 556 1991
rect 550 1986 556 1987
rect 646 1991 652 1992
rect 646 1987 647 1991
rect 651 1987 652 1991
rect 646 1986 652 1987
rect 750 1991 756 1992
rect 750 1987 751 1991
rect 755 1987 756 1991
rect 750 1986 756 1987
rect 862 1991 868 1992
rect 862 1987 863 1991
rect 867 1987 868 1991
rect 862 1986 868 1987
rect 974 1991 980 1992
rect 974 1987 975 1991
rect 979 1987 980 1991
rect 974 1986 980 1987
rect 1094 1991 1100 1992
rect 1094 1987 1095 1991
rect 1099 1987 1100 1991
rect 1094 1986 1100 1987
rect 1214 1991 1220 1992
rect 1214 1987 1215 1991
rect 1219 1987 1220 1991
rect 1286 1988 1287 1992
rect 1291 1988 1292 1992
rect 1328 1990 1330 1993
rect 1454 1992 1460 1993
rect 1286 1987 1292 1988
rect 1326 1989 1332 1990
rect 1214 1986 1220 1987
rect 248 1963 250 1986
rect 304 1963 306 1986
rect 376 1963 378 1986
rect 456 1963 458 1986
rect 552 1963 554 1986
rect 648 1963 650 1986
rect 752 1963 754 1986
rect 864 1963 866 1986
rect 976 1963 978 1986
rect 1096 1963 1098 1986
rect 1216 1963 1218 1986
rect 1288 1963 1290 1987
rect 1326 1985 1327 1989
rect 1331 1985 1332 1989
rect 1454 1988 1455 1992
rect 1459 1988 1460 1992
rect 1454 1987 1460 1988
rect 1510 1992 1516 1993
rect 1510 1988 1511 1992
rect 1515 1988 1516 1992
rect 1510 1987 1516 1988
rect 1574 1992 1580 1993
rect 1574 1988 1575 1992
rect 1579 1988 1580 1992
rect 1574 1987 1580 1988
rect 1638 1992 1644 1993
rect 1638 1988 1639 1992
rect 1643 1988 1644 1992
rect 1638 1987 1644 1988
rect 1702 1992 1708 1993
rect 1702 1988 1703 1992
rect 1707 1988 1708 1992
rect 1702 1987 1708 1988
rect 1766 1992 1772 1993
rect 1766 1988 1767 1992
rect 1771 1988 1772 1992
rect 1766 1987 1772 1988
rect 1830 1992 1836 1993
rect 1830 1988 1831 1992
rect 1835 1988 1836 1992
rect 1830 1987 1836 1988
rect 1894 1992 1900 1993
rect 1894 1988 1895 1992
rect 1899 1988 1900 1992
rect 1894 1987 1900 1988
rect 1958 1992 1964 1993
rect 1958 1988 1959 1992
rect 1963 1988 1964 1992
rect 1958 1987 1964 1988
rect 2030 1992 2036 1993
rect 2030 1988 2031 1992
rect 2035 1988 2036 1992
rect 2504 1990 2506 1993
rect 2030 1987 2036 1988
rect 2502 1989 2508 1990
rect 1326 1984 1332 1985
rect 2502 1985 2503 1989
rect 2507 1985 2508 1989
rect 2502 1984 2508 1985
rect 1326 1972 1332 1973
rect 2502 1972 2508 1973
rect 1326 1968 1327 1972
rect 1331 1968 1332 1972
rect 1326 1967 1332 1968
rect 1470 1971 1476 1972
rect 1470 1967 1471 1971
rect 1475 1967 1476 1971
rect 111 1962 115 1963
rect 111 1957 115 1958
rect 151 1962 155 1963
rect 151 1957 155 1958
rect 215 1962 219 1963
rect 215 1957 219 1958
rect 247 1962 251 1963
rect 247 1957 251 1958
rect 303 1962 307 1963
rect 303 1957 307 1958
rect 319 1962 323 1963
rect 319 1957 323 1958
rect 375 1962 379 1963
rect 375 1957 379 1958
rect 439 1962 443 1963
rect 439 1957 443 1958
rect 455 1962 459 1963
rect 455 1957 459 1958
rect 551 1962 555 1963
rect 551 1957 555 1958
rect 583 1962 587 1963
rect 583 1957 587 1958
rect 647 1962 651 1963
rect 647 1957 651 1958
rect 743 1962 747 1963
rect 743 1957 747 1958
rect 751 1962 755 1963
rect 751 1957 755 1958
rect 863 1962 867 1963
rect 863 1957 867 1958
rect 919 1962 923 1963
rect 919 1957 923 1958
rect 975 1962 979 1963
rect 975 1957 979 1958
rect 1095 1962 1099 1963
rect 1095 1957 1099 1958
rect 1215 1962 1219 1963
rect 1215 1957 1219 1958
rect 1287 1962 1291 1963
rect 1287 1957 1291 1958
rect 112 1937 114 1957
rect 152 1938 154 1957
rect 216 1938 218 1957
rect 320 1938 322 1957
rect 440 1938 442 1957
rect 584 1938 586 1957
rect 744 1938 746 1957
rect 920 1938 922 1957
rect 1096 1938 1098 1957
rect 150 1937 156 1938
rect 110 1936 116 1937
rect 110 1932 111 1936
rect 115 1932 116 1936
rect 150 1933 151 1937
rect 155 1933 156 1937
rect 150 1932 156 1933
rect 214 1937 220 1938
rect 214 1933 215 1937
rect 219 1933 220 1937
rect 214 1932 220 1933
rect 318 1937 324 1938
rect 318 1933 319 1937
rect 323 1933 324 1937
rect 318 1932 324 1933
rect 438 1937 444 1938
rect 438 1933 439 1937
rect 443 1933 444 1937
rect 438 1932 444 1933
rect 582 1937 588 1938
rect 582 1933 583 1937
rect 587 1933 588 1937
rect 582 1932 588 1933
rect 742 1937 748 1938
rect 742 1933 743 1937
rect 747 1933 748 1937
rect 742 1932 748 1933
rect 918 1937 924 1938
rect 918 1933 919 1937
rect 923 1933 924 1937
rect 918 1932 924 1933
rect 1094 1937 1100 1938
rect 1288 1937 1290 1957
rect 1328 1943 1330 1967
rect 1470 1966 1476 1967
rect 1526 1971 1532 1972
rect 1526 1967 1527 1971
rect 1531 1967 1532 1971
rect 1526 1966 1532 1967
rect 1590 1971 1596 1972
rect 1590 1967 1591 1971
rect 1595 1967 1596 1971
rect 1590 1966 1596 1967
rect 1654 1971 1660 1972
rect 1654 1967 1655 1971
rect 1659 1967 1660 1971
rect 1654 1966 1660 1967
rect 1718 1971 1724 1972
rect 1718 1967 1719 1971
rect 1723 1967 1724 1971
rect 1718 1966 1724 1967
rect 1782 1971 1788 1972
rect 1782 1967 1783 1971
rect 1787 1967 1788 1971
rect 1782 1966 1788 1967
rect 1846 1971 1852 1972
rect 1846 1967 1847 1971
rect 1851 1967 1852 1971
rect 1846 1966 1852 1967
rect 1910 1971 1916 1972
rect 1910 1967 1911 1971
rect 1915 1967 1916 1971
rect 1910 1966 1916 1967
rect 1974 1971 1980 1972
rect 1974 1967 1975 1971
rect 1979 1967 1980 1971
rect 1974 1966 1980 1967
rect 2046 1971 2052 1972
rect 2046 1967 2047 1971
rect 2051 1967 2052 1971
rect 2502 1968 2503 1972
rect 2507 1968 2508 1972
rect 2502 1967 2508 1968
rect 2046 1966 2052 1967
rect 1472 1943 1474 1966
rect 1528 1943 1530 1966
rect 1592 1943 1594 1966
rect 1656 1943 1658 1966
rect 1720 1943 1722 1966
rect 1784 1943 1786 1966
rect 1848 1943 1850 1966
rect 1912 1943 1914 1966
rect 1976 1943 1978 1966
rect 2048 1943 2050 1966
rect 2504 1943 2506 1967
rect 1327 1942 1331 1943
rect 1327 1937 1331 1938
rect 1471 1942 1475 1943
rect 1471 1937 1475 1938
rect 1527 1942 1531 1943
rect 1527 1937 1531 1938
rect 1567 1942 1571 1943
rect 1567 1937 1571 1938
rect 1591 1942 1595 1943
rect 1591 1937 1595 1938
rect 1631 1942 1635 1943
rect 1631 1937 1635 1938
rect 1655 1942 1659 1943
rect 1655 1937 1659 1938
rect 1703 1942 1707 1943
rect 1703 1937 1707 1938
rect 1719 1942 1723 1943
rect 1719 1937 1723 1938
rect 1775 1942 1779 1943
rect 1775 1937 1779 1938
rect 1783 1942 1787 1943
rect 1783 1937 1787 1938
rect 1847 1942 1851 1943
rect 1847 1937 1851 1938
rect 1911 1942 1915 1943
rect 1911 1937 1915 1938
rect 1919 1942 1923 1943
rect 1919 1937 1923 1938
rect 1975 1942 1979 1943
rect 1975 1937 1979 1938
rect 1999 1942 2003 1943
rect 1999 1937 2003 1938
rect 2047 1942 2051 1943
rect 2047 1937 2051 1938
rect 2087 1942 2091 1943
rect 2087 1937 2091 1938
rect 2183 1942 2187 1943
rect 2183 1937 2187 1938
rect 2279 1942 2283 1943
rect 2279 1937 2283 1938
rect 2375 1942 2379 1943
rect 2375 1937 2379 1938
rect 2455 1942 2459 1943
rect 2455 1937 2459 1938
rect 2503 1942 2507 1943
rect 2503 1937 2507 1938
rect 1094 1933 1095 1937
rect 1099 1933 1100 1937
rect 1094 1932 1100 1933
rect 1286 1936 1292 1937
rect 1286 1932 1287 1936
rect 1291 1932 1292 1936
rect 110 1931 116 1932
rect 1286 1931 1292 1932
rect 110 1919 116 1920
rect 110 1915 111 1919
rect 115 1915 116 1919
rect 1286 1919 1292 1920
rect 110 1914 116 1915
rect 134 1916 140 1917
rect 112 1903 114 1914
rect 134 1912 135 1916
rect 139 1912 140 1916
rect 134 1911 140 1912
rect 198 1916 204 1917
rect 198 1912 199 1916
rect 203 1912 204 1916
rect 198 1911 204 1912
rect 302 1916 308 1917
rect 302 1912 303 1916
rect 307 1912 308 1916
rect 302 1911 308 1912
rect 422 1916 428 1917
rect 422 1912 423 1916
rect 427 1912 428 1916
rect 422 1911 428 1912
rect 566 1916 572 1917
rect 566 1912 567 1916
rect 571 1912 572 1916
rect 566 1911 572 1912
rect 726 1916 732 1917
rect 726 1912 727 1916
rect 731 1912 732 1916
rect 726 1911 732 1912
rect 902 1916 908 1917
rect 902 1912 903 1916
rect 907 1912 908 1916
rect 902 1911 908 1912
rect 1078 1916 1084 1917
rect 1078 1912 1079 1916
rect 1083 1912 1084 1916
rect 1286 1915 1287 1919
rect 1291 1915 1292 1919
rect 1328 1917 1330 1937
rect 1568 1918 1570 1937
rect 1632 1918 1634 1937
rect 1704 1918 1706 1937
rect 1776 1918 1778 1937
rect 1848 1918 1850 1937
rect 1920 1918 1922 1937
rect 2000 1918 2002 1937
rect 2088 1918 2090 1937
rect 2184 1918 2186 1937
rect 2280 1918 2282 1937
rect 2376 1918 2378 1937
rect 2456 1918 2458 1937
rect 1566 1917 1572 1918
rect 1286 1914 1292 1915
rect 1326 1916 1332 1917
rect 1078 1911 1084 1912
rect 136 1903 138 1911
rect 200 1903 202 1911
rect 304 1903 306 1911
rect 424 1903 426 1911
rect 568 1903 570 1911
rect 728 1903 730 1911
rect 904 1903 906 1911
rect 1080 1903 1082 1911
rect 1288 1903 1290 1914
rect 1326 1912 1327 1916
rect 1331 1912 1332 1916
rect 1566 1913 1567 1917
rect 1571 1913 1572 1917
rect 1566 1912 1572 1913
rect 1630 1917 1636 1918
rect 1630 1913 1631 1917
rect 1635 1913 1636 1917
rect 1630 1912 1636 1913
rect 1702 1917 1708 1918
rect 1702 1913 1703 1917
rect 1707 1913 1708 1917
rect 1702 1912 1708 1913
rect 1774 1917 1780 1918
rect 1774 1913 1775 1917
rect 1779 1913 1780 1917
rect 1774 1912 1780 1913
rect 1846 1917 1852 1918
rect 1846 1913 1847 1917
rect 1851 1913 1852 1917
rect 1846 1912 1852 1913
rect 1918 1917 1924 1918
rect 1918 1913 1919 1917
rect 1923 1913 1924 1917
rect 1918 1912 1924 1913
rect 1998 1917 2004 1918
rect 1998 1913 1999 1917
rect 2003 1913 2004 1917
rect 1998 1912 2004 1913
rect 2086 1917 2092 1918
rect 2086 1913 2087 1917
rect 2091 1913 2092 1917
rect 2086 1912 2092 1913
rect 2182 1917 2188 1918
rect 2182 1913 2183 1917
rect 2187 1913 2188 1917
rect 2182 1912 2188 1913
rect 2278 1917 2284 1918
rect 2278 1913 2279 1917
rect 2283 1913 2284 1917
rect 2278 1912 2284 1913
rect 2374 1917 2380 1918
rect 2374 1913 2375 1917
rect 2379 1913 2380 1917
rect 2374 1912 2380 1913
rect 2454 1917 2460 1918
rect 2504 1917 2506 1937
rect 2454 1913 2455 1917
rect 2459 1913 2460 1917
rect 2454 1912 2460 1913
rect 2502 1916 2508 1917
rect 2502 1912 2503 1916
rect 2507 1912 2508 1916
rect 1326 1911 1332 1912
rect 2502 1911 2508 1912
rect 111 1902 115 1903
rect 111 1897 115 1898
rect 135 1902 139 1903
rect 135 1897 139 1898
rect 191 1902 195 1903
rect 191 1897 195 1898
rect 199 1902 203 1903
rect 199 1897 203 1898
rect 271 1902 275 1903
rect 271 1897 275 1898
rect 303 1902 307 1903
rect 303 1897 307 1898
rect 359 1902 363 1903
rect 359 1897 363 1898
rect 423 1902 427 1903
rect 423 1897 427 1898
rect 455 1902 459 1903
rect 455 1897 459 1898
rect 543 1902 547 1903
rect 543 1897 547 1898
rect 567 1902 571 1903
rect 567 1897 571 1898
rect 631 1902 635 1903
rect 631 1897 635 1898
rect 719 1902 723 1903
rect 719 1897 723 1898
rect 727 1902 731 1903
rect 727 1897 731 1898
rect 799 1902 803 1903
rect 799 1897 803 1898
rect 871 1902 875 1903
rect 871 1897 875 1898
rect 903 1902 907 1903
rect 903 1897 907 1898
rect 943 1902 947 1903
rect 943 1897 947 1898
rect 1015 1902 1019 1903
rect 1015 1897 1019 1898
rect 1079 1902 1083 1903
rect 1079 1897 1083 1898
rect 1087 1902 1091 1903
rect 1087 1897 1091 1898
rect 1159 1902 1163 1903
rect 1159 1897 1163 1898
rect 1287 1902 1291 1903
rect 1287 1897 1291 1898
rect 1326 1899 1332 1900
rect 112 1894 114 1897
rect 134 1896 140 1897
rect 110 1893 116 1894
rect 110 1889 111 1893
rect 115 1889 116 1893
rect 134 1892 135 1896
rect 139 1892 140 1896
rect 134 1891 140 1892
rect 190 1896 196 1897
rect 190 1892 191 1896
rect 195 1892 196 1896
rect 190 1891 196 1892
rect 270 1896 276 1897
rect 270 1892 271 1896
rect 275 1892 276 1896
rect 270 1891 276 1892
rect 358 1896 364 1897
rect 358 1892 359 1896
rect 363 1892 364 1896
rect 358 1891 364 1892
rect 454 1896 460 1897
rect 454 1892 455 1896
rect 459 1892 460 1896
rect 454 1891 460 1892
rect 542 1896 548 1897
rect 542 1892 543 1896
rect 547 1892 548 1896
rect 542 1891 548 1892
rect 630 1896 636 1897
rect 630 1892 631 1896
rect 635 1892 636 1896
rect 630 1891 636 1892
rect 718 1896 724 1897
rect 718 1892 719 1896
rect 723 1892 724 1896
rect 718 1891 724 1892
rect 798 1896 804 1897
rect 798 1892 799 1896
rect 803 1892 804 1896
rect 798 1891 804 1892
rect 870 1896 876 1897
rect 870 1892 871 1896
rect 875 1892 876 1896
rect 870 1891 876 1892
rect 942 1896 948 1897
rect 942 1892 943 1896
rect 947 1892 948 1896
rect 942 1891 948 1892
rect 1014 1896 1020 1897
rect 1014 1892 1015 1896
rect 1019 1892 1020 1896
rect 1014 1891 1020 1892
rect 1086 1896 1092 1897
rect 1086 1892 1087 1896
rect 1091 1892 1092 1896
rect 1086 1891 1092 1892
rect 1158 1896 1164 1897
rect 1158 1892 1159 1896
rect 1163 1892 1164 1896
rect 1288 1894 1290 1897
rect 1326 1895 1327 1899
rect 1331 1895 1332 1899
rect 2502 1899 2508 1900
rect 1326 1894 1332 1895
rect 1550 1896 1556 1897
rect 1158 1891 1164 1892
rect 1286 1893 1292 1894
rect 110 1888 116 1889
rect 1286 1889 1287 1893
rect 1291 1889 1292 1893
rect 1286 1888 1292 1889
rect 1328 1887 1330 1894
rect 1550 1892 1551 1896
rect 1555 1892 1556 1896
rect 1550 1891 1556 1892
rect 1614 1896 1620 1897
rect 1614 1892 1615 1896
rect 1619 1892 1620 1896
rect 1614 1891 1620 1892
rect 1686 1896 1692 1897
rect 1686 1892 1687 1896
rect 1691 1892 1692 1896
rect 1686 1891 1692 1892
rect 1758 1896 1764 1897
rect 1758 1892 1759 1896
rect 1763 1892 1764 1896
rect 1758 1891 1764 1892
rect 1830 1896 1836 1897
rect 1830 1892 1831 1896
rect 1835 1892 1836 1896
rect 1830 1891 1836 1892
rect 1902 1896 1908 1897
rect 1902 1892 1903 1896
rect 1907 1892 1908 1896
rect 1902 1891 1908 1892
rect 1982 1896 1988 1897
rect 1982 1892 1983 1896
rect 1987 1892 1988 1896
rect 1982 1891 1988 1892
rect 2070 1896 2076 1897
rect 2070 1892 2071 1896
rect 2075 1892 2076 1896
rect 2070 1891 2076 1892
rect 2166 1896 2172 1897
rect 2166 1892 2167 1896
rect 2171 1892 2172 1896
rect 2166 1891 2172 1892
rect 2262 1896 2268 1897
rect 2262 1892 2263 1896
rect 2267 1892 2268 1896
rect 2262 1891 2268 1892
rect 2358 1896 2364 1897
rect 2358 1892 2359 1896
rect 2363 1892 2364 1896
rect 2358 1891 2364 1892
rect 2438 1896 2444 1897
rect 2438 1892 2439 1896
rect 2443 1892 2444 1896
rect 2502 1895 2503 1899
rect 2507 1895 2508 1899
rect 2502 1894 2508 1895
rect 2438 1891 2444 1892
rect 1552 1887 1554 1891
rect 1616 1887 1618 1891
rect 1688 1887 1690 1891
rect 1760 1887 1762 1891
rect 1832 1887 1834 1891
rect 1904 1887 1906 1891
rect 1984 1887 1986 1891
rect 2072 1887 2074 1891
rect 2168 1887 2170 1891
rect 2264 1887 2266 1891
rect 2360 1887 2362 1891
rect 2440 1887 2442 1891
rect 2504 1887 2506 1894
rect 1327 1886 1331 1887
rect 1327 1881 1331 1882
rect 1551 1886 1555 1887
rect 1551 1881 1555 1882
rect 1607 1886 1611 1887
rect 1607 1881 1611 1882
rect 1615 1886 1619 1887
rect 1615 1881 1619 1882
rect 1663 1886 1667 1887
rect 1663 1881 1667 1882
rect 1687 1886 1691 1887
rect 1687 1881 1691 1882
rect 1727 1886 1731 1887
rect 1727 1881 1731 1882
rect 1759 1886 1763 1887
rect 1759 1881 1763 1882
rect 1799 1886 1803 1887
rect 1799 1881 1803 1882
rect 1831 1886 1835 1887
rect 1831 1881 1835 1882
rect 1871 1886 1875 1887
rect 1871 1881 1875 1882
rect 1903 1886 1907 1887
rect 1903 1881 1907 1882
rect 1943 1886 1947 1887
rect 1943 1881 1947 1882
rect 1983 1886 1987 1887
rect 1983 1881 1987 1882
rect 2007 1886 2011 1887
rect 2007 1881 2011 1882
rect 2071 1886 2075 1887
rect 2071 1881 2075 1882
rect 2135 1886 2139 1887
rect 2135 1881 2139 1882
rect 2167 1886 2171 1887
rect 2167 1881 2171 1882
rect 2199 1886 2203 1887
rect 2199 1881 2203 1882
rect 2263 1886 2267 1887
rect 2263 1881 2267 1882
rect 2327 1886 2331 1887
rect 2327 1881 2331 1882
rect 2359 1886 2363 1887
rect 2359 1881 2363 1882
rect 2383 1886 2387 1887
rect 2383 1881 2387 1882
rect 2439 1886 2443 1887
rect 2439 1881 2443 1882
rect 2503 1886 2507 1887
rect 2503 1881 2507 1882
rect 1328 1878 1330 1881
rect 1606 1880 1612 1881
rect 1326 1877 1332 1878
rect 110 1876 116 1877
rect 1286 1876 1292 1877
rect 110 1872 111 1876
rect 115 1872 116 1876
rect 110 1871 116 1872
rect 150 1875 156 1876
rect 150 1871 151 1875
rect 155 1871 156 1875
rect 112 1851 114 1871
rect 150 1870 156 1871
rect 206 1875 212 1876
rect 206 1871 207 1875
rect 211 1871 212 1875
rect 206 1870 212 1871
rect 286 1875 292 1876
rect 286 1871 287 1875
rect 291 1871 292 1875
rect 286 1870 292 1871
rect 374 1875 380 1876
rect 374 1871 375 1875
rect 379 1871 380 1875
rect 374 1870 380 1871
rect 470 1875 476 1876
rect 470 1871 471 1875
rect 475 1871 476 1875
rect 470 1870 476 1871
rect 558 1875 564 1876
rect 558 1871 559 1875
rect 563 1871 564 1875
rect 558 1870 564 1871
rect 646 1875 652 1876
rect 646 1871 647 1875
rect 651 1871 652 1875
rect 646 1870 652 1871
rect 734 1875 740 1876
rect 734 1871 735 1875
rect 739 1871 740 1875
rect 734 1870 740 1871
rect 814 1875 820 1876
rect 814 1871 815 1875
rect 819 1871 820 1875
rect 814 1870 820 1871
rect 886 1875 892 1876
rect 886 1871 887 1875
rect 891 1871 892 1875
rect 886 1870 892 1871
rect 958 1875 964 1876
rect 958 1871 959 1875
rect 963 1871 964 1875
rect 958 1870 964 1871
rect 1030 1875 1036 1876
rect 1030 1871 1031 1875
rect 1035 1871 1036 1875
rect 1030 1870 1036 1871
rect 1102 1875 1108 1876
rect 1102 1871 1103 1875
rect 1107 1871 1108 1875
rect 1102 1870 1108 1871
rect 1174 1875 1180 1876
rect 1174 1871 1175 1875
rect 1179 1871 1180 1875
rect 1286 1872 1287 1876
rect 1291 1872 1292 1876
rect 1326 1873 1327 1877
rect 1331 1873 1332 1877
rect 1606 1876 1607 1880
rect 1611 1876 1612 1880
rect 1606 1875 1612 1876
rect 1662 1880 1668 1881
rect 1662 1876 1663 1880
rect 1667 1876 1668 1880
rect 1662 1875 1668 1876
rect 1726 1880 1732 1881
rect 1726 1876 1727 1880
rect 1731 1876 1732 1880
rect 1726 1875 1732 1876
rect 1798 1880 1804 1881
rect 1798 1876 1799 1880
rect 1803 1876 1804 1880
rect 1798 1875 1804 1876
rect 1870 1880 1876 1881
rect 1870 1876 1871 1880
rect 1875 1876 1876 1880
rect 1870 1875 1876 1876
rect 1942 1880 1948 1881
rect 1942 1876 1943 1880
rect 1947 1876 1948 1880
rect 1942 1875 1948 1876
rect 2006 1880 2012 1881
rect 2006 1876 2007 1880
rect 2011 1876 2012 1880
rect 2006 1875 2012 1876
rect 2070 1880 2076 1881
rect 2070 1876 2071 1880
rect 2075 1876 2076 1880
rect 2070 1875 2076 1876
rect 2134 1880 2140 1881
rect 2134 1876 2135 1880
rect 2139 1876 2140 1880
rect 2134 1875 2140 1876
rect 2198 1880 2204 1881
rect 2198 1876 2199 1880
rect 2203 1876 2204 1880
rect 2198 1875 2204 1876
rect 2262 1880 2268 1881
rect 2262 1876 2263 1880
rect 2267 1876 2268 1880
rect 2262 1875 2268 1876
rect 2326 1880 2332 1881
rect 2326 1876 2327 1880
rect 2331 1876 2332 1880
rect 2326 1875 2332 1876
rect 2382 1880 2388 1881
rect 2382 1876 2383 1880
rect 2387 1876 2388 1880
rect 2382 1875 2388 1876
rect 2438 1880 2444 1881
rect 2438 1876 2439 1880
rect 2443 1876 2444 1880
rect 2504 1878 2506 1881
rect 2438 1875 2444 1876
rect 2502 1877 2508 1878
rect 1326 1872 1332 1873
rect 2502 1873 2503 1877
rect 2507 1873 2508 1877
rect 2502 1872 2508 1873
rect 1286 1871 1292 1872
rect 1174 1870 1180 1871
rect 152 1851 154 1870
rect 208 1851 210 1870
rect 288 1851 290 1870
rect 376 1851 378 1870
rect 472 1851 474 1870
rect 560 1851 562 1870
rect 648 1851 650 1870
rect 736 1851 738 1870
rect 816 1851 818 1870
rect 888 1851 890 1870
rect 960 1851 962 1870
rect 1032 1851 1034 1870
rect 1104 1851 1106 1870
rect 1176 1851 1178 1870
rect 1288 1851 1290 1871
rect 1326 1860 1332 1861
rect 2502 1860 2508 1861
rect 1326 1856 1327 1860
rect 1331 1856 1332 1860
rect 1326 1855 1332 1856
rect 1622 1859 1628 1860
rect 1622 1855 1623 1859
rect 1627 1855 1628 1859
rect 111 1850 115 1851
rect 111 1845 115 1846
rect 151 1850 155 1851
rect 151 1845 155 1846
rect 207 1850 211 1851
rect 207 1845 211 1846
rect 287 1850 291 1851
rect 287 1845 291 1846
rect 295 1850 299 1851
rect 295 1845 299 1846
rect 375 1850 379 1851
rect 375 1845 379 1846
rect 391 1850 395 1851
rect 391 1845 395 1846
rect 471 1850 475 1851
rect 471 1845 475 1846
rect 495 1850 499 1851
rect 495 1845 499 1846
rect 559 1850 563 1851
rect 559 1845 563 1846
rect 591 1850 595 1851
rect 591 1845 595 1846
rect 647 1850 651 1851
rect 647 1845 651 1846
rect 687 1850 691 1851
rect 687 1845 691 1846
rect 735 1850 739 1851
rect 735 1845 739 1846
rect 775 1850 779 1851
rect 775 1845 779 1846
rect 815 1850 819 1851
rect 815 1845 819 1846
rect 855 1850 859 1851
rect 855 1845 859 1846
rect 887 1850 891 1851
rect 887 1845 891 1846
rect 927 1850 931 1851
rect 927 1845 931 1846
rect 959 1850 963 1851
rect 959 1845 963 1846
rect 999 1850 1003 1851
rect 999 1845 1003 1846
rect 1031 1850 1035 1851
rect 1031 1845 1035 1846
rect 1079 1850 1083 1851
rect 1079 1845 1083 1846
rect 1103 1850 1107 1851
rect 1103 1845 1107 1846
rect 1159 1850 1163 1851
rect 1159 1845 1163 1846
rect 1175 1850 1179 1851
rect 1175 1845 1179 1846
rect 1287 1850 1291 1851
rect 1287 1845 1291 1846
rect 112 1825 114 1845
rect 152 1826 154 1845
rect 208 1826 210 1845
rect 296 1826 298 1845
rect 392 1826 394 1845
rect 496 1826 498 1845
rect 592 1826 594 1845
rect 688 1826 690 1845
rect 776 1826 778 1845
rect 856 1826 858 1845
rect 928 1826 930 1845
rect 1000 1826 1002 1845
rect 1080 1826 1082 1845
rect 1160 1826 1162 1845
rect 150 1825 156 1826
rect 110 1824 116 1825
rect 110 1820 111 1824
rect 115 1820 116 1824
rect 150 1821 151 1825
rect 155 1821 156 1825
rect 150 1820 156 1821
rect 206 1825 212 1826
rect 206 1821 207 1825
rect 211 1821 212 1825
rect 206 1820 212 1821
rect 294 1825 300 1826
rect 294 1821 295 1825
rect 299 1821 300 1825
rect 294 1820 300 1821
rect 390 1825 396 1826
rect 390 1821 391 1825
rect 395 1821 396 1825
rect 390 1820 396 1821
rect 494 1825 500 1826
rect 494 1821 495 1825
rect 499 1821 500 1825
rect 494 1820 500 1821
rect 590 1825 596 1826
rect 590 1821 591 1825
rect 595 1821 596 1825
rect 590 1820 596 1821
rect 686 1825 692 1826
rect 686 1821 687 1825
rect 691 1821 692 1825
rect 686 1820 692 1821
rect 774 1825 780 1826
rect 774 1821 775 1825
rect 779 1821 780 1825
rect 774 1820 780 1821
rect 854 1825 860 1826
rect 854 1821 855 1825
rect 859 1821 860 1825
rect 854 1820 860 1821
rect 926 1825 932 1826
rect 926 1821 927 1825
rect 931 1821 932 1825
rect 926 1820 932 1821
rect 998 1825 1004 1826
rect 998 1821 999 1825
rect 1003 1821 1004 1825
rect 998 1820 1004 1821
rect 1078 1825 1084 1826
rect 1078 1821 1079 1825
rect 1083 1821 1084 1825
rect 1078 1820 1084 1821
rect 1158 1825 1164 1826
rect 1288 1825 1290 1845
rect 1328 1831 1330 1855
rect 1622 1854 1628 1855
rect 1678 1859 1684 1860
rect 1678 1855 1679 1859
rect 1683 1855 1684 1859
rect 1678 1854 1684 1855
rect 1742 1859 1748 1860
rect 1742 1855 1743 1859
rect 1747 1855 1748 1859
rect 1742 1854 1748 1855
rect 1814 1859 1820 1860
rect 1814 1855 1815 1859
rect 1819 1855 1820 1859
rect 1814 1854 1820 1855
rect 1886 1859 1892 1860
rect 1886 1855 1887 1859
rect 1891 1855 1892 1859
rect 1886 1854 1892 1855
rect 1958 1859 1964 1860
rect 1958 1855 1959 1859
rect 1963 1855 1964 1859
rect 1958 1854 1964 1855
rect 2022 1859 2028 1860
rect 2022 1855 2023 1859
rect 2027 1855 2028 1859
rect 2022 1854 2028 1855
rect 2086 1859 2092 1860
rect 2086 1855 2087 1859
rect 2091 1855 2092 1859
rect 2086 1854 2092 1855
rect 2150 1859 2156 1860
rect 2150 1855 2151 1859
rect 2155 1855 2156 1859
rect 2150 1854 2156 1855
rect 2214 1859 2220 1860
rect 2214 1855 2215 1859
rect 2219 1855 2220 1859
rect 2214 1854 2220 1855
rect 2278 1859 2284 1860
rect 2278 1855 2279 1859
rect 2283 1855 2284 1859
rect 2278 1854 2284 1855
rect 2342 1859 2348 1860
rect 2342 1855 2343 1859
rect 2347 1855 2348 1859
rect 2342 1854 2348 1855
rect 2398 1859 2404 1860
rect 2398 1855 2399 1859
rect 2403 1855 2404 1859
rect 2398 1854 2404 1855
rect 2454 1859 2460 1860
rect 2454 1855 2455 1859
rect 2459 1855 2460 1859
rect 2502 1856 2503 1860
rect 2507 1856 2508 1860
rect 2502 1855 2508 1856
rect 2454 1854 2460 1855
rect 1624 1831 1626 1854
rect 1680 1831 1682 1854
rect 1744 1831 1746 1854
rect 1816 1831 1818 1854
rect 1888 1831 1890 1854
rect 1960 1831 1962 1854
rect 2024 1831 2026 1854
rect 2088 1831 2090 1854
rect 2152 1831 2154 1854
rect 2216 1831 2218 1854
rect 2280 1831 2282 1854
rect 2344 1831 2346 1854
rect 2400 1831 2402 1854
rect 2456 1831 2458 1854
rect 2504 1831 2506 1855
rect 1327 1830 1331 1831
rect 1327 1825 1331 1826
rect 1623 1830 1627 1831
rect 1623 1825 1627 1826
rect 1631 1830 1635 1831
rect 1631 1825 1635 1826
rect 1679 1830 1683 1831
rect 1679 1825 1683 1826
rect 1719 1830 1723 1831
rect 1719 1825 1723 1826
rect 1743 1830 1747 1831
rect 1743 1825 1747 1826
rect 1815 1830 1819 1831
rect 1815 1825 1819 1826
rect 1887 1830 1891 1831
rect 1887 1825 1891 1826
rect 1927 1830 1931 1831
rect 1927 1825 1931 1826
rect 1959 1830 1963 1831
rect 1959 1825 1963 1826
rect 2023 1830 2027 1831
rect 2023 1825 2027 1826
rect 2055 1830 2059 1831
rect 2055 1825 2059 1826
rect 2087 1830 2091 1831
rect 2087 1825 2091 1826
rect 2151 1830 2155 1831
rect 2151 1825 2155 1826
rect 2191 1830 2195 1831
rect 2191 1825 2195 1826
rect 2215 1830 2219 1831
rect 2215 1825 2219 1826
rect 2279 1830 2283 1831
rect 2279 1825 2283 1826
rect 2335 1830 2339 1831
rect 2335 1825 2339 1826
rect 2343 1830 2347 1831
rect 2343 1825 2347 1826
rect 2399 1830 2403 1831
rect 2399 1825 2403 1826
rect 2455 1830 2459 1831
rect 2455 1825 2459 1826
rect 2503 1830 2507 1831
rect 2503 1825 2507 1826
rect 1158 1821 1159 1825
rect 1163 1821 1164 1825
rect 1158 1820 1164 1821
rect 1286 1824 1292 1825
rect 1286 1820 1287 1824
rect 1291 1820 1292 1824
rect 110 1819 116 1820
rect 1286 1819 1292 1820
rect 110 1807 116 1808
rect 110 1803 111 1807
rect 115 1803 116 1807
rect 1286 1807 1292 1808
rect 110 1802 116 1803
rect 134 1804 140 1805
rect 112 1787 114 1802
rect 134 1800 135 1804
rect 139 1800 140 1804
rect 134 1799 140 1800
rect 190 1804 196 1805
rect 190 1800 191 1804
rect 195 1800 196 1804
rect 190 1799 196 1800
rect 278 1804 284 1805
rect 278 1800 279 1804
rect 283 1800 284 1804
rect 278 1799 284 1800
rect 374 1804 380 1805
rect 374 1800 375 1804
rect 379 1800 380 1804
rect 374 1799 380 1800
rect 478 1804 484 1805
rect 478 1800 479 1804
rect 483 1800 484 1804
rect 478 1799 484 1800
rect 574 1804 580 1805
rect 574 1800 575 1804
rect 579 1800 580 1804
rect 574 1799 580 1800
rect 670 1804 676 1805
rect 670 1800 671 1804
rect 675 1800 676 1804
rect 670 1799 676 1800
rect 758 1804 764 1805
rect 758 1800 759 1804
rect 763 1800 764 1804
rect 758 1799 764 1800
rect 838 1804 844 1805
rect 838 1800 839 1804
rect 843 1800 844 1804
rect 838 1799 844 1800
rect 910 1804 916 1805
rect 910 1800 911 1804
rect 915 1800 916 1804
rect 910 1799 916 1800
rect 982 1804 988 1805
rect 982 1800 983 1804
rect 987 1800 988 1804
rect 982 1799 988 1800
rect 1062 1804 1068 1805
rect 1062 1800 1063 1804
rect 1067 1800 1068 1804
rect 1062 1799 1068 1800
rect 1142 1804 1148 1805
rect 1142 1800 1143 1804
rect 1147 1800 1148 1804
rect 1286 1803 1287 1807
rect 1291 1803 1292 1807
rect 1328 1805 1330 1825
rect 1632 1806 1634 1825
rect 1720 1806 1722 1825
rect 1816 1806 1818 1825
rect 1928 1806 1930 1825
rect 2056 1806 2058 1825
rect 2192 1806 2194 1825
rect 2336 1806 2338 1825
rect 2456 1806 2458 1825
rect 1630 1805 1636 1806
rect 1286 1802 1292 1803
rect 1326 1804 1332 1805
rect 1142 1799 1148 1800
rect 136 1787 138 1799
rect 192 1787 194 1799
rect 280 1787 282 1799
rect 376 1787 378 1799
rect 480 1787 482 1799
rect 576 1787 578 1799
rect 672 1787 674 1799
rect 760 1787 762 1799
rect 840 1787 842 1799
rect 912 1787 914 1799
rect 984 1787 986 1799
rect 1064 1787 1066 1799
rect 1144 1787 1146 1799
rect 1288 1787 1290 1802
rect 1326 1800 1327 1804
rect 1331 1800 1332 1804
rect 1630 1801 1631 1805
rect 1635 1801 1636 1805
rect 1630 1800 1636 1801
rect 1718 1805 1724 1806
rect 1718 1801 1719 1805
rect 1723 1801 1724 1805
rect 1718 1800 1724 1801
rect 1814 1805 1820 1806
rect 1814 1801 1815 1805
rect 1819 1801 1820 1805
rect 1814 1800 1820 1801
rect 1926 1805 1932 1806
rect 1926 1801 1927 1805
rect 1931 1801 1932 1805
rect 1926 1800 1932 1801
rect 2054 1805 2060 1806
rect 2054 1801 2055 1805
rect 2059 1801 2060 1805
rect 2054 1800 2060 1801
rect 2190 1805 2196 1806
rect 2190 1801 2191 1805
rect 2195 1801 2196 1805
rect 2190 1800 2196 1801
rect 2334 1805 2340 1806
rect 2334 1801 2335 1805
rect 2339 1801 2340 1805
rect 2334 1800 2340 1801
rect 2454 1805 2460 1806
rect 2504 1805 2506 1825
rect 2454 1801 2455 1805
rect 2459 1801 2460 1805
rect 2454 1800 2460 1801
rect 2502 1804 2508 1805
rect 2502 1800 2503 1804
rect 2507 1800 2508 1804
rect 1326 1799 1332 1800
rect 2502 1799 2508 1800
rect 1326 1787 1332 1788
rect 111 1786 115 1787
rect 111 1781 115 1782
rect 135 1786 139 1787
rect 135 1781 139 1782
rect 191 1786 195 1787
rect 191 1781 195 1782
rect 199 1786 203 1787
rect 199 1781 203 1782
rect 279 1786 283 1787
rect 279 1781 283 1782
rect 295 1786 299 1787
rect 295 1781 299 1782
rect 375 1786 379 1787
rect 375 1781 379 1782
rect 399 1786 403 1787
rect 399 1781 403 1782
rect 479 1786 483 1787
rect 479 1781 483 1782
rect 503 1786 507 1787
rect 503 1781 507 1782
rect 575 1786 579 1787
rect 575 1781 579 1782
rect 607 1786 611 1787
rect 607 1781 611 1782
rect 671 1786 675 1787
rect 671 1781 675 1782
rect 703 1786 707 1787
rect 703 1781 707 1782
rect 759 1786 763 1787
rect 759 1781 763 1782
rect 799 1786 803 1787
rect 799 1781 803 1782
rect 839 1786 843 1787
rect 839 1781 843 1782
rect 887 1786 891 1787
rect 887 1781 891 1782
rect 911 1786 915 1787
rect 911 1781 915 1782
rect 975 1786 979 1787
rect 975 1781 979 1782
rect 983 1786 987 1787
rect 983 1781 987 1782
rect 1063 1786 1067 1787
rect 1063 1781 1067 1782
rect 1143 1786 1147 1787
rect 1143 1781 1147 1782
rect 1151 1786 1155 1787
rect 1151 1781 1155 1782
rect 1287 1786 1291 1787
rect 1326 1783 1327 1787
rect 1331 1783 1332 1787
rect 2502 1787 2508 1788
rect 1326 1782 1332 1783
rect 1614 1784 1620 1785
rect 1287 1781 1291 1782
rect 112 1778 114 1781
rect 134 1780 140 1781
rect 110 1777 116 1778
rect 110 1773 111 1777
rect 115 1773 116 1777
rect 134 1776 135 1780
rect 139 1776 140 1780
rect 134 1775 140 1776
rect 198 1780 204 1781
rect 198 1776 199 1780
rect 203 1776 204 1780
rect 198 1775 204 1776
rect 294 1780 300 1781
rect 294 1776 295 1780
rect 299 1776 300 1780
rect 294 1775 300 1776
rect 398 1780 404 1781
rect 398 1776 399 1780
rect 403 1776 404 1780
rect 398 1775 404 1776
rect 502 1780 508 1781
rect 502 1776 503 1780
rect 507 1776 508 1780
rect 502 1775 508 1776
rect 606 1780 612 1781
rect 606 1776 607 1780
rect 611 1776 612 1780
rect 606 1775 612 1776
rect 702 1780 708 1781
rect 702 1776 703 1780
rect 707 1776 708 1780
rect 702 1775 708 1776
rect 798 1780 804 1781
rect 798 1776 799 1780
rect 803 1776 804 1780
rect 798 1775 804 1776
rect 886 1780 892 1781
rect 886 1776 887 1780
rect 891 1776 892 1780
rect 886 1775 892 1776
rect 974 1780 980 1781
rect 974 1776 975 1780
rect 979 1776 980 1780
rect 974 1775 980 1776
rect 1062 1780 1068 1781
rect 1062 1776 1063 1780
rect 1067 1776 1068 1780
rect 1062 1775 1068 1776
rect 1150 1780 1156 1781
rect 1150 1776 1151 1780
rect 1155 1776 1156 1780
rect 1288 1778 1290 1781
rect 1328 1779 1330 1782
rect 1614 1780 1615 1784
rect 1619 1780 1620 1784
rect 1614 1779 1620 1780
rect 1702 1784 1708 1785
rect 1702 1780 1703 1784
rect 1707 1780 1708 1784
rect 1702 1779 1708 1780
rect 1798 1784 1804 1785
rect 1798 1780 1799 1784
rect 1803 1780 1804 1784
rect 1798 1779 1804 1780
rect 1910 1784 1916 1785
rect 1910 1780 1911 1784
rect 1915 1780 1916 1784
rect 1910 1779 1916 1780
rect 2038 1784 2044 1785
rect 2038 1780 2039 1784
rect 2043 1780 2044 1784
rect 2038 1779 2044 1780
rect 2174 1784 2180 1785
rect 2174 1780 2175 1784
rect 2179 1780 2180 1784
rect 2174 1779 2180 1780
rect 2318 1784 2324 1785
rect 2318 1780 2319 1784
rect 2323 1780 2324 1784
rect 2318 1779 2324 1780
rect 2438 1784 2444 1785
rect 2438 1780 2439 1784
rect 2443 1780 2444 1784
rect 2502 1783 2503 1787
rect 2507 1783 2508 1787
rect 2502 1782 2508 1783
rect 2438 1779 2444 1780
rect 2504 1779 2506 1782
rect 1327 1778 1331 1779
rect 1150 1775 1156 1776
rect 1286 1777 1292 1778
rect 110 1772 116 1773
rect 1286 1773 1287 1777
rect 1291 1773 1292 1777
rect 1327 1773 1331 1774
rect 1527 1778 1531 1779
rect 1527 1773 1531 1774
rect 1607 1778 1611 1779
rect 1607 1773 1611 1774
rect 1615 1778 1619 1779
rect 1615 1773 1619 1774
rect 1695 1778 1699 1779
rect 1695 1773 1699 1774
rect 1703 1778 1707 1779
rect 1703 1773 1707 1774
rect 1791 1778 1795 1779
rect 1791 1773 1795 1774
rect 1799 1778 1803 1779
rect 1799 1773 1803 1774
rect 1879 1778 1883 1779
rect 1879 1773 1883 1774
rect 1911 1778 1915 1779
rect 1911 1773 1915 1774
rect 1967 1778 1971 1779
rect 1967 1773 1971 1774
rect 2039 1778 2043 1779
rect 2039 1773 2043 1774
rect 2055 1778 2059 1779
rect 2055 1773 2059 1774
rect 2135 1778 2139 1779
rect 2135 1773 2139 1774
rect 2175 1778 2179 1779
rect 2175 1773 2179 1774
rect 2215 1778 2219 1779
rect 2215 1773 2219 1774
rect 2295 1778 2299 1779
rect 2295 1773 2299 1774
rect 2319 1778 2323 1779
rect 2319 1773 2323 1774
rect 2375 1778 2379 1779
rect 2375 1773 2379 1774
rect 2439 1778 2443 1779
rect 2439 1773 2443 1774
rect 2503 1778 2507 1779
rect 2503 1773 2507 1774
rect 1286 1772 1292 1773
rect 1328 1770 1330 1773
rect 1526 1772 1532 1773
rect 1326 1769 1332 1770
rect 1326 1765 1327 1769
rect 1331 1765 1332 1769
rect 1526 1768 1527 1772
rect 1531 1768 1532 1772
rect 1526 1767 1532 1768
rect 1606 1772 1612 1773
rect 1606 1768 1607 1772
rect 1611 1768 1612 1772
rect 1606 1767 1612 1768
rect 1694 1772 1700 1773
rect 1694 1768 1695 1772
rect 1699 1768 1700 1772
rect 1694 1767 1700 1768
rect 1790 1772 1796 1773
rect 1790 1768 1791 1772
rect 1795 1768 1796 1772
rect 1790 1767 1796 1768
rect 1878 1772 1884 1773
rect 1878 1768 1879 1772
rect 1883 1768 1884 1772
rect 1878 1767 1884 1768
rect 1966 1772 1972 1773
rect 1966 1768 1967 1772
rect 1971 1768 1972 1772
rect 1966 1767 1972 1768
rect 2054 1772 2060 1773
rect 2054 1768 2055 1772
rect 2059 1768 2060 1772
rect 2054 1767 2060 1768
rect 2134 1772 2140 1773
rect 2134 1768 2135 1772
rect 2139 1768 2140 1772
rect 2134 1767 2140 1768
rect 2214 1772 2220 1773
rect 2214 1768 2215 1772
rect 2219 1768 2220 1772
rect 2214 1767 2220 1768
rect 2294 1772 2300 1773
rect 2294 1768 2295 1772
rect 2299 1768 2300 1772
rect 2294 1767 2300 1768
rect 2374 1772 2380 1773
rect 2374 1768 2375 1772
rect 2379 1768 2380 1772
rect 2374 1767 2380 1768
rect 2438 1772 2444 1773
rect 2438 1768 2439 1772
rect 2443 1768 2444 1772
rect 2504 1770 2506 1773
rect 2438 1767 2444 1768
rect 2502 1769 2508 1770
rect 1326 1764 1332 1765
rect 2502 1765 2503 1769
rect 2507 1765 2508 1769
rect 2502 1764 2508 1765
rect 110 1760 116 1761
rect 1286 1760 1292 1761
rect 110 1756 111 1760
rect 115 1756 116 1760
rect 110 1755 116 1756
rect 150 1759 156 1760
rect 150 1755 151 1759
rect 155 1755 156 1759
rect 112 1731 114 1755
rect 150 1754 156 1755
rect 214 1759 220 1760
rect 214 1755 215 1759
rect 219 1755 220 1759
rect 214 1754 220 1755
rect 310 1759 316 1760
rect 310 1755 311 1759
rect 315 1755 316 1759
rect 310 1754 316 1755
rect 414 1759 420 1760
rect 414 1755 415 1759
rect 419 1755 420 1759
rect 414 1754 420 1755
rect 518 1759 524 1760
rect 518 1755 519 1759
rect 523 1755 524 1759
rect 518 1754 524 1755
rect 622 1759 628 1760
rect 622 1755 623 1759
rect 627 1755 628 1759
rect 622 1754 628 1755
rect 718 1759 724 1760
rect 718 1755 719 1759
rect 723 1755 724 1759
rect 718 1754 724 1755
rect 814 1759 820 1760
rect 814 1755 815 1759
rect 819 1755 820 1759
rect 814 1754 820 1755
rect 902 1759 908 1760
rect 902 1755 903 1759
rect 907 1755 908 1759
rect 902 1754 908 1755
rect 990 1759 996 1760
rect 990 1755 991 1759
rect 995 1755 996 1759
rect 990 1754 996 1755
rect 1078 1759 1084 1760
rect 1078 1755 1079 1759
rect 1083 1755 1084 1759
rect 1078 1754 1084 1755
rect 1166 1759 1172 1760
rect 1166 1755 1167 1759
rect 1171 1755 1172 1759
rect 1286 1756 1287 1760
rect 1291 1756 1292 1760
rect 1286 1755 1292 1756
rect 1166 1754 1172 1755
rect 152 1731 154 1754
rect 216 1731 218 1754
rect 312 1731 314 1754
rect 416 1731 418 1754
rect 520 1731 522 1754
rect 624 1731 626 1754
rect 720 1731 722 1754
rect 816 1731 818 1754
rect 904 1731 906 1754
rect 992 1731 994 1754
rect 1080 1731 1082 1754
rect 1168 1731 1170 1754
rect 1288 1731 1290 1755
rect 1326 1752 1332 1753
rect 2502 1752 2508 1753
rect 1326 1748 1327 1752
rect 1331 1748 1332 1752
rect 1326 1747 1332 1748
rect 1542 1751 1548 1752
rect 1542 1747 1543 1751
rect 1547 1747 1548 1751
rect 111 1730 115 1731
rect 111 1725 115 1726
rect 151 1730 155 1731
rect 151 1725 155 1726
rect 167 1730 171 1731
rect 167 1725 171 1726
rect 215 1730 219 1731
rect 215 1725 219 1726
rect 239 1730 243 1731
rect 239 1725 243 1726
rect 311 1730 315 1731
rect 311 1725 315 1726
rect 319 1730 323 1731
rect 319 1725 323 1726
rect 407 1730 411 1731
rect 407 1725 411 1726
rect 415 1730 419 1731
rect 415 1725 419 1726
rect 503 1730 507 1731
rect 503 1725 507 1726
rect 519 1730 523 1731
rect 519 1725 523 1726
rect 607 1730 611 1731
rect 607 1725 611 1726
rect 623 1730 627 1731
rect 623 1725 627 1726
rect 711 1730 715 1731
rect 711 1725 715 1726
rect 719 1730 723 1731
rect 719 1725 723 1726
rect 815 1730 819 1731
rect 815 1725 819 1726
rect 823 1730 827 1731
rect 823 1725 827 1726
rect 903 1730 907 1731
rect 903 1725 907 1726
rect 935 1730 939 1731
rect 935 1725 939 1726
rect 991 1730 995 1731
rect 991 1725 995 1726
rect 1047 1730 1051 1731
rect 1047 1725 1051 1726
rect 1079 1730 1083 1731
rect 1079 1725 1083 1726
rect 1159 1730 1163 1731
rect 1159 1725 1163 1726
rect 1167 1730 1171 1731
rect 1167 1725 1171 1726
rect 1287 1730 1291 1731
rect 1287 1725 1291 1726
rect 112 1705 114 1725
rect 168 1706 170 1725
rect 240 1706 242 1725
rect 320 1706 322 1725
rect 408 1706 410 1725
rect 504 1706 506 1725
rect 608 1706 610 1725
rect 712 1706 714 1725
rect 824 1706 826 1725
rect 936 1706 938 1725
rect 1048 1706 1050 1725
rect 1160 1706 1162 1725
rect 166 1705 172 1706
rect 110 1704 116 1705
rect 110 1700 111 1704
rect 115 1700 116 1704
rect 166 1701 167 1705
rect 171 1701 172 1705
rect 166 1700 172 1701
rect 238 1705 244 1706
rect 238 1701 239 1705
rect 243 1701 244 1705
rect 238 1700 244 1701
rect 318 1705 324 1706
rect 318 1701 319 1705
rect 323 1701 324 1705
rect 318 1700 324 1701
rect 406 1705 412 1706
rect 406 1701 407 1705
rect 411 1701 412 1705
rect 406 1700 412 1701
rect 502 1705 508 1706
rect 502 1701 503 1705
rect 507 1701 508 1705
rect 502 1700 508 1701
rect 606 1705 612 1706
rect 606 1701 607 1705
rect 611 1701 612 1705
rect 606 1700 612 1701
rect 710 1705 716 1706
rect 710 1701 711 1705
rect 715 1701 716 1705
rect 710 1700 716 1701
rect 822 1705 828 1706
rect 822 1701 823 1705
rect 827 1701 828 1705
rect 822 1700 828 1701
rect 934 1705 940 1706
rect 934 1701 935 1705
rect 939 1701 940 1705
rect 934 1700 940 1701
rect 1046 1705 1052 1706
rect 1046 1701 1047 1705
rect 1051 1701 1052 1705
rect 1046 1700 1052 1701
rect 1158 1705 1164 1706
rect 1288 1705 1290 1725
rect 1328 1723 1330 1747
rect 1542 1746 1548 1747
rect 1622 1751 1628 1752
rect 1622 1747 1623 1751
rect 1627 1747 1628 1751
rect 1622 1746 1628 1747
rect 1710 1751 1716 1752
rect 1710 1747 1711 1751
rect 1715 1747 1716 1751
rect 1710 1746 1716 1747
rect 1806 1751 1812 1752
rect 1806 1747 1807 1751
rect 1811 1747 1812 1751
rect 1806 1746 1812 1747
rect 1894 1751 1900 1752
rect 1894 1747 1895 1751
rect 1899 1747 1900 1751
rect 1894 1746 1900 1747
rect 1982 1751 1988 1752
rect 1982 1747 1983 1751
rect 1987 1747 1988 1751
rect 1982 1746 1988 1747
rect 2070 1751 2076 1752
rect 2070 1747 2071 1751
rect 2075 1747 2076 1751
rect 2070 1746 2076 1747
rect 2150 1751 2156 1752
rect 2150 1747 2151 1751
rect 2155 1747 2156 1751
rect 2150 1746 2156 1747
rect 2230 1751 2236 1752
rect 2230 1747 2231 1751
rect 2235 1747 2236 1751
rect 2230 1746 2236 1747
rect 2310 1751 2316 1752
rect 2310 1747 2311 1751
rect 2315 1747 2316 1751
rect 2310 1746 2316 1747
rect 2390 1751 2396 1752
rect 2390 1747 2391 1751
rect 2395 1747 2396 1751
rect 2390 1746 2396 1747
rect 2454 1751 2460 1752
rect 2454 1747 2455 1751
rect 2459 1747 2460 1751
rect 2502 1748 2503 1752
rect 2507 1748 2508 1752
rect 2502 1747 2508 1748
rect 2454 1746 2460 1747
rect 1544 1723 1546 1746
rect 1624 1723 1626 1746
rect 1712 1723 1714 1746
rect 1808 1723 1810 1746
rect 1896 1723 1898 1746
rect 1984 1723 1986 1746
rect 2072 1723 2074 1746
rect 2152 1723 2154 1746
rect 2232 1723 2234 1746
rect 2312 1723 2314 1746
rect 2392 1723 2394 1746
rect 2456 1723 2458 1746
rect 2504 1723 2506 1747
rect 1327 1722 1331 1723
rect 1327 1717 1331 1718
rect 1399 1722 1403 1723
rect 1399 1717 1403 1718
rect 1463 1722 1467 1723
rect 1463 1717 1467 1718
rect 1543 1722 1547 1723
rect 1543 1717 1547 1718
rect 1623 1722 1627 1723
rect 1623 1717 1627 1718
rect 1631 1722 1635 1723
rect 1631 1717 1635 1718
rect 1711 1722 1715 1723
rect 1711 1717 1715 1718
rect 1727 1722 1731 1723
rect 1727 1717 1731 1718
rect 1807 1722 1811 1723
rect 1807 1717 1811 1718
rect 1823 1722 1827 1723
rect 1823 1717 1827 1718
rect 1895 1722 1899 1723
rect 1895 1717 1899 1718
rect 1919 1722 1923 1723
rect 1919 1717 1923 1718
rect 1983 1722 1987 1723
rect 1983 1717 1987 1718
rect 2015 1722 2019 1723
rect 2015 1717 2019 1718
rect 2071 1722 2075 1723
rect 2071 1717 2075 1718
rect 2111 1722 2115 1723
rect 2111 1717 2115 1718
rect 2151 1722 2155 1723
rect 2151 1717 2155 1718
rect 2199 1722 2203 1723
rect 2199 1717 2203 1718
rect 2231 1722 2235 1723
rect 2231 1717 2235 1718
rect 2287 1722 2291 1723
rect 2287 1717 2291 1718
rect 2311 1722 2315 1723
rect 2311 1717 2315 1718
rect 2383 1722 2387 1723
rect 2383 1717 2387 1718
rect 2391 1722 2395 1723
rect 2391 1717 2395 1718
rect 2455 1722 2459 1723
rect 2455 1717 2459 1718
rect 2503 1722 2507 1723
rect 2503 1717 2507 1718
rect 1158 1701 1159 1705
rect 1163 1701 1164 1705
rect 1158 1700 1164 1701
rect 1286 1704 1292 1705
rect 1286 1700 1287 1704
rect 1291 1700 1292 1704
rect 110 1699 116 1700
rect 1286 1699 1292 1700
rect 1328 1697 1330 1717
rect 1400 1698 1402 1717
rect 1464 1698 1466 1717
rect 1544 1698 1546 1717
rect 1632 1698 1634 1717
rect 1728 1698 1730 1717
rect 1824 1698 1826 1717
rect 1920 1698 1922 1717
rect 2016 1698 2018 1717
rect 2112 1698 2114 1717
rect 2200 1698 2202 1717
rect 2288 1698 2290 1717
rect 2384 1698 2386 1717
rect 2456 1698 2458 1717
rect 1398 1697 1404 1698
rect 1326 1696 1332 1697
rect 1326 1692 1327 1696
rect 1331 1692 1332 1696
rect 1398 1693 1399 1697
rect 1403 1693 1404 1697
rect 1398 1692 1404 1693
rect 1462 1697 1468 1698
rect 1462 1693 1463 1697
rect 1467 1693 1468 1697
rect 1462 1692 1468 1693
rect 1542 1697 1548 1698
rect 1542 1693 1543 1697
rect 1547 1693 1548 1697
rect 1542 1692 1548 1693
rect 1630 1697 1636 1698
rect 1630 1693 1631 1697
rect 1635 1693 1636 1697
rect 1630 1692 1636 1693
rect 1726 1697 1732 1698
rect 1726 1693 1727 1697
rect 1731 1693 1732 1697
rect 1726 1692 1732 1693
rect 1822 1697 1828 1698
rect 1822 1693 1823 1697
rect 1827 1693 1828 1697
rect 1822 1692 1828 1693
rect 1918 1697 1924 1698
rect 1918 1693 1919 1697
rect 1923 1693 1924 1697
rect 1918 1692 1924 1693
rect 2014 1697 2020 1698
rect 2014 1693 2015 1697
rect 2019 1693 2020 1697
rect 2014 1692 2020 1693
rect 2110 1697 2116 1698
rect 2110 1693 2111 1697
rect 2115 1693 2116 1697
rect 2110 1692 2116 1693
rect 2198 1697 2204 1698
rect 2198 1693 2199 1697
rect 2203 1693 2204 1697
rect 2198 1692 2204 1693
rect 2286 1697 2292 1698
rect 2286 1693 2287 1697
rect 2291 1693 2292 1697
rect 2286 1692 2292 1693
rect 2382 1697 2388 1698
rect 2382 1693 2383 1697
rect 2387 1693 2388 1697
rect 2382 1692 2388 1693
rect 2454 1697 2460 1698
rect 2504 1697 2506 1717
rect 2454 1693 2455 1697
rect 2459 1693 2460 1697
rect 2454 1692 2460 1693
rect 2502 1696 2508 1697
rect 2502 1692 2503 1696
rect 2507 1692 2508 1696
rect 1326 1691 1332 1692
rect 2502 1691 2508 1692
rect 110 1687 116 1688
rect 110 1683 111 1687
rect 115 1683 116 1687
rect 1286 1687 1292 1688
rect 110 1682 116 1683
rect 150 1684 156 1685
rect 112 1675 114 1682
rect 150 1680 151 1684
rect 155 1680 156 1684
rect 150 1679 156 1680
rect 222 1684 228 1685
rect 222 1680 223 1684
rect 227 1680 228 1684
rect 222 1679 228 1680
rect 302 1684 308 1685
rect 302 1680 303 1684
rect 307 1680 308 1684
rect 302 1679 308 1680
rect 390 1684 396 1685
rect 390 1680 391 1684
rect 395 1680 396 1684
rect 390 1679 396 1680
rect 486 1684 492 1685
rect 486 1680 487 1684
rect 491 1680 492 1684
rect 486 1679 492 1680
rect 590 1684 596 1685
rect 590 1680 591 1684
rect 595 1680 596 1684
rect 590 1679 596 1680
rect 694 1684 700 1685
rect 694 1680 695 1684
rect 699 1680 700 1684
rect 694 1679 700 1680
rect 806 1684 812 1685
rect 806 1680 807 1684
rect 811 1680 812 1684
rect 806 1679 812 1680
rect 918 1684 924 1685
rect 918 1680 919 1684
rect 923 1680 924 1684
rect 918 1679 924 1680
rect 1030 1684 1036 1685
rect 1030 1680 1031 1684
rect 1035 1680 1036 1684
rect 1030 1679 1036 1680
rect 1142 1684 1148 1685
rect 1142 1680 1143 1684
rect 1147 1680 1148 1684
rect 1286 1683 1287 1687
rect 1291 1683 1292 1687
rect 1286 1682 1292 1683
rect 1142 1679 1148 1680
rect 152 1675 154 1679
rect 224 1675 226 1679
rect 304 1675 306 1679
rect 392 1675 394 1679
rect 488 1675 490 1679
rect 592 1675 594 1679
rect 696 1675 698 1679
rect 808 1675 810 1679
rect 920 1675 922 1679
rect 1032 1675 1034 1679
rect 1144 1675 1146 1679
rect 1288 1675 1290 1682
rect 1326 1679 1332 1680
rect 1326 1675 1327 1679
rect 1331 1675 1332 1679
rect 2502 1679 2508 1680
rect 111 1674 115 1675
rect 111 1669 115 1670
rect 151 1674 155 1675
rect 151 1669 155 1670
rect 223 1674 227 1675
rect 223 1669 227 1670
rect 255 1674 259 1675
rect 255 1669 259 1670
rect 303 1674 307 1675
rect 303 1669 307 1670
rect 319 1674 323 1675
rect 319 1669 323 1670
rect 391 1674 395 1675
rect 391 1669 395 1670
rect 399 1674 403 1675
rect 399 1669 403 1670
rect 487 1674 491 1675
rect 487 1669 491 1670
rect 575 1674 579 1675
rect 575 1669 579 1670
rect 591 1674 595 1675
rect 591 1669 595 1670
rect 671 1674 675 1675
rect 671 1669 675 1670
rect 695 1674 699 1675
rect 695 1669 699 1670
rect 767 1674 771 1675
rect 767 1669 771 1670
rect 807 1674 811 1675
rect 807 1669 811 1670
rect 863 1674 867 1675
rect 863 1669 867 1670
rect 919 1674 923 1675
rect 919 1669 923 1670
rect 959 1674 963 1675
rect 959 1669 963 1670
rect 1031 1674 1035 1675
rect 1031 1669 1035 1670
rect 1063 1674 1067 1675
rect 1063 1669 1067 1670
rect 1143 1674 1147 1675
rect 1143 1669 1147 1670
rect 1167 1674 1171 1675
rect 1167 1669 1171 1670
rect 1287 1674 1291 1675
rect 1326 1674 1332 1675
rect 1382 1676 1388 1677
rect 1287 1669 1291 1670
rect 112 1666 114 1669
rect 254 1668 260 1669
rect 110 1665 116 1666
rect 110 1661 111 1665
rect 115 1661 116 1665
rect 254 1664 255 1668
rect 259 1664 260 1668
rect 254 1663 260 1664
rect 318 1668 324 1669
rect 318 1664 319 1668
rect 323 1664 324 1668
rect 318 1663 324 1664
rect 398 1668 404 1669
rect 398 1664 399 1668
rect 403 1664 404 1668
rect 398 1663 404 1664
rect 486 1668 492 1669
rect 486 1664 487 1668
rect 491 1664 492 1668
rect 486 1663 492 1664
rect 574 1668 580 1669
rect 574 1664 575 1668
rect 579 1664 580 1668
rect 574 1663 580 1664
rect 670 1668 676 1669
rect 670 1664 671 1668
rect 675 1664 676 1668
rect 670 1663 676 1664
rect 766 1668 772 1669
rect 766 1664 767 1668
rect 771 1664 772 1668
rect 766 1663 772 1664
rect 862 1668 868 1669
rect 862 1664 863 1668
rect 867 1664 868 1668
rect 862 1663 868 1664
rect 958 1668 964 1669
rect 958 1664 959 1668
rect 963 1664 964 1668
rect 958 1663 964 1664
rect 1062 1668 1068 1669
rect 1062 1664 1063 1668
rect 1067 1664 1068 1668
rect 1062 1663 1068 1664
rect 1166 1668 1172 1669
rect 1166 1664 1167 1668
rect 1171 1664 1172 1668
rect 1288 1666 1290 1669
rect 1328 1667 1330 1674
rect 1382 1672 1383 1676
rect 1387 1672 1388 1676
rect 1382 1671 1388 1672
rect 1446 1676 1452 1677
rect 1446 1672 1447 1676
rect 1451 1672 1452 1676
rect 1446 1671 1452 1672
rect 1526 1676 1532 1677
rect 1526 1672 1527 1676
rect 1531 1672 1532 1676
rect 1526 1671 1532 1672
rect 1614 1676 1620 1677
rect 1614 1672 1615 1676
rect 1619 1672 1620 1676
rect 1614 1671 1620 1672
rect 1710 1676 1716 1677
rect 1710 1672 1711 1676
rect 1715 1672 1716 1676
rect 1710 1671 1716 1672
rect 1806 1676 1812 1677
rect 1806 1672 1807 1676
rect 1811 1672 1812 1676
rect 1806 1671 1812 1672
rect 1902 1676 1908 1677
rect 1902 1672 1903 1676
rect 1907 1672 1908 1676
rect 1902 1671 1908 1672
rect 1998 1676 2004 1677
rect 1998 1672 1999 1676
rect 2003 1672 2004 1676
rect 1998 1671 2004 1672
rect 2094 1676 2100 1677
rect 2094 1672 2095 1676
rect 2099 1672 2100 1676
rect 2094 1671 2100 1672
rect 2182 1676 2188 1677
rect 2182 1672 2183 1676
rect 2187 1672 2188 1676
rect 2182 1671 2188 1672
rect 2270 1676 2276 1677
rect 2270 1672 2271 1676
rect 2275 1672 2276 1676
rect 2270 1671 2276 1672
rect 2366 1676 2372 1677
rect 2366 1672 2367 1676
rect 2371 1672 2372 1676
rect 2366 1671 2372 1672
rect 2438 1676 2444 1677
rect 2438 1672 2439 1676
rect 2443 1672 2444 1676
rect 2502 1675 2503 1679
rect 2507 1675 2508 1679
rect 2502 1674 2508 1675
rect 2438 1671 2444 1672
rect 1384 1667 1386 1671
rect 1448 1667 1450 1671
rect 1528 1667 1530 1671
rect 1616 1667 1618 1671
rect 1712 1667 1714 1671
rect 1808 1667 1810 1671
rect 1904 1667 1906 1671
rect 2000 1667 2002 1671
rect 2096 1667 2098 1671
rect 2184 1667 2186 1671
rect 2272 1667 2274 1671
rect 2368 1667 2370 1671
rect 2440 1667 2442 1671
rect 2504 1667 2506 1674
rect 1327 1666 1331 1667
rect 1166 1663 1172 1664
rect 1286 1665 1292 1666
rect 110 1660 116 1661
rect 1286 1661 1287 1665
rect 1291 1661 1292 1665
rect 1327 1661 1331 1662
rect 1351 1666 1355 1667
rect 1351 1661 1355 1662
rect 1383 1666 1387 1667
rect 1383 1661 1387 1662
rect 1407 1666 1411 1667
rect 1407 1661 1411 1662
rect 1447 1666 1451 1667
rect 1447 1661 1451 1662
rect 1495 1666 1499 1667
rect 1495 1661 1499 1662
rect 1527 1666 1531 1667
rect 1527 1661 1531 1662
rect 1583 1666 1587 1667
rect 1583 1661 1587 1662
rect 1615 1666 1619 1667
rect 1615 1661 1619 1662
rect 1679 1666 1683 1667
rect 1679 1661 1683 1662
rect 1711 1666 1715 1667
rect 1711 1661 1715 1662
rect 1783 1666 1787 1667
rect 1783 1661 1787 1662
rect 1807 1666 1811 1667
rect 1807 1661 1811 1662
rect 1895 1666 1899 1667
rect 1895 1661 1899 1662
rect 1903 1666 1907 1667
rect 1903 1661 1907 1662
rect 1999 1666 2003 1667
rect 1999 1661 2003 1662
rect 2023 1666 2027 1667
rect 2023 1661 2027 1662
rect 2095 1666 2099 1667
rect 2095 1661 2099 1662
rect 2159 1666 2163 1667
rect 2159 1661 2163 1662
rect 2183 1666 2187 1667
rect 2183 1661 2187 1662
rect 2271 1666 2275 1667
rect 2271 1661 2275 1662
rect 2303 1666 2307 1667
rect 2303 1661 2307 1662
rect 2367 1666 2371 1667
rect 2367 1661 2371 1662
rect 2439 1666 2443 1667
rect 2439 1661 2443 1662
rect 2503 1666 2507 1667
rect 2503 1661 2507 1662
rect 1286 1660 1292 1661
rect 1328 1658 1330 1661
rect 1350 1660 1356 1661
rect 1326 1657 1332 1658
rect 1326 1653 1327 1657
rect 1331 1653 1332 1657
rect 1350 1656 1351 1660
rect 1355 1656 1356 1660
rect 1350 1655 1356 1656
rect 1406 1660 1412 1661
rect 1406 1656 1407 1660
rect 1411 1656 1412 1660
rect 1406 1655 1412 1656
rect 1494 1660 1500 1661
rect 1494 1656 1495 1660
rect 1499 1656 1500 1660
rect 1494 1655 1500 1656
rect 1582 1660 1588 1661
rect 1582 1656 1583 1660
rect 1587 1656 1588 1660
rect 1582 1655 1588 1656
rect 1678 1660 1684 1661
rect 1678 1656 1679 1660
rect 1683 1656 1684 1660
rect 1678 1655 1684 1656
rect 1782 1660 1788 1661
rect 1782 1656 1783 1660
rect 1787 1656 1788 1660
rect 1782 1655 1788 1656
rect 1894 1660 1900 1661
rect 1894 1656 1895 1660
rect 1899 1656 1900 1660
rect 1894 1655 1900 1656
rect 2022 1660 2028 1661
rect 2022 1656 2023 1660
rect 2027 1656 2028 1660
rect 2022 1655 2028 1656
rect 2158 1660 2164 1661
rect 2158 1656 2159 1660
rect 2163 1656 2164 1660
rect 2158 1655 2164 1656
rect 2302 1660 2308 1661
rect 2302 1656 2303 1660
rect 2307 1656 2308 1660
rect 2302 1655 2308 1656
rect 2438 1660 2444 1661
rect 2438 1656 2439 1660
rect 2443 1656 2444 1660
rect 2504 1658 2506 1661
rect 2438 1655 2444 1656
rect 2502 1657 2508 1658
rect 1326 1652 1332 1653
rect 2502 1653 2503 1657
rect 2507 1653 2508 1657
rect 2502 1652 2508 1653
rect 110 1648 116 1649
rect 1286 1648 1292 1649
rect 110 1644 111 1648
rect 115 1644 116 1648
rect 110 1643 116 1644
rect 270 1647 276 1648
rect 270 1643 271 1647
rect 275 1643 276 1647
rect 112 1619 114 1643
rect 270 1642 276 1643
rect 334 1647 340 1648
rect 334 1643 335 1647
rect 339 1643 340 1647
rect 334 1642 340 1643
rect 414 1647 420 1648
rect 414 1643 415 1647
rect 419 1643 420 1647
rect 414 1642 420 1643
rect 502 1647 508 1648
rect 502 1643 503 1647
rect 507 1643 508 1647
rect 502 1642 508 1643
rect 590 1647 596 1648
rect 590 1643 591 1647
rect 595 1643 596 1647
rect 590 1642 596 1643
rect 686 1647 692 1648
rect 686 1643 687 1647
rect 691 1643 692 1647
rect 686 1642 692 1643
rect 782 1647 788 1648
rect 782 1643 783 1647
rect 787 1643 788 1647
rect 782 1642 788 1643
rect 878 1647 884 1648
rect 878 1643 879 1647
rect 883 1643 884 1647
rect 878 1642 884 1643
rect 974 1647 980 1648
rect 974 1643 975 1647
rect 979 1643 980 1647
rect 974 1642 980 1643
rect 1078 1647 1084 1648
rect 1078 1643 1079 1647
rect 1083 1643 1084 1647
rect 1078 1642 1084 1643
rect 1182 1647 1188 1648
rect 1182 1643 1183 1647
rect 1187 1643 1188 1647
rect 1286 1644 1287 1648
rect 1291 1644 1292 1648
rect 1286 1643 1292 1644
rect 1182 1642 1188 1643
rect 272 1619 274 1642
rect 336 1619 338 1642
rect 416 1619 418 1642
rect 504 1619 506 1642
rect 592 1619 594 1642
rect 688 1619 690 1642
rect 784 1619 786 1642
rect 880 1619 882 1642
rect 976 1619 978 1642
rect 1080 1619 1082 1642
rect 1184 1619 1186 1642
rect 1288 1619 1290 1643
rect 1326 1640 1332 1641
rect 2502 1640 2508 1641
rect 1326 1636 1327 1640
rect 1331 1636 1332 1640
rect 1326 1635 1332 1636
rect 1366 1639 1372 1640
rect 1366 1635 1367 1639
rect 1371 1635 1372 1639
rect 111 1618 115 1619
rect 111 1613 115 1614
rect 271 1618 275 1619
rect 271 1613 275 1614
rect 303 1618 307 1619
rect 303 1613 307 1614
rect 335 1618 339 1619
rect 335 1613 339 1614
rect 359 1618 363 1619
rect 359 1613 363 1614
rect 415 1618 419 1619
rect 415 1613 419 1614
rect 431 1618 435 1619
rect 431 1613 435 1614
rect 503 1618 507 1619
rect 503 1613 507 1614
rect 511 1618 515 1619
rect 511 1613 515 1614
rect 591 1618 595 1619
rect 591 1613 595 1614
rect 599 1618 603 1619
rect 599 1613 603 1614
rect 687 1618 691 1619
rect 687 1613 691 1614
rect 695 1618 699 1619
rect 695 1613 699 1614
rect 783 1618 787 1619
rect 783 1613 787 1614
rect 791 1618 795 1619
rect 791 1613 795 1614
rect 879 1618 883 1619
rect 879 1613 883 1614
rect 895 1618 899 1619
rect 895 1613 899 1614
rect 975 1618 979 1619
rect 975 1613 979 1614
rect 1007 1618 1011 1619
rect 1007 1613 1011 1614
rect 1079 1618 1083 1619
rect 1079 1613 1083 1614
rect 1119 1618 1123 1619
rect 1119 1613 1123 1614
rect 1183 1618 1187 1619
rect 1183 1613 1187 1614
rect 1287 1618 1291 1619
rect 1328 1615 1330 1635
rect 1366 1634 1372 1635
rect 1422 1639 1428 1640
rect 1422 1635 1423 1639
rect 1427 1635 1428 1639
rect 1422 1634 1428 1635
rect 1510 1639 1516 1640
rect 1510 1635 1511 1639
rect 1515 1635 1516 1639
rect 1510 1634 1516 1635
rect 1598 1639 1604 1640
rect 1598 1635 1599 1639
rect 1603 1635 1604 1639
rect 1598 1634 1604 1635
rect 1694 1639 1700 1640
rect 1694 1635 1695 1639
rect 1699 1635 1700 1639
rect 1694 1634 1700 1635
rect 1798 1639 1804 1640
rect 1798 1635 1799 1639
rect 1803 1635 1804 1639
rect 1798 1634 1804 1635
rect 1910 1639 1916 1640
rect 1910 1635 1911 1639
rect 1915 1635 1916 1639
rect 1910 1634 1916 1635
rect 2038 1639 2044 1640
rect 2038 1635 2039 1639
rect 2043 1635 2044 1639
rect 2038 1634 2044 1635
rect 2174 1639 2180 1640
rect 2174 1635 2175 1639
rect 2179 1635 2180 1639
rect 2174 1634 2180 1635
rect 2318 1639 2324 1640
rect 2318 1635 2319 1639
rect 2323 1635 2324 1639
rect 2318 1634 2324 1635
rect 2454 1639 2460 1640
rect 2454 1635 2455 1639
rect 2459 1635 2460 1639
rect 2502 1636 2503 1640
rect 2507 1636 2508 1640
rect 2502 1635 2508 1636
rect 2454 1634 2460 1635
rect 1368 1615 1370 1634
rect 1424 1615 1426 1634
rect 1512 1615 1514 1634
rect 1600 1615 1602 1634
rect 1696 1615 1698 1634
rect 1800 1615 1802 1634
rect 1912 1615 1914 1634
rect 2040 1615 2042 1634
rect 2176 1615 2178 1634
rect 2320 1615 2322 1634
rect 2456 1615 2458 1634
rect 2504 1615 2506 1635
rect 1287 1613 1291 1614
rect 1327 1614 1331 1615
rect 112 1593 114 1613
rect 304 1594 306 1613
rect 360 1594 362 1613
rect 432 1594 434 1613
rect 512 1594 514 1613
rect 600 1594 602 1613
rect 696 1594 698 1613
rect 792 1594 794 1613
rect 896 1594 898 1613
rect 1008 1594 1010 1613
rect 1120 1594 1122 1613
rect 302 1593 308 1594
rect 110 1592 116 1593
rect 110 1588 111 1592
rect 115 1588 116 1592
rect 302 1589 303 1593
rect 307 1589 308 1593
rect 302 1588 308 1589
rect 358 1593 364 1594
rect 358 1589 359 1593
rect 363 1589 364 1593
rect 358 1588 364 1589
rect 430 1593 436 1594
rect 430 1589 431 1593
rect 435 1589 436 1593
rect 430 1588 436 1589
rect 510 1593 516 1594
rect 510 1589 511 1593
rect 515 1589 516 1593
rect 510 1588 516 1589
rect 598 1593 604 1594
rect 598 1589 599 1593
rect 603 1589 604 1593
rect 598 1588 604 1589
rect 694 1593 700 1594
rect 694 1589 695 1593
rect 699 1589 700 1593
rect 694 1588 700 1589
rect 790 1593 796 1594
rect 790 1589 791 1593
rect 795 1589 796 1593
rect 790 1588 796 1589
rect 894 1593 900 1594
rect 894 1589 895 1593
rect 899 1589 900 1593
rect 894 1588 900 1589
rect 1006 1593 1012 1594
rect 1006 1589 1007 1593
rect 1011 1589 1012 1593
rect 1006 1588 1012 1589
rect 1118 1593 1124 1594
rect 1288 1593 1290 1613
rect 1327 1609 1331 1610
rect 1367 1614 1371 1615
rect 1367 1609 1371 1610
rect 1423 1614 1427 1615
rect 1423 1609 1427 1610
rect 1479 1614 1483 1615
rect 1479 1609 1483 1610
rect 1511 1614 1515 1615
rect 1511 1609 1515 1610
rect 1559 1614 1563 1615
rect 1559 1609 1563 1610
rect 1599 1614 1603 1615
rect 1599 1609 1603 1610
rect 1639 1614 1643 1615
rect 1639 1609 1643 1610
rect 1695 1614 1699 1615
rect 1695 1609 1699 1610
rect 1719 1614 1723 1615
rect 1719 1609 1723 1610
rect 1791 1614 1795 1615
rect 1791 1609 1795 1610
rect 1799 1614 1803 1615
rect 1799 1609 1803 1610
rect 1871 1614 1875 1615
rect 1871 1609 1875 1610
rect 1911 1614 1915 1615
rect 1911 1609 1915 1610
rect 1951 1614 1955 1615
rect 1951 1609 1955 1610
rect 2031 1614 2035 1615
rect 2031 1609 2035 1610
rect 2039 1614 2043 1615
rect 2039 1609 2043 1610
rect 2175 1614 2179 1615
rect 2175 1609 2179 1610
rect 2319 1614 2323 1615
rect 2319 1609 2323 1610
rect 2455 1614 2459 1615
rect 2455 1609 2459 1610
rect 2503 1614 2507 1615
rect 2503 1609 2507 1610
rect 1118 1589 1119 1593
rect 1123 1589 1124 1593
rect 1118 1588 1124 1589
rect 1286 1592 1292 1593
rect 1286 1588 1287 1592
rect 1291 1588 1292 1592
rect 1328 1589 1330 1609
rect 1368 1590 1370 1609
rect 1424 1590 1426 1609
rect 1480 1590 1482 1609
rect 1560 1590 1562 1609
rect 1640 1590 1642 1609
rect 1720 1590 1722 1609
rect 1792 1590 1794 1609
rect 1872 1590 1874 1609
rect 1952 1590 1954 1609
rect 2032 1590 2034 1609
rect 1366 1589 1372 1590
rect 110 1587 116 1588
rect 1286 1587 1292 1588
rect 1326 1588 1332 1589
rect 1326 1584 1327 1588
rect 1331 1584 1332 1588
rect 1366 1585 1367 1589
rect 1371 1585 1372 1589
rect 1366 1584 1372 1585
rect 1422 1589 1428 1590
rect 1422 1585 1423 1589
rect 1427 1585 1428 1589
rect 1422 1584 1428 1585
rect 1478 1589 1484 1590
rect 1478 1585 1479 1589
rect 1483 1585 1484 1589
rect 1478 1584 1484 1585
rect 1558 1589 1564 1590
rect 1558 1585 1559 1589
rect 1563 1585 1564 1589
rect 1558 1584 1564 1585
rect 1638 1589 1644 1590
rect 1638 1585 1639 1589
rect 1643 1585 1644 1589
rect 1638 1584 1644 1585
rect 1718 1589 1724 1590
rect 1718 1585 1719 1589
rect 1723 1585 1724 1589
rect 1718 1584 1724 1585
rect 1790 1589 1796 1590
rect 1790 1585 1791 1589
rect 1795 1585 1796 1589
rect 1790 1584 1796 1585
rect 1870 1589 1876 1590
rect 1870 1585 1871 1589
rect 1875 1585 1876 1589
rect 1870 1584 1876 1585
rect 1950 1589 1956 1590
rect 1950 1585 1951 1589
rect 1955 1585 1956 1589
rect 1950 1584 1956 1585
rect 2030 1589 2036 1590
rect 2504 1589 2506 1609
rect 2030 1585 2031 1589
rect 2035 1585 2036 1589
rect 2030 1584 2036 1585
rect 2502 1588 2508 1589
rect 2502 1584 2503 1588
rect 2507 1584 2508 1588
rect 1326 1583 1332 1584
rect 2502 1583 2508 1584
rect 110 1575 116 1576
rect 110 1571 111 1575
rect 115 1571 116 1575
rect 1286 1575 1292 1576
rect 110 1570 116 1571
rect 286 1572 292 1573
rect 112 1567 114 1570
rect 286 1568 287 1572
rect 291 1568 292 1572
rect 286 1567 292 1568
rect 342 1572 348 1573
rect 342 1568 343 1572
rect 347 1568 348 1572
rect 342 1567 348 1568
rect 414 1572 420 1573
rect 414 1568 415 1572
rect 419 1568 420 1572
rect 414 1567 420 1568
rect 494 1572 500 1573
rect 494 1568 495 1572
rect 499 1568 500 1572
rect 494 1567 500 1568
rect 582 1572 588 1573
rect 582 1568 583 1572
rect 587 1568 588 1572
rect 582 1567 588 1568
rect 678 1572 684 1573
rect 678 1568 679 1572
rect 683 1568 684 1572
rect 678 1567 684 1568
rect 774 1572 780 1573
rect 774 1568 775 1572
rect 779 1568 780 1572
rect 774 1567 780 1568
rect 878 1572 884 1573
rect 878 1568 879 1572
rect 883 1568 884 1572
rect 878 1567 884 1568
rect 990 1572 996 1573
rect 990 1568 991 1572
rect 995 1568 996 1572
rect 990 1567 996 1568
rect 1102 1572 1108 1573
rect 1102 1568 1103 1572
rect 1107 1568 1108 1572
rect 1286 1571 1287 1575
rect 1291 1571 1292 1575
rect 1286 1570 1292 1571
rect 1326 1571 1332 1572
rect 1102 1567 1108 1568
rect 1288 1567 1290 1570
rect 1326 1567 1327 1571
rect 1331 1567 1332 1571
rect 2502 1571 2508 1572
rect 111 1566 115 1567
rect 111 1561 115 1562
rect 247 1566 251 1567
rect 247 1561 251 1562
rect 287 1566 291 1567
rect 287 1561 291 1562
rect 319 1566 323 1567
rect 319 1561 323 1562
rect 343 1566 347 1567
rect 343 1561 347 1562
rect 399 1566 403 1567
rect 399 1561 403 1562
rect 415 1566 419 1567
rect 415 1561 419 1562
rect 487 1566 491 1567
rect 487 1561 491 1562
rect 495 1566 499 1567
rect 495 1561 499 1562
rect 583 1566 587 1567
rect 583 1561 587 1562
rect 671 1566 675 1567
rect 671 1561 675 1562
rect 679 1566 683 1567
rect 679 1561 683 1562
rect 759 1566 763 1567
rect 759 1561 763 1562
rect 775 1566 779 1567
rect 775 1561 779 1562
rect 847 1566 851 1567
rect 847 1561 851 1562
rect 879 1566 883 1567
rect 879 1561 883 1562
rect 927 1566 931 1567
rect 927 1561 931 1562
rect 991 1566 995 1567
rect 991 1561 995 1562
rect 1007 1566 1011 1567
rect 1007 1561 1011 1562
rect 1087 1566 1091 1567
rect 1087 1561 1091 1562
rect 1103 1566 1107 1567
rect 1103 1561 1107 1562
rect 1167 1566 1171 1567
rect 1167 1561 1171 1562
rect 1223 1566 1227 1567
rect 1223 1561 1227 1562
rect 1287 1566 1291 1567
rect 1326 1566 1332 1567
rect 1350 1568 1356 1569
rect 1328 1563 1330 1566
rect 1350 1564 1351 1568
rect 1355 1564 1356 1568
rect 1350 1563 1356 1564
rect 1406 1568 1412 1569
rect 1406 1564 1407 1568
rect 1411 1564 1412 1568
rect 1406 1563 1412 1564
rect 1462 1568 1468 1569
rect 1462 1564 1463 1568
rect 1467 1564 1468 1568
rect 1462 1563 1468 1564
rect 1542 1568 1548 1569
rect 1542 1564 1543 1568
rect 1547 1564 1548 1568
rect 1542 1563 1548 1564
rect 1622 1568 1628 1569
rect 1622 1564 1623 1568
rect 1627 1564 1628 1568
rect 1622 1563 1628 1564
rect 1702 1568 1708 1569
rect 1702 1564 1703 1568
rect 1707 1564 1708 1568
rect 1702 1563 1708 1564
rect 1774 1568 1780 1569
rect 1774 1564 1775 1568
rect 1779 1564 1780 1568
rect 1774 1563 1780 1564
rect 1854 1568 1860 1569
rect 1854 1564 1855 1568
rect 1859 1564 1860 1568
rect 1854 1563 1860 1564
rect 1934 1568 1940 1569
rect 1934 1564 1935 1568
rect 1939 1564 1940 1568
rect 1934 1563 1940 1564
rect 2014 1568 2020 1569
rect 2014 1564 2015 1568
rect 2019 1564 2020 1568
rect 2502 1567 2503 1571
rect 2507 1567 2508 1571
rect 2502 1566 2508 1567
rect 2014 1563 2020 1564
rect 2504 1563 2506 1566
rect 1287 1561 1291 1562
rect 1327 1562 1331 1563
rect 112 1558 114 1561
rect 246 1560 252 1561
rect 110 1557 116 1558
rect 110 1553 111 1557
rect 115 1553 116 1557
rect 246 1556 247 1560
rect 251 1556 252 1560
rect 246 1555 252 1556
rect 318 1560 324 1561
rect 318 1556 319 1560
rect 323 1556 324 1560
rect 318 1555 324 1556
rect 398 1560 404 1561
rect 398 1556 399 1560
rect 403 1556 404 1560
rect 398 1555 404 1556
rect 486 1560 492 1561
rect 486 1556 487 1560
rect 491 1556 492 1560
rect 486 1555 492 1556
rect 582 1560 588 1561
rect 582 1556 583 1560
rect 587 1556 588 1560
rect 582 1555 588 1556
rect 670 1560 676 1561
rect 670 1556 671 1560
rect 675 1556 676 1560
rect 670 1555 676 1556
rect 758 1560 764 1561
rect 758 1556 759 1560
rect 763 1556 764 1560
rect 758 1555 764 1556
rect 846 1560 852 1561
rect 846 1556 847 1560
rect 851 1556 852 1560
rect 846 1555 852 1556
rect 926 1560 932 1561
rect 926 1556 927 1560
rect 931 1556 932 1560
rect 926 1555 932 1556
rect 1006 1560 1012 1561
rect 1006 1556 1007 1560
rect 1011 1556 1012 1560
rect 1006 1555 1012 1556
rect 1086 1560 1092 1561
rect 1086 1556 1087 1560
rect 1091 1556 1092 1560
rect 1086 1555 1092 1556
rect 1166 1560 1172 1561
rect 1166 1556 1167 1560
rect 1171 1556 1172 1560
rect 1166 1555 1172 1556
rect 1222 1560 1228 1561
rect 1222 1556 1223 1560
rect 1227 1556 1228 1560
rect 1288 1558 1290 1561
rect 1222 1555 1228 1556
rect 1286 1557 1292 1558
rect 1327 1557 1331 1558
rect 1351 1562 1355 1563
rect 1351 1557 1355 1558
rect 1407 1562 1411 1563
rect 1407 1557 1411 1558
rect 1463 1562 1467 1563
rect 1463 1557 1467 1558
rect 1471 1562 1475 1563
rect 1471 1557 1475 1558
rect 1543 1562 1547 1563
rect 1543 1557 1547 1558
rect 1607 1562 1611 1563
rect 1607 1557 1611 1558
rect 1623 1562 1627 1563
rect 1623 1557 1627 1558
rect 1703 1562 1707 1563
rect 1703 1557 1707 1558
rect 1735 1562 1739 1563
rect 1735 1557 1739 1558
rect 1775 1562 1779 1563
rect 1775 1557 1779 1558
rect 1855 1562 1859 1563
rect 1855 1557 1859 1558
rect 1871 1562 1875 1563
rect 1871 1557 1875 1558
rect 1935 1562 1939 1563
rect 1935 1557 1939 1558
rect 2007 1562 2011 1563
rect 2007 1557 2011 1558
rect 2015 1562 2019 1563
rect 2015 1557 2019 1558
rect 2503 1562 2507 1563
rect 2503 1557 2507 1558
rect 110 1552 116 1553
rect 1286 1553 1287 1557
rect 1291 1553 1292 1557
rect 1328 1554 1330 1557
rect 1350 1556 1356 1557
rect 1286 1552 1292 1553
rect 1326 1553 1332 1554
rect 1326 1549 1327 1553
rect 1331 1549 1332 1553
rect 1350 1552 1351 1556
rect 1355 1552 1356 1556
rect 1350 1551 1356 1552
rect 1470 1556 1476 1557
rect 1470 1552 1471 1556
rect 1475 1552 1476 1556
rect 1470 1551 1476 1552
rect 1606 1556 1612 1557
rect 1606 1552 1607 1556
rect 1611 1552 1612 1556
rect 1606 1551 1612 1552
rect 1734 1556 1740 1557
rect 1734 1552 1735 1556
rect 1739 1552 1740 1556
rect 1734 1551 1740 1552
rect 1870 1556 1876 1557
rect 1870 1552 1871 1556
rect 1875 1552 1876 1556
rect 1870 1551 1876 1552
rect 2006 1556 2012 1557
rect 2006 1552 2007 1556
rect 2011 1552 2012 1556
rect 2504 1554 2506 1557
rect 2006 1551 2012 1552
rect 2502 1553 2508 1554
rect 1326 1548 1332 1549
rect 2502 1549 2503 1553
rect 2507 1549 2508 1553
rect 2502 1548 2508 1549
rect 110 1540 116 1541
rect 1286 1540 1292 1541
rect 110 1536 111 1540
rect 115 1536 116 1540
rect 110 1535 116 1536
rect 262 1539 268 1540
rect 262 1535 263 1539
rect 267 1535 268 1539
rect 112 1507 114 1535
rect 262 1534 268 1535
rect 334 1539 340 1540
rect 334 1535 335 1539
rect 339 1535 340 1539
rect 334 1534 340 1535
rect 414 1539 420 1540
rect 414 1535 415 1539
rect 419 1535 420 1539
rect 414 1534 420 1535
rect 502 1539 508 1540
rect 502 1535 503 1539
rect 507 1535 508 1539
rect 502 1534 508 1535
rect 598 1539 604 1540
rect 598 1535 599 1539
rect 603 1535 604 1539
rect 598 1534 604 1535
rect 686 1539 692 1540
rect 686 1535 687 1539
rect 691 1535 692 1539
rect 686 1534 692 1535
rect 774 1539 780 1540
rect 774 1535 775 1539
rect 779 1535 780 1539
rect 774 1534 780 1535
rect 862 1539 868 1540
rect 862 1535 863 1539
rect 867 1535 868 1539
rect 862 1534 868 1535
rect 942 1539 948 1540
rect 942 1535 943 1539
rect 947 1535 948 1539
rect 942 1534 948 1535
rect 1022 1539 1028 1540
rect 1022 1535 1023 1539
rect 1027 1535 1028 1539
rect 1022 1534 1028 1535
rect 1102 1539 1108 1540
rect 1102 1535 1103 1539
rect 1107 1535 1108 1539
rect 1102 1534 1108 1535
rect 1182 1539 1188 1540
rect 1182 1535 1183 1539
rect 1187 1535 1188 1539
rect 1182 1534 1188 1535
rect 1238 1539 1244 1540
rect 1238 1535 1239 1539
rect 1243 1535 1244 1539
rect 1286 1536 1287 1540
rect 1291 1536 1292 1540
rect 1286 1535 1292 1536
rect 1326 1536 1332 1537
rect 2502 1536 2508 1537
rect 1238 1534 1244 1535
rect 264 1507 266 1534
rect 336 1507 338 1534
rect 416 1507 418 1534
rect 504 1507 506 1534
rect 600 1507 602 1534
rect 688 1507 690 1534
rect 776 1507 778 1534
rect 864 1507 866 1534
rect 944 1507 946 1534
rect 1024 1507 1026 1534
rect 1104 1507 1106 1534
rect 1184 1507 1186 1534
rect 1240 1507 1242 1534
rect 1288 1507 1290 1535
rect 1326 1532 1327 1536
rect 1331 1532 1332 1536
rect 1326 1531 1332 1532
rect 1366 1535 1372 1536
rect 1366 1531 1367 1535
rect 1371 1531 1372 1535
rect 1328 1511 1330 1531
rect 1366 1530 1372 1531
rect 1486 1535 1492 1536
rect 1486 1531 1487 1535
rect 1491 1531 1492 1535
rect 1486 1530 1492 1531
rect 1622 1535 1628 1536
rect 1622 1531 1623 1535
rect 1627 1531 1628 1535
rect 1622 1530 1628 1531
rect 1750 1535 1756 1536
rect 1750 1531 1751 1535
rect 1755 1531 1756 1535
rect 1750 1530 1756 1531
rect 1886 1535 1892 1536
rect 1886 1531 1887 1535
rect 1891 1531 1892 1535
rect 1886 1530 1892 1531
rect 2022 1535 2028 1536
rect 2022 1531 2023 1535
rect 2027 1531 2028 1535
rect 2502 1532 2503 1536
rect 2507 1532 2508 1536
rect 2502 1531 2508 1532
rect 2022 1530 2028 1531
rect 1368 1511 1370 1530
rect 1488 1511 1490 1530
rect 1624 1511 1626 1530
rect 1752 1511 1754 1530
rect 1888 1511 1890 1530
rect 2024 1511 2026 1530
rect 2504 1511 2506 1531
rect 1327 1510 1331 1511
rect 111 1506 115 1507
rect 111 1501 115 1502
rect 263 1506 267 1507
rect 263 1501 267 1502
rect 279 1506 283 1507
rect 279 1501 283 1502
rect 335 1506 339 1507
rect 335 1501 339 1502
rect 343 1506 347 1507
rect 343 1501 347 1502
rect 415 1506 419 1507
rect 415 1501 419 1502
rect 495 1506 499 1507
rect 495 1501 499 1502
rect 503 1506 507 1507
rect 503 1501 507 1502
rect 575 1506 579 1507
rect 575 1501 579 1502
rect 599 1506 603 1507
rect 599 1501 603 1502
rect 655 1506 659 1507
rect 655 1501 659 1502
rect 687 1506 691 1507
rect 687 1501 691 1502
rect 735 1506 739 1507
rect 735 1501 739 1502
rect 775 1506 779 1507
rect 775 1501 779 1502
rect 815 1506 819 1507
rect 815 1501 819 1502
rect 863 1506 867 1507
rect 863 1501 867 1502
rect 895 1506 899 1507
rect 895 1501 899 1502
rect 943 1506 947 1507
rect 943 1501 947 1502
rect 975 1506 979 1507
rect 975 1501 979 1502
rect 1023 1506 1027 1507
rect 1023 1501 1027 1502
rect 1055 1506 1059 1507
rect 1055 1501 1059 1502
rect 1103 1506 1107 1507
rect 1103 1501 1107 1502
rect 1143 1506 1147 1507
rect 1143 1501 1147 1502
rect 1183 1506 1187 1507
rect 1183 1501 1187 1502
rect 1239 1506 1243 1507
rect 1239 1501 1243 1502
rect 1287 1506 1291 1507
rect 1327 1505 1331 1506
rect 1367 1510 1371 1511
rect 1367 1505 1371 1506
rect 1423 1510 1427 1511
rect 1423 1505 1427 1506
rect 1479 1510 1483 1511
rect 1479 1505 1483 1506
rect 1487 1510 1491 1511
rect 1487 1505 1491 1506
rect 1551 1510 1555 1511
rect 1551 1505 1555 1506
rect 1623 1510 1627 1511
rect 1623 1505 1627 1506
rect 1631 1510 1635 1511
rect 1631 1505 1635 1506
rect 1711 1510 1715 1511
rect 1711 1505 1715 1506
rect 1751 1510 1755 1511
rect 1751 1505 1755 1506
rect 1791 1510 1795 1511
rect 1791 1505 1795 1506
rect 1871 1510 1875 1511
rect 1871 1505 1875 1506
rect 1887 1510 1891 1511
rect 1887 1505 1891 1506
rect 1951 1510 1955 1511
rect 1951 1505 1955 1506
rect 2023 1510 2027 1511
rect 2023 1505 2027 1506
rect 2031 1510 2035 1511
rect 2031 1505 2035 1506
rect 2119 1510 2123 1511
rect 2119 1505 2123 1506
rect 2503 1510 2507 1511
rect 2503 1505 2507 1506
rect 1287 1501 1291 1502
rect 112 1481 114 1501
rect 280 1482 282 1501
rect 344 1482 346 1501
rect 416 1482 418 1501
rect 496 1482 498 1501
rect 576 1482 578 1501
rect 656 1482 658 1501
rect 736 1482 738 1501
rect 816 1482 818 1501
rect 896 1482 898 1501
rect 976 1482 978 1501
rect 1056 1482 1058 1501
rect 1144 1482 1146 1501
rect 278 1481 284 1482
rect 110 1480 116 1481
rect 110 1476 111 1480
rect 115 1476 116 1480
rect 278 1477 279 1481
rect 283 1477 284 1481
rect 278 1476 284 1477
rect 342 1481 348 1482
rect 342 1477 343 1481
rect 347 1477 348 1481
rect 342 1476 348 1477
rect 414 1481 420 1482
rect 414 1477 415 1481
rect 419 1477 420 1481
rect 414 1476 420 1477
rect 494 1481 500 1482
rect 494 1477 495 1481
rect 499 1477 500 1481
rect 494 1476 500 1477
rect 574 1481 580 1482
rect 574 1477 575 1481
rect 579 1477 580 1481
rect 574 1476 580 1477
rect 654 1481 660 1482
rect 654 1477 655 1481
rect 659 1477 660 1481
rect 654 1476 660 1477
rect 734 1481 740 1482
rect 734 1477 735 1481
rect 739 1477 740 1481
rect 734 1476 740 1477
rect 814 1481 820 1482
rect 814 1477 815 1481
rect 819 1477 820 1481
rect 814 1476 820 1477
rect 894 1481 900 1482
rect 894 1477 895 1481
rect 899 1477 900 1481
rect 894 1476 900 1477
rect 974 1481 980 1482
rect 974 1477 975 1481
rect 979 1477 980 1481
rect 974 1476 980 1477
rect 1054 1481 1060 1482
rect 1054 1477 1055 1481
rect 1059 1477 1060 1481
rect 1054 1476 1060 1477
rect 1142 1481 1148 1482
rect 1288 1481 1290 1501
rect 1328 1485 1330 1505
rect 1368 1486 1370 1505
rect 1424 1486 1426 1505
rect 1480 1486 1482 1505
rect 1552 1486 1554 1505
rect 1632 1486 1634 1505
rect 1712 1486 1714 1505
rect 1792 1486 1794 1505
rect 1872 1486 1874 1505
rect 1952 1486 1954 1505
rect 2032 1486 2034 1505
rect 2120 1486 2122 1505
rect 1366 1485 1372 1486
rect 1326 1484 1332 1485
rect 1142 1477 1143 1481
rect 1147 1477 1148 1481
rect 1142 1476 1148 1477
rect 1286 1480 1292 1481
rect 1286 1476 1287 1480
rect 1291 1476 1292 1480
rect 1326 1480 1327 1484
rect 1331 1480 1332 1484
rect 1366 1481 1367 1485
rect 1371 1481 1372 1485
rect 1366 1480 1372 1481
rect 1422 1485 1428 1486
rect 1422 1481 1423 1485
rect 1427 1481 1428 1485
rect 1422 1480 1428 1481
rect 1478 1485 1484 1486
rect 1478 1481 1479 1485
rect 1483 1481 1484 1485
rect 1478 1480 1484 1481
rect 1550 1485 1556 1486
rect 1550 1481 1551 1485
rect 1555 1481 1556 1485
rect 1550 1480 1556 1481
rect 1630 1485 1636 1486
rect 1630 1481 1631 1485
rect 1635 1481 1636 1485
rect 1630 1480 1636 1481
rect 1710 1485 1716 1486
rect 1710 1481 1711 1485
rect 1715 1481 1716 1485
rect 1710 1480 1716 1481
rect 1790 1485 1796 1486
rect 1790 1481 1791 1485
rect 1795 1481 1796 1485
rect 1790 1480 1796 1481
rect 1870 1485 1876 1486
rect 1870 1481 1871 1485
rect 1875 1481 1876 1485
rect 1870 1480 1876 1481
rect 1950 1485 1956 1486
rect 1950 1481 1951 1485
rect 1955 1481 1956 1485
rect 1950 1480 1956 1481
rect 2030 1485 2036 1486
rect 2030 1481 2031 1485
rect 2035 1481 2036 1485
rect 2030 1480 2036 1481
rect 2118 1485 2124 1486
rect 2504 1485 2506 1505
rect 2118 1481 2119 1485
rect 2123 1481 2124 1485
rect 2118 1480 2124 1481
rect 2502 1484 2508 1485
rect 2502 1480 2503 1484
rect 2507 1480 2508 1484
rect 1326 1479 1332 1480
rect 2502 1479 2508 1480
rect 110 1475 116 1476
rect 1286 1475 1292 1476
rect 1326 1467 1332 1468
rect 110 1463 116 1464
rect 110 1459 111 1463
rect 115 1459 116 1463
rect 1286 1463 1292 1464
rect 110 1458 116 1459
rect 262 1460 268 1461
rect 112 1451 114 1458
rect 262 1456 263 1460
rect 267 1456 268 1460
rect 262 1455 268 1456
rect 326 1460 332 1461
rect 326 1456 327 1460
rect 331 1456 332 1460
rect 326 1455 332 1456
rect 398 1460 404 1461
rect 398 1456 399 1460
rect 403 1456 404 1460
rect 398 1455 404 1456
rect 478 1460 484 1461
rect 478 1456 479 1460
rect 483 1456 484 1460
rect 478 1455 484 1456
rect 558 1460 564 1461
rect 558 1456 559 1460
rect 563 1456 564 1460
rect 558 1455 564 1456
rect 638 1460 644 1461
rect 638 1456 639 1460
rect 643 1456 644 1460
rect 638 1455 644 1456
rect 718 1460 724 1461
rect 718 1456 719 1460
rect 723 1456 724 1460
rect 718 1455 724 1456
rect 798 1460 804 1461
rect 798 1456 799 1460
rect 803 1456 804 1460
rect 798 1455 804 1456
rect 878 1460 884 1461
rect 878 1456 879 1460
rect 883 1456 884 1460
rect 878 1455 884 1456
rect 958 1460 964 1461
rect 958 1456 959 1460
rect 963 1456 964 1460
rect 958 1455 964 1456
rect 1038 1460 1044 1461
rect 1038 1456 1039 1460
rect 1043 1456 1044 1460
rect 1038 1455 1044 1456
rect 1126 1460 1132 1461
rect 1126 1456 1127 1460
rect 1131 1456 1132 1460
rect 1286 1459 1287 1463
rect 1291 1459 1292 1463
rect 1326 1463 1327 1467
rect 1331 1463 1332 1467
rect 2502 1467 2508 1468
rect 1326 1462 1332 1463
rect 1350 1464 1356 1465
rect 1286 1458 1292 1459
rect 1126 1455 1132 1456
rect 264 1451 266 1455
rect 328 1451 330 1455
rect 400 1451 402 1455
rect 480 1451 482 1455
rect 560 1451 562 1455
rect 640 1451 642 1455
rect 720 1451 722 1455
rect 800 1451 802 1455
rect 880 1451 882 1455
rect 960 1451 962 1455
rect 1040 1451 1042 1455
rect 1128 1451 1130 1455
rect 1288 1451 1290 1458
rect 1328 1451 1330 1462
rect 1350 1460 1351 1464
rect 1355 1460 1356 1464
rect 1350 1459 1356 1460
rect 1406 1464 1412 1465
rect 1406 1460 1407 1464
rect 1411 1460 1412 1464
rect 1406 1459 1412 1460
rect 1462 1464 1468 1465
rect 1462 1460 1463 1464
rect 1467 1460 1468 1464
rect 1462 1459 1468 1460
rect 1534 1464 1540 1465
rect 1534 1460 1535 1464
rect 1539 1460 1540 1464
rect 1534 1459 1540 1460
rect 1614 1464 1620 1465
rect 1614 1460 1615 1464
rect 1619 1460 1620 1464
rect 1614 1459 1620 1460
rect 1694 1464 1700 1465
rect 1694 1460 1695 1464
rect 1699 1460 1700 1464
rect 1694 1459 1700 1460
rect 1774 1464 1780 1465
rect 1774 1460 1775 1464
rect 1779 1460 1780 1464
rect 1774 1459 1780 1460
rect 1854 1464 1860 1465
rect 1854 1460 1855 1464
rect 1859 1460 1860 1464
rect 1854 1459 1860 1460
rect 1934 1464 1940 1465
rect 1934 1460 1935 1464
rect 1939 1460 1940 1464
rect 1934 1459 1940 1460
rect 2014 1464 2020 1465
rect 2014 1460 2015 1464
rect 2019 1460 2020 1464
rect 2014 1459 2020 1460
rect 2102 1464 2108 1465
rect 2102 1460 2103 1464
rect 2107 1460 2108 1464
rect 2502 1463 2503 1467
rect 2507 1463 2508 1467
rect 2502 1462 2508 1463
rect 2102 1459 2108 1460
rect 1352 1451 1354 1459
rect 1408 1451 1410 1459
rect 1464 1451 1466 1459
rect 1536 1451 1538 1459
rect 1616 1451 1618 1459
rect 1696 1451 1698 1459
rect 1776 1451 1778 1459
rect 1856 1451 1858 1459
rect 1936 1451 1938 1459
rect 2016 1451 2018 1459
rect 2104 1451 2106 1459
rect 2504 1451 2506 1462
rect 111 1450 115 1451
rect 111 1445 115 1446
rect 191 1450 195 1451
rect 191 1445 195 1446
rect 255 1450 259 1451
rect 255 1445 259 1446
rect 263 1450 267 1451
rect 263 1445 267 1446
rect 327 1450 331 1451
rect 327 1445 331 1446
rect 399 1450 403 1451
rect 399 1445 403 1446
rect 407 1450 411 1451
rect 407 1445 411 1446
rect 479 1450 483 1451
rect 479 1445 483 1446
rect 503 1450 507 1451
rect 503 1445 507 1446
rect 559 1450 563 1451
rect 559 1445 563 1446
rect 607 1450 611 1451
rect 607 1445 611 1446
rect 639 1450 643 1451
rect 639 1445 643 1446
rect 711 1450 715 1451
rect 711 1445 715 1446
rect 719 1450 723 1451
rect 719 1445 723 1446
rect 799 1450 803 1451
rect 799 1445 803 1446
rect 815 1450 819 1451
rect 815 1445 819 1446
rect 879 1450 883 1451
rect 879 1445 883 1446
rect 919 1450 923 1451
rect 919 1445 923 1446
rect 959 1450 963 1451
rect 959 1445 963 1446
rect 1023 1450 1027 1451
rect 1023 1445 1027 1446
rect 1039 1450 1043 1451
rect 1039 1445 1043 1446
rect 1127 1450 1131 1451
rect 1127 1445 1131 1446
rect 1223 1450 1227 1451
rect 1223 1445 1227 1446
rect 1287 1450 1291 1451
rect 1287 1445 1291 1446
rect 1327 1450 1331 1451
rect 1327 1445 1331 1446
rect 1351 1450 1355 1451
rect 1351 1445 1355 1446
rect 1359 1450 1363 1451
rect 1359 1445 1363 1446
rect 1407 1450 1411 1451
rect 1407 1445 1411 1446
rect 1447 1450 1451 1451
rect 1447 1445 1451 1446
rect 1463 1450 1467 1451
rect 1463 1445 1467 1446
rect 1535 1450 1539 1451
rect 1535 1445 1539 1446
rect 1615 1450 1619 1451
rect 1615 1445 1619 1446
rect 1631 1450 1635 1451
rect 1631 1445 1635 1446
rect 1695 1450 1699 1451
rect 1695 1445 1699 1446
rect 1727 1450 1731 1451
rect 1727 1445 1731 1446
rect 1775 1450 1779 1451
rect 1775 1445 1779 1446
rect 1815 1450 1819 1451
rect 1815 1445 1819 1446
rect 1855 1450 1859 1451
rect 1855 1445 1859 1446
rect 1903 1450 1907 1451
rect 1903 1445 1907 1446
rect 1935 1450 1939 1451
rect 1935 1445 1939 1446
rect 1991 1450 1995 1451
rect 1991 1445 1995 1446
rect 2015 1450 2019 1451
rect 2015 1445 2019 1446
rect 2071 1450 2075 1451
rect 2071 1445 2075 1446
rect 2103 1450 2107 1451
rect 2103 1445 2107 1446
rect 2159 1450 2163 1451
rect 2159 1445 2163 1446
rect 2247 1450 2251 1451
rect 2247 1445 2251 1446
rect 2503 1450 2507 1451
rect 2503 1445 2507 1446
rect 112 1442 114 1445
rect 190 1444 196 1445
rect 110 1441 116 1442
rect 110 1437 111 1441
rect 115 1437 116 1441
rect 190 1440 191 1444
rect 195 1440 196 1444
rect 190 1439 196 1440
rect 254 1444 260 1445
rect 254 1440 255 1444
rect 259 1440 260 1444
rect 254 1439 260 1440
rect 326 1444 332 1445
rect 326 1440 327 1444
rect 331 1440 332 1444
rect 326 1439 332 1440
rect 406 1444 412 1445
rect 406 1440 407 1444
rect 411 1440 412 1444
rect 406 1439 412 1440
rect 502 1444 508 1445
rect 502 1440 503 1444
rect 507 1440 508 1444
rect 502 1439 508 1440
rect 606 1444 612 1445
rect 606 1440 607 1444
rect 611 1440 612 1444
rect 606 1439 612 1440
rect 710 1444 716 1445
rect 710 1440 711 1444
rect 715 1440 716 1444
rect 710 1439 716 1440
rect 814 1444 820 1445
rect 814 1440 815 1444
rect 819 1440 820 1444
rect 814 1439 820 1440
rect 918 1444 924 1445
rect 918 1440 919 1444
rect 923 1440 924 1444
rect 918 1439 924 1440
rect 1022 1444 1028 1445
rect 1022 1440 1023 1444
rect 1027 1440 1028 1444
rect 1022 1439 1028 1440
rect 1126 1444 1132 1445
rect 1126 1440 1127 1444
rect 1131 1440 1132 1444
rect 1126 1439 1132 1440
rect 1222 1444 1228 1445
rect 1222 1440 1223 1444
rect 1227 1440 1228 1444
rect 1288 1442 1290 1445
rect 1328 1442 1330 1445
rect 1358 1444 1364 1445
rect 1222 1439 1228 1440
rect 1286 1441 1292 1442
rect 110 1436 116 1437
rect 1286 1437 1287 1441
rect 1291 1437 1292 1441
rect 1286 1436 1292 1437
rect 1326 1441 1332 1442
rect 1326 1437 1327 1441
rect 1331 1437 1332 1441
rect 1358 1440 1359 1444
rect 1363 1440 1364 1444
rect 1358 1439 1364 1440
rect 1446 1444 1452 1445
rect 1446 1440 1447 1444
rect 1451 1440 1452 1444
rect 1446 1439 1452 1440
rect 1534 1444 1540 1445
rect 1534 1440 1535 1444
rect 1539 1440 1540 1444
rect 1534 1439 1540 1440
rect 1630 1444 1636 1445
rect 1630 1440 1631 1444
rect 1635 1440 1636 1444
rect 1630 1439 1636 1440
rect 1726 1444 1732 1445
rect 1726 1440 1727 1444
rect 1731 1440 1732 1444
rect 1726 1439 1732 1440
rect 1814 1444 1820 1445
rect 1814 1440 1815 1444
rect 1819 1440 1820 1444
rect 1814 1439 1820 1440
rect 1902 1444 1908 1445
rect 1902 1440 1903 1444
rect 1907 1440 1908 1444
rect 1902 1439 1908 1440
rect 1990 1444 1996 1445
rect 1990 1440 1991 1444
rect 1995 1440 1996 1444
rect 1990 1439 1996 1440
rect 2070 1444 2076 1445
rect 2070 1440 2071 1444
rect 2075 1440 2076 1444
rect 2070 1439 2076 1440
rect 2158 1444 2164 1445
rect 2158 1440 2159 1444
rect 2163 1440 2164 1444
rect 2158 1439 2164 1440
rect 2246 1444 2252 1445
rect 2246 1440 2247 1444
rect 2251 1440 2252 1444
rect 2504 1442 2506 1445
rect 2246 1439 2252 1440
rect 2502 1441 2508 1442
rect 1326 1436 1332 1437
rect 2502 1437 2503 1441
rect 2507 1437 2508 1441
rect 2502 1436 2508 1437
rect 110 1424 116 1425
rect 1286 1424 1292 1425
rect 110 1420 111 1424
rect 115 1420 116 1424
rect 110 1419 116 1420
rect 206 1423 212 1424
rect 206 1419 207 1423
rect 211 1419 212 1423
rect 112 1395 114 1419
rect 206 1418 212 1419
rect 270 1423 276 1424
rect 270 1419 271 1423
rect 275 1419 276 1423
rect 270 1418 276 1419
rect 342 1423 348 1424
rect 342 1419 343 1423
rect 347 1419 348 1423
rect 342 1418 348 1419
rect 422 1423 428 1424
rect 422 1419 423 1423
rect 427 1419 428 1423
rect 422 1418 428 1419
rect 518 1423 524 1424
rect 518 1419 519 1423
rect 523 1419 524 1423
rect 518 1418 524 1419
rect 622 1423 628 1424
rect 622 1419 623 1423
rect 627 1419 628 1423
rect 622 1418 628 1419
rect 726 1423 732 1424
rect 726 1419 727 1423
rect 731 1419 732 1423
rect 726 1418 732 1419
rect 830 1423 836 1424
rect 830 1419 831 1423
rect 835 1419 836 1423
rect 830 1418 836 1419
rect 934 1423 940 1424
rect 934 1419 935 1423
rect 939 1419 940 1423
rect 934 1418 940 1419
rect 1038 1423 1044 1424
rect 1038 1419 1039 1423
rect 1043 1419 1044 1423
rect 1038 1418 1044 1419
rect 1142 1423 1148 1424
rect 1142 1419 1143 1423
rect 1147 1419 1148 1423
rect 1142 1418 1148 1419
rect 1238 1423 1244 1424
rect 1238 1419 1239 1423
rect 1243 1419 1244 1423
rect 1286 1420 1287 1424
rect 1291 1420 1292 1424
rect 1286 1419 1292 1420
rect 1326 1424 1332 1425
rect 2502 1424 2508 1425
rect 1326 1420 1327 1424
rect 1331 1420 1332 1424
rect 1326 1419 1332 1420
rect 1374 1423 1380 1424
rect 1374 1419 1375 1423
rect 1379 1419 1380 1423
rect 1238 1418 1244 1419
rect 208 1395 210 1418
rect 272 1395 274 1418
rect 344 1395 346 1418
rect 424 1395 426 1418
rect 520 1395 522 1418
rect 624 1395 626 1418
rect 728 1395 730 1418
rect 832 1395 834 1418
rect 936 1395 938 1418
rect 1040 1395 1042 1418
rect 1144 1395 1146 1418
rect 1240 1395 1242 1418
rect 1288 1395 1290 1419
rect 1328 1399 1330 1419
rect 1374 1418 1380 1419
rect 1462 1423 1468 1424
rect 1462 1419 1463 1423
rect 1467 1419 1468 1423
rect 1462 1418 1468 1419
rect 1550 1423 1556 1424
rect 1550 1419 1551 1423
rect 1555 1419 1556 1423
rect 1550 1418 1556 1419
rect 1646 1423 1652 1424
rect 1646 1419 1647 1423
rect 1651 1419 1652 1423
rect 1646 1418 1652 1419
rect 1742 1423 1748 1424
rect 1742 1419 1743 1423
rect 1747 1419 1748 1423
rect 1742 1418 1748 1419
rect 1830 1423 1836 1424
rect 1830 1419 1831 1423
rect 1835 1419 1836 1423
rect 1830 1418 1836 1419
rect 1918 1423 1924 1424
rect 1918 1419 1919 1423
rect 1923 1419 1924 1423
rect 1918 1418 1924 1419
rect 2006 1423 2012 1424
rect 2006 1419 2007 1423
rect 2011 1419 2012 1423
rect 2006 1418 2012 1419
rect 2086 1423 2092 1424
rect 2086 1419 2087 1423
rect 2091 1419 2092 1423
rect 2086 1418 2092 1419
rect 2174 1423 2180 1424
rect 2174 1419 2175 1423
rect 2179 1419 2180 1423
rect 2174 1418 2180 1419
rect 2262 1423 2268 1424
rect 2262 1419 2263 1423
rect 2267 1419 2268 1423
rect 2502 1420 2503 1424
rect 2507 1420 2508 1424
rect 2502 1419 2508 1420
rect 2262 1418 2268 1419
rect 1376 1399 1378 1418
rect 1464 1399 1466 1418
rect 1552 1399 1554 1418
rect 1648 1399 1650 1418
rect 1744 1399 1746 1418
rect 1832 1399 1834 1418
rect 1920 1399 1922 1418
rect 2008 1399 2010 1418
rect 2088 1399 2090 1418
rect 2176 1399 2178 1418
rect 2264 1399 2266 1418
rect 2504 1399 2506 1419
rect 1327 1398 1331 1399
rect 111 1394 115 1395
rect 111 1389 115 1390
rect 151 1394 155 1395
rect 151 1389 155 1390
rect 207 1394 211 1395
rect 207 1389 211 1390
rect 223 1394 227 1395
rect 223 1389 227 1390
rect 271 1394 275 1395
rect 271 1389 275 1390
rect 295 1394 299 1395
rect 295 1389 299 1390
rect 343 1394 347 1395
rect 343 1389 347 1390
rect 359 1394 363 1395
rect 359 1389 363 1390
rect 423 1394 427 1395
rect 423 1389 427 1390
rect 431 1394 435 1395
rect 431 1389 435 1390
rect 503 1394 507 1395
rect 503 1389 507 1390
rect 519 1394 523 1395
rect 519 1389 523 1390
rect 583 1394 587 1395
rect 583 1389 587 1390
rect 623 1394 627 1395
rect 623 1389 627 1390
rect 663 1394 667 1395
rect 663 1389 667 1390
rect 727 1394 731 1395
rect 727 1389 731 1390
rect 751 1394 755 1395
rect 751 1389 755 1390
rect 831 1394 835 1395
rect 831 1389 835 1390
rect 839 1394 843 1395
rect 839 1389 843 1390
rect 927 1394 931 1395
rect 927 1389 931 1390
rect 935 1394 939 1395
rect 935 1389 939 1390
rect 1015 1394 1019 1395
rect 1015 1389 1019 1390
rect 1039 1394 1043 1395
rect 1039 1389 1043 1390
rect 1103 1394 1107 1395
rect 1103 1389 1107 1390
rect 1143 1394 1147 1395
rect 1143 1389 1147 1390
rect 1199 1394 1203 1395
rect 1199 1389 1203 1390
rect 1239 1394 1243 1395
rect 1239 1389 1243 1390
rect 1287 1394 1291 1395
rect 1327 1393 1331 1394
rect 1375 1398 1379 1399
rect 1375 1393 1379 1394
rect 1463 1398 1467 1399
rect 1463 1393 1467 1394
rect 1551 1398 1555 1399
rect 1551 1393 1555 1394
rect 1567 1398 1571 1399
rect 1567 1393 1571 1394
rect 1647 1398 1651 1399
rect 1647 1393 1651 1394
rect 1735 1398 1739 1399
rect 1735 1393 1739 1394
rect 1743 1398 1747 1399
rect 1743 1393 1747 1394
rect 1831 1398 1835 1399
rect 1831 1393 1835 1394
rect 1919 1398 1923 1399
rect 1919 1393 1923 1394
rect 2007 1398 2011 1399
rect 2007 1393 2011 1394
rect 2087 1398 2091 1399
rect 2087 1393 2091 1394
rect 2095 1398 2099 1399
rect 2095 1393 2099 1394
rect 2175 1398 2179 1399
rect 2175 1393 2179 1394
rect 2247 1398 2251 1399
rect 2247 1393 2251 1394
rect 2263 1398 2267 1399
rect 2263 1393 2267 1394
rect 2319 1398 2323 1399
rect 2319 1393 2323 1394
rect 2399 1398 2403 1399
rect 2399 1393 2403 1394
rect 2455 1398 2459 1399
rect 2455 1393 2459 1394
rect 2503 1398 2507 1399
rect 2503 1393 2507 1394
rect 1287 1389 1291 1390
rect 112 1369 114 1389
rect 152 1370 154 1389
rect 224 1370 226 1389
rect 296 1370 298 1389
rect 360 1370 362 1389
rect 432 1370 434 1389
rect 504 1370 506 1389
rect 584 1370 586 1389
rect 664 1370 666 1389
rect 752 1370 754 1389
rect 840 1370 842 1389
rect 928 1370 930 1389
rect 1016 1370 1018 1389
rect 1104 1370 1106 1389
rect 1200 1370 1202 1389
rect 150 1369 156 1370
rect 110 1368 116 1369
rect 110 1364 111 1368
rect 115 1364 116 1368
rect 150 1365 151 1369
rect 155 1365 156 1369
rect 150 1364 156 1365
rect 222 1369 228 1370
rect 222 1365 223 1369
rect 227 1365 228 1369
rect 222 1364 228 1365
rect 294 1369 300 1370
rect 294 1365 295 1369
rect 299 1365 300 1369
rect 294 1364 300 1365
rect 358 1369 364 1370
rect 358 1365 359 1369
rect 363 1365 364 1369
rect 358 1364 364 1365
rect 430 1369 436 1370
rect 430 1365 431 1369
rect 435 1365 436 1369
rect 430 1364 436 1365
rect 502 1369 508 1370
rect 502 1365 503 1369
rect 507 1365 508 1369
rect 502 1364 508 1365
rect 582 1369 588 1370
rect 582 1365 583 1369
rect 587 1365 588 1369
rect 582 1364 588 1365
rect 662 1369 668 1370
rect 662 1365 663 1369
rect 667 1365 668 1369
rect 662 1364 668 1365
rect 750 1369 756 1370
rect 750 1365 751 1369
rect 755 1365 756 1369
rect 750 1364 756 1365
rect 838 1369 844 1370
rect 838 1365 839 1369
rect 843 1365 844 1369
rect 838 1364 844 1365
rect 926 1369 932 1370
rect 926 1365 927 1369
rect 931 1365 932 1369
rect 926 1364 932 1365
rect 1014 1369 1020 1370
rect 1014 1365 1015 1369
rect 1019 1365 1020 1369
rect 1014 1364 1020 1365
rect 1102 1369 1108 1370
rect 1102 1365 1103 1369
rect 1107 1365 1108 1369
rect 1102 1364 1108 1365
rect 1198 1369 1204 1370
rect 1288 1369 1290 1389
rect 1328 1373 1330 1393
rect 1568 1374 1570 1393
rect 1648 1374 1650 1393
rect 1736 1374 1738 1393
rect 1832 1374 1834 1393
rect 1920 1374 1922 1393
rect 2008 1374 2010 1393
rect 2096 1374 2098 1393
rect 2176 1374 2178 1393
rect 2248 1374 2250 1393
rect 2320 1374 2322 1393
rect 2400 1374 2402 1393
rect 2456 1374 2458 1393
rect 1566 1373 1572 1374
rect 1326 1372 1332 1373
rect 1198 1365 1199 1369
rect 1203 1365 1204 1369
rect 1198 1364 1204 1365
rect 1286 1368 1292 1369
rect 1286 1364 1287 1368
rect 1291 1364 1292 1368
rect 1326 1368 1327 1372
rect 1331 1368 1332 1372
rect 1566 1369 1567 1373
rect 1571 1369 1572 1373
rect 1566 1368 1572 1369
rect 1646 1373 1652 1374
rect 1646 1369 1647 1373
rect 1651 1369 1652 1373
rect 1646 1368 1652 1369
rect 1734 1373 1740 1374
rect 1734 1369 1735 1373
rect 1739 1369 1740 1373
rect 1734 1368 1740 1369
rect 1830 1373 1836 1374
rect 1830 1369 1831 1373
rect 1835 1369 1836 1373
rect 1830 1368 1836 1369
rect 1918 1373 1924 1374
rect 1918 1369 1919 1373
rect 1923 1369 1924 1373
rect 1918 1368 1924 1369
rect 2006 1373 2012 1374
rect 2006 1369 2007 1373
rect 2011 1369 2012 1373
rect 2006 1368 2012 1369
rect 2094 1373 2100 1374
rect 2094 1369 2095 1373
rect 2099 1369 2100 1373
rect 2094 1368 2100 1369
rect 2174 1373 2180 1374
rect 2174 1369 2175 1373
rect 2179 1369 2180 1373
rect 2174 1368 2180 1369
rect 2246 1373 2252 1374
rect 2246 1369 2247 1373
rect 2251 1369 2252 1373
rect 2246 1368 2252 1369
rect 2318 1373 2324 1374
rect 2318 1369 2319 1373
rect 2323 1369 2324 1373
rect 2318 1368 2324 1369
rect 2398 1373 2404 1374
rect 2398 1369 2399 1373
rect 2403 1369 2404 1373
rect 2398 1368 2404 1369
rect 2454 1373 2460 1374
rect 2504 1373 2506 1393
rect 2454 1369 2455 1373
rect 2459 1369 2460 1373
rect 2454 1368 2460 1369
rect 2502 1372 2508 1373
rect 2502 1368 2503 1372
rect 2507 1368 2508 1372
rect 1326 1367 1332 1368
rect 2502 1367 2508 1368
rect 110 1363 116 1364
rect 1286 1363 1292 1364
rect 1326 1355 1332 1356
rect 110 1351 116 1352
rect 110 1347 111 1351
rect 115 1347 116 1351
rect 1286 1351 1292 1352
rect 110 1346 116 1347
rect 134 1348 140 1349
rect 112 1327 114 1346
rect 134 1344 135 1348
rect 139 1344 140 1348
rect 134 1343 140 1344
rect 206 1348 212 1349
rect 206 1344 207 1348
rect 211 1344 212 1348
rect 206 1343 212 1344
rect 278 1348 284 1349
rect 278 1344 279 1348
rect 283 1344 284 1348
rect 278 1343 284 1344
rect 342 1348 348 1349
rect 342 1344 343 1348
rect 347 1344 348 1348
rect 342 1343 348 1344
rect 414 1348 420 1349
rect 414 1344 415 1348
rect 419 1344 420 1348
rect 414 1343 420 1344
rect 486 1348 492 1349
rect 486 1344 487 1348
rect 491 1344 492 1348
rect 486 1343 492 1344
rect 566 1348 572 1349
rect 566 1344 567 1348
rect 571 1344 572 1348
rect 566 1343 572 1344
rect 646 1348 652 1349
rect 646 1344 647 1348
rect 651 1344 652 1348
rect 646 1343 652 1344
rect 734 1348 740 1349
rect 734 1344 735 1348
rect 739 1344 740 1348
rect 734 1343 740 1344
rect 822 1348 828 1349
rect 822 1344 823 1348
rect 827 1344 828 1348
rect 822 1343 828 1344
rect 910 1348 916 1349
rect 910 1344 911 1348
rect 915 1344 916 1348
rect 910 1343 916 1344
rect 998 1348 1004 1349
rect 998 1344 999 1348
rect 1003 1344 1004 1348
rect 998 1343 1004 1344
rect 1086 1348 1092 1349
rect 1086 1344 1087 1348
rect 1091 1344 1092 1348
rect 1086 1343 1092 1344
rect 1182 1348 1188 1349
rect 1182 1344 1183 1348
rect 1187 1344 1188 1348
rect 1286 1347 1287 1351
rect 1291 1347 1292 1351
rect 1326 1351 1327 1355
rect 1331 1351 1332 1355
rect 2502 1355 2508 1356
rect 1326 1350 1332 1351
rect 1550 1352 1556 1353
rect 1328 1347 1330 1350
rect 1550 1348 1551 1352
rect 1555 1348 1556 1352
rect 1550 1347 1556 1348
rect 1630 1352 1636 1353
rect 1630 1348 1631 1352
rect 1635 1348 1636 1352
rect 1630 1347 1636 1348
rect 1718 1352 1724 1353
rect 1718 1348 1719 1352
rect 1723 1348 1724 1352
rect 1718 1347 1724 1348
rect 1814 1352 1820 1353
rect 1814 1348 1815 1352
rect 1819 1348 1820 1352
rect 1814 1347 1820 1348
rect 1902 1352 1908 1353
rect 1902 1348 1903 1352
rect 1907 1348 1908 1352
rect 1902 1347 1908 1348
rect 1990 1352 1996 1353
rect 1990 1348 1991 1352
rect 1995 1348 1996 1352
rect 1990 1347 1996 1348
rect 2078 1352 2084 1353
rect 2078 1348 2079 1352
rect 2083 1348 2084 1352
rect 2078 1347 2084 1348
rect 2158 1352 2164 1353
rect 2158 1348 2159 1352
rect 2163 1348 2164 1352
rect 2158 1347 2164 1348
rect 2230 1352 2236 1353
rect 2230 1348 2231 1352
rect 2235 1348 2236 1352
rect 2230 1347 2236 1348
rect 2302 1352 2308 1353
rect 2302 1348 2303 1352
rect 2307 1348 2308 1352
rect 2302 1347 2308 1348
rect 2382 1352 2388 1353
rect 2382 1348 2383 1352
rect 2387 1348 2388 1352
rect 2382 1347 2388 1348
rect 2438 1352 2444 1353
rect 2438 1348 2439 1352
rect 2443 1348 2444 1352
rect 2502 1351 2503 1355
rect 2507 1351 2508 1355
rect 2502 1350 2508 1351
rect 2438 1347 2444 1348
rect 2504 1347 2506 1350
rect 1286 1346 1292 1347
rect 1327 1346 1331 1347
rect 1182 1343 1188 1344
rect 136 1327 138 1343
rect 208 1327 210 1343
rect 280 1327 282 1343
rect 344 1327 346 1343
rect 416 1327 418 1343
rect 488 1327 490 1343
rect 568 1327 570 1343
rect 648 1327 650 1343
rect 736 1327 738 1343
rect 824 1327 826 1343
rect 912 1327 914 1343
rect 1000 1327 1002 1343
rect 1088 1327 1090 1343
rect 1184 1327 1186 1343
rect 1288 1327 1290 1346
rect 1327 1341 1331 1342
rect 1551 1346 1555 1347
rect 1551 1341 1555 1342
rect 1583 1346 1587 1347
rect 1583 1341 1587 1342
rect 1631 1346 1635 1347
rect 1631 1341 1635 1342
rect 1647 1346 1651 1347
rect 1647 1341 1651 1342
rect 1719 1346 1723 1347
rect 1719 1341 1723 1342
rect 1727 1346 1731 1347
rect 1727 1341 1731 1342
rect 1807 1346 1811 1347
rect 1807 1341 1811 1342
rect 1815 1346 1819 1347
rect 1815 1341 1819 1342
rect 1895 1346 1899 1347
rect 1895 1341 1899 1342
rect 1903 1346 1907 1347
rect 1903 1341 1907 1342
rect 1983 1346 1987 1347
rect 1983 1341 1987 1342
rect 1991 1346 1995 1347
rect 1991 1341 1995 1342
rect 2063 1346 2067 1347
rect 2063 1341 2067 1342
rect 2079 1346 2083 1347
rect 2079 1341 2083 1342
rect 2143 1346 2147 1347
rect 2143 1341 2147 1342
rect 2159 1346 2163 1347
rect 2159 1341 2163 1342
rect 2223 1346 2227 1347
rect 2223 1341 2227 1342
rect 2231 1346 2235 1347
rect 2231 1341 2235 1342
rect 2303 1346 2307 1347
rect 2303 1341 2307 1342
rect 2383 1346 2387 1347
rect 2383 1341 2387 1342
rect 2439 1346 2443 1347
rect 2439 1341 2443 1342
rect 2503 1346 2507 1347
rect 2503 1341 2507 1342
rect 1328 1338 1330 1341
rect 1582 1340 1588 1341
rect 1326 1337 1332 1338
rect 1326 1333 1327 1337
rect 1331 1333 1332 1337
rect 1582 1336 1583 1340
rect 1587 1336 1588 1340
rect 1582 1335 1588 1336
rect 1646 1340 1652 1341
rect 1646 1336 1647 1340
rect 1651 1336 1652 1340
rect 1646 1335 1652 1336
rect 1726 1340 1732 1341
rect 1726 1336 1727 1340
rect 1731 1336 1732 1340
rect 1726 1335 1732 1336
rect 1806 1340 1812 1341
rect 1806 1336 1807 1340
rect 1811 1336 1812 1340
rect 1806 1335 1812 1336
rect 1894 1340 1900 1341
rect 1894 1336 1895 1340
rect 1899 1336 1900 1340
rect 1894 1335 1900 1336
rect 1982 1340 1988 1341
rect 1982 1336 1983 1340
rect 1987 1336 1988 1340
rect 1982 1335 1988 1336
rect 2062 1340 2068 1341
rect 2062 1336 2063 1340
rect 2067 1336 2068 1340
rect 2062 1335 2068 1336
rect 2142 1340 2148 1341
rect 2142 1336 2143 1340
rect 2147 1336 2148 1340
rect 2142 1335 2148 1336
rect 2222 1340 2228 1341
rect 2222 1336 2223 1340
rect 2227 1336 2228 1340
rect 2222 1335 2228 1336
rect 2302 1340 2308 1341
rect 2302 1336 2303 1340
rect 2307 1336 2308 1340
rect 2302 1335 2308 1336
rect 2382 1340 2388 1341
rect 2382 1336 2383 1340
rect 2387 1336 2388 1340
rect 2382 1335 2388 1336
rect 2438 1340 2444 1341
rect 2438 1336 2439 1340
rect 2443 1336 2444 1340
rect 2504 1338 2506 1341
rect 2438 1335 2444 1336
rect 2502 1337 2508 1338
rect 1326 1332 1332 1333
rect 2502 1333 2503 1337
rect 2507 1333 2508 1337
rect 2502 1332 2508 1333
rect 111 1326 115 1327
rect 111 1321 115 1322
rect 135 1326 139 1327
rect 135 1321 139 1322
rect 207 1326 211 1327
rect 207 1321 211 1322
rect 239 1326 243 1327
rect 239 1321 243 1322
rect 279 1326 283 1327
rect 279 1321 283 1322
rect 343 1326 347 1327
rect 343 1321 347 1322
rect 367 1326 371 1327
rect 367 1321 371 1322
rect 415 1326 419 1327
rect 415 1321 419 1322
rect 479 1326 483 1327
rect 479 1321 483 1322
rect 487 1326 491 1327
rect 487 1321 491 1322
rect 567 1326 571 1327
rect 567 1321 571 1322
rect 583 1326 587 1327
rect 583 1321 587 1322
rect 647 1326 651 1327
rect 647 1321 651 1322
rect 687 1326 691 1327
rect 687 1321 691 1322
rect 735 1326 739 1327
rect 735 1321 739 1322
rect 783 1326 787 1327
rect 783 1321 787 1322
rect 823 1326 827 1327
rect 823 1321 827 1322
rect 879 1326 883 1327
rect 879 1321 883 1322
rect 911 1326 915 1327
rect 911 1321 915 1322
rect 975 1326 979 1327
rect 975 1321 979 1322
rect 999 1326 1003 1327
rect 999 1321 1003 1322
rect 1087 1326 1091 1327
rect 1087 1321 1091 1322
rect 1183 1326 1187 1327
rect 1183 1321 1187 1322
rect 1287 1326 1291 1327
rect 1287 1321 1291 1322
rect 112 1318 114 1321
rect 134 1320 140 1321
rect 110 1317 116 1318
rect 110 1313 111 1317
rect 115 1313 116 1317
rect 134 1316 135 1320
rect 139 1316 140 1320
rect 134 1315 140 1316
rect 238 1320 244 1321
rect 238 1316 239 1320
rect 243 1316 244 1320
rect 238 1315 244 1316
rect 366 1320 372 1321
rect 366 1316 367 1320
rect 371 1316 372 1320
rect 366 1315 372 1316
rect 478 1320 484 1321
rect 478 1316 479 1320
rect 483 1316 484 1320
rect 478 1315 484 1316
rect 582 1320 588 1321
rect 582 1316 583 1320
rect 587 1316 588 1320
rect 582 1315 588 1316
rect 686 1320 692 1321
rect 686 1316 687 1320
rect 691 1316 692 1320
rect 686 1315 692 1316
rect 782 1320 788 1321
rect 782 1316 783 1320
rect 787 1316 788 1320
rect 782 1315 788 1316
rect 878 1320 884 1321
rect 878 1316 879 1320
rect 883 1316 884 1320
rect 878 1315 884 1316
rect 974 1320 980 1321
rect 974 1316 975 1320
rect 979 1316 980 1320
rect 1288 1318 1290 1321
rect 1326 1320 1332 1321
rect 2502 1320 2508 1321
rect 974 1315 980 1316
rect 1286 1317 1292 1318
rect 110 1312 116 1313
rect 1286 1313 1287 1317
rect 1291 1313 1292 1317
rect 1326 1316 1327 1320
rect 1331 1316 1332 1320
rect 1326 1315 1332 1316
rect 1598 1319 1604 1320
rect 1598 1315 1599 1319
rect 1603 1315 1604 1319
rect 1286 1312 1292 1313
rect 110 1300 116 1301
rect 1286 1300 1292 1301
rect 110 1296 111 1300
rect 115 1296 116 1300
rect 110 1295 116 1296
rect 150 1299 156 1300
rect 150 1295 151 1299
rect 155 1295 156 1299
rect 112 1267 114 1295
rect 150 1294 156 1295
rect 254 1299 260 1300
rect 254 1295 255 1299
rect 259 1295 260 1299
rect 254 1294 260 1295
rect 382 1299 388 1300
rect 382 1295 383 1299
rect 387 1295 388 1299
rect 382 1294 388 1295
rect 494 1299 500 1300
rect 494 1295 495 1299
rect 499 1295 500 1299
rect 494 1294 500 1295
rect 598 1299 604 1300
rect 598 1295 599 1299
rect 603 1295 604 1299
rect 598 1294 604 1295
rect 702 1299 708 1300
rect 702 1295 703 1299
rect 707 1295 708 1299
rect 702 1294 708 1295
rect 798 1299 804 1300
rect 798 1295 799 1299
rect 803 1295 804 1299
rect 798 1294 804 1295
rect 894 1299 900 1300
rect 894 1295 895 1299
rect 899 1295 900 1299
rect 894 1294 900 1295
rect 990 1299 996 1300
rect 990 1295 991 1299
rect 995 1295 996 1299
rect 1286 1296 1287 1300
rect 1291 1296 1292 1300
rect 1286 1295 1292 1296
rect 1328 1295 1330 1315
rect 1598 1314 1604 1315
rect 1662 1319 1668 1320
rect 1662 1315 1663 1319
rect 1667 1315 1668 1319
rect 1662 1314 1668 1315
rect 1742 1319 1748 1320
rect 1742 1315 1743 1319
rect 1747 1315 1748 1319
rect 1742 1314 1748 1315
rect 1822 1319 1828 1320
rect 1822 1315 1823 1319
rect 1827 1315 1828 1319
rect 1822 1314 1828 1315
rect 1910 1319 1916 1320
rect 1910 1315 1911 1319
rect 1915 1315 1916 1319
rect 1910 1314 1916 1315
rect 1998 1319 2004 1320
rect 1998 1315 1999 1319
rect 2003 1315 2004 1319
rect 1998 1314 2004 1315
rect 2078 1319 2084 1320
rect 2078 1315 2079 1319
rect 2083 1315 2084 1319
rect 2078 1314 2084 1315
rect 2158 1319 2164 1320
rect 2158 1315 2159 1319
rect 2163 1315 2164 1319
rect 2158 1314 2164 1315
rect 2238 1319 2244 1320
rect 2238 1315 2239 1319
rect 2243 1315 2244 1319
rect 2238 1314 2244 1315
rect 2318 1319 2324 1320
rect 2318 1315 2319 1319
rect 2323 1315 2324 1319
rect 2318 1314 2324 1315
rect 2398 1319 2404 1320
rect 2398 1315 2399 1319
rect 2403 1315 2404 1319
rect 2398 1314 2404 1315
rect 2454 1319 2460 1320
rect 2454 1315 2455 1319
rect 2459 1315 2460 1319
rect 2502 1316 2503 1320
rect 2507 1316 2508 1320
rect 2502 1315 2508 1316
rect 2454 1314 2460 1315
rect 1600 1295 1602 1314
rect 1664 1295 1666 1314
rect 1744 1295 1746 1314
rect 1824 1295 1826 1314
rect 1912 1295 1914 1314
rect 2000 1295 2002 1314
rect 2080 1295 2082 1314
rect 2160 1295 2162 1314
rect 2240 1295 2242 1314
rect 2320 1295 2322 1314
rect 2400 1295 2402 1314
rect 2456 1295 2458 1314
rect 2504 1295 2506 1315
rect 990 1294 996 1295
rect 152 1267 154 1294
rect 256 1267 258 1294
rect 384 1267 386 1294
rect 496 1267 498 1294
rect 600 1267 602 1294
rect 704 1267 706 1294
rect 800 1267 802 1294
rect 896 1267 898 1294
rect 992 1267 994 1294
rect 1288 1267 1290 1295
rect 1327 1294 1331 1295
rect 1327 1289 1331 1290
rect 1567 1294 1571 1295
rect 1567 1289 1571 1290
rect 1599 1294 1603 1295
rect 1599 1289 1603 1290
rect 1631 1294 1635 1295
rect 1631 1289 1635 1290
rect 1663 1294 1667 1295
rect 1663 1289 1667 1290
rect 1711 1294 1715 1295
rect 1711 1289 1715 1290
rect 1743 1294 1747 1295
rect 1743 1289 1747 1290
rect 1799 1294 1803 1295
rect 1799 1289 1803 1290
rect 1823 1294 1827 1295
rect 1823 1289 1827 1290
rect 1895 1294 1899 1295
rect 1895 1289 1899 1290
rect 1911 1294 1915 1295
rect 1911 1289 1915 1290
rect 1991 1294 1995 1295
rect 1991 1289 1995 1290
rect 1999 1294 2003 1295
rect 1999 1289 2003 1290
rect 2079 1294 2083 1295
rect 2079 1289 2083 1290
rect 2095 1294 2099 1295
rect 2095 1289 2099 1290
rect 2159 1294 2163 1295
rect 2159 1289 2163 1290
rect 2207 1294 2211 1295
rect 2207 1289 2211 1290
rect 2239 1294 2243 1295
rect 2239 1289 2243 1290
rect 2319 1294 2323 1295
rect 2319 1289 2323 1290
rect 2399 1294 2403 1295
rect 2399 1289 2403 1290
rect 2455 1294 2459 1295
rect 2455 1289 2459 1290
rect 2503 1294 2507 1295
rect 2503 1289 2507 1290
rect 1328 1269 1330 1289
rect 1568 1270 1570 1289
rect 1632 1270 1634 1289
rect 1712 1270 1714 1289
rect 1800 1270 1802 1289
rect 1896 1270 1898 1289
rect 1992 1270 1994 1289
rect 2096 1270 2098 1289
rect 2208 1270 2210 1289
rect 2320 1270 2322 1289
rect 1566 1269 1572 1270
rect 1326 1268 1332 1269
rect 111 1266 115 1267
rect 111 1261 115 1262
rect 151 1266 155 1267
rect 151 1261 155 1262
rect 215 1266 219 1267
rect 215 1261 219 1262
rect 255 1266 259 1267
rect 255 1261 259 1262
rect 303 1266 307 1267
rect 303 1261 307 1262
rect 383 1266 387 1267
rect 383 1261 387 1262
rect 391 1266 395 1267
rect 391 1261 395 1262
rect 471 1266 475 1267
rect 471 1261 475 1262
rect 495 1266 499 1267
rect 495 1261 499 1262
rect 551 1266 555 1267
rect 551 1261 555 1262
rect 599 1266 603 1267
rect 599 1261 603 1262
rect 623 1266 627 1267
rect 623 1261 627 1262
rect 695 1266 699 1267
rect 695 1261 699 1262
rect 703 1266 707 1267
rect 703 1261 707 1262
rect 767 1266 771 1267
rect 767 1261 771 1262
rect 799 1266 803 1267
rect 799 1261 803 1262
rect 839 1266 843 1267
rect 839 1261 843 1262
rect 895 1266 899 1267
rect 895 1261 899 1262
rect 919 1266 923 1267
rect 919 1261 923 1262
rect 991 1266 995 1267
rect 991 1261 995 1262
rect 1287 1266 1291 1267
rect 1326 1264 1327 1268
rect 1331 1264 1332 1268
rect 1566 1265 1567 1269
rect 1571 1265 1572 1269
rect 1566 1264 1572 1265
rect 1630 1269 1636 1270
rect 1630 1265 1631 1269
rect 1635 1265 1636 1269
rect 1630 1264 1636 1265
rect 1710 1269 1716 1270
rect 1710 1265 1711 1269
rect 1715 1265 1716 1269
rect 1710 1264 1716 1265
rect 1798 1269 1804 1270
rect 1798 1265 1799 1269
rect 1803 1265 1804 1269
rect 1798 1264 1804 1265
rect 1894 1269 1900 1270
rect 1894 1265 1895 1269
rect 1899 1265 1900 1269
rect 1894 1264 1900 1265
rect 1990 1269 1996 1270
rect 1990 1265 1991 1269
rect 1995 1265 1996 1269
rect 1990 1264 1996 1265
rect 2094 1269 2100 1270
rect 2094 1265 2095 1269
rect 2099 1265 2100 1269
rect 2094 1264 2100 1265
rect 2206 1269 2212 1270
rect 2206 1265 2207 1269
rect 2211 1265 2212 1269
rect 2206 1264 2212 1265
rect 2318 1269 2324 1270
rect 2504 1269 2506 1289
rect 2318 1265 2319 1269
rect 2323 1265 2324 1269
rect 2318 1264 2324 1265
rect 2502 1268 2508 1269
rect 2502 1264 2503 1268
rect 2507 1264 2508 1268
rect 1326 1263 1332 1264
rect 2502 1263 2508 1264
rect 1287 1261 1291 1262
rect 112 1241 114 1261
rect 152 1242 154 1261
rect 216 1242 218 1261
rect 304 1242 306 1261
rect 392 1242 394 1261
rect 472 1242 474 1261
rect 552 1242 554 1261
rect 624 1242 626 1261
rect 696 1242 698 1261
rect 768 1242 770 1261
rect 840 1242 842 1261
rect 920 1242 922 1261
rect 150 1241 156 1242
rect 110 1240 116 1241
rect 110 1236 111 1240
rect 115 1236 116 1240
rect 150 1237 151 1241
rect 155 1237 156 1241
rect 150 1236 156 1237
rect 214 1241 220 1242
rect 214 1237 215 1241
rect 219 1237 220 1241
rect 214 1236 220 1237
rect 302 1241 308 1242
rect 302 1237 303 1241
rect 307 1237 308 1241
rect 302 1236 308 1237
rect 390 1241 396 1242
rect 390 1237 391 1241
rect 395 1237 396 1241
rect 390 1236 396 1237
rect 470 1241 476 1242
rect 470 1237 471 1241
rect 475 1237 476 1241
rect 470 1236 476 1237
rect 550 1241 556 1242
rect 550 1237 551 1241
rect 555 1237 556 1241
rect 550 1236 556 1237
rect 622 1241 628 1242
rect 622 1237 623 1241
rect 627 1237 628 1241
rect 622 1236 628 1237
rect 694 1241 700 1242
rect 694 1237 695 1241
rect 699 1237 700 1241
rect 694 1236 700 1237
rect 766 1241 772 1242
rect 766 1237 767 1241
rect 771 1237 772 1241
rect 766 1236 772 1237
rect 838 1241 844 1242
rect 838 1237 839 1241
rect 843 1237 844 1241
rect 838 1236 844 1237
rect 918 1241 924 1242
rect 1288 1241 1290 1261
rect 1326 1251 1332 1252
rect 1326 1247 1327 1251
rect 1331 1247 1332 1251
rect 2502 1251 2508 1252
rect 1326 1246 1332 1247
rect 1550 1248 1556 1249
rect 918 1237 919 1241
rect 923 1237 924 1241
rect 918 1236 924 1237
rect 1286 1240 1292 1241
rect 1286 1236 1287 1240
rect 1291 1236 1292 1240
rect 1328 1239 1330 1246
rect 1550 1244 1551 1248
rect 1555 1244 1556 1248
rect 1550 1243 1556 1244
rect 1614 1248 1620 1249
rect 1614 1244 1615 1248
rect 1619 1244 1620 1248
rect 1614 1243 1620 1244
rect 1694 1248 1700 1249
rect 1694 1244 1695 1248
rect 1699 1244 1700 1248
rect 1694 1243 1700 1244
rect 1782 1248 1788 1249
rect 1782 1244 1783 1248
rect 1787 1244 1788 1248
rect 1782 1243 1788 1244
rect 1878 1248 1884 1249
rect 1878 1244 1879 1248
rect 1883 1244 1884 1248
rect 1878 1243 1884 1244
rect 1974 1248 1980 1249
rect 1974 1244 1975 1248
rect 1979 1244 1980 1248
rect 1974 1243 1980 1244
rect 2078 1248 2084 1249
rect 2078 1244 2079 1248
rect 2083 1244 2084 1248
rect 2078 1243 2084 1244
rect 2190 1248 2196 1249
rect 2190 1244 2191 1248
rect 2195 1244 2196 1248
rect 2190 1243 2196 1244
rect 2302 1248 2308 1249
rect 2302 1244 2303 1248
rect 2307 1244 2308 1248
rect 2502 1247 2503 1251
rect 2507 1247 2508 1251
rect 2502 1246 2508 1247
rect 2302 1243 2308 1244
rect 1552 1239 1554 1243
rect 1616 1239 1618 1243
rect 1696 1239 1698 1243
rect 1784 1239 1786 1243
rect 1880 1239 1882 1243
rect 1976 1239 1978 1243
rect 2080 1239 2082 1243
rect 2192 1239 2194 1243
rect 2304 1239 2306 1243
rect 2504 1239 2506 1246
rect 110 1235 116 1236
rect 1286 1235 1292 1236
rect 1327 1238 1331 1239
rect 1327 1233 1331 1234
rect 1519 1238 1523 1239
rect 1519 1233 1523 1234
rect 1551 1238 1555 1239
rect 1551 1233 1555 1234
rect 1575 1238 1579 1239
rect 1575 1233 1579 1234
rect 1615 1238 1619 1239
rect 1615 1233 1619 1234
rect 1631 1238 1635 1239
rect 1631 1233 1635 1234
rect 1687 1238 1691 1239
rect 1687 1233 1691 1234
rect 1695 1238 1699 1239
rect 1695 1233 1699 1234
rect 1743 1238 1747 1239
rect 1743 1233 1747 1234
rect 1783 1238 1787 1239
rect 1783 1233 1787 1234
rect 1799 1238 1803 1239
rect 1799 1233 1803 1234
rect 1855 1238 1859 1239
rect 1855 1233 1859 1234
rect 1879 1238 1883 1239
rect 1879 1233 1883 1234
rect 1911 1238 1915 1239
rect 1911 1233 1915 1234
rect 1967 1238 1971 1239
rect 1967 1233 1971 1234
rect 1975 1238 1979 1239
rect 1975 1233 1979 1234
rect 2031 1238 2035 1239
rect 2031 1233 2035 1234
rect 2079 1238 2083 1239
rect 2079 1233 2083 1234
rect 2103 1238 2107 1239
rect 2103 1233 2107 1234
rect 2183 1238 2187 1239
rect 2183 1233 2187 1234
rect 2191 1238 2195 1239
rect 2191 1233 2195 1234
rect 2271 1238 2275 1239
rect 2271 1233 2275 1234
rect 2303 1238 2307 1239
rect 2303 1233 2307 1234
rect 2367 1238 2371 1239
rect 2367 1233 2371 1234
rect 2439 1238 2443 1239
rect 2439 1233 2443 1234
rect 2503 1238 2507 1239
rect 2503 1233 2507 1234
rect 1328 1230 1330 1233
rect 1518 1232 1524 1233
rect 1326 1229 1332 1230
rect 1326 1225 1327 1229
rect 1331 1225 1332 1229
rect 1518 1228 1519 1232
rect 1523 1228 1524 1232
rect 1518 1227 1524 1228
rect 1574 1232 1580 1233
rect 1574 1228 1575 1232
rect 1579 1228 1580 1232
rect 1574 1227 1580 1228
rect 1630 1232 1636 1233
rect 1630 1228 1631 1232
rect 1635 1228 1636 1232
rect 1630 1227 1636 1228
rect 1686 1232 1692 1233
rect 1686 1228 1687 1232
rect 1691 1228 1692 1232
rect 1686 1227 1692 1228
rect 1742 1232 1748 1233
rect 1742 1228 1743 1232
rect 1747 1228 1748 1232
rect 1742 1227 1748 1228
rect 1798 1232 1804 1233
rect 1798 1228 1799 1232
rect 1803 1228 1804 1232
rect 1798 1227 1804 1228
rect 1854 1232 1860 1233
rect 1854 1228 1855 1232
rect 1859 1228 1860 1232
rect 1854 1227 1860 1228
rect 1910 1232 1916 1233
rect 1910 1228 1911 1232
rect 1915 1228 1916 1232
rect 1910 1227 1916 1228
rect 1966 1232 1972 1233
rect 1966 1228 1967 1232
rect 1971 1228 1972 1232
rect 1966 1227 1972 1228
rect 2030 1232 2036 1233
rect 2030 1228 2031 1232
rect 2035 1228 2036 1232
rect 2030 1227 2036 1228
rect 2102 1232 2108 1233
rect 2102 1228 2103 1232
rect 2107 1228 2108 1232
rect 2102 1227 2108 1228
rect 2182 1232 2188 1233
rect 2182 1228 2183 1232
rect 2187 1228 2188 1232
rect 2182 1227 2188 1228
rect 2270 1232 2276 1233
rect 2270 1228 2271 1232
rect 2275 1228 2276 1232
rect 2270 1227 2276 1228
rect 2366 1232 2372 1233
rect 2366 1228 2367 1232
rect 2371 1228 2372 1232
rect 2366 1227 2372 1228
rect 2438 1232 2444 1233
rect 2438 1228 2439 1232
rect 2443 1228 2444 1232
rect 2504 1230 2506 1233
rect 2438 1227 2444 1228
rect 2502 1229 2508 1230
rect 1326 1224 1332 1225
rect 2502 1225 2503 1229
rect 2507 1225 2508 1229
rect 2502 1224 2508 1225
rect 110 1223 116 1224
rect 110 1219 111 1223
rect 115 1219 116 1223
rect 1286 1223 1292 1224
rect 110 1218 116 1219
rect 134 1220 140 1221
rect 112 1211 114 1218
rect 134 1216 135 1220
rect 139 1216 140 1220
rect 134 1215 140 1216
rect 198 1220 204 1221
rect 198 1216 199 1220
rect 203 1216 204 1220
rect 198 1215 204 1216
rect 286 1220 292 1221
rect 286 1216 287 1220
rect 291 1216 292 1220
rect 286 1215 292 1216
rect 374 1220 380 1221
rect 374 1216 375 1220
rect 379 1216 380 1220
rect 374 1215 380 1216
rect 454 1220 460 1221
rect 454 1216 455 1220
rect 459 1216 460 1220
rect 454 1215 460 1216
rect 534 1220 540 1221
rect 534 1216 535 1220
rect 539 1216 540 1220
rect 534 1215 540 1216
rect 606 1220 612 1221
rect 606 1216 607 1220
rect 611 1216 612 1220
rect 606 1215 612 1216
rect 678 1220 684 1221
rect 678 1216 679 1220
rect 683 1216 684 1220
rect 678 1215 684 1216
rect 750 1220 756 1221
rect 750 1216 751 1220
rect 755 1216 756 1220
rect 750 1215 756 1216
rect 822 1220 828 1221
rect 822 1216 823 1220
rect 827 1216 828 1220
rect 822 1215 828 1216
rect 902 1220 908 1221
rect 902 1216 903 1220
rect 907 1216 908 1220
rect 1286 1219 1287 1223
rect 1291 1219 1292 1223
rect 1286 1218 1292 1219
rect 902 1215 908 1216
rect 136 1211 138 1215
rect 200 1211 202 1215
rect 288 1211 290 1215
rect 376 1211 378 1215
rect 456 1211 458 1215
rect 536 1211 538 1215
rect 608 1211 610 1215
rect 680 1211 682 1215
rect 752 1211 754 1215
rect 824 1211 826 1215
rect 904 1211 906 1215
rect 1288 1211 1290 1218
rect 1326 1212 1332 1213
rect 2502 1212 2508 1213
rect 111 1210 115 1211
rect 111 1205 115 1206
rect 135 1210 139 1211
rect 135 1205 139 1206
rect 191 1210 195 1211
rect 191 1205 195 1206
rect 199 1210 203 1211
rect 199 1205 203 1206
rect 271 1210 275 1211
rect 271 1205 275 1206
rect 287 1210 291 1211
rect 287 1205 291 1206
rect 351 1210 355 1211
rect 351 1205 355 1206
rect 375 1210 379 1211
rect 375 1205 379 1206
rect 431 1210 435 1211
rect 431 1205 435 1206
rect 455 1210 459 1211
rect 455 1205 459 1206
rect 511 1210 515 1211
rect 511 1205 515 1206
rect 535 1210 539 1211
rect 535 1205 539 1206
rect 583 1210 587 1211
rect 583 1205 587 1206
rect 607 1210 611 1211
rect 607 1205 611 1206
rect 647 1210 651 1211
rect 647 1205 651 1206
rect 679 1210 683 1211
rect 679 1205 683 1206
rect 719 1210 723 1211
rect 719 1205 723 1206
rect 751 1210 755 1211
rect 751 1205 755 1206
rect 791 1210 795 1211
rect 791 1205 795 1206
rect 823 1210 827 1211
rect 823 1205 827 1206
rect 863 1210 867 1211
rect 863 1205 867 1206
rect 903 1210 907 1211
rect 903 1205 907 1206
rect 1287 1210 1291 1211
rect 1326 1208 1327 1212
rect 1331 1208 1332 1212
rect 1326 1207 1332 1208
rect 1534 1211 1540 1212
rect 1534 1207 1535 1211
rect 1539 1207 1540 1211
rect 1287 1205 1291 1206
rect 112 1202 114 1205
rect 134 1204 140 1205
rect 110 1201 116 1202
rect 110 1197 111 1201
rect 115 1197 116 1201
rect 134 1200 135 1204
rect 139 1200 140 1204
rect 134 1199 140 1200
rect 190 1204 196 1205
rect 190 1200 191 1204
rect 195 1200 196 1204
rect 190 1199 196 1200
rect 270 1204 276 1205
rect 270 1200 271 1204
rect 275 1200 276 1204
rect 270 1199 276 1200
rect 350 1204 356 1205
rect 350 1200 351 1204
rect 355 1200 356 1204
rect 350 1199 356 1200
rect 430 1204 436 1205
rect 430 1200 431 1204
rect 435 1200 436 1204
rect 430 1199 436 1200
rect 510 1204 516 1205
rect 510 1200 511 1204
rect 515 1200 516 1204
rect 510 1199 516 1200
rect 582 1204 588 1205
rect 582 1200 583 1204
rect 587 1200 588 1204
rect 582 1199 588 1200
rect 646 1204 652 1205
rect 646 1200 647 1204
rect 651 1200 652 1204
rect 646 1199 652 1200
rect 718 1204 724 1205
rect 718 1200 719 1204
rect 723 1200 724 1204
rect 718 1199 724 1200
rect 790 1204 796 1205
rect 790 1200 791 1204
rect 795 1200 796 1204
rect 790 1199 796 1200
rect 862 1204 868 1205
rect 862 1200 863 1204
rect 867 1200 868 1204
rect 1288 1202 1290 1205
rect 862 1199 868 1200
rect 1286 1201 1292 1202
rect 110 1196 116 1197
rect 1286 1197 1287 1201
rect 1291 1197 1292 1201
rect 1286 1196 1292 1197
rect 110 1184 116 1185
rect 1286 1184 1292 1185
rect 110 1180 111 1184
rect 115 1180 116 1184
rect 110 1179 116 1180
rect 150 1183 156 1184
rect 150 1179 151 1183
rect 155 1179 156 1183
rect 112 1155 114 1179
rect 150 1178 156 1179
rect 206 1183 212 1184
rect 206 1179 207 1183
rect 211 1179 212 1183
rect 206 1178 212 1179
rect 286 1183 292 1184
rect 286 1179 287 1183
rect 291 1179 292 1183
rect 286 1178 292 1179
rect 366 1183 372 1184
rect 366 1179 367 1183
rect 371 1179 372 1183
rect 366 1178 372 1179
rect 446 1183 452 1184
rect 446 1179 447 1183
rect 451 1179 452 1183
rect 446 1178 452 1179
rect 526 1183 532 1184
rect 526 1179 527 1183
rect 531 1179 532 1183
rect 526 1178 532 1179
rect 598 1183 604 1184
rect 598 1179 599 1183
rect 603 1179 604 1183
rect 598 1178 604 1179
rect 662 1183 668 1184
rect 662 1179 663 1183
rect 667 1179 668 1183
rect 662 1178 668 1179
rect 734 1183 740 1184
rect 734 1179 735 1183
rect 739 1179 740 1183
rect 734 1178 740 1179
rect 806 1183 812 1184
rect 806 1179 807 1183
rect 811 1179 812 1183
rect 806 1178 812 1179
rect 878 1183 884 1184
rect 878 1179 879 1183
rect 883 1179 884 1183
rect 1286 1180 1287 1184
rect 1291 1180 1292 1184
rect 1328 1183 1330 1207
rect 1534 1206 1540 1207
rect 1590 1211 1596 1212
rect 1590 1207 1591 1211
rect 1595 1207 1596 1211
rect 1590 1206 1596 1207
rect 1646 1211 1652 1212
rect 1646 1207 1647 1211
rect 1651 1207 1652 1211
rect 1646 1206 1652 1207
rect 1702 1211 1708 1212
rect 1702 1207 1703 1211
rect 1707 1207 1708 1211
rect 1702 1206 1708 1207
rect 1758 1211 1764 1212
rect 1758 1207 1759 1211
rect 1763 1207 1764 1211
rect 1758 1206 1764 1207
rect 1814 1211 1820 1212
rect 1814 1207 1815 1211
rect 1819 1207 1820 1211
rect 1814 1206 1820 1207
rect 1870 1211 1876 1212
rect 1870 1207 1871 1211
rect 1875 1207 1876 1211
rect 1870 1206 1876 1207
rect 1926 1211 1932 1212
rect 1926 1207 1927 1211
rect 1931 1207 1932 1211
rect 1926 1206 1932 1207
rect 1982 1211 1988 1212
rect 1982 1207 1983 1211
rect 1987 1207 1988 1211
rect 1982 1206 1988 1207
rect 2046 1211 2052 1212
rect 2046 1207 2047 1211
rect 2051 1207 2052 1211
rect 2046 1206 2052 1207
rect 2118 1211 2124 1212
rect 2118 1207 2119 1211
rect 2123 1207 2124 1211
rect 2118 1206 2124 1207
rect 2198 1211 2204 1212
rect 2198 1207 2199 1211
rect 2203 1207 2204 1211
rect 2198 1206 2204 1207
rect 2286 1211 2292 1212
rect 2286 1207 2287 1211
rect 2291 1207 2292 1211
rect 2286 1206 2292 1207
rect 2382 1211 2388 1212
rect 2382 1207 2383 1211
rect 2387 1207 2388 1211
rect 2382 1206 2388 1207
rect 2454 1211 2460 1212
rect 2454 1207 2455 1211
rect 2459 1207 2460 1211
rect 2502 1208 2503 1212
rect 2507 1208 2508 1212
rect 2502 1207 2508 1208
rect 2454 1206 2460 1207
rect 1536 1183 1538 1206
rect 1592 1183 1594 1206
rect 1648 1183 1650 1206
rect 1704 1183 1706 1206
rect 1760 1183 1762 1206
rect 1816 1183 1818 1206
rect 1872 1183 1874 1206
rect 1928 1183 1930 1206
rect 1984 1183 1986 1206
rect 2048 1183 2050 1206
rect 2120 1183 2122 1206
rect 2200 1183 2202 1206
rect 2288 1183 2290 1206
rect 2384 1183 2386 1206
rect 2456 1183 2458 1206
rect 2504 1183 2506 1207
rect 1286 1179 1292 1180
rect 1327 1182 1331 1183
rect 878 1178 884 1179
rect 152 1155 154 1178
rect 208 1155 210 1178
rect 288 1155 290 1178
rect 368 1155 370 1178
rect 448 1155 450 1178
rect 528 1155 530 1178
rect 600 1155 602 1178
rect 664 1155 666 1178
rect 736 1155 738 1178
rect 808 1155 810 1178
rect 880 1155 882 1178
rect 1288 1155 1290 1179
rect 1327 1177 1331 1178
rect 1535 1182 1539 1183
rect 1535 1177 1539 1178
rect 1567 1182 1571 1183
rect 1567 1177 1571 1178
rect 1591 1182 1595 1183
rect 1591 1177 1595 1178
rect 1631 1182 1635 1183
rect 1631 1177 1635 1178
rect 1647 1182 1651 1183
rect 1647 1177 1651 1178
rect 1703 1182 1707 1183
rect 1703 1177 1707 1178
rect 1759 1182 1763 1183
rect 1759 1177 1763 1178
rect 1791 1182 1795 1183
rect 1791 1177 1795 1178
rect 1815 1182 1819 1183
rect 1815 1177 1819 1178
rect 1871 1182 1875 1183
rect 1871 1177 1875 1178
rect 1903 1182 1907 1183
rect 1903 1177 1907 1178
rect 1927 1182 1931 1183
rect 1927 1177 1931 1178
rect 1983 1182 1987 1183
rect 1983 1177 1987 1178
rect 2031 1182 2035 1183
rect 2031 1177 2035 1178
rect 2047 1182 2051 1183
rect 2047 1177 2051 1178
rect 2119 1182 2123 1183
rect 2119 1177 2123 1178
rect 2175 1182 2179 1183
rect 2175 1177 2179 1178
rect 2199 1182 2203 1183
rect 2199 1177 2203 1178
rect 2287 1182 2291 1183
rect 2287 1177 2291 1178
rect 2327 1182 2331 1183
rect 2327 1177 2331 1178
rect 2383 1182 2387 1183
rect 2383 1177 2387 1178
rect 2455 1182 2459 1183
rect 2455 1177 2459 1178
rect 2503 1182 2507 1183
rect 2503 1177 2507 1178
rect 1328 1157 1330 1177
rect 1568 1158 1570 1177
rect 1632 1158 1634 1177
rect 1704 1158 1706 1177
rect 1792 1158 1794 1177
rect 1904 1158 1906 1177
rect 2032 1158 2034 1177
rect 2176 1158 2178 1177
rect 2328 1158 2330 1177
rect 2456 1158 2458 1177
rect 1566 1157 1572 1158
rect 1326 1156 1332 1157
rect 111 1154 115 1155
rect 111 1149 115 1150
rect 151 1154 155 1155
rect 151 1149 155 1150
rect 183 1154 187 1155
rect 183 1149 187 1150
rect 207 1154 211 1155
rect 207 1149 211 1150
rect 279 1154 283 1155
rect 279 1149 283 1150
rect 287 1154 291 1155
rect 287 1149 291 1150
rect 367 1154 371 1155
rect 367 1149 371 1150
rect 375 1154 379 1155
rect 375 1149 379 1150
rect 447 1154 451 1155
rect 447 1149 451 1150
rect 471 1154 475 1155
rect 471 1149 475 1150
rect 527 1154 531 1155
rect 527 1149 531 1150
rect 567 1154 571 1155
rect 567 1149 571 1150
rect 599 1154 603 1155
rect 599 1149 603 1150
rect 655 1154 659 1155
rect 655 1149 659 1150
rect 663 1154 667 1155
rect 663 1149 667 1150
rect 735 1154 739 1155
rect 735 1149 739 1150
rect 807 1154 811 1155
rect 807 1149 811 1150
rect 879 1154 883 1155
rect 879 1149 883 1150
rect 959 1154 963 1155
rect 959 1149 963 1150
rect 1039 1154 1043 1155
rect 1039 1149 1043 1150
rect 1287 1154 1291 1155
rect 1326 1152 1327 1156
rect 1331 1152 1332 1156
rect 1566 1153 1567 1157
rect 1571 1153 1572 1157
rect 1566 1152 1572 1153
rect 1630 1157 1636 1158
rect 1630 1153 1631 1157
rect 1635 1153 1636 1157
rect 1630 1152 1636 1153
rect 1702 1157 1708 1158
rect 1702 1153 1703 1157
rect 1707 1153 1708 1157
rect 1702 1152 1708 1153
rect 1790 1157 1796 1158
rect 1790 1153 1791 1157
rect 1795 1153 1796 1157
rect 1790 1152 1796 1153
rect 1902 1157 1908 1158
rect 1902 1153 1903 1157
rect 1907 1153 1908 1157
rect 1902 1152 1908 1153
rect 2030 1157 2036 1158
rect 2030 1153 2031 1157
rect 2035 1153 2036 1157
rect 2030 1152 2036 1153
rect 2174 1157 2180 1158
rect 2174 1153 2175 1157
rect 2179 1153 2180 1157
rect 2174 1152 2180 1153
rect 2326 1157 2332 1158
rect 2326 1153 2327 1157
rect 2331 1153 2332 1157
rect 2326 1152 2332 1153
rect 2454 1157 2460 1158
rect 2504 1157 2506 1177
rect 2454 1153 2455 1157
rect 2459 1153 2460 1157
rect 2454 1152 2460 1153
rect 2502 1156 2508 1157
rect 2502 1152 2503 1156
rect 2507 1152 2508 1156
rect 1326 1151 1332 1152
rect 2502 1151 2508 1152
rect 1287 1149 1291 1150
rect 112 1129 114 1149
rect 184 1130 186 1149
rect 280 1130 282 1149
rect 376 1130 378 1149
rect 472 1130 474 1149
rect 568 1130 570 1149
rect 656 1130 658 1149
rect 736 1130 738 1149
rect 808 1130 810 1149
rect 880 1130 882 1149
rect 960 1130 962 1149
rect 1040 1130 1042 1149
rect 182 1129 188 1130
rect 110 1128 116 1129
rect 110 1124 111 1128
rect 115 1124 116 1128
rect 182 1125 183 1129
rect 187 1125 188 1129
rect 182 1124 188 1125
rect 278 1129 284 1130
rect 278 1125 279 1129
rect 283 1125 284 1129
rect 278 1124 284 1125
rect 374 1129 380 1130
rect 374 1125 375 1129
rect 379 1125 380 1129
rect 374 1124 380 1125
rect 470 1129 476 1130
rect 470 1125 471 1129
rect 475 1125 476 1129
rect 470 1124 476 1125
rect 566 1129 572 1130
rect 566 1125 567 1129
rect 571 1125 572 1129
rect 566 1124 572 1125
rect 654 1129 660 1130
rect 654 1125 655 1129
rect 659 1125 660 1129
rect 654 1124 660 1125
rect 734 1129 740 1130
rect 734 1125 735 1129
rect 739 1125 740 1129
rect 734 1124 740 1125
rect 806 1129 812 1130
rect 806 1125 807 1129
rect 811 1125 812 1129
rect 806 1124 812 1125
rect 878 1129 884 1130
rect 878 1125 879 1129
rect 883 1125 884 1129
rect 878 1124 884 1125
rect 958 1129 964 1130
rect 958 1125 959 1129
rect 963 1125 964 1129
rect 958 1124 964 1125
rect 1038 1129 1044 1130
rect 1288 1129 1290 1149
rect 1326 1139 1332 1140
rect 1326 1135 1327 1139
rect 1331 1135 1332 1139
rect 2502 1139 2508 1140
rect 1326 1134 1332 1135
rect 1550 1136 1556 1137
rect 1328 1131 1330 1134
rect 1550 1132 1551 1136
rect 1555 1132 1556 1136
rect 1550 1131 1556 1132
rect 1614 1136 1620 1137
rect 1614 1132 1615 1136
rect 1619 1132 1620 1136
rect 1614 1131 1620 1132
rect 1686 1136 1692 1137
rect 1686 1132 1687 1136
rect 1691 1132 1692 1136
rect 1686 1131 1692 1132
rect 1774 1136 1780 1137
rect 1774 1132 1775 1136
rect 1779 1132 1780 1136
rect 1774 1131 1780 1132
rect 1886 1136 1892 1137
rect 1886 1132 1887 1136
rect 1891 1132 1892 1136
rect 1886 1131 1892 1132
rect 2014 1136 2020 1137
rect 2014 1132 2015 1136
rect 2019 1132 2020 1136
rect 2014 1131 2020 1132
rect 2158 1136 2164 1137
rect 2158 1132 2159 1136
rect 2163 1132 2164 1136
rect 2158 1131 2164 1132
rect 2310 1136 2316 1137
rect 2310 1132 2311 1136
rect 2315 1132 2316 1136
rect 2310 1131 2316 1132
rect 2438 1136 2444 1137
rect 2438 1132 2439 1136
rect 2443 1132 2444 1136
rect 2502 1135 2503 1139
rect 2507 1135 2508 1139
rect 2502 1134 2508 1135
rect 2438 1131 2444 1132
rect 2504 1131 2506 1134
rect 1327 1130 1331 1131
rect 1038 1125 1039 1129
rect 1043 1125 1044 1129
rect 1038 1124 1044 1125
rect 1286 1128 1292 1129
rect 1286 1124 1287 1128
rect 1291 1124 1292 1128
rect 1327 1125 1331 1126
rect 1383 1130 1387 1131
rect 1383 1125 1387 1126
rect 1447 1130 1451 1131
rect 1447 1125 1451 1126
rect 1519 1130 1523 1131
rect 1519 1125 1523 1126
rect 1551 1130 1555 1131
rect 1551 1125 1555 1126
rect 1591 1130 1595 1131
rect 1591 1125 1595 1126
rect 1615 1130 1619 1131
rect 1615 1125 1619 1126
rect 1671 1130 1675 1131
rect 1671 1125 1675 1126
rect 1687 1130 1691 1131
rect 1687 1125 1691 1126
rect 1751 1130 1755 1131
rect 1751 1125 1755 1126
rect 1775 1130 1779 1131
rect 1775 1125 1779 1126
rect 1831 1130 1835 1131
rect 1831 1125 1835 1126
rect 1887 1130 1891 1131
rect 1887 1125 1891 1126
rect 1911 1130 1915 1131
rect 1911 1125 1915 1126
rect 1983 1130 1987 1131
rect 1983 1125 1987 1126
rect 2015 1130 2019 1131
rect 2015 1125 2019 1126
rect 2055 1130 2059 1131
rect 2055 1125 2059 1126
rect 2135 1130 2139 1131
rect 2135 1125 2139 1126
rect 2159 1130 2163 1131
rect 2159 1125 2163 1126
rect 2215 1130 2219 1131
rect 2215 1125 2219 1126
rect 2311 1130 2315 1131
rect 2311 1125 2315 1126
rect 2439 1130 2443 1131
rect 2439 1125 2443 1126
rect 2503 1130 2507 1131
rect 2503 1125 2507 1126
rect 110 1123 116 1124
rect 1286 1123 1292 1124
rect 1328 1122 1330 1125
rect 1382 1124 1388 1125
rect 1326 1121 1332 1122
rect 1326 1117 1327 1121
rect 1331 1117 1332 1121
rect 1382 1120 1383 1124
rect 1387 1120 1388 1124
rect 1382 1119 1388 1120
rect 1446 1124 1452 1125
rect 1446 1120 1447 1124
rect 1451 1120 1452 1124
rect 1446 1119 1452 1120
rect 1518 1124 1524 1125
rect 1518 1120 1519 1124
rect 1523 1120 1524 1124
rect 1518 1119 1524 1120
rect 1590 1124 1596 1125
rect 1590 1120 1591 1124
rect 1595 1120 1596 1124
rect 1590 1119 1596 1120
rect 1670 1124 1676 1125
rect 1670 1120 1671 1124
rect 1675 1120 1676 1124
rect 1670 1119 1676 1120
rect 1750 1124 1756 1125
rect 1750 1120 1751 1124
rect 1755 1120 1756 1124
rect 1750 1119 1756 1120
rect 1830 1124 1836 1125
rect 1830 1120 1831 1124
rect 1835 1120 1836 1124
rect 1830 1119 1836 1120
rect 1910 1124 1916 1125
rect 1910 1120 1911 1124
rect 1915 1120 1916 1124
rect 1910 1119 1916 1120
rect 1982 1124 1988 1125
rect 1982 1120 1983 1124
rect 1987 1120 1988 1124
rect 1982 1119 1988 1120
rect 2054 1124 2060 1125
rect 2054 1120 2055 1124
rect 2059 1120 2060 1124
rect 2054 1119 2060 1120
rect 2134 1124 2140 1125
rect 2134 1120 2135 1124
rect 2139 1120 2140 1124
rect 2134 1119 2140 1120
rect 2214 1124 2220 1125
rect 2214 1120 2215 1124
rect 2219 1120 2220 1124
rect 2504 1122 2506 1125
rect 2214 1119 2220 1120
rect 2502 1121 2508 1122
rect 1326 1116 1332 1117
rect 2502 1117 2503 1121
rect 2507 1117 2508 1121
rect 2502 1116 2508 1117
rect 110 1111 116 1112
rect 110 1107 111 1111
rect 115 1107 116 1111
rect 1286 1111 1292 1112
rect 110 1106 116 1107
rect 166 1108 172 1109
rect 112 1095 114 1106
rect 166 1104 167 1108
rect 171 1104 172 1108
rect 166 1103 172 1104
rect 262 1108 268 1109
rect 262 1104 263 1108
rect 267 1104 268 1108
rect 262 1103 268 1104
rect 358 1108 364 1109
rect 358 1104 359 1108
rect 363 1104 364 1108
rect 358 1103 364 1104
rect 454 1108 460 1109
rect 454 1104 455 1108
rect 459 1104 460 1108
rect 454 1103 460 1104
rect 550 1108 556 1109
rect 550 1104 551 1108
rect 555 1104 556 1108
rect 550 1103 556 1104
rect 638 1108 644 1109
rect 638 1104 639 1108
rect 643 1104 644 1108
rect 638 1103 644 1104
rect 718 1108 724 1109
rect 718 1104 719 1108
rect 723 1104 724 1108
rect 718 1103 724 1104
rect 790 1108 796 1109
rect 790 1104 791 1108
rect 795 1104 796 1108
rect 790 1103 796 1104
rect 862 1108 868 1109
rect 862 1104 863 1108
rect 867 1104 868 1108
rect 862 1103 868 1104
rect 942 1108 948 1109
rect 942 1104 943 1108
rect 947 1104 948 1108
rect 942 1103 948 1104
rect 1022 1108 1028 1109
rect 1022 1104 1023 1108
rect 1027 1104 1028 1108
rect 1286 1107 1287 1111
rect 1291 1107 1292 1111
rect 1286 1106 1292 1107
rect 1022 1103 1028 1104
rect 168 1095 170 1103
rect 264 1095 266 1103
rect 360 1095 362 1103
rect 456 1095 458 1103
rect 552 1095 554 1103
rect 640 1095 642 1103
rect 720 1095 722 1103
rect 792 1095 794 1103
rect 864 1095 866 1103
rect 944 1095 946 1103
rect 1024 1095 1026 1103
rect 1288 1095 1290 1106
rect 1326 1104 1332 1105
rect 2502 1104 2508 1105
rect 1326 1100 1327 1104
rect 1331 1100 1332 1104
rect 1326 1099 1332 1100
rect 1398 1103 1404 1104
rect 1398 1099 1399 1103
rect 1403 1099 1404 1103
rect 111 1094 115 1095
rect 111 1089 115 1090
rect 167 1094 171 1095
rect 167 1089 171 1090
rect 207 1094 211 1095
rect 207 1089 211 1090
rect 263 1094 267 1095
rect 263 1089 267 1090
rect 279 1094 283 1095
rect 279 1089 283 1090
rect 359 1094 363 1095
rect 359 1089 363 1090
rect 447 1094 451 1095
rect 447 1089 451 1090
rect 455 1094 459 1095
rect 455 1089 459 1090
rect 543 1094 547 1095
rect 543 1089 547 1090
rect 551 1094 555 1095
rect 551 1089 555 1090
rect 639 1094 643 1095
rect 639 1089 643 1090
rect 719 1094 723 1095
rect 719 1089 723 1090
rect 727 1094 731 1095
rect 727 1089 731 1090
rect 791 1094 795 1095
rect 791 1089 795 1090
rect 815 1094 819 1095
rect 815 1089 819 1090
rect 863 1094 867 1095
rect 863 1089 867 1090
rect 895 1094 899 1095
rect 895 1089 899 1090
rect 943 1094 947 1095
rect 943 1089 947 1090
rect 975 1094 979 1095
rect 975 1089 979 1090
rect 1023 1094 1027 1095
rect 1023 1089 1027 1090
rect 1055 1094 1059 1095
rect 1055 1089 1059 1090
rect 1143 1094 1147 1095
rect 1143 1089 1147 1090
rect 1287 1094 1291 1095
rect 1287 1089 1291 1090
rect 112 1086 114 1089
rect 206 1088 212 1089
rect 110 1085 116 1086
rect 110 1081 111 1085
rect 115 1081 116 1085
rect 206 1084 207 1088
rect 211 1084 212 1088
rect 206 1083 212 1084
rect 278 1088 284 1089
rect 278 1084 279 1088
rect 283 1084 284 1088
rect 278 1083 284 1084
rect 358 1088 364 1089
rect 358 1084 359 1088
rect 363 1084 364 1088
rect 358 1083 364 1084
rect 446 1088 452 1089
rect 446 1084 447 1088
rect 451 1084 452 1088
rect 446 1083 452 1084
rect 542 1088 548 1089
rect 542 1084 543 1088
rect 547 1084 548 1088
rect 542 1083 548 1084
rect 638 1088 644 1089
rect 638 1084 639 1088
rect 643 1084 644 1088
rect 638 1083 644 1084
rect 726 1088 732 1089
rect 726 1084 727 1088
rect 731 1084 732 1088
rect 726 1083 732 1084
rect 814 1088 820 1089
rect 814 1084 815 1088
rect 819 1084 820 1088
rect 814 1083 820 1084
rect 894 1088 900 1089
rect 894 1084 895 1088
rect 899 1084 900 1088
rect 894 1083 900 1084
rect 974 1088 980 1089
rect 974 1084 975 1088
rect 979 1084 980 1088
rect 974 1083 980 1084
rect 1054 1088 1060 1089
rect 1054 1084 1055 1088
rect 1059 1084 1060 1088
rect 1054 1083 1060 1084
rect 1142 1088 1148 1089
rect 1142 1084 1143 1088
rect 1147 1084 1148 1088
rect 1288 1086 1290 1089
rect 1142 1083 1148 1084
rect 1286 1085 1292 1086
rect 110 1080 116 1081
rect 1286 1081 1287 1085
rect 1291 1081 1292 1085
rect 1286 1080 1292 1081
rect 1328 1071 1330 1099
rect 1398 1098 1404 1099
rect 1462 1103 1468 1104
rect 1462 1099 1463 1103
rect 1467 1099 1468 1103
rect 1462 1098 1468 1099
rect 1534 1103 1540 1104
rect 1534 1099 1535 1103
rect 1539 1099 1540 1103
rect 1534 1098 1540 1099
rect 1606 1103 1612 1104
rect 1606 1099 1607 1103
rect 1611 1099 1612 1103
rect 1606 1098 1612 1099
rect 1686 1103 1692 1104
rect 1686 1099 1687 1103
rect 1691 1099 1692 1103
rect 1686 1098 1692 1099
rect 1766 1103 1772 1104
rect 1766 1099 1767 1103
rect 1771 1099 1772 1103
rect 1766 1098 1772 1099
rect 1846 1103 1852 1104
rect 1846 1099 1847 1103
rect 1851 1099 1852 1103
rect 1846 1098 1852 1099
rect 1926 1103 1932 1104
rect 1926 1099 1927 1103
rect 1931 1099 1932 1103
rect 1926 1098 1932 1099
rect 1998 1103 2004 1104
rect 1998 1099 1999 1103
rect 2003 1099 2004 1103
rect 1998 1098 2004 1099
rect 2070 1103 2076 1104
rect 2070 1099 2071 1103
rect 2075 1099 2076 1103
rect 2070 1098 2076 1099
rect 2150 1103 2156 1104
rect 2150 1099 2151 1103
rect 2155 1099 2156 1103
rect 2150 1098 2156 1099
rect 2230 1103 2236 1104
rect 2230 1099 2231 1103
rect 2235 1099 2236 1103
rect 2502 1100 2503 1104
rect 2507 1100 2508 1104
rect 2502 1099 2508 1100
rect 2230 1098 2236 1099
rect 1400 1071 1402 1098
rect 1464 1071 1466 1098
rect 1536 1071 1538 1098
rect 1608 1071 1610 1098
rect 1688 1071 1690 1098
rect 1768 1071 1770 1098
rect 1848 1071 1850 1098
rect 1928 1071 1930 1098
rect 2000 1071 2002 1098
rect 2072 1071 2074 1098
rect 2152 1071 2154 1098
rect 2232 1071 2234 1098
rect 2504 1071 2506 1099
rect 1327 1070 1331 1071
rect 110 1068 116 1069
rect 1286 1068 1292 1069
rect 110 1064 111 1068
rect 115 1064 116 1068
rect 110 1063 116 1064
rect 222 1067 228 1068
rect 222 1063 223 1067
rect 227 1063 228 1067
rect 112 1035 114 1063
rect 222 1062 228 1063
rect 294 1067 300 1068
rect 294 1063 295 1067
rect 299 1063 300 1067
rect 294 1062 300 1063
rect 374 1067 380 1068
rect 374 1063 375 1067
rect 379 1063 380 1067
rect 374 1062 380 1063
rect 462 1067 468 1068
rect 462 1063 463 1067
rect 467 1063 468 1067
rect 462 1062 468 1063
rect 558 1067 564 1068
rect 558 1063 559 1067
rect 563 1063 564 1067
rect 558 1062 564 1063
rect 654 1067 660 1068
rect 654 1063 655 1067
rect 659 1063 660 1067
rect 654 1062 660 1063
rect 742 1067 748 1068
rect 742 1063 743 1067
rect 747 1063 748 1067
rect 742 1062 748 1063
rect 830 1067 836 1068
rect 830 1063 831 1067
rect 835 1063 836 1067
rect 830 1062 836 1063
rect 910 1067 916 1068
rect 910 1063 911 1067
rect 915 1063 916 1067
rect 910 1062 916 1063
rect 990 1067 996 1068
rect 990 1063 991 1067
rect 995 1063 996 1067
rect 990 1062 996 1063
rect 1070 1067 1076 1068
rect 1070 1063 1071 1067
rect 1075 1063 1076 1067
rect 1070 1062 1076 1063
rect 1158 1067 1164 1068
rect 1158 1063 1159 1067
rect 1163 1063 1164 1067
rect 1286 1064 1287 1068
rect 1291 1064 1292 1068
rect 1327 1065 1331 1066
rect 1367 1070 1371 1071
rect 1367 1065 1371 1066
rect 1399 1070 1403 1071
rect 1399 1065 1403 1066
rect 1455 1070 1459 1071
rect 1455 1065 1459 1066
rect 1463 1070 1467 1071
rect 1463 1065 1467 1066
rect 1535 1070 1539 1071
rect 1535 1065 1539 1066
rect 1575 1070 1579 1071
rect 1575 1065 1579 1066
rect 1607 1070 1611 1071
rect 1607 1065 1611 1066
rect 1687 1070 1691 1071
rect 1687 1065 1691 1066
rect 1695 1070 1699 1071
rect 1695 1065 1699 1066
rect 1767 1070 1771 1071
rect 1767 1065 1771 1066
rect 1815 1070 1819 1071
rect 1815 1065 1819 1066
rect 1847 1070 1851 1071
rect 1847 1065 1851 1066
rect 1927 1070 1931 1071
rect 1927 1065 1931 1066
rect 1999 1070 2003 1071
rect 1999 1065 2003 1066
rect 2039 1070 2043 1071
rect 2039 1065 2043 1066
rect 2071 1070 2075 1071
rect 2071 1065 2075 1066
rect 2151 1070 2155 1071
rect 2151 1065 2155 1066
rect 2231 1070 2235 1071
rect 2231 1065 2235 1066
rect 2255 1070 2259 1071
rect 2255 1065 2259 1066
rect 2367 1070 2371 1071
rect 2367 1065 2371 1066
rect 2455 1070 2459 1071
rect 2455 1065 2459 1066
rect 2503 1070 2507 1071
rect 2503 1065 2507 1066
rect 1286 1063 1292 1064
rect 1158 1062 1164 1063
rect 224 1035 226 1062
rect 296 1035 298 1062
rect 376 1035 378 1062
rect 464 1035 466 1062
rect 560 1035 562 1062
rect 656 1035 658 1062
rect 744 1035 746 1062
rect 832 1035 834 1062
rect 912 1035 914 1062
rect 992 1035 994 1062
rect 1072 1035 1074 1062
rect 1160 1035 1162 1062
rect 1288 1035 1290 1063
rect 1328 1045 1330 1065
rect 1368 1046 1370 1065
rect 1456 1046 1458 1065
rect 1576 1046 1578 1065
rect 1696 1046 1698 1065
rect 1816 1046 1818 1065
rect 1928 1046 1930 1065
rect 2040 1046 2042 1065
rect 2152 1046 2154 1065
rect 2256 1046 2258 1065
rect 2368 1046 2370 1065
rect 2456 1046 2458 1065
rect 1366 1045 1372 1046
rect 1326 1044 1332 1045
rect 1326 1040 1327 1044
rect 1331 1040 1332 1044
rect 1366 1041 1367 1045
rect 1371 1041 1372 1045
rect 1366 1040 1372 1041
rect 1454 1045 1460 1046
rect 1454 1041 1455 1045
rect 1459 1041 1460 1045
rect 1454 1040 1460 1041
rect 1574 1045 1580 1046
rect 1574 1041 1575 1045
rect 1579 1041 1580 1045
rect 1574 1040 1580 1041
rect 1694 1045 1700 1046
rect 1694 1041 1695 1045
rect 1699 1041 1700 1045
rect 1694 1040 1700 1041
rect 1814 1045 1820 1046
rect 1814 1041 1815 1045
rect 1819 1041 1820 1045
rect 1814 1040 1820 1041
rect 1926 1045 1932 1046
rect 1926 1041 1927 1045
rect 1931 1041 1932 1045
rect 1926 1040 1932 1041
rect 2038 1045 2044 1046
rect 2038 1041 2039 1045
rect 2043 1041 2044 1045
rect 2038 1040 2044 1041
rect 2150 1045 2156 1046
rect 2150 1041 2151 1045
rect 2155 1041 2156 1045
rect 2150 1040 2156 1041
rect 2254 1045 2260 1046
rect 2254 1041 2255 1045
rect 2259 1041 2260 1045
rect 2254 1040 2260 1041
rect 2366 1045 2372 1046
rect 2366 1041 2367 1045
rect 2371 1041 2372 1045
rect 2366 1040 2372 1041
rect 2454 1045 2460 1046
rect 2504 1045 2506 1065
rect 2454 1041 2455 1045
rect 2459 1041 2460 1045
rect 2454 1040 2460 1041
rect 2502 1044 2508 1045
rect 2502 1040 2503 1044
rect 2507 1040 2508 1044
rect 1326 1039 1332 1040
rect 2502 1039 2508 1040
rect 111 1034 115 1035
rect 111 1029 115 1030
rect 223 1034 227 1035
rect 223 1029 227 1030
rect 295 1034 299 1035
rect 295 1029 299 1030
rect 375 1034 379 1035
rect 375 1029 379 1030
rect 383 1034 387 1035
rect 383 1029 387 1030
rect 463 1034 467 1035
rect 463 1029 467 1030
rect 479 1034 483 1035
rect 479 1029 483 1030
rect 559 1034 563 1035
rect 559 1029 563 1030
rect 575 1034 579 1035
rect 575 1029 579 1030
rect 655 1034 659 1035
rect 655 1029 659 1030
rect 671 1034 675 1035
rect 671 1029 675 1030
rect 743 1034 747 1035
rect 743 1029 747 1030
rect 767 1034 771 1035
rect 767 1029 771 1030
rect 831 1034 835 1035
rect 831 1029 835 1030
rect 855 1034 859 1035
rect 855 1029 859 1030
rect 911 1034 915 1035
rect 911 1029 915 1030
rect 943 1034 947 1035
rect 943 1029 947 1030
rect 991 1034 995 1035
rect 991 1029 995 1030
rect 1023 1034 1027 1035
rect 1023 1029 1027 1030
rect 1071 1034 1075 1035
rect 1071 1029 1075 1030
rect 1103 1034 1107 1035
rect 1103 1029 1107 1030
rect 1159 1034 1163 1035
rect 1159 1029 1163 1030
rect 1183 1034 1187 1035
rect 1183 1029 1187 1030
rect 1239 1034 1243 1035
rect 1239 1029 1243 1030
rect 1287 1034 1291 1035
rect 1287 1029 1291 1030
rect 112 1009 114 1029
rect 296 1010 298 1029
rect 384 1010 386 1029
rect 480 1010 482 1029
rect 576 1010 578 1029
rect 672 1010 674 1029
rect 768 1010 770 1029
rect 856 1010 858 1029
rect 944 1010 946 1029
rect 1024 1010 1026 1029
rect 1104 1010 1106 1029
rect 1184 1010 1186 1029
rect 1240 1010 1242 1029
rect 294 1009 300 1010
rect 110 1008 116 1009
rect 110 1004 111 1008
rect 115 1004 116 1008
rect 294 1005 295 1009
rect 299 1005 300 1009
rect 294 1004 300 1005
rect 382 1009 388 1010
rect 382 1005 383 1009
rect 387 1005 388 1009
rect 382 1004 388 1005
rect 478 1009 484 1010
rect 478 1005 479 1009
rect 483 1005 484 1009
rect 478 1004 484 1005
rect 574 1009 580 1010
rect 574 1005 575 1009
rect 579 1005 580 1009
rect 574 1004 580 1005
rect 670 1009 676 1010
rect 670 1005 671 1009
rect 675 1005 676 1009
rect 670 1004 676 1005
rect 766 1009 772 1010
rect 766 1005 767 1009
rect 771 1005 772 1009
rect 766 1004 772 1005
rect 854 1009 860 1010
rect 854 1005 855 1009
rect 859 1005 860 1009
rect 854 1004 860 1005
rect 942 1009 948 1010
rect 942 1005 943 1009
rect 947 1005 948 1009
rect 942 1004 948 1005
rect 1022 1009 1028 1010
rect 1022 1005 1023 1009
rect 1027 1005 1028 1009
rect 1022 1004 1028 1005
rect 1102 1009 1108 1010
rect 1102 1005 1103 1009
rect 1107 1005 1108 1009
rect 1102 1004 1108 1005
rect 1182 1009 1188 1010
rect 1182 1005 1183 1009
rect 1187 1005 1188 1009
rect 1182 1004 1188 1005
rect 1238 1009 1244 1010
rect 1288 1009 1290 1029
rect 1326 1027 1332 1028
rect 1326 1023 1327 1027
rect 1331 1023 1332 1027
rect 2502 1027 2508 1028
rect 1326 1022 1332 1023
rect 1350 1024 1356 1025
rect 1328 1015 1330 1022
rect 1350 1020 1351 1024
rect 1355 1020 1356 1024
rect 1350 1019 1356 1020
rect 1438 1024 1444 1025
rect 1438 1020 1439 1024
rect 1443 1020 1444 1024
rect 1438 1019 1444 1020
rect 1558 1024 1564 1025
rect 1558 1020 1559 1024
rect 1563 1020 1564 1024
rect 1558 1019 1564 1020
rect 1678 1024 1684 1025
rect 1678 1020 1679 1024
rect 1683 1020 1684 1024
rect 1678 1019 1684 1020
rect 1798 1024 1804 1025
rect 1798 1020 1799 1024
rect 1803 1020 1804 1024
rect 1798 1019 1804 1020
rect 1910 1024 1916 1025
rect 1910 1020 1911 1024
rect 1915 1020 1916 1024
rect 1910 1019 1916 1020
rect 2022 1024 2028 1025
rect 2022 1020 2023 1024
rect 2027 1020 2028 1024
rect 2022 1019 2028 1020
rect 2134 1024 2140 1025
rect 2134 1020 2135 1024
rect 2139 1020 2140 1024
rect 2134 1019 2140 1020
rect 2238 1024 2244 1025
rect 2238 1020 2239 1024
rect 2243 1020 2244 1024
rect 2238 1019 2244 1020
rect 2350 1024 2356 1025
rect 2350 1020 2351 1024
rect 2355 1020 2356 1024
rect 2350 1019 2356 1020
rect 2438 1024 2444 1025
rect 2438 1020 2439 1024
rect 2443 1020 2444 1024
rect 2502 1023 2503 1027
rect 2507 1023 2508 1027
rect 2502 1022 2508 1023
rect 2438 1019 2444 1020
rect 1352 1015 1354 1019
rect 1440 1015 1442 1019
rect 1560 1015 1562 1019
rect 1680 1015 1682 1019
rect 1800 1015 1802 1019
rect 1912 1015 1914 1019
rect 2024 1015 2026 1019
rect 2136 1015 2138 1019
rect 2240 1015 2242 1019
rect 2352 1015 2354 1019
rect 2440 1015 2442 1019
rect 2504 1015 2506 1022
rect 1327 1014 1331 1015
rect 1327 1009 1331 1010
rect 1351 1014 1355 1015
rect 1351 1009 1355 1010
rect 1439 1014 1443 1015
rect 1439 1009 1443 1010
rect 1511 1014 1515 1015
rect 1511 1009 1515 1010
rect 1559 1014 1563 1015
rect 1559 1009 1563 1010
rect 1679 1014 1683 1015
rect 1679 1009 1683 1010
rect 1799 1014 1803 1015
rect 1799 1009 1803 1010
rect 1823 1014 1827 1015
rect 1823 1009 1827 1010
rect 1911 1014 1915 1015
rect 1911 1009 1915 1010
rect 1951 1014 1955 1015
rect 1951 1009 1955 1010
rect 2023 1014 2027 1015
rect 2023 1009 2027 1010
rect 2071 1014 2075 1015
rect 2071 1009 2075 1010
rect 2135 1014 2139 1015
rect 2135 1009 2139 1010
rect 2175 1014 2179 1015
rect 2175 1009 2179 1010
rect 2239 1014 2243 1015
rect 2239 1009 2243 1010
rect 2271 1014 2275 1015
rect 2271 1009 2275 1010
rect 2351 1014 2355 1015
rect 2351 1009 2355 1010
rect 2367 1014 2371 1015
rect 2367 1009 2371 1010
rect 2439 1014 2443 1015
rect 2439 1009 2443 1010
rect 2503 1014 2507 1015
rect 2503 1009 2507 1010
rect 1238 1005 1239 1009
rect 1243 1005 1244 1009
rect 1238 1004 1244 1005
rect 1286 1008 1292 1009
rect 1286 1004 1287 1008
rect 1291 1004 1292 1008
rect 1328 1006 1330 1009
rect 1350 1008 1356 1009
rect 110 1003 116 1004
rect 1286 1003 1292 1004
rect 1326 1005 1332 1006
rect 1326 1001 1327 1005
rect 1331 1001 1332 1005
rect 1350 1004 1351 1008
rect 1355 1004 1356 1008
rect 1350 1003 1356 1004
rect 1510 1008 1516 1009
rect 1510 1004 1511 1008
rect 1515 1004 1516 1008
rect 1510 1003 1516 1004
rect 1678 1008 1684 1009
rect 1678 1004 1679 1008
rect 1683 1004 1684 1008
rect 1678 1003 1684 1004
rect 1822 1008 1828 1009
rect 1822 1004 1823 1008
rect 1827 1004 1828 1008
rect 1822 1003 1828 1004
rect 1950 1008 1956 1009
rect 1950 1004 1951 1008
rect 1955 1004 1956 1008
rect 1950 1003 1956 1004
rect 2070 1008 2076 1009
rect 2070 1004 2071 1008
rect 2075 1004 2076 1008
rect 2070 1003 2076 1004
rect 2174 1008 2180 1009
rect 2174 1004 2175 1008
rect 2179 1004 2180 1008
rect 2174 1003 2180 1004
rect 2270 1008 2276 1009
rect 2270 1004 2271 1008
rect 2275 1004 2276 1008
rect 2270 1003 2276 1004
rect 2366 1008 2372 1009
rect 2366 1004 2367 1008
rect 2371 1004 2372 1008
rect 2366 1003 2372 1004
rect 2438 1008 2444 1009
rect 2438 1004 2439 1008
rect 2443 1004 2444 1008
rect 2504 1006 2506 1009
rect 2438 1003 2444 1004
rect 2502 1005 2508 1006
rect 1326 1000 1332 1001
rect 2502 1001 2503 1005
rect 2507 1001 2508 1005
rect 2502 1000 2508 1001
rect 110 991 116 992
rect 110 987 111 991
rect 115 987 116 991
rect 1286 991 1292 992
rect 110 986 116 987
rect 278 988 284 989
rect 112 983 114 986
rect 278 984 279 988
rect 283 984 284 988
rect 278 983 284 984
rect 366 988 372 989
rect 366 984 367 988
rect 371 984 372 988
rect 366 983 372 984
rect 462 988 468 989
rect 462 984 463 988
rect 467 984 468 988
rect 462 983 468 984
rect 558 988 564 989
rect 558 984 559 988
rect 563 984 564 988
rect 558 983 564 984
rect 654 988 660 989
rect 654 984 655 988
rect 659 984 660 988
rect 654 983 660 984
rect 750 988 756 989
rect 750 984 751 988
rect 755 984 756 988
rect 750 983 756 984
rect 838 988 844 989
rect 838 984 839 988
rect 843 984 844 988
rect 838 983 844 984
rect 926 988 932 989
rect 926 984 927 988
rect 931 984 932 988
rect 926 983 932 984
rect 1006 988 1012 989
rect 1006 984 1007 988
rect 1011 984 1012 988
rect 1006 983 1012 984
rect 1086 988 1092 989
rect 1086 984 1087 988
rect 1091 984 1092 988
rect 1086 983 1092 984
rect 1166 988 1172 989
rect 1166 984 1167 988
rect 1171 984 1172 988
rect 1166 983 1172 984
rect 1222 988 1228 989
rect 1222 984 1223 988
rect 1227 984 1228 988
rect 1286 987 1287 991
rect 1291 987 1292 991
rect 1286 986 1292 987
rect 1326 988 1332 989
rect 2502 988 2508 989
rect 1222 983 1228 984
rect 1288 983 1290 986
rect 1326 984 1327 988
rect 1331 984 1332 988
rect 1326 983 1332 984
rect 1366 987 1372 988
rect 1366 983 1367 987
rect 1371 983 1372 987
rect 111 982 115 983
rect 111 977 115 978
rect 271 982 275 983
rect 271 977 275 978
rect 279 982 283 983
rect 279 977 283 978
rect 359 982 363 983
rect 359 977 363 978
rect 367 982 371 983
rect 367 977 371 978
rect 455 982 459 983
rect 455 977 459 978
rect 463 982 467 983
rect 463 977 467 978
rect 551 982 555 983
rect 551 977 555 978
rect 559 982 563 983
rect 559 977 563 978
rect 655 982 659 983
rect 655 977 659 978
rect 751 982 755 983
rect 751 977 755 978
rect 839 982 843 983
rect 839 977 843 978
rect 927 982 931 983
rect 927 977 931 978
rect 1007 982 1011 983
rect 1007 977 1011 978
rect 1087 982 1091 983
rect 1087 977 1091 978
rect 1167 982 1171 983
rect 1167 977 1171 978
rect 1223 982 1227 983
rect 1223 977 1227 978
rect 1287 982 1291 983
rect 1287 977 1291 978
rect 112 974 114 977
rect 270 976 276 977
rect 110 973 116 974
rect 110 969 111 973
rect 115 969 116 973
rect 270 972 271 976
rect 275 972 276 976
rect 270 971 276 972
rect 358 976 364 977
rect 358 972 359 976
rect 363 972 364 976
rect 358 971 364 972
rect 454 976 460 977
rect 454 972 455 976
rect 459 972 460 976
rect 454 971 460 972
rect 550 976 556 977
rect 550 972 551 976
rect 555 972 556 976
rect 550 971 556 972
rect 654 976 660 977
rect 654 972 655 976
rect 659 972 660 976
rect 654 971 660 972
rect 750 976 756 977
rect 750 972 751 976
rect 755 972 756 976
rect 750 971 756 972
rect 838 976 844 977
rect 838 972 839 976
rect 843 972 844 976
rect 838 971 844 972
rect 926 976 932 977
rect 926 972 927 976
rect 931 972 932 976
rect 926 971 932 972
rect 1006 976 1012 977
rect 1006 972 1007 976
rect 1011 972 1012 976
rect 1006 971 1012 972
rect 1086 976 1092 977
rect 1086 972 1087 976
rect 1091 972 1092 976
rect 1086 971 1092 972
rect 1166 976 1172 977
rect 1166 972 1167 976
rect 1171 972 1172 976
rect 1166 971 1172 972
rect 1222 976 1228 977
rect 1222 972 1223 976
rect 1227 972 1228 976
rect 1288 974 1290 977
rect 1222 971 1228 972
rect 1286 973 1292 974
rect 110 968 116 969
rect 1286 969 1287 973
rect 1291 969 1292 973
rect 1286 968 1292 969
rect 110 956 116 957
rect 1286 956 1292 957
rect 110 952 111 956
rect 115 952 116 956
rect 110 951 116 952
rect 286 955 292 956
rect 286 951 287 955
rect 291 951 292 955
rect 112 923 114 951
rect 286 950 292 951
rect 374 955 380 956
rect 374 951 375 955
rect 379 951 380 955
rect 374 950 380 951
rect 470 955 476 956
rect 470 951 471 955
rect 475 951 476 955
rect 470 950 476 951
rect 566 955 572 956
rect 566 951 567 955
rect 571 951 572 955
rect 566 950 572 951
rect 670 955 676 956
rect 670 951 671 955
rect 675 951 676 955
rect 670 950 676 951
rect 766 955 772 956
rect 766 951 767 955
rect 771 951 772 955
rect 766 950 772 951
rect 854 955 860 956
rect 854 951 855 955
rect 859 951 860 955
rect 854 950 860 951
rect 942 955 948 956
rect 942 951 943 955
rect 947 951 948 955
rect 942 950 948 951
rect 1022 955 1028 956
rect 1022 951 1023 955
rect 1027 951 1028 955
rect 1022 950 1028 951
rect 1102 955 1108 956
rect 1102 951 1103 955
rect 1107 951 1108 955
rect 1102 950 1108 951
rect 1182 955 1188 956
rect 1182 951 1183 955
rect 1187 951 1188 955
rect 1182 950 1188 951
rect 1238 955 1244 956
rect 1238 951 1239 955
rect 1243 951 1244 955
rect 1286 952 1287 956
rect 1291 952 1292 956
rect 1286 951 1292 952
rect 1328 951 1330 983
rect 1366 982 1372 983
rect 1526 987 1532 988
rect 1526 983 1527 987
rect 1531 983 1532 987
rect 1526 982 1532 983
rect 1694 987 1700 988
rect 1694 983 1695 987
rect 1699 983 1700 987
rect 1694 982 1700 983
rect 1838 987 1844 988
rect 1838 983 1839 987
rect 1843 983 1844 987
rect 1838 982 1844 983
rect 1966 987 1972 988
rect 1966 983 1967 987
rect 1971 983 1972 987
rect 1966 982 1972 983
rect 2086 987 2092 988
rect 2086 983 2087 987
rect 2091 983 2092 987
rect 2086 982 2092 983
rect 2190 987 2196 988
rect 2190 983 2191 987
rect 2195 983 2196 987
rect 2190 982 2196 983
rect 2286 987 2292 988
rect 2286 983 2287 987
rect 2291 983 2292 987
rect 2286 982 2292 983
rect 2382 987 2388 988
rect 2382 983 2383 987
rect 2387 983 2388 987
rect 2382 982 2388 983
rect 2454 987 2460 988
rect 2454 983 2455 987
rect 2459 983 2460 987
rect 2502 984 2503 988
rect 2507 984 2508 988
rect 2502 983 2508 984
rect 2454 982 2460 983
rect 1368 951 1370 982
rect 1528 951 1530 982
rect 1696 951 1698 982
rect 1840 951 1842 982
rect 1968 951 1970 982
rect 2088 951 2090 982
rect 2192 951 2194 982
rect 2288 951 2290 982
rect 2384 951 2386 982
rect 2456 951 2458 982
rect 2504 951 2506 983
rect 1238 950 1244 951
rect 288 923 290 950
rect 376 923 378 950
rect 472 923 474 950
rect 568 923 570 950
rect 672 923 674 950
rect 768 923 770 950
rect 856 923 858 950
rect 944 923 946 950
rect 1024 923 1026 950
rect 1104 923 1106 950
rect 1184 923 1186 950
rect 1240 923 1242 950
rect 1288 923 1290 951
rect 1327 950 1331 951
rect 1327 945 1331 946
rect 1367 950 1371 951
rect 1367 945 1371 946
rect 1423 950 1427 951
rect 1423 945 1427 946
rect 1503 950 1507 951
rect 1503 945 1507 946
rect 1527 950 1531 951
rect 1527 945 1531 946
rect 1607 950 1611 951
rect 1607 945 1611 946
rect 1695 950 1699 951
rect 1695 945 1699 946
rect 1719 950 1723 951
rect 1719 945 1723 946
rect 1831 950 1835 951
rect 1831 945 1835 946
rect 1839 950 1843 951
rect 1839 945 1843 946
rect 1935 950 1939 951
rect 1935 945 1939 946
rect 1967 950 1971 951
rect 1967 945 1971 946
rect 2031 950 2035 951
rect 2031 945 2035 946
rect 2087 950 2091 951
rect 2087 945 2091 946
rect 2127 950 2131 951
rect 2127 945 2131 946
rect 2191 950 2195 951
rect 2191 945 2195 946
rect 2215 950 2219 951
rect 2215 945 2219 946
rect 2287 950 2291 951
rect 2287 945 2291 946
rect 2295 950 2299 951
rect 2295 945 2299 946
rect 2375 950 2379 951
rect 2375 945 2379 946
rect 2383 950 2387 951
rect 2383 945 2387 946
rect 2455 950 2459 951
rect 2455 945 2459 946
rect 2503 950 2507 951
rect 2503 945 2507 946
rect 1328 925 1330 945
rect 1368 926 1370 945
rect 1424 926 1426 945
rect 1504 926 1506 945
rect 1608 926 1610 945
rect 1720 926 1722 945
rect 1832 926 1834 945
rect 1936 926 1938 945
rect 2032 926 2034 945
rect 2128 926 2130 945
rect 2216 926 2218 945
rect 2296 926 2298 945
rect 2376 926 2378 945
rect 2456 926 2458 945
rect 1366 925 1372 926
rect 1326 924 1332 925
rect 111 922 115 923
rect 111 917 115 918
rect 271 922 275 923
rect 271 917 275 918
rect 287 922 291 923
rect 287 917 291 918
rect 343 922 347 923
rect 343 917 347 918
rect 375 922 379 923
rect 375 917 379 918
rect 423 922 427 923
rect 423 917 427 918
rect 471 922 475 923
rect 471 917 475 918
rect 519 922 523 923
rect 519 917 523 918
rect 567 922 571 923
rect 567 917 571 918
rect 615 922 619 923
rect 615 917 619 918
rect 671 922 675 923
rect 671 917 675 918
rect 711 922 715 923
rect 711 917 715 918
rect 767 922 771 923
rect 767 917 771 918
rect 807 922 811 923
rect 807 917 811 918
rect 855 922 859 923
rect 855 917 859 918
rect 903 922 907 923
rect 903 917 907 918
rect 943 922 947 923
rect 943 917 947 918
rect 991 922 995 923
rect 991 917 995 918
rect 1023 922 1027 923
rect 1023 917 1027 918
rect 1087 922 1091 923
rect 1087 917 1091 918
rect 1103 922 1107 923
rect 1103 917 1107 918
rect 1183 922 1187 923
rect 1183 917 1187 918
rect 1239 922 1243 923
rect 1239 917 1243 918
rect 1287 922 1291 923
rect 1326 920 1327 924
rect 1331 920 1332 924
rect 1366 921 1367 925
rect 1371 921 1372 925
rect 1366 920 1372 921
rect 1422 925 1428 926
rect 1422 921 1423 925
rect 1427 921 1428 925
rect 1422 920 1428 921
rect 1502 925 1508 926
rect 1502 921 1503 925
rect 1507 921 1508 925
rect 1502 920 1508 921
rect 1606 925 1612 926
rect 1606 921 1607 925
rect 1611 921 1612 925
rect 1606 920 1612 921
rect 1718 925 1724 926
rect 1718 921 1719 925
rect 1723 921 1724 925
rect 1718 920 1724 921
rect 1830 925 1836 926
rect 1830 921 1831 925
rect 1835 921 1836 925
rect 1830 920 1836 921
rect 1934 925 1940 926
rect 1934 921 1935 925
rect 1939 921 1940 925
rect 1934 920 1940 921
rect 2030 925 2036 926
rect 2030 921 2031 925
rect 2035 921 2036 925
rect 2030 920 2036 921
rect 2126 925 2132 926
rect 2126 921 2127 925
rect 2131 921 2132 925
rect 2126 920 2132 921
rect 2214 925 2220 926
rect 2214 921 2215 925
rect 2219 921 2220 925
rect 2214 920 2220 921
rect 2294 925 2300 926
rect 2294 921 2295 925
rect 2299 921 2300 925
rect 2294 920 2300 921
rect 2374 925 2380 926
rect 2374 921 2375 925
rect 2379 921 2380 925
rect 2374 920 2380 921
rect 2454 925 2460 926
rect 2504 925 2506 945
rect 2454 921 2455 925
rect 2459 921 2460 925
rect 2454 920 2460 921
rect 2502 924 2508 925
rect 2502 920 2503 924
rect 2507 920 2508 924
rect 1326 919 1332 920
rect 2502 919 2508 920
rect 1287 917 1291 918
rect 112 897 114 917
rect 272 898 274 917
rect 344 898 346 917
rect 424 898 426 917
rect 520 898 522 917
rect 616 898 618 917
rect 712 898 714 917
rect 808 898 810 917
rect 904 898 906 917
rect 992 898 994 917
rect 1088 898 1090 917
rect 1184 898 1186 917
rect 270 897 276 898
rect 110 896 116 897
rect 110 892 111 896
rect 115 892 116 896
rect 270 893 271 897
rect 275 893 276 897
rect 270 892 276 893
rect 342 897 348 898
rect 342 893 343 897
rect 347 893 348 897
rect 342 892 348 893
rect 422 897 428 898
rect 422 893 423 897
rect 427 893 428 897
rect 422 892 428 893
rect 518 897 524 898
rect 518 893 519 897
rect 523 893 524 897
rect 518 892 524 893
rect 614 897 620 898
rect 614 893 615 897
rect 619 893 620 897
rect 614 892 620 893
rect 710 897 716 898
rect 710 893 711 897
rect 715 893 716 897
rect 710 892 716 893
rect 806 897 812 898
rect 806 893 807 897
rect 811 893 812 897
rect 806 892 812 893
rect 902 897 908 898
rect 902 893 903 897
rect 907 893 908 897
rect 902 892 908 893
rect 990 897 996 898
rect 990 893 991 897
rect 995 893 996 897
rect 990 892 996 893
rect 1086 897 1092 898
rect 1086 893 1087 897
rect 1091 893 1092 897
rect 1086 892 1092 893
rect 1182 897 1188 898
rect 1288 897 1290 917
rect 1326 907 1332 908
rect 1326 903 1327 907
rect 1331 903 1332 907
rect 2502 907 2508 908
rect 1326 902 1332 903
rect 1350 904 1356 905
rect 1182 893 1183 897
rect 1187 893 1188 897
rect 1182 892 1188 893
rect 1286 896 1292 897
rect 1286 892 1287 896
rect 1291 892 1292 896
rect 1328 895 1330 902
rect 1350 900 1351 904
rect 1355 900 1356 904
rect 1350 899 1356 900
rect 1406 904 1412 905
rect 1406 900 1407 904
rect 1411 900 1412 904
rect 1406 899 1412 900
rect 1486 904 1492 905
rect 1486 900 1487 904
rect 1491 900 1492 904
rect 1486 899 1492 900
rect 1590 904 1596 905
rect 1590 900 1591 904
rect 1595 900 1596 904
rect 1590 899 1596 900
rect 1702 904 1708 905
rect 1702 900 1703 904
rect 1707 900 1708 904
rect 1702 899 1708 900
rect 1814 904 1820 905
rect 1814 900 1815 904
rect 1819 900 1820 904
rect 1814 899 1820 900
rect 1918 904 1924 905
rect 1918 900 1919 904
rect 1923 900 1924 904
rect 1918 899 1924 900
rect 2014 904 2020 905
rect 2014 900 2015 904
rect 2019 900 2020 904
rect 2014 899 2020 900
rect 2110 904 2116 905
rect 2110 900 2111 904
rect 2115 900 2116 904
rect 2110 899 2116 900
rect 2198 904 2204 905
rect 2198 900 2199 904
rect 2203 900 2204 904
rect 2198 899 2204 900
rect 2278 904 2284 905
rect 2278 900 2279 904
rect 2283 900 2284 904
rect 2278 899 2284 900
rect 2358 904 2364 905
rect 2358 900 2359 904
rect 2363 900 2364 904
rect 2358 899 2364 900
rect 2438 904 2444 905
rect 2438 900 2439 904
rect 2443 900 2444 904
rect 2502 903 2503 907
rect 2507 903 2508 907
rect 2502 902 2508 903
rect 2438 899 2444 900
rect 1352 895 1354 899
rect 1408 895 1410 899
rect 1488 895 1490 899
rect 1592 895 1594 899
rect 1704 895 1706 899
rect 1816 895 1818 899
rect 1920 895 1922 899
rect 2016 895 2018 899
rect 2112 895 2114 899
rect 2200 895 2202 899
rect 2280 895 2282 899
rect 2360 895 2362 899
rect 2440 895 2442 899
rect 2504 895 2506 902
rect 110 891 116 892
rect 1286 891 1292 892
rect 1327 894 1331 895
rect 1327 889 1331 890
rect 1351 894 1355 895
rect 1351 889 1355 890
rect 1407 894 1411 895
rect 1407 889 1411 890
rect 1431 894 1435 895
rect 1431 889 1435 890
rect 1487 894 1491 895
rect 1487 889 1491 890
rect 1551 894 1555 895
rect 1551 889 1555 890
rect 1591 894 1595 895
rect 1591 889 1595 890
rect 1623 894 1627 895
rect 1623 889 1627 890
rect 1703 894 1707 895
rect 1703 889 1707 890
rect 1791 894 1795 895
rect 1791 889 1795 890
rect 1815 894 1819 895
rect 1815 889 1819 890
rect 1895 894 1899 895
rect 1895 889 1899 890
rect 1919 894 1923 895
rect 1919 889 1923 890
rect 2015 894 2019 895
rect 2015 889 2019 890
rect 2111 894 2115 895
rect 2111 889 2115 890
rect 2143 894 2147 895
rect 2143 889 2147 890
rect 2199 894 2203 895
rect 2199 889 2203 890
rect 2279 894 2283 895
rect 2279 889 2283 890
rect 2359 894 2363 895
rect 2359 889 2363 890
rect 2423 894 2427 895
rect 2423 889 2427 890
rect 2439 894 2443 895
rect 2439 889 2443 890
rect 2503 894 2507 895
rect 2503 889 2507 890
rect 1328 886 1330 889
rect 1430 888 1436 889
rect 1326 885 1332 886
rect 1326 881 1327 885
rect 1331 881 1332 885
rect 1430 884 1431 888
rect 1435 884 1436 888
rect 1430 883 1436 884
rect 1486 888 1492 889
rect 1486 884 1487 888
rect 1491 884 1492 888
rect 1486 883 1492 884
rect 1550 888 1556 889
rect 1550 884 1551 888
rect 1555 884 1556 888
rect 1550 883 1556 884
rect 1622 888 1628 889
rect 1622 884 1623 888
rect 1627 884 1628 888
rect 1622 883 1628 884
rect 1702 888 1708 889
rect 1702 884 1703 888
rect 1707 884 1708 888
rect 1702 883 1708 884
rect 1790 888 1796 889
rect 1790 884 1791 888
rect 1795 884 1796 888
rect 1790 883 1796 884
rect 1894 888 1900 889
rect 1894 884 1895 888
rect 1899 884 1900 888
rect 1894 883 1900 884
rect 2014 888 2020 889
rect 2014 884 2015 888
rect 2019 884 2020 888
rect 2014 883 2020 884
rect 2142 888 2148 889
rect 2142 884 2143 888
rect 2147 884 2148 888
rect 2142 883 2148 884
rect 2278 888 2284 889
rect 2278 884 2279 888
rect 2283 884 2284 888
rect 2278 883 2284 884
rect 2422 888 2428 889
rect 2422 884 2423 888
rect 2427 884 2428 888
rect 2504 886 2506 889
rect 2422 883 2428 884
rect 2502 885 2508 886
rect 1326 880 1332 881
rect 2502 881 2503 885
rect 2507 881 2508 885
rect 2502 880 2508 881
rect 110 879 116 880
rect 110 875 111 879
rect 115 875 116 879
rect 1286 879 1292 880
rect 110 874 116 875
rect 254 876 260 877
rect 112 867 114 874
rect 254 872 255 876
rect 259 872 260 876
rect 254 871 260 872
rect 326 876 332 877
rect 326 872 327 876
rect 331 872 332 876
rect 326 871 332 872
rect 406 876 412 877
rect 406 872 407 876
rect 411 872 412 876
rect 406 871 412 872
rect 502 876 508 877
rect 502 872 503 876
rect 507 872 508 876
rect 502 871 508 872
rect 598 876 604 877
rect 598 872 599 876
rect 603 872 604 876
rect 598 871 604 872
rect 694 876 700 877
rect 694 872 695 876
rect 699 872 700 876
rect 694 871 700 872
rect 790 876 796 877
rect 790 872 791 876
rect 795 872 796 876
rect 790 871 796 872
rect 886 876 892 877
rect 886 872 887 876
rect 891 872 892 876
rect 886 871 892 872
rect 974 876 980 877
rect 974 872 975 876
rect 979 872 980 876
rect 974 871 980 872
rect 1070 876 1076 877
rect 1070 872 1071 876
rect 1075 872 1076 876
rect 1070 871 1076 872
rect 1166 876 1172 877
rect 1166 872 1167 876
rect 1171 872 1172 876
rect 1286 875 1287 879
rect 1291 875 1292 879
rect 1286 874 1292 875
rect 1166 871 1172 872
rect 256 867 258 871
rect 328 867 330 871
rect 408 867 410 871
rect 504 867 506 871
rect 600 867 602 871
rect 696 867 698 871
rect 792 867 794 871
rect 888 867 890 871
rect 976 867 978 871
rect 1072 867 1074 871
rect 1168 867 1170 871
rect 1288 867 1290 874
rect 1326 868 1332 869
rect 2502 868 2508 869
rect 111 866 115 867
rect 111 861 115 862
rect 247 866 251 867
rect 247 861 251 862
rect 255 866 259 867
rect 255 861 259 862
rect 311 866 315 867
rect 311 861 315 862
rect 327 866 331 867
rect 327 861 331 862
rect 375 866 379 867
rect 375 861 379 862
rect 407 866 411 867
rect 407 861 411 862
rect 439 866 443 867
rect 439 861 443 862
rect 503 866 507 867
rect 503 861 507 862
rect 567 866 571 867
rect 567 861 571 862
rect 599 866 603 867
rect 599 861 603 862
rect 631 866 635 867
rect 631 861 635 862
rect 695 866 699 867
rect 695 861 699 862
rect 759 866 763 867
rect 759 861 763 862
rect 791 866 795 867
rect 791 861 795 862
rect 831 866 835 867
rect 831 861 835 862
rect 887 866 891 867
rect 887 861 891 862
rect 903 866 907 867
rect 903 861 907 862
rect 975 866 979 867
rect 975 861 979 862
rect 1071 866 1075 867
rect 1071 861 1075 862
rect 1167 866 1171 867
rect 1167 861 1171 862
rect 1287 866 1291 867
rect 1326 864 1327 868
rect 1331 864 1332 868
rect 1326 863 1332 864
rect 1446 867 1452 868
rect 1446 863 1447 867
rect 1451 863 1452 867
rect 1287 861 1291 862
rect 112 858 114 861
rect 246 860 252 861
rect 110 857 116 858
rect 110 853 111 857
rect 115 853 116 857
rect 246 856 247 860
rect 251 856 252 860
rect 246 855 252 856
rect 310 860 316 861
rect 310 856 311 860
rect 315 856 316 860
rect 310 855 316 856
rect 374 860 380 861
rect 374 856 375 860
rect 379 856 380 860
rect 374 855 380 856
rect 438 860 444 861
rect 438 856 439 860
rect 443 856 444 860
rect 438 855 444 856
rect 502 860 508 861
rect 502 856 503 860
rect 507 856 508 860
rect 502 855 508 856
rect 566 860 572 861
rect 566 856 567 860
rect 571 856 572 860
rect 566 855 572 856
rect 630 860 636 861
rect 630 856 631 860
rect 635 856 636 860
rect 630 855 636 856
rect 694 860 700 861
rect 694 856 695 860
rect 699 856 700 860
rect 694 855 700 856
rect 758 860 764 861
rect 758 856 759 860
rect 763 856 764 860
rect 758 855 764 856
rect 830 860 836 861
rect 830 856 831 860
rect 835 856 836 860
rect 830 855 836 856
rect 902 860 908 861
rect 902 856 903 860
rect 907 856 908 860
rect 1288 858 1290 861
rect 902 855 908 856
rect 1286 857 1292 858
rect 110 852 116 853
rect 1286 853 1287 857
rect 1291 853 1292 857
rect 1286 852 1292 853
rect 110 840 116 841
rect 1286 840 1292 841
rect 110 836 111 840
rect 115 836 116 840
rect 110 835 116 836
rect 262 839 268 840
rect 262 835 263 839
rect 267 835 268 839
rect 112 811 114 835
rect 262 834 268 835
rect 326 839 332 840
rect 326 835 327 839
rect 331 835 332 839
rect 326 834 332 835
rect 390 839 396 840
rect 390 835 391 839
rect 395 835 396 839
rect 390 834 396 835
rect 454 839 460 840
rect 454 835 455 839
rect 459 835 460 839
rect 454 834 460 835
rect 518 839 524 840
rect 518 835 519 839
rect 523 835 524 839
rect 518 834 524 835
rect 582 839 588 840
rect 582 835 583 839
rect 587 835 588 839
rect 582 834 588 835
rect 646 839 652 840
rect 646 835 647 839
rect 651 835 652 839
rect 646 834 652 835
rect 710 839 716 840
rect 710 835 711 839
rect 715 835 716 839
rect 710 834 716 835
rect 774 839 780 840
rect 774 835 775 839
rect 779 835 780 839
rect 774 834 780 835
rect 846 839 852 840
rect 846 835 847 839
rect 851 835 852 839
rect 846 834 852 835
rect 918 839 924 840
rect 918 835 919 839
rect 923 835 924 839
rect 1286 836 1287 840
rect 1291 836 1292 840
rect 1328 839 1330 863
rect 1446 862 1452 863
rect 1502 867 1508 868
rect 1502 863 1503 867
rect 1507 863 1508 867
rect 1502 862 1508 863
rect 1566 867 1572 868
rect 1566 863 1567 867
rect 1571 863 1572 867
rect 1566 862 1572 863
rect 1638 867 1644 868
rect 1638 863 1639 867
rect 1643 863 1644 867
rect 1638 862 1644 863
rect 1718 867 1724 868
rect 1718 863 1719 867
rect 1723 863 1724 867
rect 1718 862 1724 863
rect 1806 867 1812 868
rect 1806 863 1807 867
rect 1811 863 1812 867
rect 1806 862 1812 863
rect 1910 867 1916 868
rect 1910 863 1911 867
rect 1915 863 1916 867
rect 1910 862 1916 863
rect 2030 867 2036 868
rect 2030 863 2031 867
rect 2035 863 2036 867
rect 2030 862 2036 863
rect 2158 867 2164 868
rect 2158 863 2159 867
rect 2163 863 2164 867
rect 2158 862 2164 863
rect 2294 867 2300 868
rect 2294 863 2295 867
rect 2299 863 2300 867
rect 2294 862 2300 863
rect 2438 867 2444 868
rect 2438 863 2439 867
rect 2443 863 2444 867
rect 2502 864 2503 868
rect 2507 864 2508 868
rect 2502 863 2508 864
rect 2438 862 2444 863
rect 1448 839 1450 862
rect 1504 839 1506 862
rect 1568 839 1570 862
rect 1640 839 1642 862
rect 1720 839 1722 862
rect 1808 839 1810 862
rect 1912 839 1914 862
rect 2032 839 2034 862
rect 2160 839 2162 862
rect 2296 839 2298 862
rect 2440 839 2442 862
rect 2504 839 2506 863
rect 1286 835 1292 836
rect 1327 838 1331 839
rect 918 834 924 835
rect 264 811 266 834
rect 328 811 330 834
rect 392 811 394 834
rect 456 811 458 834
rect 520 811 522 834
rect 584 811 586 834
rect 648 811 650 834
rect 712 811 714 834
rect 776 811 778 834
rect 848 811 850 834
rect 920 811 922 834
rect 1288 811 1290 835
rect 1327 833 1331 834
rect 1447 838 1451 839
rect 1447 833 1451 834
rect 1503 838 1507 839
rect 1503 833 1507 834
rect 1567 838 1571 839
rect 1567 833 1571 834
rect 1591 838 1595 839
rect 1591 833 1595 834
rect 1639 838 1643 839
rect 1639 833 1643 834
rect 1647 838 1651 839
rect 1647 833 1651 834
rect 1703 838 1707 839
rect 1703 833 1707 834
rect 1719 838 1723 839
rect 1719 833 1723 834
rect 1767 838 1771 839
rect 1767 833 1771 834
rect 1807 838 1811 839
rect 1807 833 1811 834
rect 1847 838 1851 839
rect 1847 833 1851 834
rect 1911 838 1915 839
rect 1911 833 1915 834
rect 1927 838 1931 839
rect 1927 833 1931 834
rect 2015 838 2019 839
rect 2015 833 2019 834
rect 2031 838 2035 839
rect 2031 833 2035 834
rect 2103 838 2107 839
rect 2103 833 2107 834
rect 2159 838 2163 839
rect 2159 833 2163 834
rect 2191 838 2195 839
rect 2191 833 2195 834
rect 2287 838 2291 839
rect 2287 833 2291 834
rect 2295 838 2299 839
rect 2295 833 2299 834
rect 2383 838 2387 839
rect 2383 833 2387 834
rect 2439 838 2443 839
rect 2439 833 2443 834
rect 2455 838 2459 839
rect 2455 833 2459 834
rect 2503 838 2507 839
rect 2503 833 2507 834
rect 1328 813 1330 833
rect 1592 814 1594 833
rect 1648 814 1650 833
rect 1704 814 1706 833
rect 1768 814 1770 833
rect 1848 814 1850 833
rect 1928 814 1930 833
rect 2016 814 2018 833
rect 2104 814 2106 833
rect 2192 814 2194 833
rect 2288 814 2290 833
rect 2384 814 2386 833
rect 2456 814 2458 833
rect 1590 813 1596 814
rect 1326 812 1332 813
rect 111 810 115 811
rect 111 805 115 806
rect 215 810 219 811
rect 215 805 219 806
rect 263 810 267 811
rect 263 805 267 806
rect 303 810 307 811
rect 303 805 307 806
rect 327 810 331 811
rect 327 805 331 806
rect 391 810 395 811
rect 391 805 395 806
rect 455 810 459 811
rect 455 805 459 806
rect 479 810 483 811
rect 479 805 483 806
rect 519 810 523 811
rect 519 805 523 806
rect 559 810 563 811
rect 559 805 563 806
rect 583 810 587 811
rect 583 805 587 806
rect 631 810 635 811
rect 631 805 635 806
rect 647 810 651 811
rect 647 805 651 806
rect 703 810 707 811
rect 703 805 707 806
rect 711 810 715 811
rect 711 805 715 806
rect 767 810 771 811
rect 767 805 771 806
rect 775 810 779 811
rect 775 805 779 806
rect 831 810 835 811
rect 831 805 835 806
rect 847 810 851 811
rect 847 805 851 806
rect 895 810 899 811
rect 895 805 899 806
rect 919 810 923 811
rect 919 805 923 806
rect 967 810 971 811
rect 967 805 971 806
rect 1039 810 1043 811
rect 1039 805 1043 806
rect 1287 810 1291 811
rect 1326 808 1327 812
rect 1331 808 1332 812
rect 1590 809 1591 813
rect 1595 809 1596 813
rect 1590 808 1596 809
rect 1646 813 1652 814
rect 1646 809 1647 813
rect 1651 809 1652 813
rect 1646 808 1652 809
rect 1702 813 1708 814
rect 1702 809 1703 813
rect 1707 809 1708 813
rect 1702 808 1708 809
rect 1766 813 1772 814
rect 1766 809 1767 813
rect 1771 809 1772 813
rect 1766 808 1772 809
rect 1846 813 1852 814
rect 1846 809 1847 813
rect 1851 809 1852 813
rect 1846 808 1852 809
rect 1926 813 1932 814
rect 1926 809 1927 813
rect 1931 809 1932 813
rect 1926 808 1932 809
rect 2014 813 2020 814
rect 2014 809 2015 813
rect 2019 809 2020 813
rect 2014 808 2020 809
rect 2102 813 2108 814
rect 2102 809 2103 813
rect 2107 809 2108 813
rect 2102 808 2108 809
rect 2190 813 2196 814
rect 2190 809 2191 813
rect 2195 809 2196 813
rect 2190 808 2196 809
rect 2286 813 2292 814
rect 2286 809 2287 813
rect 2291 809 2292 813
rect 2286 808 2292 809
rect 2382 813 2388 814
rect 2382 809 2383 813
rect 2387 809 2388 813
rect 2382 808 2388 809
rect 2454 813 2460 814
rect 2504 813 2506 833
rect 2454 809 2455 813
rect 2459 809 2460 813
rect 2454 808 2460 809
rect 2502 812 2508 813
rect 2502 808 2503 812
rect 2507 808 2508 812
rect 1326 807 1332 808
rect 2502 807 2508 808
rect 1287 805 1291 806
rect 112 785 114 805
rect 216 786 218 805
rect 304 786 306 805
rect 392 786 394 805
rect 480 786 482 805
rect 560 786 562 805
rect 632 786 634 805
rect 704 786 706 805
rect 768 786 770 805
rect 832 786 834 805
rect 896 786 898 805
rect 968 786 970 805
rect 1040 786 1042 805
rect 214 785 220 786
rect 110 784 116 785
rect 110 780 111 784
rect 115 780 116 784
rect 214 781 215 785
rect 219 781 220 785
rect 214 780 220 781
rect 302 785 308 786
rect 302 781 303 785
rect 307 781 308 785
rect 302 780 308 781
rect 390 785 396 786
rect 390 781 391 785
rect 395 781 396 785
rect 390 780 396 781
rect 478 785 484 786
rect 478 781 479 785
rect 483 781 484 785
rect 478 780 484 781
rect 558 785 564 786
rect 558 781 559 785
rect 563 781 564 785
rect 558 780 564 781
rect 630 785 636 786
rect 630 781 631 785
rect 635 781 636 785
rect 630 780 636 781
rect 702 785 708 786
rect 702 781 703 785
rect 707 781 708 785
rect 702 780 708 781
rect 766 785 772 786
rect 766 781 767 785
rect 771 781 772 785
rect 766 780 772 781
rect 830 785 836 786
rect 830 781 831 785
rect 835 781 836 785
rect 830 780 836 781
rect 894 785 900 786
rect 894 781 895 785
rect 899 781 900 785
rect 894 780 900 781
rect 966 785 972 786
rect 966 781 967 785
rect 971 781 972 785
rect 966 780 972 781
rect 1038 785 1044 786
rect 1288 785 1290 805
rect 1326 795 1332 796
rect 1326 791 1327 795
rect 1331 791 1332 795
rect 2502 795 2508 796
rect 1326 790 1332 791
rect 1574 792 1580 793
rect 1038 781 1039 785
rect 1043 781 1044 785
rect 1038 780 1044 781
rect 1286 784 1292 785
rect 1286 780 1287 784
rect 1291 780 1292 784
rect 1328 783 1330 790
rect 1574 788 1575 792
rect 1579 788 1580 792
rect 1574 787 1580 788
rect 1630 792 1636 793
rect 1630 788 1631 792
rect 1635 788 1636 792
rect 1630 787 1636 788
rect 1686 792 1692 793
rect 1686 788 1687 792
rect 1691 788 1692 792
rect 1686 787 1692 788
rect 1750 792 1756 793
rect 1750 788 1751 792
rect 1755 788 1756 792
rect 1750 787 1756 788
rect 1830 792 1836 793
rect 1830 788 1831 792
rect 1835 788 1836 792
rect 1830 787 1836 788
rect 1910 792 1916 793
rect 1910 788 1911 792
rect 1915 788 1916 792
rect 1910 787 1916 788
rect 1998 792 2004 793
rect 1998 788 1999 792
rect 2003 788 2004 792
rect 1998 787 2004 788
rect 2086 792 2092 793
rect 2086 788 2087 792
rect 2091 788 2092 792
rect 2086 787 2092 788
rect 2174 792 2180 793
rect 2174 788 2175 792
rect 2179 788 2180 792
rect 2174 787 2180 788
rect 2270 792 2276 793
rect 2270 788 2271 792
rect 2275 788 2276 792
rect 2270 787 2276 788
rect 2366 792 2372 793
rect 2366 788 2367 792
rect 2371 788 2372 792
rect 2366 787 2372 788
rect 2438 792 2444 793
rect 2438 788 2439 792
rect 2443 788 2444 792
rect 2502 791 2503 795
rect 2507 791 2508 795
rect 2502 790 2508 791
rect 2438 787 2444 788
rect 1576 783 1578 787
rect 1632 783 1634 787
rect 1688 783 1690 787
rect 1752 783 1754 787
rect 1832 783 1834 787
rect 1912 783 1914 787
rect 2000 783 2002 787
rect 2088 783 2090 787
rect 2176 783 2178 787
rect 2272 783 2274 787
rect 2368 783 2370 787
rect 2440 783 2442 787
rect 2504 783 2506 790
rect 110 779 116 780
rect 1286 779 1292 780
rect 1327 782 1331 783
rect 1327 777 1331 778
rect 1567 782 1571 783
rect 1567 777 1571 778
rect 1575 782 1579 783
rect 1575 777 1579 778
rect 1623 782 1627 783
rect 1623 777 1627 778
rect 1631 782 1635 783
rect 1631 777 1635 778
rect 1687 782 1691 783
rect 1687 777 1691 778
rect 1751 782 1755 783
rect 1751 777 1755 778
rect 1759 782 1763 783
rect 1759 777 1763 778
rect 1831 782 1835 783
rect 1831 777 1835 778
rect 1911 782 1915 783
rect 1911 777 1915 778
rect 1919 782 1923 783
rect 1919 777 1923 778
rect 1999 782 2003 783
rect 1999 777 2003 778
rect 2015 782 2019 783
rect 2015 777 2019 778
rect 2087 782 2091 783
rect 2087 777 2091 778
rect 2119 782 2123 783
rect 2119 777 2123 778
rect 2175 782 2179 783
rect 2175 777 2179 778
rect 2231 782 2235 783
rect 2231 777 2235 778
rect 2271 782 2275 783
rect 2271 777 2275 778
rect 2343 782 2347 783
rect 2343 777 2347 778
rect 2367 782 2371 783
rect 2367 777 2371 778
rect 2439 782 2443 783
rect 2439 777 2443 778
rect 2503 782 2507 783
rect 2503 777 2507 778
rect 1328 774 1330 777
rect 1566 776 1572 777
rect 1326 773 1332 774
rect 1326 769 1327 773
rect 1331 769 1332 773
rect 1566 772 1567 776
rect 1571 772 1572 776
rect 1566 771 1572 772
rect 1622 776 1628 777
rect 1622 772 1623 776
rect 1627 772 1628 776
rect 1622 771 1628 772
rect 1686 776 1692 777
rect 1686 772 1687 776
rect 1691 772 1692 776
rect 1686 771 1692 772
rect 1758 776 1764 777
rect 1758 772 1759 776
rect 1763 772 1764 776
rect 1758 771 1764 772
rect 1830 776 1836 777
rect 1830 772 1831 776
rect 1835 772 1836 776
rect 1830 771 1836 772
rect 1918 776 1924 777
rect 1918 772 1919 776
rect 1923 772 1924 776
rect 1918 771 1924 772
rect 2014 776 2020 777
rect 2014 772 2015 776
rect 2019 772 2020 776
rect 2014 771 2020 772
rect 2118 776 2124 777
rect 2118 772 2119 776
rect 2123 772 2124 776
rect 2118 771 2124 772
rect 2230 776 2236 777
rect 2230 772 2231 776
rect 2235 772 2236 776
rect 2230 771 2236 772
rect 2342 776 2348 777
rect 2342 772 2343 776
rect 2347 772 2348 776
rect 2342 771 2348 772
rect 2438 776 2444 777
rect 2438 772 2439 776
rect 2443 772 2444 776
rect 2504 774 2506 777
rect 2438 771 2444 772
rect 2502 773 2508 774
rect 1326 768 1332 769
rect 2502 769 2503 773
rect 2507 769 2508 773
rect 2502 768 2508 769
rect 110 767 116 768
rect 110 763 111 767
rect 115 763 116 767
rect 1286 767 1292 768
rect 110 762 116 763
rect 198 764 204 765
rect 112 759 114 762
rect 198 760 199 764
rect 203 760 204 764
rect 198 759 204 760
rect 286 764 292 765
rect 286 760 287 764
rect 291 760 292 764
rect 286 759 292 760
rect 374 764 380 765
rect 374 760 375 764
rect 379 760 380 764
rect 374 759 380 760
rect 462 764 468 765
rect 462 760 463 764
rect 467 760 468 764
rect 462 759 468 760
rect 542 764 548 765
rect 542 760 543 764
rect 547 760 548 764
rect 542 759 548 760
rect 614 764 620 765
rect 614 760 615 764
rect 619 760 620 764
rect 614 759 620 760
rect 686 764 692 765
rect 686 760 687 764
rect 691 760 692 764
rect 686 759 692 760
rect 750 764 756 765
rect 750 760 751 764
rect 755 760 756 764
rect 750 759 756 760
rect 814 764 820 765
rect 814 760 815 764
rect 819 760 820 764
rect 814 759 820 760
rect 878 764 884 765
rect 878 760 879 764
rect 883 760 884 764
rect 878 759 884 760
rect 950 764 956 765
rect 950 760 951 764
rect 955 760 956 764
rect 950 759 956 760
rect 1022 764 1028 765
rect 1022 760 1023 764
rect 1027 760 1028 764
rect 1286 763 1287 767
rect 1291 763 1292 767
rect 1286 762 1292 763
rect 1022 759 1028 760
rect 1288 759 1290 762
rect 111 758 115 759
rect 111 753 115 754
rect 135 758 139 759
rect 135 753 139 754
rect 199 758 203 759
rect 199 753 203 754
rect 255 758 259 759
rect 255 753 259 754
rect 287 758 291 759
rect 287 753 291 754
rect 375 758 379 759
rect 375 753 379 754
rect 391 758 395 759
rect 391 753 395 754
rect 463 758 467 759
rect 463 753 467 754
rect 519 758 523 759
rect 519 753 523 754
rect 543 758 547 759
rect 543 753 547 754
rect 615 758 619 759
rect 615 753 619 754
rect 647 758 651 759
rect 647 753 651 754
rect 687 758 691 759
rect 687 753 691 754
rect 751 758 755 759
rect 751 753 755 754
rect 775 758 779 759
rect 775 753 779 754
rect 815 758 819 759
rect 815 753 819 754
rect 879 758 883 759
rect 879 753 883 754
rect 903 758 907 759
rect 903 753 907 754
rect 951 758 955 759
rect 951 753 955 754
rect 1023 758 1027 759
rect 1023 753 1027 754
rect 1039 758 1043 759
rect 1039 753 1043 754
rect 1287 758 1291 759
rect 1287 753 1291 754
rect 1326 756 1332 757
rect 2502 756 2508 757
rect 112 750 114 753
rect 134 752 140 753
rect 110 749 116 750
rect 110 745 111 749
rect 115 745 116 749
rect 134 748 135 752
rect 139 748 140 752
rect 134 747 140 748
rect 254 752 260 753
rect 254 748 255 752
rect 259 748 260 752
rect 254 747 260 748
rect 390 752 396 753
rect 390 748 391 752
rect 395 748 396 752
rect 390 747 396 748
rect 518 752 524 753
rect 518 748 519 752
rect 523 748 524 752
rect 518 747 524 748
rect 646 752 652 753
rect 646 748 647 752
rect 651 748 652 752
rect 646 747 652 748
rect 774 752 780 753
rect 774 748 775 752
rect 779 748 780 752
rect 774 747 780 748
rect 902 752 908 753
rect 902 748 903 752
rect 907 748 908 752
rect 902 747 908 748
rect 1038 752 1044 753
rect 1038 748 1039 752
rect 1043 748 1044 752
rect 1288 750 1290 753
rect 1326 752 1327 756
rect 1331 752 1332 756
rect 1326 751 1332 752
rect 1582 755 1588 756
rect 1582 751 1583 755
rect 1587 751 1588 755
rect 1038 747 1044 748
rect 1286 749 1292 750
rect 110 744 116 745
rect 1286 745 1287 749
rect 1291 745 1292 749
rect 1286 744 1292 745
rect 110 732 116 733
rect 1286 732 1292 733
rect 110 728 111 732
rect 115 728 116 732
rect 110 727 116 728
rect 150 731 156 732
rect 150 727 151 731
rect 155 727 156 731
rect 112 707 114 727
rect 150 726 156 727
rect 270 731 276 732
rect 270 727 271 731
rect 275 727 276 731
rect 270 726 276 727
rect 406 731 412 732
rect 406 727 407 731
rect 411 727 412 731
rect 406 726 412 727
rect 534 731 540 732
rect 534 727 535 731
rect 539 727 540 731
rect 534 726 540 727
rect 662 731 668 732
rect 662 727 663 731
rect 667 727 668 731
rect 662 726 668 727
rect 790 731 796 732
rect 790 727 791 731
rect 795 727 796 731
rect 790 726 796 727
rect 918 731 924 732
rect 918 727 919 731
rect 923 727 924 731
rect 918 726 924 727
rect 1054 731 1060 732
rect 1054 727 1055 731
rect 1059 727 1060 731
rect 1286 728 1287 732
rect 1291 728 1292 732
rect 1328 731 1330 751
rect 1582 750 1588 751
rect 1638 755 1644 756
rect 1638 751 1639 755
rect 1643 751 1644 755
rect 1638 750 1644 751
rect 1702 755 1708 756
rect 1702 751 1703 755
rect 1707 751 1708 755
rect 1702 750 1708 751
rect 1774 755 1780 756
rect 1774 751 1775 755
rect 1779 751 1780 755
rect 1774 750 1780 751
rect 1846 755 1852 756
rect 1846 751 1847 755
rect 1851 751 1852 755
rect 1846 750 1852 751
rect 1934 755 1940 756
rect 1934 751 1935 755
rect 1939 751 1940 755
rect 1934 750 1940 751
rect 2030 755 2036 756
rect 2030 751 2031 755
rect 2035 751 2036 755
rect 2030 750 2036 751
rect 2134 755 2140 756
rect 2134 751 2135 755
rect 2139 751 2140 755
rect 2134 750 2140 751
rect 2246 755 2252 756
rect 2246 751 2247 755
rect 2251 751 2252 755
rect 2246 750 2252 751
rect 2358 755 2364 756
rect 2358 751 2359 755
rect 2363 751 2364 755
rect 2358 750 2364 751
rect 2454 755 2460 756
rect 2454 751 2455 755
rect 2459 751 2460 755
rect 2502 752 2503 756
rect 2507 752 2508 756
rect 2502 751 2508 752
rect 2454 750 2460 751
rect 1584 731 1586 750
rect 1640 731 1642 750
rect 1704 731 1706 750
rect 1776 731 1778 750
rect 1848 731 1850 750
rect 1936 731 1938 750
rect 2032 731 2034 750
rect 2136 731 2138 750
rect 2248 731 2250 750
rect 2360 731 2362 750
rect 2456 731 2458 750
rect 2504 731 2506 751
rect 1286 727 1292 728
rect 1327 730 1331 731
rect 1054 726 1060 727
rect 152 707 154 726
rect 272 707 274 726
rect 408 707 410 726
rect 536 707 538 726
rect 664 707 666 726
rect 792 707 794 726
rect 920 707 922 726
rect 1056 707 1058 726
rect 1288 707 1290 727
rect 1327 725 1331 726
rect 1367 730 1371 731
rect 1367 725 1371 726
rect 1431 730 1435 731
rect 1431 725 1435 726
rect 1527 730 1531 731
rect 1527 725 1531 726
rect 1583 730 1587 731
rect 1583 725 1587 726
rect 1631 730 1635 731
rect 1631 725 1635 726
rect 1639 730 1643 731
rect 1639 725 1643 726
rect 1703 730 1707 731
rect 1703 725 1707 726
rect 1735 730 1739 731
rect 1735 725 1739 726
rect 1775 730 1779 731
rect 1775 725 1779 726
rect 1839 730 1843 731
rect 1839 725 1843 726
rect 1847 730 1851 731
rect 1847 725 1851 726
rect 1935 730 1939 731
rect 1935 725 1939 726
rect 1943 730 1947 731
rect 1943 725 1947 726
rect 2031 730 2035 731
rect 2031 725 2035 726
rect 2047 730 2051 731
rect 2047 725 2051 726
rect 2135 730 2139 731
rect 2135 725 2139 726
rect 2151 730 2155 731
rect 2151 725 2155 726
rect 2247 730 2251 731
rect 2247 725 2251 726
rect 2255 730 2259 731
rect 2255 725 2259 726
rect 2359 730 2363 731
rect 2359 725 2363 726
rect 2367 730 2371 731
rect 2367 725 2371 726
rect 2455 730 2459 731
rect 2455 725 2459 726
rect 2503 730 2507 731
rect 2503 725 2507 726
rect 111 706 115 707
rect 111 701 115 702
rect 151 706 155 707
rect 151 701 155 702
rect 207 706 211 707
rect 207 701 211 702
rect 271 706 275 707
rect 271 701 275 702
rect 295 706 299 707
rect 295 701 299 702
rect 391 706 395 707
rect 391 701 395 702
rect 407 706 411 707
rect 407 701 411 702
rect 503 706 507 707
rect 503 701 507 702
rect 535 706 539 707
rect 535 701 539 702
rect 623 706 627 707
rect 623 701 627 702
rect 663 706 667 707
rect 663 701 667 702
rect 743 706 747 707
rect 743 701 747 702
rect 791 706 795 707
rect 791 701 795 702
rect 871 706 875 707
rect 871 701 875 702
rect 919 706 923 707
rect 919 701 923 702
rect 999 706 1003 707
rect 999 701 1003 702
rect 1055 706 1059 707
rect 1055 701 1059 702
rect 1127 706 1131 707
rect 1127 701 1131 702
rect 1239 706 1243 707
rect 1239 701 1243 702
rect 1287 706 1291 707
rect 1328 705 1330 725
rect 1368 706 1370 725
rect 1432 706 1434 725
rect 1528 706 1530 725
rect 1632 706 1634 725
rect 1736 706 1738 725
rect 1840 706 1842 725
rect 1944 706 1946 725
rect 2048 706 2050 725
rect 2152 706 2154 725
rect 2256 706 2258 725
rect 2368 706 2370 725
rect 2456 706 2458 725
rect 1366 705 1372 706
rect 1287 701 1291 702
rect 1326 704 1332 705
rect 112 681 114 701
rect 152 682 154 701
rect 208 682 210 701
rect 296 682 298 701
rect 392 682 394 701
rect 504 682 506 701
rect 624 682 626 701
rect 744 682 746 701
rect 872 682 874 701
rect 1000 682 1002 701
rect 1128 682 1130 701
rect 1240 682 1242 701
rect 150 681 156 682
rect 110 680 116 681
rect 110 676 111 680
rect 115 676 116 680
rect 150 677 151 681
rect 155 677 156 681
rect 150 676 156 677
rect 206 681 212 682
rect 206 677 207 681
rect 211 677 212 681
rect 206 676 212 677
rect 294 681 300 682
rect 294 677 295 681
rect 299 677 300 681
rect 294 676 300 677
rect 390 681 396 682
rect 390 677 391 681
rect 395 677 396 681
rect 390 676 396 677
rect 502 681 508 682
rect 502 677 503 681
rect 507 677 508 681
rect 502 676 508 677
rect 622 681 628 682
rect 622 677 623 681
rect 627 677 628 681
rect 622 676 628 677
rect 742 681 748 682
rect 742 677 743 681
rect 747 677 748 681
rect 742 676 748 677
rect 870 681 876 682
rect 870 677 871 681
rect 875 677 876 681
rect 870 676 876 677
rect 998 681 1004 682
rect 998 677 999 681
rect 1003 677 1004 681
rect 998 676 1004 677
rect 1126 681 1132 682
rect 1126 677 1127 681
rect 1131 677 1132 681
rect 1126 676 1132 677
rect 1238 681 1244 682
rect 1288 681 1290 701
rect 1326 700 1327 704
rect 1331 700 1332 704
rect 1366 701 1367 705
rect 1371 701 1372 705
rect 1366 700 1372 701
rect 1430 705 1436 706
rect 1430 701 1431 705
rect 1435 701 1436 705
rect 1430 700 1436 701
rect 1526 705 1532 706
rect 1526 701 1527 705
rect 1531 701 1532 705
rect 1526 700 1532 701
rect 1630 705 1636 706
rect 1630 701 1631 705
rect 1635 701 1636 705
rect 1630 700 1636 701
rect 1734 705 1740 706
rect 1734 701 1735 705
rect 1739 701 1740 705
rect 1734 700 1740 701
rect 1838 705 1844 706
rect 1838 701 1839 705
rect 1843 701 1844 705
rect 1838 700 1844 701
rect 1942 705 1948 706
rect 1942 701 1943 705
rect 1947 701 1948 705
rect 1942 700 1948 701
rect 2046 705 2052 706
rect 2046 701 2047 705
rect 2051 701 2052 705
rect 2046 700 2052 701
rect 2150 705 2156 706
rect 2150 701 2151 705
rect 2155 701 2156 705
rect 2150 700 2156 701
rect 2254 705 2260 706
rect 2254 701 2255 705
rect 2259 701 2260 705
rect 2254 700 2260 701
rect 2366 705 2372 706
rect 2366 701 2367 705
rect 2371 701 2372 705
rect 2366 700 2372 701
rect 2454 705 2460 706
rect 2504 705 2506 725
rect 2454 701 2455 705
rect 2459 701 2460 705
rect 2454 700 2460 701
rect 2502 704 2508 705
rect 2502 700 2503 704
rect 2507 700 2508 704
rect 1326 699 1332 700
rect 2502 699 2508 700
rect 1326 687 1332 688
rect 1326 683 1327 687
rect 1331 683 1332 687
rect 2502 687 2508 688
rect 1326 682 1332 683
rect 1350 684 1356 685
rect 1238 677 1239 681
rect 1243 677 1244 681
rect 1238 676 1244 677
rect 1286 680 1292 681
rect 1286 676 1287 680
rect 1291 676 1292 680
rect 110 675 116 676
rect 1286 675 1292 676
rect 1328 667 1330 682
rect 1350 680 1351 684
rect 1355 680 1356 684
rect 1350 679 1356 680
rect 1414 684 1420 685
rect 1414 680 1415 684
rect 1419 680 1420 684
rect 1414 679 1420 680
rect 1510 684 1516 685
rect 1510 680 1511 684
rect 1515 680 1516 684
rect 1510 679 1516 680
rect 1614 684 1620 685
rect 1614 680 1615 684
rect 1619 680 1620 684
rect 1614 679 1620 680
rect 1718 684 1724 685
rect 1718 680 1719 684
rect 1723 680 1724 684
rect 1718 679 1724 680
rect 1822 684 1828 685
rect 1822 680 1823 684
rect 1827 680 1828 684
rect 1822 679 1828 680
rect 1926 684 1932 685
rect 1926 680 1927 684
rect 1931 680 1932 684
rect 1926 679 1932 680
rect 2030 684 2036 685
rect 2030 680 2031 684
rect 2035 680 2036 684
rect 2030 679 2036 680
rect 2134 684 2140 685
rect 2134 680 2135 684
rect 2139 680 2140 684
rect 2134 679 2140 680
rect 2238 684 2244 685
rect 2238 680 2239 684
rect 2243 680 2244 684
rect 2238 679 2244 680
rect 2350 684 2356 685
rect 2350 680 2351 684
rect 2355 680 2356 684
rect 2350 679 2356 680
rect 2438 684 2444 685
rect 2438 680 2439 684
rect 2443 680 2444 684
rect 2502 683 2503 687
rect 2507 683 2508 687
rect 2502 682 2508 683
rect 2438 679 2444 680
rect 1352 667 1354 679
rect 1416 667 1418 679
rect 1512 667 1514 679
rect 1616 667 1618 679
rect 1720 667 1722 679
rect 1824 667 1826 679
rect 1928 667 1930 679
rect 2032 667 2034 679
rect 2136 667 2138 679
rect 2240 667 2242 679
rect 2352 667 2354 679
rect 2440 667 2442 679
rect 2504 667 2506 682
rect 1327 666 1331 667
rect 110 663 116 664
rect 110 659 111 663
rect 115 659 116 663
rect 1286 663 1292 664
rect 110 658 116 659
rect 134 660 140 661
rect 112 651 114 658
rect 134 656 135 660
rect 139 656 140 660
rect 134 655 140 656
rect 190 660 196 661
rect 190 656 191 660
rect 195 656 196 660
rect 190 655 196 656
rect 278 660 284 661
rect 278 656 279 660
rect 283 656 284 660
rect 278 655 284 656
rect 374 660 380 661
rect 374 656 375 660
rect 379 656 380 660
rect 374 655 380 656
rect 486 660 492 661
rect 486 656 487 660
rect 491 656 492 660
rect 486 655 492 656
rect 606 660 612 661
rect 606 656 607 660
rect 611 656 612 660
rect 606 655 612 656
rect 726 660 732 661
rect 726 656 727 660
rect 731 656 732 660
rect 726 655 732 656
rect 854 660 860 661
rect 854 656 855 660
rect 859 656 860 660
rect 854 655 860 656
rect 982 660 988 661
rect 982 656 983 660
rect 987 656 988 660
rect 982 655 988 656
rect 1110 660 1116 661
rect 1110 656 1111 660
rect 1115 656 1116 660
rect 1110 655 1116 656
rect 1222 660 1228 661
rect 1222 656 1223 660
rect 1227 656 1228 660
rect 1286 659 1287 663
rect 1291 659 1292 663
rect 1327 661 1331 662
rect 1351 666 1355 667
rect 1351 661 1355 662
rect 1415 666 1419 667
rect 1415 661 1419 662
rect 1511 666 1515 667
rect 1511 661 1515 662
rect 1607 666 1611 667
rect 1607 661 1611 662
rect 1615 666 1619 667
rect 1615 661 1619 662
rect 1711 666 1715 667
rect 1711 661 1715 662
rect 1719 666 1723 667
rect 1719 661 1723 662
rect 1823 666 1827 667
rect 1823 661 1827 662
rect 1927 666 1931 667
rect 1927 661 1931 662
rect 1935 666 1939 667
rect 1935 661 1939 662
rect 2031 666 2035 667
rect 2031 661 2035 662
rect 2055 666 2059 667
rect 2055 661 2059 662
rect 2135 666 2139 667
rect 2135 661 2139 662
rect 2183 666 2187 667
rect 2183 661 2187 662
rect 2239 666 2243 667
rect 2239 661 2243 662
rect 2319 666 2323 667
rect 2319 661 2323 662
rect 2351 666 2355 667
rect 2351 661 2355 662
rect 2439 666 2443 667
rect 2439 661 2443 662
rect 2503 666 2507 667
rect 2503 661 2507 662
rect 1286 658 1292 659
rect 1328 658 1330 661
rect 1350 660 1356 661
rect 1222 655 1228 656
rect 136 651 138 655
rect 192 651 194 655
rect 280 651 282 655
rect 376 651 378 655
rect 488 651 490 655
rect 608 651 610 655
rect 728 651 730 655
rect 856 651 858 655
rect 984 651 986 655
rect 1112 651 1114 655
rect 1224 651 1226 655
rect 1288 651 1290 658
rect 1326 657 1332 658
rect 1326 653 1327 657
rect 1331 653 1332 657
rect 1350 656 1351 660
rect 1355 656 1356 660
rect 1350 655 1356 656
rect 1414 660 1420 661
rect 1414 656 1415 660
rect 1419 656 1420 660
rect 1414 655 1420 656
rect 1510 660 1516 661
rect 1510 656 1511 660
rect 1515 656 1516 660
rect 1510 655 1516 656
rect 1606 660 1612 661
rect 1606 656 1607 660
rect 1611 656 1612 660
rect 1606 655 1612 656
rect 1710 660 1716 661
rect 1710 656 1711 660
rect 1715 656 1716 660
rect 1710 655 1716 656
rect 1822 660 1828 661
rect 1822 656 1823 660
rect 1827 656 1828 660
rect 1822 655 1828 656
rect 1934 660 1940 661
rect 1934 656 1935 660
rect 1939 656 1940 660
rect 1934 655 1940 656
rect 2054 660 2060 661
rect 2054 656 2055 660
rect 2059 656 2060 660
rect 2054 655 2060 656
rect 2182 660 2188 661
rect 2182 656 2183 660
rect 2187 656 2188 660
rect 2182 655 2188 656
rect 2318 660 2324 661
rect 2318 656 2319 660
rect 2323 656 2324 660
rect 2318 655 2324 656
rect 2438 660 2444 661
rect 2438 656 2439 660
rect 2443 656 2444 660
rect 2504 658 2506 661
rect 2438 655 2444 656
rect 2502 657 2508 658
rect 1326 652 1332 653
rect 2502 653 2503 657
rect 2507 653 2508 657
rect 2502 652 2508 653
rect 111 650 115 651
rect 111 645 115 646
rect 135 650 139 651
rect 135 645 139 646
rect 151 650 155 651
rect 151 645 155 646
rect 191 650 195 651
rect 191 645 195 646
rect 263 650 267 651
rect 263 645 267 646
rect 279 650 283 651
rect 279 645 283 646
rect 367 650 371 651
rect 367 645 371 646
rect 375 650 379 651
rect 375 645 379 646
rect 463 650 467 651
rect 463 645 467 646
rect 487 650 491 651
rect 487 645 491 646
rect 559 650 563 651
rect 559 645 563 646
rect 607 650 611 651
rect 607 645 611 646
rect 655 650 659 651
rect 655 645 659 646
rect 727 650 731 651
rect 727 645 731 646
rect 751 650 755 651
rect 751 645 755 646
rect 847 650 851 651
rect 847 645 851 646
rect 855 650 859 651
rect 855 645 859 646
rect 943 650 947 651
rect 943 645 947 646
rect 983 650 987 651
rect 983 645 987 646
rect 1039 650 1043 651
rect 1039 645 1043 646
rect 1111 650 1115 651
rect 1111 645 1115 646
rect 1143 650 1147 651
rect 1143 645 1147 646
rect 1223 650 1227 651
rect 1223 645 1227 646
rect 1287 650 1291 651
rect 1287 645 1291 646
rect 112 642 114 645
rect 150 644 156 645
rect 110 641 116 642
rect 110 637 111 641
rect 115 637 116 641
rect 150 640 151 644
rect 155 640 156 644
rect 150 639 156 640
rect 262 644 268 645
rect 262 640 263 644
rect 267 640 268 644
rect 262 639 268 640
rect 366 644 372 645
rect 366 640 367 644
rect 371 640 372 644
rect 366 639 372 640
rect 462 644 468 645
rect 462 640 463 644
rect 467 640 468 644
rect 462 639 468 640
rect 558 644 564 645
rect 558 640 559 644
rect 563 640 564 644
rect 558 639 564 640
rect 654 644 660 645
rect 654 640 655 644
rect 659 640 660 644
rect 654 639 660 640
rect 750 644 756 645
rect 750 640 751 644
rect 755 640 756 644
rect 750 639 756 640
rect 846 644 852 645
rect 846 640 847 644
rect 851 640 852 644
rect 846 639 852 640
rect 942 644 948 645
rect 942 640 943 644
rect 947 640 948 644
rect 942 639 948 640
rect 1038 644 1044 645
rect 1038 640 1039 644
rect 1043 640 1044 644
rect 1038 639 1044 640
rect 1142 644 1148 645
rect 1142 640 1143 644
rect 1147 640 1148 644
rect 1142 639 1148 640
rect 1222 644 1228 645
rect 1222 640 1223 644
rect 1227 640 1228 644
rect 1288 642 1290 645
rect 1222 639 1228 640
rect 1286 641 1292 642
rect 110 636 116 637
rect 1286 637 1287 641
rect 1291 637 1292 641
rect 1286 636 1292 637
rect 1326 640 1332 641
rect 2502 640 2508 641
rect 1326 636 1327 640
rect 1331 636 1332 640
rect 1326 635 1332 636
rect 1366 639 1372 640
rect 1366 635 1367 639
rect 1371 635 1372 639
rect 110 624 116 625
rect 1286 624 1292 625
rect 110 620 111 624
rect 115 620 116 624
rect 110 619 116 620
rect 166 623 172 624
rect 166 619 167 623
rect 171 619 172 623
rect 112 599 114 619
rect 166 618 172 619
rect 278 623 284 624
rect 278 619 279 623
rect 283 619 284 623
rect 278 618 284 619
rect 382 623 388 624
rect 382 619 383 623
rect 387 619 388 623
rect 382 618 388 619
rect 478 623 484 624
rect 478 619 479 623
rect 483 619 484 623
rect 478 618 484 619
rect 574 623 580 624
rect 574 619 575 623
rect 579 619 580 623
rect 574 618 580 619
rect 670 623 676 624
rect 670 619 671 623
rect 675 619 676 623
rect 670 618 676 619
rect 766 623 772 624
rect 766 619 767 623
rect 771 619 772 623
rect 766 618 772 619
rect 862 623 868 624
rect 862 619 863 623
rect 867 619 868 623
rect 862 618 868 619
rect 958 623 964 624
rect 958 619 959 623
rect 963 619 964 623
rect 958 618 964 619
rect 1054 623 1060 624
rect 1054 619 1055 623
rect 1059 619 1060 623
rect 1054 618 1060 619
rect 1158 623 1164 624
rect 1158 619 1159 623
rect 1163 619 1164 623
rect 1158 618 1164 619
rect 1238 623 1244 624
rect 1238 619 1239 623
rect 1243 619 1244 623
rect 1286 620 1287 624
rect 1291 620 1292 624
rect 1286 619 1292 620
rect 1238 618 1244 619
rect 168 599 170 618
rect 280 599 282 618
rect 384 599 386 618
rect 480 599 482 618
rect 576 599 578 618
rect 672 599 674 618
rect 768 599 770 618
rect 864 599 866 618
rect 960 599 962 618
rect 1056 599 1058 618
rect 1160 599 1162 618
rect 1240 599 1242 618
rect 1288 599 1290 619
rect 1328 615 1330 635
rect 1366 634 1372 635
rect 1430 639 1436 640
rect 1430 635 1431 639
rect 1435 635 1436 639
rect 1430 634 1436 635
rect 1526 639 1532 640
rect 1526 635 1527 639
rect 1531 635 1532 639
rect 1526 634 1532 635
rect 1622 639 1628 640
rect 1622 635 1623 639
rect 1627 635 1628 639
rect 1622 634 1628 635
rect 1726 639 1732 640
rect 1726 635 1727 639
rect 1731 635 1732 639
rect 1726 634 1732 635
rect 1838 639 1844 640
rect 1838 635 1839 639
rect 1843 635 1844 639
rect 1838 634 1844 635
rect 1950 639 1956 640
rect 1950 635 1951 639
rect 1955 635 1956 639
rect 1950 634 1956 635
rect 2070 639 2076 640
rect 2070 635 2071 639
rect 2075 635 2076 639
rect 2070 634 2076 635
rect 2198 639 2204 640
rect 2198 635 2199 639
rect 2203 635 2204 639
rect 2198 634 2204 635
rect 2334 639 2340 640
rect 2334 635 2335 639
rect 2339 635 2340 639
rect 2334 634 2340 635
rect 2454 639 2460 640
rect 2454 635 2455 639
rect 2459 635 2460 639
rect 2502 636 2503 640
rect 2507 636 2508 640
rect 2502 635 2508 636
rect 2454 634 2460 635
rect 1368 615 1370 634
rect 1432 615 1434 634
rect 1528 615 1530 634
rect 1624 615 1626 634
rect 1728 615 1730 634
rect 1840 615 1842 634
rect 1952 615 1954 634
rect 2072 615 2074 634
rect 2200 615 2202 634
rect 2336 615 2338 634
rect 2456 615 2458 634
rect 2504 615 2506 635
rect 1327 614 1331 615
rect 1327 609 1331 610
rect 1367 614 1371 615
rect 1367 609 1371 610
rect 1383 614 1387 615
rect 1383 609 1387 610
rect 1431 614 1435 615
rect 1431 609 1435 610
rect 1463 614 1467 615
rect 1463 609 1467 610
rect 1527 614 1531 615
rect 1527 609 1531 610
rect 1551 614 1555 615
rect 1551 609 1555 610
rect 1623 614 1627 615
rect 1623 609 1627 610
rect 1647 614 1651 615
rect 1647 609 1651 610
rect 1727 614 1731 615
rect 1727 609 1731 610
rect 1743 614 1747 615
rect 1743 609 1747 610
rect 1839 614 1843 615
rect 1839 609 1843 610
rect 1847 614 1851 615
rect 1847 609 1851 610
rect 1951 614 1955 615
rect 1951 609 1955 610
rect 1959 614 1963 615
rect 1959 609 1963 610
rect 2071 614 2075 615
rect 2071 609 2075 610
rect 2079 614 2083 615
rect 2079 609 2083 610
rect 2199 614 2203 615
rect 2199 609 2203 610
rect 2207 614 2211 615
rect 2207 609 2211 610
rect 2335 614 2339 615
rect 2335 609 2339 610
rect 2343 614 2347 615
rect 2343 609 2347 610
rect 2455 614 2459 615
rect 2455 609 2459 610
rect 2503 614 2507 615
rect 2503 609 2507 610
rect 111 598 115 599
rect 111 593 115 594
rect 151 598 155 599
rect 151 593 155 594
rect 167 598 171 599
rect 167 593 171 594
rect 239 598 243 599
rect 239 593 243 594
rect 279 598 283 599
rect 279 593 283 594
rect 335 598 339 599
rect 335 593 339 594
rect 383 598 387 599
rect 383 593 387 594
rect 431 598 435 599
rect 431 593 435 594
rect 479 598 483 599
rect 479 593 483 594
rect 535 598 539 599
rect 535 593 539 594
rect 575 598 579 599
rect 575 593 579 594
rect 631 598 635 599
rect 631 593 635 594
rect 671 598 675 599
rect 671 593 675 594
rect 727 598 731 599
rect 727 593 731 594
rect 767 598 771 599
rect 767 593 771 594
rect 823 598 827 599
rect 823 593 827 594
rect 863 598 867 599
rect 863 593 867 594
rect 911 598 915 599
rect 911 593 915 594
rect 959 598 963 599
rect 959 593 963 594
rect 999 598 1003 599
rect 999 593 1003 594
rect 1055 598 1059 599
rect 1055 593 1059 594
rect 1087 598 1091 599
rect 1087 593 1091 594
rect 1159 598 1163 599
rect 1159 593 1163 594
rect 1183 598 1187 599
rect 1183 593 1187 594
rect 1239 598 1243 599
rect 1239 593 1243 594
rect 1287 598 1291 599
rect 1287 593 1291 594
rect 112 573 114 593
rect 152 574 154 593
rect 240 574 242 593
rect 336 574 338 593
rect 432 574 434 593
rect 536 574 538 593
rect 632 574 634 593
rect 728 574 730 593
rect 824 574 826 593
rect 912 574 914 593
rect 1000 574 1002 593
rect 1088 574 1090 593
rect 1184 574 1186 593
rect 150 573 156 574
rect 110 572 116 573
rect 110 568 111 572
rect 115 568 116 572
rect 150 569 151 573
rect 155 569 156 573
rect 150 568 156 569
rect 238 573 244 574
rect 238 569 239 573
rect 243 569 244 573
rect 238 568 244 569
rect 334 573 340 574
rect 334 569 335 573
rect 339 569 340 573
rect 334 568 340 569
rect 430 573 436 574
rect 430 569 431 573
rect 435 569 436 573
rect 430 568 436 569
rect 534 573 540 574
rect 534 569 535 573
rect 539 569 540 573
rect 534 568 540 569
rect 630 573 636 574
rect 630 569 631 573
rect 635 569 636 573
rect 630 568 636 569
rect 726 573 732 574
rect 726 569 727 573
rect 731 569 732 573
rect 726 568 732 569
rect 822 573 828 574
rect 822 569 823 573
rect 827 569 828 573
rect 822 568 828 569
rect 910 573 916 574
rect 910 569 911 573
rect 915 569 916 573
rect 910 568 916 569
rect 998 573 1004 574
rect 998 569 999 573
rect 1003 569 1004 573
rect 998 568 1004 569
rect 1086 573 1092 574
rect 1086 569 1087 573
rect 1091 569 1092 573
rect 1086 568 1092 569
rect 1182 573 1188 574
rect 1288 573 1290 593
rect 1328 589 1330 609
rect 1384 590 1386 609
rect 1464 590 1466 609
rect 1552 590 1554 609
rect 1648 590 1650 609
rect 1744 590 1746 609
rect 1848 590 1850 609
rect 1960 590 1962 609
rect 2080 590 2082 609
rect 2208 590 2210 609
rect 2344 590 2346 609
rect 2456 590 2458 609
rect 1382 589 1388 590
rect 1326 588 1332 589
rect 1326 584 1327 588
rect 1331 584 1332 588
rect 1382 585 1383 589
rect 1387 585 1388 589
rect 1382 584 1388 585
rect 1462 589 1468 590
rect 1462 585 1463 589
rect 1467 585 1468 589
rect 1462 584 1468 585
rect 1550 589 1556 590
rect 1550 585 1551 589
rect 1555 585 1556 589
rect 1550 584 1556 585
rect 1646 589 1652 590
rect 1646 585 1647 589
rect 1651 585 1652 589
rect 1646 584 1652 585
rect 1742 589 1748 590
rect 1742 585 1743 589
rect 1747 585 1748 589
rect 1742 584 1748 585
rect 1846 589 1852 590
rect 1846 585 1847 589
rect 1851 585 1852 589
rect 1846 584 1852 585
rect 1958 589 1964 590
rect 1958 585 1959 589
rect 1963 585 1964 589
rect 1958 584 1964 585
rect 2078 589 2084 590
rect 2078 585 2079 589
rect 2083 585 2084 589
rect 2078 584 2084 585
rect 2206 589 2212 590
rect 2206 585 2207 589
rect 2211 585 2212 589
rect 2206 584 2212 585
rect 2342 589 2348 590
rect 2342 585 2343 589
rect 2347 585 2348 589
rect 2342 584 2348 585
rect 2454 589 2460 590
rect 2504 589 2506 609
rect 2454 585 2455 589
rect 2459 585 2460 589
rect 2454 584 2460 585
rect 2502 588 2508 589
rect 2502 584 2503 588
rect 2507 584 2508 588
rect 1326 583 1332 584
rect 2502 583 2508 584
rect 1182 569 1183 573
rect 1187 569 1188 573
rect 1182 568 1188 569
rect 1286 572 1292 573
rect 1286 568 1287 572
rect 1291 568 1292 572
rect 110 567 116 568
rect 1286 567 1292 568
rect 1326 571 1332 572
rect 1326 567 1327 571
rect 1331 567 1332 571
rect 2502 571 2508 572
rect 1326 566 1332 567
rect 1366 568 1372 569
rect 1328 563 1330 566
rect 1366 564 1367 568
rect 1371 564 1372 568
rect 1366 563 1372 564
rect 1446 568 1452 569
rect 1446 564 1447 568
rect 1451 564 1452 568
rect 1446 563 1452 564
rect 1534 568 1540 569
rect 1534 564 1535 568
rect 1539 564 1540 568
rect 1534 563 1540 564
rect 1630 568 1636 569
rect 1630 564 1631 568
rect 1635 564 1636 568
rect 1630 563 1636 564
rect 1726 568 1732 569
rect 1726 564 1727 568
rect 1731 564 1732 568
rect 1726 563 1732 564
rect 1830 568 1836 569
rect 1830 564 1831 568
rect 1835 564 1836 568
rect 1830 563 1836 564
rect 1942 568 1948 569
rect 1942 564 1943 568
rect 1947 564 1948 568
rect 1942 563 1948 564
rect 2062 568 2068 569
rect 2062 564 2063 568
rect 2067 564 2068 568
rect 2062 563 2068 564
rect 2190 568 2196 569
rect 2190 564 2191 568
rect 2195 564 2196 568
rect 2190 563 2196 564
rect 2326 568 2332 569
rect 2326 564 2327 568
rect 2331 564 2332 568
rect 2326 563 2332 564
rect 2438 568 2444 569
rect 2438 564 2439 568
rect 2443 564 2444 568
rect 2502 567 2503 571
rect 2507 567 2508 571
rect 2502 566 2508 567
rect 2438 563 2444 564
rect 2504 563 2506 566
rect 1327 562 1331 563
rect 1327 557 1331 558
rect 1367 562 1371 563
rect 1367 557 1371 558
rect 1375 562 1379 563
rect 1375 557 1379 558
rect 1447 562 1451 563
rect 1447 557 1451 558
rect 1455 562 1459 563
rect 1455 557 1459 558
rect 1535 562 1539 563
rect 1535 557 1539 558
rect 1551 562 1555 563
rect 1551 557 1555 558
rect 1631 562 1635 563
rect 1631 557 1635 558
rect 1647 562 1651 563
rect 1647 557 1651 558
rect 1727 562 1731 563
rect 1727 557 1731 558
rect 1751 562 1755 563
rect 1751 557 1755 558
rect 1831 562 1835 563
rect 1831 557 1835 558
rect 1855 562 1859 563
rect 1855 557 1859 558
rect 1943 562 1947 563
rect 1943 557 1947 558
rect 1959 562 1963 563
rect 1959 557 1963 558
rect 2055 562 2059 563
rect 2055 557 2059 558
rect 2063 562 2067 563
rect 2063 557 2067 558
rect 2151 562 2155 563
rect 2151 557 2155 558
rect 2191 562 2195 563
rect 2191 557 2195 558
rect 2255 562 2259 563
rect 2255 557 2259 558
rect 2327 562 2331 563
rect 2327 557 2331 558
rect 2359 562 2363 563
rect 2359 557 2363 558
rect 2439 562 2443 563
rect 2439 557 2443 558
rect 2503 562 2507 563
rect 2503 557 2507 558
rect 110 555 116 556
rect 110 551 111 555
rect 115 551 116 555
rect 1286 555 1292 556
rect 110 550 116 551
rect 134 552 140 553
rect 112 539 114 550
rect 134 548 135 552
rect 139 548 140 552
rect 134 547 140 548
rect 222 552 228 553
rect 222 548 223 552
rect 227 548 228 552
rect 222 547 228 548
rect 318 552 324 553
rect 318 548 319 552
rect 323 548 324 552
rect 318 547 324 548
rect 414 552 420 553
rect 414 548 415 552
rect 419 548 420 552
rect 414 547 420 548
rect 518 552 524 553
rect 518 548 519 552
rect 523 548 524 552
rect 518 547 524 548
rect 614 552 620 553
rect 614 548 615 552
rect 619 548 620 552
rect 614 547 620 548
rect 710 552 716 553
rect 710 548 711 552
rect 715 548 716 552
rect 710 547 716 548
rect 806 552 812 553
rect 806 548 807 552
rect 811 548 812 552
rect 806 547 812 548
rect 894 552 900 553
rect 894 548 895 552
rect 899 548 900 552
rect 894 547 900 548
rect 982 552 988 553
rect 982 548 983 552
rect 987 548 988 552
rect 982 547 988 548
rect 1070 552 1076 553
rect 1070 548 1071 552
rect 1075 548 1076 552
rect 1070 547 1076 548
rect 1166 552 1172 553
rect 1166 548 1167 552
rect 1171 548 1172 552
rect 1286 551 1287 555
rect 1291 551 1292 555
rect 1328 554 1330 557
rect 1374 556 1380 557
rect 1286 550 1292 551
rect 1326 553 1332 554
rect 1166 547 1172 548
rect 136 539 138 547
rect 224 539 226 547
rect 320 539 322 547
rect 416 539 418 547
rect 520 539 522 547
rect 616 539 618 547
rect 712 539 714 547
rect 808 539 810 547
rect 896 539 898 547
rect 984 539 986 547
rect 1072 539 1074 547
rect 1168 539 1170 547
rect 1288 539 1290 550
rect 1326 549 1327 553
rect 1331 549 1332 553
rect 1374 552 1375 556
rect 1379 552 1380 556
rect 1374 551 1380 552
rect 1454 556 1460 557
rect 1454 552 1455 556
rect 1459 552 1460 556
rect 1454 551 1460 552
rect 1550 556 1556 557
rect 1550 552 1551 556
rect 1555 552 1556 556
rect 1550 551 1556 552
rect 1646 556 1652 557
rect 1646 552 1647 556
rect 1651 552 1652 556
rect 1646 551 1652 552
rect 1750 556 1756 557
rect 1750 552 1751 556
rect 1755 552 1756 556
rect 1750 551 1756 552
rect 1854 556 1860 557
rect 1854 552 1855 556
rect 1859 552 1860 556
rect 1854 551 1860 552
rect 1958 556 1964 557
rect 1958 552 1959 556
rect 1963 552 1964 556
rect 1958 551 1964 552
rect 2054 556 2060 557
rect 2054 552 2055 556
rect 2059 552 2060 556
rect 2054 551 2060 552
rect 2150 556 2156 557
rect 2150 552 2151 556
rect 2155 552 2156 556
rect 2150 551 2156 552
rect 2254 556 2260 557
rect 2254 552 2255 556
rect 2259 552 2260 556
rect 2254 551 2260 552
rect 2358 556 2364 557
rect 2358 552 2359 556
rect 2363 552 2364 556
rect 2358 551 2364 552
rect 2438 556 2444 557
rect 2438 552 2439 556
rect 2443 552 2444 556
rect 2504 554 2506 557
rect 2438 551 2444 552
rect 2502 553 2508 554
rect 1326 548 1332 549
rect 2502 549 2503 553
rect 2507 549 2508 553
rect 2502 548 2508 549
rect 111 538 115 539
rect 111 533 115 534
rect 135 538 139 539
rect 135 533 139 534
rect 143 538 147 539
rect 143 533 147 534
rect 223 538 227 539
rect 223 533 227 534
rect 239 538 243 539
rect 239 533 243 534
rect 319 538 323 539
rect 319 533 323 534
rect 335 538 339 539
rect 335 533 339 534
rect 415 538 419 539
rect 415 533 419 534
rect 431 538 435 539
rect 431 533 435 534
rect 519 538 523 539
rect 519 533 523 534
rect 527 538 531 539
rect 527 533 531 534
rect 615 538 619 539
rect 615 533 619 534
rect 623 538 627 539
rect 623 533 627 534
rect 711 538 715 539
rect 711 533 715 534
rect 791 538 795 539
rect 791 533 795 534
rect 807 538 811 539
rect 807 533 811 534
rect 871 538 875 539
rect 871 533 875 534
rect 895 538 899 539
rect 895 533 899 534
rect 951 538 955 539
rect 951 533 955 534
rect 983 538 987 539
rect 983 533 987 534
rect 1031 538 1035 539
rect 1031 533 1035 534
rect 1071 538 1075 539
rect 1071 533 1075 534
rect 1167 538 1171 539
rect 1167 533 1171 534
rect 1287 538 1291 539
rect 1287 533 1291 534
rect 1326 536 1332 537
rect 2502 536 2508 537
rect 112 530 114 533
rect 142 532 148 533
rect 110 529 116 530
rect 110 525 111 529
rect 115 525 116 529
rect 142 528 143 532
rect 147 528 148 532
rect 142 527 148 528
rect 238 532 244 533
rect 238 528 239 532
rect 243 528 244 532
rect 238 527 244 528
rect 334 532 340 533
rect 334 528 335 532
rect 339 528 340 532
rect 334 527 340 528
rect 430 532 436 533
rect 430 528 431 532
rect 435 528 436 532
rect 430 527 436 528
rect 526 532 532 533
rect 526 528 527 532
rect 531 528 532 532
rect 526 527 532 528
rect 622 532 628 533
rect 622 528 623 532
rect 627 528 628 532
rect 622 527 628 528
rect 710 532 716 533
rect 710 528 711 532
rect 715 528 716 532
rect 710 527 716 528
rect 790 532 796 533
rect 790 528 791 532
rect 795 528 796 532
rect 790 527 796 528
rect 870 532 876 533
rect 870 528 871 532
rect 875 528 876 532
rect 870 527 876 528
rect 950 532 956 533
rect 950 528 951 532
rect 955 528 956 532
rect 950 527 956 528
rect 1030 532 1036 533
rect 1030 528 1031 532
rect 1035 528 1036 532
rect 1288 530 1290 533
rect 1326 532 1327 536
rect 1331 532 1332 536
rect 1326 531 1332 532
rect 1390 535 1396 536
rect 1390 531 1391 535
rect 1395 531 1396 535
rect 1030 527 1036 528
rect 1286 529 1292 530
rect 110 524 116 525
rect 1286 525 1287 529
rect 1291 525 1292 529
rect 1286 524 1292 525
rect 110 512 116 513
rect 1286 512 1292 513
rect 110 508 111 512
rect 115 508 116 512
rect 110 507 116 508
rect 158 511 164 512
rect 158 507 159 511
rect 163 507 164 511
rect 112 483 114 507
rect 158 506 164 507
rect 254 511 260 512
rect 254 507 255 511
rect 259 507 260 511
rect 254 506 260 507
rect 350 511 356 512
rect 350 507 351 511
rect 355 507 356 511
rect 350 506 356 507
rect 446 511 452 512
rect 446 507 447 511
rect 451 507 452 511
rect 446 506 452 507
rect 542 511 548 512
rect 542 507 543 511
rect 547 507 548 511
rect 542 506 548 507
rect 638 511 644 512
rect 638 507 639 511
rect 643 507 644 511
rect 638 506 644 507
rect 726 511 732 512
rect 726 507 727 511
rect 731 507 732 511
rect 726 506 732 507
rect 806 511 812 512
rect 806 507 807 511
rect 811 507 812 511
rect 806 506 812 507
rect 886 511 892 512
rect 886 507 887 511
rect 891 507 892 511
rect 886 506 892 507
rect 966 511 972 512
rect 966 507 967 511
rect 971 507 972 511
rect 966 506 972 507
rect 1046 511 1052 512
rect 1046 507 1047 511
rect 1051 507 1052 511
rect 1286 508 1287 512
rect 1291 508 1292 512
rect 1286 507 1292 508
rect 1328 507 1330 531
rect 1390 530 1396 531
rect 1470 535 1476 536
rect 1470 531 1471 535
rect 1475 531 1476 535
rect 1470 530 1476 531
rect 1566 535 1572 536
rect 1566 531 1567 535
rect 1571 531 1572 535
rect 1566 530 1572 531
rect 1662 535 1668 536
rect 1662 531 1663 535
rect 1667 531 1668 535
rect 1662 530 1668 531
rect 1766 535 1772 536
rect 1766 531 1767 535
rect 1771 531 1772 535
rect 1766 530 1772 531
rect 1870 535 1876 536
rect 1870 531 1871 535
rect 1875 531 1876 535
rect 1870 530 1876 531
rect 1974 535 1980 536
rect 1974 531 1975 535
rect 1979 531 1980 535
rect 1974 530 1980 531
rect 2070 535 2076 536
rect 2070 531 2071 535
rect 2075 531 2076 535
rect 2070 530 2076 531
rect 2166 535 2172 536
rect 2166 531 2167 535
rect 2171 531 2172 535
rect 2166 530 2172 531
rect 2270 535 2276 536
rect 2270 531 2271 535
rect 2275 531 2276 535
rect 2270 530 2276 531
rect 2374 535 2380 536
rect 2374 531 2375 535
rect 2379 531 2380 535
rect 2374 530 2380 531
rect 2454 535 2460 536
rect 2454 531 2455 535
rect 2459 531 2460 535
rect 2502 532 2503 536
rect 2507 532 2508 536
rect 2502 531 2508 532
rect 2454 530 2460 531
rect 1392 507 1394 530
rect 1472 507 1474 530
rect 1568 507 1570 530
rect 1664 507 1666 530
rect 1768 507 1770 530
rect 1872 507 1874 530
rect 1976 507 1978 530
rect 2072 507 2074 530
rect 2168 507 2170 530
rect 2272 507 2274 530
rect 2376 507 2378 530
rect 2456 507 2458 530
rect 2504 507 2506 531
rect 1046 506 1052 507
rect 160 483 162 506
rect 256 483 258 506
rect 352 483 354 506
rect 448 483 450 506
rect 544 483 546 506
rect 640 483 642 506
rect 728 483 730 506
rect 808 483 810 506
rect 888 483 890 506
rect 968 483 970 506
rect 1048 483 1050 506
rect 1288 483 1290 507
rect 1327 506 1331 507
rect 1327 501 1331 502
rect 1367 506 1371 507
rect 1367 501 1371 502
rect 1391 506 1395 507
rect 1391 501 1395 502
rect 1455 506 1459 507
rect 1455 501 1459 502
rect 1471 506 1475 507
rect 1471 501 1475 502
rect 1567 506 1571 507
rect 1567 501 1571 502
rect 1575 506 1579 507
rect 1575 501 1579 502
rect 1663 506 1667 507
rect 1663 501 1667 502
rect 1695 506 1699 507
rect 1695 501 1699 502
rect 1767 506 1771 507
rect 1767 501 1771 502
rect 1807 506 1811 507
rect 1807 501 1811 502
rect 1871 506 1875 507
rect 1871 501 1875 502
rect 1919 506 1923 507
rect 1919 501 1923 502
rect 1975 506 1979 507
rect 1975 501 1979 502
rect 2023 506 2027 507
rect 2023 501 2027 502
rect 2071 506 2075 507
rect 2071 501 2075 502
rect 2119 506 2123 507
rect 2119 501 2123 502
rect 2167 506 2171 507
rect 2167 501 2171 502
rect 2207 506 2211 507
rect 2207 501 2211 502
rect 2271 506 2275 507
rect 2271 501 2275 502
rect 2295 506 2299 507
rect 2295 501 2299 502
rect 2375 506 2379 507
rect 2375 501 2379 502
rect 2383 506 2387 507
rect 2383 501 2387 502
rect 2455 506 2459 507
rect 2455 501 2459 502
rect 2503 506 2507 507
rect 2503 501 2507 502
rect 111 482 115 483
rect 111 477 115 478
rect 151 482 155 483
rect 151 477 155 478
rect 159 482 163 483
rect 159 477 163 478
rect 207 482 211 483
rect 207 477 211 478
rect 255 482 259 483
rect 255 477 259 478
rect 287 482 291 483
rect 287 477 291 478
rect 351 482 355 483
rect 351 477 355 478
rect 375 482 379 483
rect 375 477 379 478
rect 447 482 451 483
rect 447 477 451 478
rect 463 482 467 483
rect 463 477 467 478
rect 543 482 547 483
rect 543 477 547 478
rect 559 482 563 483
rect 559 477 563 478
rect 639 482 643 483
rect 639 477 643 478
rect 655 482 659 483
rect 655 477 659 478
rect 727 482 731 483
rect 727 477 731 478
rect 751 482 755 483
rect 751 477 755 478
rect 807 482 811 483
rect 807 477 811 478
rect 847 482 851 483
rect 847 477 851 478
rect 887 482 891 483
rect 887 477 891 478
rect 951 482 955 483
rect 951 477 955 478
rect 967 482 971 483
rect 967 477 971 478
rect 1047 482 1051 483
rect 1047 477 1051 478
rect 1055 482 1059 483
rect 1055 477 1059 478
rect 1159 482 1163 483
rect 1159 477 1163 478
rect 1239 482 1243 483
rect 1239 477 1243 478
rect 1287 482 1291 483
rect 1328 481 1330 501
rect 1368 482 1370 501
rect 1456 482 1458 501
rect 1576 482 1578 501
rect 1696 482 1698 501
rect 1808 482 1810 501
rect 1920 482 1922 501
rect 2024 482 2026 501
rect 2120 482 2122 501
rect 2208 482 2210 501
rect 2296 482 2298 501
rect 2384 482 2386 501
rect 2456 482 2458 501
rect 1366 481 1372 482
rect 1287 477 1291 478
rect 1326 480 1332 481
rect 112 457 114 477
rect 152 458 154 477
rect 208 458 210 477
rect 288 458 290 477
rect 376 458 378 477
rect 464 458 466 477
rect 560 458 562 477
rect 656 458 658 477
rect 752 458 754 477
rect 848 458 850 477
rect 952 458 954 477
rect 1056 458 1058 477
rect 1160 458 1162 477
rect 1240 458 1242 477
rect 150 457 156 458
rect 110 456 116 457
rect 110 452 111 456
rect 115 452 116 456
rect 150 453 151 457
rect 155 453 156 457
rect 150 452 156 453
rect 206 457 212 458
rect 206 453 207 457
rect 211 453 212 457
rect 206 452 212 453
rect 286 457 292 458
rect 286 453 287 457
rect 291 453 292 457
rect 286 452 292 453
rect 374 457 380 458
rect 374 453 375 457
rect 379 453 380 457
rect 374 452 380 453
rect 462 457 468 458
rect 462 453 463 457
rect 467 453 468 457
rect 462 452 468 453
rect 558 457 564 458
rect 558 453 559 457
rect 563 453 564 457
rect 558 452 564 453
rect 654 457 660 458
rect 654 453 655 457
rect 659 453 660 457
rect 654 452 660 453
rect 750 457 756 458
rect 750 453 751 457
rect 755 453 756 457
rect 750 452 756 453
rect 846 457 852 458
rect 846 453 847 457
rect 851 453 852 457
rect 846 452 852 453
rect 950 457 956 458
rect 950 453 951 457
rect 955 453 956 457
rect 950 452 956 453
rect 1054 457 1060 458
rect 1054 453 1055 457
rect 1059 453 1060 457
rect 1054 452 1060 453
rect 1158 457 1164 458
rect 1158 453 1159 457
rect 1163 453 1164 457
rect 1158 452 1164 453
rect 1238 457 1244 458
rect 1288 457 1290 477
rect 1326 476 1327 480
rect 1331 476 1332 480
rect 1366 477 1367 481
rect 1371 477 1372 481
rect 1366 476 1372 477
rect 1454 481 1460 482
rect 1454 477 1455 481
rect 1459 477 1460 481
rect 1454 476 1460 477
rect 1574 481 1580 482
rect 1574 477 1575 481
rect 1579 477 1580 481
rect 1574 476 1580 477
rect 1694 481 1700 482
rect 1694 477 1695 481
rect 1699 477 1700 481
rect 1694 476 1700 477
rect 1806 481 1812 482
rect 1806 477 1807 481
rect 1811 477 1812 481
rect 1806 476 1812 477
rect 1918 481 1924 482
rect 1918 477 1919 481
rect 1923 477 1924 481
rect 1918 476 1924 477
rect 2022 481 2028 482
rect 2022 477 2023 481
rect 2027 477 2028 481
rect 2022 476 2028 477
rect 2118 481 2124 482
rect 2118 477 2119 481
rect 2123 477 2124 481
rect 2118 476 2124 477
rect 2206 481 2212 482
rect 2206 477 2207 481
rect 2211 477 2212 481
rect 2206 476 2212 477
rect 2294 481 2300 482
rect 2294 477 2295 481
rect 2299 477 2300 481
rect 2294 476 2300 477
rect 2382 481 2388 482
rect 2382 477 2383 481
rect 2387 477 2388 481
rect 2382 476 2388 477
rect 2454 481 2460 482
rect 2504 481 2506 501
rect 2454 477 2455 481
rect 2459 477 2460 481
rect 2454 476 2460 477
rect 2502 480 2508 481
rect 2502 476 2503 480
rect 2507 476 2508 480
rect 1326 475 1332 476
rect 2502 475 2508 476
rect 1326 463 1332 464
rect 1326 459 1327 463
rect 1331 459 1332 463
rect 2502 463 2508 464
rect 1326 458 1332 459
rect 1350 460 1356 461
rect 1238 453 1239 457
rect 1243 453 1244 457
rect 1238 452 1244 453
rect 1286 456 1292 457
rect 1286 452 1287 456
rect 1291 452 1292 456
rect 110 451 116 452
rect 1286 451 1292 452
rect 1328 443 1330 458
rect 1350 456 1351 460
rect 1355 456 1356 460
rect 1350 455 1356 456
rect 1438 460 1444 461
rect 1438 456 1439 460
rect 1443 456 1444 460
rect 1438 455 1444 456
rect 1558 460 1564 461
rect 1558 456 1559 460
rect 1563 456 1564 460
rect 1558 455 1564 456
rect 1678 460 1684 461
rect 1678 456 1679 460
rect 1683 456 1684 460
rect 1678 455 1684 456
rect 1790 460 1796 461
rect 1790 456 1791 460
rect 1795 456 1796 460
rect 1790 455 1796 456
rect 1902 460 1908 461
rect 1902 456 1903 460
rect 1907 456 1908 460
rect 1902 455 1908 456
rect 2006 460 2012 461
rect 2006 456 2007 460
rect 2011 456 2012 460
rect 2006 455 2012 456
rect 2102 460 2108 461
rect 2102 456 2103 460
rect 2107 456 2108 460
rect 2102 455 2108 456
rect 2190 460 2196 461
rect 2190 456 2191 460
rect 2195 456 2196 460
rect 2190 455 2196 456
rect 2278 460 2284 461
rect 2278 456 2279 460
rect 2283 456 2284 460
rect 2278 455 2284 456
rect 2366 460 2372 461
rect 2366 456 2367 460
rect 2371 456 2372 460
rect 2366 455 2372 456
rect 2438 460 2444 461
rect 2438 456 2439 460
rect 2443 456 2444 460
rect 2502 459 2503 463
rect 2507 459 2508 463
rect 2502 458 2508 459
rect 2438 455 2444 456
rect 1352 443 1354 455
rect 1440 443 1442 455
rect 1560 443 1562 455
rect 1680 443 1682 455
rect 1792 443 1794 455
rect 1904 443 1906 455
rect 2008 443 2010 455
rect 2104 443 2106 455
rect 2192 443 2194 455
rect 2280 443 2282 455
rect 2368 443 2370 455
rect 2440 443 2442 455
rect 2504 443 2506 458
rect 1327 442 1331 443
rect 110 439 116 440
rect 110 435 111 439
rect 115 435 116 439
rect 1286 439 1292 440
rect 110 434 116 435
rect 134 436 140 437
rect 112 431 114 434
rect 134 432 135 436
rect 139 432 140 436
rect 134 431 140 432
rect 190 436 196 437
rect 190 432 191 436
rect 195 432 196 436
rect 190 431 196 432
rect 270 436 276 437
rect 270 432 271 436
rect 275 432 276 436
rect 270 431 276 432
rect 358 436 364 437
rect 358 432 359 436
rect 363 432 364 436
rect 358 431 364 432
rect 446 436 452 437
rect 446 432 447 436
rect 451 432 452 436
rect 446 431 452 432
rect 542 436 548 437
rect 542 432 543 436
rect 547 432 548 436
rect 542 431 548 432
rect 638 436 644 437
rect 638 432 639 436
rect 643 432 644 436
rect 638 431 644 432
rect 734 436 740 437
rect 734 432 735 436
rect 739 432 740 436
rect 734 431 740 432
rect 830 436 836 437
rect 830 432 831 436
rect 835 432 836 436
rect 830 431 836 432
rect 934 436 940 437
rect 934 432 935 436
rect 939 432 940 436
rect 934 431 940 432
rect 1038 436 1044 437
rect 1038 432 1039 436
rect 1043 432 1044 436
rect 1038 431 1044 432
rect 1142 436 1148 437
rect 1142 432 1143 436
rect 1147 432 1148 436
rect 1142 431 1148 432
rect 1222 436 1228 437
rect 1222 432 1223 436
rect 1227 432 1228 436
rect 1286 435 1287 439
rect 1291 435 1292 439
rect 1327 437 1331 438
rect 1351 442 1355 443
rect 1351 437 1355 438
rect 1439 442 1443 443
rect 1439 437 1443 438
rect 1559 442 1563 443
rect 1559 437 1563 438
rect 1583 442 1587 443
rect 1583 437 1587 438
rect 1639 442 1643 443
rect 1639 437 1643 438
rect 1679 442 1683 443
rect 1679 437 1683 438
rect 1695 442 1699 443
rect 1695 437 1699 438
rect 1759 442 1763 443
rect 1759 437 1763 438
rect 1791 442 1795 443
rect 1791 437 1795 438
rect 1831 442 1835 443
rect 1831 437 1835 438
rect 1903 442 1907 443
rect 1903 437 1907 438
rect 1911 442 1915 443
rect 1911 437 1915 438
rect 1991 442 1995 443
rect 1991 437 1995 438
rect 2007 442 2011 443
rect 2007 437 2011 438
rect 2079 442 2083 443
rect 2079 437 2083 438
rect 2103 442 2107 443
rect 2103 437 2107 438
rect 2175 442 2179 443
rect 2175 437 2179 438
rect 2191 442 2195 443
rect 2191 437 2195 438
rect 2271 442 2275 443
rect 2271 437 2275 438
rect 2279 442 2283 443
rect 2279 437 2283 438
rect 2367 442 2371 443
rect 2367 437 2371 438
rect 2439 442 2443 443
rect 2439 437 2443 438
rect 2503 442 2507 443
rect 2503 437 2507 438
rect 1286 434 1292 435
rect 1328 434 1330 437
rect 1582 436 1588 437
rect 1222 431 1228 432
rect 1288 431 1290 434
rect 1326 433 1332 434
rect 111 430 115 431
rect 111 425 115 426
rect 135 430 139 431
rect 135 425 139 426
rect 191 430 195 431
rect 191 425 195 426
rect 271 430 275 431
rect 271 425 275 426
rect 279 430 283 431
rect 279 425 283 426
rect 359 430 363 431
rect 359 425 363 426
rect 383 430 387 431
rect 383 425 387 426
rect 447 430 451 431
rect 447 425 451 426
rect 495 430 499 431
rect 495 425 499 426
rect 543 430 547 431
rect 543 425 547 426
rect 607 430 611 431
rect 607 425 611 426
rect 639 430 643 431
rect 639 425 643 426
rect 719 430 723 431
rect 719 425 723 426
rect 735 430 739 431
rect 735 425 739 426
rect 831 430 835 431
rect 831 425 835 426
rect 935 430 939 431
rect 935 425 939 426
rect 1039 430 1043 431
rect 1039 425 1043 426
rect 1143 430 1147 431
rect 1143 425 1147 426
rect 1223 430 1227 431
rect 1223 425 1227 426
rect 1287 430 1291 431
rect 1326 429 1327 433
rect 1331 429 1332 433
rect 1582 432 1583 436
rect 1587 432 1588 436
rect 1582 431 1588 432
rect 1638 436 1644 437
rect 1638 432 1639 436
rect 1643 432 1644 436
rect 1638 431 1644 432
rect 1694 436 1700 437
rect 1694 432 1695 436
rect 1699 432 1700 436
rect 1694 431 1700 432
rect 1758 436 1764 437
rect 1758 432 1759 436
rect 1763 432 1764 436
rect 1758 431 1764 432
rect 1830 436 1836 437
rect 1830 432 1831 436
rect 1835 432 1836 436
rect 1830 431 1836 432
rect 1910 436 1916 437
rect 1910 432 1911 436
rect 1915 432 1916 436
rect 1910 431 1916 432
rect 1990 436 1996 437
rect 1990 432 1991 436
rect 1995 432 1996 436
rect 1990 431 1996 432
rect 2078 436 2084 437
rect 2078 432 2079 436
rect 2083 432 2084 436
rect 2078 431 2084 432
rect 2174 436 2180 437
rect 2174 432 2175 436
rect 2179 432 2180 436
rect 2174 431 2180 432
rect 2270 436 2276 437
rect 2270 432 2271 436
rect 2275 432 2276 436
rect 2270 431 2276 432
rect 2366 436 2372 437
rect 2366 432 2367 436
rect 2371 432 2372 436
rect 2366 431 2372 432
rect 2438 436 2444 437
rect 2438 432 2439 436
rect 2443 432 2444 436
rect 2504 434 2506 437
rect 2438 431 2444 432
rect 2502 433 2508 434
rect 1326 428 1332 429
rect 2502 429 2503 433
rect 2507 429 2508 433
rect 2502 428 2508 429
rect 1287 425 1291 426
rect 112 422 114 425
rect 134 424 140 425
rect 110 421 116 422
rect 110 417 111 421
rect 115 417 116 421
rect 134 420 135 424
rect 139 420 140 424
rect 134 419 140 420
rect 190 424 196 425
rect 190 420 191 424
rect 195 420 196 424
rect 190 419 196 420
rect 278 424 284 425
rect 278 420 279 424
rect 283 420 284 424
rect 278 419 284 420
rect 382 424 388 425
rect 382 420 383 424
rect 387 420 388 424
rect 382 419 388 420
rect 494 424 500 425
rect 494 420 495 424
rect 499 420 500 424
rect 494 419 500 420
rect 606 424 612 425
rect 606 420 607 424
rect 611 420 612 424
rect 606 419 612 420
rect 718 424 724 425
rect 718 420 719 424
rect 723 420 724 424
rect 718 419 724 420
rect 830 424 836 425
rect 830 420 831 424
rect 835 420 836 424
rect 830 419 836 420
rect 934 424 940 425
rect 934 420 935 424
rect 939 420 940 424
rect 934 419 940 420
rect 1038 424 1044 425
rect 1038 420 1039 424
rect 1043 420 1044 424
rect 1038 419 1044 420
rect 1142 424 1148 425
rect 1142 420 1143 424
rect 1147 420 1148 424
rect 1142 419 1148 420
rect 1222 424 1228 425
rect 1222 420 1223 424
rect 1227 420 1228 424
rect 1288 422 1290 425
rect 1222 419 1228 420
rect 1286 421 1292 422
rect 110 416 116 417
rect 1286 417 1287 421
rect 1291 417 1292 421
rect 1286 416 1292 417
rect 1326 416 1332 417
rect 2502 416 2508 417
rect 1326 412 1327 416
rect 1331 412 1332 416
rect 1326 411 1332 412
rect 1598 415 1604 416
rect 1598 411 1599 415
rect 1603 411 1604 415
rect 110 404 116 405
rect 1286 404 1292 405
rect 110 400 111 404
rect 115 400 116 404
rect 110 399 116 400
rect 150 403 156 404
rect 150 399 151 403
rect 155 399 156 403
rect 112 375 114 399
rect 150 398 156 399
rect 206 403 212 404
rect 206 399 207 403
rect 211 399 212 403
rect 206 398 212 399
rect 294 403 300 404
rect 294 399 295 403
rect 299 399 300 403
rect 294 398 300 399
rect 398 403 404 404
rect 398 399 399 403
rect 403 399 404 403
rect 398 398 404 399
rect 510 403 516 404
rect 510 399 511 403
rect 515 399 516 403
rect 510 398 516 399
rect 622 403 628 404
rect 622 399 623 403
rect 627 399 628 403
rect 622 398 628 399
rect 734 403 740 404
rect 734 399 735 403
rect 739 399 740 403
rect 734 398 740 399
rect 846 403 852 404
rect 846 399 847 403
rect 851 399 852 403
rect 846 398 852 399
rect 950 403 956 404
rect 950 399 951 403
rect 955 399 956 403
rect 950 398 956 399
rect 1054 403 1060 404
rect 1054 399 1055 403
rect 1059 399 1060 403
rect 1054 398 1060 399
rect 1158 403 1164 404
rect 1158 399 1159 403
rect 1163 399 1164 403
rect 1158 398 1164 399
rect 1238 403 1244 404
rect 1238 399 1239 403
rect 1243 399 1244 403
rect 1286 400 1287 404
rect 1291 400 1292 404
rect 1286 399 1292 400
rect 1238 398 1244 399
rect 152 375 154 398
rect 208 375 210 398
rect 296 375 298 398
rect 400 375 402 398
rect 512 375 514 398
rect 624 375 626 398
rect 736 375 738 398
rect 848 375 850 398
rect 952 375 954 398
rect 1056 375 1058 398
rect 1160 375 1162 398
rect 1240 375 1242 398
rect 1288 375 1290 399
rect 1328 387 1330 411
rect 1598 410 1604 411
rect 1654 415 1660 416
rect 1654 411 1655 415
rect 1659 411 1660 415
rect 1654 410 1660 411
rect 1710 415 1716 416
rect 1710 411 1711 415
rect 1715 411 1716 415
rect 1710 410 1716 411
rect 1774 415 1780 416
rect 1774 411 1775 415
rect 1779 411 1780 415
rect 1774 410 1780 411
rect 1846 415 1852 416
rect 1846 411 1847 415
rect 1851 411 1852 415
rect 1846 410 1852 411
rect 1926 415 1932 416
rect 1926 411 1927 415
rect 1931 411 1932 415
rect 1926 410 1932 411
rect 2006 415 2012 416
rect 2006 411 2007 415
rect 2011 411 2012 415
rect 2006 410 2012 411
rect 2094 415 2100 416
rect 2094 411 2095 415
rect 2099 411 2100 415
rect 2094 410 2100 411
rect 2190 415 2196 416
rect 2190 411 2191 415
rect 2195 411 2196 415
rect 2190 410 2196 411
rect 2286 415 2292 416
rect 2286 411 2287 415
rect 2291 411 2292 415
rect 2286 410 2292 411
rect 2382 415 2388 416
rect 2382 411 2383 415
rect 2387 411 2388 415
rect 2382 410 2388 411
rect 2454 415 2460 416
rect 2454 411 2455 415
rect 2459 411 2460 415
rect 2502 412 2503 416
rect 2507 412 2508 416
rect 2502 411 2508 412
rect 2454 410 2460 411
rect 1600 387 1602 410
rect 1656 387 1658 410
rect 1712 387 1714 410
rect 1776 387 1778 410
rect 1848 387 1850 410
rect 1928 387 1930 410
rect 2008 387 2010 410
rect 2096 387 2098 410
rect 2192 387 2194 410
rect 2288 387 2290 410
rect 2384 387 2386 410
rect 2456 387 2458 410
rect 2504 387 2506 411
rect 1327 386 1331 387
rect 1327 381 1331 382
rect 1599 386 1603 387
rect 1599 381 1603 382
rect 1655 386 1659 387
rect 1655 381 1659 382
rect 1679 386 1683 387
rect 1679 381 1683 382
rect 1711 386 1715 387
rect 1711 381 1715 382
rect 1735 386 1739 387
rect 1735 381 1739 382
rect 1775 386 1779 387
rect 1775 381 1779 382
rect 1799 386 1803 387
rect 1799 381 1803 382
rect 1847 386 1851 387
rect 1847 381 1851 382
rect 1871 386 1875 387
rect 1871 381 1875 382
rect 1927 386 1931 387
rect 1927 381 1931 382
rect 1943 386 1947 387
rect 1943 381 1947 382
rect 2007 386 2011 387
rect 2007 381 2011 382
rect 2023 386 2027 387
rect 2023 381 2027 382
rect 2095 386 2099 387
rect 2095 381 2099 382
rect 2111 386 2115 387
rect 2111 381 2115 382
rect 2191 386 2195 387
rect 2191 381 2195 382
rect 2199 386 2203 387
rect 2199 381 2203 382
rect 2287 386 2291 387
rect 2287 381 2291 382
rect 2375 386 2379 387
rect 2375 381 2379 382
rect 2383 386 2387 387
rect 2383 381 2387 382
rect 2455 386 2459 387
rect 2455 381 2459 382
rect 2503 386 2507 387
rect 2503 381 2507 382
rect 111 374 115 375
rect 111 369 115 370
rect 151 374 155 375
rect 151 369 155 370
rect 207 374 211 375
rect 207 369 211 370
rect 231 374 235 375
rect 231 369 235 370
rect 295 374 299 375
rect 295 369 299 370
rect 335 374 339 375
rect 335 369 339 370
rect 399 374 403 375
rect 399 369 403 370
rect 439 374 443 375
rect 439 369 443 370
rect 511 374 515 375
rect 511 369 515 370
rect 543 374 547 375
rect 543 369 547 370
rect 623 374 627 375
rect 623 369 627 370
rect 647 374 651 375
rect 647 369 651 370
rect 735 374 739 375
rect 735 369 739 370
rect 751 374 755 375
rect 751 369 755 370
rect 847 374 851 375
rect 847 369 851 370
rect 935 374 939 375
rect 935 369 939 370
rect 951 374 955 375
rect 951 369 955 370
rect 1015 374 1019 375
rect 1015 369 1019 370
rect 1055 374 1059 375
rect 1055 369 1059 370
rect 1095 374 1099 375
rect 1095 369 1099 370
rect 1159 374 1163 375
rect 1159 369 1163 370
rect 1175 374 1179 375
rect 1175 369 1179 370
rect 1239 374 1243 375
rect 1239 369 1243 370
rect 1287 374 1291 375
rect 1287 369 1291 370
rect 112 349 114 369
rect 152 350 154 369
rect 232 350 234 369
rect 336 350 338 369
rect 440 350 442 369
rect 544 350 546 369
rect 648 350 650 369
rect 752 350 754 369
rect 848 350 850 369
rect 936 350 938 369
rect 1016 350 1018 369
rect 1096 350 1098 369
rect 1176 350 1178 369
rect 1240 350 1242 369
rect 150 349 156 350
rect 110 348 116 349
rect 110 344 111 348
rect 115 344 116 348
rect 150 345 151 349
rect 155 345 156 349
rect 150 344 156 345
rect 230 349 236 350
rect 230 345 231 349
rect 235 345 236 349
rect 230 344 236 345
rect 334 349 340 350
rect 334 345 335 349
rect 339 345 340 349
rect 334 344 340 345
rect 438 349 444 350
rect 438 345 439 349
rect 443 345 444 349
rect 438 344 444 345
rect 542 349 548 350
rect 542 345 543 349
rect 547 345 548 349
rect 542 344 548 345
rect 646 349 652 350
rect 646 345 647 349
rect 651 345 652 349
rect 646 344 652 345
rect 750 349 756 350
rect 750 345 751 349
rect 755 345 756 349
rect 750 344 756 345
rect 846 349 852 350
rect 846 345 847 349
rect 851 345 852 349
rect 846 344 852 345
rect 934 349 940 350
rect 934 345 935 349
rect 939 345 940 349
rect 934 344 940 345
rect 1014 349 1020 350
rect 1014 345 1015 349
rect 1019 345 1020 349
rect 1014 344 1020 345
rect 1094 349 1100 350
rect 1094 345 1095 349
rect 1099 345 1100 349
rect 1094 344 1100 345
rect 1174 349 1180 350
rect 1174 345 1175 349
rect 1179 345 1180 349
rect 1174 344 1180 345
rect 1238 349 1244 350
rect 1288 349 1290 369
rect 1328 361 1330 381
rect 1680 362 1682 381
rect 1736 362 1738 381
rect 1800 362 1802 381
rect 1872 362 1874 381
rect 1944 362 1946 381
rect 2024 362 2026 381
rect 2112 362 2114 381
rect 2200 362 2202 381
rect 2288 362 2290 381
rect 2376 362 2378 381
rect 2456 362 2458 381
rect 1678 361 1684 362
rect 1326 360 1332 361
rect 1326 356 1327 360
rect 1331 356 1332 360
rect 1678 357 1679 361
rect 1683 357 1684 361
rect 1678 356 1684 357
rect 1734 361 1740 362
rect 1734 357 1735 361
rect 1739 357 1740 361
rect 1734 356 1740 357
rect 1798 361 1804 362
rect 1798 357 1799 361
rect 1803 357 1804 361
rect 1798 356 1804 357
rect 1870 361 1876 362
rect 1870 357 1871 361
rect 1875 357 1876 361
rect 1870 356 1876 357
rect 1942 361 1948 362
rect 1942 357 1943 361
rect 1947 357 1948 361
rect 1942 356 1948 357
rect 2022 361 2028 362
rect 2022 357 2023 361
rect 2027 357 2028 361
rect 2022 356 2028 357
rect 2110 361 2116 362
rect 2110 357 2111 361
rect 2115 357 2116 361
rect 2110 356 2116 357
rect 2198 361 2204 362
rect 2198 357 2199 361
rect 2203 357 2204 361
rect 2198 356 2204 357
rect 2286 361 2292 362
rect 2286 357 2287 361
rect 2291 357 2292 361
rect 2286 356 2292 357
rect 2374 361 2380 362
rect 2374 357 2375 361
rect 2379 357 2380 361
rect 2374 356 2380 357
rect 2454 361 2460 362
rect 2504 361 2506 381
rect 2454 357 2455 361
rect 2459 357 2460 361
rect 2454 356 2460 357
rect 2502 360 2508 361
rect 2502 356 2503 360
rect 2507 356 2508 360
rect 1326 355 1332 356
rect 2502 355 2508 356
rect 1238 345 1239 349
rect 1243 345 1244 349
rect 1238 344 1244 345
rect 1286 348 1292 349
rect 1286 344 1287 348
rect 1291 344 1292 348
rect 110 343 116 344
rect 1286 343 1292 344
rect 1326 343 1332 344
rect 1326 339 1327 343
rect 1331 339 1332 343
rect 2502 343 2508 344
rect 1326 338 1332 339
rect 1662 340 1668 341
rect 110 331 116 332
rect 110 327 111 331
rect 115 327 116 331
rect 1286 331 1292 332
rect 110 326 116 327
rect 134 328 140 329
rect 112 319 114 326
rect 134 324 135 328
rect 139 324 140 328
rect 134 323 140 324
rect 214 328 220 329
rect 214 324 215 328
rect 219 324 220 328
rect 214 323 220 324
rect 318 328 324 329
rect 318 324 319 328
rect 323 324 324 328
rect 318 323 324 324
rect 422 328 428 329
rect 422 324 423 328
rect 427 324 428 328
rect 422 323 428 324
rect 526 328 532 329
rect 526 324 527 328
rect 531 324 532 328
rect 526 323 532 324
rect 630 328 636 329
rect 630 324 631 328
rect 635 324 636 328
rect 630 323 636 324
rect 734 328 740 329
rect 734 324 735 328
rect 739 324 740 328
rect 734 323 740 324
rect 830 328 836 329
rect 830 324 831 328
rect 835 324 836 328
rect 830 323 836 324
rect 918 328 924 329
rect 918 324 919 328
rect 923 324 924 328
rect 918 323 924 324
rect 998 328 1004 329
rect 998 324 999 328
rect 1003 324 1004 328
rect 998 323 1004 324
rect 1078 328 1084 329
rect 1078 324 1079 328
rect 1083 324 1084 328
rect 1078 323 1084 324
rect 1158 328 1164 329
rect 1158 324 1159 328
rect 1163 324 1164 328
rect 1158 323 1164 324
rect 1222 328 1228 329
rect 1222 324 1223 328
rect 1227 324 1228 328
rect 1286 327 1287 331
rect 1291 327 1292 331
rect 1328 327 1330 338
rect 1662 336 1663 340
rect 1667 336 1668 340
rect 1662 335 1668 336
rect 1718 340 1724 341
rect 1718 336 1719 340
rect 1723 336 1724 340
rect 1718 335 1724 336
rect 1782 340 1788 341
rect 1782 336 1783 340
rect 1787 336 1788 340
rect 1782 335 1788 336
rect 1854 340 1860 341
rect 1854 336 1855 340
rect 1859 336 1860 340
rect 1854 335 1860 336
rect 1926 340 1932 341
rect 1926 336 1927 340
rect 1931 336 1932 340
rect 1926 335 1932 336
rect 2006 340 2012 341
rect 2006 336 2007 340
rect 2011 336 2012 340
rect 2006 335 2012 336
rect 2094 340 2100 341
rect 2094 336 2095 340
rect 2099 336 2100 340
rect 2094 335 2100 336
rect 2182 340 2188 341
rect 2182 336 2183 340
rect 2187 336 2188 340
rect 2182 335 2188 336
rect 2270 340 2276 341
rect 2270 336 2271 340
rect 2275 336 2276 340
rect 2270 335 2276 336
rect 2358 340 2364 341
rect 2358 336 2359 340
rect 2363 336 2364 340
rect 2358 335 2364 336
rect 2438 340 2444 341
rect 2438 336 2439 340
rect 2443 336 2444 340
rect 2502 339 2503 343
rect 2507 339 2508 343
rect 2502 338 2508 339
rect 2438 335 2444 336
rect 1664 327 1666 335
rect 1720 327 1722 335
rect 1784 327 1786 335
rect 1856 327 1858 335
rect 1928 327 1930 335
rect 2008 327 2010 335
rect 2096 327 2098 335
rect 2184 327 2186 335
rect 2272 327 2274 335
rect 2360 327 2362 335
rect 2440 327 2442 335
rect 2504 327 2506 338
rect 1286 326 1292 327
rect 1327 326 1331 327
rect 1222 323 1228 324
rect 136 319 138 323
rect 216 319 218 323
rect 320 319 322 323
rect 424 319 426 323
rect 528 319 530 323
rect 632 319 634 323
rect 736 319 738 323
rect 832 319 834 323
rect 920 319 922 323
rect 1000 319 1002 323
rect 1080 319 1082 323
rect 1160 319 1162 323
rect 1224 319 1226 323
rect 1288 319 1290 326
rect 1327 321 1331 322
rect 1351 326 1355 327
rect 1351 321 1355 322
rect 1455 326 1459 327
rect 1455 321 1459 322
rect 1583 326 1587 327
rect 1583 321 1587 322
rect 1663 326 1667 327
rect 1663 321 1667 322
rect 1711 326 1715 327
rect 1711 321 1715 322
rect 1719 326 1723 327
rect 1719 321 1723 322
rect 1783 326 1787 327
rect 1783 321 1787 322
rect 1839 326 1843 327
rect 1839 321 1843 322
rect 1855 326 1859 327
rect 1855 321 1859 322
rect 1927 326 1931 327
rect 1927 321 1931 322
rect 1951 326 1955 327
rect 1951 321 1955 322
rect 2007 326 2011 327
rect 2007 321 2011 322
rect 2063 326 2067 327
rect 2063 321 2067 322
rect 2095 326 2099 327
rect 2095 321 2099 322
rect 2167 326 2171 327
rect 2167 321 2171 322
rect 2183 326 2187 327
rect 2183 321 2187 322
rect 2263 326 2267 327
rect 2263 321 2267 322
rect 2271 326 2275 327
rect 2271 321 2275 322
rect 2359 326 2363 327
rect 2359 321 2363 322
rect 2439 326 2443 327
rect 2439 321 2443 322
rect 2503 326 2507 327
rect 2503 321 2507 322
rect 111 318 115 319
rect 111 313 115 314
rect 135 318 139 319
rect 135 313 139 314
rect 215 318 219 319
rect 215 313 219 314
rect 319 318 323 319
rect 319 313 323 314
rect 423 318 427 319
rect 423 313 427 314
rect 527 318 531 319
rect 527 313 531 314
rect 535 318 539 319
rect 535 313 539 314
rect 631 318 635 319
rect 631 313 635 314
rect 639 318 643 319
rect 639 313 643 314
rect 735 318 739 319
rect 735 313 739 314
rect 743 318 747 319
rect 743 313 747 314
rect 831 318 835 319
rect 831 313 835 314
rect 847 318 851 319
rect 847 313 851 314
rect 919 318 923 319
rect 919 313 923 314
rect 943 318 947 319
rect 943 313 947 314
rect 999 318 1003 319
rect 999 313 1003 314
rect 1039 318 1043 319
rect 1039 313 1043 314
rect 1079 318 1083 319
rect 1079 313 1083 314
rect 1143 318 1147 319
rect 1143 313 1147 314
rect 1159 318 1163 319
rect 1159 313 1163 314
rect 1223 318 1227 319
rect 1223 313 1227 314
rect 1287 318 1291 319
rect 1328 318 1330 321
rect 1350 320 1356 321
rect 1287 313 1291 314
rect 1326 317 1332 318
rect 1326 313 1327 317
rect 1331 313 1332 317
rect 1350 316 1351 320
rect 1355 316 1356 320
rect 1350 315 1356 316
rect 1454 320 1460 321
rect 1454 316 1455 320
rect 1459 316 1460 320
rect 1454 315 1460 316
rect 1582 320 1588 321
rect 1582 316 1583 320
rect 1587 316 1588 320
rect 1582 315 1588 316
rect 1710 320 1716 321
rect 1710 316 1711 320
rect 1715 316 1716 320
rect 1710 315 1716 316
rect 1838 320 1844 321
rect 1838 316 1839 320
rect 1843 316 1844 320
rect 1838 315 1844 316
rect 1950 320 1956 321
rect 1950 316 1951 320
rect 1955 316 1956 320
rect 1950 315 1956 316
rect 2062 320 2068 321
rect 2062 316 2063 320
rect 2067 316 2068 320
rect 2062 315 2068 316
rect 2166 320 2172 321
rect 2166 316 2167 320
rect 2171 316 2172 320
rect 2166 315 2172 316
rect 2262 320 2268 321
rect 2262 316 2263 320
rect 2267 316 2268 320
rect 2262 315 2268 316
rect 2358 320 2364 321
rect 2358 316 2359 320
rect 2363 316 2364 320
rect 2358 315 2364 316
rect 2438 320 2444 321
rect 2438 316 2439 320
rect 2443 316 2444 320
rect 2504 318 2506 321
rect 2438 315 2444 316
rect 2502 317 2508 318
rect 112 310 114 313
rect 134 312 140 313
rect 110 309 116 310
rect 110 305 111 309
rect 115 305 116 309
rect 134 308 135 312
rect 139 308 140 312
rect 134 307 140 308
rect 214 312 220 313
rect 214 308 215 312
rect 219 308 220 312
rect 214 307 220 308
rect 318 312 324 313
rect 318 308 319 312
rect 323 308 324 312
rect 318 307 324 308
rect 422 312 428 313
rect 422 308 423 312
rect 427 308 428 312
rect 422 307 428 308
rect 534 312 540 313
rect 534 308 535 312
rect 539 308 540 312
rect 534 307 540 308
rect 638 312 644 313
rect 638 308 639 312
rect 643 308 644 312
rect 638 307 644 308
rect 742 312 748 313
rect 742 308 743 312
rect 747 308 748 312
rect 742 307 748 308
rect 846 312 852 313
rect 846 308 847 312
rect 851 308 852 312
rect 846 307 852 308
rect 942 312 948 313
rect 942 308 943 312
rect 947 308 948 312
rect 942 307 948 308
rect 1038 312 1044 313
rect 1038 308 1039 312
rect 1043 308 1044 312
rect 1038 307 1044 308
rect 1142 312 1148 313
rect 1142 308 1143 312
rect 1147 308 1148 312
rect 1142 307 1148 308
rect 1222 312 1228 313
rect 1222 308 1223 312
rect 1227 308 1228 312
rect 1288 310 1290 313
rect 1326 312 1332 313
rect 2502 313 2503 317
rect 2507 313 2508 317
rect 2502 312 2508 313
rect 1222 307 1228 308
rect 1286 309 1292 310
rect 110 304 116 305
rect 1286 305 1287 309
rect 1291 305 1292 309
rect 1286 304 1292 305
rect 1326 300 1332 301
rect 2502 300 2508 301
rect 1326 296 1327 300
rect 1331 296 1332 300
rect 1326 295 1332 296
rect 1366 299 1372 300
rect 1366 295 1367 299
rect 1371 295 1372 299
rect 110 292 116 293
rect 1286 292 1292 293
rect 110 288 111 292
rect 115 288 116 292
rect 110 287 116 288
rect 150 291 156 292
rect 150 287 151 291
rect 155 287 156 291
rect 112 267 114 287
rect 150 286 156 287
rect 230 291 236 292
rect 230 287 231 291
rect 235 287 236 291
rect 230 286 236 287
rect 334 291 340 292
rect 334 287 335 291
rect 339 287 340 291
rect 334 286 340 287
rect 438 291 444 292
rect 438 287 439 291
rect 443 287 444 291
rect 438 286 444 287
rect 550 291 556 292
rect 550 287 551 291
rect 555 287 556 291
rect 550 286 556 287
rect 654 291 660 292
rect 654 287 655 291
rect 659 287 660 291
rect 654 286 660 287
rect 758 291 764 292
rect 758 287 759 291
rect 763 287 764 291
rect 758 286 764 287
rect 862 291 868 292
rect 862 287 863 291
rect 867 287 868 291
rect 862 286 868 287
rect 958 291 964 292
rect 958 287 959 291
rect 963 287 964 291
rect 958 286 964 287
rect 1054 291 1060 292
rect 1054 287 1055 291
rect 1059 287 1060 291
rect 1054 286 1060 287
rect 1158 291 1164 292
rect 1158 287 1159 291
rect 1163 287 1164 291
rect 1158 286 1164 287
rect 1238 291 1244 292
rect 1238 287 1239 291
rect 1243 287 1244 291
rect 1286 288 1287 292
rect 1291 288 1292 292
rect 1286 287 1292 288
rect 1238 286 1244 287
rect 152 267 154 286
rect 232 267 234 286
rect 336 267 338 286
rect 440 267 442 286
rect 552 267 554 286
rect 656 267 658 286
rect 760 267 762 286
rect 864 267 866 286
rect 960 267 962 286
rect 1056 267 1058 286
rect 1160 267 1162 286
rect 1240 267 1242 286
rect 1288 267 1290 287
rect 1328 267 1330 295
rect 1366 294 1372 295
rect 1470 299 1476 300
rect 1470 295 1471 299
rect 1475 295 1476 299
rect 1470 294 1476 295
rect 1598 299 1604 300
rect 1598 295 1599 299
rect 1603 295 1604 299
rect 1598 294 1604 295
rect 1726 299 1732 300
rect 1726 295 1727 299
rect 1731 295 1732 299
rect 1726 294 1732 295
rect 1854 299 1860 300
rect 1854 295 1855 299
rect 1859 295 1860 299
rect 1854 294 1860 295
rect 1966 299 1972 300
rect 1966 295 1967 299
rect 1971 295 1972 299
rect 1966 294 1972 295
rect 2078 299 2084 300
rect 2078 295 2079 299
rect 2083 295 2084 299
rect 2078 294 2084 295
rect 2182 299 2188 300
rect 2182 295 2183 299
rect 2187 295 2188 299
rect 2182 294 2188 295
rect 2278 299 2284 300
rect 2278 295 2279 299
rect 2283 295 2284 299
rect 2278 294 2284 295
rect 2374 299 2380 300
rect 2374 295 2375 299
rect 2379 295 2380 299
rect 2374 294 2380 295
rect 2454 299 2460 300
rect 2454 295 2455 299
rect 2459 295 2460 299
rect 2502 296 2503 300
rect 2507 296 2508 300
rect 2502 295 2508 296
rect 2454 294 2460 295
rect 1368 267 1370 294
rect 1472 267 1474 294
rect 1600 267 1602 294
rect 1728 267 1730 294
rect 1856 267 1858 294
rect 1968 267 1970 294
rect 2080 267 2082 294
rect 2184 267 2186 294
rect 2280 267 2282 294
rect 2376 267 2378 294
rect 2456 267 2458 294
rect 2504 267 2506 295
rect 111 266 115 267
rect 111 261 115 262
rect 151 266 155 267
rect 151 261 155 262
rect 223 266 227 267
rect 223 261 227 262
rect 231 266 235 267
rect 231 261 235 262
rect 319 266 323 267
rect 319 261 323 262
rect 335 266 339 267
rect 335 261 339 262
rect 423 266 427 267
rect 423 261 427 262
rect 439 266 443 267
rect 439 261 443 262
rect 535 266 539 267
rect 535 261 539 262
rect 551 266 555 267
rect 551 261 555 262
rect 647 266 651 267
rect 647 261 651 262
rect 655 266 659 267
rect 655 261 659 262
rect 759 266 763 267
rect 759 261 763 262
rect 863 266 867 267
rect 863 261 867 262
rect 871 266 875 267
rect 871 261 875 262
rect 959 266 963 267
rect 959 261 963 262
rect 983 266 987 267
rect 983 261 987 262
rect 1055 266 1059 267
rect 1055 261 1059 262
rect 1103 266 1107 267
rect 1103 261 1107 262
rect 1159 266 1163 267
rect 1159 261 1163 262
rect 1223 266 1227 267
rect 1223 261 1227 262
rect 1239 266 1243 267
rect 1239 261 1243 262
rect 1287 266 1291 267
rect 1287 261 1291 262
rect 1327 266 1331 267
rect 1327 261 1331 262
rect 1367 266 1371 267
rect 1367 261 1371 262
rect 1447 266 1451 267
rect 1447 261 1451 262
rect 1471 266 1475 267
rect 1471 261 1475 262
rect 1551 266 1555 267
rect 1551 261 1555 262
rect 1599 266 1603 267
rect 1599 261 1603 262
rect 1655 266 1659 267
rect 1655 261 1659 262
rect 1727 266 1731 267
rect 1727 261 1731 262
rect 1759 266 1763 267
rect 1759 261 1763 262
rect 1855 266 1859 267
rect 1855 261 1859 262
rect 1863 266 1867 267
rect 1863 261 1867 262
rect 1967 266 1971 267
rect 1967 261 1971 262
rect 2071 266 2075 267
rect 2071 261 2075 262
rect 2079 266 2083 267
rect 2079 261 2083 262
rect 2175 266 2179 267
rect 2175 261 2179 262
rect 2183 266 2187 267
rect 2183 261 2187 262
rect 2271 266 2275 267
rect 2271 261 2275 262
rect 2279 266 2283 267
rect 2279 261 2283 262
rect 2375 266 2379 267
rect 2375 261 2379 262
rect 2455 266 2459 267
rect 2455 261 2459 262
rect 2503 266 2507 267
rect 2503 261 2507 262
rect 112 241 114 261
rect 152 242 154 261
rect 224 242 226 261
rect 320 242 322 261
rect 424 242 426 261
rect 536 242 538 261
rect 648 242 650 261
rect 760 242 762 261
rect 872 242 874 261
rect 984 242 986 261
rect 1104 242 1106 261
rect 1224 242 1226 261
rect 150 241 156 242
rect 110 240 116 241
rect 110 236 111 240
rect 115 236 116 240
rect 150 237 151 241
rect 155 237 156 241
rect 150 236 156 237
rect 222 241 228 242
rect 222 237 223 241
rect 227 237 228 241
rect 222 236 228 237
rect 318 241 324 242
rect 318 237 319 241
rect 323 237 324 241
rect 318 236 324 237
rect 422 241 428 242
rect 422 237 423 241
rect 427 237 428 241
rect 422 236 428 237
rect 534 241 540 242
rect 534 237 535 241
rect 539 237 540 241
rect 534 236 540 237
rect 646 241 652 242
rect 646 237 647 241
rect 651 237 652 241
rect 646 236 652 237
rect 758 241 764 242
rect 758 237 759 241
rect 763 237 764 241
rect 758 236 764 237
rect 870 241 876 242
rect 870 237 871 241
rect 875 237 876 241
rect 870 236 876 237
rect 982 241 988 242
rect 982 237 983 241
rect 987 237 988 241
rect 982 236 988 237
rect 1102 241 1108 242
rect 1102 237 1103 241
rect 1107 237 1108 241
rect 1102 236 1108 237
rect 1222 241 1228 242
rect 1288 241 1290 261
rect 1328 241 1330 261
rect 1368 242 1370 261
rect 1448 242 1450 261
rect 1552 242 1554 261
rect 1656 242 1658 261
rect 1760 242 1762 261
rect 1864 242 1866 261
rect 1968 242 1970 261
rect 2072 242 2074 261
rect 2176 242 2178 261
rect 2272 242 2274 261
rect 2376 242 2378 261
rect 2456 242 2458 261
rect 1366 241 1372 242
rect 1222 237 1223 241
rect 1227 237 1228 241
rect 1222 236 1228 237
rect 1286 240 1292 241
rect 1286 236 1287 240
rect 1291 236 1292 240
rect 110 235 116 236
rect 1286 235 1292 236
rect 1326 240 1332 241
rect 1326 236 1327 240
rect 1331 236 1332 240
rect 1366 237 1367 241
rect 1371 237 1372 241
rect 1366 236 1372 237
rect 1446 241 1452 242
rect 1446 237 1447 241
rect 1451 237 1452 241
rect 1446 236 1452 237
rect 1550 241 1556 242
rect 1550 237 1551 241
rect 1555 237 1556 241
rect 1550 236 1556 237
rect 1654 241 1660 242
rect 1654 237 1655 241
rect 1659 237 1660 241
rect 1654 236 1660 237
rect 1758 241 1764 242
rect 1758 237 1759 241
rect 1763 237 1764 241
rect 1758 236 1764 237
rect 1862 241 1868 242
rect 1862 237 1863 241
rect 1867 237 1868 241
rect 1862 236 1868 237
rect 1966 241 1972 242
rect 1966 237 1967 241
rect 1971 237 1972 241
rect 1966 236 1972 237
rect 2070 241 2076 242
rect 2070 237 2071 241
rect 2075 237 2076 241
rect 2070 236 2076 237
rect 2174 241 2180 242
rect 2174 237 2175 241
rect 2179 237 2180 241
rect 2174 236 2180 237
rect 2270 241 2276 242
rect 2270 237 2271 241
rect 2275 237 2276 241
rect 2270 236 2276 237
rect 2374 241 2380 242
rect 2374 237 2375 241
rect 2379 237 2380 241
rect 2374 236 2380 237
rect 2454 241 2460 242
rect 2504 241 2506 261
rect 2454 237 2455 241
rect 2459 237 2460 241
rect 2454 236 2460 237
rect 2502 240 2508 241
rect 2502 236 2503 240
rect 2507 236 2508 240
rect 1326 235 1332 236
rect 2502 235 2508 236
rect 110 223 116 224
rect 110 219 111 223
rect 115 219 116 223
rect 1286 223 1292 224
rect 110 218 116 219
rect 134 220 140 221
rect 112 211 114 218
rect 134 216 135 220
rect 139 216 140 220
rect 134 215 140 216
rect 206 220 212 221
rect 206 216 207 220
rect 211 216 212 220
rect 206 215 212 216
rect 302 220 308 221
rect 302 216 303 220
rect 307 216 308 220
rect 302 215 308 216
rect 406 220 412 221
rect 406 216 407 220
rect 411 216 412 220
rect 406 215 412 216
rect 518 220 524 221
rect 518 216 519 220
rect 523 216 524 220
rect 518 215 524 216
rect 630 220 636 221
rect 630 216 631 220
rect 635 216 636 220
rect 630 215 636 216
rect 742 220 748 221
rect 742 216 743 220
rect 747 216 748 220
rect 742 215 748 216
rect 854 220 860 221
rect 854 216 855 220
rect 859 216 860 220
rect 854 215 860 216
rect 966 220 972 221
rect 966 216 967 220
rect 971 216 972 220
rect 966 215 972 216
rect 1086 220 1092 221
rect 1086 216 1087 220
rect 1091 216 1092 220
rect 1086 215 1092 216
rect 1206 220 1212 221
rect 1206 216 1207 220
rect 1211 216 1212 220
rect 1286 219 1287 223
rect 1291 219 1292 223
rect 1286 218 1292 219
rect 1326 223 1332 224
rect 1326 219 1327 223
rect 1331 219 1332 223
rect 2502 223 2508 224
rect 1326 218 1332 219
rect 1350 220 1356 221
rect 1206 215 1212 216
rect 136 211 138 215
rect 208 211 210 215
rect 304 211 306 215
rect 408 211 410 215
rect 520 211 522 215
rect 632 211 634 215
rect 744 211 746 215
rect 856 211 858 215
rect 968 211 970 215
rect 1088 211 1090 215
rect 1208 211 1210 215
rect 1288 211 1290 218
rect 1328 211 1330 218
rect 1350 216 1351 220
rect 1355 216 1356 220
rect 1350 215 1356 216
rect 1430 220 1436 221
rect 1430 216 1431 220
rect 1435 216 1436 220
rect 1430 215 1436 216
rect 1534 220 1540 221
rect 1534 216 1535 220
rect 1539 216 1540 220
rect 1534 215 1540 216
rect 1638 220 1644 221
rect 1638 216 1639 220
rect 1643 216 1644 220
rect 1638 215 1644 216
rect 1742 220 1748 221
rect 1742 216 1743 220
rect 1747 216 1748 220
rect 1742 215 1748 216
rect 1846 220 1852 221
rect 1846 216 1847 220
rect 1851 216 1852 220
rect 1846 215 1852 216
rect 1950 220 1956 221
rect 1950 216 1951 220
rect 1955 216 1956 220
rect 1950 215 1956 216
rect 2054 220 2060 221
rect 2054 216 2055 220
rect 2059 216 2060 220
rect 2054 215 2060 216
rect 2158 220 2164 221
rect 2158 216 2159 220
rect 2163 216 2164 220
rect 2158 215 2164 216
rect 2254 220 2260 221
rect 2254 216 2255 220
rect 2259 216 2260 220
rect 2254 215 2260 216
rect 2358 220 2364 221
rect 2358 216 2359 220
rect 2363 216 2364 220
rect 2358 215 2364 216
rect 2438 220 2444 221
rect 2438 216 2439 220
rect 2443 216 2444 220
rect 2502 219 2503 223
rect 2507 219 2508 223
rect 2502 218 2508 219
rect 2438 215 2444 216
rect 1352 211 1354 215
rect 1432 211 1434 215
rect 1536 211 1538 215
rect 1640 211 1642 215
rect 1744 211 1746 215
rect 1848 211 1850 215
rect 1952 211 1954 215
rect 2056 211 2058 215
rect 2160 211 2162 215
rect 2256 211 2258 215
rect 2360 211 2362 215
rect 2440 211 2442 215
rect 2504 211 2506 218
rect 111 210 115 211
rect 111 205 115 206
rect 135 210 139 211
rect 135 205 139 206
rect 183 210 187 211
rect 183 205 187 206
rect 207 210 211 211
rect 207 205 211 206
rect 279 210 283 211
rect 279 205 283 206
rect 303 210 307 211
rect 303 205 307 206
rect 383 210 387 211
rect 383 205 387 206
rect 407 210 411 211
rect 407 205 411 206
rect 487 210 491 211
rect 487 205 491 206
rect 519 210 523 211
rect 519 205 523 206
rect 591 210 595 211
rect 591 205 595 206
rect 631 210 635 211
rect 631 205 635 206
rect 695 210 699 211
rect 695 205 699 206
rect 743 210 747 211
rect 743 205 747 206
rect 799 210 803 211
rect 799 205 803 206
rect 855 210 859 211
rect 855 205 859 206
rect 895 210 899 211
rect 895 205 899 206
rect 967 210 971 211
rect 967 205 971 206
rect 999 210 1003 211
rect 999 205 1003 206
rect 1087 210 1091 211
rect 1087 205 1091 206
rect 1103 210 1107 211
rect 1103 205 1107 206
rect 1207 210 1211 211
rect 1207 205 1211 206
rect 1287 210 1291 211
rect 1287 205 1291 206
rect 1327 210 1331 211
rect 1327 205 1331 206
rect 1351 210 1355 211
rect 1351 205 1355 206
rect 1407 210 1411 211
rect 1407 205 1411 206
rect 1431 210 1435 211
rect 1431 205 1435 206
rect 1471 210 1475 211
rect 1471 205 1475 206
rect 1535 210 1539 211
rect 1535 205 1539 206
rect 1551 210 1555 211
rect 1551 205 1555 206
rect 1639 210 1643 211
rect 1639 205 1643 206
rect 1719 210 1723 211
rect 1719 205 1723 206
rect 1743 210 1747 211
rect 1743 205 1747 206
rect 1807 210 1811 211
rect 1807 205 1811 206
rect 1847 210 1851 211
rect 1847 205 1851 206
rect 1895 210 1899 211
rect 1895 205 1899 206
rect 1951 210 1955 211
rect 1951 205 1955 206
rect 1991 210 1995 211
rect 1991 205 1995 206
rect 2055 210 2059 211
rect 2055 205 2059 206
rect 2103 210 2107 211
rect 2103 205 2107 206
rect 2159 210 2163 211
rect 2159 205 2163 206
rect 2215 210 2219 211
rect 2215 205 2219 206
rect 2255 210 2259 211
rect 2255 205 2259 206
rect 2335 210 2339 211
rect 2335 205 2339 206
rect 2359 210 2363 211
rect 2359 205 2363 206
rect 2439 210 2443 211
rect 2439 205 2443 206
rect 2503 210 2507 211
rect 2503 205 2507 206
rect 112 202 114 205
rect 182 204 188 205
rect 110 201 116 202
rect 110 197 111 201
rect 115 197 116 201
rect 182 200 183 204
rect 187 200 188 204
rect 182 199 188 200
rect 278 204 284 205
rect 278 200 279 204
rect 283 200 284 204
rect 278 199 284 200
rect 382 204 388 205
rect 382 200 383 204
rect 387 200 388 204
rect 382 199 388 200
rect 486 204 492 205
rect 486 200 487 204
rect 491 200 492 204
rect 486 199 492 200
rect 590 204 596 205
rect 590 200 591 204
rect 595 200 596 204
rect 590 199 596 200
rect 694 204 700 205
rect 694 200 695 204
rect 699 200 700 204
rect 694 199 700 200
rect 798 204 804 205
rect 798 200 799 204
rect 803 200 804 204
rect 798 199 804 200
rect 894 204 900 205
rect 894 200 895 204
rect 899 200 900 204
rect 894 199 900 200
rect 998 204 1004 205
rect 998 200 999 204
rect 1003 200 1004 204
rect 998 199 1004 200
rect 1102 204 1108 205
rect 1102 200 1103 204
rect 1107 200 1108 204
rect 1288 202 1290 205
rect 1328 202 1330 205
rect 1350 204 1356 205
rect 1102 199 1108 200
rect 1286 201 1292 202
rect 110 196 116 197
rect 1286 197 1287 201
rect 1291 197 1292 201
rect 1286 196 1292 197
rect 1326 201 1332 202
rect 1326 197 1327 201
rect 1331 197 1332 201
rect 1350 200 1351 204
rect 1355 200 1356 204
rect 1350 199 1356 200
rect 1406 204 1412 205
rect 1406 200 1407 204
rect 1411 200 1412 204
rect 1406 199 1412 200
rect 1470 204 1476 205
rect 1470 200 1471 204
rect 1475 200 1476 204
rect 1470 199 1476 200
rect 1550 204 1556 205
rect 1550 200 1551 204
rect 1555 200 1556 204
rect 1550 199 1556 200
rect 1638 204 1644 205
rect 1638 200 1639 204
rect 1643 200 1644 204
rect 1638 199 1644 200
rect 1718 204 1724 205
rect 1718 200 1719 204
rect 1723 200 1724 204
rect 1718 199 1724 200
rect 1806 204 1812 205
rect 1806 200 1807 204
rect 1811 200 1812 204
rect 1806 199 1812 200
rect 1894 204 1900 205
rect 1894 200 1895 204
rect 1899 200 1900 204
rect 1894 199 1900 200
rect 1990 204 1996 205
rect 1990 200 1991 204
rect 1995 200 1996 204
rect 1990 199 1996 200
rect 2102 204 2108 205
rect 2102 200 2103 204
rect 2107 200 2108 204
rect 2102 199 2108 200
rect 2214 204 2220 205
rect 2214 200 2215 204
rect 2219 200 2220 204
rect 2214 199 2220 200
rect 2334 204 2340 205
rect 2334 200 2335 204
rect 2339 200 2340 204
rect 2334 199 2340 200
rect 2438 204 2444 205
rect 2438 200 2439 204
rect 2443 200 2444 204
rect 2504 202 2506 205
rect 2438 199 2444 200
rect 2502 201 2508 202
rect 1326 196 1332 197
rect 2502 197 2503 201
rect 2507 197 2508 201
rect 2502 196 2508 197
rect 110 184 116 185
rect 1286 184 1292 185
rect 110 180 111 184
rect 115 180 116 184
rect 110 179 116 180
rect 198 183 204 184
rect 198 179 199 183
rect 203 179 204 183
rect 112 151 114 179
rect 198 178 204 179
rect 294 183 300 184
rect 294 179 295 183
rect 299 179 300 183
rect 294 178 300 179
rect 398 183 404 184
rect 398 179 399 183
rect 403 179 404 183
rect 398 178 404 179
rect 502 183 508 184
rect 502 179 503 183
rect 507 179 508 183
rect 502 178 508 179
rect 606 183 612 184
rect 606 179 607 183
rect 611 179 612 183
rect 606 178 612 179
rect 710 183 716 184
rect 710 179 711 183
rect 715 179 716 183
rect 710 178 716 179
rect 814 183 820 184
rect 814 179 815 183
rect 819 179 820 183
rect 814 178 820 179
rect 910 183 916 184
rect 910 179 911 183
rect 915 179 916 183
rect 910 178 916 179
rect 1014 183 1020 184
rect 1014 179 1015 183
rect 1019 179 1020 183
rect 1014 178 1020 179
rect 1118 183 1124 184
rect 1118 179 1119 183
rect 1123 179 1124 183
rect 1286 180 1287 184
rect 1291 180 1292 184
rect 1286 179 1292 180
rect 1326 184 1332 185
rect 2502 184 2508 185
rect 1326 180 1327 184
rect 1331 180 1332 184
rect 1326 179 1332 180
rect 1366 183 1372 184
rect 1366 179 1367 183
rect 1371 179 1372 183
rect 1118 178 1124 179
rect 200 151 202 178
rect 296 151 298 178
rect 400 151 402 178
rect 504 151 506 178
rect 608 151 610 178
rect 712 151 714 178
rect 816 151 818 178
rect 912 151 914 178
rect 1016 151 1018 178
rect 1120 151 1122 178
rect 1288 151 1290 179
rect 111 150 115 151
rect 111 145 115 146
rect 151 150 155 151
rect 151 145 155 146
rect 199 150 203 151
rect 199 145 203 146
rect 207 150 211 151
rect 207 145 211 146
rect 263 150 267 151
rect 263 145 267 146
rect 295 150 299 151
rect 295 145 299 146
rect 319 150 323 151
rect 319 145 323 146
rect 375 150 379 151
rect 375 145 379 146
rect 399 150 403 151
rect 399 145 403 146
rect 431 150 435 151
rect 431 145 435 146
rect 487 150 491 151
rect 487 145 491 146
rect 503 150 507 151
rect 503 145 507 146
rect 543 150 547 151
rect 543 145 547 146
rect 599 150 603 151
rect 599 145 603 146
rect 607 150 611 151
rect 607 145 611 146
rect 655 150 659 151
rect 655 145 659 146
rect 711 150 715 151
rect 711 145 715 146
rect 767 150 771 151
rect 767 145 771 146
rect 815 150 819 151
rect 815 145 819 146
rect 831 150 835 151
rect 831 145 835 146
rect 895 150 899 151
rect 895 145 899 146
rect 911 150 915 151
rect 911 145 915 146
rect 959 150 963 151
rect 959 145 963 146
rect 1015 150 1019 151
rect 1015 145 1019 146
rect 1023 150 1027 151
rect 1023 145 1027 146
rect 1087 150 1091 151
rect 1087 145 1091 146
rect 1119 150 1123 151
rect 1119 145 1123 146
rect 1151 150 1155 151
rect 1151 145 1155 146
rect 1287 150 1291 151
rect 1287 145 1291 146
rect 112 125 114 145
rect 152 126 154 145
rect 208 126 210 145
rect 264 126 266 145
rect 320 126 322 145
rect 376 126 378 145
rect 432 126 434 145
rect 488 126 490 145
rect 544 126 546 145
rect 600 126 602 145
rect 656 126 658 145
rect 712 126 714 145
rect 768 126 770 145
rect 832 126 834 145
rect 896 126 898 145
rect 960 126 962 145
rect 1024 126 1026 145
rect 1088 126 1090 145
rect 1152 126 1154 145
rect 150 125 156 126
rect 110 124 116 125
rect 110 120 111 124
rect 115 120 116 124
rect 150 121 151 125
rect 155 121 156 125
rect 150 120 156 121
rect 206 125 212 126
rect 206 121 207 125
rect 211 121 212 125
rect 206 120 212 121
rect 262 125 268 126
rect 262 121 263 125
rect 267 121 268 125
rect 262 120 268 121
rect 318 125 324 126
rect 318 121 319 125
rect 323 121 324 125
rect 318 120 324 121
rect 374 125 380 126
rect 374 121 375 125
rect 379 121 380 125
rect 374 120 380 121
rect 430 125 436 126
rect 430 121 431 125
rect 435 121 436 125
rect 430 120 436 121
rect 486 125 492 126
rect 486 121 487 125
rect 491 121 492 125
rect 486 120 492 121
rect 542 125 548 126
rect 542 121 543 125
rect 547 121 548 125
rect 542 120 548 121
rect 598 125 604 126
rect 598 121 599 125
rect 603 121 604 125
rect 598 120 604 121
rect 654 125 660 126
rect 654 121 655 125
rect 659 121 660 125
rect 654 120 660 121
rect 710 125 716 126
rect 710 121 711 125
rect 715 121 716 125
rect 710 120 716 121
rect 766 125 772 126
rect 766 121 767 125
rect 771 121 772 125
rect 766 120 772 121
rect 830 125 836 126
rect 830 121 831 125
rect 835 121 836 125
rect 830 120 836 121
rect 894 125 900 126
rect 894 121 895 125
rect 899 121 900 125
rect 894 120 900 121
rect 958 125 964 126
rect 958 121 959 125
rect 963 121 964 125
rect 958 120 964 121
rect 1022 125 1028 126
rect 1022 121 1023 125
rect 1027 121 1028 125
rect 1022 120 1028 121
rect 1086 125 1092 126
rect 1086 121 1087 125
rect 1091 121 1092 125
rect 1086 120 1092 121
rect 1150 125 1156 126
rect 1288 125 1290 145
rect 1328 139 1330 179
rect 1366 178 1372 179
rect 1422 183 1428 184
rect 1422 179 1423 183
rect 1427 179 1428 183
rect 1422 178 1428 179
rect 1486 183 1492 184
rect 1486 179 1487 183
rect 1491 179 1492 183
rect 1486 178 1492 179
rect 1566 183 1572 184
rect 1566 179 1567 183
rect 1571 179 1572 183
rect 1566 178 1572 179
rect 1654 183 1660 184
rect 1654 179 1655 183
rect 1659 179 1660 183
rect 1654 178 1660 179
rect 1734 183 1740 184
rect 1734 179 1735 183
rect 1739 179 1740 183
rect 1734 178 1740 179
rect 1822 183 1828 184
rect 1822 179 1823 183
rect 1827 179 1828 183
rect 1822 178 1828 179
rect 1910 183 1916 184
rect 1910 179 1911 183
rect 1915 179 1916 183
rect 1910 178 1916 179
rect 2006 183 2012 184
rect 2006 179 2007 183
rect 2011 179 2012 183
rect 2006 178 2012 179
rect 2118 183 2124 184
rect 2118 179 2119 183
rect 2123 179 2124 183
rect 2118 178 2124 179
rect 2230 183 2236 184
rect 2230 179 2231 183
rect 2235 179 2236 183
rect 2230 178 2236 179
rect 2350 183 2356 184
rect 2350 179 2351 183
rect 2355 179 2356 183
rect 2350 178 2356 179
rect 2454 183 2460 184
rect 2454 179 2455 183
rect 2459 179 2460 183
rect 2502 180 2503 184
rect 2507 180 2508 184
rect 2502 179 2508 180
rect 2454 178 2460 179
rect 1368 139 1370 178
rect 1424 139 1426 178
rect 1488 139 1490 178
rect 1568 139 1570 178
rect 1656 139 1658 178
rect 1736 139 1738 178
rect 1824 139 1826 178
rect 1912 139 1914 178
rect 2008 139 2010 178
rect 2120 139 2122 178
rect 2232 139 2234 178
rect 2352 139 2354 178
rect 2456 139 2458 178
rect 2504 139 2506 179
rect 1327 138 1331 139
rect 1327 133 1331 134
rect 1367 138 1371 139
rect 1367 133 1371 134
rect 1423 138 1427 139
rect 1423 133 1427 134
rect 1479 138 1483 139
rect 1479 133 1483 134
rect 1487 138 1491 139
rect 1487 133 1491 134
rect 1535 138 1539 139
rect 1535 133 1539 134
rect 1567 138 1571 139
rect 1567 133 1571 134
rect 1591 138 1595 139
rect 1591 133 1595 134
rect 1647 138 1651 139
rect 1647 133 1651 134
rect 1655 138 1659 139
rect 1655 133 1659 134
rect 1703 138 1707 139
rect 1703 133 1707 134
rect 1735 138 1739 139
rect 1735 133 1739 134
rect 1759 138 1763 139
rect 1759 133 1763 134
rect 1823 138 1827 139
rect 1823 133 1827 134
rect 1879 138 1883 139
rect 1879 133 1883 134
rect 1911 138 1915 139
rect 1911 133 1915 134
rect 1943 138 1947 139
rect 1943 133 1947 134
rect 2007 138 2011 139
rect 2007 133 2011 134
rect 2071 138 2075 139
rect 2071 133 2075 134
rect 2119 138 2123 139
rect 2119 133 2123 134
rect 2143 138 2147 139
rect 2143 133 2147 134
rect 2223 138 2227 139
rect 2223 133 2227 134
rect 2231 138 2235 139
rect 2231 133 2235 134
rect 2303 138 2307 139
rect 2303 133 2307 134
rect 2351 138 2355 139
rect 2351 133 2355 134
rect 2391 138 2395 139
rect 2391 133 2395 134
rect 2455 138 2459 139
rect 2455 133 2459 134
rect 2503 138 2507 139
rect 2503 133 2507 134
rect 1150 121 1151 125
rect 1155 121 1156 125
rect 1150 120 1156 121
rect 1286 124 1292 125
rect 1286 120 1287 124
rect 1291 120 1292 124
rect 110 119 116 120
rect 1286 119 1292 120
rect 1328 113 1330 133
rect 1368 114 1370 133
rect 1424 114 1426 133
rect 1480 114 1482 133
rect 1536 114 1538 133
rect 1592 114 1594 133
rect 1648 114 1650 133
rect 1704 114 1706 133
rect 1760 114 1762 133
rect 1824 114 1826 133
rect 1880 114 1882 133
rect 1944 114 1946 133
rect 2008 114 2010 133
rect 2072 114 2074 133
rect 2144 114 2146 133
rect 2224 114 2226 133
rect 2304 114 2306 133
rect 2392 114 2394 133
rect 2456 114 2458 133
rect 1366 113 1372 114
rect 1326 112 1332 113
rect 1326 108 1327 112
rect 1331 108 1332 112
rect 1366 109 1367 113
rect 1371 109 1372 113
rect 1366 108 1372 109
rect 1422 113 1428 114
rect 1422 109 1423 113
rect 1427 109 1428 113
rect 1422 108 1428 109
rect 1478 113 1484 114
rect 1478 109 1479 113
rect 1483 109 1484 113
rect 1478 108 1484 109
rect 1534 113 1540 114
rect 1534 109 1535 113
rect 1539 109 1540 113
rect 1534 108 1540 109
rect 1590 113 1596 114
rect 1590 109 1591 113
rect 1595 109 1596 113
rect 1590 108 1596 109
rect 1646 113 1652 114
rect 1646 109 1647 113
rect 1651 109 1652 113
rect 1646 108 1652 109
rect 1702 113 1708 114
rect 1702 109 1703 113
rect 1707 109 1708 113
rect 1702 108 1708 109
rect 1758 113 1764 114
rect 1758 109 1759 113
rect 1763 109 1764 113
rect 1758 108 1764 109
rect 1822 113 1828 114
rect 1822 109 1823 113
rect 1827 109 1828 113
rect 1822 108 1828 109
rect 1878 113 1884 114
rect 1878 109 1879 113
rect 1883 109 1884 113
rect 1878 108 1884 109
rect 1942 113 1948 114
rect 1942 109 1943 113
rect 1947 109 1948 113
rect 1942 108 1948 109
rect 2006 113 2012 114
rect 2006 109 2007 113
rect 2011 109 2012 113
rect 2006 108 2012 109
rect 2070 113 2076 114
rect 2070 109 2071 113
rect 2075 109 2076 113
rect 2070 108 2076 109
rect 2142 113 2148 114
rect 2142 109 2143 113
rect 2147 109 2148 113
rect 2142 108 2148 109
rect 2222 113 2228 114
rect 2222 109 2223 113
rect 2227 109 2228 113
rect 2222 108 2228 109
rect 2302 113 2308 114
rect 2302 109 2303 113
rect 2307 109 2308 113
rect 2302 108 2308 109
rect 2390 113 2396 114
rect 2390 109 2391 113
rect 2395 109 2396 113
rect 2390 108 2396 109
rect 2454 113 2460 114
rect 2504 113 2506 133
rect 2454 109 2455 113
rect 2459 109 2460 113
rect 2454 108 2460 109
rect 2502 112 2508 113
rect 2502 108 2503 112
rect 2507 108 2508 112
rect 110 107 116 108
rect 110 103 111 107
rect 115 103 116 107
rect 1286 107 1292 108
rect 1326 107 1332 108
rect 2502 107 2508 108
rect 110 102 116 103
rect 134 104 140 105
rect 112 99 114 102
rect 134 100 135 104
rect 139 100 140 104
rect 134 99 140 100
rect 190 104 196 105
rect 190 100 191 104
rect 195 100 196 104
rect 190 99 196 100
rect 246 104 252 105
rect 246 100 247 104
rect 251 100 252 104
rect 246 99 252 100
rect 302 104 308 105
rect 302 100 303 104
rect 307 100 308 104
rect 302 99 308 100
rect 358 104 364 105
rect 358 100 359 104
rect 363 100 364 104
rect 358 99 364 100
rect 414 104 420 105
rect 414 100 415 104
rect 419 100 420 104
rect 414 99 420 100
rect 470 104 476 105
rect 470 100 471 104
rect 475 100 476 104
rect 470 99 476 100
rect 526 104 532 105
rect 526 100 527 104
rect 531 100 532 104
rect 526 99 532 100
rect 582 104 588 105
rect 582 100 583 104
rect 587 100 588 104
rect 582 99 588 100
rect 638 104 644 105
rect 638 100 639 104
rect 643 100 644 104
rect 638 99 644 100
rect 694 104 700 105
rect 694 100 695 104
rect 699 100 700 104
rect 694 99 700 100
rect 750 104 756 105
rect 750 100 751 104
rect 755 100 756 104
rect 750 99 756 100
rect 814 104 820 105
rect 814 100 815 104
rect 819 100 820 104
rect 814 99 820 100
rect 878 104 884 105
rect 878 100 879 104
rect 883 100 884 104
rect 878 99 884 100
rect 942 104 948 105
rect 942 100 943 104
rect 947 100 948 104
rect 942 99 948 100
rect 1006 104 1012 105
rect 1006 100 1007 104
rect 1011 100 1012 104
rect 1006 99 1012 100
rect 1070 104 1076 105
rect 1070 100 1071 104
rect 1075 100 1076 104
rect 1070 99 1076 100
rect 1134 104 1140 105
rect 1134 100 1135 104
rect 1139 100 1140 104
rect 1286 103 1287 107
rect 1291 103 1292 107
rect 1286 102 1292 103
rect 1134 99 1140 100
rect 1288 99 1290 102
rect 111 98 115 99
rect 111 93 115 94
rect 135 98 139 99
rect 135 93 139 94
rect 191 98 195 99
rect 191 93 195 94
rect 247 98 251 99
rect 247 93 251 94
rect 303 98 307 99
rect 303 93 307 94
rect 359 98 363 99
rect 359 93 363 94
rect 415 98 419 99
rect 415 93 419 94
rect 471 98 475 99
rect 471 93 475 94
rect 527 98 531 99
rect 527 93 531 94
rect 583 98 587 99
rect 583 93 587 94
rect 639 98 643 99
rect 639 93 643 94
rect 695 98 699 99
rect 695 93 699 94
rect 751 98 755 99
rect 751 93 755 94
rect 815 98 819 99
rect 815 93 819 94
rect 879 98 883 99
rect 879 93 883 94
rect 943 98 947 99
rect 943 93 947 94
rect 1007 98 1011 99
rect 1007 93 1011 94
rect 1071 98 1075 99
rect 1071 93 1075 94
rect 1135 98 1139 99
rect 1135 93 1139 94
rect 1287 98 1291 99
rect 1287 93 1291 94
rect 1326 95 1332 96
rect 1326 91 1327 95
rect 1331 91 1332 95
rect 2502 95 2508 96
rect 1326 90 1332 91
rect 1350 92 1356 93
rect 1328 87 1330 90
rect 1350 88 1351 92
rect 1355 88 1356 92
rect 1350 87 1356 88
rect 1406 92 1412 93
rect 1406 88 1407 92
rect 1411 88 1412 92
rect 1406 87 1412 88
rect 1462 92 1468 93
rect 1462 88 1463 92
rect 1467 88 1468 92
rect 1462 87 1468 88
rect 1518 92 1524 93
rect 1518 88 1519 92
rect 1523 88 1524 92
rect 1518 87 1524 88
rect 1574 92 1580 93
rect 1574 88 1575 92
rect 1579 88 1580 92
rect 1574 87 1580 88
rect 1630 92 1636 93
rect 1630 88 1631 92
rect 1635 88 1636 92
rect 1630 87 1636 88
rect 1686 92 1692 93
rect 1686 88 1687 92
rect 1691 88 1692 92
rect 1686 87 1692 88
rect 1742 92 1748 93
rect 1742 88 1743 92
rect 1747 88 1748 92
rect 1742 87 1748 88
rect 1806 92 1812 93
rect 1806 88 1807 92
rect 1811 88 1812 92
rect 1806 87 1812 88
rect 1862 92 1868 93
rect 1862 88 1863 92
rect 1867 88 1868 92
rect 1862 87 1868 88
rect 1926 92 1932 93
rect 1926 88 1927 92
rect 1931 88 1932 92
rect 1926 87 1932 88
rect 1990 92 1996 93
rect 1990 88 1991 92
rect 1995 88 1996 92
rect 1990 87 1996 88
rect 2054 92 2060 93
rect 2054 88 2055 92
rect 2059 88 2060 92
rect 2054 87 2060 88
rect 2126 92 2132 93
rect 2126 88 2127 92
rect 2131 88 2132 92
rect 2126 87 2132 88
rect 2206 92 2212 93
rect 2206 88 2207 92
rect 2211 88 2212 92
rect 2206 87 2212 88
rect 2286 92 2292 93
rect 2286 88 2287 92
rect 2291 88 2292 92
rect 2286 87 2292 88
rect 2374 92 2380 93
rect 2374 88 2375 92
rect 2379 88 2380 92
rect 2374 87 2380 88
rect 2438 92 2444 93
rect 2438 88 2439 92
rect 2443 88 2444 92
rect 2502 91 2503 95
rect 2507 91 2508 95
rect 2502 90 2508 91
rect 2438 87 2444 88
rect 2504 87 2506 90
rect 1327 86 1331 87
rect 1327 81 1331 82
rect 1351 86 1355 87
rect 1351 81 1355 82
rect 1407 86 1411 87
rect 1407 81 1411 82
rect 1463 86 1467 87
rect 1463 81 1467 82
rect 1519 86 1523 87
rect 1519 81 1523 82
rect 1575 86 1579 87
rect 1575 81 1579 82
rect 1631 86 1635 87
rect 1631 81 1635 82
rect 1687 86 1691 87
rect 1687 81 1691 82
rect 1743 86 1747 87
rect 1743 81 1747 82
rect 1807 86 1811 87
rect 1807 81 1811 82
rect 1863 86 1867 87
rect 1863 81 1867 82
rect 1927 86 1931 87
rect 1927 81 1931 82
rect 1991 86 1995 87
rect 1991 81 1995 82
rect 2055 86 2059 87
rect 2055 81 2059 82
rect 2127 86 2131 87
rect 2127 81 2131 82
rect 2207 86 2211 87
rect 2207 81 2211 82
rect 2287 86 2291 87
rect 2287 81 2291 82
rect 2375 86 2379 87
rect 2375 81 2379 82
rect 2439 86 2443 87
rect 2439 81 2443 82
rect 2503 86 2507 87
rect 2503 81 2507 82
<< m4c >>
rect 111 2578 115 2582
rect 135 2578 139 2582
rect 191 2578 195 2582
rect 247 2578 251 2582
rect 303 2578 307 2582
rect 359 2578 363 2582
rect 1287 2578 1291 2582
rect 1327 2558 1331 2562
rect 1495 2558 1499 2562
rect 1551 2558 1555 2562
rect 1607 2558 1611 2562
rect 1663 2558 1667 2562
rect 1719 2558 1723 2562
rect 1775 2558 1779 2562
rect 1831 2558 1835 2562
rect 1887 2558 1891 2562
rect 1943 2558 1947 2562
rect 1999 2558 2003 2562
rect 2055 2558 2059 2562
rect 2111 2558 2115 2562
rect 2167 2558 2171 2562
rect 2503 2558 2507 2562
rect 111 2526 115 2530
rect 151 2526 155 2530
rect 207 2526 211 2530
rect 223 2526 227 2530
rect 263 2526 267 2530
rect 279 2526 283 2530
rect 319 2526 323 2530
rect 343 2526 347 2530
rect 375 2526 379 2530
rect 415 2526 419 2530
rect 487 2526 491 2530
rect 551 2526 555 2530
rect 615 2526 619 2530
rect 679 2526 683 2530
rect 743 2526 747 2530
rect 807 2526 811 2530
rect 871 2526 875 2530
rect 935 2526 939 2530
rect 999 2526 1003 2530
rect 1063 2526 1067 2530
rect 1287 2526 1291 2530
rect 1327 2506 1331 2510
rect 1511 2506 1515 2510
rect 1543 2506 1547 2510
rect 1567 2506 1571 2510
rect 1607 2506 1611 2510
rect 1623 2506 1627 2510
rect 1679 2506 1683 2510
rect 1735 2506 1739 2510
rect 1751 2506 1755 2510
rect 1791 2506 1795 2510
rect 1823 2506 1827 2510
rect 1847 2506 1851 2510
rect 1895 2506 1899 2510
rect 1903 2506 1907 2510
rect 1959 2506 1963 2510
rect 1967 2506 1971 2510
rect 2015 2506 2019 2510
rect 2039 2506 2043 2510
rect 2071 2506 2075 2510
rect 2111 2506 2115 2510
rect 2127 2506 2131 2510
rect 2183 2506 2187 2510
rect 2503 2506 2507 2510
rect 111 2466 115 2470
rect 167 2466 171 2470
rect 207 2466 211 2470
rect 223 2466 227 2470
rect 263 2466 267 2470
rect 279 2466 283 2470
rect 327 2466 331 2470
rect 335 2466 339 2470
rect 391 2466 395 2470
rect 399 2466 403 2470
rect 447 2466 451 2470
rect 471 2466 475 2470
rect 503 2466 507 2470
rect 535 2466 539 2470
rect 559 2466 563 2470
rect 599 2466 603 2470
rect 615 2466 619 2470
rect 663 2466 667 2470
rect 671 2466 675 2470
rect 727 2466 731 2470
rect 783 2466 787 2470
rect 791 2466 795 2470
rect 839 2466 843 2470
rect 855 2466 859 2470
rect 895 2466 899 2470
rect 919 2466 923 2470
rect 951 2466 955 2470
rect 983 2466 987 2470
rect 1007 2466 1011 2470
rect 1047 2466 1051 2470
rect 1063 2466 1067 2470
rect 1287 2466 1291 2470
rect 1327 2450 1331 2454
rect 1527 2450 1531 2454
rect 1543 2450 1547 2454
rect 1591 2450 1595 2454
rect 1607 2450 1611 2454
rect 1663 2450 1667 2454
rect 1671 2450 1675 2454
rect 1735 2450 1739 2454
rect 1743 2450 1747 2454
rect 1807 2450 1811 2454
rect 1815 2450 1819 2454
rect 1879 2450 1883 2454
rect 1951 2450 1955 2454
rect 2023 2450 2027 2454
rect 2095 2450 2099 2454
rect 2167 2450 2171 2454
rect 2503 2450 2507 2454
rect 111 2402 115 2406
rect 183 2402 187 2406
rect 239 2402 243 2406
rect 295 2402 299 2406
rect 351 2402 355 2406
rect 407 2402 411 2406
rect 463 2402 467 2406
rect 519 2402 523 2406
rect 575 2402 579 2406
rect 631 2402 635 2406
rect 687 2402 691 2406
rect 743 2402 747 2406
rect 799 2402 803 2406
rect 855 2402 859 2406
rect 911 2402 915 2406
rect 967 2402 971 2406
rect 1023 2402 1027 2406
rect 1079 2402 1083 2406
rect 1287 2402 1291 2406
rect 1327 2394 1331 2398
rect 1559 2394 1563 2398
rect 1567 2394 1571 2398
rect 1623 2394 1627 2398
rect 1679 2394 1683 2398
rect 1687 2394 1691 2398
rect 1735 2394 1739 2398
rect 1759 2394 1763 2398
rect 1791 2394 1795 2398
rect 1831 2394 1835 2398
rect 1855 2394 1859 2398
rect 1895 2394 1899 2398
rect 1919 2394 1923 2398
rect 1967 2394 1971 2398
rect 1983 2394 1987 2398
rect 2039 2394 2043 2398
rect 2047 2394 2051 2398
rect 2111 2394 2115 2398
rect 2183 2394 2187 2398
rect 2503 2394 2507 2398
rect 111 2342 115 2346
rect 319 2342 323 2346
rect 391 2342 395 2346
rect 463 2342 467 2346
rect 503 2342 507 2346
rect 535 2342 539 2346
rect 559 2342 563 2346
rect 607 2342 611 2346
rect 615 2342 619 2346
rect 671 2342 675 2346
rect 679 2342 683 2346
rect 743 2342 747 2346
rect 807 2342 811 2346
rect 863 2342 867 2346
rect 927 2342 931 2346
rect 991 2342 995 2346
rect 1055 2342 1059 2346
rect 1111 2342 1115 2346
rect 1167 2342 1171 2346
rect 1223 2342 1227 2346
rect 1287 2342 1291 2346
rect 1327 2334 1331 2338
rect 1471 2334 1475 2338
rect 1535 2334 1539 2338
rect 1551 2334 1555 2338
rect 1607 2334 1611 2338
rect 1663 2334 1667 2338
rect 1687 2334 1691 2338
rect 1719 2334 1723 2338
rect 1759 2334 1763 2338
rect 1775 2334 1779 2338
rect 1831 2334 1835 2338
rect 1839 2334 1843 2338
rect 1903 2334 1907 2338
rect 1967 2334 1971 2338
rect 1983 2334 1987 2338
rect 2031 2334 2035 2338
rect 2063 2334 2067 2338
rect 2095 2334 2099 2338
rect 2143 2334 2147 2338
rect 2503 2334 2507 2338
rect 111 2282 115 2286
rect 175 2282 179 2286
rect 271 2282 275 2286
rect 335 2282 339 2286
rect 375 2282 379 2286
rect 407 2282 411 2286
rect 479 2282 483 2286
rect 551 2282 555 2286
rect 591 2282 595 2286
rect 623 2282 627 2286
rect 695 2282 699 2286
rect 703 2282 707 2286
rect 759 2282 763 2286
rect 807 2282 811 2286
rect 823 2282 827 2286
rect 879 2282 883 2286
rect 911 2282 915 2286
rect 943 2282 947 2286
rect 1007 2282 1011 2286
rect 1015 2282 1019 2286
rect 1071 2282 1075 2286
rect 1127 2282 1131 2286
rect 1183 2282 1187 2286
rect 1239 2282 1243 2286
rect 1287 2282 1291 2286
rect 1327 2282 1331 2286
rect 1383 2282 1387 2286
rect 1479 2282 1483 2286
rect 1487 2282 1491 2286
rect 1551 2282 1555 2286
rect 1583 2282 1587 2286
rect 1623 2282 1627 2286
rect 1687 2282 1691 2286
rect 1703 2282 1707 2286
rect 1775 2282 1779 2286
rect 1791 2282 1795 2286
rect 1847 2282 1851 2286
rect 1903 2282 1907 2286
rect 1919 2282 1923 2286
rect 1999 2282 2003 2286
rect 2015 2282 2019 2286
rect 2079 2282 2083 2286
rect 2127 2282 2131 2286
rect 2159 2282 2163 2286
rect 2239 2282 2243 2286
rect 2503 2282 2507 2286
rect 111 2230 115 2234
rect 143 2230 147 2234
rect 159 2230 163 2234
rect 231 2230 235 2234
rect 255 2230 259 2234
rect 319 2230 323 2234
rect 359 2230 363 2234
rect 415 2230 419 2234
rect 463 2230 467 2234
rect 519 2230 523 2234
rect 575 2230 579 2234
rect 623 2230 627 2234
rect 687 2230 691 2234
rect 727 2230 731 2234
rect 791 2230 795 2234
rect 831 2230 835 2234
rect 895 2230 899 2234
rect 935 2230 939 2234
rect 999 2230 1003 2234
rect 1039 2230 1043 2234
rect 1111 2230 1115 2234
rect 1143 2230 1147 2234
rect 1223 2230 1227 2234
rect 1287 2230 1291 2234
rect 1327 2230 1331 2234
rect 1367 2230 1371 2234
rect 1463 2230 1467 2234
rect 1487 2230 1491 2234
rect 1567 2230 1571 2234
rect 1607 2230 1611 2234
rect 1671 2230 1675 2234
rect 1719 2230 1723 2234
rect 1775 2230 1779 2234
rect 1815 2230 1819 2234
rect 1887 2230 1891 2234
rect 1903 2230 1907 2234
rect 1983 2230 1987 2234
rect 1999 2230 2003 2234
rect 2055 2230 2059 2234
rect 2111 2230 2115 2234
rect 2127 2230 2131 2234
rect 2191 2230 2195 2234
rect 2223 2230 2227 2234
rect 2255 2230 2259 2234
rect 2319 2230 2323 2234
rect 2383 2230 2387 2234
rect 2439 2230 2443 2234
rect 2503 2230 2507 2234
rect 111 2178 115 2182
rect 159 2178 163 2182
rect 247 2178 251 2182
rect 255 2178 259 2182
rect 335 2178 339 2182
rect 351 2178 355 2182
rect 431 2178 435 2182
rect 455 2178 459 2182
rect 535 2178 539 2182
rect 559 2178 563 2182
rect 639 2178 643 2182
rect 663 2178 667 2182
rect 743 2178 747 2182
rect 767 2178 771 2182
rect 847 2178 851 2182
rect 863 2178 867 2182
rect 951 2178 955 2182
rect 959 2178 963 2182
rect 1055 2178 1059 2182
rect 1159 2178 1163 2182
rect 1239 2178 1243 2182
rect 1287 2178 1291 2182
rect 1327 2158 1331 2162
rect 1383 2158 1387 2162
rect 1407 2158 1411 2162
rect 1503 2158 1507 2162
rect 1623 2158 1627 2162
rect 1735 2158 1739 2162
rect 1815 2158 1819 2162
rect 1831 2158 1835 2162
rect 1919 2158 1923 2162
rect 1991 2158 1995 2162
rect 1999 2158 2003 2162
rect 2071 2158 2075 2162
rect 2143 2158 2147 2162
rect 2159 2158 2163 2162
rect 2207 2158 2211 2162
rect 2271 2158 2275 2162
rect 2319 2158 2323 2162
rect 2335 2158 2339 2162
rect 2399 2158 2403 2162
rect 2455 2158 2459 2162
rect 2503 2158 2507 2162
rect 111 2126 115 2130
rect 239 2126 243 2130
rect 303 2126 307 2130
rect 335 2126 339 2130
rect 359 2126 363 2130
rect 423 2126 427 2130
rect 439 2126 443 2130
rect 487 2126 491 2130
rect 543 2126 547 2130
rect 559 2126 563 2130
rect 631 2126 635 2130
rect 647 2126 651 2130
rect 711 2126 715 2130
rect 751 2126 755 2130
rect 799 2126 803 2130
rect 847 2126 851 2130
rect 887 2126 891 2130
rect 943 2126 947 2130
rect 975 2126 979 2130
rect 1039 2126 1043 2130
rect 1063 2126 1067 2130
rect 1143 2126 1147 2130
rect 1151 2126 1155 2130
rect 1223 2126 1227 2130
rect 1287 2126 1291 2130
rect 1327 2106 1331 2110
rect 1383 2106 1387 2110
rect 1391 2106 1395 2110
rect 1551 2106 1555 2110
rect 1607 2106 1611 2110
rect 1711 2106 1715 2110
rect 1799 2106 1803 2110
rect 1855 2106 1859 2110
rect 1975 2106 1979 2110
rect 1991 2106 1995 2110
rect 2119 2106 2123 2110
rect 2143 2106 2147 2110
rect 2239 2106 2243 2110
rect 2303 2106 2307 2110
rect 2367 2106 2371 2110
rect 2439 2106 2443 2110
rect 2503 2106 2507 2110
rect 111 2070 115 2074
rect 319 2070 323 2074
rect 375 2070 379 2074
rect 399 2070 403 2074
rect 439 2070 443 2074
rect 455 2070 459 2074
rect 503 2070 507 2074
rect 511 2070 515 2074
rect 575 2070 579 2074
rect 639 2070 643 2074
rect 647 2070 651 2074
rect 711 2070 715 2074
rect 727 2070 731 2074
rect 791 2070 795 2074
rect 815 2070 819 2074
rect 863 2070 867 2074
rect 903 2070 907 2074
rect 943 2070 947 2074
rect 991 2070 995 2074
rect 1023 2070 1027 2074
rect 1079 2070 1083 2074
rect 1103 2070 1107 2074
rect 1167 2070 1171 2074
rect 1183 2070 1187 2074
rect 1239 2070 1243 2074
rect 1287 2070 1291 2074
rect 1327 2050 1331 2054
rect 1399 2050 1403 2054
rect 1447 2050 1451 2054
rect 1551 2050 1555 2054
rect 1567 2050 1571 2054
rect 1655 2050 1659 2054
rect 1727 2050 1731 2054
rect 1751 2050 1755 2054
rect 1839 2050 1843 2054
rect 1871 2050 1875 2054
rect 1927 2050 1931 2054
rect 2007 2050 2011 2054
rect 2023 2050 2027 2054
rect 2119 2050 2123 2054
rect 2135 2050 2139 2054
rect 2255 2050 2259 2054
rect 2383 2050 2387 2054
rect 2503 2050 2507 2054
rect 111 2014 115 2018
rect 231 2014 235 2018
rect 287 2014 291 2018
rect 359 2014 363 2018
rect 383 2014 387 2018
rect 439 2014 443 2018
rect 495 2014 499 2018
rect 535 2014 539 2018
rect 559 2014 563 2018
rect 623 2014 627 2018
rect 631 2014 635 2018
rect 695 2014 699 2018
rect 735 2014 739 2018
rect 775 2014 779 2018
rect 847 2014 851 2018
rect 927 2014 931 2018
rect 959 2014 963 2018
rect 1007 2014 1011 2018
rect 1079 2014 1083 2018
rect 1087 2014 1091 2018
rect 1167 2014 1171 2018
rect 1199 2014 1203 2018
rect 1223 2014 1227 2018
rect 1287 2014 1291 2018
rect 1327 1994 1331 1998
rect 1431 1994 1435 1998
rect 1455 1994 1459 1998
rect 1511 1994 1515 1998
rect 1535 1994 1539 1998
rect 1575 1994 1579 1998
rect 1639 1994 1643 1998
rect 1703 1994 1707 1998
rect 1735 1994 1739 1998
rect 1767 1994 1771 1998
rect 1823 1994 1827 1998
rect 1831 1994 1835 1998
rect 1895 1994 1899 1998
rect 1911 1994 1915 1998
rect 1959 1994 1963 1998
rect 2007 1994 2011 1998
rect 2031 1994 2035 1998
rect 2103 1994 2107 1998
rect 2503 1994 2507 1998
rect 111 1958 115 1962
rect 151 1958 155 1962
rect 215 1958 219 1962
rect 247 1958 251 1962
rect 303 1958 307 1962
rect 319 1958 323 1962
rect 375 1958 379 1962
rect 439 1958 443 1962
rect 455 1958 459 1962
rect 551 1958 555 1962
rect 583 1958 587 1962
rect 647 1958 651 1962
rect 743 1958 747 1962
rect 751 1958 755 1962
rect 863 1958 867 1962
rect 919 1958 923 1962
rect 975 1958 979 1962
rect 1095 1958 1099 1962
rect 1215 1958 1219 1962
rect 1287 1958 1291 1962
rect 1327 1938 1331 1942
rect 1471 1938 1475 1942
rect 1527 1938 1531 1942
rect 1567 1938 1571 1942
rect 1591 1938 1595 1942
rect 1631 1938 1635 1942
rect 1655 1938 1659 1942
rect 1703 1938 1707 1942
rect 1719 1938 1723 1942
rect 1775 1938 1779 1942
rect 1783 1938 1787 1942
rect 1847 1938 1851 1942
rect 1911 1938 1915 1942
rect 1919 1938 1923 1942
rect 1975 1938 1979 1942
rect 1999 1938 2003 1942
rect 2047 1938 2051 1942
rect 2087 1938 2091 1942
rect 2183 1938 2187 1942
rect 2279 1938 2283 1942
rect 2375 1938 2379 1942
rect 2455 1938 2459 1942
rect 2503 1938 2507 1942
rect 111 1898 115 1902
rect 135 1898 139 1902
rect 191 1898 195 1902
rect 199 1898 203 1902
rect 271 1898 275 1902
rect 303 1898 307 1902
rect 359 1898 363 1902
rect 423 1898 427 1902
rect 455 1898 459 1902
rect 543 1898 547 1902
rect 567 1898 571 1902
rect 631 1898 635 1902
rect 719 1898 723 1902
rect 727 1898 731 1902
rect 799 1898 803 1902
rect 871 1898 875 1902
rect 903 1898 907 1902
rect 943 1898 947 1902
rect 1015 1898 1019 1902
rect 1079 1898 1083 1902
rect 1087 1898 1091 1902
rect 1159 1898 1163 1902
rect 1287 1898 1291 1902
rect 1327 1882 1331 1886
rect 1551 1882 1555 1886
rect 1607 1882 1611 1886
rect 1615 1882 1619 1886
rect 1663 1882 1667 1886
rect 1687 1882 1691 1886
rect 1727 1882 1731 1886
rect 1759 1882 1763 1886
rect 1799 1882 1803 1886
rect 1831 1882 1835 1886
rect 1871 1882 1875 1886
rect 1903 1882 1907 1886
rect 1943 1882 1947 1886
rect 1983 1882 1987 1886
rect 2007 1882 2011 1886
rect 2071 1882 2075 1886
rect 2135 1882 2139 1886
rect 2167 1882 2171 1886
rect 2199 1882 2203 1886
rect 2263 1882 2267 1886
rect 2327 1882 2331 1886
rect 2359 1882 2363 1886
rect 2383 1882 2387 1886
rect 2439 1882 2443 1886
rect 2503 1882 2507 1886
rect 111 1846 115 1850
rect 151 1846 155 1850
rect 207 1846 211 1850
rect 287 1846 291 1850
rect 295 1846 299 1850
rect 375 1846 379 1850
rect 391 1846 395 1850
rect 471 1846 475 1850
rect 495 1846 499 1850
rect 559 1846 563 1850
rect 591 1846 595 1850
rect 647 1846 651 1850
rect 687 1846 691 1850
rect 735 1846 739 1850
rect 775 1846 779 1850
rect 815 1846 819 1850
rect 855 1846 859 1850
rect 887 1846 891 1850
rect 927 1846 931 1850
rect 959 1846 963 1850
rect 999 1846 1003 1850
rect 1031 1846 1035 1850
rect 1079 1846 1083 1850
rect 1103 1846 1107 1850
rect 1159 1846 1163 1850
rect 1175 1846 1179 1850
rect 1287 1846 1291 1850
rect 1327 1826 1331 1830
rect 1623 1826 1627 1830
rect 1631 1826 1635 1830
rect 1679 1826 1683 1830
rect 1719 1826 1723 1830
rect 1743 1826 1747 1830
rect 1815 1826 1819 1830
rect 1887 1826 1891 1830
rect 1927 1826 1931 1830
rect 1959 1826 1963 1830
rect 2023 1826 2027 1830
rect 2055 1826 2059 1830
rect 2087 1826 2091 1830
rect 2151 1826 2155 1830
rect 2191 1826 2195 1830
rect 2215 1826 2219 1830
rect 2279 1826 2283 1830
rect 2335 1826 2339 1830
rect 2343 1826 2347 1830
rect 2399 1826 2403 1830
rect 2455 1826 2459 1830
rect 2503 1826 2507 1830
rect 111 1782 115 1786
rect 135 1782 139 1786
rect 191 1782 195 1786
rect 199 1782 203 1786
rect 279 1782 283 1786
rect 295 1782 299 1786
rect 375 1782 379 1786
rect 399 1782 403 1786
rect 479 1782 483 1786
rect 503 1782 507 1786
rect 575 1782 579 1786
rect 607 1782 611 1786
rect 671 1782 675 1786
rect 703 1782 707 1786
rect 759 1782 763 1786
rect 799 1782 803 1786
rect 839 1782 843 1786
rect 887 1782 891 1786
rect 911 1782 915 1786
rect 975 1782 979 1786
rect 983 1782 987 1786
rect 1063 1782 1067 1786
rect 1143 1782 1147 1786
rect 1151 1782 1155 1786
rect 1287 1782 1291 1786
rect 1327 1774 1331 1778
rect 1527 1774 1531 1778
rect 1607 1774 1611 1778
rect 1615 1774 1619 1778
rect 1695 1774 1699 1778
rect 1703 1774 1707 1778
rect 1791 1774 1795 1778
rect 1799 1774 1803 1778
rect 1879 1774 1883 1778
rect 1911 1774 1915 1778
rect 1967 1774 1971 1778
rect 2039 1774 2043 1778
rect 2055 1774 2059 1778
rect 2135 1774 2139 1778
rect 2175 1774 2179 1778
rect 2215 1774 2219 1778
rect 2295 1774 2299 1778
rect 2319 1774 2323 1778
rect 2375 1774 2379 1778
rect 2439 1774 2443 1778
rect 2503 1774 2507 1778
rect 111 1726 115 1730
rect 151 1726 155 1730
rect 167 1726 171 1730
rect 215 1726 219 1730
rect 239 1726 243 1730
rect 311 1726 315 1730
rect 319 1726 323 1730
rect 407 1726 411 1730
rect 415 1726 419 1730
rect 503 1726 507 1730
rect 519 1726 523 1730
rect 607 1726 611 1730
rect 623 1726 627 1730
rect 711 1726 715 1730
rect 719 1726 723 1730
rect 815 1726 819 1730
rect 823 1726 827 1730
rect 903 1726 907 1730
rect 935 1726 939 1730
rect 991 1726 995 1730
rect 1047 1726 1051 1730
rect 1079 1726 1083 1730
rect 1159 1726 1163 1730
rect 1167 1726 1171 1730
rect 1287 1726 1291 1730
rect 1327 1718 1331 1722
rect 1399 1718 1403 1722
rect 1463 1718 1467 1722
rect 1543 1718 1547 1722
rect 1623 1718 1627 1722
rect 1631 1718 1635 1722
rect 1711 1718 1715 1722
rect 1727 1718 1731 1722
rect 1807 1718 1811 1722
rect 1823 1718 1827 1722
rect 1895 1718 1899 1722
rect 1919 1718 1923 1722
rect 1983 1718 1987 1722
rect 2015 1718 2019 1722
rect 2071 1718 2075 1722
rect 2111 1718 2115 1722
rect 2151 1718 2155 1722
rect 2199 1718 2203 1722
rect 2231 1718 2235 1722
rect 2287 1718 2291 1722
rect 2311 1718 2315 1722
rect 2383 1718 2387 1722
rect 2391 1718 2395 1722
rect 2455 1718 2459 1722
rect 2503 1718 2507 1722
rect 111 1670 115 1674
rect 151 1670 155 1674
rect 223 1670 227 1674
rect 255 1670 259 1674
rect 303 1670 307 1674
rect 319 1670 323 1674
rect 391 1670 395 1674
rect 399 1670 403 1674
rect 487 1670 491 1674
rect 575 1670 579 1674
rect 591 1670 595 1674
rect 671 1670 675 1674
rect 695 1670 699 1674
rect 767 1670 771 1674
rect 807 1670 811 1674
rect 863 1670 867 1674
rect 919 1670 923 1674
rect 959 1670 963 1674
rect 1031 1670 1035 1674
rect 1063 1670 1067 1674
rect 1143 1670 1147 1674
rect 1167 1670 1171 1674
rect 1287 1670 1291 1674
rect 1327 1662 1331 1666
rect 1351 1662 1355 1666
rect 1383 1662 1387 1666
rect 1407 1662 1411 1666
rect 1447 1662 1451 1666
rect 1495 1662 1499 1666
rect 1527 1662 1531 1666
rect 1583 1662 1587 1666
rect 1615 1662 1619 1666
rect 1679 1662 1683 1666
rect 1711 1662 1715 1666
rect 1783 1662 1787 1666
rect 1807 1662 1811 1666
rect 1895 1662 1899 1666
rect 1903 1662 1907 1666
rect 1999 1662 2003 1666
rect 2023 1662 2027 1666
rect 2095 1662 2099 1666
rect 2159 1662 2163 1666
rect 2183 1662 2187 1666
rect 2271 1662 2275 1666
rect 2303 1662 2307 1666
rect 2367 1662 2371 1666
rect 2439 1662 2443 1666
rect 2503 1662 2507 1666
rect 111 1614 115 1618
rect 271 1614 275 1618
rect 303 1614 307 1618
rect 335 1614 339 1618
rect 359 1614 363 1618
rect 415 1614 419 1618
rect 431 1614 435 1618
rect 503 1614 507 1618
rect 511 1614 515 1618
rect 591 1614 595 1618
rect 599 1614 603 1618
rect 687 1614 691 1618
rect 695 1614 699 1618
rect 783 1614 787 1618
rect 791 1614 795 1618
rect 879 1614 883 1618
rect 895 1614 899 1618
rect 975 1614 979 1618
rect 1007 1614 1011 1618
rect 1079 1614 1083 1618
rect 1119 1614 1123 1618
rect 1183 1614 1187 1618
rect 1287 1614 1291 1618
rect 1327 1610 1331 1614
rect 1367 1610 1371 1614
rect 1423 1610 1427 1614
rect 1479 1610 1483 1614
rect 1511 1610 1515 1614
rect 1559 1610 1563 1614
rect 1599 1610 1603 1614
rect 1639 1610 1643 1614
rect 1695 1610 1699 1614
rect 1719 1610 1723 1614
rect 1791 1610 1795 1614
rect 1799 1610 1803 1614
rect 1871 1610 1875 1614
rect 1911 1610 1915 1614
rect 1951 1610 1955 1614
rect 2031 1610 2035 1614
rect 2039 1610 2043 1614
rect 2175 1610 2179 1614
rect 2319 1610 2323 1614
rect 2455 1610 2459 1614
rect 2503 1610 2507 1614
rect 111 1562 115 1566
rect 247 1562 251 1566
rect 287 1562 291 1566
rect 319 1562 323 1566
rect 343 1562 347 1566
rect 399 1562 403 1566
rect 415 1562 419 1566
rect 487 1562 491 1566
rect 495 1562 499 1566
rect 583 1562 587 1566
rect 671 1562 675 1566
rect 679 1562 683 1566
rect 759 1562 763 1566
rect 775 1562 779 1566
rect 847 1562 851 1566
rect 879 1562 883 1566
rect 927 1562 931 1566
rect 991 1562 995 1566
rect 1007 1562 1011 1566
rect 1087 1562 1091 1566
rect 1103 1562 1107 1566
rect 1167 1562 1171 1566
rect 1223 1562 1227 1566
rect 1287 1562 1291 1566
rect 1327 1558 1331 1562
rect 1351 1558 1355 1562
rect 1407 1558 1411 1562
rect 1463 1558 1467 1562
rect 1471 1558 1475 1562
rect 1543 1558 1547 1562
rect 1607 1558 1611 1562
rect 1623 1558 1627 1562
rect 1703 1558 1707 1562
rect 1735 1558 1739 1562
rect 1775 1558 1779 1562
rect 1855 1558 1859 1562
rect 1871 1558 1875 1562
rect 1935 1558 1939 1562
rect 2007 1558 2011 1562
rect 2015 1558 2019 1562
rect 2503 1558 2507 1562
rect 111 1502 115 1506
rect 263 1502 267 1506
rect 279 1502 283 1506
rect 335 1502 339 1506
rect 343 1502 347 1506
rect 415 1502 419 1506
rect 495 1502 499 1506
rect 503 1502 507 1506
rect 575 1502 579 1506
rect 599 1502 603 1506
rect 655 1502 659 1506
rect 687 1502 691 1506
rect 735 1502 739 1506
rect 775 1502 779 1506
rect 815 1502 819 1506
rect 863 1502 867 1506
rect 895 1502 899 1506
rect 943 1502 947 1506
rect 975 1502 979 1506
rect 1023 1502 1027 1506
rect 1055 1502 1059 1506
rect 1103 1502 1107 1506
rect 1143 1502 1147 1506
rect 1183 1502 1187 1506
rect 1239 1502 1243 1506
rect 1287 1502 1291 1506
rect 1327 1506 1331 1510
rect 1367 1506 1371 1510
rect 1423 1506 1427 1510
rect 1479 1506 1483 1510
rect 1487 1506 1491 1510
rect 1551 1506 1555 1510
rect 1623 1506 1627 1510
rect 1631 1506 1635 1510
rect 1711 1506 1715 1510
rect 1751 1506 1755 1510
rect 1791 1506 1795 1510
rect 1871 1506 1875 1510
rect 1887 1506 1891 1510
rect 1951 1506 1955 1510
rect 2023 1506 2027 1510
rect 2031 1506 2035 1510
rect 2119 1506 2123 1510
rect 2503 1506 2507 1510
rect 111 1446 115 1450
rect 191 1446 195 1450
rect 255 1446 259 1450
rect 263 1446 267 1450
rect 327 1446 331 1450
rect 399 1446 403 1450
rect 407 1446 411 1450
rect 479 1446 483 1450
rect 503 1446 507 1450
rect 559 1446 563 1450
rect 607 1446 611 1450
rect 639 1446 643 1450
rect 711 1446 715 1450
rect 719 1446 723 1450
rect 799 1446 803 1450
rect 815 1446 819 1450
rect 879 1446 883 1450
rect 919 1446 923 1450
rect 959 1446 963 1450
rect 1023 1446 1027 1450
rect 1039 1446 1043 1450
rect 1127 1446 1131 1450
rect 1223 1446 1227 1450
rect 1287 1446 1291 1450
rect 1327 1446 1331 1450
rect 1351 1446 1355 1450
rect 1359 1446 1363 1450
rect 1407 1446 1411 1450
rect 1447 1446 1451 1450
rect 1463 1446 1467 1450
rect 1535 1446 1539 1450
rect 1615 1446 1619 1450
rect 1631 1446 1635 1450
rect 1695 1446 1699 1450
rect 1727 1446 1731 1450
rect 1775 1446 1779 1450
rect 1815 1446 1819 1450
rect 1855 1446 1859 1450
rect 1903 1446 1907 1450
rect 1935 1446 1939 1450
rect 1991 1446 1995 1450
rect 2015 1446 2019 1450
rect 2071 1446 2075 1450
rect 2103 1446 2107 1450
rect 2159 1446 2163 1450
rect 2247 1446 2251 1450
rect 2503 1446 2507 1450
rect 111 1390 115 1394
rect 151 1390 155 1394
rect 207 1390 211 1394
rect 223 1390 227 1394
rect 271 1390 275 1394
rect 295 1390 299 1394
rect 343 1390 347 1394
rect 359 1390 363 1394
rect 423 1390 427 1394
rect 431 1390 435 1394
rect 503 1390 507 1394
rect 519 1390 523 1394
rect 583 1390 587 1394
rect 623 1390 627 1394
rect 663 1390 667 1394
rect 727 1390 731 1394
rect 751 1390 755 1394
rect 831 1390 835 1394
rect 839 1390 843 1394
rect 927 1390 931 1394
rect 935 1390 939 1394
rect 1015 1390 1019 1394
rect 1039 1390 1043 1394
rect 1103 1390 1107 1394
rect 1143 1390 1147 1394
rect 1199 1390 1203 1394
rect 1239 1390 1243 1394
rect 1287 1390 1291 1394
rect 1327 1394 1331 1398
rect 1375 1394 1379 1398
rect 1463 1394 1467 1398
rect 1551 1394 1555 1398
rect 1567 1394 1571 1398
rect 1647 1394 1651 1398
rect 1735 1394 1739 1398
rect 1743 1394 1747 1398
rect 1831 1394 1835 1398
rect 1919 1394 1923 1398
rect 2007 1394 2011 1398
rect 2087 1394 2091 1398
rect 2095 1394 2099 1398
rect 2175 1394 2179 1398
rect 2247 1394 2251 1398
rect 2263 1394 2267 1398
rect 2319 1394 2323 1398
rect 2399 1394 2403 1398
rect 2455 1394 2459 1398
rect 2503 1394 2507 1398
rect 1327 1342 1331 1346
rect 1551 1342 1555 1346
rect 1583 1342 1587 1346
rect 1631 1342 1635 1346
rect 1647 1342 1651 1346
rect 1719 1342 1723 1346
rect 1727 1342 1731 1346
rect 1807 1342 1811 1346
rect 1815 1342 1819 1346
rect 1895 1342 1899 1346
rect 1903 1342 1907 1346
rect 1983 1342 1987 1346
rect 1991 1342 1995 1346
rect 2063 1342 2067 1346
rect 2079 1342 2083 1346
rect 2143 1342 2147 1346
rect 2159 1342 2163 1346
rect 2223 1342 2227 1346
rect 2231 1342 2235 1346
rect 2303 1342 2307 1346
rect 2383 1342 2387 1346
rect 2439 1342 2443 1346
rect 2503 1342 2507 1346
rect 111 1322 115 1326
rect 135 1322 139 1326
rect 207 1322 211 1326
rect 239 1322 243 1326
rect 279 1322 283 1326
rect 343 1322 347 1326
rect 367 1322 371 1326
rect 415 1322 419 1326
rect 479 1322 483 1326
rect 487 1322 491 1326
rect 567 1322 571 1326
rect 583 1322 587 1326
rect 647 1322 651 1326
rect 687 1322 691 1326
rect 735 1322 739 1326
rect 783 1322 787 1326
rect 823 1322 827 1326
rect 879 1322 883 1326
rect 911 1322 915 1326
rect 975 1322 979 1326
rect 999 1322 1003 1326
rect 1087 1322 1091 1326
rect 1183 1322 1187 1326
rect 1287 1322 1291 1326
rect 1327 1290 1331 1294
rect 1567 1290 1571 1294
rect 1599 1290 1603 1294
rect 1631 1290 1635 1294
rect 1663 1290 1667 1294
rect 1711 1290 1715 1294
rect 1743 1290 1747 1294
rect 1799 1290 1803 1294
rect 1823 1290 1827 1294
rect 1895 1290 1899 1294
rect 1911 1290 1915 1294
rect 1991 1290 1995 1294
rect 1999 1290 2003 1294
rect 2079 1290 2083 1294
rect 2095 1290 2099 1294
rect 2159 1290 2163 1294
rect 2207 1290 2211 1294
rect 2239 1290 2243 1294
rect 2319 1290 2323 1294
rect 2399 1290 2403 1294
rect 2455 1290 2459 1294
rect 2503 1290 2507 1294
rect 111 1262 115 1266
rect 151 1262 155 1266
rect 215 1262 219 1266
rect 255 1262 259 1266
rect 303 1262 307 1266
rect 383 1262 387 1266
rect 391 1262 395 1266
rect 471 1262 475 1266
rect 495 1262 499 1266
rect 551 1262 555 1266
rect 599 1262 603 1266
rect 623 1262 627 1266
rect 695 1262 699 1266
rect 703 1262 707 1266
rect 767 1262 771 1266
rect 799 1262 803 1266
rect 839 1262 843 1266
rect 895 1262 899 1266
rect 919 1262 923 1266
rect 991 1262 995 1266
rect 1287 1262 1291 1266
rect 1327 1234 1331 1238
rect 1519 1234 1523 1238
rect 1551 1234 1555 1238
rect 1575 1234 1579 1238
rect 1615 1234 1619 1238
rect 1631 1234 1635 1238
rect 1687 1234 1691 1238
rect 1695 1234 1699 1238
rect 1743 1234 1747 1238
rect 1783 1234 1787 1238
rect 1799 1234 1803 1238
rect 1855 1234 1859 1238
rect 1879 1234 1883 1238
rect 1911 1234 1915 1238
rect 1967 1234 1971 1238
rect 1975 1234 1979 1238
rect 2031 1234 2035 1238
rect 2079 1234 2083 1238
rect 2103 1234 2107 1238
rect 2183 1234 2187 1238
rect 2191 1234 2195 1238
rect 2271 1234 2275 1238
rect 2303 1234 2307 1238
rect 2367 1234 2371 1238
rect 2439 1234 2443 1238
rect 2503 1234 2507 1238
rect 111 1206 115 1210
rect 135 1206 139 1210
rect 191 1206 195 1210
rect 199 1206 203 1210
rect 271 1206 275 1210
rect 287 1206 291 1210
rect 351 1206 355 1210
rect 375 1206 379 1210
rect 431 1206 435 1210
rect 455 1206 459 1210
rect 511 1206 515 1210
rect 535 1206 539 1210
rect 583 1206 587 1210
rect 607 1206 611 1210
rect 647 1206 651 1210
rect 679 1206 683 1210
rect 719 1206 723 1210
rect 751 1206 755 1210
rect 791 1206 795 1210
rect 823 1206 827 1210
rect 863 1206 867 1210
rect 903 1206 907 1210
rect 1287 1206 1291 1210
rect 1327 1178 1331 1182
rect 1535 1178 1539 1182
rect 1567 1178 1571 1182
rect 1591 1178 1595 1182
rect 1631 1178 1635 1182
rect 1647 1178 1651 1182
rect 1703 1178 1707 1182
rect 1759 1178 1763 1182
rect 1791 1178 1795 1182
rect 1815 1178 1819 1182
rect 1871 1178 1875 1182
rect 1903 1178 1907 1182
rect 1927 1178 1931 1182
rect 1983 1178 1987 1182
rect 2031 1178 2035 1182
rect 2047 1178 2051 1182
rect 2119 1178 2123 1182
rect 2175 1178 2179 1182
rect 2199 1178 2203 1182
rect 2287 1178 2291 1182
rect 2327 1178 2331 1182
rect 2383 1178 2387 1182
rect 2455 1178 2459 1182
rect 2503 1178 2507 1182
rect 111 1150 115 1154
rect 151 1150 155 1154
rect 183 1150 187 1154
rect 207 1150 211 1154
rect 279 1150 283 1154
rect 287 1150 291 1154
rect 367 1150 371 1154
rect 375 1150 379 1154
rect 447 1150 451 1154
rect 471 1150 475 1154
rect 527 1150 531 1154
rect 567 1150 571 1154
rect 599 1150 603 1154
rect 655 1150 659 1154
rect 663 1150 667 1154
rect 735 1150 739 1154
rect 807 1150 811 1154
rect 879 1150 883 1154
rect 959 1150 963 1154
rect 1039 1150 1043 1154
rect 1287 1150 1291 1154
rect 1327 1126 1331 1130
rect 1383 1126 1387 1130
rect 1447 1126 1451 1130
rect 1519 1126 1523 1130
rect 1551 1126 1555 1130
rect 1591 1126 1595 1130
rect 1615 1126 1619 1130
rect 1671 1126 1675 1130
rect 1687 1126 1691 1130
rect 1751 1126 1755 1130
rect 1775 1126 1779 1130
rect 1831 1126 1835 1130
rect 1887 1126 1891 1130
rect 1911 1126 1915 1130
rect 1983 1126 1987 1130
rect 2015 1126 2019 1130
rect 2055 1126 2059 1130
rect 2135 1126 2139 1130
rect 2159 1126 2163 1130
rect 2215 1126 2219 1130
rect 2311 1126 2315 1130
rect 2439 1126 2443 1130
rect 2503 1126 2507 1130
rect 111 1090 115 1094
rect 167 1090 171 1094
rect 207 1090 211 1094
rect 263 1090 267 1094
rect 279 1090 283 1094
rect 359 1090 363 1094
rect 447 1090 451 1094
rect 455 1090 459 1094
rect 543 1090 547 1094
rect 551 1090 555 1094
rect 639 1090 643 1094
rect 719 1090 723 1094
rect 727 1090 731 1094
rect 791 1090 795 1094
rect 815 1090 819 1094
rect 863 1090 867 1094
rect 895 1090 899 1094
rect 943 1090 947 1094
rect 975 1090 979 1094
rect 1023 1090 1027 1094
rect 1055 1090 1059 1094
rect 1143 1090 1147 1094
rect 1287 1090 1291 1094
rect 1327 1066 1331 1070
rect 1367 1066 1371 1070
rect 1399 1066 1403 1070
rect 1455 1066 1459 1070
rect 1463 1066 1467 1070
rect 1535 1066 1539 1070
rect 1575 1066 1579 1070
rect 1607 1066 1611 1070
rect 1687 1066 1691 1070
rect 1695 1066 1699 1070
rect 1767 1066 1771 1070
rect 1815 1066 1819 1070
rect 1847 1066 1851 1070
rect 1927 1066 1931 1070
rect 1999 1066 2003 1070
rect 2039 1066 2043 1070
rect 2071 1066 2075 1070
rect 2151 1066 2155 1070
rect 2231 1066 2235 1070
rect 2255 1066 2259 1070
rect 2367 1066 2371 1070
rect 2455 1066 2459 1070
rect 2503 1066 2507 1070
rect 111 1030 115 1034
rect 223 1030 227 1034
rect 295 1030 299 1034
rect 375 1030 379 1034
rect 383 1030 387 1034
rect 463 1030 467 1034
rect 479 1030 483 1034
rect 559 1030 563 1034
rect 575 1030 579 1034
rect 655 1030 659 1034
rect 671 1030 675 1034
rect 743 1030 747 1034
rect 767 1030 771 1034
rect 831 1030 835 1034
rect 855 1030 859 1034
rect 911 1030 915 1034
rect 943 1030 947 1034
rect 991 1030 995 1034
rect 1023 1030 1027 1034
rect 1071 1030 1075 1034
rect 1103 1030 1107 1034
rect 1159 1030 1163 1034
rect 1183 1030 1187 1034
rect 1239 1030 1243 1034
rect 1287 1030 1291 1034
rect 1327 1010 1331 1014
rect 1351 1010 1355 1014
rect 1439 1010 1443 1014
rect 1511 1010 1515 1014
rect 1559 1010 1563 1014
rect 1679 1010 1683 1014
rect 1799 1010 1803 1014
rect 1823 1010 1827 1014
rect 1911 1010 1915 1014
rect 1951 1010 1955 1014
rect 2023 1010 2027 1014
rect 2071 1010 2075 1014
rect 2135 1010 2139 1014
rect 2175 1010 2179 1014
rect 2239 1010 2243 1014
rect 2271 1010 2275 1014
rect 2351 1010 2355 1014
rect 2367 1010 2371 1014
rect 2439 1010 2443 1014
rect 2503 1010 2507 1014
rect 111 978 115 982
rect 271 978 275 982
rect 279 978 283 982
rect 359 978 363 982
rect 367 978 371 982
rect 455 978 459 982
rect 463 978 467 982
rect 551 978 555 982
rect 559 978 563 982
rect 655 978 659 982
rect 751 978 755 982
rect 839 978 843 982
rect 927 978 931 982
rect 1007 978 1011 982
rect 1087 978 1091 982
rect 1167 978 1171 982
rect 1223 978 1227 982
rect 1287 978 1291 982
rect 1327 946 1331 950
rect 1367 946 1371 950
rect 1423 946 1427 950
rect 1503 946 1507 950
rect 1527 946 1531 950
rect 1607 946 1611 950
rect 1695 946 1699 950
rect 1719 946 1723 950
rect 1831 946 1835 950
rect 1839 946 1843 950
rect 1935 946 1939 950
rect 1967 946 1971 950
rect 2031 946 2035 950
rect 2087 946 2091 950
rect 2127 946 2131 950
rect 2191 946 2195 950
rect 2215 946 2219 950
rect 2287 946 2291 950
rect 2295 946 2299 950
rect 2375 946 2379 950
rect 2383 946 2387 950
rect 2455 946 2459 950
rect 2503 946 2507 950
rect 111 918 115 922
rect 271 918 275 922
rect 287 918 291 922
rect 343 918 347 922
rect 375 918 379 922
rect 423 918 427 922
rect 471 918 475 922
rect 519 918 523 922
rect 567 918 571 922
rect 615 918 619 922
rect 671 918 675 922
rect 711 918 715 922
rect 767 918 771 922
rect 807 918 811 922
rect 855 918 859 922
rect 903 918 907 922
rect 943 918 947 922
rect 991 918 995 922
rect 1023 918 1027 922
rect 1087 918 1091 922
rect 1103 918 1107 922
rect 1183 918 1187 922
rect 1239 918 1243 922
rect 1287 918 1291 922
rect 1327 890 1331 894
rect 1351 890 1355 894
rect 1407 890 1411 894
rect 1431 890 1435 894
rect 1487 890 1491 894
rect 1551 890 1555 894
rect 1591 890 1595 894
rect 1623 890 1627 894
rect 1703 890 1707 894
rect 1791 890 1795 894
rect 1815 890 1819 894
rect 1895 890 1899 894
rect 1919 890 1923 894
rect 2015 890 2019 894
rect 2111 890 2115 894
rect 2143 890 2147 894
rect 2199 890 2203 894
rect 2279 890 2283 894
rect 2359 890 2363 894
rect 2423 890 2427 894
rect 2439 890 2443 894
rect 2503 890 2507 894
rect 111 862 115 866
rect 247 862 251 866
rect 255 862 259 866
rect 311 862 315 866
rect 327 862 331 866
rect 375 862 379 866
rect 407 862 411 866
rect 439 862 443 866
rect 503 862 507 866
rect 567 862 571 866
rect 599 862 603 866
rect 631 862 635 866
rect 695 862 699 866
rect 759 862 763 866
rect 791 862 795 866
rect 831 862 835 866
rect 887 862 891 866
rect 903 862 907 866
rect 975 862 979 866
rect 1071 862 1075 866
rect 1167 862 1171 866
rect 1287 862 1291 866
rect 1327 834 1331 838
rect 1447 834 1451 838
rect 1503 834 1507 838
rect 1567 834 1571 838
rect 1591 834 1595 838
rect 1639 834 1643 838
rect 1647 834 1651 838
rect 1703 834 1707 838
rect 1719 834 1723 838
rect 1767 834 1771 838
rect 1807 834 1811 838
rect 1847 834 1851 838
rect 1911 834 1915 838
rect 1927 834 1931 838
rect 2015 834 2019 838
rect 2031 834 2035 838
rect 2103 834 2107 838
rect 2159 834 2163 838
rect 2191 834 2195 838
rect 2287 834 2291 838
rect 2295 834 2299 838
rect 2383 834 2387 838
rect 2439 834 2443 838
rect 2455 834 2459 838
rect 2503 834 2507 838
rect 111 806 115 810
rect 215 806 219 810
rect 263 806 267 810
rect 303 806 307 810
rect 327 806 331 810
rect 391 806 395 810
rect 455 806 459 810
rect 479 806 483 810
rect 519 806 523 810
rect 559 806 563 810
rect 583 806 587 810
rect 631 806 635 810
rect 647 806 651 810
rect 703 806 707 810
rect 711 806 715 810
rect 767 806 771 810
rect 775 806 779 810
rect 831 806 835 810
rect 847 806 851 810
rect 895 806 899 810
rect 919 806 923 810
rect 967 806 971 810
rect 1039 806 1043 810
rect 1287 806 1291 810
rect 1327 778 1331 782
rect 1567 778 1571 782
rect 1575 778 1579 782
rect 1623 778 1627 782
rect 1631 778 1635 782
rect 1687 778 1691 782
rect 1751 778 1755 782
rect 1759 778 1763 782
rect 1831 778 1835 782
rect 1911 778 1915 782
rect 1919 778 1923 782
rect 1999 778 2003 782
rect 2015 778 2019 782
rect 2087 778 2091 782
rect 2119 778 2123 782
rect 2175 778 2179 782
rect 2231 778 2235 782
rect 2271 778 2275 782
rect 2343 778 2347 782
rect 2367 778 2371 782
rect 2439 778 2443 782
rect 2503 778 2507 782
rect 111 754 115 758
rect 135 754 139 758
rect 199 754 203 758
rect 255 754 259 758
rect 287 754 291 758
rect 375 754 379 758
rect 391 754 395 758
rect 463 754 467 758
rect 519 754 523 758
rect 543 754 547 758
rect 615 754 619 758
rect 647 754 651 758
rect 687 754 691 758
rect 751 754 755 758
rect 775 754 779 758
rect 815 754 819 758
rect 879 754 883 758
rect 903 754 907 758
rect 951 754 955 758
rect 1023 754 1027 758
rect 1039 754 1043 758
rect 1287 754 1291 758
rect 1327 726 1331 730
rect 1367 726 1371 730
rect 1431 726 1435 730
rect 1527 726 1531 730
rect 1583 726 1587 730
rect 1631 726 1635 730
rect 1639 726 1643 730
rect 1703 726 1707 730
rect 1735 726 1739 730
rect 1775 726 1779 730
rect 1839 726 1843 730
rect 1847 726 1851 730
rect 1935 726 1939 730
rect 1943 726 1947 730
rect 2031 726 2035 730
rect 2047 726 2051 730
rect 2135 726 2139 730
rect 2151 726 2155 730
rect 2247 726 2251 730
rect 2255 726 2259 730
rect 2359 726 2363 730
rect 2367 726 2371 730
rect 2455 726 2459 730
rect 2503 726 2507 730
rect 111 702 115 706
rect 151 702 155 706
rect 207 702 211 706
rect 271 702 275 706
rect 295 702 299 706
rect 391 702 395 706
rect 407 702 411 706
rect 503 702 507 706
rect 535 702 539 706
rect 623 702 627 706
rect 663 702 667 706
rect 743 702 747 706
rect 791 702 795 706
rect 871 702 875 706
rect 919 702 923 706
rect 999 702 1003 706
rect 1055 702 1059 706
rect 1127 702 1131 706
rect 1239 702 1243 706
rect 1287 702 1291 706
rect 1327 662 1331 666
rect 1351 662 1355 666
rect 1415 662 1419 666
rect 1511 662 1515 666
rect 1607 662 1611 666
rect 1615 662 1619 666
rect 1711 662 1715 666
rect 1719 662 1723 666
rect 1823 662 1827 666
rect 1927 662 1931 666
rect 1935 662 1939 666
rect 2031 662 2035 666
rect 2055 662 2059 666
rect 2135 662 2139 666
rect 2183 662 2187 666
rect 2239 662 2243 666
rect 2319 662 2323 666
rect 2351 662 2355 666
rect 2439 662 2443 666
rect 2503 662 2507 666
rect 111 646 115 650
rect 135 646 139 650
rect 151 646 155 650
rect 191 646 195 650
rect 263 646 267 650
rect 279 646 283 650
rect 367 646 371 650
rect 375 646 379 650
rect 463 646 467 650
rect 487 646 491 650
rect 559 646 563 650
rect 607 646 611 650
rect 655 646 659 650
rect 727 646 731 650
rect 751 646 755 650
rect 847 646 851 650
rect 855 646 859 650
rect 943 646 947 650
rect 983 646 987 650
rect 1039 646 1043 650
rect 1111 646 1115 650
rect 1143 646 1147 650
rect 1223 646 1227 650
rect 1287 646 1291 650
rect 1327 610 1331 614
rect 1367 610 1371 614
rect 1383 610 1387 614
rect 1431 610 1435 614
rect 1463 610 1467 614
rect 1527 610 1531 614
rect 1551 610 1555 614
rect 1623 610 1627 614
rect 1647 610 1651 614
rect 1727 610 1731 614
rect 1743 610 1747 614
rect 1839 610 1843 614
rect 1847 610 1851 614
rect 1951 610 1955 614
rect 1959 610 1963 614
rect 2071 610 2075 614
rect 2079 610 2083 614
rect 2199 610 2203 614
rect 2207 610 2211 614
rect 2335 610 2339 614
rect 2343 610 2347 614
rect 2455 610 2459 614
rect 2503 610 2507 614
rect 111 594 115 598
rect 151 594 155 598
rect 167 594 171 598
rect 239 594 243 598
rect 279 594 283 598
rect 335 594 339 598
rect 383 594 387 598
rect 431 594 435 598
rect 479 594 483 598
rect 535 594 539 598
rect 575 594 579 598
rect 631 594 635 598
rect 671 594 675 598
rect 727 594 731 598
rect 767 594 771 598
rect 823 594 827 598
rect 863 594 867 598
rect 911 594 915 598
rect 959 594 963 598
rect 999 594 1003 598
rect 1055 594 1059 598
rect 1087 594 1091 598
rect 1159 594 1163 598
rect 1183 594 1187 598
rect 1239 594 1243 598
rect 1287 594 1291 598
rect 1327 558 1331 562
rect 1367 558 1371 562
rect 1375 558 1379 562
rect 1447 558 1451 562
rect 1455 558 1459 562
rect 1535 558 1539 562
rect 1551 558 1555 562
rect 1631 558 1635 562
rect 1647 558 1651 562
rect 1727 558 1731 562
rect 1751 558 1755 562
rect 1831 558 1835 562
rect 1855 558 1859 562
rect 1943 558 1947 562
rect 1959 558 1963 562
rect 2055 558 2059 562
rect 2063 558 2067 562
rect 2151 558 2155 562
rect 2191 558 2195 562
rect 2255 558 2259 562
rect 2327 558 2331 562
rect 2359 558 2363 562
rect 2439 558 2443 562
rect 2503 558 2507 562
rect 111 534 115 538
rect 135 534 139 538
rect 143 534 147 538
rect 223 534 227 538
rect 239 534 243 538
rect 319 534 323 538
rect 335 534 339 538
rect 415 534 419 538
rect 431 534 435 538
rect 519 534 523 538
rect 527 534 531 538
rect 615 534 619 538
rect 623 534 627 538
rect 711 534 715 538
rect 791 534 795 538
rect 807 534 811 538
rect 871 534 875 538
rect 895 534 899 538
rect 951 534 955 538
rect 983 534 987 538
rect 1031 534 1035 538
rect 1071 534 1075 538
rect 1167 534 1171 538
rect 1287 534 1291 538
rect 1327 502 1331 506
rect 1367 502 1371 506
rect 1391 502 1395 506
rect 1455 502 1459 506
rect 1471 502 1475 506
rect 1567 502 1571 506
rect 1575 502 1579 506
rect 1663 502 1667 506
rect 1695 502 1699 506
rect 1767 502 1771 506
rect 1807 502 1811 506
rect 1871 502 1875 506
rect 1919 502 1923 506
rect 1975 502 1979 506
rect 2023 502 2027 506
rect 2071 502 2075 506
rect 2119 502 2123 506
rect 2167 502 2171 506
rect 2207 502 2211 506
rect 2271 502 2275 506
rect 2295 502 2299 506
rect 2375 502 2379 506
rect 2383 502 2387 506
rect 2455 502 2459 506
rect 2503 502 2507 506
rect 111 478 115 482
rect 151 478 155 482
rect 159 478 163 482
rect 207 478 211 482
rect 255 478 259 482
rect 287 478 291 482
rect 351 478 355 482
rect 375 478 379 482
rect 447 478 451 482
rect 463 478 467 482
rect 543 478 547 482
rect 559 478 563 482
rect 639 478 643 482
rect 655 478 659 482
rect 727 478 731 482
rect 751 478 755 482
rect 807 478 811 482
rect 847 478 851 482
rect 887 478 891 482
rect 951 478 955 482
rect 967 478 971 482
rect 1047 478 1051 482
rect 1055 478 1059 482
rect 1159 478 1163 482
rect 1239 478 1243 482
rect 1287 478 1291 482
rect 1327 438 1331 442
rect 1351 438 1355 442
rect 1439 438 1443 442
rect 1559 438 1563 442
rect 1583 438 1587 442
rect 1639 438 1643 442
rect 1679 438 1683 442
rect 1695 438 1699 442
rect 1759 438 1763 442
rect 1791 438 1795 442
rect 1831 438 1835 442
rect 1903 438 1907 442
rect 1911 438 1915 442
rect 1991 438 1995 442
rect 2007 438 2011 442
rect 2079 438 2083 442
rect 2103 438 2107 442
rect 2175 438 2179 442
rect 2191 438 2195 442
rect 2271 438 2275 442
rect 2279 438 2283 442
rect 2367 438 2371 442
rect 2439 438 2443 442
rect 2503 438 2507 442
rect 111 426 115 430
rect 135 426 139 430
rect 191 426 195 430
rect 271 426 275 430
rect 279 426 283 430
rect 359 426 363 430
rect 383 426 387 430
rect 447 426 451 430
rect 495 426 499 430
rect 543 426 547 430
rect 607 426 611 430
rect 639 426 643 430
rect 719 426 723 430
rect 735 426 739 430
rect 831 426 835 430
rect 935 426 939 430
rect 1039 426 1043 430
rect 1143 426 1147 430
rect 1223 426 1227 430
rect 1287 426 1291 430
rect 1327 382 1331 386
rect 1599 382 1603 386
rect 1655 382 1659 386
rect 1679 382 1683 386
rect 1711 382 1715 386
rect 1735 382 1739 386
rect 1775 382 1779 386
rect 1799 382 1803 386
rect 1847 382 1851 386
rect 1871 382 1875 386
rect 1927 382 1931 386
rect 1943 382 1947 386
rect 2007 382 2011 386
rect 2023 382 2027 386
rect 2095 382 2099 386
rect 2111 382 2115 386
rect 2191 382 2195 386
rect 2199 382 2203 386
rect 2287 382 2291 386
rect 2375 382 2379 386
rect 2383 382 2387 386
rect 2455 382 2459 386
rect 2503 382 2507 386
rect 111 370 115 374
rect 151 370 155 374
rect 207 370 211 374
rect 231 370 235 374
rect 295 370 299 374
rect 335 370 339 374
rect 399 370 403 374
rect 439 370 443 374
rect 511 370 515 374
rect 543 370 547 374
rect 623 370 627 374
rect 647 370 651 374
rect 735 370 739 374
rect 751 370 755 374
rect 847 370 851 374
rect 935 370 939 374
rect 951 370 955 374
rect 1015 370 1019 374
rect 1055 370 1059 374
rect 1095 370 1099 374
rect 1159 370 1163 374
rect 1175 370 1179 374
rect 1239 370 1243 374
rect 1287 370 1291 374
rect 1327 322 1331 326
rect 1351 322 1355 326
rect 1455 322 1459 326
rect 1583 322 1587 326
rect 1663 322 1667 326
rect 1711 322 1715 326
rect 1719 322 1723 326
rect 1783 322 1787 326
rect 1839 322 1843 326
rect 1855 322 1859 326
rect 1927 322 1931 326
rect 1951 322 1955 326
rect 2007 322 2011 326
rect 2063 322 2067 326
rect 2095 322 2099 326
rect 2167 322 2171 326
rect 2183 322 2187 326
rect 2263 322 2267 326
rect 2271 322 2275 326
rect 2359 322 2363 326
rect 2439 322 2443 326
rect 2503 322 2507 326
rect 111 314 115 318
rect 135 314 139 318
rect 215 314 219 318
rect 319 314 323 318
rect 423 314 427 318
rect 527 314 531 318
rect 535 314 539 318
rect 631 314 635 318
rect 639 314 643 318
rect 735 314 739 318
rect 743 314 747 318
rect 831 314 835 318
rect 847 314 851 318
rect 919 314 923 318
rect 943 314 947 318
rect 999 314 1003 318
rect 1039 314 1043 318
rect 1079 314 1083 318
rect 1143 314 1147 318
rect 1159 314 1163 318
rect 1223 314 1227 318
rect 1287 314 1291 318
rect 111 262 115 266
rect 151 262 155 266
rect 223 262 227 266
rect 231 262 235 266
rect 319 262 323 266
rect 335 262 339 266
rect 423 262 427 266
rect 439 262 443 266
rect 535 262 539 266
rect 551 262 555 266
rect 647 262 651 266
rect 655 262 659 266
rect 759 262 763 266
rect 863 262 867 266
rect 871 262 875 266
rect 959 262 963 266
rect 983 262 987 266
rect 1055 262 1059 266
rect 1103 262 1107 266
rect 1159 262 1163 266
rect 1223 262 1227 266
rect 1239 262 1243 266
rect 1287 262 1291 266
rect 1327 262 1331 266
rect 1367 262 1371 266
rect 1447 262 1451 266
rect 1471 262 1475 266
rect 1551 262 1555 266
rect 1599 262 1603 266
rect 1655 262 1659 266
rect 1727 262 1731 266
rect 1759 262 1763 266
rect 1855 262 1859 266
rect 1863 262 1867 266
rect 1967 262 1971 266
rect 2071 262 2075 266
rect 2079 262 2083 266
rect 2175 262 2179 266
rect 2183 262 2187 266
rect 2271 262 2275 266
rect 2279 262 2283 266
rect 2375 262 2379 266
rect 2455 262 2459 266
rect 2503 262 2507 266
rect 111 206 115 210
rect 135 206 139 210
rect 183 206 187 210
rect 207 206 211 210
rect 279 206 283 210
rect 303 206 307 210
rect 383 206 387 210
rect 407 206 411 210
rect 487 206 491 210
rect 519 206 523 210
rect 591 206 595 210
rect 631 206 635 210
rect 695 206 699 210
rect 743 206 747 210
rect 799 206 803 210
rect 855 206 859 210
rect 895 206 899 210
rect 967 206 971 210
rect 999 206 1003 210
rect 1087 206 1091 210
rect 1103 206 1107 210
rect 1207 206 1211 210
rect 1287 206 1291 210
rect 1327 206 1331 210
rect 1351 206 1355 210
rect 1407 206 1411 210
rect 1431 206 1435 210
rect 1471 206 1475 210
rect 1535 206 1539 210
rect 1551 206 1555 210
rect 1639 206 1643 210
rect 1719 206 1723 210
rect 1743 206 1747 210
rect 1807 206 1811 210
rect 1847 206 1851 210
rect 1895 206 1899 210
rect 1951 206 1955 210
rect 1991 206 1995 210
rect 2055 206 2059 210
rect 2103 206 2107 210
rect 2159 206 2163 210
rect 2215 206 2219 210
rect 2255 206 2259 210
rect 2335 206 2339 210
rect 2359 206 2363 210
rect 2439 206 2443 210
rect 2503 206 2507 210
rect 111 146 115 150
rect 151 146 155 150
rect 199 146 203 150
rect 207 146 211 150
rect 263 146 267 150
rect 295 146 299 150
rect 319 146 323 150
rect 375 146 379 150
rect 399 146 403 150
rect 431 146 435 150
rect 487 146 491 150
rect 503 146 507 150
rect 543 146 547 150
rect 599 146 603 150
rect 607 146 611 150
rect 655 146 659 150
rect 711 146 715 150
rect 767 146 771 150
rect 815 146 819 150
rect 831 146 835 150
rect 895 146 899 150
rect 911 146 915 150
rect 959 146 963 150
rect 1015 146 1019 150
rect 1023 146 1027 150
rect 1087 146 1091 150
rect 1119 146 1123 150
rect 1151 146 1155 150
rect 1287 146 1291 150
rect 1327 134 1331 138
rect 1367 134 1371 138
rect 1423 134 1427 138
rect 1479 134 1483 138
rect 1487 134 1491 138
rect 1535 134 1539 138
rect 1567 134 1571 138
rect 1591 134 1595 138
rect 1647 134 1651 138
rect 1655 134 1659 138
rect 1703 134 1707 138
rect 1735 134 1739 138
rect 1759 134 1763 138
rect 1823 134 1827 138
rect 1879 134 1883 138
rect 1911 134 1915 138
rect 1943 134 1947 138
rect 2007 134 2011 138
rect 2071 134 2075 138
rect 2119 134 2123 138
rect 2143 134 2147 138
rect 2223 134 2227 138
rect 2231 134 2235 138
rect 2303 134 2307 138
rect 2351 134 2355 138
rect 2391 134 2395 138
rect 2455 134 2459 138
rect 2503 134 2507 138
rect 111 94 115 98
rect 135 94 139 98
rect 191 94 195 98
rect 247 94 251 98
rect 303 94 307 98
rect 359 94 363 98
rect 415 94 419 98
rect 471 94 475 98
rect 527 94 531 98
rect 583 94 587 98
rect 639 94 643 98
rect 695 94 699 98
rect 751 94 755 98
rect 815 94 819 98
rect 879 94 883 98
rect 943 94 947 98
rect 1007 94 1011 98
rect 1071 94 1075 98
rect 1135 94 1139 98
rect 1287 94 1291 98
rect 1327 82 1331 86
rect 1351 82 1355 86
rect 1407 82 1411 86
rect 1463 82 1467 86
rect 1519 82 1523 86
rect 1575 82 1579 86
rect 1631 82 1635 86
rect 1687 82 1691 86
rect 1743 82 1747 86
rect 1807 82 1811 86
rect 1863 82 1867 86
rect 1927 82 1931 86
rect 1991 82 1995 86
rect 2055 82 2059 86
rect 2127 82 2131 86
rect 2207 82 2211 86
rect 2287 82 2291 86
rect 2375 82 2379 86
rect 2439 82 2443 86
rect 2503 82 2507 86
<< m4 >>
rect 84 2577 85 2583
rect 91 2582 1299 2583
rect 91 2578 111 2582
rect 115 2578 135 2582
rect 139 2578 191 2582
rect 195 2578 247 2582
rect 251 2578 303 2582
rect 307 2578 359 2582
rect 363 2578 1287 2582
rect 1291 2578 1299 2582
rect 91 2577 1299 2578
rect 1305 2577 1306 2583
rect 1298 2557 1299 2563
rect 1305 2562 2527 2563
rect 1305 2558 1327 2562
rect 1331 2558 1495 2562
rect 1499 2558 1551 2562
rect 1555 2558 1607 2562
rect 1611 2558 1663 2562
rect 1667 2558 1719 2562
rect 1723 2558 1775 2562
rect 1779 2558 1831 2562
rect 1835 2558 1887 2562
rect 1891 2558 1943 2562
rect 1947 2558 1999 2562
rect 2003 2558 2055 2562
rect 2059 2558 2111 2562
rect 2115 2558 2167 2562
rect 2171 2558 2503 2562
rect 2507 2558 2527 2562
rect 1305 2557 2527 2558
rect 2533 2557 2534 2563
rect 96 2525 97 2531
rect 103 2530 1311 2531
rect 103 2526 111 2530
rect 115 2526 151 2530
rect 155 2526 207 2530
rect 211 2526 223 2530
rect 227 2526 263 2530
rect 267 2526 279 2530
rect 283 2526 319 2530
rect 323 2526 343 2530
rect 347 2526 375 2530
rect 379 2526 415 2530
rect 419 2526 487 2530
rect 491 2526 551 2530
rect 555 2526 615 2530
rect 619 2526 679 2530
rect 683 2526 743 2530
rect 747 2526 807 2530
rect 811 2526 871 2530
rect 875 2526 935 2530
rect 939 2526 999 2530
rect 1003 2526 1063 2530
rect 1067 2526 1287 2530
rect 1291 2526 1311 2530
rect 103 2525 1311 2526
rect 1317 2525 1318 2531
rect 1310 2505 1311 2511
rect 1317 2510 2539 2511
rect 1317 2506 1327 2510
rect 1331 2506 1511 2510
rect 1515 2506 1543 2510
rect 1547 2506 1567 2510
rect 1571 2506 1607 2510
rect 1611 2506 1623 2510
rect 1627 2506 1679 2510
rect 1683 2506 1735 2510
rect 1739 2506 1751 2510
rect 1755 2506 1791 2510
rect 1795 2506 1823 2510
rect 1827 2506 1847 2510
rect 1851 2506 1895 2510
rect 1899 2506 1903 2510
rect 1907 2506 1959 2510
rect 1963 2506 1967 2510
rect 1971 2506 2015 2510
rect 2019 2506 2039 2510
rect 2043 2506 2071 2510
rect 2075 2506 2111 2510
rect 2115 2506 2127 2510
rect 2131 2506 2183 2510
rect 2187 2506 2503 2510
rect 2507 2506 2539 2510
rect 1317 2505 2539 2506
rect 2545 2505 2546 2511
rect 84 2465 85 2471
rect 91 2470 1299 2471
rect 91 2466 111 2470
rect 115 2466 167 2470
rect 171 2466 207 2470
rect 211 2466 223 2470
rect 227 2466 263 2470
rect 267 2466 279 2470
rect 283 2466 327 2470
rect 331 2466 335 2470
rect 339 2466 391 2470
rect 395 2466 399 2470
rect 403 2466 447 2470
rect 451 2466 471 2470
rect 475 2466 503 2470
rect 507 2466 535 2470
rect 539 2466 559 2470
rect 563 2466 599 2470
rect 603 2466 615 2470
rect 619 2466 663 2470
rect 667 2466 671 2470
rect 675 2466 727 2470
rect 731 2466 783 2470
rect 787 2466 791 2470
rect 795 2466 839 2470
rect 843 2466 855 2470
rect 859 2466 895 2470
rect 899 2466 919 2470
rect 923 2466 951 2470
rect 955 2466 983 2470
rect 987 2466 1007 2470
rect 1011 2466 1047 2470
rect 1051 2466 1063 2470
rect 1067 2466 1287 2470
rect 1291 2466 1299 2470
rect 91 2465 1299 2466
rect 1305 2465 1306 2471
rect 1298 2449 1299 2455
rect 1305 2454 2527 2455
rect 1305 2450 1327 2454
rect 1331 2450 1527 2454
rect 1531 2450 1543 2454
rect 1547 2450 1591 2454
rect 1595 2450 1607 2454
rect 1611 2450 1663 2454
rect 1667 2450 1671 2454
rect 1675 2450 1735 2454
rect 1739 2450 1743 2454
rect 1747 2450 1807 2454
rect 1811 2450 1815 2454
rect 1819 2450 1879 2454
rect 1883 2450 1951 2454
rect 1955 2450 2023 2454
rect 2027 2450 2095 2454
rect 2099 2450 2167 2454
rect 2171 2450 2503 2454
rect 2507 2450 2527 2454
rect 1305 2449 2527 2450
rect 2533 2449 2534 2455
rect 96 2401 97 2407
rect 103 2406 1311 2407
rect 103 2402 111 2406
rect 115 2402 183 2406
rect 187 2402 239 2406
rect 243 2402 295 2406
rect 299 2402 351 2406
rect 355 2402 407 2406
rect 411 2402 463 2406
rect 467 2402 519 2406
rect 523 2402 575 2406
rect 579 2402 631 2406
rect 635 2402 687 2406
rect 691 2402 743 2406
rect 747 2402 799 2406
rect 803 2402 855 2406
rect 859 2402 911 2406
rect 915 2402 967 2406
rect 971 2402 1023 2406
rect 1027 2402 1079 2406
rect 1083 2402 1287 2406
rect 1291 2402 1311 2406
rect 103 2401 1311 2402
rect 1317 2401 1318 2407
rect 1310 2399 1318 2401
rect 1310 2393 1311 2399
rect 1317 2398 2539 2399
rect 1317 2394 1327 2398
rect 1331 2394 1559 2398
rect 1563 2394 1567 2398
rect 1571 2394 1623 2398
rect 1627 2394 1679 2398
rect 1683 2394 1687 2398
rect 1691 2394 1735 2398
rect 1739 2394 1759 2398
rect 1763 2394 1791 2398
rect 1795 2394 1831 2398
rect 1835 2394 1855 2398
rect 1859 2394 1895 2398
rect 1899 2394 1919 2398
rect 1923 2394 1967 2398
rect 1971 2394 1983 2398
rect 1987 2394 2039 2398
rect 2043 2394 2047 2398
rect 2051 2394 2111 2398
rect 2115 2394 2183 2398
rect 2187 2394 2503 2398
rect 2507 2394 2539 2398
rect 1317 2393 2539 2394
rect 2545 2393 2546 2399
rect 84 2341 85 2347
rect 91 2346 1299 2347
rect 91 2342 111 2346
rect 115 2342 319 2346
rect 323 2342 391 2346
rect 395 2342 463 2346
rect 467 2342 503 2346
rect 507 2342 535 2346
rect 539 2342 559 2346
rect 563 2342 607 2346
rect 611 2342 615 2346
rect 619 2342 671 2346
rect 675 2342 679 2346
rect 683 2342 743 2346
rect 747 2342 807 2346
rect 811 2342 863 2346
rect 867 2342 927 2346
rect 931 2342 991 2346
rect 995 2342 1055 2346
rect 1059 2342 1111 2346
rect 1115 2342 1167 2346
rect 1171 2342 1223 2346
rect 1227 2342 1287 2346
rect 1291 2342 1299 2346
rect 91 2341 1299 2342
rect 1305 2341 1306 2347
rect 1298 2339 1306 2341
rect 1298 2333 1299 2339
rect 1305 2338 2527 2339
rect 1305 2334 1327 2338
rect 1331 2334 1471 2338
rect 1475 2334 1535 2338
rect 1539 2334 1551 2338
rect 1555 2334 1607 2338
rect 1611 2334 1663 2338
rect 1667 2334 1687 2338
rect 1691 2334 1719 2338
rect 1723 2334 1759 2338
rect 1763 2334 1775 2338
rect 1779 2334 1831 2338
rect 1835 2334 1839 2338
rect 1843 2334 1903 2338
rect 1907 2334 1967 2338
rect 1971 2334 1983 2338
rect 1987 2334 2031 2338
rect 2035 2334 2063 2338
rect 2067 2334 2095 2338
rect 2099 2334 2143 2338
rect 2147 2334 2503 2338
rect 2507 2334 2527 2338
rect 1305 2333 2527 2334
rect 2533 2333 2534 2339
rect 96 2281 97 2287
rect 103 2286 1311 2287
rect 103 2282 111 2286
rect 115 2282 175 2286
rect 179 2282 271 2286
rect 275 2282 335 2286
rect 339 2282 375 2286
rect 379 2282 407 2286
rect 411 2282 479 2286
rect 483 2282 551 2286
rect 555 2282 591 2286
rect 595 2282 623 2286
rect 627 2282 695 2286
rect 699 2282 703 2286
rect 707 2282 759 2286
rect 763 2282 807 2286
rect 811 2282 823 2286
rect 827 2282 879 2286
rect 883 2282 911 2286
rect 915 2282 943 2286
rect 947 2282 1007 2286
rect 1011 2282 1015 2286
rect 1019 2282 1071 2286
rect 1075 2282 1127 2286
rect 1131 2282 1183 2286
rect 1187 2282 1239 2286
rect 1243 2282 1287 2286
rect 1291 2282 1311 2286
rect 103 2281 1311 2282
rect 1317 2286 2546 2287
rect 1317 2282 1327 2286
rect 1331 2282 1383 2286
rect 1387 2282 1479 2286
rect 1483 2282 1487 2286
rect 1491 2282 1551 2286
rect 1555 2282 1583 2286
rect 1587 2282 1623 2286
rect 1627 2282 1687 2286
rect 1691 2282 1703 2286
rect 1707 2282 1775 2286
rect 1779 2282 1791 2286
rect 1795 2282 1847 2286
rect 1851 2282 1903 2286
rect 1907 2282 1919 2286
rect 1923 2282 1999 2286
rect 2003 2282 2015 2286
rect 2019 2282 2079 2286
rect 2083 2282 2127 2286
rect 2131 2282 2159 2286
rect 2163 2282 2239 2286
rect 2243 2282 2503 2286
rect 2507 2282 2546 2286
rect 1317 2281 2546 2282
rect 84 2229 85 2235
rect 91 2234 1299 2235
rect 91 2230 111 2234
rect 115 2230 143 2234
rect 147 2230 159 2234
rect 163 2230 231 2234
rect 235 2230 255 2234
rect 259 2230 319 2234
rect 323 2230 359 2234
rect 363 2230 415 2234
rect 419 2230 463 2234
rect 467 2230 519 2234
rect 523 2230 575 2234
rect 579 2230 623 2234
rect 627 2230 687 2234
rect 691 2230 727 2234
rect 731 2230 791 2234
rect 795 2230 831 2234
rect 835 2230 895 2234
rect 899 2230 935 2234
rect 939 2230 999 2234
rect 1003 2230 1039 2234
rect 1043 2230 1111 2234
rect 1115 2230 1143 2234
rect 1147 2230 1223 2234
rect 1227 2230 1287 2234
rect 1291 2230 1299 2234
rect 91 2229 1299 2230
rect 1305 2234 2534 2235
rect 1305 2230 1327 2234
rect 1331 2230 1367 2234
rect 1371 2230 1463 2234
rect 1467 2230 1487 2234
rect 1491 2230 1567 2234
rect 1571 2230 1607 2234
rect 1611 2230 1671 2234
rect 1675 2230 1719 2234
rect 1723 2230 1775 2234
rect 1779 2230 1815 2234
rect 1819 2230 1887 2234
rect 1891 2230 1903 2234
rect 1907 2230 1983 2234
rect 1987 2230 1999 2234
rect 2003 2230 2055 2234
rect 2059 2230 2111 2234
rect 2115 2230 2127 2234
rect 2131 2230 2191 2234
rect 2195 2230 2223 2234
rect 2227 2230 2255 2234
rect 2259 2230 2319 2234
rect 2323 2230 2383 2234
rect 2387 2230 2439 2234
rect 2443 2230 2503 2234
rect 2507 2230 2534 2234
rect 1305 2229 2534 2230
rect 96 2177 97 2183
rect 103 2182 1311 2183
rect 103 2178 111 2182
rect 115 2178 159 2182
rect 163 2178 247 2182
rect 251 2178 255 2182
rect 259 2178 335 2182
rect 339 2178 351 2182
rect 355 2178 431 2182
rect 435 2178 455 2182
rect 459 2178 535 2182
rect 539 2178 559 2182
rect 563 2178 639 2182
rect 643 2178 663 2182
rect 667 2178 743 2182
rect 747 2178 767 2182
rect 771 2178 847 2182
rect 851 2178 863 2182
rect 867 2178 951 2182
rect 955 2178 959 2182
rect 963 2178 1055 2182
rect 1059 2178 1159 2182
rect 1163 2178 1239 2182
rect 1243 2178 1287 2182
rect 1291 2178 1311 2182
rect 103 2177 1311 2178
rect 1317 2177 1318 2183
rect 1310 2157 1311 2163
rect 1317 2162 2539 2163
rect 1317 2158 1327 2162
rect 1331 2158 1383 2162
rect 1387 2158 1407 2162
rect 1411 2158 1503 2162
rect 1507 2158 1623 2162
rect 1627 2158 1735 2162
rect 1739 2158 1815 2162
rect 1819 2158 1831 2162
rect 1835 2158 1919 2162
rect 1923 2158 1991 2162
rect 1995 2158 1999 2162
rect 2003 2158 2071 2162
rect 2075 2158 2143 2162
rect 2147 2158 2159 2162
rect 2163 2158 2207 2162
rect 2211 2158 2271 2162
rect 2275 2158 2319 2162
rect 2323 2158 2335 2162
rect 2339 2158 2399 2162
rect 2403 2158 2455 2162
rect 2459 2158 2503 2162
rect 2507 2158 2539 2162
rect 1317 2157 2539 2158
rect 2545 2157 2546 2163
rect 84 2125 85 2131
rect 91 2130 1299 2131
rect 91 2126 111 2130
rect 115 2126 239 2130
rect 243 2126 303 2130
rect 307 2126 335 2130
rect 339 2126 359 2130
rect 363 2126 423 2130
rect 427 2126 439 2130
rect 443 2126 487 2130
rect 491 2126 543 2130
rect 547 2126 559 2130
rect 563 2126 631 2130
rect 635 2126 647 2130
rect 651 2126 711 2130
rect 715 2126 751 2130
rect 755 2126 799 2130
rect 803 2126 847 2130
rect 851 2126 887 2130
rect 891 2126 943 2130
rect 947 2126 975 2130
rect 979 2126 1039 2130
rect 1043 2126 1063 2130
rect 1067 2126 1143 2130
rect 1147 2126 1151 2130
rect 1155 2126 1223 2130
rect 1227 2126 1287 2130
rect 1291 2126 1299 2130
rect 91 2125 1299 2126
rect 1305 2125 1306 2131
rect 1298 2105 1299 2111
rect 1305 2110 2527 2111
rect 1305 2106 1327 2110
rect 1331 2106 1383 2110
rect 1387 2106 1391 2110
rect 1395 2106 1551 2110
rect 1555 2106 1607 2110
rect 1611 2106 1711 2110
rect 1715 2106 1799 2110
rect 1803 2106 1855 2110
rect 1859 2106 1975 2110
rect 1979 2106 1991 2110
rect 1995 2106 2119 2110
rect 2123 2106 2143 2110
rect 2147 2106 2239 2110
rect 2243 2106 2303 2110
rect 2307 2106 2367 2110
rect 2371 2106 2439 2110
rect 2443 2106 2503 2110
rect 2507 2106 2527 2110
rect 1305 2105 2527 2106
rect 2533 2105 2534 2111
rect 96 2069 97 2075
rect 103 2074 1311 2075
rect 103 2070 111 2074
rect 115 2070 319 2074
rect 323 2070 375 2074
rect 379 2070 399 2074
rect 403 2070 439 2074
rect 443 2070 455 2074
rect 459 2070 503 2074
rect 507 2070 511 2074
rect 515 2070 575 2074
rect 579 2070 639 2074
rect 643 2070 647 2074
rect 651 2070 711 2074
rect 715 2070 727 2074
rect 731 2070 791 2074
rect 795 2070 815 2074
rect 819 2070 863 2074
rect 867 2070 903 2074
rect 907 2070 943 2074
rect 947 2070 991 2074
rect 995 2070 1023 2074
rect 1027 2070 1079 2074
rect 1083 2070 1103 2074
rect 1107 2070 1167 2074
rect 1171 2070 1183 2074
rect 1187 2070 1239 2074
rect 1243 2070 1287 2074
rect 1291 2070 1311 2074
rect 103 2069 1311 2070
rect 1317 2069 1318 2075
rect 1310 2049 1311 2055
rect 1317 2054 2539 2055
rect 1317 2050 1327 2054
rect 1331 2050 1399 2054
rect 1403 2050 1447 2054
rect 1451 2050 1551 2054
rect 1555 2050 1567 2054
rect 1571 2050 1655 2054
rect 1659 2050 1727 2054
rect 1731 2050 1751 2054
rect 1755 2050 1839 2054
rect 1843 2050 1871 2054
rect 1875 2050 1927 2054
rect 1931 2050 2007 2054
rect 2011 2050 2023 2054
rect 2027 2050 2119 2054
rect 2123 2050 2135 2054
rect 2139 2050 2255 2054
rect 2259 2050 2383 2054
rect 2387 2050 2503 2054
rect 2507 2050 2539 2054
rect 1317 2049 2539 2050
rect 2545 2049 2546 2055
rect 84 2013 85 2019
rect 91 2018 1299 2019
rect 91 2014 111 2018
rect 115 2014 231 2018
rect 235 2014 287 2018
rect 291 2014 359 2018
rect 363 2014 383 2018
rect 387 2014 439 2018
rect 443 2014 495 2018
rect 499 2014 535 2018
rect 539 2014 559 2018
rect 563 2014 623 2018
rect 627 2014 631 2018
rect 635 2014 695 2018
rect 699 2014 735 2018
rect 739 2014 775 2018
rect 779 2014 847 2018
rect 851 2014 927 2018
rect 931 2014 959 2018
rect 963 2014 1007 2018
rect 1011 2014 1079 2018
rect 1083 2014 1087 2018
rect 1091 2014 1167 2018
rect 1171 2014 1199 2018
rect 1203 2014 1223 2018
rect 1227 2014 1287 2018
rect 1291 2014 1299 2018
rect 91 2013 1299 2014
rect 1305 2013 1306 2019
rect 1298 1993 1299 1999
rect 1305 1998 2527 1999
rect 1305 1994 1327 1998
rect 1331 1994 1431 1998
rect 1435 1994 1455 1998
rect 1459 1994 1511 1998
rect 1515 1994 1535 1998
rect 1539 1994 1575 1998
rect 1579 1994 1639 1998
rect 1643 1994 1703 1998
rect 1707 1994 1735 1998
rect 1739 1994 1767 1998
rect 1771 1994 1823 1998
rect 1827 1994 1831 1998
rect 1835 1994 1895 1998
rect 1899 1994 1911 1998
rect 1915 1994 1959 1998
rect 1963 1994 2007 1998
rect 2011 1994 2031 1998
rect 2035 1994 2103 1998
rect 2107 1994 2503 1998
rect 2507 1994 2527 1998
rect 1305 1993 2527 1994
rect 2533 1993 2534 1999
rect 96 1957 97 1963
rect 103 1962 1311 1963
rect 103 1958 111 1962
rect 115 1958 151 1962
rect 155 1958 215 1962
rect 219 1958 247 1962
rect 251 1958 303 1962
rect 307 1958 319 1962
rect 323 1958 375 1962
rect 379 1958 439 1962
rect 443 1958 455 1962
rect 459 1958 551 1962
rect 555 1958 583 1962
rect 587 1958 647 1962
rect 651 1958 743 1962
rect 747 1958 751 1962
rect 755 1958 863 1962
rect 867 1958 919 1962
rect 923 1958 975 1962
rect 979 1958 1095 1962
rect 1099 1958 1215 1962
rect 1219 1958 1287 1962
rect 1291 1958 1311 1962
rect 103 1957 1311 1958
rect 1317 1957 1318 1963
rect 1310 1937 1311 1943
rect 1317 1942 2539 1943
rect 1317 1938 1327 1942
rect 1331 1938 1471 1942
rect 1475 1938 1527 1942
rect 1531 1938 1567 1942
rect 1571 1938 1591 1942
rect 1595 1938 1631 1942
rect 1635 1938 1655 1942
rect 1659 1938 1703 1942
rect 1707 1938 1719 1942
rect 1723 1938 1775 1942
rect 1779 1938 1783 1942
rect 1787 1938 1847 1942
rect 1851 1938 1911 1942
rect 1915 1938 1919 1942
rect 1923 1938 1975 1942
rect 1979 1938 1999 1942
rect 2003 1938 2047 1942
rect 2051 1938 2087 1942
rect 2091 1938 2183 1942
rect 2187 1938 2279 1942
rect 2283 1938 2375 1942
rect 2379 1938 2455 1942
rect 2459 1938 2503 1942
rect 2507 1938 2539 1942
rect 1317 1937 2539 1938
rect 2545 1937 2546 1943
rect 84 1897 85 1903
rect 91 1902 1299 1903
rect 91 1898 111 1902
rect 115 1898 135 1902
rect 139 1898 191 1902
rect 195 1898 199 1902
rect 203 1898 271 1902
rect 275 1898 303 1902
rect 307 1898 359 1902
rect 363 1898 423 1902
rect 427 1898 455 1902
rect 459 1898 543 1902
rect 547 1898 567 1902
rect 571 1898 631 1902
rect 635 1898 719 1902
rect 723 1898 727 1902
rect 731 1898 799 1902
rect 803 1898 871 1902
rect 875 1898 903 1902
rect 907 1898 943 1902
rect 947 1898 1015 1902
rect 1019 1898 1079 1902
rect 1083 1898 1087 1902
rect 1091 1898 1159 1902
rect 1163 1898 1287 1902
rect 1291 1898 1299 1902
rect 91 1897 1299 1898
rect 1305 1897 1306 1903
rect 1298 1881 1299 1887
rect 1305 1886 2527 1887
rect 1305 1882 1327 1886
rect 1331 1882 1551 1886
rect 1555 1882 1607 1886
rect 1611 1882 1615 1886
rect 1619 1882 1663 1886
rect 1667 1882 1687 1886
rect 1691 1882 1727 1886
rect 1731 1882 1759 1886
rect 1763 1882 1799 1886
rect 1803 1882 1831 1886
rect 1835 1882 1871 1886
rect 1875 1882 1903 1886
rect 1907 1882 1943 1886
rect 1947 1882 1983 1886
rect 1987 1882 2007 1886
rect 2011 1882 2071 1886
rect 2075 1882 2135 1886
rect 2139 1882 2167 1886
rect 2171 1882 2199 1886
rect 2203 1882 2263 1886
rect 2267 1882 2327 1886
rect 2331 1882 2359 1886
rect 2363 1882 2383 1886
rect 2387 1882 2439 1886
rect 2443 1882 2503 1886
rect 2507 1882 2527 1886
rect 1305 1881 2527 1882
rect 2533 1881 2534 1887
rect 96 1845 97 1851
rect 103 1850 1311 1851
rect 103 1846 111 1850
rect 115 1846 151 1850
rect 155 1846 207 1850
rect 211 1846 287 1850
rect 291 1846 295 1850
rect 299 1846 375 1850
rect 379 1846 391 1850
rect 395 1846 471 1850
rect 475 1846 495 1850
rect 499 1846 559 1850
rect 563 1846 591 1850
rect 595 1846 647 1850
rect 651 1846 687 1850
rect 691 1846 735 1850
rect 739 1846 775 1850
rect 779 1846 815 1850
rect 819 1846 855 1850
rect 859 1846 887 1850
rect 891 1846 927 1850
rect 931 1846 959 1850
rect 963 1846 999 1850
rect 1003 1846 1031 1850
rect 1035 1846 1079 1850
rect 1083 1846 1103 1850
rect 1107 1846 1159 1850
rect 1163 1846 1175 1850
rect 1179 1846 1287 1850
rect 1291 1846 1311 1850
rect 103 1845 1311 1846
rect 1317 1845 1318 1851
rect 1310 1825 1311 1831
rect 1317 1830 2539 1831
rect 1317 1826 1327 1830
rect 1331 1826 1623 1830
rect 1627 1826 1631 1830
rect 1635 1826 1679 1830
rect 1683 1826 1719 1830
rect 1723 1826 1743 1830
rect 1747 1826 1815 1830
rect 1819 1826 1887 1830
rect 1891 1826 1927 1830
rect 1931 1826 1959 1830
rect 1963 1826 2023 1830
rect 2027 1826 2055 1830
rect 2059 1826 2087 1830
rect 2091 1826 2151 1830
rect 2155 1826 2191 1830
rect 2195 1826 2215 1830
rect 2219 1826 2279 1830
rect 2283 1826 2335 1830
rect 2339 1826 2343 1830
rect 2347 1826 2399 1830
rect 2403 1826 2455 1830
rect 2459 1826 2503 1830
rect 2507 1826 2539 1830
rect 1317 1825 2539 1826
rect 2545 1825 2546 1831
rect 84 1781 85 1787
rect 91 1786 1299 1787
rect 91 1782 111 1786
rect 115 1782 135 1786
rect 139 1782 191 1786
rect 195 1782 199 1786
rect 203 1782 279 1786
rect 283 1782 295 1786
rect 299 1782 375 1786
rect 379 1782 399 1786
rect 403 1782 479 1786
rect 483 1782 503 1786
rect 507 1782 575 1786
rect 579 1782 607 1786
rect 611 1782 671 1786
rect 675 1782 703 1786
rect 707 1782 759 1786
rect 763 1782 799 1786
rect 803 1782 839 1786
rect 843 1782 887 1786
rect 891 1782 911 1786
rect 915 1782 975 1786
rect 979 1782 983 1786
rect 987 1782 1063 1786
rect 1067 1782 1143 1786
rect 1147 1782 1151 1786
rect 1155 1782 1287 1786
rect 1291 1782 1299 1786
rect 91 1781 1299 1782
rect 1305 1781 1306 1787
rect 1298 1779 1306 1781
rect 1298 1773 1299 1779
rect 1305 1778 2527 1779
rect 1305 1774 1327 1778
rect 1331 1774 1527 1778
rect 1531 1774 1607 1778
rect 1611 1774 1615 1778
rect 1619 1774 1695 1778
rect 1699 1774 1703 1778
rect 1707 1774 1791 1778
rect 1795 1774 1799 1778
rect 1803 1774 1879 1778
rect 1883 1774 1911 1778
rect 1915 1774 1967 1778
rect 1971 1774 2039 1778
rect 2043 1774 2055 1778
rect 2059 1774 2135 1778
rect 2139 1774 2175 1778
rect 2179 1774 2215 1778
rect 2219 1774 2295 1778
rect 2299 1774 2319 1778
rect 2323 1774 2375 1778
rect 2379 1774 2439 1778
rect 2443 1774 2503 1778
rect 2507 1774 2527 1778
rect 1305 1773 2527 1774
rect 2533 1773 2534 1779
rect 96 1725 97 1731
rect 103 1730 1311 1731
rect 103 1726 111 1730
rect 115 1726 151 1730
rect 155 1726 167 1730
rect 171 1726 215 1730
rect 219 1726 239 1730
rect 243 1726 311 1730
rect 315 1726 319 1730
rect 323 1726 407 1730
rect 411 1726 415 1730
rect 419 1726 503 1730
rect 507 1726 519 1730
rect 523 1726 607 1730
rect 611 1726 623 1730
rect 627 1726 711 1730
rect 715 1726 719 1730
rect 723 1726 815 1730
rect 819 1726 823 1730
rect 827 1726 903 1730
rect 907 1726 935 1730
rect 939 1726 991 1730
rect 995 1726 1047 1730
rect 1051 1726 1079 1730
rect 1083 1726 1159 1730
rect 1163 1726 1167 1730
rect 1171 1726 1287 1730
rect 1291 1726 1311 1730
rect 103 1725 1311 1726
rect 1317 1725 1318 1731
rect 1310 1723 1318 1725
rect 1310 1717 1311 1723
rect 1317 1722 2539 1723
rect 1317 1718 1327 1722
rect 1331 1718 1399 1722
rect 1403 1718 1463 1722
rect 1467 1718 1543 1722
rect 1547 1718 1623 1722
rect 1627 1718 1631 1722
rect 1635 1718 1711 1722
rect 1715 1718 1727 1722
rect 1731 1718 1807 1722
rect 1811 1718 1823 1722
rect 1827 1718 1895 1722
rect 1899 1718 1919 1722
rect 1923 1718 1983 1722
rect 1987 1718 2015 1722
rect 2019 1718 2071 1722
rect 2075 1718 2111 1722
rect 2115 1718 2151 1722
rect 2155 1718 2199 1722
rect 2203 1718 2231 1722
rect 2235 1718 2287 1722
rect 2291 1718 2311 1722
rect 2315 1718 2383 1722
rect 2387 1718 2391 1722
rect 2395 1718 2455 1722
rect 2459 1718 2503 1722
rect 2507 1718 2539 1722
rect 1317 1717 2539 1718
rect 2545 1717 2546 1723
rect 84 1669 85 1675
rect 91 1674 1299 1675
rect 91 1670 111 1674
rect 115 1670 151 1674
rect 155 1670 223 1674
rect 227 1670 255 1674
rect 259 1670 303 1674
rect 307 1670 319 1674
rect 323 1670 391 1674
rect 395 1670 399 1674
rect 403 1670 487 1674
rect 491 1670 575 1674
rect 579 1670 591 1674
rect 595 1670 671 1674
rect 675 1670 695 1674
rect 699 1670 767 1674
rect 771 1670 807 1674
rect 811 1670 863 1674
rect 867 1670 919 1674
rect 923 1670 959 1674
rect 963 1670 1031 1674
rect 1035 1670 1063 1674
rect 1067 1670 1143 1674
rect 1147 1670 1167 1674
rect 1171 1670 1287 1674
rect 1291 1670 1299 1674
rect 91 1669 1299 1670
rect 1305 1669 1306 1675
rect 1298 1667 1306 1669
rect 1298 1661 1299 1667
rect 1305 1666 2527 1667
rect 1305 1662 1327 1666
rect 1331 1662 1351 1666
rect 1355 1662 1383 1666
rect 1387 1662 1407 1666
rect 1411 1662 1447 1666
rect 1451 1662 1495 1666
rect 1499 1662 1527 1666
rect 1531 1662 1583 1666
rect 1587 1662 1615 1666
rect 1619 1662 1679 1666
rect 1683 1662 1711 1666
rect 1715 1662 1783 1666
rect 1787 1662 1807 1666
rect 1811 1662 1895 1666
rect 1899 1662 1903 1666
rect 1907 1662 1999 1666
rect 2003 1662 2023 1666
rect 2027 1662 2095 1666
rect 2099 1662 2159 1666
rect 2163 1662 2183 1666
rect 2187 1662 2271 1666
rect 2275 1662 2303 1666
rect 2307 1662 2367 1666
rect 2371 1662 2439 1666
rect 2443 1662 2503 1666
rect 2507 1662 2527 1666
rect 1305 1661 2527 1662
rect 2533 1661 2534 1667
rect 96 1613 97 1619
rect 103 1618 1311 1619
rect 103 1614 111 1618
rect 115 1614 271 1618
rect 275 1614 303 1618
rect 307 1614 335 1618
rect 339 1614 359 1618
rect 363 1614 415 1618
rect 419 1614 431 1618
rect 435 1614 503 1618
rect 507 1614 511 1618
rect 515 1614 591 1618
rect 595 1614 599 1618
rect 603 1614 687 1618
rect 691 1614 695 1618
rect 699 1614 783 1618
rect 787 1614 791 1618
rect 795 1614 879 1618
rect 883 1614 895 1618
rect 899 1614 975 1618
rect 979 1614 1007 1618
rect 1011 1614 1079 1618
rect 1083 1614 1119 1618
rect 1123 1614 1183 1618
rect 1187 1614 1287 1618
rect 1291 1614 1311 1618
rect 103 1613 1311 1614
rect 1317 1615 1318 1619
rect 1317 1614 2546 1615
rect 1317 1613 1327 1614
rect 1310 1610 1327 1613
rect 1331 1610 1367 1614
rect 1371 1610 1423 1614
rect 1427 1610 1479 1614
rect 1483 1610 1511 1614
rect 1515 1610 1559 1614
rect 1563 1610 1599 1614
rect 1603 1610 1639 1614
rect 1643 1610 1695 1614
rect 1699 1610 1719 1614
rect 1723 1610 1791 1614
rect 1795 1610 1799 1614
rect 1803 1610 1871 1614
rect 1875 1610 1911 1614
rect 1915 1610 1951 1614
rect 1955 1610 2031 1614
rect 2035 1610 2039 1614
rect 2043 1610 2175 1614
rect 2179 1610 2319 1614
rect 2323 1610 2455 1614
rect 2459 1610 2503 1614
rect 2507 1610 2546 1614
rect 1310 1609 2546 1610
rect 84 1561 85 1567
rect 91 1566 1299 1567
rect 91 1562 111 1566
rect 115 1562 247 1566
rect 251 1562 287 1566
rect 291 1562 319 1566
rect 323 1562 343 1566
rect 347 1562 399 1566
rect 403 1562 415 1566
rect 419 1562 487 1566
rect 491 1562 495 1566
rect 499 1562 583 1566
rect 587 1562 671 1566
rect 675 1562 679 1566
rect 683 1562 759 1566
rect 763 1562 775 1566
rect 779 1562 847 1566
rect 851 1562 879 1566
rect 883 1562 927 1566
rect 931 1562 991 1566
rect 995 1562 1007 1566
rect 1011 1562 1087 1566
rect 1091 1562 1103 1566
rect 1107 1562 1167 1566
rect 1171 1562 1223 1566
rect 1227 1562 1287 1566
rect 1291 1562 1299 1566
rect 91 1561 1299 1562
rect 1305 1563 1306 1567
rect 1305 1562 2534 1563
rect 1305 1561 1327 1562
rect 1298 1558 1327 1561
rect 1331 1558 1351 1562
rect 1355 1558 1407 1562
rect 1411 1558 1463 1562
rect 1467 1558 1471 1562
rect 1475 1558 1543 1562
rect 1547 1558 1607 1562
rect 1611 1558 1623 1562
rect 1627 1558 1703 1562
rect 1707 1558 1735 1562
rect 1739 1558 1775 1562
rect 1779 1558 1855 1562
rect 1859 1558 1871 1562
rect 1875 1558 1935 1562
rect 1939 1558 2007 1562
rect 2011 1558 2015 1562
rect 2019 1558 2503 1562
rect 2507 1558 2534 1562
rect 1298 1557 2534 1558
rect 1310 1510 2546 1511
rect 1310 1507 1327 1510
rect 96 1501 97 1507
rect 103 1506 1311 1507
rect 103 1502 111 1506
rect 115 1502 263 1506
rect 267 1502 279 1506
rect 283 1502 335 1506
rect 339 1502 343 1506
rect 347 1502 415 1506
rect 419 1502 495 1506
rect 499 1502 503 1506
rect 507 1502 575 1506
rect 579 1502 599 1506
rect 603 1502 655 1506
rect 659 1502 687 1506
rect 691 1502 735 1506
rect 739 1502 775 1506
rect 779 1502 815 1506
rect 819 1502 863 1506
rect 867 1502 895 1506
rect 899 1502 943 1506
rect 947 1502 975 1506
rect 979 1502 1023 1506
rect 1027 1502 1055 1506
rect 1059 1502 1103 1506
rect 1107 1502 1143 1506
rect 1147 1502 1183 1506
rect 1187 1502 1239 1506
rect 1243 1502 1287 1506
rect 1291 1502 1311 1506
rect 103 1501 1311 1502
rect 1317 1506 1327 1507
rect 1331 1506 1367 1510
rect 1371 1506 1423 1510
rect 1427 1506 1479 1510
rect 1483 1506 1487 1510
rect 1491 1506 1551 1510
rect 1555 1506 1623 1510
rect 1627 1506 1631 1510
rect 1635 1506 1711 1510
rect 1715 1506 1751 1510
rect 1755 1506 1791 1510
rect 1795 1506 1871 1510
rect 1875 1506 1887 1510
rect 1891 1506 1951 1510
rect 1955 1506 2023 1510
rect 2027 1506 2031 1510
rect 2035 1506 2119 1510
rect 2123 1506 2503 1510
rect 2507 1506 2546 1510
rect 1317 1505 2546 1506
rect 1317 1501 1318 1505
rect 84 1445 85 1451
rect 91 1450 1299 1451
rect 91 1446 111 1450
rect 115 1446 191 1450
rect 195 1446 255 1450
rect 259 1446 263 1450
rect 267 1446 327 1450
rect 331 1446 399 1450
rect 403 1446 407 1450
rect 411 1446 479 1450
rect 483 1446 503 1450
rect 507 1446 559 1450
rect 563 1446 607 1450
rect 611 1446 639 1450
rect 643 1446 711 1450
rect 715 1446 719 1450
rect 723 1446 799 1450
rect 803 1446 815 1450
rect 819 1446 879 1450
rect 883 1446 919 1450
rect 923 1446 959 1450
rect 963 1446 1023 1450
rect 1027 1446 1039 1450
rect 1043 1446 1127 1450
rect 1131 1446 1223 1450
rect 1227 1446 1287 1450
rect 1291 1446 1299 1450
rect 91 1445 1299 1446
rect 1305 1450 2534 1451
rect 1305 1446 1327 1450
rect 1331 1446 1351 1450
rect 1355 1446 1359 1450
rect 1363 1446 1407 1450
rect 1411 1446 1447 1450
rect 1451 1446 1463 1450
rect 1467 1446 1535 1450
rect 1539 1446 1615 1450
rect 1619 1446 1631 1450
rect 1635 1446 1695 1450
rect 1699 1446 1727 1450
rect 1731 1446 1775 1450
rect 1779 1446 1815 1450
rect 1819 1446 1855 1450
rect 1859 1446 1903 1450
rect 1907 1446 1935 1450
rect 1939 1446 1991 1450
rect 1995 1446 2015 1450
rect 2019 1446 2071 1450
rect 2075 1446 2103 1450
rect 2107 1446 2159 1450
rect 2163 1446 2247 1450
rect 2251 1446 2503 1450
rect 2507 1446 2534 1450
rect 1305 1445 2534 1446
rect 1310 1398 2546 1399
rect 1310 1395 1327 1398
rect 96 1389 97 1395
rect 103 1394 1311 1395
rect 103 1390 111 1394
rect 115 1390 151 1394
rect 155 1390 207 1394
rect 211 1390 223 1394
rect 227 1390 271 1394
rect 275 1390 295 1394
rect 299 1390 343 1394
rect 347 1390 359 1394
rect 363 1390 423 1394
rect 427 1390 431 1394
rect 435 1390 503 1394
rect 507 1390 519 1394
rect 523 1390 583 1394
rect 587 1390 623 1394
rect 627 1390 663 1394
rect 667 1390 727 1394
rect 731 1390 751 1394
rect 755 1390 831 1394
rect 835 1390 839 1394
rect 843 1390 927 1394
rect 931 1390 935 1394
rect 939 1390 1015 1394
rect 1019 1390 1039 1394
rect 1043 1390 1103 1394
rect 1107 1390 1143 1394
rect 1147 1390 1199 1394
rect 1203 1390 1239 1394
rect 1243 1390 1287 1394
rect 1291 1390 1311 1394
rect 103 1389 1311 1390
rect 1317 1394 1327 1395
rect 1331 1394 1375 1398
rect 1379 1394 1463 1398
rect 1467 1394 1551 1398
rect 1555 1394 1567 1398
rect 1571 1394 1647 1398
rect 1651 1394 1735 1398
rect 1739 1394 1743 1398
rect 1747 1394 1831 1398
rect 1835 1394 1919 1398
rect 1923 1394 2007 1398
rect 2011 1394 2087 1398
rect 2091 1394 2095 1398
rect 2099 1394 2175 1398
rect 2179 1394 2247 1398
rect 2251 1394 2263 1398
rect 2267 1394 2319 1398
rect 2323 1394 2399 1398
rect 2403 1394 2455 1398
rect 2459 1394 2503 1398
rect 2507 1394 2546 1398
rect 1317 1393 2546 1394
rect 1317 1389 1318 1393
rect 1298 1341 1299 1347
rect 1305 1346 2527 1347
rect 1305 1342 1327 1346
rect 1331 1342 1551 1346
rect 1555 1342 1583 1346
rect 1587 1342 1631 1346
rect 1635 1342 1647 1346
rect 1651 1342 1719 1346
rect 1723 1342 1727 1346
rect 1731 1342 1807 1346
rect 1811 1342 1815 1346
rect 1819 1342 1895 1346
rect 1899 1342 1903 1346
rect 1907 1342 1983 1346
rect 1987 1342 1991 1346
rect 1995 1342 2063 1346
rect 2067 1342 2079 1346
rect 2083 1342 2143 1346
rect 2147 1342 2159 1346
rect 2163 1342 2223 1346
rect 2227 1342 2231 1346
rect 2235 1342 2303 1346
rect 2307 1342 2383 1346
rect 2387 1342 2439 1346
rect 2443 1342 2503 1346
rect 2507 1342 2527 1346
rect 1305 1341 2527 1342
rect 2533 1341 2534 1347
rect 84 1321 85 1327
rect 91 1326 1299 1327
rect 91 1322 111 1326
rect 115 1322 135 1326
rect 139 1322 207 1326
rect 211 1322 239 1326
rect 243 1322 279 1326
rect 283 1322 343 1326
rect 347 1322 367 1326
rect 371 1322 415 1326
rect 419 1322 479 1326
rect 483 1322 487 1326
rect 491 1322 567 1326
rect 571 1322 583 1326
rect 587 1322 647 1326
rect 651 1322 687 1326
rect 691 1322 735 1326
rect 739 1322 783 1326
rect 787 1322 823 1326
rect 827 1322 879 1326
rect 883 1322 911 1326
rect 915 1322 975 1326
rect 979 1322 999 1326
rect 1003 1322 1087 1326
rect 1091 1322 1183 1326
rect 1187 1322 1287 1326
rect 1291 1322 1299 1326
rect 91 1321 1299 1322
rect 1305 1321 1306 1327
rect 1310 1289 1311 1295
rect 1317 1294 2539 1295
rect 1317 1290 1327 1294
rect 1331 1290 1567 1294
rect 1571 1290 1599 1294
rect 1603 1290 1631 1294
rect 1635 1290 1663 1294
rect 1667 1290 1711 1294
rect 1715 1290 1743 1294
rect 1747 1290 1799 1294
rect 1803 1290 1823 1294
rect 1827 1290 1895 1294
rect 1899 1290 1911 1294
rect 1915 1290 1991 1294
rect 1995 1290 1999 1294
rect 2003 1290 2079 1294
rect 2083 1290 2095 1294
rect 2099 1290 2159 1294
rect 2163 1290 2207 1294
rect 2211 1290 2239 1294
rect 2243 1290 2319 1294
rect 2323 1290 2399 1294
rect 2403 1290 2455 1294
rect 2459 1290 2503 1294
rect 2507 1290 2539 1294
rect 1317 1289 2539 1290
rect 2545 1289 2546 1295
rect 96 1261 97 1267
rect 103 1266 1311 1267
rect 103 1262 111 1266
rect 115 1262 151 1266
rect 155 1262 215 1266
rect 219 1262 255 1266
rect 259 1262 303 1266
rect 307 1262 383 1266
rect 387 1262 391 1266
rect 395 1262 471 1266
rect 475 1262 495 1266
rect 499 1262 551 1266
rect 555 1262 599 1266
rect 603 1262 623 1266
rect 627 1262 695 1266
rect 699 1262 703 1266
rect 707 1262 767 1266
rect 771 1262 799 1266
rect 803 1262 839 1266
rect 843 1262 895 1266
rect 899 1262 919 1266
rect 923 1262 991 1266
rect 995 1262 1287 1266
rect 1291 1262 1311 1266
rect 103 1261 1311 1262
rect 1317 1261 1318 1267
rect 1298 1233 1299 1239
rect 1305 1238 2527 1239
rect 1305 1234 1327 1238
rect 1331 1234 1519 1238
rect 1523 1234 1551 1238
rect 1555 1234 1575 1238
rect 1579 1234 1615 1238
rect 1619 1234 1631 1238
rect 1635 1234 1687 1238
rect 1691 1234 1695 1238
rect 1699 1234 1743 1238
rect 1747 1234 1783 1238
rect 1787 1234 1799 1238
rect 1803 1234 1855 1238
rect 1859 1234 1879 1238
rect 1883 1234 1911 1238
rect 1915 1234 1967 1238
rect 1971 1234 1975 1238
rect 1979 1234 2031 1238
rect 2035 1234 2079 1238
rect 2083 1234 2103 1238
rect 2107 1234 2183 1238
rect 2187 1234 2191 1238
rect 2195 1234 2271 1238
rect 2275 1234 2303 1238
rect 2307 1234 2367 1238
rect 2371 1234 2439 1238
rect 2443 1234 2503 1238
rect 2507 1234 2527 1238
rect 1305 1233 2527 1234
rect 2533 1233 2534 1239
rect 84 1205 85 1211
rect 91 1210 1299 1211
rect 91 1206 111 1210
rect 115 1206 135 1210
rect 139 1206 191 1210
rect 195 1206 199 1210
rect 203 1206 271 1210
rect 275 1206 287 1210
rect 291 1206 351 1210
rect 355 1206 375 1210
rect 379 1206 431 1210
rect 435 1206 455 1210
rect 459 1206 511 1210
rect 515 1206 535 1210
rect 539 1206 583 1210
rect 587 1206 607 1210
rect 611 1206 647 1210
rect 651 1206 679 1210
rect 683 1206 719 1210
rect 723 1206 751 1210
rect 755 1206 791 1210
rect 795 1206 823 1210
rect 827 1206 863 1210
rect 867 1206 903 1210
rect 907 1206 1287 1210
rect 1291 1206 1299 1210
rect 91 1205 1299 1206
rect 1305 1205 1306 1211
rect 1310 1177 1311 1183
rect 1317 1182 2539 1183
rect 1317 1178 1327 1182
rect 1331 1178 1535 1182
rect 1539 1178 1567 1182
rect 1571 1178 1591 1182
rect 1595 1178 1631 1182
rect 1635 1178 1647 1182
rect 1651 1178 1703 1182
rect 1707 1178 1759 1182
rect 1763 1178 1791 1182
rect 1795 1178 1815 1182
rect 1819 1178 1871 1182
rect 1875 1178 1903 1182
rect 1907 1178 1927 1182
rect 1931 1178 1983 1182
rect 1987 1178 2031 1182
rect 2035 1178 2047 1182
rect 2051 1178 2119 1182
rect 2123 1178 2175 1182
rect 2179 1178 2199 1182
rect 2203 1178 2287 1182
rect 2291 1178 2327 1182
rect 2331 1178 2383 1182
rect 2387 1178 2455 1182
rect 2459 1178 2503 1182
rect 2507 1178 2539 1182
rect 1317 1177 2539 1178
rect 2545 1177 2546 1183
rect 96 1149 97 1155
rect 103 1154 1311 1155
rect 103 1150 111 1154
rect 115 1150 151 1154
rect 155 1150 183 1154
rect 187 1150 207 1154
rect 211 1150 279 1154
rect 283 1150 287 1154
rect 291 1150 367 1154
rect 371 1150 375 1154
rect 379 1150 447 1154
rect 451 1150 471 1154
rect 475 1150 527 1154
rect 531 1150 567 1154
rect 571 1150 599 1154
rect 603 1150 655 1154
rect 659 1150 663 1154
rect 667 1150 735 1154
rect 739 1150 807 1154
rect 811 1150 879 1154
rect 883 1150 959 1154
rect 963 1150 1039 1154
rect 1043 1150 1287 1154
rect 1291 1150 1311 1154
rect 103 1149 1311 1150
rect 1317 1149 1318 1155
rect 1298 1125 1299 1131
rect 1305 1130 2527 1131
rect 1305 1126 1327 1130
rect 1331 1126 1383 1130
rect 1387 1126 1447 1130
rect 1451 1126 1519 1130
rect 1523 1126 1551 1130
rect 1555 1126 1591 1130
rect 1595 1126 1615 1130
rect 1619 1126 1671 1130
rect 1675 1126 1687 1130
rect 1691 1126 1751 1130
rect 1755 1126 1775 1130
rect 1779 1126 1831 1130
rect 1835 1126 1887 1130
rect 1891 1126 1911 1130
rect 1915 1126 1983 1130
rect 1987 1126 2015 1130
rect 2019 1126 2055 1130
rect 2059 1126 2135 1130
rect 2139 1126 2159 1130
rect 2163 1126 2215 1130
rect 2219 1126 2311 1130
rect 2315 1126 2439 1130
rect 2443 1126 2503 1130
rect 2507 1126 2527 1130
rect 1305 1125 2527 1126
rect 2533 1125 2534 1131
rect 84 1089 85 1095
rect 91 1094 1299 1095
rect 91 1090 111 1094
rect 115 1090 167 1094
rect 171 1090 207 1094
rect 211 1090 263 1094
rect 267 1090 279 1094
rect 283 1090 359 1094
rect 363 1090 447 1094
rect 451 1090 455 1094
rect 459 1090 543 1094
rect 547 1090 551 1094
rect 555 1090 639 1094
rect 643 1090 719 1094
rect 723 1090 727 1094
rect 731 1090 791 1094
rect 795 1090 815 1094
rect 819 1090 863 1094
rect 867 1090 895 1094
rect 899 1090 943 1094
rect 947 1090 975 1094
rect 979 1090 1023 1094
rect 1027 1090 1055 1094
rect 1059 1090 1143 1094
rect 1147 1090 1287 1094
rect 1291 1090 1299 1094
rect 91 1089 1299 1090
rect 1305 1089 1306 1095
rect 1310 1065 1311 1071
rect 1317 1070 2539 1071
rect 1317 1066 1327 1070
rect 1331 1066 1367 1070
rect 1371 1066 1399 1070
rect 1403 1066 1455 1070
rect 1459 1066 1463 1070
rect 1467 1066 1535 1070
rect 1539 1066 1575 1070
rect 1579 1066 1607 1070
rect 1611 1066 1687 1070
rect 1691 1066 1695 1070
rect 1699 1066 1767 1070
rect 1771 1066 1815 1070
rect 1819 1066 1847 1070
rect 1851 1066 1927 1070
rect 1931 1066 1999 1070
rect 2003 1066 2039 1070
rect 2043 1066 2071 1070
rect 2075 1066 2151 1070
rect 2155 1066 2231 1070
rect 2235 1066 2255 1070
rect 2259 1066 2367 1070
rect 2371 1066 2455 1070
rect 2459 1066 2503 1070
rect 2507 1066 2539 1070
rect 1317 1065 2539 1066
rect 2545 1065 2546 1071
rect 96 1029 97 1035
rect 103 1034 1311 1035
rect 103 1030 111 1034
rect 115 1030 223 1034
rect 227 1030 295 1034
rect 299 1030 375 1034
rect 379 1030 383 1034
rect 387 1030 463 1034
rect 467 1030 479 1034
rect 483 1030 559 1034
rect 563 1030 575 1034
rect 579 1030 655 1034
rect 659 1030 671 1034
rect 675 1030 743 1034
rect 747 1030 767 1034
rect 771 1030 831 1034
rect 835 1030 855 1034
rect 859 1030 911 1034
rect 915 1030 943 1034
rect 947 1030 991 1034
rect 995 1030 1023 1034
rect 1027 1030 1071 1034
rect 1075 1030 1103 1034
rect 1107 1030 1159 1034
rect 1163 1030 1183 1034
rect 1187 1030 1239 1034
rect 1243 1030 1287 1034
rect 1291 1030 1311 1034
rect 103 1029 1311 1030
rect 1317 1029 1318 1035
rect 1298 1009 1299 1015
rect 1305 1014 2527 1015
rect 1305 1010 1327 1014
rect 1331 1010 1351 1014
rect 1355 1010 1439 1014
rect 1443 1010 1511 1014
rect 1515 1010 1559 1014
rect 1563 1010 1679 1014
rect 1683 1010 1799 1014
rect 1803 1010 1823 1014
rect 1827 1010 1911 1014
rect 1915 1010 1951 1014
rect 1955 1010 2023 1014
rect 2027 1010 2071 1014
rect 2075 1010 2135 1014
rect 2139 1010 2175 1014
rect 2179 1010 2239 1014
rect 2243 1010 2271 1014
rect 2275 1010 2351 1014
rect 2355 1010 2367 1014
rect 2371 1010 2439 1014
rect 2443 1010 2503 1014
rect 2507 1010 2527 1014
rect 1305 1009 2527 1010
rect 2533 1009 2534 1015
rect 84 977 85 983
rect 91 982 1299 983
rect 91 978 111 982
rect 115 978 271 982
rect 275 978 279 982
rect 283 978 359 982
rect 363 978 367 982
rect 371 978 455 982
rect 459 978 463 982
rect 467 978 551 982
rect 555 978 559 982
rect 563 978 655 982
rect 659 978 751 982
rect 755 978 839 982
rect 843 978 927 982
rect 931 978 1007 982
rect 1011 978 1087 982
rect 1091 978 1167 982
rect 1171 978 1223 982
rect 1227 978 1287 982
rect 1291 978 1299 982
rect 91 977 1299 978
rect 1305 977 1306 983
rect 1310 945 1311 951
rect 1317 950 2539 951
rect 1317 946 1327 950
rect 1331 946 1367 950
rect 1371 946 1423 950
rect 1427 946 1503 950
rect 1507 946 1527 950
rect 1531 946 1607 950
rect 1611 946 1695 950
rect 1699 946 1719 950
rect 1723 946 1831 950
rect 1835 946 1839 950
rect 1843 946 1935 950
rect 1939 946 1967 950
rect 1971 946 2031 950
rect 2035 946 2087 950
rect 2091 946 2127 950
rect 2131 946 2191 950
rect 2195 946 2215 950
rect 2219 946 2287 950
rect 2291 946 2295 950
rect 2299 946 2375 950
rect 2379 946 2383 950
rect 2387 946 2455 950
rect 2459 946 2503 950
rect 2507 946 2539 950
rect 1317 945 2539 946
rect 2545 945 2546 951
rect 96 917 97 923
rect 103 922 1311 923
rect 103 918 111 922
rect 115 918 271 922
rect 275 918 287 922
rect 291 918 343 922
rect 347 918 375 922
rect 379 918 423 922
rect 427 918 471 922
rect 475 918 519 922
rect 523 918 567 922
rect 571 918 615 922
rect 619 918 671 922
rect 675 918 711 922
rect 715 918 767 922
rect 771 918 807 922
rect 811 918 855 922
rect 859 918 903 922
rect 907 918 943 922
rect 947 918 991 922
rect 995 918 1023 922
rect 1027 918 1087 922
rect 1091 918 1103 922
rect 1107 918 1183 922
rect 1187 918 1239 922
rect 1243 918 1287 922
rect 1291 918 1311 922
rect 103 917 1311 918
rect 1317 917 1318 923
rect 1298 889 1299 895
rect 1305 894 2527 895
rect 1305 890 1327 894
rect 1331 890 1351 894
rect 1355 890 1407 894
rect 1411 890 1431 894
rect 1435 890 1487 894
rect 1491 890 1551 894
rect 1555 890 1591 894
rect 1595 890 1623 894
rect 1627 890 1703 894
rect 1707 890 1791 894
rect 1795 890 1815 894
rect 1819 890 1895 894
rect 1899 890 1919 894
rect 1923 890 2015 894
rect 2019 890 2111 894
rect 2115 890 2143 894
rect 2147 890 2199 894
rect 2203 890 2279 894
rect 2283 890 2359 894
rect 2363 890 2423 894
rect 2427 890 2439 894
rect 2443 890 2503 894
rect 2507 890 2527 894
rect 1305 889 2527 890
rect 2533 889 2534 895
rect 84 861 85 867
rect 91 866 1299 867
rect 91 862 111 866
rect 115 862 247 866
rect 251 862 255 866
rect 259 862 311 866
rect 315 862 327 866
rect 331 862 375 866
rect 379 862 407 866
rect 411 862 439 866
rect 443 862 503 866
rect 507 862 567 866
rect 571 862 599 866
rect 603 862 631 866
rect 635 862 695 866
rect 699 862 759 866
rect 763 862 791 866
rect 795 862 831 866
rect 835 862 887 866
rect 891 862 903 866
rect 907 862 975 866
rect 979 862 1071 866
rect 1075 862 1167 866
rect 1171 862 1287 866
rect 1291 862 1299 866
rect 91 861 1299 862
rect 1305 861 1306 867
rect 1310 833 1311 839
rect 1317 838 2539 839
rect 1317 834 1327 838
rect 1331 834 1447 838
rect 1451 834 1503 838
rect 1507 834 1567 838
rect 1571 834 1591 838
rect 1595 834 1639 838
rect 1643 834 1647 838
rect 1651 834 1703 838
rect 1707 834 1719 838
rect 1723 834 1767 838
rect 1771 834 1807 838
rect 1811 834 1847 838
rect 1851 834 1911 838
rect 1915 834 1927 838
rect 1931 834 2015 838
rect 2019 834 2031 838
rect 2035 834 2103 838
rect 2107 834 2159 838
rect 2163 834 2191 838
rect 2195 834 2287 838
rect 2291 834 2295 838
rect 2299 834 2383 838
rect 2387 834 2439 838
rect 2443 834 2455 838
rect 2459 834 2503 838
rect 2507 834 2539 838
rect 1317 833 2539 834
rect 2545 833 2546 839
rect 96 805 97 811
rect 103 810 1311 811
rect 103 806 111 810
rect 115 806 215 810
rect 219 806 263 810
rect 267 806 303 810
rect 307 806 327 810
rect 331 806 391 810
rect 395 806 455 810
rect 459 806 479 810
rect 483 806 519 810
rect 523 806 559 810
rect 563 806 583 810
rect 587 806 631 810
rect 635 806 647 810
rect 651 806 703 810
rect 707 806 711 810
rect 715 806 767 810
rect 771 806 775 810
rect 779 806 831 810
rect 835 806 847 810
rect 851 806 895 810
rect 899 806 919 810
rect 923 806 967 810
rect 971 806 1039 810
rect 1043 806 1287 810
rect 1291 806 1311 810
rect 103 805 1311 806
rect 1317 805 1318 811
rect 1298 777 1299 783
rect 1305 782 2527 783
rect 1305 778 1327 782
rect 1331 778 1567 782
rect 1571 778 1575 782
rect 1579 778 1623 782
rect 1627 778 1631 782
rect 1635 778 1687 782
rect 1691 778 1751 782
rect 1755 778 1759 782
rect 1763 778 1831 782
rect 1835 778 1911 782
rect 1915 778 1919 782
rect 1923 778 1999 782
rect 2003 778 2015 782
rect 2019 778 2087 782
rect 2091 778 2119 782
rect 2123 778 2175 782
rect 2179 778 2231 782
rect 2235 778 2271 782
rect 2275 778 2343 782
rect 2347 778 2367 782
rect 2371 778 2439 782
rect 2443 778 2503 782
rect 2507 778 2527 782
rect 1305 777 2527 778
rect 2533 777 2534 783
rect 84 753 85 759
rect 91 758 1299 759
rect 91 754 111 758
rect 115 754 135 758
rect 139 754 199 758
rect 203 754 255 758
rect 259 754 287 758
rect 291 754 375 758
rect 379 754 391 758
rect 395 754 463 758
rect 467 754 519 758
rect 523 754 543 758
rect 547 754 615 758
rect 619 754 647 758
rect 651 754 687 758
rect 691 754 751 758
rect 755 754 775 758
rect 779 754 815 758
rect 819 754 879 758
rect 883 754 903 758
rect 907 754 951 758
rect 955 754 1023 758
rect 1027 754 1039 758
rect 1043 754 1287 758
rect 1291 754 1299 758
rect 91 753 1299 754
rect 1305 753 1306 759
rect 1310 725 1311 731
rect 1317 730 2539 731
rect 1317 726 1327 730
rect 1331 726 1367 730
rect 1371 726 1431 730
rect 1435 726 1527 730
rect 1531 726 1583 730
rect 1587 726 1631 730
rect 1635 726 1639 730
rect 1643 726 1703 730
rect 1707 726 1735 730
rect 1739 726 1775 730
rect 1779 726 1839 730
rect 1843 726 1847 730
rect 1851 726 1935 730
rect 1939 726 1943 730
rect 1947 726 2031 730
rect 2035 726 2047 730
rect 2051 726 2135 730
rect 2139 726 2151 730
rect 2155 726 2247 730
rect 2251 726 2255 730
rect 2259 726 2359 730
rect 2363 726 2367 730
rect 2371 726 2455 730
rect 2459 726 2503 730
rect 2507 726 2539 730
rect 1317 725 2539 726
rect 2545 725 2546 731
rect 96 701 97 707
rect 103 706 1311 707
rect 103 702 111 706
rect 115 702 151 706
rect 155 702 207 706
rect 211 702 271 706
rect 275 702 295 706
rect 299 702 391 706
rect 395 702 407 706
rect 411 702 503 706
rect 507 702 535 706
rect 539 702 623 706
rect 627 702 663 706
rect 667 702 743 706
rect 747 702 791 706
rect 795 702 871 706
rect 875 702 919 706
rect 923 702 999 706
rect 1003 702 1055 706
rect 1059 702 1127 706
rect 1131 702 1239 706
rect 1243 702 1287 706
rect 1291 702 1311 706
rect 103 701 1311 702
rect 1317 701 1318 707
rect 1298 661 1299 667
rect 1305 666 2527 667
rect 1305 662 1327 666
rect 1331 662 1351 666
rect 1355 662 1415 666
rect 1419 662 1511 666
rect 1515 662 1607 666
rect 1611 662 1615 666
rect 1619 662 1711 666
rect 1715 662 1719 666
rect 1723 662 1823 666
rect 1827 662 1927 666
rect 1931 662 1935 666
rect 1939 662 2031 666
rect 2035 662 2055 666
rect 2059 662 2135 666
rect 2139 662 2183 666
rect 2187 662 2239 666
rect 2243 662 2319 666
rect 2323 662 2351 666
rect 2355 662 2439 666
rect 2443 662 2503 666
rect 2507 662 2527 666
rect 1305 661 2527 662
rect 2533 661 2534 667
rect 84 645 85 651
rect 91 650 1299 651
rect 91 646 111 650
rect 115 646 135 650
rect 139 646 151 650
rect 155 646 191 650
rect 195 646 263 650
rect 267 646 279 650
rect 283 646 367 650
rect 371 646 375 650
rect 379 646 463 650
rect 467 646 487 650
rect 491 646 559 650
rect 563 646 607 650
rect 611 646 655 650
rect 659 646 727 650
rect 731 646 751 650
rect 755 646 847 650
rect 851 646 855 650
rect 859 646 943 650
rect 947 646 983 650
rect 987 646 1039 650
rect 1043 646 1111 650
rect 1115 646 1143 650
rect 1147 646 1223 650
rect 1227 646 1287 650
rect 1291 646 1299 650
rect 91 645 1299 646
rect 1305 645 1306 651
rect 1310 609 1311 615
rect 1317 614 2539 615
rect 1317 610 1327 614
rect 1331 610 1367 614
rect 1371 610 1383 614
rect 1387 610 1431 614
rect 1435 610 1463 614
rect 1467 610 1527 614
rect 1531 610 1551 614
rect 1555 610 1623 614
rect 1627 610 1647 614
rect 1651 610 1727 614
rect 1731 610 1743 614
rect 1747 610 1839 614
rect 1843 610 1847 614
rect 1851 610 1951 614
rect 1955 610 1959 614
rect 1963 610 2071 614
rect 2075 610 2079 614
rect 2083 610 2199 614
rect 2203 610 2207 614
rect 2211 610 2335 614
rect 2339 610 2343 614
rect 2347 610 2455 614
rect 2459 610 2503 614
rect 2507 610 2539 614
rect 1317 609 2539 610
rect 2545 609 2546 615
rect 96 593 97 599
rect 103 598 1311 599
rect 103 594 111 598
rect 115 594 151 598
rect 155 594 167 598
rect 171 594 239 598
rect 243 594 279 598
rect 283 594 335 598
rect 339 594 383 598
rect 387 594 431 598
rect 435 594 479 598
rect 483 594 535 598
rect 539 594 575 598
rect 579 594 631 598
rect 635 594 671 598
rect 675 594 727 598
rect 731 594 767 598
rect 771 594 823 598
rect 827 594 863 598
rect 867 594 911 598
rect 915 594 959 598
rect 963 594 999 598
rect 1003 594 1055 598
rect 1059 594 1087 598
rect 1091 594 1159 598
rect 1163 594 1183 598
rect 1187 594 1239 598
rect 1243 594 1287 598
rect 1291 594 1311 598
rect 103 593 1311 594
rect 1317 593 1318 599
rect 1298 557 1299 563
rect 1305 562 2527 563
rect 1305 558 1327 562
rect 1331 558 1367 562
rect 1371 558 1375 562
rect 1379 558 1447 562
rect 1451 558 1455 562
rect 1459 558 1535 562
rect 1539 558 1551 562
rect 1555 558 1631 562
rect 1635 558 1647 562
rect 1651 558 1727 562
rect 1731 558 1751 562
rect 1755 558 1831 562
rect 1835 558 1855 562
rect 1859 558 1943 562
rect 1947 558 1959 562
rect 1963 558 2055 562
rect 2059 558 2063 562
rect 2067 558 2151 562
rect 2155 558 2191 562
rect 2195 558 2255 562
rect 2259 558 2327 562
rect 2331 558 2359 562
rect 2363 558 2439 562
rect 2443 558 2503 562
rect 2507 558 2527 562
rect 1305 557 2527 558
rect 2533 557 2534 563
rect 84 533 85 539
rect 91 538 1299 539
rect 91 534 111 538
rect 115 534 135 538
rect 139 534 143 538
rect 147 534 223 538
rect 227 534 239 538
rect 243 534 319 538
rect 323 534 335 538
rect 339 534 415 538
rect 419 534 431 538
rect 435 534 519 538
rect 523 534 527 538
rect 531 534 615 538
rect 619 534 623 538
rect 627 534 711 538
rect 715 534 791 538
rect 795 534 807 538
rect 811 534 871 538
rect 875 534 895 538
rect 899 534 951 538
rect 955 534 983 538
rect 987 534 1031 538
rect 1035 534 1071 538
rect 1075 534 1167 538
rect 1171 534 1287 538
rect 1291 534 1299 538
rect 91 533 1299 534
rect 1305 533 1306 539
rect 1310 501 1311 507
rect 1317 506 2539 507
rect 1317 502 1327 506
rect 1331 502 1367 506
rect 1371 502 1391 506
rect 1395 502 1455 506
rect 1459 502 1471 506
rect 1475 502 1567 506
rect 1571 502 1575 506
rect 1579 502 1663 506
rect 1667 502 1695 506
rect 1699 502 1767 506
rect 1771 502 1807 506
rect 1811 502 1871 506
rect 1875 502 1919 506
rect 1923 502 1975 506
rect 1979 502 2023 506
rect 2027 502 2071 506
rect 2075 502 2119 506
rect 2123 502 2167 506
rect 2171 502 2207 506
rect 2211 502 2271 506
rect 2275 502 2295 506
rect 2299 502 2375 506
rect 2379 502 2383 506
rect 2387 502 2455 506
rect 2459 502 2503 506
rect 2507 502 2539 506
rect 1317 501 2539 502
rect 2545 501 2546 507
rect 96 477 97 483
rect 103 482 1311 483
rect 103 478 111 482
rect 115 478 151 482
rect 155 478 159 482
rect 163 478 207 482
rect 211 478 255 482
rect 259 478 287 482
rect 291 478 351 482
rect 355 478 375 482
rect 379 478 447 482
rect 451 478 463 482
rect 467 478 543 482
rect 547 478 559 482
rect 563 478 639 482
rect 643 478 655 482
rect 659 478 727 482
rect 731 478 751 482
rect 755 478 807 482
rect 811 478 847 482
rect 851 478 887 482
rect 891 478 951 482
rect 955 478 967 482
rect 971 478 1047 482
rect 1051 478 1055 482
rect 1059 478 1159 482
rect 1163 478 1239 482
rect 1243 478 1287 482
rect 1291 478 1311 482
rect 103 477 1311 478
rect 1317 477 1318 483
rect 1298 437 1299 443
rect 1305 442 2527 443
rect 1305 438 1327 442
rect 1331 438 1351 442
rect 1355 438 1439 442
rect 1443 438 1559 442
rect 1563 438 1583 442
rect 1587 438 1639 442
rect 1643 438 1679 442
rect 1683 438 1695 442
rect 1699 438 1759 442
rect 1763 438 1791 442
rect 1795 438 1831 442
rect 1835 438 1903 442
rect 1907 438 1911 442
rect 1915 438 1991 442
rect 1995 438 2007 442
rect 2011 438 2079 442
rect 2083 438 2103 442
rect 2107 438 2175 442
rect 2179 438 2191 442
rect 2195 438 2271 442
rect 2275 438 2279 442
rect 2283 438 2367 442
rect 2371 438 2439 442
rect 2443 438 2503 442
rect 2507 438 2527 442
rect 1305 437 2527 438
rect 2533 437 2534 443
rect 84 425 85 431
rect 91 430 1299 431
rect 91 426 111 430
rect 115 426 135 430
rect 139 426 191 430
rect 195 426 271 430
rect 275 426 279 430
rect 283 426 359 430
rect 363 426 383 430
rect 387 426 447 430
rect 451 426 495 430
rect 499 426 543 430
rect 547 426 607 430
rect 611 426 639 430
rect 643 426 719 430
rect 723 426 735 430
rect 739 426 831 430
rect 835 426 935 430
rect 939 426 1039 430
rect 1043 426 1143 430
rect 1147 426 1223 430
rect 1227 426 1287 430
rect 1291 426 1299 430
rect 91 425 1299 426
rect 1305 425 1306 431
rect 1310 381 1311 387
rect 1317 386 2539 387
rect 1317 382 1327 386
rect 1331 382 1599 386
rect 1603 382 1655 386
rect 1659 382 1679 386
rect 1683 382 1711 386
rect 1715 382 1735 386
rect 1739 382 1775 386
rect 1779 382 1799 386
rect 1803 382 1847 386
rect 1851 382 1871 386
rect 1875 382 1927 386
rect 1931 382 1943 386
rect 1947 382 2007 386
rect 2011 382 2023 386
rect 2027 382 2095 386
rect 2099 382 2111 386
rect 2115 382 2191 386
rect 2195 382 2199 386
rect 2203 382 2287 386
rect 2291 382 2375 386
rect 2379 382 2383 386
rect 2387 382 2455 386
rect 2459 382 2503 386
rect 2507 382 2539 386
rect 1317 381 2539 382
rect 2545 381 2546 387
rect 96 369 97 375
rect 103 374 1311 375
rect 103 370 111 374
rect 115 370 151 374
rect 155 370 207 374
rect 211 370 231 374
rect 235 370 295 374
rect 299 370 335 374
rect 339 370 399 374
rect 403 370 439 374
rect 443 370 511 374
rect 515 370 543 374
rect 547 370 623 374
rect 627 370 647 374
rect 651 370 735 374
rect 739 370 751 374
rect 755 370 847 374
rect 851 370 935 374
rect 939 370 951 374
rect 955 370 1015 374
rect 1019 370 1055 374
rect 1059 370 1095 374
rect 1099 370 1159 374
rect 1163 370 1175 374
rect 1179 370 1239 374
rect 1243 370 1287 374
rect 1291 370 1311 374
rect 103 369 1311 370
rect 1317 369 1318 375
rect 1298 321 1299 327
rect 1305 326 2527 327
rect 1305 322 1327 326
rect 1331 322 1351 326
rect 1355 322 1455 326
rect 1459 322 1583 326
rect 1587 322 1663 326
rect 1667 322 1711 326
rect 1715 322 1719 326
rect 1723 322 1783 326
rect 1787 322 1839 326
rect 1843 322 1855 326
rect 1859 322 1927 326
rect 1931 322 1951 326
rect 1955 322 2007 326
rect 2011 322 2063 326
rect 2067 322 2095 326
rect 2099 322 2167 326
rect 2171 322 2183 326
rect 2187 322 2263 326
rect 2267 322 2271 326
rect 2275 322 2359 326
rect 2363 322 2439 326
rect 2443 322 2503 326
rect 2507 322 2527 326
rect 1305 321 2527 322
rect 2533 321 2534 327
rect 1298 319 1306 321
rect 84 313 85 319
rect 91 318 1299 319
rect 91 314 111 318
rect 115 314 135 318
rect 139 314 215 318
rect 219 314 319 318
rect 323 314 423 318
rect 427 314 527 318
rect 531 314 535 318
rect 539 314 631 318
rect 635 314 639 318
rect 643 314 735 318
rect 739 314 743 318
rect 747 314 831 318
rect 835 314 847 318
rect 851 314 919 318
rect 923 314 943 318
rect 947 314 999 318
rect 1003 314 1039 318
rect 1043 314 1079 318
rect 1083 314 1143 318
rect 1147 314 1159 318
rect 1163 314 1223 318
rect 1227 314 1287 318
rect 1291 314 1299 318
rect 91 313 1299 314
rect 1305 313 1306 319
rect 96 261 97 267
rect 103 266 1311 267
rect 103 262 111 266
rect 115 262 151 266
rect 155 262 223 266
rect 227 262 231 266
rect 235 262 319 266
rect 323 262 335 266
rect 339 262 423 266
rect 427 262 439 266
rect 443 262 535 266
rect 539 262 551 266
rect 555 262 647 266
rect 651 262 655 266
rect 659 262 759 266
rect 763 262 863 266
rect 867 262 871 266
rect 875 262 959 266
rect 963 262 983 266
rect 987 262 1055 266
rect 1059 262 1103 266
rect 1107 262 1159 266
rect 1163 262 1223 266
rect 1227 262 1239 266
rect 1243 262 1287 266
rect 1291 262 1311 266
rect 103 261 1311 262
rect 1317 266 2546 267
rect 1317 262 1327 266
rect 1331 262 1367 266
rect 1371 262 1447 266
rect 1451 262 1471 266
rect 1475 262 1551 266
rect 1555 262 1599 266
rect 1603 262 1655 266
rect 1659 262 1727 266
rect 1731 262 1759 266
rect 1763 262 1855 266
rect 1859 262 1863 266
rect 1867 262 1967 266
rect 1971 262 2071 266
rect 2075 262 2079 266
rect 2083 262 2175 266
rect 2179 262 2183 266
rect 2187 262 2271 266
rect 2275 262 2279 266
rect 2283 262 2375 266
rect 2379 262 2455 266
rect 2459 262 2503 266
rect 2507 262 2546 266
rect 1317 261 2546 262
rect 84 205 85 211
rect 91 210 1299 211
rect 91 206 111 210
rect 115 206 135 210
rect 139 206 183 210
rect 187 206 207 210
rect 211 206 279 210
rect 283 206 303 210
rect 307 206 383 210
rect 387 206 407 210
rect 411 206 487 210
rect 491 206 519 210
rect 523 206 591 210
rect 595 206 631 210
rect 635 206 695 210
rect 699 206 743 210
rect 747 206 799 210
rect 803 206 855 210
rect 859 206 895 210
rect 899 206 967 210
rect 971 206 999 210
rect 1003 206 1087 210
rect 1091 206 1103 210
rect 1107 206 1207 210
rect 1211 206 1287 210
rect 1291 206 1299 210
rect 91 205 1299 206
rect 1305 210 2534 211
rect 1305 206 1327 210
rect 1331 206 1351 210
rect 1355 206 1407 210
rect 1411 206 1431 210
rect 1435 206 1471 210
rect 1475 206 1535 210
rect 1539 206 1551 210
rect 1555 206 1639 210
rect 1643 206 1719 210
rect 1723 206 1743 210
rect 1747 206 1807 210
rect 1811 206 1847 210
rect 1851 206 1895 210
rect 1899 206 1951 210
rect 1955 206 1991 210
rect 1995 206 2055 210
rect 2059 206 2103 210
rect 2107 206 2159 210
rect 2163 206 2215 210
rect 2219 206 2255 210
rect 2259 206 2335 210
rect 2339 206 2359 210
rect 2363 206 2439 210
rect 2443 206 2503 210
rect 2507 206 2534 210
rect 1305 205 2534 206
rect 96 145 97 151
rect 103 150 1311 151
rect 103 146 111 150
rect 115 146 151 150
rect 155 146 199 150
rect 203 146 207 150
rect 211 146 263 150
rect 267 146 295 150
rect 299 146 319 150
rect 323 146 375 150
rect 379 146 399 150
rect 403 146 431 150
rect 435 146 487 150
rect 491 146 503 150
rect 507 146 543 150
rect 547 146 599 150
rect 603 146 607 150
rect 611 146 655 150
rect 659 146 711 150
rect 715 146 767 150
rect 771 146 815 150
rect 819 146 831 150
rect 835 146 895 150
rect 899 146 911 150
rect 915 146 959 150
rect 963 146 1015 150
rect 1019 146 1023 150
rect 1027 146 1087 150
rect 1091 146 1119 150
rect 1123 146 1151 150
rect 1155 146 1287 150
rect 1291 146 1311 150
rect 103 145 1311 146
rect 1317 145 1318 151
rect 1310 133 1311 139
rect 1317 138 2539 139
rect 1317 134 1327 138
rect 1331 134 1367 138
rect 1371 134 1423 138
rect 1427 134 1479 138
rect 1483 134 1487 138
rect 1491 134 1535 138
rect 1539 134 1567 138
rect 1571 134 1591 138
rect 1595 134 1647 138
rect 1651 134 1655 138
rect 1659 134 1703 138
rect 1707 134 1735 138
rect 1739 134 1759 138
rect 1763 134 1823 138
rect 1827 134 1879 138
rect 1883 134 1911 138
rect 1915 134 1943 138
rect 1947 134 2007 138
rect 2011 134 2071 138
rect 2075 134 2119 138
rect 2123 134 2143 138
rect 2147 134 2223 138
rect 2227 134 2231 138
rect 2235 134 2303 138
rect 2307 134 2351 138
rect 2355 134 2391 138
rect 2395 134 2455 138
rect 2459 134 2503 138
rect 2507 134 2539 138
rect 1317 133 2539 134
rect 2545 133 2546 139
rect 84 93 85 99
rect 91 98 1299 99
rect 91 94 111 98
rect 115 94 135 98
rect 139 94 191 98
rect 195 94 247 98
rect 251 94 303 98
rect 307 94 359 98
rect 363 94 415 98
rect 419 94 471 98
rect 475 94 527 98
rect 531 94 583 98
rect 587 94 639 98
rect 643 94 695 98
rect 699 94 751 98
rect 755 94 815 98
rect 819 94 879 98
rect 883 94 943 98
rect 947 94 1007 98
rect 1011 94 1071 98
rect 1075 94 1135 98
rect 1139 94 1287 98
rect 1291 94 1299 98
rect 91 93 1299 94
rect 1305 93 1306 99
rect 1298 81 1299 87
rect 1305 86 2527 87
rect 1305 82 1327 86
rect 1331 82 1351 86
rect 1355 82 1407 86
rect 1411 82 1463 86
rect 1467 82 1519 86
rect 1523 82 1575 86
rect 1579 82 1631 86
rect 1635 82 1687 86
rect 1691 82 1743 86
rect 1747 82 1807 86
rect 1811 82 1863 86
rect 1867 82 1927 86
rect 1931 82 1991 86
rect 1995 82 2055 86
rect 2059 82 2127 86
rect 2131 82 2207 86
rect 2211 82 2287 86
rect 2291 82 2375 86
rect 2379 82 2439 86
rect 2443 82 2503 86
rect 2507 82 2527 86
rect 1305 81 2527 82
rect 2533 81 2534 87
<< m5c >>
rect 85 2577 91 2583
rect 1299 2577 1305 2583
rect 1299 2557 1305 2563
rect 2527 2557 2533 2563
rect 97 2525 103 2531
rect 1311 2525 1317 2531
rect 1311 2505 1317 2511
rect 2539 2505 2545 2511
rect 85 2465 91 2471
rect 1299 2465 1305 2471
rect 1299 2449 1305 2455
rect 2527 2449 2533 2455
rect 97 2401 103 2407
rect 1311 2401 1317 2407
rect 1311 2393 1317 2399
rect 2539 2393 2545 2399
rect 85 2341 91 2347
rect 1299 2341 1305 2347
rect 1299 2333 1305 2339
rect 2527 2333 2533 2339
rect 97 2281 103 2287
rect 1311 2281 1317 2287
rect 85 2229 91 2235
rect 1299 2229 1305 2235
rect 97 2177 103 2183
rect 1311 2177 1317 2183
rect 1311 2157 1317 2163
rect 2539 2157 2545 2163
rect 85 2125 91 2131
rect 1299 2125 1305 2131
rect 1299 2105 1305 2111
rect 2527 2105 2533 2111
rect 97 2069 103 2075
rect 1311 2069 1317 2075
rect 1311 2049 1317 2055
rect 2539 2049 2545 2055
rect 85 2013 91 2019
rect 1299 2013 1305 2019
rect 1299 1993 1305 1999
rect 2527 1993 2533 1999
rect 97 1957 103 1963
rect 1311 1957 1317 1963
rect 1311 1937 1317 1943
rect 2539 1937 2545 1943
rect 85 1897 91 1903
rect 1299 1897 1305 1903
rect 1299 1881 1305 1887
rect 2527 1881 2533 1887
rect 97 1845 103 1851
rect 1311 1845 1317 1851
rect 1311 1825 1317 1831
rect 2539 1825 2545 1831
rect 85 1781 91 1787
rect 1299 1781 1305 1787
rect 1299 1773 1305 1779
rect 2527 1773 2533 1779
rect 97 1725 103 1731
rect 1311 1725 1317 1731
rect 1311 1717 1317 1723
rect 2539 1717 2545 1723
rect 85 1669 91 1675
rect 1299 1669 1305 1675
rect 1299 1661 1305 1667
rect 2527 1661 2533 1667
rect 97 1613 103 1619
rect 1311 1613 1317 1619
rect 85 1561 91 1567
rect 1299 1561 1305 1567
rect 97 1501 103 1507
rect 1311 1501 1317 1507
rect 85 1445 91 1451
rect 1299 1445 1305 1451
rect 97 1389 103 1395
rect 1311 1389 1317 1395
rect 1299 1341 1305 1347
rect 2527 1341 2533 1347
rect 85 1321 91 1327
rect 1299 1321 1305 1327
rect 1311 1289 1317 1295
rect 2539 1289 2545 1295
rect 97 1261 103 1267
rect 1311 1261 1317 1267
rect 1299 1233 1305 1239
rect 2527 1233 2533 1239
rect 85 1205 91 1211
rect 1299 1205 1305 1211
rect 1311 1177 1317 1183
rect 2539 1177 2545 1183
rect 97 1149 103 1155
rect 1311 1149 1317 1155
rect 1299 1125 1305 1131
rect 2527 1125 2533 1131
rect 85 1089 91 1095
rect 1299 1089 1305 1095
rect 1311 1065 1317 1071
rect 2539 1065 2545 1071
rect 97 1029 103 1035
rect 1311 1029 1317 1035
rect 1299 1009 1305 1015
rect 2527 1009 2533 1015
rect 85 977 91 983
rect 1299 977 1305 983
rect 1311 945 1317 951
rect 2539 945 2545 951
rect 97 917 103 923
rect 1311 917 1317 923
rect 1299 889 1305 895
rect 2527 889 2533 895
rect 85 861 91 867
rect 1299 861 1305 867
rect 1311 833 1317 839
rect 2539 833 2545 839
rect 97 805 103 811
rect 1311 805 1317 811
rect 1299 777 1305 783
rect 2527 777 2533 783
rect 85 753 91 759
rect 1299 753 1305 759
rect 1311 725 1317 731
rect 2539 725 2545 731
rect 97 701 103 707
rect 1311 701 1317 707
rect 1299 661 1305 667
rect 2527 661 2533 667
rect 85 645 91 651
rect 1299 645 1305 651
rect 1311 609 1317 615
rect 2539 609 2545 615
rect 97 593 103 599
rect 1311 593 1317 599
rect 1299 557 1305 563
rect 2527 557 2533 563
rect 85 533 91 539
rect 1299 533 1305 539
rect 1311 501 1317 507
rect 2539 501 2545 507
rect 97 477 103 483
rect 1311 477 1317 483
rect 1299 437 1305 443
rect 2527 437 2533 443
rect 85 425 91 431
rect 1299 425 1305 431
rect 1311 381 1317 387
rect 2539 381 2545 387
rect 97 369 103 375
rect 1311 369 1317 375
rect 1299 321 1305 327
rect 2527 321 2533 327
rect 85 313 91 319
rect 1299 313 1305 319
rect 97 261 103 267
rect 1311 261 1317 267
rect 85 205 91 211
rect 1299 205 1305 211
rect 97 145 103 151
rect 1311 145 1317 151
rect 1311 133 1317 139
rect 2539 133 2545 139
rect 85 93 91 99
rect 1299 93 1305 99
rect 1299 81 1305 87
rect 2527 81 2533 87
<< m5 >>
rect 84 2583 92 2592
rect 84 2577 85 2583
rect 91 2577 92 2583
rect 84 2471 92 2577
rect 84 2465 85 2471
rect 91 2465 92 2471
rect 84 2347 92 2465
rect 84 2341 85 2347
rect 91 2341 92 2347
rect 84 2235 92 2341
rect 84 2229 85 2235
rect 91 2229 92 2235
rect 84 2131 92 2229
rect 84 2125 85 2131
rect 91 2125 92 2131
rect 84 2019 92 2125
rect 84 2013 85 2019
rect 91 2013 92 2019
rect 84 1903 92 2013
rect 84 1897 85 1903
rect 91 1897 92 1903
rect 84 1787 92 1897
rect 84 1781 85 1787
rect 91 1781 92 1787
rect 84 1675 92 1781
rect 84 1669 85 1675
rect 91 1669 92 1675
rect 84 1567 92 1669
rect 84 1561 85 1567
rect 91 1561 92 1567
rect 84 1451 92 1561
rect 84 1445 85 1451
rect 91 1445 92 1451
rect 84 1327 92 1445
rect 84 1321 85 1327
rect 91 1321 92 1327
rect 84 1211 92 1321
rect 84 1205 85 1211
rect 91 1205 92 1211
rect 84 1095 92 1205
rect 84 1089 85 1095
rect 91 1089 92 1095
rect 84 983 92 1089
rect 84 977 85 983
rect 91 977 92 983
rect 84 867 92 977
rect 84 861 85 867
rect 91 861 92 867
rect 84 759 92 861
rect 84 753 85 759
rect 91 753 92 759
rect 84 651 92 753
rect 84 645 85 651
rect 91 645 92 651
rect 84 539 92 645
rect 84 533 85 539
rect 91 533 92 539
rect 84 431 92 533
rect 84 425 85 431
rect 91 425 92 431
rect 84 319 92 425
rect 84 313 85 319
rect 91 313 92 319
rect 84 211 92 313
rect 84 205 85 211
rect 91 205 92 211
rect 84 99 92 205
rect 84 93 85 99
rect 91 93 92 99
rect 84 72 92 93
rect 96 2531 104 2592
rect 96 2525 97 2531
rect 103 2525 104 2531
rect 96 2407 104 2525
rect 96 2401 97 2407
rect 103 2401 104 2407
rect 96 2287 104 2401
rect 96 2281 97 2287
rect 103 2281 104 2287
rect 96 2183 104 2281
rect 96 2177 97 2183
rect 103 2177 104 2183
rect 96 2075 104 2177
rect 96 2069 97 2075
rect 103 2069 104 2075
rect 96 1963 104 2069
rect 96 1957 97 1963
rect 103 1957 104 1963
rect 96 1851 104 1957
rect 96 1845 97 1851
rect 103 1845 104 1851
rect 96 1731 104 1845
rect 96 1725 97 1731
rect 103 1725 104 1731
rect 96 1619 104 1725
rect 96 1613 97 1619
rect 103 1613 104 1619
rect 96 1507 104 1613
rect 96 1501 97 1507
rect 103 1501 104 1507
rect 96 1395 104 1501
rect 96 1389 97 1395
rect 103 1389 104 1395
rect 96 1267 104 1389
rect 96 1261 97 1267
rect 103 1261 104 1267
rect 96 1155 104 1261
rect 96 1149 97 1155
rect 103 1149 104 1155
rect 96 1035 104 1149
rect 96 1029 97 1035
rect 103 1029 104 1035
rect 96 923 104 1029
rect 96 917 97 923
rect 103 917 104 923
rect 96 811 104 917
rect 96 805 97 811
rect 103 805 104 811
rect 96 707 104 805
rect 96 701 97 707
rect 103 701 104 707
rect 96 599 104 701
rect 96 593 97 599
rect 103 593 104 599
rect 96 483 104 593
rect 96 477 97 483
rect 103 477 104 483
rect 96 375 104 477
rect 96 369 97 375
rect 103 369 104 375
rect 96 267 104 369
rect 96 261 97 267
rect 103 261 104 267
rect 96 151 104 261
rect 96 145 97 151
rect 103 145 104 151
rect 96 72 104 145
rect 1298 2583 1306 2592
rect 1298 2577 1299 2583
rect 1305 2577 1306 2583
rect 1298 2563 1306 2577
rect 1298 2557 1299 2563
rect 1305 2557 1306 2563
rect 1298 2471 1306 2557
rect 1298 2465 1299 2471
rect 1305 2465 1306 2471
rect 1298 2455 1306 2465
rect 1298 2449 1299 2455
rect 1305 2449 1306 2455
rect 1298 2347 1306 2449
rect 1298 2341 1299 2347
rect 1305 2341 1306 2347
rect 1298 2339 1306 2341
rect 1298 2333 1299 2339
rect 1305 2333 1306 2339
rect 1298 2235 1306 2333
rect 1298 2229 1299 2235
rect 1305 2229 1306 2235
rect 1298 2131 1306 2229
rect 1298 2125 1299 2131
rect 1305 2125 1306 2131
rect 1298 2111 1306 2125
rect 1298 2105 1299 2111
rect 1305 2105 1306 2111
rect 1298 2019 1306 2105
rect 1298 2013 1299 2019
rect 1305 2013 1306 2019
rect 1298 1999 1306 2013
rect 1298 1993 1299 1999
rect 1305 1993 1306 1999
rect 1298 1903 1306 1993
rect 1298 1897 1299 1903
rect 1305 1897 1306 1903
rect 1298 1887 1306 1897
rect 1298 1881 1299 1887
rect 1305 1881 1306 1887
rect 1298 1787 1306 1881
rect 1298 1781 1299 1787
rect 1305 1781 1306 1787
rect 1298 1779 1306 1781
rect 1298 1773 1299 1779
rect 1305 1773 1306 1779
rect 1298 1675 1306 1773
rect 1298 1669 1299 1675
rect 1305 1669 1306 1675
rect 1298 1667 1306 1669
rect 1298 1661 1299 1667
rect 1305 1661 1306 1667
rect 1298 1567 1306 1661
rect 1298 1561 1299 1567
rect 1305 1561 1306 1567
rect 1298 1451 1306 1561
rect 1298 1445 1299 1451
rect 1305 1445 1306 1451
rect 1298 1347 1306 1445
rect 1298 1341 1299 1347
rect 1305 1341 1306 1347
rect 1298 1327 1306 1341
rect 1298 1321 1299 1327
rect 1305 1321 1306 1327
rect 1298 1239 1306 1321
rect 1298 1233 1299 1239
rect 1305 1233 1306 1239
rect 1298 1211 1306 1233
rect 1298 1205 1299 1211
rect 1305 1205 1306 1211
rect 1298 1131 1306 1205
rect 1298 1125 1299 1131
rect 1305 1125 1306 1131
rect 1298 1095 1306 1125
rect 1298 1089 1299 1095
rect 1305 1089 1306 1095
rect 1298 1015 1306 1089
rect 1298 1009 1299 1015
rect 1305 1009 1306 1015
rect 1298 983 1306 1009
rect 1298 977 1299 983
rect 1305 977 1306 983
rect 1298 895 1306 977
rect 1298 889 1299 895
rect 1305 889 1306 895
rect 1298 867 1306 889
rect 1298 861 1299 867
rect 1305 861 1306 867
rect 1298 783 1306 861
rect 1298 777 1299 783
rect 1305 777 1306 783
rect 1298 759 1306 777
rect 1298 753 1299 759
rect 1305 753 1306 759
rect 1298 667 1306 753
rect 1298 661 1299 667
rect 1305 661 1306 667
rect 1298 651 1306 661
rect 1298 645 1299 651
rect 1305 645 1306 651
rect 1298 563 1306 645
rect 1298 557 1299 563
rect 1305 557 1306 563
rect 1298 539 1306 557
rect 1298 533 1299 539
rect 1305 533 1306 539
rect 1298 443 1306 533
rect 1298 437 1299 443
rect 1305 437 1306 443
rect 1298 431 1306 437
rect 1298 425 1299 431
rect 1305 425 1306 431
rect 1298 327 1306 425
rect 1298 321 1299 327
rect 1305 321 1306 327
rect 1298 319 1306 321
rect 1298 313 1299 319
rect 1305 313 1306 319
rect 1298 211 1306 313
rect 1298 205 1299 211
rect 1305 205 1306 211
rect 1298 99 1306 205
rect 1298 93 1299 99
rect 1305 93 1306 99
rect 1298 87 1306 93
rect 1298 81 1299 87
rect 1305 81 1306 87
rect 1298 72 1306 81
rect 1310 2531 1318 2592
rect 1310 2525 1311 2531
rect 1317 2525 1318 2531
rect 1310 2511 1318 2525
rect 1310 2505 1311 2511
rect 1317 2505 1318 2511
rect 1310 2407 1318 2505
rect 1310 2401 1311 2407
rect 1317 2401 1318 2407
rect 1310 2399 1318 2401
rect 1310 2393 1311 2399
rect 1317 2393 1318 2399
rect 1310 2287 1318 2393
rect 1310 2281 1311 2287
rect 1317 2281 1318 2287
rect 1310 2183 1318 2281
rect 1310 2177 1311 2183
rect 1317 2177 1318 2183
rect 1310 2163 1318 2177
rect 1310 2157 1311 2163
rect 1317 2157 1318 2163
rect 1310 2075 1318 2157
rect 1310 2069 1311 2075
rect 1317 2069 1318 2075
rect 1310 2055 1318 2069
rect 1310 2049 1311 2055
rect 1317 2049 1318 2055
rect 1310 1963 1318 2049
rect 1310 1957 1311 1963
rect 1317 1957 1318 1963
rect 1310 1943 1318 1957
rect 1310 1937 1311 1943
rect 1317 1937 1318 1943
rect 1310 1851 1318 1937
rect 1310 1845 1311 1851
rect 1317 1845 1318 1851
rect 1310 1831 1318 1845
rect 1310 1825 1311 1831
rect 1317 1825 1318 1831
rect 1310 1731 1318 1825
rect 1310 1725 1311 1731
rect 1317 1725 1318 1731
rect 1310 1723 1318 1725
rect 1310 1717 1311 1723
rect 1317 1717 1318 1723
rect 1310 1619 1318 1717
rect 1310 1613 1311 1619
rect 1317 1613 1318 1619
rect 1310 1507 1318 1613
rect 1310 1501 1311 1507
rect 1317 1501 1318 1507
rect 1310 1395 1318 1501
rect 1310 1389 1311 1395
rect 1317 1389 1318 1395
rect 1310 1295 1318 1389
rect 1310 1289 1311 1295
rect 1317 1289 1318 1295
rect 1310 1267 1318 1289
rect 1310 1261 1311 1267
rect 1317 1261 1318 1267
rect 1310 1183 1318 1261
rect 1310 1177 1311 1183
rect 1317 1177 1318 1183
rect 1310 1155 1318 1177
rect 1310 1149 1311 1155
rect 1317 1149 1318 1155
rect 1310 1071 1318 1149
rect 1310 1065 1311 1071
rect 1317 1065 1318 1071
rect 1310 1035 1318 1065
rect 1310 1029 1311 1035
rect 1317 1029 1318 1035
rect 1310 951 1318 1029
rect 1310 945 1311 951
rect 1317 945 1318 951
rect 1310 923 1318 945
rect 1310 917 1311 923
rect 1317 917 1318 923
rect 1310 839 1318 917
rect 1310 833 1311 839
rect 1317 833 1318 839
rect 1310 811 1318 833
rect 1310 805 1311 811
rect 1317 805 1318 811
rect 1310 731 1318 805
rect 1310 725 1311 731
rect 1317 725 1318 731
rect 1310 707 1318 725
rect 1310 701 1311 707
rect 1317 701 1318 707
rect 1310 615 1318 701
rect 1310 609 1311 615
rect 1317 609 1318 615
rect 1310 599 1318 609
rect 1310 593 1311 599
rect 1317 593 1318 599
rect 1310 507 1318 593
rect 1310 501 1311 507
rect 1317 501 1318 507
rect 1310 483 1318 501
rect 1310 477 1311 483
rect 1317 477 1318 483
rect 1310 387 1318 477
rect 1310 381 1311 387
rect 1317 381 1318 387
rect 1310 375 1318 381
rect 1310 369 1311 375
rect 1317 369 1318 375
rect 1310 267 1318 369
rect 1310 261 1311 267
rect 1317 261 1318 267
rect 1310 151 1318 261
rect 1310 145 1311 151
rect 1317 145 1318 151
rect 1310 139 1318 145
rect 1310 133 1311 139
rect 1317 133 1318 139
rect 1310 72 1318 133
rect 2526 2563 2534 2592
rect 2526 2557 2527 2563
rect 2533 2557 2534 2563
rect 2526 2455 2534 2557
rect 2526 2449 2527 2455
rect 2533 2449 2534 2455
rect 2526 2339 2534 2449
rect 2526 2333 2527 2339
rect 2533 2333 2534 2339
rect 2526 2111 2534 2333
rect 2526 2105 2527 2111
rect 2533 2105 2534 2111
rect 2526 1999 2534 2105
rect 2526 1993 2527 1999
rect 2533 1993 2534 1999
rect 2526 1887 2534 1993
rect 2526 1881 2527 1887
rect 2533 1881 2534 1887
rect 2526 1779 2534 1881
rect 2526 1773 2527 1779
rect 2533 1773 2534 1779
rect 2526 1667 2534 1773
rect 2526 1661 2527 1667
rect 2533 1661 2534 1667
rect 2526 1347 2534 1661
rect 2526 1341 2527 1347
rect 2533 1341 2534 1347
rect 2526 1239 2534 1341
rect 2526 1233 2527 1239
rect 2533 1233 2534 1239
rect 2526 1131 2534 1233
rect 2526 1125 2527 1131
rect 2533 1125 2534 1131
rect 2526 1015 2534 1125
rect 2526 1009 2527 1015
rect 2533 1009 2534 1015
rect 2526 895 2534 1009
rect 2526 889 2527 895
rect 2533 889 2534 895
rect 2526 783 2534 889
rect 2526 777 2527 783
rect 2533 777 2534 783
rect 2526 667 2534 777
rect 2526 661 2527 667
rect 2533 661 2534 667
rect 2526 563 2534 661
rect 2526 557 2527 563
rect 2533 557 2534 563
rect 2526 443 2534 557
rect 2526 437 2527 443
rect 2533 437 2534 443
rect 2526 327 2534 437
rect 2526 321 2527 327
rect 2533 321 2534 327
rect 2526 87 2534 321
rect 2526 81 2527 87
rect 2533 81 2534 87
rect 2526 72 2534 81
rect 2538 2511 2546 2592
rect 2538 2505 2539 2511
rect 2545 2505 2546 2511
rect 2538 2399 2546 2505
rect 2538 2393 2539 2399
rect 2545 2393 2546 2399
rect 2538 2163 2546 2393
rect 2538 2157 2539 2163
rect 2545 2157 2546 2163
rect 2538 2055 2546 2157
rect 2538 2049 2539 2055
rect 2545 2049 2546 2055
rect 2538 1943 2546 2049
rect 2538 1937 2539 1943
rect 2545 1937 2546 1943
rect 2538 1831 2546 1937
rect 2538 1825 2539 1831
rect 2545 1825 2546 1831
rect 2538 1723 2546 1825
rect 2538 1717 2539 1723
rect 2545 1717 2546 1723
rect 2538 1295 2546 1717
rect 2538 1289 2539 1295
rect 2545 1289 2546 1295
rect 2538 1183 2546 1289
rect 2538 1177 2539 1183
rect 2545 1177 2546 1183
rect 2538 1071 2546 1177
rect 2538 1065 2539 1071
rect 2545 1065 2546 1071
rect 2538 951 2546 1065
rect 2538 945 2539 951
rect 2545 945 2546 951
rect 2538 839 2546 945
rect 2538 833 2539 839
rect 2545 833 2546 839
rect 2538 731 2546 833
rect 2538 725 2539 731
rect 2545 725 2546 731
rect 2538 615 2546 725
rect 2538 609 2539 615
rect 2545 609 2546 615
rect 2538 507 2546 609
rect 2538 501 2539 507
rect 2545 501 2546 507
rect 2538 387 2546 501
rect 2538 381 2539 387
rect 2545 381 2546 387
rect 2538 139 2546 381
rect 2538 133 2539 139
rect 2545 133 2546 139
rect 2538 72 2546 133
use circuitwell  npwells
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use circuitppnp  ppnps
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use welltap_svt  __well_tap__175
timestamp 1731220653
transform 1 0 2496 0 -1 2556
box 7 3 12 24
use welltap_svt  __well_tap__174
timestamp 1731220653
transform 1 0 1320 0 -1 2556
box 7 3 12 24
use welltap_svt  __well_tap__173
timestamp 1731220653
transform 1 0 2496 0 1 2460
box 7 3 12 24
use welltap_svt  __well_tap__172
timestamp 1731220653
transform 1 0 1320 0 1 2460
box 7 3 12 24
use welltap_svt  __well_tap__171
timestamp 1731220653
transform 1 0 2496 0 -1 2448
box 7 3 12 24
use welltap_svt  __well_tap__170
timestamp 1731220653
transform 1 0 1320 0 -1 2448
box 7 3 12 24
use welltap_svt  __well_tap__169
timestamp 1731220653
transform 1 0 2496 0 1 2348
box 7 3 12 24
use welltap_svt  __well_tap__168
timestamp 1731220653
transform 1 0 1320 0 1 2348
box 7 3 12 24
use welltap_svt  __well_tap__167
timestamp 1731220653
transform 1 0 2496 0 -1 2332
box 7 3 12 24
use welltap_svt  __well_tap__166
timestamp 1731220653
transform 1 0 1320 0 -1 2332
box 7 3 12 24
use welltap_svt  __well_tap__165
timestamp 1731220653
transform 1 0 2496 0 1 2236
box 7 3 12 24
use welltap_svt  __well_tap__164
timestamp 1731220653
transform 1 0 1320 0 1 2236
box 7 3 12 24
use welltap_svt  __well_tap__163
timestamp 1731220653
transform 1 0 2496 0 -1 2228
box 7 3 12 24
use welltap_svt  __well_tap__162
timestamp 1731220653
transform 1 0 1320 0 -1 2228
box 7 3 12 24
use welltap_svt  __well_tap__161
timestamp 1731220653
transform 1 0 2496 0 1 2112
box 7 3 12 24
use welltap_svt  __well_tap__160
timestamp 1731220653
transform 1 0 1320 0 1 2112
box 7 3 12 24
use welltap_svt  __well_tap__159
timestamp 1731220653
transform 1 0 2496 0 -1 2104
box 7 3 12 24
use welltap_svt  __well_tap__158
timestamp 1731220653
transform 1 0 1320 0 -1 2104
box 7 3 12 24
use welltap_svt  __well_tap__157
timestamp 1731220653
transform 1 0 2496 0 1 2004
box 7 3 12 24
use welltap_svt  __well_tap__156
timestamp 1731220653
transform 1 0 1320 0 1 2004
box 7 3 12 24
use welltap_svt  __well_tap__155
timestamp 1731220653
transform 1 0 2496 0 -1 1992
box 7 3 12 24
use welltap_svt  __well_tap__154
timestamp 1731220653
transform 1 0 1320 0 -1 1992
box 7 3 12 24
use welltap_svt  __well_tap__153
timestamp 1731220653
transform 1 0 2496 0 1 1892
box 7 3 12 24
use welltap_svt  __well_tap__152
timestamp 1731220653
transform 1 0 1320 0 1 1892
box 7 3 12 24
use welltap_svt  __well_tap__151
timestamp 1731220653
transform 1 0 2496 0 -1 1880
box 7 3 12 24
use welltap_svt  __well_tap__150
timestamp 1731220653
transform 1 0 1320 0 -1 1880
box 7 3 12 24
use welltap_svt  __well_tap__149
timestamp 1731220653
transform 1 0 2496 0 1 1780
box 7 3 12 24
use welltap_svt  __well_tap__148
timestamp 1731220653
transform 1 0 1320 0 1 1780
box 7 3 12 24
use welltap_svt  __well_tap__147
timestamp 1731220653
transform 1 0 2496 0 -1 1772
box 7 3 12 24
use welltap_svt  __well_tap__146
timestamp 1731220653
transform 1 0 1320 0 -1 1772
box 7 3 12 24
use welltap_svt  __well_tap__145
timestamp 1731220653
transform 1 0 2496 0 1 1672
box 7 3 12 24
use welltap_svt  __well_tap__144
timestamp 1731220653
transform 1 0 1320 0 1 1672
box 7 3 12 24
use welltap_svt  __well_tap__143
timestamp 1731220653
transform 1 0 2496 0 -1 1660
box 7 3 12 24
use welltap_svt  __well_tap__142
timestamp 1731220653
transform 1 0 1320 0 -1 1660
box 7 3 12 24
use welltap_svt  __well_tap__141
timestamp 1731220653
transform 1 0 2496 0 1 1564
box 7 3 12 24
use welltap_svt  __well_tap__140
timestamp 1731220653
transform 1 0 1320 0 1 1564
box 7 3 12 24
use welltap_svt  __well_tap__139
timestamp 1731220653
transform 1 0 2496 0 -1 1556
box 7 3 12 24
use welltap_svt  __well_tap__138
timestamp 1731220653
transform 1 0 1320 0 -1 1556
box 7 3 12 24
use welltap_svt  __well_tap__137
timestamp 1731220653
transform 1 0 2496 0 1 1460
box 7 3 12 24
use welltap_svt  __well_tap__136
timestamp 1731220653
transform 1 0 1320 0 1 1460
box 7 3 12 24
use welltap_svt  __well_tap__135
timestamp 1731220653
transform 1 0 2496 0 -1 1444
box 7 3 12 24
use welltap_svt  __well_tap__134
timestamp 1731220653
transform 1 0 1320 0 -1 1444
box 7 3 12 24
use welltap_svt  __well_tap__133
timestamp 1731220653
transform 1 0 2496 0 1 1348
box 7 3 12 24
use welltap_svt  __well_tap__132
timestamp 1731220653
transform 1 0 1320 0 1 1348
box 7 3 12 24
use welltap_svt  __well_tap__131
timestamp 1731220653
transform 1 0 2496 0 -1 1340
box 7 3 12 24
use welltap_svt  __well_tap__130
timestamp 1731220653
transform 1 0 1320 0 -1 1340
box 7 3 12 24
use welltap_svt  __well_tap__129
timestamp 1731220653
transform 1 0 2496 0 1 1244
box 7 3 12 24
use welltap_svt  __well_tap__128
timestamp 1731220653
transform 1 0 1320 0 1 1244
box 7 3 12 24
use welltap_svt  __well_tap__127
timestamp 1731220653
transform 1 0 2496 0 -1 1232
box 7 3 12 24
use welltap_svt  __well_tap__126
timestamp 1731220653
transform 1 0 1320 0 -1 1232
box 7 3 12 24
use welltap_svt  __well_tap__125
timestamp 1731220653
transform 1 0 2496 0 1 1132
box 7 3 12 24
use welltap_svt  __well_tap__124
timestamp 1731220653
transform 1 0 1320 0 1 1132
box 7 3 12 24
use welltap_svt  __well_tap__123
timestamp 1731220653
transform 1 0 2496 0 -1 1124
box 7 3 12 24
use welltap_svt  __well_tap__122
timestamp 1731220653
transform 1 0 1320 0 -1 1124
box 7 3 12 24
use welltap_svt  __well_tap__121
timestamp 1731220653
transform 1 0 2496 0 1 1020
box 7 3 12 24
use welltap_svt  __well_tap__120
timestamp 1731220653
transform 1 0 1320 0 1 1020
box 7 3 12 24
use welltap_svt  __well_tap__119
timestamp 1731220653
transform 1 0 2496 0 -1 1008
box 7 3 12 24
use welltap_svt  __well_tap__118
timestamp 1731220653
transform 1 0 1320 0 -1 1008
box 7 3 12 24
use welltap_svt  __well_tap__117
timestamp 1731220653
transform 1 0 2496 0 1 900
box 7 3 12 24
use welltap_svt  __well_tap__116
timestamp 1731220653
transform 1 0 1320 0 1 900
box 7 3 12 24
use welltap_svt  __well_tap__115
timestamp 1731220653
transform 1 0 2496 0 -1 888
box 7 3 12 24
use welltap_svt  __well_tap__114
timestamp 1731220653
transform 1 0 1320 0 -1 888
box 7 3 12 24
use welltap_svt  __well_tap__113
timestamp 1731220653
transform 1 0 2496 0 1 788
box 7 3 12 24
use welltap_svt  __well_tap__112
timestamp 1731220653
transform 1 0 1320 0 1 788
box 7 3 12 24
use welltap_svt  __well_tap__111
timestamp 1731220653
transform 1 0 2496 0 -1 776
box 7 3 12 24
use welltap_svt  __well_tap__110
timestamp 1731220653
transform 1 0 1320 0 -1 776
box 7 3 12 24
use welltap_svt  __well_tap__109
timestamp 1731220653
transform 1 0 2496 0 1 680
box 7 3 12 24
use welltap_svt  __well_tap__108
timestamp 1731220653
transform 1 0 1320 0 1 680
box 7 3 12 24
use welltap_svt  __well_tap__107
timestamp 1731220653
transform 1 0 2496 0 -1 660
box 7 3 12 24
use welltap_svt  __well_tap__106
timestamp 1731220653
transform 1 0 1320 0 -1 660
box 7 3 12 24
use welltap_svt  __well_tap__105
timestamp 1731220653
transform 1 0 2496 0 1 564
box 7 3 12 24
use welltap_svt  __well_tap__104
timestamp 1731220653
transform 1 0 1320 0 1 564
box 7 3 12 24
use welltap_svt  __well_tap__103
timestamp 1731220653
transform 1 0 2496 0 -1 556
box 7 3 12 24
use welltap_svt  __well_tap__102
timestamp 1731220653
transform 1 0 1320 0 -1 556
box 7 3 12 24
use welltap_svt  __well_tap__101
timestamp 1731220653
transform 1 0 2496 0 1 456
box 7 3 12 24
use welltap_svt  __well_tap__100
timestamp 1731220653
transform 1 0 1320 0 1 456
box 7 3 12 24
use welltap_svt  __well_tap__99
timestamp 1731220653
transform 1 0 2496 0 -1 436
box 7 3 12 24
use welltap_svt  __well_tap__98
timestamp 1731220653
transform 1 0 1320 0 -1 436
box 7 3 12 24
use welltap_svt  __well_tap__97
timestamp 1731220653
transform 1 0 2496 0 1 336
box 7 3 12 24
use welltap_svt  __well_tap__96
timestamp 1731220653
transform 1 0 1320 0 1 336
box 7 3 12 24
use welltap_svt  __well_tap__95
timestamp 1731220653
transform 1 0 2496 0 -1 320
box 7 3 12 24
use welltap_svt  __well_tap__94
timestamp 1731220653
transform 1 0 1320 0 -1 320
box 7 3 12 24
use welltap_svt  __well_tap__93
timestamp 1731220653
transform 1 0 2496 0 1 216
box 7 3 12 24
use welltap_svt  __well_tap__92
timestamp 1731220653
transform 1 0 1320 0 1 216
box 7 3 12 24
use welltap_svt  __well_tap__91
timestamp 1731220653
transform 1 0 2496 0 -1 204
box 7 3 12 24
use welltap_svt  __well_tap__90
timestamp 1731220653
transform 1 0 1320 0 -1 204
box 7 3 12 24
use welltap_svt  __well_tap__89
timestamp 1731220653
transform 1 0 2496 0 1 88
box 7 3 12 24
use welltap_svt  __well_tap__88
timestamp 1731220653
transform 1 0 1320 0 1 88
box 7 3 12 24
use welltap_svt  __well_tap__87
timestamp 1731220653
transform 1 0 1280 0 -1 2576
box 7 3 12 24
use welltap_svt  __well_tap__86
timestamp 1731220653
transform 1 0 104 0 -1 2576
box 7 3 12 24
use welltap_svt  __well_tap__85
timestamp 1731220653
transform 1 0 1280 0 1 2480
box 7 3 12 24
use welltap_svt  __well_tap__84
timestamp 1731220653
transform 1 0 104 0 1 2480
box 7 3 12 24
use welltap_svt  __well_tap__83
timestamp 1731220653
transform 1 0 1280 0 -1 2464
box 7 3 12 24
use welltap_svt  __well_tap__82
timestamp 1731220653
transform 1 0 104 0 -1 2464
box 7 3 12 24
use welltap_svt  __well_tap__81
timestamp 1731220653
transform 1 0 1280 0 1 2356
box 7 3 12 24
use welltap_svt  __well_tap__80
timestamp 1731220653
transform 1 0 104 0 1 2356
box 7 3 12 24
use welltap_svt  __well_tap__79
timestamp 1731220653
transform 1 0 1280 0 -1 2340
box 7 3 12 24
use welltap_svt  __well_tap__78
timestamp 1731220653
transform 1 0 104 0 -1 2340
box 7 3 12 24
use welltap_svt  __well_tap__77
timestamp 1731220653
transform 1 0 1280 0 1 2236
box 7 3 12 24
use welltap_svt  __well_tap__76
timestamp 1731220653
transform 1 0 104 0 1 2236
box 7 3 12 24
use welltap_svt  __well_tap__75
timestamp 1731220653
transform 1 0 1280 0 -1 2228
box 7 3 12 24
use welltap_svt  __well_tap__74
timestamp 1731220653
transform 1 0 104 0 -1 2228
box 7 3 12 24
use welltap_svt  __well_tap__73
timestamp 1731220653
transform 1 0 1280 0 1 2132
box 7 3 12 24
use welltap_svt  __well_tap__72
timestamp 1731220653
transform 1 0 104 0 1 2132
box 7 3 12 24
use welltap_svt  __well_tap__71
timestamp 1731220653
transform 1 0 1280 0 -1 2124
box 7 3 12 24
use welltap_svt  __well_tap__70
timestamp 1731220653
transform 1 0 104 0 -1 2124
box 7 3 12 24
use welltap_svt  __well_tap__69
timestamp 1731220653
transform 1 0 1280 0 1 2024
box 7 3 12 24
use welltap_svt  __well_tap__68
timestamp 1731220653
transform 1 0 104 0 1 2024
box 7 3 12 24
use welltap_svt  __well_tap__67
timestamp 1731220653
transform 1 0 1280 0 -1 2012
box 7 3 12 24
use welltap_svt  __well_tap__66
timestamp 1731220653
transform 1 0 104 0 -1 2012
box 7 3 12 24
use welltap_svt  __well_tap__65
timestamp 1731220653
transform 1 0 1280 0 1 1912
box 7 3 12 24
use welltap_svt  __well_tap__64
timestamp 1731220653
transform 1 0 104 0 1 1912
box 7 3 12 24
use welltap_svt  __well_tap__63
timestamp 1731220653
transform 1 0 1280 0 -1 1896
box 7 3 12 24
use welltap_svt  __well_tap__62
timestamp 1731220653
transform 1 0 104 0 -1 1896
box 7 3 12 24
use welltap_svt  __well_tap__61
timestamp 1731220653
transform 1 0 1280 0 1 1800
box 7 3 12 24
use welltap_svt  __well_tap__60
timestamp 1731220653
transform 1 0 104 0 1 1800
box 7 3 12 24
use welltap_svt  __well_tap__59
timestamp 1731220653
transform 1 0 1280 0 -1 1780
box 7 3 12 24
use welltap_svt  __well_tap__58
timestamp 1731220653
transform 1 0 104 0 -1 1780
box 7 3 12 24
use welltap_svt  __well_tap__57
timestamp 1731220653
transform 1 0 1280 0 1 1680
box 7 3 12 24
use welltap_svt  __well_tap__56
timestamp 1731220653
transform 1 0 104 0 1 1680
box 7 3 12 24
use welltap_svt  __well_tap__55
timestamp 1731220653
transform 1 0 1280 0 -1 1668
box 7 3 12 24
use welltap_svt  __well_tap__54
timestamp 1731220653
transform 1 0 104 0 -1 1668
box 7 3 12 24
use welltap_svt  __well_tap__53
timestamp 1731220653
transform 1 0 1280 0 1 1568
box 7 3 12 24
use welltap_svt  __well_tap__52
timestamp 1731220653
transform 1 0 104 0 1 1568
box 7 3 12 24
use welltap_svt  __well_tap__51
timestamp 1731220653
transform 1 0 1280 0 -1 1560
box 7 3 12 24
use welltap_svt  __well_tap__50
timestamp 1731220653
transform 1 0 104 0 -1 1560
box 7 3 12 24
use welltap_svt  __well_tap__49
timestamp 1731220653
transform 1 0 1280 0 1 1456
box 7 3 12 24
use welltap_svt  __well_tap__48
timestamp 1731220653
transform 1 0 104 0 1 1456
box 7 3 12 24
use welltap_svt  __well_tap__47
timestamp 1731220653
transform 1 0 1280 0 -1 1444
box 7 3 12 24
use welltap_svt  __well_tap__46
timestamp 1731220653
transform 1 0 104 0 -1 1444
box 7 3 12 24
use welltap_svt  __well_tap__45
timestamp 1731220653
transform 1 0 1280 0 1 1344
box 7 3 12 24
use welltap_svt  __well_tap__44
timestamp 1731220653
transform 1 0 104 0 1 1344
box 7 3 12 24
use welltap_svt  __well_tap__43
timestamp 1731220653
transform 1 0 1280 0 -1 1320
box 7 3 12 24
use welltap_svt  __well_tap__42
timestamp 1731220653
transform 1 0 104 0 -1 1320
box 7 3 12 24
use welltap_svt  __well_tap__41
timestamp 1731220653
transform 1 0 1280 0 1 1216
box 7 3 12 24
use welltap_svt  __well_tap__40
timestamp 1731220653
transform 1 0 104 0 1 1216
box 7 3 12 24
use welltap_svt  __well_tap__39
timestamp 1731220653
transform 1 0 1280 0 -1 1204
box 7 3 12 24
use welltap_svt  __well_tap__38
timestamp 1731220653
transform 1 0 104 0 -1 1204
box 7 3 12 24
use welltap_svt  __well_tap__37
timestamp 1731220653
transform 1 0 1280 0 1 1104
box 7 3 12 24
use welltap_svt  __well_tap__36
timestamp 1731220653
transform 1 0 104 0 1 1104
box 7 3 12 24
use welltap_svt  __well_tap__35
timestamp 1731220653
transform 1 0 1280 0 -1 1088
box 7 3 12 24
use welltap_svt  __well_tap__34
timestamp 1731220653
transform 1 0 104 0 -1 1088
box 7 3 12 24
use welltap_svt  __well_tap__33
timestamp 1731220653
transform 1 0 1280 0 1 984
box 7 3 12 24
use welltap_svt  __well_tap__32
timestamp 1731220653
transform 1 0 104 0 1 984
box 7 3 12 24
use welltap_svt  __well_tap__31
timestamp 1731220653
transform 1 0 1280 0 -1 976
box 7 3 12 24
use welltap_svt  __well_tap__30
timestamp 1731220653
transform 1 0 104 0 -1 976
box 7 3 12 24
use welltap_svt  __well_tap__29
timestamp 1731220653
transform 1 0 1280 0 1 872
box 7 3 12 24
use welltap_svt  __well_tap__28
timestamp 1731220653
transform 1 0 104 0 1 872
box 7 3 12 24
use welltap_svt  __well_tap__27
timestamp 1731220653
transform 1 0 1280 0 -1 860
box 7 3 12 24
use welltap_svt  __well_tap__26
timestamp 1731220653
transform 1 0 104 0 -1 860
box 7 3 12 24
use welltap_svt  __well_tap__25
timestamp 1731220653
transform 1 0 1280 0 1 760
box 7 3 12 24
use welltap_svt  __well_tap__24
timestamp 1731220653
transform 1 0 104 0 1 760
box 7 3 12 24
use welltap_svt  __well_tap__23
timestamp 1731220653
transform 1 0 1280 0 -1 752
box 7 3 12 24
use welltap_svt  __well_tap__22
timestamp 1731220653
transform 1 0 104 0 -1 752
box 7 3 12 24
use welltap_svt  __well_tap__21
timestamp 1731220653
transform 1 0 1280 0 1 656
box 7 3 12 24
use welltap_svt  __well_tap__20
timestamp 1731220653
transform 1 0 104 0 1 656
box 7 3 12 24
use welltap_svt  __well_tap__19
timestamp 1731220653
transform 1 0 1280 0 -1 644
box 7 3 12 24
use welltap_svt  __well_tap__18
timestamp 1731220653
transform 1 0 104 0 -1 644
box 7 3 12 24
use welltap_svt  __well_tap__17
timestamp 1731220653
transform 1 0 1280 0 1 548
box 7 3 12 24
use welltap_svt  __well_tap__16
timestamp 1731220653
transform 1 0 104 0 1 548
box 7 3 12 24
use welltap_svt  __well_tap__15
timestamp 1731220653
transform 1 0 1280 0 -1 532
box 7 3 12 24
use welltap_svt  __well_tap__14
timestamp 1731220653
transform 1 0 104 0 -1 532
box 7 3 12 24
use welltap_svt  __well_tap__13
timestamp 1731220653
transform 1 0 1280 0 1 432
box 7 3 12 24
use welltap_svt  __well_tap__12
timestamp 1731220653
transform 1 0 104 0 1 432
box 7 3 12 24
use welltap_svt  __well_tap__11
timestamp 1731220653
transform 1 0 1280 0 -1 424
box 7 3 12 24
use welltap_svt  __well_tap__10
timestamp 1731220653
transform 1 0 104 0 -1 424
box 7 3 12 24
use welltap_svt  __well_tap__9
timestamp 1731220653
transform 1 0 1280 0 1 324
box 7 3 12 24
use welltap_svt  __well_tap__8
timestamp 1731220653
transform 1 0 104 0 1 324
box 7 3 12 24
use welltap_svt  __well_tap__7
timestamp 1731220653
transform 1 0 1280 0 -1 312
box 7 3 12 24
use welltap_svt  __well_tap__6
timestamp 1731220653
transform 1 0 104 0 -1 312
box 7 3 12 24
use welltap_svt  __well_tap__5
timestamp 1731220653
transform 1 0 1280 0 1 216
box 7 3 12 24
use welltap_svt  __well_tap__4
timestamp 1731220653
transform 1 0 104 0 1 216
box 7 3 12 24
use welltap_svt  __well_tap__3
timestamp 1731220653
transform 1 0 1280 0 -1 204
box 7 3 12 24
use welltap_svt  __well_tap__2
timestamp 1731220653
transform 1 0 104 0 -1 204
box 7 3 12 24
use welltap_svt  __well_tap__1
timestamp 1731220653
transform 1 0 1280 0 1 100
box 7 3 12 24
use welltap_svt  __well_tap__0
timestamp 1731220653
transform 1 0 104 0 1 100
box 7 3 12 24
use _0_0std_0_0cells_0_0OR2X1  tst_5999_6
timestamp 1731220653
transform 1 0 2368 0 1 84
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5998_6
timestamp 1731220653
transform 1 0 2432 0 1 84
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5997_6
timestamp 1731220653
transform 1 0 2432 0 -1 208
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5996_6
timestamp 1731220653
transform 1 0 2432 0 1 212
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5995_6
timestamp 1731220653
transform 1 0 2352 0 1 212
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5994_6
timestamp 1731220653
transform 1 0 2256 0 -1 324
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5993_6
timestamp 1731220653
transform 1 0 2352 0 -1 324
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5992_6
timestamp 1731220653
transform 1 0 2352 0 1 332
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5991_6
timestamp 1731220653
transform 1 0 2360 0 -1 440
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5990_6
timestamp 1731220653
transform 1 0 2360 0 1 452
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5989_6
timestamp 1731220653
transform 1 0 2272 0 1 452
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5988_6
timestamp 1731220653
transform 1 0 2248 0 -1 560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5987_6
timestamp 1731220653
transform 1 0 2144 0 -1 560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5986_6
timestamp 1731220653
transform 1 0 2048 0 -1 560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5985_6
timestamp 1731220653
transform 1 0 2184 0 1 560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5984_6
timestamp 1731220653
transform 1 0 2320 0 1 560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5983_6
timestamp 1731220653
transform 1 0 2312 0 -1 664
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5982_6
timestamp 1731220653
transform 1 0 2176 0 -1 664
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5981_6
timestamp 1731220653
transform 1 0 2048 0 -1 664
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5980_6
timestamp 1731220653
transform 1 0 2024 0 1 676
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5979_6
timestamp 1731220653
transform 1 0 1920 0 1 676
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5978_6
timestamp 1731220653
transform 1 0 1816 0 1 676
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5977_6
timestamp 1731220653
transform 1 0 1816 0 -1 664
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5976_6
timestamp 1731220653
transform 1 0 1928 0 -1 664
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5975_6
timestamp 1731220653
transform 1 0 2056 0 1 560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5974_6
timestamp 1731220653
transform 1 0 1936 0 1 560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5973_6
timestamp 1731220653
transform 1 0 1824 0 1 560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5972_6
timestamp 1731220653
transform 1 0 1848 0 -1 560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5971_6
timestamp 1731220653
transform 1 0 1952 0 -1 560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5970_6
timestamp 1731220653
transform 1 0 1896 0 1 452
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5969_6
timestamp 1731220653
transform 1 0 1920 0 1 332
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5968_6
timestamp 1731220653
transform 1 0 1832 0 -1 324
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5967_6
timestamp 1731220653
transform 1 0 1944 0 -1 324
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5966_6
timestamp 1731220653
transform 1 0 1944 0 1 212
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5965_6
timestamp 1731220653
transform 1 0 1840 0 1 212
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5964_6
timestamp 1731220653
transform 1 0 1800 0 -1 208
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5963_6
timestamp 1731220653
transform 1 0 1888 0 -1 208
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5962_6
timestamp 1731220653
transform 1 0 1984 0 -1 208
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5961_6
timestamp 1731220653
transform 1 0 1920 0 1 84
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5960_6
timestamp 1731220653
transform 1 0 1856 0 1 84
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5959_6
timestamp 1731220653
transform 1 0 1800 0 1 84
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5958_6
timestamp 1731220653
transform 1 0 1984 0 1 84
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5957_6
timestamp 1731220653
transform 1 0 2048 0 1 84
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5956_6
timestamp 1731220653
transform 1 0 2280 0 1 84
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5955_6
timestamp 1731220653
transform 1 0 2200 0 1 84
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5954_6
timestamp 1731220653
transform 1 0 2120 0 1 84
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5953_6
timestamp 1731220653
transform 1 0 2096 0 -1 208
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5952_6
timestamp 1731220653
transform 1 0 2208 0 -1 208
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5951_6
timestamp 1731220653
transform 1 0 2328 0 -1 208
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5950_6
timestamp 1731220653
transform 1 0 2248 0 1 212
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5949_6
timestamp 1731220653
transform 1 0 2152 0 1 212
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5948_6
timestamp 1731220653
transform 1 0 2048 0 1 212
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5947_6
timestamp 1731220653
transform 1 0 2056 0 -1 324
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5946_6
timestamp 1731220653
transform 1 0 2160 0 -1 324
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5945_6
timestamp 1731220653
transform 1 0 2176 0 1 332
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5944_6
timestamp 1731220653
transform 1 0 2264 0 1 332
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5943_6
timestamp 1731220653
transform 1 0 2264 0 -1 440
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5942_6
timestamp 1731220653
transform 1 0 2168 0 -1 440
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5941_6
timestamp 1731220653
transform 1 0 2096 0 1 452
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5940_6
timestamp 1731220653
transform 1 0 2000 0 1 452
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5939_6
timestamp 1731220653
transform 1 0 2184 0 1 452
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5938_6
timestamp 1731220653
transform 1 0 2352 0 -1 560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5937_6
timestamp 1731220653
transform 1 0 2432 0 1 452
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5936_6
timestamp 1731220653
transform 1 0 2432 0 1 332
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5935_6
timestamp 1731220653
transform 1 0 2432 0 -1 324
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5934_6
timestamp 1731220653
transform 1 0 2432 0 -1 440
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5933_6
timestamp 1731220653
transform 1 0 2432 0 -1 560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5932_6
timestamp 1731220653
transform 1 0 2432 0 1 560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5931_6
timestamp 1731220653
transform 1 0 2432 0 -1 664
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5930_6
timestamp 1731220653
transform 1 0 2432 0 1 676
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5929_6
timestamp 1731220653
transform 1 0 2432 0 -1 780
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5928_6
timestamp 1731220653
transform 1 0 2432 0 1 784
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5927_6
timestamp 1731220653
transform 1 0 2432 0 1 896
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5926_6
timestamp 1731220653
transform 1 0 2432 0 1 1016
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5925_6
timestamp 1731220653
transform 1 0 2432 0 1 1128
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5924_6
timestamp 1731220653
transform 1 0 2432 0 -1 1236
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5923_6
timestamp 1731220653
transform 1 0 2432 0 -1 1344
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5922_6
timestamp 1731220653
transform 1 0 2432 0 1 1344
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5921_6
timestamp 1731220653
transform 1 0 2376 0 1 1344
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5920_6
timestamp 1731220653
transform 1 0 2376 0 -1 1344
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5919_6
timestamp 1731220653
transform 1 0 2360 0 -1 1236
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5918_6
timestamp 1731220653
transform 1 0 2432 0 -1 1012
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5917_6
timestamp 1731220653
transform 1 0 2416 0 -1 892
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5916_6
timestamp 1731220653
transform 1 0 2360 0 1 784
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5915_6
timestamp 1731220653
transform 1 0 2264 0 1 784
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5914_6
timestamp 1731220653
transform 1 0 2168 0 1 784
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5913_6
timestamp 1731220653
transform 1 0 2336 0 -1 780
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5912_6
timestamp 1731220653
transform 1 0 2344 0 1 676
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5911_6
timestamp 1731220653
transform 1 0 2232 0 1 676
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5910_6
timestamp 1731220653
transform 1 0 2128 0 1 676
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5909_6
timestamp 1731220653
transform 1 0 2224 0 -1 780
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5908_6
timestamp 1731220653
transform 1 0 2112 0 -1 780
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5907_6
timestamp 1731220653
transform 1 0 2008 0 -1 780
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5906_6
timestamp 1731220653
transform 1 0 1912 0 -1 780
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5905_6
timestamp 1731220653
transform 1 0 2080 0 1 784
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5904_6
timestamp 1731220653
transform 1 0 1992 0 1 784
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5903_6
timestamp 1731220653
transform 1 0 1904 0 1 784
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5902_6
timestamp 1731220653
transform 1 0 1888 0 -1 892
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5901_6
timestamp 1731220653
transform 1 0 1784 0 -1 892
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5900_6
timestamp 1731220653
transform 1 0 2008 0 -1 892
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5899_6
timestamp 1731220653
transform 1 0 2272 0 -1 892
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5898_6
timestamp 1731220653
transform 1 0 2136 0 -1 892
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5897_6
timestamp 1731220653
transform 1 0 2104 0 1 896
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5896_6
timestamp 1731220653
transform 1 0 2008 0 1 896
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5895_6
timestamp 1731220653
transform 1 0 1912 0 1 896
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5894_6
timestamp 1731220653
transform 1 0 2192 0 1 896
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5893_6
timestamp 1731220653
transform 1 0 2272 0 1 896
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5892_6
timestamp 1731220653
transform 1 0 2352 0 1 896
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5891_6
timestamp 1731220653
transform 1 0 2360 0 -1 1012
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5890_6
timestamp 1731220653
transform 1 0 2264 0 -1 1012
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5889_6
timestamp 1731220653
transform 1 0 2168 0 -1 1012
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5888_6
timestamp 1731220653
transform 1 0 2064 0 -1 1012
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5887_6
timestamp 1731220653
transform 1 0 1944 0 -1 1012
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5886_6
timestamp 1731220653
transform 1 0 1816 0 -1 1012
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5885_6
timestamp 1731220653
transform 1 0 2344 0 1 1016
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5884_6
timestamp 1731220653
transform 1 0 2232 0 1 1016
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5883_6
timestamp 1731220653
transform 1 0 2128 0 1 1016
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5882_6
timestamp 1731220653
transform 1 0 2016 0 1 1016
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5881_6
timestamp 1731220653
transform 1 0 1904 0 1 1016
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5880_6
timestamp 1731220653
transform 1 0 2208 0 -1 1128
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5879_6
timestamp 1731220653
transform 1 0 2128 0 -1 1128
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5878_6
timestamp 1731220653
transform 1 0 2048 0 -1 1128
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5877_6
timestamp 1731220653
transform 1 0 1976 0 -1 1128
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5876_6
timestamp 1731220653
transform 1 0 1904 0 -1 1128
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5875_6
timestamp 1731220653
transform 1 0 1824 0 -1 1128
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5874_6
timestamp 1731220653
transform 1 0 1880 0 1 1128
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5873_6
timestamp 1731220653
transform 1 0 2008 0 1 1128
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5872_6
timestamp 1731220653
transform 1 0 2152 0 1 1128
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5871_6
timestamp 1731220653
transform 1 0 2304 0 1 1128
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5870_6
timestamp 1731220653
transform 1 0 2264 0 -1 1236
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5869_6
timestamp 1731220653
transform 1 0 2176 0 -1 1236
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5868_6
timestamp 1731220653
transform 1 0 2096 0 -1 1236
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5867_6
timestamp 1731220653
transform 1 0 2072 0 1 1240
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5866_6
timestamp 1731220653
transform 1 0 2184 0 1 1240
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5865_6
timestamp 1731220653
transform 1 0 2296 0 1 1240
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5864_6
timestamp 1731220653
transform 1 0 2216 0 -1 1344
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5863_6
timestamp 1731220653
transform 1 0 2136 0 -1 1344
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5862_6
timestamp 1731220653
transform 1 0 2056 0 -1 1344
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5861_6
timestamp 1731220653
transform 1 0 2296 0 -1 1344
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5860_6
timestamp 1731220653
transform 1 0 2296 0 1 1344
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5859_6
timestamp 1731220653
transform 1 0 2224 0 1 1344
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5858_6
timestamp 1731220653
transform 1 0 2152 0 1 1344
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5857_6
timestamp 1731220653
transform 1 0 2072 0 1 1344
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5856_6
timestamp 1731220653
transform 1 0 1984 0 1 1344
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5855_6
timestamp 1731220653
transform 1 0 2240 0 -1 1448
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5854_6
timestamp 1731220653
transform 1 0 2152 0 -1 1448
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5853_6
timestamp 1731220653
transform 1 0 2064 0 -1 1448
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5852_6
timestamp 1731220653
transform 1 0 1984 0 -1 1448
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5851_6
timestamp 1731220653
transform 1 0 1896 0 -1 1448
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5850_6
timestamp 1731220653
transform 1 0 1808 0 -1 1448
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5849_6
timestamp 1731220653
transform 1 0 2096 0 1 1456
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5848_6
timestamp 1731220653
transform 1 0 2008 0 1 1456
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5847_6
timestamp 1731220653
transform 1 0 1928 0 1 1456
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5846_6
timestamp 1731220653
transform 1 0 1848 0 1 1456
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5845_6
timestamp 1731220653
transform 1 0 1768 0 1 1456
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5844_6
timestamp 1731220653
transform 1 0 2000 0 -1 1560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5843_6
timestamp 1731220653
transform 1 0 1864 0 -1 1560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5842_6
timestamp 1731220653
transform 1 0 1728 0 -1 1560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5841_6
timestamp 1731220653
transform 1 0 1600 0 -1 1560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5840_6
timestamp 1731220653
transform 1 0 1464 0 -1 1560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5839_6
timestamp 1731220653
transform 1 0 1696 0 1 1560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5838_6
timestamp 1731220653
transform 1 0 1768 0 1 1560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5837_6
timestamp 1731220653
transform 1 0 1848 0 1 1560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5836_6
timestamp 1731220653
transform 1 0 2008 0 1 1560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5835_6
timestamp 1731220653
transform 1 0 1928 0 1 1560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5834_6
timestamp 1731220653
transform 1 0 1888 0 -1 1664
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5833_6
timestamp 1731220653
transform 1 0 1776 0 -1 1664
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5832_6
timestamp 1731220653
transform 1 0 2296 0 -1 1664
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5831_6
timestamp 1731220653
transform 1 0 2152 0 -1 1664
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5830_6
timestamp 1731220653
transform 1 0 2016 0 -1 1664
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5829_6
timestamp 1731220653
transform 1 0 1992 0 1 1668
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5828_6
timestamp 1731220653
transform 1 0 1896 0 1 1668
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5827_6
timestamp 1731220653
transform 1 0 2176 0 1 1668
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5826_6
timestamp 1731220653
transform 1 0 2088 0 1 1668
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5825_6
timestamp 1731220653
transform 1 0 2048 0 -1 1776
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5824_6
timestamp 1731220653
transform 1 0 1960 0 -1 1776
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5823_6
timestamp 1731220653
transform 1 0 2128 0 -1 1776
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5822_6
timestamp 1731220653
transform 1 0 2208 0 -1 1776
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5821_6
timestamp 1731220653
transform 1 0 2168 0 1 1776
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5820_6
timestamp 1731220653
transform 1 0 2312 0 1 1776
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5819_6
timestamp 1731220653
transform 1 0 2288 0 -1 1776
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5818_6
timestamp 1731220653
transform 1 0 2368 0 -1 1776
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5817_6
timestamp 1731220653
transform 1 0 2360 0 1 1668
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5816_6
timestamp 1731220653
transform 1 0 2264 0 1 1668
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5815_6
timestamp 1731220653
transform 1 0 2432 0 -1 1664
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5814_6
timestamp 1731220653
transform 1 0 2432 0 1 1668
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5813_6
timestamp 1731220653
transform 1 0 2432 0 -1 1776
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5812_6
timestamp 1731220653
transform 1 0 2432 0 1 1776
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5811_6
timestamp 1731220653
transform 1 0 2432 0 -1 1884
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5810_6
timestamp 1731220653
transform 1 0 2432 0 1 1888
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5809_6
timestamp 1731220653
transform 1 0 2352 0 1 1888
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5808_6
timestamp 1731220653
transform 1 0 2376 0 -1 1884
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5807_6
timestamp 1731220653
transform 1 0 2320 0 -1 1884
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5806_6
timestamp 1731220653
transform 1 0 2256 0 -1 1884
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5805_6
timestamp 1731220653
transform 1 0 2192 0 -1 1884
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5804_6
timestamp 1731220653
transform 1 0 2128 0 -1 1884
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5803_6
timestamp 1731220653
transform 1 0 2064 0 -1 1884
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5802_6
timestamp 1731220653
transform 1 0 2000 0 -1 1884
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5801_6
timestamp 1731220653
transform 1 0 2256 0 1 1888
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5800_6
timestamp 1731220653
transform 1 0 2160 0 1 1888
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5799_6
timestamp 1731220653
transform 1 0 2064 0 1 1888
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5798_6
timestamp 1731220653
transform 1 0 1976 0 1 1888
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5797_6
timestamp 1731220653
transform 1 0 1896 0 1 1888
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5796_6
timestamp 1731220653
transform 1 0 2024 0 -1 1996
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5795_6
timestamp 1731220653
transform 1 0 1952 0 -1 1996
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5794_6
timestamp 1731220653
transform 1 0 1888 0 -1 1996
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5793_6
timestamp 1731220653
transform 1 0 1824 0 -1 1996
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5792_6
timestamp 1731220653
transform 1 0 1760 0 -1 1996
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5791_6
timestamp 1731220653
transform 1 0 1728 0 1 2000
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5790_6
timestamp 1731220653
transform 1 0 1816 0 1 2000
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5789_6
timestamp 1731220653
transform 1 0 2096 0 1 2000
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5788_6
timestamp 1731220653
transform 1 0 2000 0 1 2000
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5787_6
timestamp 1731220653
transform 1 0 1904 0 1 2000
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5786_6
timestamp 1731220653
transform 1 0 1848 0 -1 2108
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5785_6
timestamp 1731220653
transform 1 0 1984 0 -1 2108
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5784_6
timestamp 1731220653
transform 1 0 2360 0 -1 2108
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5783_6
timestamp 1731220653
transform 1 0 2232 0 -1 2108
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5782_6
timestamp 1731220653
transform 1 0 2112 0 -1 2108
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5781_6
timestamp 1731220653
transform 1 0 1968 0 1 2108
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5780_6
timestamp 1731220653
transform 1 0 1792 0 1 2108
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5779_6
timestamp 1731220653
transform 1 0 2136 0 1 2108
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5778_6
timestamp 1731220653
transform 1 0 2296 0 1 2108
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5777_6
timestamp 1731220653
transform 1 0 2432 0 1 2108
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5776_6
timestamp 1731220653
transform 1 0 2432 0 -1 2232
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5775_6
timestamp 1731220653
transform 1 0 2376 0 -1 2232
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5774_6
timestamp 1731220653
transform 1 0 2312 0 -1 2232
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5773_6
timestamp 1731220653
transform 1 0 2248 0 -1 2232
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5772_6
timestamp 1731220653
transform 1 0 2184 0 -1 2232
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5771_6
timestamp 1731220653
transform 1 0 2120 0 -1 2232
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5770_6
timestamp 1731220653
transform 1 0 2048 0 -1 2232
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5769_6
timestamp 1731220653
transform 1 0 1976 0 -1 2232
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5768_6
timestamp 1731220653
transform 1 0 1896 0 -1 2232
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5767_6
timestamp 1731220653
transform 1 0 1808 0 -1 2232
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5766_6
timestamp 1731220653
transform 1 0 1712 0 -1 2232
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5765_6
timestamp 1731220653
transform 1 0 2216 0 1 2232
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5764_6
timestamp 1731220653
transform 1 0 2104 0 1 2232
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5763_6
timestamp 1731220653
transform 1 0 1992 0 1 2232
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5762_6
timestamp 1731220653
transform 1 0 1880 0 1 2232
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5761_6
timestamp 1731220653
transform 1 0 2136 0 -1 2336
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5760_6
timestamp 1731220653
transform 1 0 2056 0 -1 2336
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5759_6
timestamp 1731220653
transform 1 0 1976 0 -1 2336
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5758_6
timestamp 1731220653
transform 1 0 1896 0 -1 2336
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5757_6
timestamp 1731220653
transform 1 0 1824 0 -1 2336
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5756_6
timestamp 1731220653
transform 1 0 1832 0 1 2344
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5755_6
timestamp 1731220653
transform 1 0 1896 0 1 2344
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5754_6
timestamp 1731220653
transform 1 0 2088 0 1 2344
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5753_6
timestamp 1731220653
transform 1 0 2024 0 1 2344
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5752_6
timestamp 1731220653
transform 1 0 1960 0 1 2344
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5751_6
timestamp 1731220653
transform 1 0 1944 0 -1 2452
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5750_6
timestamp 1731220653
transform 1 0 1872 0 -1 2452
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5749_6
timestamp 1731220653
transform 1 0 2016 0 -1 2452
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5748_6
timestamp 1731220653
transform 1 0 2088 0 -1 2452
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5747_6
timestamp 1731220653
transform 1 0 2160 0 -1 2452
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5746_6
timestamp 1731220653
transform 1 0 2160 0 1 2456
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5745_6
timestamp 1731220653
transform 1 0 2088 0 1 2456
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5744_6
timestamp 1731220653
transform 1 0 2016 0 1 2456
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5743_6
timestamp 1731220653
transform 1 0 1944 0 1 2456
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5742_6
timestamp 1731220653
transform 1 0 1872 0 1 2456
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5741_6
timestamp 1731220653
transform 1 0 2160 0 -1 2560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5740_6
timestamp 1731220653
transform 1 0 2104 0 -1 2560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5739_6
timestamp 1731220653
transform 1 0 2048 0 -1 2560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5738_6
timestamp 1731220653
transform 1 0 1992 0 -1 2560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5737_6
timestamp 1731220653
transform 1 0 1936 0 -1 2560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5736_6
timestamp 1731220653
transform 1 0 1880 0 -1 2560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5735_6
timestamp 1731220653
transform 1 0 1824 0 -1 2560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5734_6
timestamp 1731220653
transform 1 0 1768 0 -1 2560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5733_6
timestamp 1731220653
transform 1 0 1712 0 -1 2560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5732_6
timestamp 1731220653
transform 1 0 1656 0 -1 2560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5731_6
timestamp 1731220653
transform 1 0 1600 0 -1 2560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5730_6
timestamp 1731220653
transform 1 0 1544 0 -1 2560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5729_6
timestamp 1731220653
transform 1 0 1488 0 -1 2560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5728_6
timestamp 1731220653
transform 1 0 1800 0 1 2456
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5727_6
timestamp 1731220653
transform 1 0 1728 0 1 2456
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5726_6
timestamp 1731220653
transform 1 0 1656 0 1 2456
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5725_6
timestamp 1731220653
transform 1 0 1584 0 1 2456
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5724_6
timestamp 1731220653
transform 1 0 1520 0 1 2456
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5723_6
timestamp 1731220653
transform 1 0 1536 0 -1 2452
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5722_6
timestamp 1731220653
transform 1 0 1600 0 -1 2452
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5721_6
timestamp 1731220653
transform 1 0 1664 0 -1 2452
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5720_6
timestamp 1731220653
transform 1 0 1736 0 -1 2452
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5719_6
timestamp 1731220653
transform 1 0 1808 0 -1 2452
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5718_6
timestamp 1731220653
transform 1 0 1768 0 1 2344
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5717_6
timestamp 1731220653
transform 1 0 1712 0 1 2344
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5716_6
timestamp 1731220653
transform 1 0 1656 0 1 2344
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5715_6
timestamp 1731220653
transform 1 0 1600 0 1 2344
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5714_6
timestamp 1731220653
transform 1 0 1544 0 1 2344
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5713_6
timestamp 1731220653
transform 1 0 1752 0 -1 2336
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5712_6
timestamp 1731220653
transform 1 0 1680 0 -1 2336
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5711_6
timestamp 1731220653
transform 1 0 1600 0 -1 2336
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5710_6
timestamp 1731220653
transform 1 0 1528 0 -1 2336
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5709_6
timestamp 1731220653
transform 1 0 1464 0 -1 2336
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5708_6
timestamp 1731220653
transform 1 0 1768 0 1 2232
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5707_6
timestamp 1731220653
transform 1 0 1664 0 1 2232
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5706_6
timestamp 1731220653
transform 1 0 1560 0 1 2232
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5705_6
timestamp 1731220653
transform 1 0 1456 0 1 2232
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5704_6
timestamp 1731220653
transform 1 0 1360 0 1 2232
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5703_6
timestamp 1731220653
transform 1 0 1360 0 -1 2232
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5702_6
timestamp 1731220653
transform 1 0 1600 0 -1 2232
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5701_6
timestamp 1731220653
transform 1 0 1480 0 -1 2232
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5700_6
timestamp 1731220653
transform 1 0 1384 0 1 2108
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5699_6
timestamp 1731220653
transform 1 0 1600 0 1 2108
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5698_6
timestamp 1731220653
transform 1 0 1704 0 -1 2108
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5697_6
timestamp 1731220653
transform 1 0 1544 0 -1 2108
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5696_6
timestamp 1731220653
transform 1 0 1376 0 -1 2108
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5695_6
timestamp 1731220653
transform 1 0 1424 0 1 2000
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5694_6
timestamp 1731220653
transform 1 0 1632 0 1 2000
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5693_6
timestamp 1731220653
transform 1 0 1528 0 1 2000
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5692_6
timestamp 1731220653
transform 1 0 1504 0 -1 1996
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5691_6
timestamp 1731220653
transform 1 0 1448 0 -1 1996
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5690_6
timestamp 1731220653
transform 1 0 1568 0 -1 1996
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5689_6
timestamp 1731220653
transform 1 0 1632 0 -1 1996
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5688_6
timestamp 1731220653
transform 1 0 1696 0 -1 1996
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5687_6
timestamp 1731220653
transform 1 0 1680 0 1 1888
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5686_6
timestamp 1731220653
transform 1 0 1608 0 1 1888
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5685_6
timestamp 1731220653
transform 1 0 1544 0 1 1888
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5684_6
timestamp 1731220653
transform 1 0 1824 0 1 1888
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5683_6
timestamp 1731220653
transform 1 0 1752 0 1 1888
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5682_6
timestamp 1731220653
transform 1 0 1720 0 -1 1884
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5681_6
timestamp 1731220653
transform 1 0 1656 0 -1 1884
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5680_6
timestamp 1731220653
transform 1 0 1600 0 -1 1884
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5679_6
timestamp 1731220653
transform 1 0 1792 0 -1 1884
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5678_6
timestamp 1731220653
transform 1 0 1864 0 -1 1884
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5677_6
timestamp 1731220653
transform 1 0 1936 0 -1 1884
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5676_6
timestamp 1731220653
transform 1 0 2032 0 1 1776
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5675_6
timestamp 1731220653
transform 1 0 1904 0 1 1776
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5674_6
timestamp 1731220653
transform 1 0 1792 0 1 1776
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5673_6
timestamp 1731220653
transform 1 0 1696 0 1 1776
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5672_6
timestamp 1731220653
transform 1 0 1608 0 1 1776
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5671_6
timestamp 1731220653
transform 1 0 1872 0 -1 1776
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5670_6
timestamp 1731220653
transform 1 0 1784 0 -1 1776
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5669_6
timestamp 1731220653
transform 1 0 1688 0 -1 1776
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5668_6
timestamp 1731220653
transform 1 0 1600 0 -1 1776
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5667_6
timestamp 1731220653
transform 1 0 1520 0 -1 1776
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5666_6
timestamp 1731220653
transform 1 0 1800 0 1 1668
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5665_6
timestamp 1731220653
transform 1 0 1704 0 1 1668
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5664_6
timestamp 1731220653
transform 1 0 1608 0 1 1668
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5663_6
timestamp 1731220653
transform 1 0 1520 0 1 1668
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5662_6
timestamp 1731220653
transform 1 0 1440 0 1 1668
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5661_6
timestamp 1731220653
transform 1 0 1376 0 1 1668
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5660_6
timestamp 1731220653
transform 1 0 1672 0 -1 1664
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5659_6
timestamp 1731220653
transform 1 0 1576 0 -1 1664
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5658_6
timestamp 1731220653
transform 1 0 1488 0 -1 1664
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5657_6
timestamp 1731220653
transform 1 0 1400 0 -1 1664
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5656_6
timestamp 1731220653
transform 1 0 1344 0 -1 1664
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5655_6
timestamp 1731220653
transform 1 0 1616 0 1 1560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5654_6
timestamp 1731220653
transform 1 0 1536 0 1 1560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5653_6
timestamp 1731220653
transform 1 0 1456 0 1 1560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5652_6
timestamp 1731220653
transform 1 0 1400 0 1 1560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5651_6
timestamp 1731220653
transform 1 0 1344 0 1 1560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5650_6
timestamp 1731220653
transform 1 0 1216 0 -1 1564
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5649_6
timestamp 1731220653
transform 1 0 1160 0 -1 1564
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5648_6
timestamp 1731220653
transform 1 0 1080 0 -1 1564
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5647_6
timestamp 1731220653
transform 1 0 1344 0 -1 1560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5646_6
timestamp 1731220653
transform 1 0 1344 0 1 1456
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5645_6
timestamp 1731220653
transform 1 0 1400 0 1 1456
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5644_6
timestamp 1731220653
transform 1 0 1456 0 1 1456
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5643_6
timestamp 1731220653
transform 1 0 1688 0 1 1456
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5642_6
timestamp 1731220653
transform 1 0 1608 0 1 1456
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5641_6
timestamp 1731220653
transform 1 0 1528 0 1 1456
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5640_6
timestamp 1731220653
transform 1 0 1528 0 -1 1448
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5639_6
timestamp 1731220653
transform 1 0 1440 0 -1 1448
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5638_6
timestamp 1731220653
transform 1 0 1352 0 -1 1448
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5637_6
timestamp 1731220653
transform 1 0 1624 0 -1 1448
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5636_6
timestamp 1731220653
transform 1 0 1720 0 -1 1448
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5635_6
timestamp 1731220653
transform 1 0 1712 0 1 1344
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5634_6
timestamp 1731220653
transform 1 0 1624 0 1 1344
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5633_6
timestamp 1731220653
transform 1 0 1544 0 1 1344
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5632_6
timestamp 1731220653
transform 1 0 1808 0 1 1344
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5631_6
timestamp 1731220653
transform 1 0 1896 0 1 1344
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5630_6
timestamp 1731220653
transform 1 0 1888 0 -1 1344
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5629_6
timestamp 1731220653
transform 1 0 1800 0 -1 1344
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5628_6
timestamp 1731220653
transform 1 0 1976 0 -1 1344
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5627_6
timestamp 1731220653
transform 1 0 1968 0 1 1240
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5626_6
timestamp 1731220653
transform 1 0 2024 0 -1 1236
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5625_6
timestamp 1731220653
transform 1 0 1960 0 -1 1236
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5624_6
timestamp 1731220653
transform 1 0 1904 0 -1 1236
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5623_6
timestamp 1731220653
transform 1 0 1848 0 -1 1236
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5622_6
timestamp 1731220653
transform 1 0 1792 0 -1 1236
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5621_6
timestamp 1731220653
transform 1 0 1736 0 -1 1236
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5620_6
timestamp 1731220653
transform 1 0 1680 0 -1 1236
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5619_6
timestamp 1731220653
transform 1 0 1624 0 -1 1236
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5618_6
timestamp 1731220653
transform 1 0 1688 0 1 1240
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5617_6
timestamp 1731220653
transform 1 0 1872 0 1 1240
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5616_6
timestamp 1731220653
transform 1 0 1776 0 1 1240
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5615_6
timestamp 1731220653
transform 1 0 1720 0 -1 1344
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5614_6
timestamp 1731220653
transform 1 0 1640 0 -1 1344
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5613_6
timestamp 1731220653
transform 1 0 1576 0 -1 1344
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5612_6
timestamp 1731220653
transform 1 0 1544 0 1 1240
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5611_6
timestamp 1731220653
transform 1 0 1608 0 1 1240
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5610_6
timestamp 1731220653
transform 1 0 1568 0 -1 1236
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5609_6
timestamp 1731220653
transform 1 0 1512 0 -1 1236
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5608_6
timestamp 1731220653
transform 1 0 1768 0 1 1128
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5607_6
timestamp 1731220653
transform 1 0 1680 0 1 1128
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5606_6
timestamp 1731220653
transform 1 0 1608 0 1 1128
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5605_6
timestamp 1731220653
transform 1 0 1544 0 1 1128
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5604_6
timestamp 1731220653
transform 1 0 1744 0 -1 1128
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5603_6
timestamp 1731220653
transform 1 0 1664 0 -1 1128
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5602_6
timestamp 1731220653
transform 1 0 1584 0 -1 1128
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5601_6
timestamp 1731220653
transform 1 0 1512 0 -1 1128
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5600_6
timestamp 1731220653
transform 1 0 1440 0 -1 1128
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5599_6
timestamp 1731220653
transform 1 0 1376 0 -1 1128
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5598_6
timestamp 1731220653
transform 1 0 1792 0 1 1016
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5597_6
timestamp 1731220653
transform 1 0 1672 0 1 1016
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5596_6
timestamp 1731220653
transform 1 0 1552 0 1 1016
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5595_6
timestamp 1731220653
transform 1 0 1432 0 1 1016
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5594_6
timestamp 1731220653
transform 1 0 1344 0 1 1016
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5593_6
timestamp 1731220653
transform 1 0 1672 0 -1 1012
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5592_6
timestamp 1731220653
transform 1 0 1504 0 -1 1012
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5591_6
timestamp 1731220653
transform 1 0 1216 0 1 980
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5590_6
timestamp 1731220653
transform 1 0 1160 0 1 980
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5589_6
timestamp 1731220653
transform 1 0 1080 0 1 980
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5588_6
timestamp 1731220653
transform 1 0 1000 0 -1 980
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5587_6
timestamp 1731220653
transform 1 0 920 0 -1 980
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5586_6
timestamp 1731220653
transform 1 0 832 0 -1 980
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5585_6
timestamp 1731220653
transform 1 0 744 0 -1 980
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5584_6
timestamp 1731220653
transform 1 0 1080 0 -1 980
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5583_6
timestamp 1731220653
transform 1 0 1160 0 -1 980
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5582_6
timestamp 1731220653
transform 1 0 1160 0 1 868
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5581_6
timestamp 1731220653
transform 1 0 1064 0 1 868
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5580_6
timestamp 1731220653
transform 1 0 968 0 1 868
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5579_6
timestamp 1731220653
transform 1 0 880 0 1 868
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5578_6
timestamp 1731220653
transform 1 0 784 0 1 868
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5577_6
timestamp 1731220653
transform 1 0 896 0 -1 864
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5576_6
timestamp 1731220653
transform 1 0 824 0 -1 864
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5575_6
timestamp 1731220653
transform 1 0 752 0 -1 864
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5574_6
timestamp 1731220653
transform 1 0 688 0 -1 864
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5573_6
timestamp 1731220653
transform 1 0 624 0 -1 864
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5572_6
timestamp 1731220653
transform 1 0 680 0 1 756
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5571_6
timestamp 1731220653
transform 1 0 608 0 1 756
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5570_6
timestamp 1731220653
transform 1 0 536 0 1 756
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5569_6
timestamp 1731220653
transform 1 0 456 0 1 756
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5568_6
timestamp 1731220653
transform 1 0 368 0 1 756
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5567_6
timestamp 1731220653
transform 1 0 560 0 -1 864
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5566_6
timestamp 1731220653
transform 1 0 496 0 -1 864
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5565_6
timestamp 1731220653
transform 1 0 432 0 -1 864
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5564_6
timestamp 1731220653
transform 1 0 368 0 -1 864
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5563_6
timestamp 1731220653
transform 1 0 688 0 1 868
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5562_6
timestamp 1731220653
transform 1 0 592 0 1 868
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5561_6
timestamp 1731220653
transform 1 0 496 0 1 868
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5560_6
timestamp 1731220653
transform 1 0 400 0 1 868
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5559_6
timestamp 1731220653
transform 1 0 448 0 -1 980
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5558_6
timestamp 1731220653
transform 1 0 352 0 -1 980
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5557_6
timestamp 1731220653
transform 1 0 264 0 -1 980
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5556_6
timestamp 1731220653
transform 1 0 272 0 1 980
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5555_6
timestamp 1731220653
transform 1 0 360 0 1 980
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5554_6
timestamp 1731220653
transform 1 0 456 0 1 980
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5553_6
timestamp 1731220653
transform 1 0 440 0 -1 1092
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5552_6
timestamp 1731220653
transform 1 0 352 0 -1 1092
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5551_6
timestamp 1731220653
transform 1 0 272 0 -1 1092
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5550_6
timestamp 1731220653
transform 1 0 200 0 -1 1092
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5549_6
timestamp 1731220653
transform 1 0 160 0 1 1100
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5548_6
timestamp 1731220653
transform 1 0 256 0 1 1100
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5547_6
timestamp 1731220653
transform 1 0 352 0 1 1100
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5546_6
timestamp 1731220653
transform 1 0 344 0 -1 1208
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5545_6
timestamp 1731220653
transform 1 0 264 0 -1 1208
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5544_6
timestamp 1731220653
transform 1 0 184 0 -1 1208
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5543_6
timestamp 1731220653
transform 1 0 128 0 -1 1208
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5542_6
timestamp 1731220653
transform 1 0 368 0 1 1212
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5541_6
timestamp 1731220653
transform 1 0 280 0 1 1212
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5540_6
timestamp 1731220653
transform 1 0 192 0 1 1212
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5539_6
timestamp 1731220653
transform 1 0 128 0 1 1212
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5538_6
timestamp 1731220653
transform 1 0 128 0 -1 1324
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5537_6
timestamp 1731220653
transform 1 0 360 0 -1 1324
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5536_6
timestamp 1731220653
transform 1 0 232 0 -1 1324
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5535_6
timestamp 1731220653
transform 1 0 200 0 1 1340
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5534_6
timestamp 1731220653
transform 1 0 128 0 1 1340
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5533_6
timestamp 1731220653
transform 1 0 184 0 -1 1448
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5532_6
timestamp 1731220653
transform 1 0 248 0 -1 1448
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5531_6
timestamp 1731220653
transform 1 0 256 0 1 1452
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5530_6
timestamp 1731220653
transform 1 0 240 0 -1 1564
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5529_6
timestamp 1731220653
transform 1 0 488 0 1 1564
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5528_6
timestamp 1731220653
transform 1 0 576 0 1 1564
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5527_6
timestamp 1731220653
transform 1 0 568 0 -1 1672
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5526_6
timestamp 1731220653
transform 1 0 584 0 1 1676
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5525_6
timestamp 1731220653
transform 1 0 496 0 -1 1784
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5524_6
timestamp 1731220653
transform 1 0 600 0 -1 1784
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5523_6
timestamp 1731220653
transform 1 0 568 0 1 1796
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5522_6
timestamp 1731220653
transform 1 0 536 0 -1 1900
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5521_6
timestamp 1731220653
transform 1 0 624 0 -1 1900
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5520_6
timestamp 1731220653
transform 1 0 720 0 1 1908
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5519_6
timestamp 1731220653
transform 1 0 896 0 1 1908
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5518_6
timestamp 1731220653
transform 1 0 840 0 -1 2016
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5517_6
timestamp 1731220653
transform 1 0 728 0 -1 2016
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5516_6
timestamp 1731220653
transform 1 0 688 0 1 2020
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5515_6
timestamp 1731220653
transform 1 0 768 0 1 2020
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5514_6
timestamp 1731220653
transform 1 0 920 0 1 2020
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5513_6
timestamp 1731220653
transform 1 0 840 0 1 2020
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5512_6
timestamp 1731220653
transform 1 0 792 0 -1 2128
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5511_6
timestamp 1731220653
transform 1 0 704 0 -1 2128
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5510_6
timestamp 1731220653
transform 1 0 880 0 -1 2128
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5509_6
timestamp 1731220653
transform 1 0 968 0 -1 2128
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5508_6
timestamp 1731220653
transform 1 0 936 0 1 2128
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5507_6
timestamp 1731220653
transform 1 0 840 0 1 2128
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5506_6
timestamp 1731220653
transform 1 0 744 0 1 2128
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5505_6
timestamp 1731220653
transform 1 0 640 0 1 2128
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5504_6
timestamp 1731220653
transform 1 0 616 0 -1 2232
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5503_6
timestamp 1731220653
transform 1 0 720 0 -1 2232
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5502_6
timestamp 1731220653
transform 1 0 824 0 -1 2232
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5501_6
timestamp 1731220653
transform 1 0 928 0 -1 2232
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5500_6
timestamp 1731220653
transform 1 0 888 0 1 2232
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5499_6
timestamp 1731220653
transform 1 0 784 0 1 2232
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5498_6
timestamp 1731220653
transform 1 0 680 0 1 2232
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5497_6
timestamp 1731220653
transform 1 0 672 0 -1 2344
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5496_6
timestamp 1731220653
transform 1 0 600 0 -1 2344
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5495_6
timestamp 1731220653
transform 1 0 736 0 -1 2344
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5494_6
timestamp 1731220653
transform 1 0 800 0 -1 2344
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5493_6
timestamp 1731220653
transform 1 0 856 0 -1 2344
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5492_6
timestamp 1731220653
transform 1 0 920 0 -1 2344
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5491_6
timestamp 1731220653
transform 1 0 984 0 -1 2344
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5490_6
timestamp 1731220653
transform 1 0 1048 0 -1 2344
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5489_6
timestamp 1731220653
transform 1 0 1104 0 -1 2344
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5488_6
timestamp 1731220653
transform 1 0 1160 0 -1 2344
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5487_6
timestamp 1731220653
transform 1 0 1216 0 -1 2344
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5486_6
timestamp 1731220653
transform 1 0 1216 0 1 2232
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5485_6
timestamp 1731220653
transform 1 0 1104 0 1 2232
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5484_6
timestamp 1731220653
transform 1 0 992 0 1 2232
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5483_6
timestamp 1731220653
transform 1 0 1032 0 -1 2232
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5482_6
timestamp 1731220653
transform 1 0 1216 0 -1 2232
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5481_6
timestamp 1731220653
transform 1 0 1136 0 -1 2232
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5480_6
timestamp 1731220653
transform 1 0 1032 0 1 2128
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5479_6
timestamp 1731220653
transform 1 0 1136 0 1 2128
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5478_6
timestamp 1731220653
transform 1 0 1216 0 1 2128
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5477_6
timestamp 1731220653
transform 1 0 1216 0 -1 2128
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5476_6
timestamp 1731220653
transform 1 0 1144 0 -1 2128
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5475_6
timestamp 1731220653
transform 1 0 1056 0 -1 2128
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5474_6
timestamp 1731220653
transform 1 0 1216 0 1 2020
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5473_6
timestamp 1731220653
transform 1 0 1160 0 1 2020
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5472_6
timestamp 1731220653
transform 1 0 1080 0 1 2020
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5471_6
timestamp 1731220653
transform 1 0 1000 0 1 2020
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5470_6
timestamp 1731220653
transform 1 0 952 0 -1 2016
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5469_6
timestamp 1731220653
transform 1 0 1192 0 -1 2016
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5468_6
timestamp 1731220653
transform 1 0 1072 0 -1 2016
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5467_6
timestamp 1731220653
transform 1 0 1072 0 1 1908
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5466_6
timestamp 1731220653
transform 1 0 1008 0 -1 1900
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5465_6
timestamp 1731220653
transform 1 0 904 0 1 1796
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5464_6
timestamp 1731220653
transform 1 0 880 0 -1 1784
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5463_6
timestamp 1731220653
transform 1 0 912 0 1 1676
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5462_6
timestamp 1731220653
transform 1 0 856 0 -1 1672
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5461_6
timestamp 1731220653
transform 1 0 872 0 1 1564
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5460_6
timestamp 1731220653
transform 1 0 752 0 -1 1564
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5459_6
timestamp 1731220653
transform 1 0 712 0 1 1452
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5458_6
timestamp 1731220653
transform 1 0 792 0 1 1452
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5457_6
timestamp 1731220653
transform 1 0 808 0 -1 1448
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5456_6
timestamp 1731220653
transform 1 0 816 0 1 1340
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5455_6
timestamp 1731220653
transform 1 0 728 0 1 1340
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5454_6
timestamp 1731220653
transform 1 0 576 0 -1 1324
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5453_6
timestamp 1731220653
transform 1 0 472 0 -1 1324
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5452_6
timestamp 1731220653
transform 1 0 528 0 1 1212
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5451_6
timestamp 1731220653
transform 1 0 448 0 1 1212
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5450_6
timestamp 1731220653
transform 1 0 424 0 -1 1208
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5449_6
timestamp 1731220653
transform 1 0 504 0 -1 1208
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5448_6
timestamp 1731220653
transform 1 0 448 0 1 1100
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5447_6
timestamp 1731220653
transform 1 0 544 0 1 1100
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5446_6
timestamp 1731220653
transform 1 0 536 0 -1 1092
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5445_6
timestamp 1731220653
transform 1 0 632 0 -1 1092
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5444_6
timestamp 1731220653
transform 1 0 552 0 1 980
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5443_6
timestamp 1731220653
transform 1 0 648 0 1 980
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5442_6
timestamp 1731220653
transform 1 0 648 0 -1 980
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5441_6
timestamp 1731220653
transform 1 0 544 0 -1 980
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5440_6
timestamp 1731220653
transform 1 0 320 0 1 868
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5439_6
timestamp 1731220653
transform 1 0 248 0 1 868
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5438_6
timestamp 1731220653
transform 1 0 240 0 -1 864
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5437_6
timestamp 1731220653
transform 1 0 304 0 -1 864
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5436_6
timestamp 1731220653
transform 1 0 280 0 1 756
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5435_6
timestamp 1731220653
transform 1 0 192 0 1 756
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5434_6
timestamp 1731220653
transform 1 0 128 0 -1 756
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5433_6
timestamp 1731220653
transform 1 0 248 0 -1 756
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5432_6
timestamp 1731220653
transform 1 0 384 0 -1 756
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5431_6
timestamp 1731220653
transform 1 0 480 0 1 652
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5430_6
timestamp 1731220653
transform 1 0 368 0 1 652
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5429_6
timestamp 1731220653
transform 1 0 272 0 1 652
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5428_6
timestamp 1731220653
transform 1 0 184 0 1 652
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5427_6
timestamp 1731220653
transform 1 0 128 0 1 652
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5426_6
timestamp 1731220653
transform 1 0 256 0 -1 648
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5425_6
timestamp 1731220653
transform 1 0 144 0 -1 648
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5424_6
timestamp 1731220653
transform 1 0 128 0 1 544
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5423_6
timestamp 1731220653
transform 1 0 216 0 1 544
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5422_6
timestamp 1731220653
transform 1 0 312 0 1 544
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5421_6
timestamp 1731220653
transform 1 0 232 0 -1 536
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5420_6
timestamp 1731220653
transform 1 0 136 0 -1 536
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5419_6
timestamp 1731220653
transform 1 0 128 0 1 428
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5418_6
timestamp 1731220653
transform 1 0 184 0 1 428
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5417_6
timestamp 1731220653
transform 1 0 272 0 -1 428
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5416_6
timestamp 1731220653
transform 1 0 184 0 -1 428
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5415_6
timestamp 1731220653
transform 1 0 128 0 -1 428
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5414_6
timestamp 1731220653
transform 1 0 128 0 1 320
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5413_6
timestamp 1731220653
transform 1 0 208 0 1 320
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5412_6
timestamp 1731220653
transform 1 0 208 0 -1 316
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5411_6
timestamp 1731220653
transform 1 0 128 0 -1 316
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5410_6
timestamp 1731220653
transform 1 0 128 0 1 212
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5409_6
timestamp 1731220653
transform 1 0 200 0 1 212
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5408_6
timestamp 1731220653
transform 1 0 296 0 1 212
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5407_6
timestamp 1731220653
transform 1 0 272 0 -1 208
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5406_6
timestamp 1731220653
transform 1 0 176 0 -1 208
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5405_6
timestamp 1731220653
transform 1 0 184 0 1 96
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5404_6
timestamp 1731220653
transform 1 0 128 0 1 96
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5403_6
timestamp 1731220653
transform 1 0 240 0 1 96
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5402_6
timestamp 1731220653
transform 1 0 296 0 1 96
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5401_6
timestamp 1731220653
transform 1 0 352 0 1 96
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5400_6
timestamp 1731220653
transform 1 0 408 0 1 96
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5399_6
timestamp 1731220653
transform 1 0 576 0 1 96
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5398_6
timestamp 1731220653
transform 1 0 520 0 1 96
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5397_6
timestamp 1731220653
transform 1 0 464 0 1 96
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5396_6
timestamp 1731220653
transform 1 0 376 0 -1 208
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5395_6
timestamp 1731220653
transform 1 0 480 0 -1 208
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5394_6
timestamp 1731220653
transform 1 0 584 0 -1 208
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5393_6
timestamp 1731220653
transform 1 0 624 0 1 212
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5392_6
timestamp 1731220653
transform 1 0 512 0 1 212
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5391_6
timestamp 1731220653
transform 1 0 400 0 1 212
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5390_6
timestamp 1731220653
transform 1 0 312 0 -1 316
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5389_6
timestamp 1731220653
transform 1 0 416 0 -1 316
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5388_6
timestamp 1731220653
transform 1 0 528 0 -1 316
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5387_6
timestamp 1731220653
transform 1 0 520 0 1 320
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5386_6
timestamp 1731220653
transform 1 0 416 0 1 320
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5385_6
timestamp 1731220653
transform 1 0 312 0 1 320
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5384_6
timestamp 1731220653
transform 1 0 600 0 -1 428
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5383_6
timestamp 1731220653
transform 1 0 488 0 -1 428
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5382_6
timestamp 1731220653
transform 1 0 376 0 -1 428
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5381_6
timestamp 1731220653
transform 1 0 352 0 1 428
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5380_6
timestamp 1731220653
transform 1 0 264 0 1 428
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5379_6
timestamp 1731220653
transform 1 0 536 0 1 428
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5378_6
timestamp 1731220653
transform 1 0 440 0 1 428
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5377_6
timestamp 1731220653
transform 1 0 424 0 -1 536
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5376_6
timestamp 1731220653
transform 1 0 328 0 -1 536
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5375_6
timestamp 1731220653
transform 1 0 520 0 -1 536
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5374_6
timestamp 1731220653
transform 1 0 608 0 1 544
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5373_6
timestamp 1731220653
transform 1 0 512 0 1 544
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5372_6
timestamp 1731220653
transform 1 0 408 0 1 544
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5371_6
timestamp 1731220653
transform 1 0 360 0 -1 648
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5370_6
timestamp 1731220653
transform 1 0 456 0 -1 648
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5369_6
timestamp 1731220653
transform 1 0 552 0 -1 648
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5368_6
timestamp 1731220653
transform 1 0 648 0 -1 648
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5367_6
timestamp 1731220653
transform 1 0 600 0 1 652
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5366_6
timestamp 1731220653
transform 1 0 720 0 1 652
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5365_6
timestamp 1731220653
transform 1 0 640 0 -1 756
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5364_6
timestamp 1731220653
transform 1 0 512 0 -1 756
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5363_6
timestamp 1731220653
transform 1 0 768 0 -1 756
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5362_6
timestamp 1731220653
transform 1 0 744 0 1 756
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5361_6
timestamp 1731220653
transform 1 0 808 0 1 756
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5360_6
timestamp 1731220653
transform 1 0 872 0 1 756
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5359_6
timestamp 1731220653
transform 1 0 944 0 1 756
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5358_6
timestamp 1731220653
transform 1 0 1016 0 1 756
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5357_6
timestamp 1731220653
transform 1 0 1032 0 -1 756
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5356_6
timestamp 1731220653
transform 1 0 896 0 -1 756
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5355_6
timestamp 1731220653
transform 1 0 848 0 1 652
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5354_6
timestamp 1731220653
transform 1 0 976 0 1 652
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5353_6
timestamp 1731220653
transform 1 0 936 0 -1 648
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5352_6
timestamp 1731220653
transform 1 0 840 0 -1 648
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5351_6
timestamp 1731220653
transform 1 0 744 0 -1 648
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5350_6
timestamp 1731220653
transform 1 0 800 0 1 544
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5349_6
timestamp 1731220653
transform 1 0 704 0 1 544
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5348_6
timestamp 1731220653
transform 1 0 704 0 -1 536
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5347_6
timestamp 1731220653
transform 1 0 616 0 -1 536
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5346_6
timestamp 1731220653
transform 1 0 632 0 1 428
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5345_6
timestamp 1731220653
transform 1 0 728 0 1 428
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5344_6
timestamp 1731220653
transform 1 0 712 0 -1 428
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5343_6
timestamp 1731220653
transform 1 0 728 0 1 320
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5342_6
timestamp 1731220653
transform 1 0 624 0 1 320
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5341_6
timestamp 1731220653
transform 1 0 632 0 -1 316
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5340_6
timestamp 1731220653
transform 1 0 736 0 -1 316
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5339_6
timestamp 1731220653
transform 1 0 840 0 -1 316
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5338_6
timestamp 1731220653
transform 1 0 848 0 1 212
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5337_6
timestamp 1731220653
transform 1 0 736 0 1 212
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5336_6
timestamp 1731220653
transform 1 0 688 0 -1 208
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5335_6
timestamp 1731220653
transform 1 0 792 0 -1 208
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5334_6
timestamp 1731220653
transform 1 0 744 0 1 96
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5333_6
timestamp 1731220653
transform 1 0 688 0 1 96
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5332_6
timestamp 1731220653
transform 1 0 632 0 1 96
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5331_6
timestamp 1731220653
transform 1 0 808 0 1 96
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5330_6
timestamp 1731220653
transform 1 0 872 0 1 96
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5329_6
timestamp 1731220653
transform 1 0 936 0 1 96
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5328_6
timestamp 1731220653
transform 1 0 1000 0 1 96
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5327_6
timestamp 1731220653
transform 1 0 1064 0 1 96
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5326_6
timestamp 1731220653
transform 1 0 1128 0 1 96
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5325_6
timestamp 1731220653
transform 1 0 1096 0 -1 208
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5324_6
timestamp 1731220653
transform 1 0 992 0 -1 208
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5323_6
timestamp 1731220653
transform 1 0 888 0 -1 208
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5322_6
timestamp 1731220653
transform 1 0 960 0 1 212
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5321_6
timestamp 1731220653
transform 1 0 1080 0 1 212
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5320_6
timestamp 1731220653
transform 1 0 1200 0 1 212
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5319_6
timestamp 1731220653
transform 1 0 1136 0 -1 316
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5318_6
timestamp 1731220653
transform 1 0 1032 0 -1 316
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5317_6
timestamp 1731220653
transform 1 0 936 0 -1 316
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5316_6
timestamp 1731220653
transform 1 0 912 0 1 320
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5315_6
timestamp 1731220653
transform 1 0 824 0 1 320
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5314_6
timestamp 1731220653
transform 1 0 992 0 1 320
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5313_6
timestamp 1731220653
transform 1 0 928 0 -1 428
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5312_6
timestamp 1731220653
transform 1 0 824 0 -1 428
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5311_6
timestamp 1731220653
transform 1 0 1032 0 1 428
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5310_6
timestamp 1731220653
transform 1 0 928 0 1 428
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5309_6
timestamp 1731220653
transform 1 0 824 0 1 428
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5308_6
timestamp 1731220653
transform 1 0 784 0 -1 536
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5307_6
timestamp 1731220653
transform 1 0 864 0 -1 536
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5306_6
timestamp 1731220653
transform 1 0 1024 0 -1 536
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5305_6
timestamp 1731220653
transform 1 0 944 0 -1 536
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5304_6
timestamp 1731220653
transform 1 0 888 0 1 544
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5303_6
timestamp 1731220653
transform 1 0 976 0 1 544
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5302_6
timestamp 1731220653
transform 1 0 1064 0 1 544
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5301_6
timestamp 1731220653
transform 1 0 1160 0 1 544
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5300_6
timestamp 1731220653
transform 1 0 1136 0 -1 648
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5299_6
timestamp 1731220653
transform 1 0 1032 0 -1 648
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5298_6
timestamp 1731220653
transform 1 0 1216 0 -1 648
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5297_6
timestamp 1731220653
transform 1 0 1600 0 -1 664
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5296_6
timestamp 1731220653
transform 1 0 1704 0 -1 664
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5295_6
timestamp 1731220653
transform 1 0 1720 0 1 560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5294_6
timestamp 1731220653
transform 1 0 1624 0 1 560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5293_6
timestamp 1731220653
transform 1 0 1528 0 1 560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5292_6
timestamp 1731220653
transform 1 0 1544 0 -1 560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5291_6
timestamp 1731220653
transform 1 0 1640 0 -1 560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5290_6
timestamp 1731220653
transform 1 0 1744 0 -1 560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5289_6
timestamp 1731220653
transform 1 0 1784 0 1 452
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5288_6
timestamp 1731220653
transform 1 0 1672 0 1 452
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5287_6
timestamp 1731220653
transform 1 0 1552 0 1 452
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5286_6
timestamp 1731220653
transform 1 0 1576 0 -1 440
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5285_6
timestamp 1731220653
transform 1 0 1632 0 -1 440
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5284_6
timestamp 1731220653
transform 1 0 1688 0 -1 440
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5283_6
timestamp 1731220653
transform 1 0 1752 0 -1 440
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5282_6
timestamp 1731220653
transform 1 0 1824 0 -1 440
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5281_6
timestamp 1731220653
transform 1 0 2000 0 1 332
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5280_6
timestamp 1731220653
transform 1 0 2088 0 1 332
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5279_6
timestamp 1731220653
transform 1 0 2072 0 -1 440
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5278_6
timestamp 1731220653
transform 1 0 1984 0 -1 440
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5277_6
timestamp 1731220653
transform 1 0 1904 0 -1 440
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5276_6
timestamp 1731220653
transform 1 0 1848 0 1 332
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5275_6
timestamp 1731220653
transform 1 0 1776 0 1 332
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5274_6
timestamp 1731220653
transform 1 0 1712 0 1 332
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5273_6
timestamp 1731220653
transform 1 0 1656 0 1 332
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5272_6
timestamp 1731220653
transform 1 0 1576 0 -1 324
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5271_6
timestamp 1731220653
transform 1 0 1448 0 -1 324
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5270_6
timestamp 1731220653
transform 1 0 1704 0 -1 324
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5269_6
timestamp 1731220653
transform 1 0 1736 0 1 212
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5268_6
timestamp 1731220653
transform 1 0 1632 0 1 212
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5267_6
timestamp 1731220653
transform 1 0 1528 0 1 212
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5266_6
timestamp 1731220653
transform 1 0 1544 0 -1 208
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5265_6
timestamp 1731220653
transform 1 0 1632 0 -1 208
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5264_6
timestamp 1731220653
transform 1 0 1712 0 -1 208
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5263_6
timestamp 1731220653
transform 1 0 1736 0 1 84
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5262_6
timestamp 1731220653
transform 1 0 1680 0 1 84
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5261_6
timestamp 1731220653
transform 1 0 1624 0 1 84
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5260_6
timestamp 1731220653
transform 1 0 1568 0 1 84
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5259_6
timestamp 1731220653
transform 1 0 1512 0 1 84
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5258_6
timestamp 1731220653
transform 1 0 1456 0 1 84
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5257_6
timestamp 1731220653
transform 1 0 1400 0 1 84
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5256_6
timestamp 1731220653
transform 1 0 1344 0 1 84
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5255_6
timestamp 1731220653
transform 1 0 1344 0 -1 208
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5254_6
timestamp 1731220653
transform 1 0 1400 0 -1 208
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5253_6
timestamp 1731220653
transform 1 0 1464 0 -1 208
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5252_6
timestamp 1731220653
transform 1 0 1424 0 1 212
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5251_6
timestamp 1731220653
transform 1 0 1344 0 1 212
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5250_6
timestamp 1731220653
transform 1 0 1344 0 -1 324
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5249_6
timestamp 1731220653
transform 1 0 1216 0 -1 316
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5248_6
timestamp 1731220653
transform 1 0 1216 0 1 320
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5247_6
timestamp 1731220653
transform 1 0 1152 0 1 320
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5246_6
timestamp 1731220653
transform 1 0 1072 0 1 320
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5245_6
timestamp 1731220653
transform 1 0 1032 0 -1 428
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5244_6
timestamp 1731220653
transform 1 0 1216 0 -1 428
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5243_6
timestamp 1731220653
transform 1 0 1136 0 -1 428
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5242_6
timestamp 1731220653
transform 1 0 1136 0 1 428
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5241_6
timestamp 1731220653
transform 1 0 1216 0 1 428
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5240_6
timestamp 1731220653
transform 1 0 1344 0 1 452
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5239_6
timestamp 1731220653
transform 1 0 1432 0 1 452
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5238_6
timestamp 1731220653
transform 1 0 1448 0 -1 560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5237_6
timestamp 1731220653
transform 1 0 1368 0 -1 560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5236_6
timestamp 1731220653
transform 1 0 1360 0 1 560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5235_6
timestamp 1731220653
transform 1 0 1440 0 1 560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5234_6
timestamp 1731220653
transform 1 0 1504 0 -1 664
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5233_6
timestamp 1731220653
transform 1 0 1408 0 -1 664
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5232_6
timestamp 1731220653
transform 1 0 1344 0 -1 664
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5231_6
timestamp 1731220653
transform 1 0 1216 0 1 652
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5230_6
timestamp 1731220653
transform 1 0 1104 0 1 652
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5229_6
timestamp 1731220653
transform 1 0 1344 0 1 676
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5228_6
timestamp 1731220653
transform 1 0 1408 0 1 676
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5227_6
timestamp 1731220653
transform 1 0 1504 0 1 676
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5226_6
timestamp 1731220653
transform 1 0 1608 0 1 676
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5225_6
timestamp 1731220653
transform 1 0 1712 0 1 676
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5224_6
timestamp 1731220653
transform 1 0 1680 0 -1 780
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5223_6
timestamp 1731220653
transform 1 0 1616 0 -1 780
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5222_6
timestamp 1731220653
transform 1 0 1560 0 -1 780
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5221_6
timestamp 1731220653
transform 1 0 1752 0 -1 780
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5220_6
timestamp 1731220653
transform 1 0 1824 0 -1 780
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5219_6
timestamp 1731220653
transform 1 0 1824 0 1 784
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5218_6
timestamp 1731220653
transform 1 0 1744 0 1 784
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5217_6
timestamp 1731220653
transform 1 0 1680 0 1 784
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5216_6
timestamp 1731220653
transform 1 0 1624 0 1 784
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5215_6
timestamp 1731220653
transform 1 0 1568 0 1 784
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5214_6
timestamp 1731220653
transform 1 0 1696 0 -1 892
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5213_6
timestamp 1731220653
transform 1 0 1616 0 -1 892
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5212_6
timestamp 1731220653
transform 1 0 1544 0 -1 892
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5211_6
timestamp 1731220653
transform 1 0 1480 0 -1 892
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5210_6
timestamp 1731220653
transform 1 0 1424 0 -1 892
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5209_6
timestamp 1731220653
transform 1 0 1808 0 1 896
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5208_6
timestamp 1731220653
transform 1 0 1696 0 1 896
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5207_6
timestamp 1731220653
transform 1 0 1584 0 1 896
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5206_6
timestamp 1731220653
transform 1 0 1480 0 1 896
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5205_6
timestamp 1731220653
transform 1 0 1400 0 1 896
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5204_6
timestamp 1731220653
transform 1 0 1344 0 1 896
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5203_6
timestamp 1731220653
transform 1 0 1344 0 -1 1012
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5202_6
timestamp 1731220653
transform 1 0 1216 0 -1 980
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5201_6
timestamp 1731220653
transform 1 0 1000 0 1 980
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5200_6
timestamp 1731220653
transform 1 0 920 0 1 980
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5199_6
timestamp 1731220653
transform 1 0 832 0 1 980
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5198_6
timestamp 1731220653
transform 1 0 744 0 1 980
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5197_6
timestamp 1731220653
transform 1 0 1136 0 -1 1092
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5196_6
timestamp 1731220653
transform 1 0 1048 0 -1 1092
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5195_6
timestamp 1731220653
transform 1 0 968 0 -1 1092
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5194_6
timestamp 1731220653
transform 1 0 888 0 -1 1092
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5193_6
timestamp 1731220653
transform 1 0 808 0 -1 1092
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5192_6
timestamp 1731220653
transform 1 0 720 0 -1 1092
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5191_6
timestamp 1731220653
transform 1 0 1016 0 1 1100
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5190_6
timestamp 1731220653
transform 1 0 936 0 1 1100
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5189_6
timestamp 1731220653
transform 1 0 856 0 1 1100
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5188_6
timestamp 1731220653
transform 1 0 784 0 1 1100
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5187_6
timestamp 1731220653
transform 1 0 712 0 1 1100
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5186_6
timestamp 1731220653
transform 1 0 632 0 1 1100
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5185_6
timestamp 1731220653
transform 1 0 856 0 -1 1208
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5184_6
timestamp 1731220653
transform 1 0 784 0 -1 1208
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5183_6
timestamp 1731220653
transform 1 0 712 0 -1 1208
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5182_6
timestamp 1731220653
transform 1 0 640 0 -1 1208
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5181_6
timestamp 1731220653
transform 1 0 576 0 -1 1208
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5180_6
timestamp 1731220653
transform 1 0 600 0 1 1212
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5179_6
timestamp 1731220653
transform 1 0 672 0 1 1212
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5178_6
timestamp 1731220653
transform 1 0 896 0 1 1212
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5177_6
timestamp 1731220653
transform 1 0 816 0 1 1212
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5176_6
timestamp 1731220653
transform 1 0 744 0 1 1212
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5175_6
timestamp 1731220653
transform 1 0 680 0 -1 1324
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5174_6
timestamp 1731220653
transform 1 0 776 0 -1 1324
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5173_6
timestamp 1731220653
transform 1 0 872 0 -1 1324
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5172_6
timestamp 1731220653
transform 1 0 968 0 -1 1324
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5171_6
timestamp 1731220653
transform 1 0 904 0 1 1340
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5170_6
timestamp 1731220653
transform 1 0 992 0 1 1340
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5169_6
timestamp 1731220653
transform 1 0 1080 0 1 1340
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5168_6
timestamp 1731220653
transform 1 0 1176 0 1 1340
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5167_6
timestamp 1731220653
transform 1 0 1216 0 -1 1448
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5166_6
timestamp 1731220653
transform 1 0 1120 0 -1 1448
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5165_6
timestamp 1731220653
transform 1 0 1016 0 -1 1448
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5164_6
timestamp 1731220653
transform 1 0 912 0 -1 1448
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5163_6
timestamp 1731220653
transform 1 0 1120 0 1 1452
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5162_6
timestamp 1731220653
transform 1 0 1032 0 1 1452
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5161_6
timestamp 1731220653
transform 1 0 952 0 1 1452
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5160_6
timestamp 1731220653
transform 1 0 872 0 1 1452
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5159_6
timestamp 1731220653
transform 1 0 840 0 -1 1564
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5158_6
timestamp 1731220653
transform 1 0 920 0 -1 1564
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5157_6
timestamp 1731220653
transform 1 0 1000 0 -1 1564
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5156_6
timestamp 1731220653
transform 1 0 984 0 1 1564
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5155_6
timestamp 1731220653
transform 1 0 1096 0 1 1564
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5154_6
timestamp 1731220653
transform 1 0 1056 0 -1 1672
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5153_6
timestamp 1731220653
transform 1 0 952 0 -1 1672
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5152_6
timestamp 1731220653
transform 1 0 1160 0 -1 1672
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5151_6
timestamp 1731220653
transform 1 0 1136 0 1 1676
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5150_6
timestamp 1731220653
transform 1 0 1024 0 1 1676
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5149_6
timestamp 1731220653
transform 1 0 968 0 -1 1784
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5148_6
timestamp 1731220653
transform 1 0 1056 0 -1 1784
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5147_6
timestamp 1731220653
transform 1 0 1144 0 -1 1784
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5146_6
timestamp 1731220653
transform 1 0 1136 0 1 1796
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5145_6
timestamp 1731220653
transform 1 0 1056 0 1 1796
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5144_6
timestamp 1731220653
transform 1 0 976 0 1 1796
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5143_6
timestamp 1731220653
transform 1 0 1152 0 -1 1900
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5142_6
timestamp 1731220653
transform 1 0 1080 0 -1 1900
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5141_6
timestamp 1731220653
transform 1 0 936 0 -1 1900
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5140_6
timestamp 1731220653
transform 1 0 864 0 -1 1900
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5139_6
timestamp 1731220653
transform 1 0 792 0 -1 1900
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5138_6
timestamp 1731220653
transform 1 0 712 0 -1 1900
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5137_6
timestamp 1731220653
transform 1 0 664 0 1 1796
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5136_6
timestamp 1731220653
transform 1 0 752 0 1 1796
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5135_6
timestamp 1731220653
transform 1 0 832 0 1 1796
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5134_6
timestamp 1731220653
transform 1 0 792 0 -1 1784
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5133_6
timestamp 1731220653
transform 1 0 696 0 -1 1784
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5132_6
timestamp 1731220653
transform 1 0 688 0 1 1676
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5131_6
timestamp 1731220653
transform 1 0 800 0 1 1676
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5130_6
timestamp 1731220653
transform 1 0 760 0 -1 1672
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5129_6
timestamp 1731220653
transform 1 0 664 0 -1 1672
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5128_6
timestamp 1731220653
transform 1 0 768 0 1 1564
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5127_6
timestamp 1731220653
transform 1 0 672 0 1 1564
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5126_6
timestamp 1731220653
transform 1 0 664 0 -1 1564
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5125_6
timestamp 1731220653
transform 1 0 632 0 1 1452
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5124_6
timestamp 1731220653
transform 1 0 552 0 1 1452
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5123_6
timestamp 1731220653
transform 1 0 600 0 -1 1448
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5122_6
timestamp 1731220653
transform 1 0 704 0 -1 1448
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5121_6
timestamp 1731220653
transform 1 0 640 0 1 1340
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5120_6
timestamp 1731220653
transform 1 0 560 0 1 1340
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5119_6
timestamp 1731220653
transform 1 0 480 0 1 1340
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5118_6
timestamp 1731220653
transform 1 0 408 0 1 1340
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5117_6
timestamp 1731220653
transform 1 0 336 0 1 1340
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5116_6
timestamp 1731220653
transform 1 0 272 0 1 1340
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5115_6
timestamp 1731220653
transform 1 0 320 0 -1 1448
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5114_6
timestamp 1731220653
transform 1 0 400 0 -1 1448
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5113_6
timestamp 1731220653
transform 1 0 496 0 -1 1448
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5112_6
timestamp 1731220653
transform 1 0 472 0 1 1452
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5111_6
timestamp 1731220653
transform 1 0 392 0 1 1452
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5110_6
timestamp 1731220653
transform 1 0 320 0 1 1452
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5109_6
timestamp 1731220653
transform 1 0 312 0 -1 1564
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5108_6
timestamp 1731220653
transform 1 0 392 0 -1 1564
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5107_6
timestamp 1731220653
transform 1 0 576 0 -1 1564
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5106_6
timestamp 1731220653
transform 1 0 480 0 -1 1564
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5105_6
timestamp 1731220653
transform 1 0 408 0 1 1564
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5104_6
timestamp 1731220653
transform 1 0 336 0 1 1564
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5103_6
timestamp 1731220653
transform 1 0 280 0 1 1564
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5102_6
timestamp 1731220653
transform 1 0 480 0 -1 1672
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5101_6
timestamp 1731220653
transform 1 0 392 0 -1 1672
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5100_6
timestamp 1731220653
transform 1 0 312 0 -1 1672
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_599_6
timestamp 1731220653
transform 1 0 248 0 -1 1672
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_598_6
timestamp 1731220653
transform 1 0 480 0 1 1676
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_597_6
timestamp 1731220653
transform 1 0 384 0 1 1676
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_596_6
timestamp 1731220653
transform 1 0 296 0 1 1676
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_595_6
timestamp 1731220653
transform 1 0 216 0 1 1676
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_594_6
timestamp 1731220653
transform 1 0 144 0 1 1676
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_593_6
timestamp 1731220653
transform 1 0 392 0 -1 1784
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_592_6
timestamp 1731220653
transform 1 0 288 0 -1 1784
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_591_6
timestamp 1731220653
transform 1 0 192 0 -1 1784
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_590_6
timestamp 1731220653
transform 1 0 128 0 -1 1784
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_589_6
timestamp 1731220653
transform 1 0 472 0 1 1796
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_588_6
timestamp 1731220653
transform 1 0 368 0 1 1796
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_587_6
timestamp 1731220653
transform 1 0 272 0 1 1796
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_586_6
timestamp 1731220653
transform 1 0 184 0 1 1796
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_585_6
timestamp 1731220653
transform 1 0 128 0 1 1796
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_584_6
timestamp 1731220653
transform 1 0 128 0 -1 1900
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_583_6
timestamp 1731220653
transform 1 0 184 0 -1 1900
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_582_6
timestamp 1731220653
transform 1 0 264 0 -1 1900
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_581_6
timestamp 1731220653
transform 1 0 448 0 -1 1900
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_580_6
timestamp 1731220653
transform 1 0 352 0 -1 1900
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_579_6
timestamp 1731220653
transform 1 0 296 0 1 1908
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_578_6
timestamp 1731220653
transform 1 0 192 0 1 1908
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_577_6
timestamp 1731220653
transform 1 0 128 0 1 1908
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_576_6
timestamp 1731220653
transform 1 0 560 0 1 1908
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_575_6
timestamp 1731220653
transform 1 0 416 0 1 1908
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_574_6
timestamp 1731220653
transform 1 0 352 0 -1 2016
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_573_6
timestamp 1731220653
transform 1 0 280 0 -1 2016
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_572_6
timestamp 1731220653
transform 1 0 224 0 -1 2016
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_571_6
timestamp 1731220653
transform 1 0 624 0 -1 2016
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_570_6
timestamp 1731220653
transform 1 0 528 0 -1 2016
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_569_6
timestamp 1731220653
transform 1 0 432 0 -1 2016
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_568_6
timestamp 1731220653
transform 1 0 376 0 1 2020
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_567_6
timestamp 1731220653
transform 1 0 432 0 1 2020
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_566_6
timestamp 1731220653
transform 1 0 488 0 1 2020
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_565_6
timestamp 1731220653
transform 1 0 552 0 1 2020
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_564_6
timestamp 1731220653
transform 1 0 616 0 1 2020
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_563_6
timestamp 1731220653
transform 1 0 624 0 -1 2128
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_562_6
timestamp 1731220653
transform 1 0 552 0 -1 2128
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_561_6
timestamp 1731220653
transform 1 0 480 0 -1 2128
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_560_6
timestamp 1731220653
transform 1 0 416 0 -1 2128
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_559_6
timestamp 1731220653
transform 1 0 352 0 -1 2128
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_558_6
timestamp 1731220653
transform 1 0 296 0 -1 2128
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_557_6
timestamp 1731220653
transform 1 0 536 0 1 2128
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_556_6
timestamp 1731220653
transform 1 0 432 0 1 2128
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_555_6
timestamp 1731220653
transform 1 0 328 0 1 2128
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_554_6
timestamp 1731220653
transform 1 0 232 0 1 2128
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_553_6
timestamp 1731220653
transform 1 0 512 0 -1 2232
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_552_6
timestamp 1731220653
transform 1 0 408 0 -1 2232
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_551_6
timestamp 1731220653
transform 1 0 312 0 -1 2232
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_550_6
timestamp 1731220653
transform 1 0 224 0 -1 2232
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_549_6
timestamp 1731220653
transform 1 0 136 0 -1 2232
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_548_6
timestamp 1731220653
transform 1 0 152 0 1 2232
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_547_6
timestamp 1731220653
transform 1 0 248 0 1 2232
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_546_6
timestamp 1731220653
transform 1 0 352 0 1 2232
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_545_6
timestamp 1731220653
transform 1 0 568 0 1 2232
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_544_6
timestamp 1731220653
transform 1 0 456 0 1 2232
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_543_6
timestamp 1731220653
transform 1 0 384 0 -1 2344
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_542_6
timestamp 1731220653
transform 1 0 312 0 -1 2344
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_541_6
timestamp 1731220653
transform 1 0 456 0 -1 2344
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_540_6
timestamp 1731220653
transform 1 0 528 0 -1 2344
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_539_6
timestamp 1731220653
transform 1 0 496 0 1 2352
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_538_6
timestamp 1731220653
transform 1 0 552 0 1 2352
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_537_6
timestamp 1731220653
transform 1 0 608 0 1 2352
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_536_6
timestamp 1731220653
transform 1 0 664 0 1 2352
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_535_6
timestamp 1731220653
transform 1 0 888 0 -1 2468
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_534_6
timestamp 1731220653
transform 1 0 944 0 -1 2468
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_533_6
timestamp 1731220653
transform 1 0 1000 0 -1 2468
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_532_6
timestamp 1731220653
transform 1 0 1056 0 -1 2468
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_531_6
timestamp 1731220653
transform 1 0 1040 0 1 2476
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_530_6
timestamp 1731220653
transform 1 0 976 0 1 2476
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_529_6
timestamp 1731220653
transform 1 0 912 0 1 2476
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_528_6
timestamp 1731220653
transform 1 0 848 0 1 2476
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_527_6
timestamp 1731220653
transform 1 0 784 0 1 2476
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_526_6
timestamp 1731220653
transform 1 0 720 0 1 2476
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_525_6
timestamp 1731220653
transform 1 0 656 0 1 2476
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_524_6
timestamp 1731220653
transform 1 0 592 0 1 2476
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_523_6
timestamp 1731220653
transform 1 0 528 0 1 2476
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_522_6
timestamp 1731220653
transform 1 0 832 0 -1 2468
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_521_6
timestamp 1731220653
transform 1 0 776 0 -1 2468
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_520_6
timestamp 1731220653
transform 1 0 720 0 -1 2468
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_519_6
timestamp 1731220653
transform 1 0 664 0 -1 2468
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_518_6
timestamp 1731220653
transform 1 0 608 0 -1 2468
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_517_6
timestamp 1731220653
transform 1 0 552 0 -1 2468
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_516_6
timestamp 1731220653
transform 1 0 496 0 -1 2468
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_515_6
timestamp 1731220653
transform 1 0 440 0 -1 2468
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_514_6
timestamp 1731220653
transform 1 0 384 0 -1 2468
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_513_6
timestamp 1731220653
transform 1 0 328 0 -1 2468
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_512_6
timestamp 1731220653
transform 1 0 272 0 -1 2468
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_511_6
timestamp 1731220653
transform 1 0 216 0 -1 2468
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_510_6
timestamp 1731220653
transform 1 0 160 0 -1 2468
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_59_6
timestamp 1731220653
transform 1 0 464 0 1 2476
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_58_6
timestamp 1731220653
transform 1 0 392 0 1 2476
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_57_6
timestamp 1731220653
transform 1 0 320 0 1 2476
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_56_6
timestamp 1731220653
transform 1 0 256 0 1 2476
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_55_6
timestamp 1731220653
transform 1 0 200 0 1 2476
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_54_6
timestamp 1731220653
transform 1 0 352 0 -1 2580
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_53_6
timestamp 1731220653
transform 1 0 296 0 -1 2580
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_52_6
timestamp 1731220653
transform 1 0 240 0 -1 2580
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_51_6
timestamp 1731220653
transform 1 0 184 0 -1 2580
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_50_6
timestamp 1731220653
transform 1 0 128 0 -1 2580
box 4 4 48 48
<< end >>
