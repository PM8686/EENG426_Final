magic
tech sky130l
timestamp 1731220329
<< m1 >>
rect 2168 3463 2172 3483
rect 2312 3427 2316 3447
rect 2928 3427 2932 3467
rect 2912 3283 2916 3323
rect 3192 3283 3196 3303
rect 808 3255 812 3275
rect 1976 3183 1980 3203
rect 2448 3171 2452 3207
rect 2656 3147 2660 3167
rect 3360 3147 3364 3167
rect 592 3111 596 3131
rect 1184 2971 1188 2991
rect 2168 2871 2172 2891
rect 2568 2871 2572 2891
rect 2568 2775 2572 2799
rect 2848 2735 2852 2771
rect 1088 2691 1092 2711
rect 2600 2603 2604 2623
rect 2752 2603 2756 2623
rect 3240 2603 3244 2623
rect 1488 2563 1496 2567
rect 1488 2543 1492 2563
rect 232 2399 236 2419
rect 1576 2399 1580 2419
rect 2840 2355 2844 2379
rect 1272 2255 1276 2275
rect 1384 2255 1388 2275
rect 1408 2191 1412 2275
rect 2560 2251 2564 2339
rect 2600 2319 2604 2339
rect 944 2111 948 2131
rect 872 1983 876 2003
rect 1248 1983 1252 2015
rect 560 1891 564 1911
rect 792 1731 796 1779
rect 1472 1755 1476 1779
rect 1960 1739 1964 1759
rect 2616 1595 2620 1615
rect 408 1571 412 1591
rect 1048 1571 1052 1591
rect 736 1475 740 1499
rect 2024 1451 2028 1471
rect 216 1431 220 1451
rect 3056 1451 3060 1471
rect 3112 1351 3116 1375
rect 2504 1311 2508 1331
rect 1528 1051 1532 1087
rect 2328 1079 2332 1103
rect 3360 1079 3364 1103
rect 688 883 692 903
rect 976 883 980 903
rect 1448 883 1452 903
rect 2408 895 2412 915
rect 1504 675 1508 767
rect 1960 759 1964 779
rect 568 607 572 635
rect 1472 471 1476 491
rect 2568 487 2572 507
rect 728 335 732 355
rect 3248 235 3252 275
<< m2c >>
rect 2168 3483 2172 3487
rect 2928 3467 2932 3471
rect 2060 3459 2064 3463
rect 2168 3459 2172 3463
rect 2292 3459 2296 3463
rect 2508 3459 2512 3463
rect 2708 3461 2712 3465
rect 2908 3459 2912 3463
rect 1884 3447 1888 3451
rect 1996 3447 2000 3451
rect 2132 3447 2136 3451
rect 2268 3447 2272 3451
rect 2312 3447 2316 3451
rect 2404 3447 2408 3451
rect 2532 3447 2536 3451
rect 2652 3447 2656 3451
rect 2772 3447 2776 3451
rect 2900 3447 2904 3451
rect 508 3425 512 3429
rect 596 3423 600 3427
rect 684 3423 688 3427
rect 772 3423 776 3427
rect 860 3423 864 3427
rect 948 3423 952 3427
rect 1036 3425 1040 3429
rect 1124 3423 1128 3427
rect 1212 3423 1216 3427
rect 2312 3423 2316 3427
rect 3100 3459 3104 3463
rect 3300 3459 3304 3463
rect 3028 3447 3032 3451
rect 2928 3423 2932 3427
rect 468 3411 472 3415
rect 556 3411 560 3415
rect 644 3411 648 3415
rect 732 3411 736 3415
rect 820 3411 824 3415
rect 908 3411 912 3415
rect 996 3411 1000 3415
rect 1084 3411 1088 3415
rect 1172 3411 1176 3415
rect 1260 3411 1264 3415
rect 1356 3411 1360 3415
rect 1884 3323 1888 3327
rect 2004 3323 2008 3327
rect 2148 3323 2152 3327
rect 2292 3323 2296 3327
rect 2436 3323 2440 3327
rect 2572 3323 2576 3327
rect 2700 3323 2704 3327
rect 2828 3325 2832 3329
rect 2912 3323 2916 3327
rect 2956 3323 2960 3327
rect 3092 3323 3096 3327
rect 1884 3303 1888 3307
rect 2028 3303 2032 3307
rect 2204 3303 2208 3307
rect 2388 3303 2392 3307
rect 2564 3303 2568 3307
rect 2732 3303 2736 3307
rect 2884 3303 2888 3307
rect 452 3291 456 3295
rect 548 3291 552 3295
rect 652 3291 656 3295
rect 756 3291 760 3295
rect 860 3291 864 3295
rect 964 3293 968 3297
rect 1068 3291 1072 3295
rect 1172 3291 1176 3295
rect 1276 3291 1280 3295
rect 1380 3291 1384 3295
rect 3028 3303 3032 3307
rect 3164 3303 3168 3307
rect 3192 3303 3196 3307
rect 3300 3303 3304 3307
rect 3420 3303 3424 3307
rect 2912 3279 2916 3283
rect 3192 3279 3196 3283
rect 436 3275 440 3279
rect 548 3275 552 3279
rect 660 3275 664 3279
rect 780 3275 784 3279
rect 808 3275 812 3279
rect 900 3275 904 3279
rect 1020 3275 1024 3279
rect 1140 3275 1144 3279
rect 1260 3275 1264 3279
rect 1388 3275 1392 3279
rect 808 3251 812 3255
rect 2448 3207 2452 3211
rect 1976 3203 1980 3207
rect 1884 3179 1888 3183
rect 1976 3179 1980 3183
rect 2084 3179 2088 3183
rect 2300 3179 2304 3183
rect 2508 3179 2512 3183
rect 2708 3179 2712 3183
rect 2892 3179 2896 3183
rect 3076 3179 3080 3183
rect 3260 3179 3264 3183
rect 3420 3179 3424 3183
rect 1892 3167 1896 3171
rect 2084 3167 2088 3171
rect 2276 3167 2280 3171
rect 2448 3167 2452 3171
rect 2460 3167 2464 3171
rect 2628 3167 2632 3171
rect 2656 3167 2660 3171
rect 2788 3167 2792 3171
rect 2932 3167 2936 3171
rect 3060 3167 3064 3171
rect 3188 3167 3192 3171
rect 3316 3167 3320 3171
rect 3360 3167 3364 3171
rect 3420 3167 3424 3171
rect 356 3157 360 3161
rect 476 3155 480 3159
rect 596 3155 600 3159
rect 724 3155 728 3159
rect 852 3155 856 3159
rect 980 3155 984 3159
rect 1108 3155 1112 3159
rect 1228 3157 1232 3161
rect 1356 3155 1360 3159
rect 1484 3155 1488 3159
rect 2656 3143 2660 3147
rect 3360 3143 3364 3147
rect 228 3131 232 3135
rect 372 3131 376 3135
rect 524 3131 528 3135
rect 592 3131 596 3135
rect 676 3131 680 3135
rect 828 3131 832 3135
rect 972 3131 976 3135
rect 1116 3131 1120 3135
rect 1252 3131 1256 3135
rect 1396 3131 1400 3135
rect 1540 3131 1544 3135
rect 592 3107 596 3111
rect 1988 3047 1992 3051
rect 2108 3047 2112 3051
rect 2228 3047 2232 3051
rect 2356 3047 2360 3051
rect 2484 3047 2488 3051
rect 2620 3047 2624 3051
rect 2772 3047 2776 3051
rect 2924 3047 2928 3051
rect 3084 3047 3088 3051
rect 3252 3047 3256 3051
rect 3420 3047 3424 3051
rect 2076 3027 2080 3031
rect 2180 3027 2184 3031
rect 2284 3027 2288 3031
rect 2388 3027 2392 3031
rect 2492 3027 2496 3031
rect 2596 3027 2600 3031
rect 2700 3027 2704 3031
rect 2812 3027 2816 3031
rect 188 3009 192 3013
rect 316 3007 320 3011
rect 484 3007 488 3011
rect 660 3007 664 3011
rect 844 3007 848 3011
rect 1020 3007 1024 3011
rect 1196 3007 1200 3011
rect 1380 3007 1384 3011
rect 1564 3007 1568 3011
rect 188 2991 192 2995
rect 380 2991 384 2995
rect 588 2991 592 2995
rect 788 2991 792 2995
rect 980 2991 984 2995
rect 1156 2991 1160 2995
rect 1184 2991 1188 2995
rect 1332 2991 1336 2995
rect 1500 2991 1504 2995
rect 1676 2991 1680 2995
rect 1184 2967 1188 2971
rect 2108 2911 2112 2915
rect 2196 2911 2200 2915
rect 2284 2913 2288 2917
rect 2372 2911 2376 2915
rect 2460 2911 2464 2915
rect 2548 2911 2552 2915
rect 2636 2911 2640 2915
rect 2724 2911 2728 2915
rect 2812 2911 2816 2915
rect 2900 2911 2904 2915
rect 2124 2891 2128 2895
rect 2168 2891 2172 2895
rect 2228 2891 2232 2895
rect 2324 2891 2328 2895
rect 2420 2891 2424 2895
rect 2524 2891 2528 2895
rect 2568 2891 2572 2895
rect 2628 2891 2632 2895
rect 2732 2891 2736 2895
rect 2836 2891 2840 2895
rect 188 2867 192 2871
rect 316 2867 320 2871
rect 484 2867 488 2871
rect 660 2867 664 2871
rect 836 2867 840 2871
rect 1004 2867 1008 2871
rect 1164 2867 1168 2871
rect 1324 2867 1328 2871
rect 1484 2867 1488 2871
rect 1644 2867 1648 2871
rect 2168 2867 2172 2871
rect 2568 2867 2572 2871
rect 188 2853 192 2857
rect 308 2851 312 2855
rect 460 2851 464 2855
rect 620 2851 624 2855
rect 780 2851 784 2855
rect 932 2851 936 2855
rect 1076 2851 1080 2855
rect 1220 2851 1224 2855
rect 1364 2851 1368 2855
rect 1516 2851 1520 2855
rect 2568 2799 2572 2803
rect 2036 2771 2040 2775
rect 2164 2771 2168 2775
rect 2292 2771 2296 2775
rect 2420 2771 2424 2775
rect 2540 2771 2544 2775
rect 2568 2771 2572 2775
rect 2660 2771 2664 2775
rect 2772 2773 2776 2777
rect 2848 2771 2852 2775
rect 2892 2771 2896 2775
rect 3012 2771 3016 2775
rect 1940 2755 1944 2759
rect 2084 2755 2088 2759
rect 2236 2755 2240 2759
rect 2388 2755 2392 2759
rect 2532 2755 2536 2759
rect 2676 2755 2680 2759
rect 2820 2755 2824 2759
rect 2964 2755 2968 2759
rect 3108 2755 3112 2759
rect 340 2729 344 2733
rect 2848 2731 2852 2735
rect 444 2727 448 2731
rect 556 2727 560 2731
rect 676 2727 680 2731
rect 796 2727 800 2731
rect 908 2727 912 2731
rect 1020 2727 1024 2731
rect 1132 2727 1136 2731
rect 1252 2727 1256 2731
rect 1372 2727 1376 2731
rect 532 2713 536 2717
rect 620 2711 624 2715
rect 708 2711 712 2715
rect 796 2711 800 2715
rect 884 2711 888 2715
rect 972 2711 976 2715
rect 1060 2711 1064 2715
rect 1088 2711 1092 2715
rect 1148 2711 1152 2715
rect 1236 2711 1240 2715
rect 1088 2687 1092 2691
rect 1884 2639 1888 2643
rect 2076 2639 2080 2643
rect 2284 2639 2288 2643
rect 2484 2639 2488 2643
rect 2668 2639 2672 2643
rect 2836 2639 2840 2643
rect 2996 2639 3000 2643
rect 3148 2639 3152 2643
rect 3292 2639 3296 2643
rect 3420 2639 3424 2643
rect 1884 2623 1888 2627
rect 2052 2623 2056 2627
rect 2236 2623 2240 2627
rect 2412 2623 2416 2627
rect 2572 2623 2576 2627
rect 2600 2623 2604 2627
rect 2724 2623 2728 2627
rect 2752 2623 2756 2627
rect 2860 2623 2864 2627
rect 2980 2623 2984 2627
rect 3100 2623 3104 2627
rect 3212 2623 3216 2627
rect 3240 2623 3244 2627
rect 3324 2623 3328 2627
rect 3420 2623 3424 2627
rect 2600 2599 2604 2603
rect 2752 2599 2756 2603
rect 3240 2599 3244 2603
rect 524 2587 528 2591
rect 612 2587 616 2591
rect 700 2587 704 2591
rect 788 2587 792 2591
rect 876 2587 880 2591
rect 964 2587 968 2591
rect 1052 2587 1056 2591
rect 1140 2587 1144 2591
rect 276 2563 280 2567
rect 364 2563 368 2567
rect 460 2563 464 2567
rect 556 2563 560 2567
rect 644 2563 648 2567
rect 732 2563 736 2567
rect 820 2563 824 2567
rect 908 2563 912 2567
rect 996 2563 1000 2567
rect 1084 2563 1088 2567
rect 1172 2563 1176 2567
rect 1268 2563 1272 2567
rect 1364 2563 1368 2567
rect 1460 2563 1464 2567
rect 1496 2563 1500 2567
rect 1548 2563 1552 2567
rect 1636 2563 1640 2567
rect 1724 2563 1728 2567
rect 1488 2539 1492 2543
rect 2260 2499 2264 2503
rect 2852 2499 2856 2503
rect 3420 2499 3424 2503
rect 2068 2471 2072 2475
rect 2252 2471 2256 2475
rect 2420 2471 2424 2475
rect 2580 2471 2584 2475
rect 2724 2471 2728 2475
rect 2860 2471 2864 2475
rect 2980 2471 2984 2475
rect 3100 2471 3104 2475
rect 3212 2471 3216 2475
rect 3324 2471 3328 2475
rect 3420 2471 3424 2475
rect 188 2447 192 2451
rect 300 2449 304 2453
rect 444 2447 448 2451
rect 596 2447 600 2451
rect 748 2447 752 2451
rect 892 2447 896 2451
rect 1028 2447 1032 2451
rect 1156 2447 1160 2451
rect 1284 2447 1288 2451
rect 1404 2447 1408 2451
rect 1516 2449 1520 2453
rect 1628 2447 1632 2451
rect 1724 2447 1728 2451
rect 188 2419 192 2423
rect 232 2419 236 2423
rect 292 2419 296 2423
rect 444 2419 448 2423
rect 604 2419 608 2423
rect 772 2419 776 2423
rect 948 2419 952 2423
rect 1116 2419 1120 2423
rect 1292 2419 1296 2423
rect 1468 2419 1472 2423
rect 1576 2419 1580 2423
rect 1644 2419 1648 2423
rect 232 2395 236 2399
rect 1576 2395 1580 2399
rect 2840 2379 2844 2383
rect 1892 2351 1896 2355
rect 2060 2351 2064 2355
rect 2236 2351 2240 2355
rect 2420 2351 2424 2355
rect 2612 2351 2616 2355
rect 2812 2351 2816 2355
rect 2840 2351 2844 2355
rect 3020 2351 3024 2355
rect 3228 2351 3232 2355
rect 3420 2351 3424 2355
rect 1940 2339 1944 2343
rect 2068 2339 2072 2343
rect 2204 2339 2208 2343
rect 2356 2339 2360 2343
rect 2516 2339 2520 2343
rect 2560 2339 2564 2343
rect 428 2297 432 2301
rect 532 2295 536 2299
rect 652 2295 656 2299
rect 772 2295 776 2299
rect 900 2295 904 2299
rect 1028 2295 1032 2299
rect 1156 2295 1160 2299
rect 1292 2295 1296 2299
rect 1428 2295 1432 2299
rect 1564 2295 1568 2299
rect 628 2277 632 2281
rect 716 2275 720 2279
rect 812 2275 816 2279
rect 916 2275 920 2279
rect 1020 2275 1024 2279
rect 1132 2275 1136 2279
rect 1244 2275 1248 2279
rect 1272 2275 1276 2279
rect 1356 2275 1360 2279
rect 1384 2275 1388 2279
rect 1272 2251 1276 2255
rect 1384 2251 1388 2255
rect 1408 2275 1412 2279
rect 1468 2275 1472 2279
rect 2600 2339 2604 2343
rect 2700 2339 2704 2343
rect 2892 2339 2896 2343
rect 3100 2339 3104 2343
rect 3308 2339 3312 2343
rect 2600 2315 2604 2319
rect 2560 2247 2564 2251
rect 2092 2221 2096 2225
rect 2188 2219 2192 2223
rect 2292 2219 2296 2223
rect 2396 2219 2400 2223
rect 2516 2219 2520 2223
rect 2644 2219 2648 2223
rect 2788 2219 2792 2223
rect 2940 2219 2944 2223
rect 3100 2219 3104 2223
rect 3268 2219 3272 2223
rect 3420 2219 3424 2223
rect 2236 2197 2240 2201
rect 2332 2195 2336 2199
rect 2436 2195 2440 2199
rect 2548 2195 2552 2199
rect 2660 2195 2664 2199
rect 2772 2195 2776 2199
rect 2892 2195 2896 2199
rect 3020 2195 3024 2199
rect 3156 2195 3160 2199
rect 3300 2195 3304 2199
rect 3420 2195 3424 2199
rect 1408 2187 1412 2191
rect 492 2159 496 2163
rect 580 2159 584 2163
rect 668 2159 672 2163
rect 756 2159 760 2163
rect 844 2159 848 2163
rect 932 2161 936 2165
rect 1020 2159 1024 2163
rect 1108 2159 1112 2163
rect 1196 2159 1200 2163
rect 1284 2159 1288 2163
rect 1372 2159 1376 2163
rect 356 2131 360 2135
rect 460 2131 464 2135
rect 572 2131 576 2135
rect 684 2131 688 2135
rect 796 2131 800 2135
rect 916 2131 920 2135
rect 944 2131 948 2135
rect 1036 2131 1040 2135
rect 944 2107 948 2111
rect 2188 2071 2192 2075
rect 2308 2071 2312 2075
rect 2436 2071 2440 2075
rect 2572 2071 2576 2075
rect 2708 2071 2712 2075
rect 2836 2073 2840 2077
rect 2964 2071 2968 2075
rect 3084 2071 3088 2075
rect 3204 2071 3208 2075
rect 3324 2071 3328 2075
rect 3420 2071 3424 2075
rect 2300 2051 2304 2055
rect 2468 2051 2472 2055
rect 2628 2051 2632 2055
rect 2780 2051 2784 2055
rect 2924 2051 2928 2055
rect 3060 2051 3064 2055
rect 3188 2051 3192 2055
rect 3316 2051 3320 2055
rect 3420 2051 3424 2055
rect 308 2015 312 2019
rect 428 2015 432 2019
rect 548 2015 552 2019
rect 668 2017 672 2021
rect 780 2015 784 2019
rect 884 2017 888 2021
rect 988 2015 992 2019
rect 1092 2015 1096 2019
rect 1196 2015 1200 2019
rect 1248 2015 1252 2019
rect 1308 2015 1312 2019
rect 412 2003 416 2007
rect 540 2003 544 2007
rect 676 2003 680 2007
rect 812 2003 816 2007
rect 872 2003 876 2007
rect 948 2003 952 2007
rect 1076 2003 1080 2007
rect 1204 2003 1208 2007
rect 872 1979 876 1983
rect 1324 2003 1328 2007
rect 1452 2003 1456 2007
rect 1580 2003 1584 2007
rect 1248 1979 1252 1983
rect 1884 1919 1888 1923
rect 1972 1919 1976 1923
rect 2100 1919 2104 1923
rect 2236 1919 2240 1923
rect 2380 1919 2384 1923
rect 2524 1919 2528 1923
rect 2668 1919 2672 1923
rect 2804 1919 2808 1923
rect 2940 1919 2944 1923
rect 3084 1919 3088 1923
rect 3228 1919 3232 1923
rect 3372 1919 3376 1923
rect 560 1911 564 1915
rect 1884 1903 1888 1907
rect 1972 1905 1976 1909
rect 2092 1903 2096 1907
rect 2220 1903 2224 1907
rect 2356 1903 2360 1907
rect 2508 1903 2512 1907
rect 2668 1903 2672 1907
rect 2844 1903 2848 1907
rect 3036 1903 3040 1907
rect 3236 1903 3240 1907
rect 3420 1903 3424 1907
rect 500 1887 504 1891
rect 560 1887 564 1891
rect 628 1887 632 1891
rect 764 1887 768 1891
rect 900 1887 904 1891
rect 1036 1887 1040 1891
rect 1172 1889 1176 1893
rect 1308 1887 1312 1891
rect 1436 1887 1440 1891
rect 1572 1887 1576 1891
rect 1708 1887 1712 1891
rect 612 1875 616 1879
rect 748 1875 752 1879
rect 884 1875 888 1879
rect 1012 1875 1016 1879
rect 1132 1875 1136 1879
rect 1252 1875 1256 1879
rect 1380 1875 1384 1879
rect 1508 1875 1512 1879
rect 1884 1783 1888 1787
rect 2012 1783 2016 1787
rect 2164 1783 2168 1787
rect 2308 1783 2312 1787
rect 2460 1783 2464 1787
rect 2620 1783 2624 1787
rect 2796 1783 2800 1787
rect 2988 1783 2992 1787
rect 3188 1783 3192 1787
rect 3396 1783 3400 1787
rect 792 1779 796 1783
rect 188 1751 192 1755
rect 276 1751 280 1755
rect 364 1751 368 1755
rect 460 1751 464 1755
rect 580 1751 584 1755
rect 708 1751 712 1755
rect 1472 1779 1476 1783
rect 1932 1759 1936 1763
rect 1960 1759 1964 1763
rect 2068 1759 2072 1763
rect 2204 1759 2208 1763
rect 2356 1759 2360 1763
rect 2532 1759 2536 1763
rect 2740 1759 2744 1763
rect 2964 1761 2968 1765
rect 3204 1759 3208 1763
rect 3420 1759 3424 1763
rect 852 1751 856 1755
rect 996 1751 1000 1755
rect 1140 1751 1144 1755
rect 1292 1751 1296 1755
rect 1444 1751 1448 1755
rect 1472 1751 1476 1755
rect 1596 1751 1600 1755
rect 1724 1751 1728 1755
rect 1960 1735 1964 1739
rect 188 1727 192 1731
rect 300 1727 304 1731
rect 452 1727 456 1731
rect 620 1727 624 1731
rect 792 1727 796 1731
rect 804 1727 808 1731
rect 988 1727 992 1731
rect 1172 1727 1176 1731
rect 1364 1727 1368 1731
rect 1556 1727 1560 1731
rect 1724 1727 1728 1731
rect 1884 1635 1888 1639
rect 1988 1635 1992 1639
rect 2116 1635 2120 1639
rect 2236 1635 2240 1639
rect 2364 1635 2368 1639
rect 2492 1637 2496 1641
rect 2628 1635 2632 1639
rect 2780 1635 2784 1639
rect 2940 1635 2944 1639
rect 3100 1635 3104 1639
rect 3268 1635 3272 1639
rect 3420 1635 3424 1639
rect 1884 1615 1888 1619
rect 1996 1615 2000 1619
rect 2140 1615 2144 1619
rect 2284 1615 2288 1619
rect 2420 1615 2424 1619
rect 2556 1615 2560 1619
rect 2616 1615 2620 1619
rect 2692 1615 2696 1619
rect 2820 1615 2824 1619
rect 2948 1615 2952 1619
rect 3068 1615 3072 1619
rect 3188 1615 3192 1619
rect 3316 1615 3320 1619
rect 3420 1615 3424 1619
rect 244 1607 248 1611
rect 348 1607 352 1611
rect 460 1607 464 1611
rect 588 1607 592 1611
rect 740 1607 744 1611
rect 908 1607 912 1611
rect 1092 1607 1096 1611
rect 1284 1607 1288 1611
rect 1484 1607 1488 1611
rect 1692 1607 1696 1611
rect 380 1591 384 1595
rect 408 1591 412 1595
rect 484 1591 488 1595
rect 596 1591 600 1595
rect 724 1591 728 1595
rect 868 1591 872 1595
rect 1020 1591 1024 1595
rect 1048 1591 1052 1595
rect 1172 1591 1176 1595
rect 1332 1591 1336 1595
rect 1492 1591 1496 1595
rect 1660 1591 1664 1595
rect 2616 1591 2620 1595
rect 408 1567 412 1571
rect 1048 1567 1052 1571
rect 736 1499 740 1503
rect 1892 1491 1896 1495
rect 2044 1491 2048 1495
rect 2204 1491 2208 1495
rect 2356 1491 2360 1495
rect 2508 1491 2512 1495
rect 2652 1491 2656 1495
rect 2788 1491 2792 1495
rect 2924 1491 2928 1495
rect 3060 1491 3064 1495
rect 3196 1491 3200 1495
rect 276 1471 280 1475
rect 396 1471 400 1475
rect 524 1471 528 1475
rect 660 1471 664 1475
rect 736 1471 740 1475
rect 804 1471 808 1475
rect 948 1471 952 1475
rect 1100 1471 1104 1475
rect 1252 1471 1256 1475
rect 1404 1471 1408 1475
rect 1556 1471 1560 1475
rect 1996 1471 2000 1475
rect 2024 1471 2028 1475
rect 2108 1471 2112 1475
rect 2244 1471 2248 1475
rect 2388 1471 2392 1475
rect 2532 1471 2536 1475
rect 2684 1471 2688 1475
rect 2836 1471 2840 1475
rect 2988 1471 2992 1475
rect 3056 1471 3060 1475
rect 3140 1471 3144 1475
rect 3292 1471 3296 1475
rect 188 1451 192 1455
rect 216 1451 220 1455
rect 356 1451 360 1455
rect 524 1451 528 1455
rect 684 1451 688 1455
rect 836 1451 840 1455
rect 980 1451 984 1455
rect 1116 1451 1120 1455
rect 1252 1451 1256 1455
rect 1388 1451 1392 1455
rect 1524 1451 1528 1455
rect 2024 1447 2028 1451
rect 3056 1447 3060 1451
rect 216 1427 220 1431
rect 3112 1375 3116 1379
rect 2148 1349 2152 1353
rect 2252 1347 2256 1351
rect 2372 1347 2376 1351
rect 2508 1347 2512 1351
rect 2652 1347 2656 1351
rect 2796 1347 2800 1351
rect 2940 1347 2944 1351
rect 3084 1347 3088 1351
rect 3112 1347 3116 1351
rect 3228 1347 3232 1351
rect 3380 1347 3384 1351
rect 188 1331 192 1335
rect 332 1331 336 1335
rect 500 1331 504 1335
rect 660 1331 664 1335
rect 812 1331 816 1335
rect 956 1331 960 1335
rect 1084 1331 1088 1335
rect 1212 1331 1216 1335
rect 1340 1331 1344 1335
rect 1468 1331 1472 1335
rect 2156 1331 2160 1335
rect 2292 1331 2296 1335
rect 2436 1331 2440 1335
rect 2504 1331 2508 1335
rect 2588 1331 2592 1335
rect 2740 1331 2744 1335
rect 2892 1331 2896 1335
rect 3044 1331 3048 1335
rect 3196 1331 3200 1335
rect 3356 1331 3360 1335
rect 188 1315 192 1319
rect 332 1317 336 1321
rect 492 1315 496 1319
rect 636 1315 640 1319
rect 772 1315 776 1319
rect 900 1315 904 1319
rect 1020 1315 1024 1319
rect 1132 1315 1136 1319
rect 1244 1315 1248 1319
rect 1364 1315 1368 1319
rect 2504 1307 2508 1311
rect 1988 1217 1992 1221
rect 2116 1215 2120 1219
rect 2252 1215 2256 1219
rect 2396 1215 2400 1219
rect 2548 1215 2552 1219
rect 2708 1215 2712 1219
rect 2868 1215 2872 1219
rect 3028 1215 3032 1219
rect 3196 1215 3200 1219
rect 1884 1203 1888 1207
rect 1988 1203 1992 1207
rect 2132 1203 2136 1207
rect 2284 1203 2288 1207
rect 2444 1203 2448 1207
rect 2596 1203 2600 1207
rect 2748 1203 2752 1207
rect 2900 1203 2904 1207
rect 3052 1203 3056 1207
rect 3212 1203 3216 1207
rect 188 1195 192 1199
rect 292 1195 296 1199
rect 420 1195 424 1199
rect 548 1195 552 1199
rect 668 1195 672 1199
rect 788 1197 792 1201
rect 900 1195 904 1199
rect 1012 1195 1016 1199
rect 1124 1195 1128 1199
rect 1244 1195 1248 1199
rect 188 1179 192 1183
rect 292 1179 296 1183
rect 428 1179 432 1183
rect 564 1179 568 1183
rect 708 1179 712 1183
rect 844 1181 848 1185
rect 980 1179 984 1183
rect 1116 1179 1120 1183
rect 1252 1179 1256 1183
rect 1388 1179 1392 1183
rect 2328 1103 2332 1107
rect 1528 1087 1532 1091
rect 244 1059 248 1063
rect 388 1059 392 1063
rect 548 1061 552 1065
rect 708 1059 712 1063
rect 868 1059 872 1063
rect 1020 1061 1024 1065
rect 1172 1059 1176 1063
rect 1316 1059 1320 1063
rect 1460 1059 1464 1063
rect 3360 1103 3364 1107
rect 1916 1075 1920 1079
rect 2036 1075 2040 1079
rect 2164 1075 2168 1079
rect 2300 1075 2304 1079
rect 2328 1075 2332 1079
rect 2436 1075 2440 1079
rect 2564 1075 2568 1079
rect 2692 1077 2696 1081
rect 2812 1075 2816 1079
rect 2924 1075 2928 1079
rect 3028 1075 3032 1079
rect 3132 1075 3136 1079
rect 3236 1075 3240 1079
rect 3332 1075 3336 1079
rect 3360 1075 3364 1079
rect 3420 1075 3424 1079
rect 1612 1059 1616 1063
rect 2156 1055 2160 1059
rect 2244 1057 2248 1061
rect 2332 1055 2336 1059
rect 2420 1055 2424 1059
rect 2508 1055 2512 1059
rect 2596 1055 2600 1059
rect 2684 1055 2688 1059
rect 2772 1055 2776 1059
rect 2860 1055 2864 1059
rect 1528 1047 1532 1051
rect 380 1039 384 1043
rect 516 1041 520 1045
rect 660 1039 664 1043
rect 820 1039 824 1043
rect 980 1039 984 1043
rect 1132 1039 1136 1043
rect 1284 1041 1288 1045
rect 1436 1039 1440 1043
rect 1588 1039 1592 1043
rect 1724 1039 1728 1043
rect 2364 939 2368 943
rect 2460 939 2464 943
rect 2564 939 2568 943
rect 2676 941 2680 945
rect 2804 939 2808 943
rect 2948 939 2952 943
rect 3108 939 3112 943
rect 3276 939 3280 943
rect 3420 939 3424 943
rect 524 919 528 923
rect 620 919 624 923
rect 724 919 728 923
rect 836 919 840 923
rect 940 919 944 923
rect 1044 919 1048 923
rect 1148 919 1152 923
rect 1252 919 1256 923
rect 1348 919 1352 923
rect 1444 919 1448 923
rect 1540 921 1544 925
rect 1636 919 1640 923
rect 1724 919 1728 923
rect 1884 915 1888 919
rect 2036 915 2040 919
rect 2204 915 2208 919
rect 2380 915 2384 919
rect 2408 915 2412 919
rect 2572 915 2576 919
rect 2772 915 2776 919
rect 2988 917 2992 921
rect 3212 915 3216 919
rect 3420 915 3424 919
rect 660 903 664 907
rect 688 903 692 907
rect 748 903 752 907
rect 844 903 848 907
rect 948 903 952 907
rect 976 903 980 907
rect 1052 903 1056 907
rect 1164 903 1168 907
rect 1276 903 1280 907
rect 1396 903 1400 907
rect 1448 903 1452 907
rect 1516 903 1520 907
rect 1636 903 1640 907
rect 688 879 692 883
rect 976 879 980 883
rect 2408 891 2412 895
rect 1448 879 1452 883
rect 1884 795 1888 799
rect 2012 795 2016 799
rect 2140 797 2144 801
rect 2260 795 2264 799
rect 2380 795 2384 799
rect 2516 795 2520 799
rect 2668 795 2672 799
rect 2844 795 2848 799
rect 3036 795 3040 799
rect 3236 795 3240 799
rect 3420 795 3424 799
rect 572 783 576 787
rect 668 785 672 789
rect 772 783 776 787
rect 884 783 888 787
rect 1004 783 1008 787
rect 1124 783 1128 787
rect 1244 783 1248 787
rect 1364 783 1368 787
rect 1484 783 1488 787
rect 1612 783 1616 787
rect 1932 779 1936 783
rect 1960 779 1964 783
rect 2068 779 2072 783
rect 2204 779 2208 783
rect 2340 779 2344 783
rect 2476 779 2480 783
rect 2612 781 2616 785
rect 2764 779 2768 783
rect 2924 779 2928 783
rect 3092 779 3096 783
rect 3268 779 3272 783
rect 3420 779 3424 783
rect 436 767 440 771
rect 524 767 528 771
rect 628 767 632 771
rect 732 767 736 771
rect 844 767 848 771
rect 964 767 968 771
rect 1084 767 1088 771
rect 1212 767 1216 771
rect 1340 767 1344 771
rect 1468 767 1472 771
rect 1504 767 1508 771
rect 984 735 988 739
rect 1960 755 1964 759
rect 1952 747 1956 751
rect 1504 671 1508 675
rect 1884 659 1888 663
rect 2004 659 2008 663
rect 2156 659 2160 663
rect 2316 659 2320 663
rect 2468 659 2472 663
rect 2620 659 2624 663
rect 2772 659 2776 663
rect 2932 661 2936 665
rect 3092 659 3096 663
rect 3252 659 3256 663
rect 2028 647 2032 651
rect 2292 647 2296 651
rect 2532 647 2536 651
rect 2740 647 2744 651
rect 2932 647 2936 651
rect 3108 647 3112 651
rect 3276 647 3280 651
rect 3420 647 3424 651
rect 300 643 304 647
rect 396 643 400 647
rect 508 643 512 647
rect 620 643 624 647
rect 748 643 752 647
rect 884 643 888 647
rect 1036 643 1040 647
rect 1204 643 1208 647
rect 1380 643 1384 647
rect 1564 643 1568 647
rect 1724 643 1728 647
rect 568 635 572 639
rect 188 627 192 631
rect 284 627 288 631
rect 412 627 416 631
rect 540 627 544 631
rect 676 627 680 631
rect 820 627 824 631
rect 964 627 968 631
rect 1108 627 1112 631
rect 1260 627 1264 631
rect 1420 627 1424 631
rect 1580 627 1584 631
rect 1724 627 1728 631
rect 568 603 572 607
rect 1948 523 1952 527
rect 2068 523 2072 527
rect 2196 523 2200 527
rect 2332 523 2336 527
rect 2476 523 2480 527
rect 2620 523 2624 527
rect 2772 523 2776 527
rect 2924 525 2928 529
rect 3084 523 3088 527
rect 3252 523 3256 527
rect 3420 523 3424 527
rect 188 507 192 511
rect 300 507 304 511
rect 460 509 464 513
rect 636 507 640 511
rect 820 507 824 511
rect 1004 507 1008 511
rect 1188 507 1192 511
rect 1372 509 1376 513
rect 1556 507 1560 511
rect 1724 507 1728 511
rect 2188 507 2192 511
rect 2292 509 2296 513
rect 2412 507 2416 511
rect 2540 507 2544 511
rect 2568 507 2572 511
rect 2668 507 2672 511
rect 2804 507 2808 511
rect 2932 507 2936 511
rect 3060 507 3064 511
rect 3188 507 3192 511
rect 3316 507 3320 511
rect 3420 507 3424 511
rect 300 491 304 495
rect 452 491 456 495
rect 620 491 624 495
rect 788 491 792 495
rect 956 491 960 495
rect 1116 491 1120 495
rect 1276 491 1280 495
rect 1428 491 1432 495
rect 1472 491 1476 495
rect 1580 491 1584 495
rect 1724 491 1728 495
rect 2568 483 2572 487
rect 1472 467 1476 471
rect 2292 383 2296 387
rect 2388 385 2392 389
rect 2500 383 2504 387
rect 2612 383 2616 387
rect 2732 383 2736 387
rect 2852 383 2856 387
rect 2964 383 2968 387
rect 3076 383 3080 387
rect 3196 383 3200 387
rect 3316 383 3320 387
rect 3420 383 3424 387
rect 572 373 576 377
rect 668 371 672 375
rect 772 371 776 375
rect 876 371 880 375
rect 980 373 984 377
rect 1076 373 1080 377
rect 1180 371 1184 375
rect 1284 373 1288 377
rect 1388 371 1392 375
rect 1492 371 1496 375
rect 2116 367 2120 371
rect 2204 367 2208 371
rect 2300 367 2304 371
rect 2412 367 2416 371
rect 2532 367 2536 371
rect 2668 367 2672 371
rect 2812 367 2816 371
rect 2964 367 2968 371
rect 3116 367 3120 371
rect 3276 367 3280 371
rect 3420 367 3424 371
rect 524 355 528 359
rect 612 355 616 359
rect 700 355 704 359
rect 728 355 732 359
rect 788 355 792 359
rect 876 355 880 359
rect 964 355 968 359
rect 1052 355 1056 359
rect 1140 355 1144 359
rect 1228 355 1232 359
rect 1316 355 1320 359
rect 728 331 732 335
rect 3248 275 3252 279
rect 1980 247 1984 251
rect 2092 247 2096 251
rect 2220 247 2224 251
rect 2356 247 2360 251
rect 2500 247 2504 251
rect 2652 247 2656 251
rect 2812 247 2816 251
rect 2972 247 2976 251
rect 3140 247 3144 251
rect 332 235 336 239
rect 420 235 424 239
rect 516 235 520 239
rect 612 235 616 239
rect 708 235 712 239
rect 804 237 808 241
rect 900 235 904 239
rect 996 235 1000 239
rect 1100 235 1104 239
rect 1204 235 1208 239
rect 3308 247 3312 251
rect 1884 231 1888 235
rect 1980 231 1984 235
rect 2108 231 2112 235
rect 2252 231 2256 235
rect 2404 231 2408 235
rect 2564 231 2568 235
rect 2732 231 2736 235
rect 2900 231 2904 235
rect 3076 231 3080 235
rect 3248 231 3252 235
rect 3260 231 3264 235
rect 3420 231 3424 235
rect 220 219 224 223
rect 396 219 400 223
rect 564 219 568 223
rect 732 219 736 223
rect 892 221 896 225
rect 1044 219 1048 223
rect 1188 219 1192 223
rect 1332 219 1336 223
rect 1484 219 1488 223
rect 1884 97 1888 101
rect 1972 95 1976 99
rect 2092 95 2096 99
rect 2212 95 2216 99
rect 2332 95 2336 99
rect 2452 95 2456 99
rect 2564 95 2568 99
rect 2676 95 2680 99
rect 2788 95 2792 99
rect 2892 95 2896 99
rect 2996 95 3000 99
rect 3108 95 3112 99
rect 3220 95 3224 99
rect 3332 97 3336 101
rect 3420 95 3424 99
rect 276 79 280 83
rect 364 79 368 83
rect 452 79 456 83
rect 540 79 544 83
rect 628 79 632 83
rect 716 79 720 83
rect 804 79 808 83
rect 900 79 904 83
rect 996 79 1000 83
rect 1084 79 1088 83
rect 1172 79 1176 83
rect 1268 79 1272 83
rect 1364 79 1368 83
rect 1460 79 1464 83
rect 1548 79 1552 83
rect 1636 79 1640 83
rect 1724 79 1728 83
<< m2 >>
rect 1806 3500 1812 3501
rect 3462 3500 3468 3501
rect 1806 3496 1807 3500
rect 1811 3496 1812 3500
rect 1806 3495 1812 3496
rect 2006 3499 2012 3500
rect 2006 3495 2007 3499
rect 2011 3495 2012 3499
rect 2006 3494 2012 3495
rect 2238 3499 2244 3500
rect 2238 3495 2239 3499
rect 2243 3495 2244 3499
rect 2238 3494 2244 3495
rect 2454 3499 2460 3500
rect 2454 3495 2455 3499
rect 2459 3495 2460 3499
rect 2454 3494 2460 3495
rect 2654 3499 2660 3500
rect 2654 3495 2655 3499
rect 2659 3495 2660 3499
rect 2654 3494 2660 3495
rect 2854 3499 2860 3500
rect 2854 3495 2855 3499
rect 2859 3495 2860 3499
rect 2854 3494 2860 3495
rect 3046 3499 3052 3500
rect 3046 3495 3047 3499
rect 3051 3495 3052 3499
rect 3046 3494 3052 3495
rect 3246 3499 3252 3500
rect 3246 3495 3247 3499
rect 3251 3495 3252 3499
rect 3462 3496 3463 3500
rect 3467 3496 3468 3500
rect 3462 3495 3468 3496
rect 3246 3494 3252 3495
rect 2406 3491 2412 3492
rect 2167 3487 2173 3488
rect 2167 3486 2168 3487
rect 2081 3484 2168 3486
rect 1806 3483 1812 3484
rect 1806 3479 1807 3483
rect 1811 3479 1812 3483
rect 2167 3483 2168 3484
rect 2172 3483 2173 3487
rect 2167 3482 2173 3483
rect 2310 3487 2316 3488
rect 2310 3483 2311 3487
rect 2315 3483 2316 3487
rect 2406 3487 2407 3491
rect 2411 3490 2412 3491
rect 2411 3488 2497 3490
rect 2411 3487 2412 3488
rect 2406 3486 2412 3487
rect 2726 3487 2732 3488
rect 2310 3482 2316 3483
rect 2726 3483 2727 3487
rect 2731 3483 2732 3487
rect 2726 3482 2732 3483
rect 2926 3487 2932 3488
rect 2926 3483 2927 3487
rect 2931 3483 2932 3487
rect 2926 3482 2932 3483
rect 3118 3487 3124 3488
rect 3118 3483 3119 3487
rect 3123 3483 3124 3487
rect 3118 3482 3124 3483
rect 3462 3483 3468 3484
rect 1806 3478 1812 3479
rect 2006 3480 2012 3481
rect 2006 3476 2007 3480
rect 2011 3476 2012 3480
rect 2006 3475 2012 3476
rect 2238 3480 2244 3481
rect 2238 3476 2239 3480
rect 2243 3476 2244 3480
rect 2238 3475 2244 3476
rect 2454 3480 2460 3481
rect 2454 3476 2455 3480
rect 2459 3476 2460 3480
rect 2454 3475 2460 3476
rect 2654 3480 2660 3481
rect 2654 3476 2655 3480
rect 2659 3476 2660 3480
rect 2654 3475 2660 3476
rect 2854 3480 2860 3481
rect 2854 3476 2855 3480
rect 2859 3476 2860 3480
rect 2854 3475 2860 3476
rect 3046 3480 3052 3481
rect 3046 3476 3047 3480
rect 3051 3476 3052 3480
rect 3046 3475 3052 3476
rect 3246 3480 3252 3481
rect 3246 3476 3247 3480
rect 3251 3476 3252 3480
rect 3462 3479 3463 3483
rect 3467 3479 3468 3483
rect 3462 3478 3468 3479
rect 3246 3475 3252 3476
rect 2927 3471 2933 3472
rect 2927 3470 2928 3471
rect 2708 3468 2928 3470
rect 2708 3466 2710 3468
rect 2927 3467 2928 3468
rect 2932 3467 2933 3471
rect 2927 3466 2933 3467
rect 2707 3465 2713 3466
rect 110 3464 116 3465
rect 1766 3464 1772 3465
rect 110 3460 111 3464
rect 115 3460 116 3464
rect 110 3459 116 3460
rect 454 3463 460 3464
rect 454 3459 455 3463
rect 459 3459 460 3463
rect 454 3458 460 3459
rect 542 3463 548 3464
rect 542 3459 543 3463
rect 547 3459 548 3463
rect 542 3458 548 3459
rect 630 3463 636 3464
rect 630 3459 631 3463
rect 635 3459 636 3463
rect 630 3458 636 3459
rect 718 3463 724 3464
rect 718 3459 719 3463
rect 723 3459 724 3463
rect 718 3458 724 3459
rect 806 3463 812 3464
rect 806 3459 807 3463
rect 811 3459 812 3463
rect 806 3458 812 3459
rect 894 3463 900 3464
rect 894 3459 895 3463
rect 899 3459 900 3463
rect 894 3458 900 3459
rect 982 3463 988 3464
rect 982 3459 983 3463
rect 987 3459 988 3463
rect 982 3458 988 3459
rect 1070 3463 1076 3464
rect 1070 3459 1071 3463
rect 1075 3459 1076 3463
rect 1070 3458 1076 3459
rect 1158 3463 1164 3464
rect 1158 3459 1159 3463
rect 1163 3459 1164 3463
rect 1766 3460 1767 3464
rect 1771 3460 1772 3464
rect 1766 3459 1772 3460
rect 2014 3463 2020 3464
rect 2014 3459 2015 3463
rect 2019 3462 2020 3463
rect 2059 3463 2065 3464
rect 2059 3462 2060 3463
rect 2019 3460 2060 3462
rect 2019 3459 2020 3460
rect 1158 3458 1164 3459
rect 2014 3458 2020 3459
rect 2059 3459 2060 3460
rect 2064 3459 2065 3463
rect 2059 3458 2065 3459
rect 2167 3463 2173 3464
rect 2167 3459 2168 3463
rect 2172 3462 2173 3463
rect 2291 3463 2297 3464
rect 2291 3462 2292 3463
rect 2172 3460 2292 3462
rect 2172 3459 2173 3460
rect 2167 3458 2173 3459
rect 2291 3459 2292 3460
rect 2296 3459 2297 3463
rect 2291 3458 2297 3459
rect 2310 3463 2316 3464
rect 2310 3459 2311 3463
rect 2315 3462 2316 3463
rect 2507 3463 2513 3464
rect 2507 3462 2508 3463
rect 2315 3460 2508 3462
rect 2315 3459 2316 3460
rect 2310 3458 2316 3459
rect 2507 3459 2508 3460
rect 2512 3459 2513 3463
rect 2707 3461 2708 3465
rect 2712 3461 2713 3465
rect 2707 3460 2713 3461
rect 2726 3463 2732 3464
rect 2507 3458 2513 3459
rect 2726 3459 2727 3463
rect 2731 3462 2732 3463
rect 2907 3463 2913 3464
rect 2907 3462 2908 3463
rect 2731 3460 2908 3462
rect 2731 3459 2732 3460
rect 2726 3458 2732 3459
rect 2907 3459 2908 3460
rect 2912 3459 2913 3463
rect 2907 3458 2913 3459
rect 2926 3463 2932 3464
rect 2926 3459 2927 3463
rect 2931 3462 2932 3463
rect 3099 3463 3105 3464
rect 3099 3462 3100 3463
rect 2931 3460 3100 3462
rect 2931 3459 2932 3460
rect 2926 3458 2932 3459
rect 3099 3459 3100 3460
rect 3104 3459 3105 3463
rect 3099 3458 3105 3459
rect 3118 3463 3124 3464
rect 3118 3459 3119 3463
rect 3123 3462 3124 3463
rect 3299 3463 3305 3464
rect 3299 3462 3300 3463
rect 3123 3460 3300 3462
rect 3123 3459 3124 3460
rect 3118 3458 3124 3459
rect 3299 3459 3300 3460
rect 3304 3459 3305 3463
rect 3299 3458 3305 3459
rect 622 3455 628 3456
rect 526 3451 532 3452
rect 110 3447 116 3448
rect 110 3443 111 3447
rect 115 3443 116 3447
rect 526 3447 527 3451
rect 531 3447 532 3451
rect 526 3446 532 3447
rect 614 3451 620 3452
rect 614 3447 615 3451
rect 619 3447 620 3451
rect 622 3451 623 3455
rect 627 3454 628 3455
rect 710 3455 716 3456
rect 627 3452 673 3454
rect 627 3451 628 3452
rect 622 3450 628 3451
rect 710 3451 711 3455
rect 715 3454 716 3455
rect 798 3455 804 3456
rect 715 3452 761 3454
rect 715 3451 716 3452
rect 710 3450 716 3451
rect 798 3451 799 3455
rect 803 3454 804 3455
rect 886 3455 892 3456
rect 803 3452 849 3454
rect 803 3451 804 3452
rect 798 3450 804 3451
rect 886 3451 887 3455
rect 891 3454 892 3455
rect 974 3455 980 3456
rect 891 3452 937 3454
rect 891 3451 892 3452
rect 886 3450 892 3451
rect 974 3451 975 3455
rect 979 3454 980 3455
rect 1150 3455 1156 3456
rect 979 3452 1025 3454
rect 979 3451 980 3452
rect 974 3450 980 3451
rect 1142 3451 1148 3452
rect 614 3446 620 3447
rect 1142 3447 1143 3451
rect 1147 3447 1148 3451
rect 1150 3451 1151 3455
rect 1155 3454 1156 3455
rect 1155 3452 1201 3454
rect 1155 3451 1156 3452
rect 1150 3450 1156 3451
rect 1883 3451 1889 3452
rect 1142 3446 1148 3447
rect 1766 3447 1772 3448
rect 110 3442 116 3443
rect 454 3444 460 3445
rect 454 3440 455 3444
rect 459 3440 460 3444
rect 454 3439 460 3440
rect 542 3444 548 3445
rect 542 3440 543 3444
rect 547 3440 548 3444
rect 542 3439 548 3440
rect 630 3444 636 3445
rect 630 3440 631 3444
rect 635 3440 636 3444
rect 630 3439 636 3440
rect 718 3444 724 3445
rect 718 3440 719 3444
rect 723 3440 724 3444
rect 718 3439 724 3440
rect 806 3444 812 3445
rect 806 3440 807 3444
rect 811 3440 812 3444
rect 806 3439 812 3440
rect 894 3444 900 3445
rect 894 3440 895 3444
rect 899 3440 900 3444
rect 894 3439 900 3440
rect 982 3444 988 3445
rect 982 3440 983 3444
rect 987 3440 988 3444
rect 982 3439 988 3440
rect 1070 3444 1076 3445
rect 1070 3440 1071 3444
rect 1075 3440 1076 3444
rect 1070 3439 1076 3440
rect 1158 3444 1164 3445
rect 1158 3440 1159 3444
rect 1163 3440 1164 3444
rect 1766 3443 1767 3447
rect 1771 3443 1772 3447
rect 1883 3447 1884 3451
rect 1888 3450 1889 3451
rect 1902 3451 1908 3452
rect 1888 3448 1898 3450
rect 1888 3447 1889 3448
rect 1883 3446 1889 3447
rect 1766 3442 1772 3443
rect 1896 3442 1898 3448
rect 1902 3447 1903 3451
rect 1907 3450 1908 3451
rect 1995 3451 2001 3452
rect 1995 3450 1996 3451
rect 1907 3448 1996 3450
rect 1907 3447 1908 3448
rect 1902 3446 1908 3447
rect 1995 3447 1996 3448
rect 2000 3447 2001 3451
rect 1995 3446 2001 3447
rect 2131 3451 2137 3452
rect 2131 3447 2132 3451
rect 2136 3450 2137 3451
rect 2166 3451 2172 3452
rect 2166 3450 2167 3451
rect 2136 3448 2167 3450
rect 2136 3447 2137 3448
rect 2131 3446 2137 3447
rect 2166 3447 2167 3448
rect 2171 3447 2172 3451
rect 2166 3446 2172 3447
rect 2267 3451 2273 3452
rect 2267 3447 2268 3451
rect 2272 3450 2273 3451
rect 2311 3451 2317 3452
rect 2311 3450 2312 3451
rect 2272 3448 2312 3450
rect 2272 3447 2273 3448
rect 2267 3446 2273 3447
rect 2311 3447 2312 3448
rect 2316 3447 2317 3451
rect 2311 3446 2317 3447
rect 2403 3451 2412 3452
rect 2403 3447 2404 3451
rect 2411 3447 2412 3451
rect 2403 3446 2412 3447
rect 2531 3451 2537 3452
rect 2531 3447 2532 3451
rect 2536 3450 2537 3451
rect 2590 3451 2596 3452
rect 2590 3450 2591 3451
rect 2536 3448 2591 3450
rect 2536 3447 2537 3448
rect 2531 3446 2537 3447
rect 2590 3447 2591 3448
rect 2595 3447 2596 3451
rect 2651 3451 2657 3452
rect 2651 3450 2652 3451
rect 2590 3446 2596 3447
rect 2600 3448 2652 3450
rect 2600 3442 2602 3448
rect 2651 3447 2652 3448
rect 2656 3447 2657 3451
rect 2651 3446 2657 3447
rect 2670 3451 2676 3452
rect 2670 3447 2671 3451
rect 2675 3450 2676 3451
rect 2771 3451 2777 3452
rect 2771 3450 2772 3451
rect 2675 3448 2772 3450
rect 2675 3447 2676 3448
rect 2670 3446 2676 3447
rect 2771 3447 2772 3448
rect 2776 3447 2777 3451
rect 2771 3446 2777 3447
rect 2790 3451 2796 3452
rect 2790 3447 2791 3451
rect 2795 3450 2796 3451
rect 2899 3451 2905 3452
rect 2899 3450 2900 3451
rect 2795 3448 2900 3450
rect 2795 3447 2796 3448
rect 2790 3446 2796 3447
rect 2899 3447 2900 3448
rect 2904 3447 2905 3451
rect 2899 3446 2905 3447
rect 2918 3451 2924 3452
rect 2918 3447 2919 3451
rect 2923 3450 2924 3451
rect 3027 3451 3033 3452
rect 3027 3450 3028 3451
rect 2923 3448 3028 3450
rect 2923 3447 2924 3448
rect 2918 3446 2924 3447
rect 3027 3447 3028 3448
rect 3032 3447 3033 3451
rect 3027 3446 3033 3447
rect 1896 3440 2026 3442
rect 1158 3439 1164 3440
rect 1830 3436 1836 3437
rect 622 3435 628 3436
rect 622 3434 623 3435
rect 508 3432 623 3434
rect 508 3430 510 3432
rect 622 3431 623 3432
rect 627 3431 628 3435
rect 1150 3435 1156 3436
rect 1150 3434 1151 3435
rect 622 3430 628 3431
rect 1036 3432 1151 3434
rect 1036 3430 1038 3432
rect 1150 3431 1151 3432
rect 1155 3431 1156 3435
rect 1150 3430 1156 3431
rect 1806 3433 1812 3434
rect 507 3429 513 3430
rect 507 3425 508 3429
rect 512 3425 513 3429
rect 1035 3429 1041 3430
rect 507 3424 513 3425
rect 526 3427 532 3428
rect 526 3423 527 3427
rect 531 3426 532 3427
rect 595 3427 601 3428
rect 595 3426 596 3427
rect 531 3424 596 3426
rect 531 3423 532 3424
rect 526 3422 532 3423
rect 595 3423 596 3424
rect 600 3423 601 3427
rect 595 3422 601 3423
rect 683 3427 689 3428
rect 683 3423 684 3427
rect 688 3426 689 3427
rect 710 3427 716 3428
rect 710 3426 711 3427
rect 688 3424 711 3426
rect 688 3423 689 3424
rect 683 3422 689 3423
rect 710 3423 711 3424
rect 715 3423 716 3427
rect 710 3422 716 3423
rect 771 3427 777 3428
rect 771 3423 772 3427
rect 776 3426 777 3427
rect 798 3427 804 3428
rect 798 3426 799 3427
rect 776 3424 799 3426
rect 776 3423 777 3424
rect 771 3422 777 3423
rect 798 3423 799 3424
rect 803 3423 804 3427
rect 798 3422 804 3423
rect 859 3427 865 3428
rect 859 3423 860 3427
rect 864 3426 865 3427
rect 886 3427 892 3428
rect 886 3426 887 3427
rect 864 3424 887 3426
rect 864 3423 865 3424
rect 859 3422 865 3423
rect 886 3423 887 3424
rect 891 3423 892 3427
rect 886 3422 892 3423
rect 947 3427 953 3428
rect 947 3423 948 3427
rect 952 3426 953 3427
rect 974 3427 980 3428
rect 974 3426 975 3427
rect 952 3424 975 3426
rect 952 3423 953 3424
rect 947 3422 953 3423
rect 974 3423 975 3424
rect 979 3423 980 3427
rect 1035 3425 1036 3429
rect 1040 3425 1041 3429
rect 1806 3429 1807 3433
rect 1811 3429 1812 3433
rect 1830 3432 1831 3436
rect 1835 3432 1836 3436
rect 1830 3431 1836 3432
rect 1942 3436 1948 3437
rect 1942 3432 1943 3436
rect 1947 3432 1948 3436
rect 1942 3431 1948 3432
rect 1806 3428 1812 3429
rect 1035 3424 1041 3425
rect 1102 3427 1108 3428
rect 974 3422 980 3423
rect 1102 3423 1103 3427
rect 1107 3426 1108 3427
rect 1123 3427 1129 3428
rect 1123 3426 1124 3427
rect 1107 3424 1124 3426
rect 1107 3423 1108 3424
rect 1102 3422 1108 3423
rect 1123 3423 1124 3424
rect 1128 3423 1129 3427
rect 1123 3422 1129 3423
rect 1142 3427 1148 3428
rect 1142 3423 1143 3427
rect 1147 3426 1148 3427
rect 1211 3427 1217 3428
rect 1211 3426 1212 3427
rect 1147 3424 1212 3426
rect 1147 3423 1148 3424
rect 1142 3422 1148 3423
rect 1211 3423 1212 3424
rect 1216 3423 1217 3427
rect 1211 3422 1217 3423
rect 1902 3427 1908 3428
rect 1902 3423 1903 3427
rect 1907 3423 1908 3427
rect 1902 3422 1908 3423
rect 2014 3427 2020 3428
rect 2014 3423 2015 3427
rect 2019 3423 2020 3427
rect 2024 3426 2026 3440
rect 2588 3440 2602 3442
rect 2078 3436 2084 3437
rect 2078 3432 2079 3436
rect 2083 3432 2084 3436
rect 2078 3431 2084 3432
rect 2214 3436 2220 3437
rect 2214 3432 2215 3436
rect 2219 3432 2220 3436
rect 2214 3431 2220 3432
rect 2350 3436 2356 3437
rect 2350 3432 2351 3436
rect 2355 3432 2356 3436
rect 2350 3431 2356 3432
rect 2478 3436 2484 3437
rect 2478 3432 2479 3436
rect 2483 3432 2484 3436
rect 2478 3431 2484 3432
rect 2286 3427 2292 3428
rect 2024 3424 2121 3426
rect 2014 3422 2020 3423
rect 2286 3423 2287 3427
rect 2291 3423 2292 3427
rect 2286 3422 2292 3423
rect 2311 3427 2317 3428
rect 2311 3423 2312 3427
rect 2316 3426 2317 3427
rect 2588 3426 2590 3440
rect 2598 3436 2604 3437
rect 2598 3432 2599 3436
rect 2603 3432 2604 3436
rect 2598 3431 2604 3432
rect 2718 3436 2724 3437
rect 2718 3432 2719 3436
rect 2723 3432 2724 3436
rect 2718 3431 2724 3432
rect 2846 3436 2852 3437
rect 2846 3432 2847 3436
rect 2851 3432 2852 3436
rect 2846 3431 2852 3432
rect 2974 3436 2980 3437
rect 2974 3432 2975 3436
rect 2979 3432 2980 3436
rect 2974 3431 2980 3432
rect 3462 3433 3468 3434
rect 3462 3429 3463 3433
rect 3467 3429 3468 3433
rect 3462 3428 3468 3429
rect 2316 3424 2393 3426
rect 2553 3424 2590 3426
rect 2670 3427 2676 3428
rect 2316 3423 2317 3424
rect 2311 3422 2317 3423
rect 2670 3423 2671 3427
rect 2675 3423 2676 3427
rect 2670 3422 2676 3423
rect 2790 3427 2796 3428
rect 2790 3423 2791 3427
rect 2795 3423 2796 3427
rect 2790 3422 2796 3423
rect 2918 3427 2924 3428
rect 2918 3423 2919 3427
rect 2923 3423 2924 3427
rect 2918 3422 2924 3423
rect 2927 3427 2933 3428
rect 2927 3423 2928 3427
rect 2932 3426 2933 3427
rect 2932 3424 3017 3426
rect 2932 3423 2933 3424
rect 2927 3422 2933 3423
rect 1830 3417 1836 3418
rect 1806 3416 1812 3417
rect 467 3415 473 3416
rect 467 3411 468 3415
rect 472 3414 473 3415
rect 494 3415 500 3416
rect 494 3414 495 3415
rect 472 3412 495 3414
rect 472 3411 473 3412
rect 467 3410 473 3411
rect 494 3411 495 3412
rect 499 3411 500 3415
rect 494 3410 500 3411
rect 555 3415 561 3416
rect 555 3411 556 3415
rect 560 3414 561 3415
rect 614 3415 620 3416
rect 560 3412 610 3414
rect 560 3411 561 3412
rect 555 3410 561 3411
rect 608 3406 610 3412
rect 614 3411 615 3415
rect 619 3414 620 3415
rect 643 3415 649 3416
rect 643 3414 644 3415
rect 619 3412 644 3414
rect 619 3411 620 3412
rect 614 3410 620 3411
rect 643 3411 644 3412
rect 648 3411 649 3415
rect 643 3410 649 3411
rect 662 3415 668 3416
rect 662 3411 663 3415
rect 667 3414 668 3415
rect 731 3415 737 3416
rect 731 3414 732 3415
rect 667 3412 732 3414
rect 667 3411 668 3412
rect 662 3410 668 3411
rect 731 3411 732 3412
rect 736 3411 737 3415
rect 731 3410 737 3411
rect 750 3415 756 3416
rect 750 3411 751 3415
rect 755 3414 756 3415
rect 819 3415 825 3416
rect 819 3414 820 3415
rect 755 3412 820 3414
rect 755 3411 756 3412
rect 750 3410 756 3411
rect 819 3411 820 3412
rect 824 3411 825 3415
rect 819 3410 825 3411
rect 907 3415 913 3416
rect 907 3411 908 3415
rect 912 3414 913 3415
rect 926 3415 932 3416
rect 912 3412 922 3414
rect 912 3411 913 3412
rect 907 3410 913 3411
rect 920 3406 922 3412
rect 926 3411 927 3415
rect 931 3414 932 3415
rect 995 3415 1001 3416
rect 995 3414 996 3415
rect 931 3412 996 3414
rect 931 3411 932 3412
rect 926 3410 932 3411
rect 995 3411 996 3412
rect 1000 3411 1001 3415
rect 995 3410 1001 3411
rect 1014 3415 1020 3416
rect 1014 3411 1015 3415
rect 1019 3414 1020 3415
rect 1083 3415 1089 3416
rect 1083 3414 1084 3415
rect 1019 3412 1084 3414
rect 1019 3411 1020 3412
rect 1014 3410 1020 3411
rect 1083 3411 1084 3412
rect 1088 3411 1089 3415
rect 1083 3410 1089 3411
rect 1171 3415 1177 3416
rect 1171 3411 1172 3415
rect 1176 3414 1177 3415
rect 1258 3415 1265 3416
rect 1176 3412 1254 3414
rect 1176 3411 1177 3412
rect 1171 3410 1177 3411
rect 1252 3406 1254 3412
rect 1258 3411 1259 3415
rect 1264 3411 1265 3415
rect 1258 3410 1265 3411
rect 1278 3415 1284 3416
rect 1278 3411 1279 3415
rect 1283 3414 1284 3415
rect 1355 3415 1361 3416
rect 1355 3414 1356 3415
rect 1283 3412 1356 3414
rect 1283 3411 1284 3412
rect 1278 3410 1284 3411
rect 1355 3411 1356 3412
rect 1360 3411 1361 3415
rect 1806 3412 1807 3416
rect 1811 3412 1812 3416
rect 1830 3413 1831 3417
rect 1835 3413 1836 3417
rect 1830 3412 1836 3413
rect 1942 3417 1948 3418
rect 1942 3413 1943 3417
rect 1947 3413 1948 3417
rect 1942 3412 1948 3413
rect 2078 3417 2084 3418
rect 2078 3413 2079 3417
rect 2083 3413 2084 3417
rect 2078 3412 2084 3413
rect 2214 3417 2220 3418
rect 2214 3413 2215 3417
rect 2219 3413 2220 3417
rect 2214 3412 2220 3413
rect 2350 3417 2356 3418
rect 2350 3413 2351 3417
rect 2355 3413 2356 3417
rect 2350 3412 2356 3413
rect 2478 3417 2484 3418
rect 2478 3413 2479 3417
rect 2483 3413 2484 3417
rect 2478 3412 2484 3413
rect 2598 3417 2604 3418
rect 2598 3413 2599 3417
rect 2603 3413 2604 3417
rect 2598 3412 2604 3413
rect 2718 3417 2724 3418
rect 2718 3413 2719 3417
rect 2723 3413 2724 3417
rect 2718 3412 2724 3413
rect 2846 3417 2852 3418
rect 2846 3413 2847 3417
rect 2851 3413 2852 3417
rect 2846 3412 2852 3413
rect 2974 3417 2980 3418
rect 2974 3413 2975 3417
rect 2979 3413 2980 3417
rect 2974 3412 2980 3413
rect 3462 3416 3468 3417
rect 3462 3412 3463 3416
rect 3467 3412 3468 3416
rect 1806 3411 1812 3412
rect 3462 3411 3468 3412
rect 1355 3410 1361 3411
rect 608 3404 762 3406
rect 920 3404 1114 3406
rect 1252 3404 1290 3406
rect 414 3400 420 3401
rect 110 3397 116 3398
rect 110 3393 111 3397
rect 115 3393 116 3397
rect 414 3396 415 3400
rect 419 3396 420 3400
rect 414 3395 420 3396
rect 502 3400 508 3401
rect 502 3396 503 3400
rect 507 3396 508 3400
rect 502 3395 508 3396
rect 590 3400 596 3401
rect 590 3396 591 3400
rect 595 3396 596 3400
rect 590 3395 596 3396
rect 678 3400 684 3401
rect 678 3396 679 3400
rect 683 3396 684 3400
rect 678 3395 684 3396
rect 110 3392 116 3393
rect 478 3391 484 3392
rect 478 3387 479 3391
rect 483 3387 484 3391
rect 478 3386 484 3387
rect 494 3391 500 3392
rect 494 3387 495 3391
rect 499 3390 500 3391
rect 662 3391 668 3392
rect 499 3388 545 3390
rect 499 3387 500 3388
rect 494 3386 500 3387
rect 662 3387 663 3391
rect 667 3387 668 3391
rect 662 3386 668 3387
rect 750 3391 756 3392
rect 750 3387 751 3391
rect 755 3387 756 3391
rect 760 3390 762 3404
rect 766 3400 772 3401
rect 766 3396 767 3400
rect 771 3396 772 3400
rect 766 3395 772 3396
rect 854 3400 860 3401
rect 854 3396 855 3400
rect 859 3396 860 3400
rect 854 3395 860 3396
rect 942 3400 948 3401
rect 942 3396 943 3400
rect 947 3396 948 3400
rect 942 3395 948 3396
rect 1030 3400 1036 3401
rect 1030 3396 1031 3400
rect 1035 3396 1036 3400
rect 1030 3395 1036 3396
rect 926 3391 932 3392
rect 760 3388 809 3390
rect 750 3386 756 3387
rect 926 3387 927 3391
rect 931 3387 932 3391
rect 926 3386 932 3387
rect 1014 3391 1020 3392
rect 1014 3387 1015 3391
rect 1019 3387 1020 3391
rect 1014 3386 1020 3387
rect 1102 3391 1108 3392
rect 1102 3387 1103 3391
rect 1107 3387 1108 3391
rect 1112 3390 1114 3404
rect 1118 3400 1124 3401
rect 1118 3396 1119 3400
rect 1123 3396 1124 3400
rect 1118 3395 1124 3396
rect 1206 3400 1212 3401
rect 1206 3396 1207 3400
rect 1211 3396 1212 3400
rect 1206 3395 1212 3396
rect 1278 3391 1284 3392
rect 1112 3388 1161 3390
rect 1102 3386 1108 3387
rect 1278 3387 1279 3391
rect 1283 3387 1284 3391
rect 1288 3390 1290 3404
rect 1302 3400 1308 3401
rect 1302 3396 1303 3400
rect 1307 3396 1308 3400
rect 1302 3395 1308 3396
rect 1766 3397 1772 3398
rect 1766 3393 1767 3397
rect 1771 3393 1772 3397
rect 1766 3392 1772 3393
rect 1288 3388 1345 3390
rect 1278 3386 1284 3387
rect 414 3381 420 3382
rect 110 3380 116 3381
rect 110 3376 111 3380
rect 115 3376 116 3380
rect 414 3377 415 3381
rect 419 3377 420 3381
rect 414 3376 420 3377
rect 502 3381 508 3382
rect 502 3377 503 3381
rect 507 3377 508 3381
rect 502 3376 508 3377
rect 590 3381 596 3382
rect 590 3377 591 3381
rect 595 3377 596 3381
rect 590 3376 596 3377
rect 678 3381 684 3382
rect 678 3377 679 3381
rect 683 3377 684 3381
rect 678 3376 684 3377
rect 766 3381 772 3382
rect 766 3377 767 3381
rect 771 3377 772 3381
rect 766 3376 772 3377
rect 854 3381 860 3382
rect 854 3377 855 3381
rect 859 3377 860 3381
rect 854 3376 860 3377
rect 942 3381 948 3382
rect 942 3377 943 3381
rect 947 3377 948 3381
rect 942 3376 948 3377
rect 1030 3381 1036 3382
rect 1030 3377 1031 3381
rect 1035 3377 1036 3381
rect 1030 3376 1036 3377
rect 1118 3381 1124 3382
rect 1118 3377 1119 3381
rect 1123 3377 1124 3381
rect 1118 3376 1124 3377
rect 1206 3381 1212 3382
rect 1206 3377 1207 3381
rect 1211 3377 1212 3381
rect 1206 3376 1212 3377
rect 1302 3381 1308 3382
rect 1302 3377 1303 3381
rect 1307 3377 1308 3381
rect 1302 3376 1308 3377
rect 1766 3380 1772 3381
rect 1766 3376 1767 3380
rect 1771 3376 1772 3380
rect 110 3375 116 3376
rect 1766 3375 1772 3376
rect 1806 3364 1812 3365
rect 3462 3364 3468 3365
rect 1806 3360 1807 3364
rect 1811 3360 1812 3364
rect 1806 3359 1812 3360
rect 1830 3363 1836 3364
rect 1830 3359 1831 3363
rect 1835 3359 1836 3363
rect 1830 3358 1836 3359
rect 1950 3363 1956 3364
rect 1950 3359 1951 3363
rect 1955 3359 1956 3363
rect 1950 3358 1956 3359
rect 2094 3363 2100 3364
rect 2094 3359 2095 3363
rect 2099 3359 2100 3363
rect 2094 3358 2100 3359
rect 2238 3363 2244 3364
rect 2238 3359 2239 3363
rect 2243 3359 2244 3363
rect 2238 3358 2244 3359
rect 2382 3363 2388 3364
rect 2382 3359 2383 3363
rect 2387 3359 2388 3363
rect 2382 3358 2388 3359
rect 2518 3363 2524 3364
rect 2518 3359 2519 3363
rect 2523 3359 2524 3363
rect 2518 3358 2524 3359
rect 2646 3363 2652 3364
rect 2646 3359 2647 3363
rect 2651 3359 2652 3363
rect 2646 3358 2652 3359
rect 2774 3363 2780 3364
rect 2774 3359 2775 3363
rect 2779 3359 2780 3363
rect 2774 3358 2780 3359
rect 2902 3363 2908 3364
rect 2902 3359 2903 3363
rect 2907 3359 2908 3363
rect 2902 3358 2908 3359
rect 3038 3363 3044 3364
rect 3038 3359 3039 3363
rect 3043 3359 3044 3363
rect 3462 3360 3463 3364
rect 3467 3360 3468 3364
rect 3462 3359 3468 3360
rect 3038 3358 3044 3359
rect 2166 3355 2172 3356
rect 1902 3351 1908 3352
rect 1190 3347 1196 3348
rect 1190 3343 1191 3347
rect 1195 3346 1196 3347
rect 1258 3347 1264 3348
rect 1258 3346 1259 3347
rect 1195 3344 1259 3346
rect 1195 3343 1196 3344
rect 1190 3342 1196 3343
rect 1258 3343 1259 3344
rect 1263 3343 1264 3347
rect 1258 3342 1264 3343
rect 1806 3347 1812 3348
rect 1806 3343 1807 3347
rect 1811 3343 1812 3347
rect 1902 3347 1903 3351
rect 1907 3347 1908 3351
rect 1902 3346 1908 3347
rect 2022 3351 2028 3352
rect 2022 3347 2023 3351
rect 2027 3347 2028 3351
rect 2166 3351 2167 3355
rect 2171 3351 2172 3355
rect 2590 3355 2596 3356
rect 2166 3350 2172 3351
rect 2310 3351 2316 3352
rect 2022 3346 2028 3347
rect 2310 3347 2311 3351
rect 2315 3347 2316 3351
rect 2310 3346 2316 3347
rect 2454 3351 2460 3352
rect 2454 3347 2455 3351
rect 2459 3347 2460 3351
rect 2590 3351 2591 3355
rect 2595 3351 2596 3355
rect 2590 3350 2596 3351
rect 2598 3355 2604 3356
rect 2598 3351 2599 3355
rect 2603 3354 2604 3355
rect 2726 3355 2732 3356
rect 2603 3352 2689 3354
rect 2603 3351 2604 3352
rect 2598 3350 2604 3351
rect 2726 3351 2727 3355
rect 2731 3354 2732 3355
rect 2982 3355 2988 3356
rect 2731 3352 2817 3354
rect 2731 3351 2732 3352
rect 2726 3350 2732 3351
rect 2974 3351 2980 3352
rect 2454 3346 2460 3347
rect 2974 3347 2975 3351
rect 2979 3347 2980 3351
rect 2982 3351 2983 3355
rect 2987 3354 2988 3355
rect 2987 3352 3081 3354
rect 2987 3351 2988 3352
rect 2982 3350 2988 3351
rect 2974 3346 2980 3347
rect 3462 3347 3468 3348
rect 1806 3342 1812 3343
rect 1830 3344 1836 3345
rect 1830 3340 1831 3344
rect 1835 3340 1836 3344
rect 1830 3339 1836 3340
rect 1950 3344 1956 3345
rect 1950 3340 1951 3344
rect 1955 3340 1956 3344
rect 1950 3339 1956 3340
rect 2094 3344 2100 3345
rect 2094 3340 2095 3344
rect 2099 3340 2100 3344
rect 2094 3339 2100 3340
rect 2238 3344 2244 3345
rect 2238 3340 2239 3344
rect 2243 3340 2244 3344
rect 2238 3339 2244 3340
rect 2382 3344 2388 3345
rect 2382 3340 2383 3344
rect 2387 3340 2388 3344
rect 2382 3339 2388 3340
rect 2518 3344 2524 3345
rect 2518 3340 2519 3344
rect 2523 3340 2524 3344
rect 2518 3339 2524 3340
rect 2646 3344 2652 3345
rect 2646 3340 2647 3344
rect 2651 3340 2652 3344
rect 2646 3339 2652 3340
rect 2774 3344 2780 3345
rect 2774 3340 2775 3344
rect 2779 3340 2780 3344
rect 2774 3339 2780 3340
rect 2902 3344 2908 3345
rect 2902 3340 2903 3344
rect 2907 3340 2908 3344
rect 2902 3339 2908 3340
rect 3038 3344 3044 3345
rect 3038 3340 3039 3344
rect 3043 3340 3044 3344
rect 3462 3343 3463 3347
rect 3467 3343 3468 3347
rect 3462 3342 3468 3343
rect 3038 3339 3044 3340
rect 2982 3335 2988 3336
rect 2982 3334 2983 3335
rect 110 3332 116 3333
rect 1766 3332 1772 3333
rect 110 3328 111 3332
rect 115 3328 116 3332
rect 110 3327 116 3328
rect 398 3331 404 3332
rect 398 3327 399 3331
rect 403 3327 404 3331
rect 398 3326 404 3327
rect 494 3331 500 3332
rect 494 3327 495 3331
rect 499 3327 500 3331
rect 494 3326 500 3327
rect 598 3331 604 3332
rect 598 3327 599 3331
rect 603 3327 604 3331
rect 598 3326 604 3327
rect 702 3331 708 3332
rect 702 3327 703 3331
rect 707 3327 708 3331
rect 702 3326 708 3327
rect 806 3331 812 3332
rect 806 3327 807 3331
rect 811 3327 812 3331
rect 806 3326 812 3327
rect 910 3331 916 3332
rect 910 3327 911 3331
rect 915 3327 916 3331
rect 910 3326 916 3327
rect 1014 3331 1020 3332
rect 1014 3327 1015 3331
rect 1019 3327 1020 3331
rect 1014 3326 1020 3327
rect 1118 3331 1124 3332
rect 1118 3327 1119 3331
rect 1123 3327 1124 3331
rect 1118 3326 1124 3327
rect 1222 3331 1228 3332
rect 1222 3327 1223 3331
rect 1227 3327 1228 3331
rect 1222 3326 1228 3327
rect 1326 3331 1332 3332
rect 1326 3327 1327 3331
rect 1331 3327 1332 3331
rect 1766 3328 1767 3332
rect 1771 3328 1772 3332
rect 2828 3332 2983 3334
rect 2828 3330 2830 3332
rect 2982 3331 2983 3332
rect 2987 3331 2988 3335
rect 2982 3330 2988 3331
rect 2827 3329 2833 3330
rect 1766 3327 1772 3328
rect 1883 3327 1889 3328
rect 1326 3326 1332 3327
rect 1190 3323 1196 3324
rect 486 3319 492 3320
rect 486 3318 487 3319
rect 473 3316 487 3318
rect 110 3315 116 3316
rect 110 3311 111 3315
rect 115 3311 116 3315
rect 486 3315 487 3316
rect 491 3315 492 3319
rect 486 3314 492 3315
rect 566 3319 572 3320
rect 566 3315 567 3319
rect 571 3315 572 3319
rect 566 3314 572 3315
rect 670 3319 676 3320
rect 670 3315 671 3319
rect 675 3315 676 3319
rect 670 3314 676 3315
rect 774 3319 780 3320
rect 774 3315 775 3319
rect 779 3315 780 3319
rect 774 3314 780 3315
rect 878 3319 884 3320
rect 878 3315 879 3319
rect 883 3315 884 3319
rect 878 3314 884 3315
rect 982 3319 988 3320
rect 982 3315 983 3319
rect 987 3315 988 3319
rect 982 3314 988 3315
rect 1086 3319 1092 3320
rect 1086 3315 1087 3319
rect 1091 3315 1092 3319
rect 1190 3319 1191 3323
rect 1195 3319 1196 3323
rect 1190 3318 1196 3319
rect 1198 3323 1204 3324
rect 1198 3319 1199 3323
rect 1203 3322 1204 3323
rect 1302 3323 1308 3324
rect 1203 3320 1265 3322
rect 1203 3319 1204 3320
rect 1198 3318 1204 3319
rect 1302 3319 1303 3323
rect 1307 3322 1308 3323
rect 1883 3323 1884 3327
rect 1888 3326 1889 3327
rect 1894 3327 1900 3328
rect 1894 3326 1895 3327
rect 1888 3324 1895 3326
rect 1888 3323 1889 3324
rect 1883 3322 1889 3323
rect 1894 3323 1895 3324
rect 1899 3323 1900 3327
rect 1894 3322 1900 3323
rect 1902 3327 1908 3328
rect 1902 3323 1903 3327
rect 1907 3326 1908 3327
rect 2003 3327 2009 3328
rect 2003 3326 2004 3327
rect 1907 3324 2004 3326
rect 1907 3323 1908 3324
rect 1902 3322 1908 3323
rect 2003 3323 2004 3324
rect 2008 3323 2009 3327
rect 2003 3322 2009 3323
rect 2022 3327 2028 3328
rect 2022 3323 2023 3327
rect 2027 3326 2028 3327
rect 2147 3327 2153 3328
rect 2147 3326 2148 3327
rect 2027 3324 2148 3326
rect 2027 3323 2028 3324
rect 2022 3322 2028 3323
rect 2147 3323 2148 3324
rect 2152 3323 2153 3327
rect 2147 3322 2153 3323
rect 2286 3327 2297 3328
rect 2286 3323 2287 3327
rect 2291 3323 2292 3327
rect 2296 3323 2297 3327
rect 2286 3322 2297 3323
rect 2310 3327 2316 3328
rect 2310 3323 2311 3327
rect 2315 3326 2316 3327
rect 2435 3327 2441 3328
rect 2435 3326 2436 3327
rect 2315 3324 2436 3326
rect 2315 3323 2316 3324
rect 2310 3322 2316 3323
rect 2435 3323 2436 3324
rect 2440 3323 2441 3327
rect 2435 3322 2441 3323
rect 2571 3327 2577 3328
rect 2571 3323 2572 3327
rect 2576 3326 2577 3327
rect 2598 3327 2604 3328
rect 2598 3326 2599 3327
rect 2576 3324 2599 3326
rect 2576 3323 2577 3324
rect 2571 3322 2577 3323
rect 2598 3323 2599 3324
rect 2603 3323 2604 3327
rect 2598 3322 2604 3323
rect 2699 3327 2705 3328
rect 2699 3323 2700 3327
rect 2704 3326 2705 3327
rect 2726 3327 2732 3328
rect 2726 3326 2727 3327
rect 2704 3324 2727 3326
rect 2704 3323 2705 3324
rect 2699 3322 2705 3323
rect 2726 3323 2727 3324
rect 2731 3323 2732 3327
rect 2827 3325 2828 3329
rect 2832 3325 2833 3329
rect 2827 3324 2833 3325
rect 2911 3327 2917 3328
rect 2726 3322 2732 3323
rect 2911 3323 2912 3327
rect 2916 3326 2917 3327
rect 2955 3327 2961 3328
rect 2955 3326 2956 3327
rect 2916 3324 2956 3326
rect 2916 3323 2917 3324
rect 2911 3322 2917 3323
rect 2955 3323 2956 3324
rect 2960 3323 2961 3327
rect 2955 3322 2961 3323
rect 2974 3327 2980 3328
rect 2974 3323 2975 3327
rect 2979 3326 2980 3327
rect 3091 3327 3097 3328
rect 3091 3326 3092 3327
rect 2979 3324 3092 3326
rect 2979 3323 2980 3324
rect 2974 3322 2980 3323
rect 3091 3323 3092 3324
rect 3096 3323 3097 3327
rect 3091 3322 3097 3323
rect 1307 3320 1369 3322
rect 1307 3319 1308 3320
rect 1302 3318 1308 3319
rect 1086 3314 1092 3315
rect 1766 3315 1772 3316
rect 110 3310 116 3311
rect 398 3312 404 3313
rect 398 3308 399 3312
rect 403 3308 404 3312
rect 398 3307 404 3308
rect 494 3312 500 3313
rect 494 3308 495 3312
rect 499 3308 500 3312
rect 494 3307 500 3308
rect 598 3312 604 3313
rect 598 3308 599 3312
rect 603 3308 604 3312
rect 598 3307 604 3308
rect 702 3312 708 3313
rect 702 3308 703 3312
rect 707 3308 708 3312
rect 702 3307 708 3308
rect 806 3312 812 3313
rect 806 3308 807 3312
rect 811 3308 812 3312
rect 806 3307 812 3308
rect 910 3312 916 3313
rect 910 3308 911 3312
rect 915 3308 916 3312
rect 910 3307 916 3308
rect 1014 3312 1020 3313
rect 1014 3308 1015 3312
rect 1019 3308 1020 3312
rect 1014 3307 1020 3308
rect 1118 3312 1124 3313
rect 1118 3308 1119 3312
rect 1123 3308 1124 3312
rect 1118 3307 1124 3308
rect 1222 3312 1228 3313
rect 1222 3308 1223 3312
rect 1227 3308 1228 3312
rect 1222 3307 1228 3308
rect 1326 3312 1332 3313
rect 1326 3308 1327 3312
rect 1331 3308 1332 3312
rect 1766 3311 1767 3315
rect 1771 3311 1772 3315
rect 1766 3310 1772 3311
rect 1326 3307 1332 3308
rect 1883 3307 1889 3308
rect 1198 3303 1204 3304
rect 1198 3302 1199 3303
rect 964 3300 1199 3302
rect 964 3298 966 3300
rect 1198 3299 1199 3300
rect 1203 3299 1204 3303
rect 1883 3303 1884 3307
rect 1888 3306 1889 3307
rect 1910 3307 1916 3308
rect 1910 3306 1911 3307
rect 1888 3304 1911 3306
rect 1888 3303 1889 3304
rect 1883 3302 1889 3303
rect 1910 3303 1911 3304
rect 1915 3303 1916 3307
rect 1910 3302 1916 3303
rect 2027 3307 2033 3308
rect 2027 3303 2028 3307
rect 2032 3306 2033 3307
rect 2054 3307 2060 3308
rect 2054 3306 2055 3307
rect 2032 3304 2055 3306
rect 2032 3303 2033 3304
rect 2027 3302 2033 3303
rect 2054 3303 2055 3304
rect 2059 3303 2060 3307
rect 2054 3302 2060 3303
rect 2102 3307 2108 3308
rect 2102 3303 2103 3307
rect 2107 3306 2108 3307
rect 2203 3307 2209 3308
rect 2203 3306 2204 3307
rect 2107 3304 2204 3306
rect 2107 3303 2108 3304
rect 2102 3302 2108 3303
rect 2203 3303 2204 3304
rect 2208 3303 2209 3307
rect 2203 3302 2209 3303
rect 2387 3307 2393 3308
rect 2387 3303 2388 3307
rect 2392 3306 2393 3307
rect 2414 3307 2420 3308
rect 2414 3306 2415 3307
rect 2392 3304 2415 3306
rect 2392 3303 2393 3304
rect 2387 3302 2393 3303
rect 2414 3303 2415 3304
rect 2419 3303 2420 3307
rect 2414 3302 2420 3303
rect 2454 3307 2460 3308
rect 2454 3303 2455 3307
rect 2459 3306 2460 3307
rect 2563 3307 2569 3308
rect 2563 3306 2564 3307
rect 2459 3304 2564 3306
rect 2459 3303 2460 3304
rect 2454 3302 2460 3303
rect 2563 3303 2564 3304
rect 2568 3303 2569 3307
rect 2563 3302 2569 3303
rect 2731 3307 2737 3308
rect 2731 3303 2732 3307
rect 2736 3306 2737 3307
rect 2750 3307 2756 3308
rect 2736 3304 2746 3306
rect 2736 3303 2737 3304
rect 2731 3302 2737 3303
rect 1198 3298 1204 3299
rect 2744 3298 2746 3304
rect 2750 3303 2751 3307
rect 2755 3306 2756 3307
rect 2883 3307 2889 3308
rect 2883 3306 2884 3307
rect 2755 3304 2884 3306
rect 2755 3303 2756 3304
rect 2750 3302 2756 3303
rect 2883 3303 2884 3304
rect 2888 3303 2889 3307
rect 2883 3302 2889 3303
rect 3027 3307 3033 3308
rect 3027 3303 3028 3307
rect 3032 3306 3033 3307
rect 3054 3307 3060 3308
rect 3054 3306 3055 3307
rect 3032 3304 3055 3306
rect 3032 3303 3033 3304
rect 3027 3302 3033 3303
rect 3054 3303 3055 3304
rect 3059 3303 3060 3307
rect 3054 3302 3060 3303
rect 3163 3307 3169 3308
rect 3163 3303 3164 3307
rect 3168 3306 3169 3307
rect 3191 3307 3197 3308
rect 3191 3306 3192 3307
rect 3168 3304 3192 3306
rect 3168 3303 3169 3304
rect 3163 3302 3169 3303
rect 3191 3303 3192 3304
rect 3196 3303 3197 3307
rect 3191 3302 3197 3303
rect 3299 3307 3305 3308
rect 3299 3303 3300 3307
rect 3304 3306 3305 3307
rect 3326 3307 3332 3308
rect 3326 3306 3327 3307
rect 3304 3304 3327 3306
rect 3304 3303 3305 3304
rect 3299 3302 3305 3303
rect 3326 3303 3327 3304
rect 3331 3303 3332 3307
rect 3326 3302 3332 3303
rect 3419 3307 3425 3308
rect 3419 3303 3420 3307
rect 3424 3306 3425 3307
rect 3438 3307 3444 3308
rect 3438 3306 3439 3307
rect 3424 3304 3439 3306
rect 3424 3303 3425 3304
rect 3419 3302 3425 3303
rect 3438 3303 3439 3304
rect 3443 3303 3444 3307
rect 3438 3302 3444 3303
rect 963 3297 969 3298
rect 451 3295 457 3296
rect 451 3291 452 3295
rect 456 3294 457 3295
rect 478 3295 484 3296
rect 478 3294 479 3295
rect 456 3292 479 3294
rect 456 3291 457 3292
rect 451 3290 457 3291
rect 478 3291 479 3292
rect 483 3291 484 3295
rect 478 3290 484 3291
rect 486 3295 492 3296
rect 486 3291 487 3295
rect 491 3294 492 3295
rect 547 3295 553 3296
rect 547 3294 548 3295
rect 491 3292 548 3294
rect 491 3291 492 3292
rect 486 3290 492 3291
rect 547 3291 548 3292
rect 552 3291 553 3295
rect 547 3290 553 3291
rect 566 3295 572 3296
rect 566 3291 567 3295
rect 571 3294 572 3295
rect 651 3295 657 3296
rect 651 3294 652 3295
rect 571 3292 652 3294
rect 571 3291 572 3292
rect 566 3290 572 3291
rect 651 3291 652 3292
rect 656 3291 657 3295
rect 651 3290 657 3291
rect 670 3295 676 3296
rect 670 3291 671 3295
rect 675 3294 676 3295
rect 755 3295 761 3296
rect 755 3294 756 3295
rect 675 3292 756 3294
rect 675 3291 676 3292
rect 670 3290 676 3291
rect 755 3291 756 3292
rect 760 3291 761 3295
rect 755 3290 761 3291
rect 774 3295 780 3296
rect 774 3291 775 3295
rect 779 3294 780 3295
rect 859 3295 865 3296
rect 859 3294 860 3295
rect 779 3292 860 3294
rect 779 3291 780 3292
rect 774 3290 780 3291
rect 859 3291 860 3292
rect 864 3291 865 3295
rect 963 3293 964 3297
rect 968 3293 969 3297
rect 2744 3296 2922 3298
rect 963 3292 969 3293
rect 982 3295 988 3296
rect 859 3290 865 3291
rect 982 3291 983 3295
rect 987 3294 988 3295
rect 1067 3295 1073 3296
rect 1067 3294 1068 3295
rect 987 3292 1068 3294
rect 987 3291 988 3292
rect 982 3290 988 3291
rect 1067 3291 1068 3292
rect 1072 3291 1073 3295
rect 1067 3290 1073 3291
rect 1086 3295 1092 3296
rect 1086 3291 1087 3295
rect 1091 3294 1092 3295
rect 1171 3295 1177 3296
rect 1171 3294 1172 3295
rect 1091 3292 1172 3294
rect 1091 3291 1092 3292
rect 1086 3290 1092 3291
rect 1171 3291 1172 3292
rect 1176 3291 1177 3295
rect 1171 3290 1177 3291
rect 1275 3295 1281 3296
rect 1275 3291 1276 3295
rect 1280 3294 1281 3295
rect 1302 3295 1308 3296
rect 1302 3294 1303 3295
rect 1280 3292 1303 3294
rect 1280 3291 1281 3292
rect 1275 3290 1281 3291
rect 1302 3291 1303 3292
rect 1307 3291 1308 3295
rect 1302 3290 1308 3291
rect 1379 3295 1385 3296
rect 1379 3291 1380 3295
rect 1384 3294 1385 3295
rect 1398 3295 1404 3296
rect 1398 3294 1399 3295
rect 1384 3292 1399 3294
rect 1384 3291 1385 3292
rect 1379 3290 1385 3291
rect 1398 3291 1399 3292
rect 1403 3291 1404 3295
rect 1398 3290 1404 3291
rect 1830 3292 1836 3293
rect 1806 3289 1812 3290
rect 1806 3285 1807 3289
rect 1811 3285 1812 3289
rect 1830 3288 1831 3292
rect 1835 3288 1836 3292
rect 1830 3287 1836 3288
rect 1974 3292 1980 3293
rect 1974 3288 1975 3292
rect 1979 3288 1980 3292
rect 1974 3287 1980 3288
rect 2150 3292 2156 3293
rect 2150 3288 2151 3292
rect 2155 3288 2156 3292
rect 2150 3287 2156 3288
rect 2334 3292 2340 3293
rect 2334 3288 2335 3292
rect 2339 3288 2340 3292
rect 2334 3287 2340 3288
rect 2510 3292 2516 3293
rect 2510 3288 2511 3292
rect 2515 3288 2516 3292
rect 2510 3287 2516 3288
rect 2678 3292 2684 3293
rect 2678 3288 2679 3292
rect 2683 3288 2684 3292
rect 2678 3287 2684 3288
rect 2830 3292 2836 3293
rect 2830 3288 2831 3292
rect 2835 3288 2836 3292
rect 2830 3287 2836 3288
rect 1806 3284 1812 3285
rect 1894 3283 1900 3284
rect 435 3279 441 3280
rect 435 3275 436 3279
rect 440 3278 441 3279
rect 454 3279 460 3280
rect 440 3276 450 3278
rect 440 3275 441 3276
rect 435 3274 441 3275
rect 448 3270 450 3276
rect 454 3275 455 3279
rect 459 3278 460 3279
rect 547 3279 553 3280
rect 547 3278 548 3279
rect 459 3276 548 3278
rect 459 3275 460 3276
rect 454 3274 460 3275
rect 547 3275 548 3276
rect 552 3275 553 3279
rect 547 3274 553 3275
rect 659 3279 665 3280
rect 659 3275 660 3279
rect 664 3278 665 3279
rect 694 3279 700 3280
rect 694 3278 695 3279
rect 664 3276 695 3278
rect 664 3275 665 3276
rect 659 3274 665 3275
rect 694 3275 695 3276
rect 699 3275 700 3279
rect 694 3274 700 3275
rect 779 3279 785 3280
rect 779 3275 780 3279
rect 784 3278 785 3279
rect 807 3279 813 3280
rect 807 3278 808 3279
rect 784 3276 808 3278
rect 784 3275 785 3276
rect 779 3274 785 3275
rect 807 3275 808 3276
rect 812 3275 813 3279
rect 807 3274 813 3275
rect 878 3279 884 3280
rect 878 3275 879 3279
rect 883 3278 884 3279
rect 899 3279 905 3280
rect 899 3278 900 3279
rect 883 3276 900 3278
rect 883 3275 884 3276
rect 878 3274 884 3275
rect 899 3275 900 3276
rect 904 3275 905 3279
rect 899 3274 905 3275
rect 998 3279 1004 3280
rect 998 3275 999 3279
rect 1003 3278 1004 3279
rect 1019 3279 1025 3280
rect 1019 3278 1020 3279
rect 1003 3276 1020 3278
rect 1003 3275 1004 3276
rect 998 3274 1004 3275
rect 1019 3275 1020 3276
rect 1024 3275 1025 3279
rect 1019 3274 1025 3275
rect 1038 3279 1044 3280
rect 1038 3275 1039 3279
rect 1043 3278 1044 3279
rect 1139 3279 1145 3280
rect 1139 3278 1140 3279
rect 1043 3276 1140 3278
rect 1043 3275 1044 3276
rect 1038 3274 1044 3275
rect 1139 3275 1140 3276
rect 1144 3275 1145 3279
rect 1139 3274 1145 3275
rect 1158 3279 1164 3280
rect 1158 3275 1159 3279
rect 1163 3278 1164 3279
rect 1259 3279 1265 3280
rect 1259 3278 1260 3279
rect 1163 3276 1260 3278
rect 1163 3275 1164 3276
rect 1158 3274 1164 3275
rect 1259 3275 1260 3276
rect 1264 3275 1265 3279
rect 1259 3274 1265 3275
rect 1278 3279 1284 3280
rect 1278 3275 1279 3279
rect 1283 3278 1284 3279
rect 1387 3279 1393 3280
rect 1387 3278 1388 3279
rect 1283 3276 1388 3278
rect 1283 3275 1284 3276
rect 1278 3274 1284 3275
rect 1387 3275 1388 3276
rect 1392 3275 1393 3279
rect 1894 3279 1895 3283
rect 1899 3279 1900 3283
rect 1894 3278 1900 3279
rect 1910 3283 1916 3284
rect 1910 3279 1911 3283
rect 1915 3282 1916 3283
rect 2054 3283 2060 3284
rect 1915 3280 2017 3282
rect 1915 3279 1916 3280
rect 1910 3278 1916 3279
rect 2054 3279 2055 3283
rect 2059 3282 2060 3283
rect 2302 3283 2308 3284
rect 2059 3280 2193 3282
rect 2059 3279 2060 3280
rect 2054 3278 2060 3279
rect 2302 3279 2303 3283
rect 2307 3282 2308 3283
rect 2414 3283 2420 3284
rect 2307 3280 2377 3282
rect 2307 3279 2308 3280
rect 2302 3278 2308 3279
rect 2414 3279 2415 3283
rect 2419 3282 2420 3283
rect 2750 3283 2756 3284
rect 2419 3280 2553 3282
rect 2419 3279 2420 3280
rect 2414 3278 2420 3279
rect 2750 3279 2751 3283
rect 2755 3279 2756 3283
rect 2911 3283 2917 3284
rect 2911 3282 2912 3283
rect 2905 3280 2912 3282
rect 2750 3278 2756 3279
rect 2911 3279 2912 3280
rect 2916 3279 2917 3283
rect 2920 3282 2922 3296
rect 2974 3292 2980 3293
rect 2974 3288 2975 3292
rect 2979 3288 2980 3292
rect 2974 3287 2980 3288
rect 3110 3292 3116 3293
rect 3110 3288 3111 3292
rect 3115 3288 3116 3292
rect 3110 3287 3116 3288
rect 3246 3292 3252 3293
rect 3246 3288 3247 3292
rect 3251 3288 3252 3292
rect 3246 3287 3252 3288
rect 3366 3292 3372 3293
rect 3366 3288 3367 3292
rect 3371 3288 3372 3292
rect 3366 3287 3372 3288
rect 3462 3289 3468 3290
rect 3462 3285 3463 3289
rect 3467 3285 3468 3289
rect 3462 3284 3468 3285
rect 3054 3283 3060 3284
rect 2920 3280 3017 3282
rect 2911 3278 2917 3279
rect 3054 3279 3055 3283
rect 3059 3282 3060 3283
rect 3191 3283 3197 3284
rect 3059 3280 3153 3282
rect 3059 3279 3060 3280
rect 3054 3278 3060 3279
rect 3191 3279 3192 3283
rect 3196 3282 3197 3283
rect 3326 3283 3332 3284
rect 3196 3280 3289 3282
rect 3196 3279 3197 3280
rect 3191 3278 3197 3279
rect 3326 3279 3327 3283
rect 3331 3282 3332 3283
rect 3331 3280 3409 3282
rect 3331 3279 3332 3280
rect 3326 3278 3332 3279
rect 1387 3274 1393 3275
rect 1830 3273 1836 3274
rect 1806 3272 1812 3273
rect 448 3268 578 3270
rect 382 3264 388 3265
rect 110 3261 116 3262
rect 110 3257 111 3261
rect 115 3257 116 3261
rect 382 3260 383 3264
rect 387 3260 388 3264
rect 382 3259 388 3260
rect 494 3264 500 3265
rect 494 3260 495 3264
rect 499 3260 500 3264
rect 494 3259 500 3260
rect 110 3256 116 3257
rect 454 3255 460 3256
rect 454 3251 455 3255
rect 459 3251 460 3255
rect 454 3250 460 3251
rect 566 3255 572 3256
rect 566 3251 567 3255
rect 571 3251 572 3255
rect 576 3254 578 3268
rect 1806 3268 1807 3272
rect 1811 3268 1812 3272
rect 1830 3269 1831 3273
rect 1835 3269 1836 3273
rect 1830 3268 1836 3269
rect 1974 3273 1980 3274
rect 1974 3269 1975 3273
rect 1979 3269 1980 3273
rect 1974 3268 1980 3269
rect 2150 3273 2156 3274
rect 2150 3269 2151 3273
rect 2155 3269 2156 3273
rect 2150 3268 2156 3269
rect 2334 3273 2340 3274
rect 2334 3269 2335 3273
rect 2339 3269 2340 3273
rect 2334 3268 2340 3269
rect 2510 3273 2516 3274
rect 2510 3269 2511 3273
rect 2515 3269 2516 3273
rect 2510 3268 2516 3269
rect 2678 3273 2684 3274
rect 2678 3269 2679 3273
rect 2683 3269 2684 3273
rect 2678 3268 2684 3269
rect 2830 3273 2836 3274
rect 2830 3269 2831 3273
rect 2835 3269 2836 3273
rect 2830 3268 2836 3269
rect 2974 3273 2980 3274
rect 2974 3269 2975 3273
rect 2979 3269 2980 3273
rect 2974 3268 2980 3269
rect 3110 3273 3116 3274
rect 3110 3269 3111 3273
rect 3115 3269 3116 3273
rect 3110 3268 3116 3269
rect 3246 3273 3252 3274
rect 3246 3269 3247 3273
rect 3251 3269 3252 3273
rect 3246 3268 3252 3269
rect 3366 3273 3372 3274
rect 3366 3269 3367 3273
rect 3371 3269 3372 3273
rect 3366 3268 3372 3269
rect 3462 3272 3468 3273
rect 3462 3268 3463 3272
rect 3467 3268 3468 3272
rect 1806 3267 1812 3268
rect 3462 3267 3468 3268
rect 606 3264 612 3265
rect 606 3260 607 3264
rect 611 3260 612 3264
rect 606 3259 612 3260
rect 726 3264 732 3265
rect 726 3260 727 3264
rect 731 3260 732 3264
rect 726 3259 732 3260
rect 846 3264 852 3265
rect 846 3260 847 3264
rect 851 3260 852 3264
rect 846 3259 852 3260
rect 966 3264 972 3265
rect 966 3260 967 3264
rect 971 3260 972 3264
rect 966 3259 972 3260
rect 1086 3264 1092 3265
rect 1086 3260 1087 3264
rect 1091 3260 1092 3264
rect 1086 3259 1092 3260
rect 1206 3264 1212 3265
rect 1206 3260 1207 3264
rect 1211 3260 1212 3264
rect 1206 3259 1212 3260
rect 1334 3264 1340 3265
rect 1334 3260 1335 3264
rect 1339 3260 1340 3264
rect 1334 3259 1340 3260
rect 1766 3261 1772 3262
rect 1766 3257 1767 3261
rect 1771 3257 1772 3261
rect 1766 3256 1772 3257
rect 694 3255 700 3256
rect 576 3252 649 3254
rect 566 3250 572 3251
rect 694 3251 695 3255
rect 699 3254 700 3255
rect 807 3255 813 3256
rect 699 3252 769 3254
rect 699 3251 700 3252
rect 694 3250 700 3251
rect 807 3251 808 3255
rect 812 3254 813 3255
rect 1038 3255 1044 3256
rect 812 3252 889 3254
rect 812 3251 813 3252
rect 807 3250 813 3251
rect 1038 3251 1039 3255
rect 1043 3251 1044 3255
rect 1038 3250 1044 3251
rect 1158 3255 1164 3256
rect 1158 3251 1159 3255
rect 1163 3251 1164 3255
rect 1158 3250 1164 3251
rect 1278 3255 1284 3256
rect 1278 3251 1279 3255
rect 1283 3251 1284 3255
rect 1278 3250 1284 3251
rect 1398 3255 1404 3256
rect 1398 3251 1399 3255
rect 1403 3251 1404 3255
rect 1398 3250 1404 3251
rect 382 3245 388 3246
rect 110 3244 116 3245
rect 110 3240 111 3244
rect 115 3240 116 3244
rect 382 3241 383 3245
rect 387 3241 388 3245
rect 382 3240 388 3241
rect 494 3245 500 3246
rect 494 3241 495 3245
rect 499 3241 500 3245
rect 494 3240 500 3241
rect 606 3245 612 3246
rect 606 3241 607 3245
rect 611 3241 612 3245
rect 606 3240 612 3241
rect 726 3245 732 3246
rect 726 3241 727 3245
rect 731 3241 732 3245
rect 726 3240 732 3241
rect 846 3245 852 3246
rect 846 3241 847 3245
rect 851 3241 852 3245
rect 846 3240 852 3241
rect 966 3245 972 3246
rect 966 3241 967 3245
rect 971 3241 972 3245
rect 966 3240 972 3241
rect 1086 3245 1092 3246
rect 1086 3241 1087 3245
rect 1091 3241 1092 3245
rect 1086 3240 1092 3241
rect 1206 3245 1212 3246
rect 1206 3241 1207 3245
rect 1211 3241 1212 3245
rect 1206 3240 1212 3241
rect 1334 3245 1340 3246
rect 1334 3241 1335 3245
rect 1339 3241 1340 3245
rect 1334 3240 1340 3241
rect 1766 3244 1772 3245
rect 1766 3240 1767 3244
rect 1771 3240 1772 3244
rect 110 3239 116 3240
rect 1766 3239 1772 3240
rect 1806 3220 1812 3221
rect 3462 3220 3468 3221
rect 1806 3216 1807 3220
rect 1811 3216 1812 3220
rect 1806 3215 1812 3216
rect 1830 3219 1836 3220
rect 1830 3215 1831 3219
rect 1835 3215 1836 3219
rect 1830 3214 1836 3215
rect 2030 3219 2036 3220
rect 2030 3215 2031 3219
rect 2035 3215 2036 3219
rect 2030 3214 2036 3215
rect 2246 3219 2252 3220
rect 2246 3215 2247 3219
rect 2251 3215 2252 3219
rect 2246 3214 2252 3215
rect 2454 3219 2460 3220
rect 2454 3215 2455 3219
rect 2459 3215 2460 3219
rect 2454 3214 2460 3215
rect 2654 3219 2660 3220
rect 2654 3215 2655 3219
rect 2659 3215 2660 3219
rect 2654 3214 2660 3215
rect 2838 3219 2844 3220
rect 2838 3215 2839 3219
rect 2843 3215 2844 3219
rect 2838 3214 2844 3215
rect 3022 3219 3028 3220
rect 3022 3215 3023 3219
rect 3027 3215 3028 3219
rect 3022 3214 3028 3215
rect 3206 3219 3212 3220
rect 3206 3215 3207 3219
rect 3211 3215 3212 3219
rect 3206 3214 3212 3215
rect 3366 3219 3372 3220
rect 3366 3215 3367 3219
rect 3371 3215 3372 3219
rect 3462 3216 3463 3220
rect 3467 3216 3468 3220
rect 3462 3215 3468 3216
rect 3366 3214 3372 3215
rect 2102 3211 2108 3212
rect 1975 3207 1981 3208
rect 1975 3206 1976 3207
rect 1905 3204 1976 3206
rect 1806 3203 1812 3204
rect 1806 3199 1807 3203
rect 1811 3199 1812 3203
rect 1975 3203 1976 3204
rect 1980 3203 1981 3207
rect 2102 3207 2103 3211
rect 2107 3207 2108 3211
rect 2447 3211 2453 3212
rect 2102 3206 2108 3207
rect 2318 3207 2324 3208
rect 1975 3202 1981 3203
rect 2318 3203 2319 3207
rect 2323 3203 2324 3207
rect 2447 3207 2448 3211
rect 2452 3210 2453 3211
rect 3438 3211 3444 3212
rect 2452 3208 2497 3210
rect 3199 3208 3249 3210
rect 2452 3207 2453 3208
rect 2447 3206 2453 3207
rect 2726 3207 2732 3208
rect 2318 3202 2324 3203
rect 2726 3203 2727 3207
rect 2731 3203 2732 3207
rect 2726 3202 2732 3203
rect 2910 3207 2916 3208
rect 2910 3203 2911 3207
rect 2915 3203 2916 3207
rect 2910 3202 2916 3203
rect 3094 3207 3100 3208
rect 3094 3203 3095 3207
rect 3099 3203 3100 3207
rect 3094 3202 3100 3203
rect 1806 3198 1812 3199
rect 1830 3200 1836 3201
rect 110 3196 116 3197
rect 1766 3196 1772 3197
rect 110 3192 111 3196
rect 115 3192 116 3196
rect 110 3191 116 3192
rect 302 3195 308 3196
rect 302 3191 303 3195
rect 307 3191 308 3195
rect 302 3190 308 3191
rect 422 3195 428 3196
rect 422 3191 423 3195
rect 427 3191 428 3195
rect 422 3190 428 3191
rect 542 3195 548 3196
rect 542 3191 543 3195
rect 547 3191 548 3195
rect 542 3190 548 3191
rect 670 3195 676 3196
rect 670 3191 671 3195
rect 675 3191 676 3195
rect 670 3190 676 3191
rect 798 3195 804 3196
rect 798 3191 799 3195
rect 803 3191 804 3195
rect 798 3190 804 3191
rect 926 3195 932 3196
rect 926 3191 927 3195
rect 931 3191 932 3195
rect 926 3190 932 3191
rect 1054 3195 1060 3196
rect 1054 3191 1055 3195
rect 1059 3191 1060 3195
rect 1054 3190 1060 3191
rect 1174 3195 1180 3196
rect 1174 3191 1175 3195
rect 1179 3191 1180 3195
rect 1174 3190 1180 3191
rect 1302 3195 1308 3196
rect 1302 3191 1303 3195
rect 1307 3191 1308 3195
rect 1302 3190 1308 3191
rect 1430 3195 1436 3196
rect 1430 3191 1431 3195
rect 1435 3191 1436 3195
rect 1766 3192 1767 3196
rect 1771 3192 1772 3196
rect 1830 3196 1831 3200
rect 1835 3196 1836 3200
rect 1830 3195 1836 3196
rect 2030 3200 2036 3201
rect 2030 3196 2031 3200
rect 2035 3196 2036 3200
rect 2030 3195 2036 3196
rect 2246 3200 2252 3201
rect 2246 3196 2247 3200
rect 2251 3196 2252 3200
rect 2246 3195 2252 3196
rect 2454 3200 2460 3201
rect 2454 3196 2455 3200
rect 2459 3196 2460 3200
rect 2454 3195 2460 3196
rect 2654 3200 2660 3201
rect 2654 3196 2655 3200
rect 2659 3196 2660 3200
rect 2654 3195 2660 3196
rect 2838 3200 2844 3201
rect 2838 3196 2839 3200
rect 2843 3196 2844 3200
rect 2838 3195 2844 3196
rect 3022 3200 3028 3201
rect 3022 3196 3023 3200
rect 3027 3196 3028 3200
rect 3022 3195 3028 3196
rect 3062 3195 3068 3196
rect 1766 3191 1772 3192
rect 3062 3191 3063 3195
rect 3067 3194 3068 3195
rect 3199 3194 3201 3208
rect 3438 3207 3439 3211
rect 3443 3207 3444 3211
rect 3438 3206 3444 3207
rect 3462 3203 3468 3204
rect 3206 3200 3212 3201
rect 3206 3196 3207 3200
rect 3211 3196 3212 3200
rect 3206 3195 3212 3196
rect 3366 3200 3372 3201
rect 3366 3196 3367 3200
rect 3371 3196 3372 3200
rect 3462 3199 3463 3203
rect 3467 3199 3468 3203
rect 3462 3198 3468 3199
rect 3366 3195 3372 3196
rect 3067 3192 3201 3194
rect 3067 3191 3068 3192
rect 1430 3190 1436 3191
rect 3062 3190 3068 3191
rect 758 3187 764 3188
rect 374 3183 380 3184
rect 110 3179 116 3180
rect 110 3175 111 3179
rect 115 3175 116 3179
rect 374 3179 375 3183
rect 379 3179 380 3183
rect 374 3178 380 3179
rect 494 3183 500 3184
rect 494 3179 495 3183
rect 499 3179 500 3183
rect 494 3178 500 3179
rect 614 3183 620 3184
rect 614 3179 615 3183
rect 619 3179 620 3183
rect 614 3178 620 3179
rect 742 3183 748 3184
rect 742 3179 743 3183
rect 747 3179 748 3183
rect 758 3183 759 3187
rect 763 3186 764 3187
rect 998 3187 1004 3188
rect 763 3184 841 3186
rect 763 3183 764 3184
rect 758 3182 764 3183
rect 998 3183 999 3187
rect 1003 3183 1004 3187
rect 998 3182 1004 3183
rect 1006 3187 1012 3188
rect 1006 3183 1007 3187
rect 1011 3186 1012 3187
rect 1134 3187 1140 3188
rect 1011 3184 1097 3186
rect 1011 3183 1012 3184
rect 1006 3182 1012 3183
rect 1134 3183 1135 3187
rect 1139 3186 1140 3187
rect 1382 3187 1388 3188
rect 1139 3184 1217 3186
rect 1139 3183 1140 3184
rect 1134 3182 1140 3183
rect 1374 3183 1380 3184
rect 742 3178 748 3179
rect 1374 3179 1375 3183
rect 1379 3179 1380 3183
rect 1382 3183 1383 3187
rect 1387 3186 1388 3187
rect 1387 3184 1473 3186
rect 1387 3183 1388 3184
rect 1382 3182 1388 3183
rect 1883 3183 1889 3184
rect 1374 3178 1380 3179
rect 1766 3179 1772 3180
rect 110 3174 116 3175
rect 302 3176 308 3177
rect 302 3172 303 3176
rect 307 3172 308 3176
rect 302 3171 308 3172
rect 422 3176 428 3177
rect 422 3172 423 3176
rect 427 3172 428 3176
rect 422 3171 428 3172
rect 542 3176 548 3177
rect 542 3172 543 3176
rect 547 3172 548 3176
rect 542 3171 548 3172
rect 670 3176 676 3177
rect 670 3172 671 3176
rect 675 3172 676 3176
rect 670 3171 676 3172
rect 798 3176 804 3177
rect 798 3172 799 3176
rect 803 3172 804 3176
rect 798 3171 804 3172
rect 926 3176 932 3177
rect 926 3172 927 3176
rect 931 3172 932 3176
rect 926 3171 932 3172
rect 1054 3176 1060 3177
rect 1054 3172 1055 3176
rect 1059 3172 1060 3176
rect 1054 3171 1060 3172
rect 1174 3176 1180 3177
rect 1174 3172 1175 3176
rect 1179 3172 1180 3176
rect 1174 3171 1180 3172
rect 1302 3176 1308 3177
rect 1302 3172 1303 3176
rect 1307 3172 1308 3176
rect 1302 3171 1308 3172
rect 1430 3176 1436 3177
rect 1430 3172 1431 3176
rect 1435 3172 1436 3176
rect 1766 3175 1767 3179
rect 1771 3175 1772 3179
rect 1883 3179 1884 3183
rect 1888 3182 1889 3183
rect 1902 3183 1908 3184
rect 1902 3182 1903 3183
rect 1888 3180 1903 3182
rect 1888 3179 1889 3180
rect 1883 3178 1889 3179
rect 1902 3179 1903 3180
rect 1907 3179 1908 3183
rect 1902 3178 1908 3179
rect 1975 3183 1981 3184
rect 1975 3179 1976 3183
rect 1980 3182 1981 3183
rect 2083 3183 2089 3184
rect 2083 3182 2084 3183
rect 1980 3180 2084 3182
rect 1980 3179 1981 3180
rect 1975 3178 1981 3179
rect 2083 3179 2084 3180
rect 2088 3179 2089 3183
rect 2083 3178 2089 3179
rect 2299 3183 2308 3184
rect 2299 3179 2300 3183
rect 2307 3179 2308 3183
rect 2299 3178 2308 3179
rect 2318 3183 2324 3184
rect 2318 3179 2319 3183
rect 2323 3182 2324 3183
rect 2507 3183 2513 3184
rect 2507 3182 2508 3183
rect 2323 3180 2508 3182
rect 2323 3179 2324 3180
rect 2318 3178 2324 3179
rect 2507 3179 2508 3180
rect 2512 3179 2513 3183
rect 2507 3178 2513 3179
rect 2646 3183 2652 3184
rect 2646 3179 2647 3183
rect 2651 3182 2652 3183
rect 2707 3183 2713 3184
rect 2707 3182 2708 3183
rect 2651 3180 2708 3182
rect 2651 3179 2652 3180
rect 2646 3178 2652 3179
rect 2707 3179 2708 3180
rect 2712 3179 2713 3183
rect 2707 3178 2713 3179
rect 2726 3183 2732 3184
rect 2726 3179 2727 3183
rect 2731 3182 2732 3183
rect 2891 3183 2897 3184
rect 2891 3182 2892 3183
rect 2731 3180 2892 3182
rect 2731 3179 2732 3180
rect 2726 3178 2732 3179
rect 2891 3179 2892 3180
rect 2896 3179 2897 3183
rect 2891 3178 2897 3179
rect 2910 3183 2916 3184
rect 2910 3179 2911 3183
rect 2915 3182 2916 3183
rect 3075 3183 3081 3184
rect 3075 3182 3076 3183
rect 2915 3180 3076 3182
rect 2915 3179 2916 3180
rect 2910 3178 2916 3179
rect 3075 3179 3076 3180
rect 3080 3179 3081 3183
rect 3075 3178 3081 3179
rect 3094 3183 3100 3184
rect 3094 3179 3095 3183
rect 3099 3182 3100 3183
rect 3259 3183 3265 3184
rect 3259 3182 3260 3183
rect 3099 3180 3260 3182
rect 3099 3179 3100 3180
rect 3094 3178 3100 3179
rect 3259 3179 3260 3180
rect 3264 3179 3265 3183
rect 3259 3178 3265 3179
rect 3419 3183 3425 3184
rect 3419 3179 3420 3183
rect 3424 3182 3425 3183
rect 3430 3183 3436 3184
rect 3430 3182 3431 3183
rect 3424 3180 3431 3182
rect 3424 3179 3425 3180
rect 3419 3178 3425 3179
rect 3430 3179 3431 3180
rect 3435 3179 3436 3183
rect 3430 3178 3436 3179
rect 1766 3174 1772 3175
rect 1430 3171 1436 3172
rect 1891 3171 1897 3172
rect 758 3167 764 3168
rect 758 3166 759 3167
rect 356 3164 759 3166
rect 356 3162 358 3164
rect 758 3163 759 3164
rect 763 3163 764 3167
rect 1382 3167 1388 3168
rect 1382 3166 1383 3167
rect 758 3162 764 3163
rect 1228 3164 1383 3166
rect 1228 3162 1230 3164
rect 1382 3163 1383 3164
rect 1387 3163 1388 3167
rect 1891 3167 1892 3171
rect 1896 3170 1897 3171
rect 1918 3171 1924 3172
rect 1918 3170 1919 3171
rect 1896 3168 1919 3170
rect 1896 3167 1897 3168
rect 1891 3166 1897 3167
rect 1918 3167 1919 3168
rect 1923 3167 1924 3171
rect 1918 3166 1924 3167
rect 2083 3171 2089 3172
rect 2083 3167 2084 3171
rect 2088 3170 2089 3171
rect 2110 3171 2116 3172
rect 2110 3170 2111 3171
rect 2088 3168 2111 3170
rect 2088 3167 2089 3168
rect 2083 3166 2089 3167
rect 2110 3167 2111 3168
rect 2115 3167 2116 3171
rect 2110 3166 2116 3167
rect 2254 3171 2260 3172
rect 2254 3167 2255 3171
rect 2259 3170 2260 3171
rect 2275 3171 2281 3172
rect 2275 3170 2276 3171
rect 2259 3168 2276 3170
rect 2259 3167 2260 3168
rect 2254 3166 2260 3167
rect 2275 3167 2276 3168
rect 2280 3167 2281 3171
rect 2275 3166 2281 3167
rect 2447 3171 2453 3172
rect 2447 3167 2448 3171
rect 2452 3170 2453 3171
rect 2459 3171 2465 3172
rect 2459 3170 2460 3171
rect 2452 3168 2460 3170
rect 2452 3167 2453 3168
rect 2447 3166 2453 3167
rect 2459 3167 2460 3168
rect 2464 3167 2465 3171
rect 2459 3166 2465 3167
rect 2627 3171 2633 3172
rect 2627 3167 2628 3171
rect 2632 3170 2633 3171
rect 2655 3171 2661 3172
rect 2655 3170 2656 3171
rect 2632 3168 2656 3170
rect 2632 3167 2633 3168
rect 2627 3166 2633 3167
rect 2655 3167 2656 3168
rect 2660 3167 2661 3171
rect 2655 3166 2661 3167
rect 2787 3171 2793 3172
rect 2787 3167 2788 3171
rect 2792 3170 2793 3171
rect 2814 3171 2820 3172
rect 2814 3170 2815 3171
rect 2792 3168 2815 3170
rect 2792 3167 2793 3168
rect 2787 3166 2793 3167
rect 2814 3167 2815 3168
rect 2819 3167 2820 3171
rect 2814 3166 2820 3167
rect 2931 3171 2937 3172
rect 2931 3167 2932 3171
rect 2936 3170 2937 3171
rect 2974 3171 2980 3172
rect 2974 3170 2975 3171
rect 2936 3168 2975 3170
rect 2936 3167 2937 3168
rect 2931 3166 2937 3167
rect 2974 3167 2975 3168
rect 2979 3167 2980 3171
rect 2974 3166 2980 3167
rect 3059 3171 3068 3172
rect 3059 3167 3060 3171
rect 3067 3167 3068 3171
rect 3059 3166 3068 3167
rect 3078 3171 3084 3172
rect 3078 3167 3079 3171
rect 3083 3170 3084 3171
rect 3187 3171 3193 3172
rect 3187 3170 3188 3171
rect 3083 3168 3188 3170
rect 3083 3167 3084 3168
rect 3078 3166 3084 3167
rect 3187 3167 3188 3168
rect 3192 3167 3193 3171
rect 3187 3166 3193 3167
rect 3315 3171 3321 3172
rect 3315 3167 3316 3171
rect 3320 3170 3321 3171
rect 3350 3171 3356 3172
rect 3350 3170 3351 3171
rect 3320 3168 3351 3170
rect 3320 3167 3321 3168
rect 3315 3166 3321 3167
rect 3350 3167 3351 3168
rect 3355 3167 3356 3171
rect 3350 3166 3356 3167
rect 3359 3171 3365 3172
rect 3359 3167 3360 3171
rect 3364 3170 3365 3171
rect 3419 3171 3425 3172
rect 3419 3170 3420 3171
rect 3364 3168 3420 3170
rect 3364 3167 3365 3168
rect 3359 3166 3365 3167
rect 3419 3167 3420 3168
rect 3424 3167 3425 3171
rect 3419 3166 3425 3167
rect 1382 3162 1388 3163
rect 355 3161 361 3162
rect 355 3157 356 3161
rect 360 3157 361 3161
rect 1227 3161 1233 3162
rect 355 3156 361 3157
rect 374 3159 380 3160
rect 374 3155 375 3159
rect 379 3158 380 3159
rect 475 3159 481 3160
rect 475 3158 476 3159
rect 379 3156 476 3158
rect 379 3155 380 3156
rect 374 3154 380 3155
rect 475 3155 476 3156
rect 480 3155 481 3159
rect 475 3154 481 3155
rect 566 3159 572 3160
rect 566 3155 567 3159
rect 571 3158 572 3159
rect 595 3159 601 3160
rect 595 3158 596 3159
rect 571 3156 596 3158
rect 571 3155 572 3156
rect 566 3154 572 3155
rect 595 3155 596 3156
rect 600 3155 601 3159
rect 595 3154 601 3155
rect 614 3159 620 3160
rect 614 3155 615 3159
rect 619 3158 620 3159
rect 723 3159 729 3160
rect 723 3158 724 3159
rect 619 3156 724 3158
rect 619 3155 620 3156
rect 614 3154 620 3155
rect 723 3155 724 3156
rect 728 3155 729 3159
rect 723 3154 729 3155
rect 742 3159 748 3160
rect 742 3155 743 3159
rect 747 3158 748 3159
rect 851 3159 857 3160
rect 851 3158 852 3159
rect 747 3156 852 3158
rect 747 3155 748 3156
rect 742 3154 748 3155
rect 851 3155 852 3156
rect 856 3155 857 3159
rect 851 3154 857 3155
rect 979 3159 985 3160
rect 979 3155 980 3159
rect 984 3158 985 3159
rect 1006 3159 1012 3160
rect 1006 3158 1007 3159
rect 984 3156 1007 3158
rect 984 3155 985 3156
rect 979 3154 985 3155
rect 1006 3155 1007 3156
rect 1011 3155 1012 3159
rect 1006 3154 1012 3155
rect 1107 3159 1113 3160
rect 1107 3155 1108 3159
rect 1112 3158 1113 3159
rect 1134 3159 1140 3160
rect 1134 3158 1135 3159
rect 1112 3156 1135 3158
rect 1112 3155 1113 3156
rect 1107 3154 1113 3155
rect 1134 3155 1135 3156
rect 1139 3155 1140 3159
rect 1227 3157 1228 3161
rect 1232 3157 1233 3161
rect 1227 3156 1233 3157
rect 1270 3159 1276 3160
rect 1134 3154 1140 3155
rect 1270 3155 1271 3159
rect 1275 3158 1276 3159
rect 1355 3159 1361 3160
rect 1355 3158 1356 3159
rect 1275 3156 1356 3158
rect 1275 3155 1276 3156
rect 1270 3154 1276 3155
rect 1355 3155 1356 3156
rect 1360 3155 1361 3159
rect 1355 3154 1361 3155
rect 1374 3159 1380 3160
rect 1374 3155 1375 3159
rect 1379 3158 1380 3159
rect 1483 3159 1489 3160
rect 1483 3158 1484 3159
rect 1379 3156 1484 3158
rect 1379 3155 1380 3156
rect 1374 3154 1380 3155
rect 1483 3155 1484 3156
rect 1488 3155 1489 3159
rect 1483 3154 1489 3155
rect 1838 3156 1844 3157
rect 1806 3153 1812 3154
rect 1806 3149 1807 3153
rect 1811 3149 1812 3153
rect 1838 3152 1839 3156
rect 1843 3152 1844 3156
rect 1838 3151 1844 3152
rect 2030 3156 2036 3157
rect 2030 3152 2031 3156
rect 2035 3152 2036 3156
rect 2030 3151 2036 3152
rect 2222 3156 2228 3157
rect 2222 3152 2223 3156
rect 2227 3152 2228 3156
rect 2222 3151 2228 3152
rect 2406 3156 2412 3157
rect 2406 3152 2407 3156
rect 2411 3152 2412 3156
rect 2406 3151 2412 3152
rect 2574 3156 2580 3157
rect 2574 3152 2575 3156
rect 2579 3152 2580 3156
rect 2574 3151 2580 3152
rect 2734 3156 2740 3157
rect 2734 3152 2735 3156
rect 2739 3152 2740 3156
rect 2734 3151 2740 3152
rect 2878 3156 2884 3157
rect 2878 3152 2879 3156
rect 2883 3152 2884 3156
rect 2878 3151 2884 3152
rect 3006 3156 3012 3157
rect 3006 3152 3007 3156
rect 3011 3152 3012 3156
rect 3006 3151 3012 3152
rect 3134 3156 3140 3157
rect 3134 3152 3135 3156
rect 3139 3152 3140 3156
rect 3134 3151 3140 3152
rect 3262 3156 3268 3157
rect 3262 3152 3263 3156
rect 3267 3152 3268 3156
rect 3262 3151 3268 3152
rect 3366 3156 3372 3157
rect 3366 3152 3367 3156
rect 3371 3152 3372 3156
rect 3366 3151 3372 3152
rect 3462 3153 3468 3154
rect 1806 3148 1812 3149
rect 3462 3149 3463 3153
rect 3467 3149 3468 3153
rect 3462 3148 3468 3149
rect 1902 3147 1908 3148
rect 1902 3143 1903 3147
rect 1907 3143 1908 3147
rect 1902 3142 1908 3143
rect 1918 3147 1924 3148
rect 1918 3143 1919 3147
rect 1923 3146 1924 3147
rect 2110 3147 2116 3148
rect 1923 3144 2073 3146
rect 1923 3143 1924 3144
rect 1918 3142 1924 3143
rect 2110 3143 2111 3147
rect 2115 3146 2116 3147
rect 2478 3147 2484 3148
rect 2115 3144 2265 3146
rect 2115 3143 2116 3144
rect 2110 3142 2116 3143
rect 2478 3143 2479 3147
rect 2483 3143 2484 3147
rect 2478 3142 2484 3143
rect 2646 3147 2652 3148
rect 2646 3143 2647 3147
rect 2651 3143 2652 3147
rect 2646 3142 2652 3143
rect 2655 3147 2661 3148
rect 2655 3143 2656 3147
rect 2660 3146 2661 3147
rect 2814 3147 2820 3148
rect 2660 3144 2777 3146
rect 2660 3143 2661 3144
rect 2655 3142 2661 3143
rect 2814 3143 2815 3147
rect 2819 3146 2820 3147
rect 3078 3147 3084 3148
rect 2819 3144 2921 3146
rect 2819 3143 2820 3144
rect 2814 3142 2820 3143
rect 3078 3143 3079 3147
rect 3083 3143 3084 3147
rect 3078 3142 3084 3143
rect 3206 3147 3212 3148
rect 3206 3143 3207 3147
rect 3211 3143 3212 3147
rect 3359 3147 3365 3148
rect 3359 3146 3360 3147
rect 3337 3144 3360 3146
rect 3206 3142 3212 3143
rect 3359 3143 3360 3144
rect 3364 3143 3365 3147
rect 3359 3142 3365 3143
rect 3430 3147 3436 3148
rect 3430 3143 3431 3147
rect 3435 3143 3436 3147
rect 3430 3142 3436 3143
rect 1838 3137 1844 3138
rect 1806 3136 1812 3137
rect 227 3135 233 3136
rect 227 3131 228 3135
rect 232 3134 233 3135
rect 246 3135 252 3136
rect 232 3132 242 3134
rect 232 3131 233 3132
rect 227 3130 233 3131
rect 240 3126 242 3132
rect 246 3131 247 3135
rect 251 3134 252 3135
rect 371 3135 377 3136
rect 371 3134 372 3135
rect 251 3132 372 3134
rect 251 3131 252 3132
rect 246 3130 252 3131
rect 371 3131 372 3132
rect 376 3131 377 3135
rect 371 3130 377 3131
rect 494 3135 500 3136
rect 494 3131 495 3135
rect 499 3134 500 3135
rect 523 3135 529 3136
rect 523 3134 524 3135
rect 499 3132 524 3134
rect 499 3131 500 3132
rect 494 3130 500 3131
rect 523 3131 524 3132
rect 528 3131 529 3135
rect 523 3130 529 3131
rect 591 3135 597 3136
rect 591 3131 592 3135
rect 596 3134 597 3135
rect 675 3135 681 3136
rect 675 3134 676 3135
rect 596 3132 676 3134
rect 596 3131 597 3132
rect 591 3130 597 3131
rect 675 3131 676 3132
rect 680 3131 681 3135
rect 675 3130 681 3131
rect 694 3135 700 3136
rect 694 3131 695 3135
rect 699 3134 700 3135
rect 827 3135 833 3136
rect 827 3134 828 3135
rect 699 3132 828 3134
rect 699 3131 700 3132
rect 694 3130 700 3131
rect 827 3131 828 3132
rect 832 3131 833 3135
rect 827 3130 833 3131
rect 971 3135 977 3136
rect 971 3131 972 3135
rect 976 3134 977 3135
rect 990 3135 996 3136
rect 976 3132 986 3134
rect 976 3131 977 3132
rect 971 3130 977 3131
rect 984 3126 986 3132
rect 990 3131 991 3135
rect 995 3134 996 3135
rect 1115 3135 1121 3136
rect 1115 3134 1116 3135
rect 995 3132 1116 3134
rect 995 3131 996 3132
rect 990 3130 996 3131
rect 1115 3131 1116 3132
rect 1120 3131 1121 3135
rect 1115 3130 1121 3131
rect 1134 3135 1140 3136
rect 1134 3131 1135 3135
rect 1139 3134 1140 3135
rect 1251 3135 1257 3136
rect 1251 3134 1252 3135
rect 1139 3132 1252 3134
rect 1139 3131 1140 3132
rect 1134 3130 1140 3131
rect 1251 3131 1252 3132
rect 1256 3131 1257 3135
rect 1251 3130 1257 3131
rect 1395 3135 1401 3136
rect 1395 3131 1396 3135
rect 1400 3134 1401 3135
rect 1422 3135 1428 3136
rect 1422 3134 1423 3135
rect 1400 3132 1423 3134
rect 1400 3131 1401 3132
rect 1395 3130 1401 3131
rect 1422 3131 1423 3132
rect 1427 3131 1428 3135
rect 1422 3130 1428 3131
rect 1539 3135 1545 3136
rect 1539 3131 1540 3135
rect 1544 3134 1545 3135
rect 1582 3135 1588 3136
rect 1582 3134 1583 3135
rect 1544 3132 1583 3134
rect 1544 3131 1545 3132
rect 1539 3130 1545 3131
rect 1582 3131 1583 3132
rect 1587 3131 1588 3135
rect 1806 3132 1807 3136
rect 1811 3132 1812 3136
rect 1838 3133 1839 3137
rect 1843 3133 1844 3137
rect 1838 3132 1844 3133
rect 2030 3137 2036 3138
rect 2030 3133 2031 3137
rect 2035 3133 2036 3137
rect 2030 3132 2036 3133
rect 2222 3137 2228 3138
rect 2222 3133 2223 3137
rect 2227 3133 2228 3137
rect 2222 3132 2228 3133
rect 2406 3137 2412 3138
rect 2406 3133 2407 3137
rect 2411 3133 2412 3137
rect 2406 3132 2412 3133
rect 2574 3137 2580 3138
rect 2574 3133 2575 3137
rect 2579 3133 2580 3137
rect 2574 3132 2580 3133
rect 2734 3137 2740 3138
rect 2734 3133 2735 3137
rect 2739 3133 2740 3137
rect 2734 3132 2740 3133
rect 2878 3137 2884 3138
rect 2878 3133 2879 3137
rect 2883 3133 2884 3137
rect 2878 3132 2884 3133
rect 3006 3137 3012 3138
rect 3006 3133 3007 3137
rect 3011 3133 3012 3137
rect 3006 3132 3012 3133
rect 3134 3137 3140 3138
rect 3134 3133 3135 3137
rect 3139 3133 3140 3137
rect 3134 3132 3140 3133
rect 3262 3137 3268 3138
rect 3262 3133 3263 3137
rect 3267 3133 3268 3137
rect 3262 3132 3268 3133
rect 3366 3137 3372 3138
rect 3366 3133 3367 3137
rect 3371 3133 3372 3137
rect 3366 3132 3372 3133
rect 3462 3136 3468 3137
rect 3462 3132 3463 3136
rect 3467 3132 3468 3136
rect 1806 3131 1812 3132
rect 3462 3131 3468 3132
rect 1582 3130 1588 3131
rect 240 3124 750 3126
rect 984 3124 1282 3126
rect 174 3120 180 3121
rect 110 3117 116 3118
rect 110 3113 111 3117
rect 115 3113 116 3117
rect 174 3116 175 3120
rect 179 3116 180 3120
rect 174 3115 180 3116
rect 318 3120 324 3121
rect 318 3116 319 3120
rect 323 3116 324 3120
rect 318 3115 324 3116
rect 470 3120 476 3121
rect 470 3116 471 3120
rect 475 3116 476 3120
rect 470 3115 476 3116
rect 622 3120 628 3121
rect 622 3116 623 3120
rect 627 3116 628 3120
rect 622 3115 628 3116
rect 110 3112 116 3113
rect 246 3111 252 3112
rect 246 3107 247 3111
rect 251 3107 252 3111
rect 246 3106 252 3107
rect 390 3111 396 3112
rect 390 3107 391 3111
rect 395 3107 396 3111
rect 591 3111 597 3112
rect 591 3110 592 3111
rect 545 3108 592 3110
rect 390 3106 396 3107
rect 591 3107 592 3108
rect 596 3107 597 3111
rect 591 3106 597 3107
rect 694 3111 700 3112
rect 694 3107 695 3111
rect 699 3107 700 3111
rect 748 3110 750 3124
rect 774 3120 780 3121
rect 774 3116 775 3120
rect 779 3116 780 3120
rect 774 3115 780 3116
rect 918 3120 924 3121
rect 918 3116 919 3120
rect 923 3116 924 3120
rect 918 3115 924 3116
rect 1062 3120 1068 3121
rect 1062 3116 1063 3120
rect 1067 3116 1068 3120
rect 1062 3115 1068 3116
rect 1198 3120 1204 3121
rect 1198 3116 1199 3120
rect 1203 3116 1204 3120
rect 1198 3115 1204 3116
rect 990 3111 996 3112
rect 748 3108 817 3110
rect 694 3106 700 3107
rect 990 3107 991 3111
rect 995 3107 996 3111
rect 990 3106 996 3107
rect 1134 3111 1140 3112
rect 1134 3107 1135 3111
rect 1139 3107 1140 3111
rect 1134 3106 1140 3107
rect 1270 3111 1276 3112
rect 1270 3107 1271 3111
rect 1275 3107 1276 3111
rect 1280 3110 1282 3124
rect 1342 3120 1348 3121
rect 1342 3116 1343 3120
rect 1347 3116 1348 3120
rect 1342 3115 1348 3116
rect 1486 3120 1492 3121
rect 1486 3116 1487 3120
rect 1491 3116 1492 3120
rect 1486 3115 1492 3116
rect 1766 3117 1772 3118
rect 1766 3113 1767 3117
rect 1771 3113 1772 3117
rect 1766 3112 1772 3113
rect 1422 3111 1428 3112
rect 1280 3108 1385 3110
rect 1270 3106 1276 3107
rect 1422 3107 1423 3111
rect 1427 3110 1428 3111
rect 1427 3108 1529 3110
rect 1427 3107 1428 3108
rect 1422 3106 1428 3107
rect 174 3101 180 3102
rect 110 3100 116 3101
rect 110 3096 111 3100
rect 115 3096 116 3100
rect 174 3097 175 3101
rect 179 3097 180 3101
rect 174 3096 180 3097
rect 318 3101 324 3102
rect 318 3097 319 3101
rect 323 3097 324 3101
rect 318 3096 324 3097
rect 470 3101 476 3102
rect 470 3097 471 3101
rect 475 3097 476 3101
rect 470 3096 476 3097
rect 622 3101 628 3102
rect 622 3097 623 3101
rect 627 3097 628 3101
rect 622 3096 628 3097
rect 774 3101 780 3102
rect 774 3097 775 3101
rect 779 3097 780 3101
rect 774 3096 780 3097
rect 918 3101 924 3102
rect 918 3097 919 3101
rect 923 3097 924 3101
rect 918 3096 924 3097
rect 1062 3101 1068 3102
rect 1062 3097 1063 3101
rect 1067 3097 1068 3101
rect 1062 3096 1068 3097
rect 1198 3101 1204 3102
rect 1198 3097 1199 3101
rect 1203 3097 1204 3101
rect 1198 3096 1204 3097
rect 1342 3101 1348 3102
rect 1342 3097 1343 3101
rect 1347 3097 1348 3101
rect 1342 3096 1348 3097
rect 1486 3101 1492 3102
rect 1486 3097 1487 3101
rect 1491 3097 1492 3101
rect 1486 3096 1492 3097
rect 1766 3100 1772 3101
rect 1766 3096 1767 3100
rect 1771 3096 1772 3100
rect 110 3095 116 3096
rect 1766 3095 1772 3096
rect 1806 3088 1812 3089
rect 3462 3088 3468 3089
rect 1806 3084 1807 3088
rect 1811 3084 1812 3088
rect 1806 3083 1812 3084
rect 1934 3087 1940 3088
rect 1934 3083 1935 3087
rect 1939 3083 1940 3087
rect 1934 3082 1940 3083
rect 2054 3087 2060 3088
rect 2054 3083 2055 3087
rect 2059 3083 2060 3087
rect 2054 3082 2060 3083
rect 2174 3087 2180 3088
rect 2174 3083 2175 3087
rect 2179 3083 2180 3087
rect 2174 3082 2180 3083
rect 2302 3087 2308 3088
rect 2302 3083 2303 3087
rect 2307 3083 2308 3087
rect 2302 3082 2308 3083
rect 2430 3087 2436 3088
rect 2430 3083 2431 3087
rect 2435 3083 2436 3087
rect 2430 3082 2436 3083
rect 2566 3087 2572 3088
rect 2566 3083 2567 3087
rect 2571 3083 2572 3087
rect 2566 3082 2572 3083
rect 2718 3087 2724 3088
rect 2718 3083 2719 3087
rect 2723 3083 2724 3087
rect 2718 3082 2724 3083
rect 2870 3087 2876 3088
rect 2870 3083 2871 3087
rect 2875 3083 2876 3087
rect 2870 3082 2876 3083
rect 3030 3087 3036 3088
rect 3030 3083 3031 3087
rect 3035 3083 3036 3087
rect 3030 3082 3036 3083
rect 3198 3087 3204 3088
rect 3198 3083 3199 3087
rect 3203 3083 3204 3087
rect 3198 3082 3204 3083
rect 3366 3087 3372 3088
rect 3366 3083 3367 3087
rect 3371 3083 3372 3087
rect 3462 3084 3463 3088
rect 3467 3084 3468 3088
rect 3462 3083 3468 3084
rect 3366 3082 3372 3083
rect 2254 3079 2260 3080
rect 2254 3078 2255 3079
rect 2249 3076 2255 3078
rect 2006 3075 2012 3076
rect 1806 3071 1812 3072
rect 1806 3067 1807 3071
rect 1811 3067 1812 3071
rect 2006 3071 2007 3075
rect 2011 3071 2012 3075
rect 2006 3070 2012 3071
rect 2126 3075 2132 3076
rect 2126 3071 2127 3075
rect 2131 3071 2132 3075
rect 2254 3075 2255 3076
rect 2259 3075 2260 3079
rect 2414 3079 2420 3080
rect 2254 3074 2260 3075
rect 2374 3075 2380 3076
rect 2126 3070 2132 3071
rect 2374 3071 2375 3075
rect 2379 3071 2380 3075
rect 2414 3075 2415 3079
rect 2419 3078 2420 3079
rect 2974 3079 2980 3080
rect 2419 3076 2473 3078
rect 2419 3075 2420 3076
rect 2414 3074 2420 3075
rect 2638 3075 2644 3076
rect 2374 3070 2380 3071
rect 2638 3071 2639 3075
rect 2643 3071 2644 3075
rect 2638 3070 2644 3071
rect 2790 3075 2796 3076
rect 2790 3071 2791 3075
rect 2795 3071 2796 3075
rect 2790 3070 2796 3071
rect 2942 3075 2948 3076
rect 2942 3071 2943 3075
rect 2947 3071 2948 3075
rect 2974 3075 2975 3079
rect 2979 3078 2980 3079
rect 3350 3079 3356 3080
rect 2979 3076 3073 3078
rect 2979 3075 2980 3076
rect 2974 3074 2980 3075
rect 3270 3075 3276 3076
rect 2942 3070 2948 3071
rect 3270 3071 3271 3075
rect 3275 3071 3276 3075
rect 3350 3075 3351 3079
rect 3355 3078 3356 3079
rect 3355 3076 3409 3078
rect 3355 3075 3356 3076
rect 3350 3074 3356 3075
rect 3270 3070 3276 3071
rect 3462 3071 3468 3072
rect 1806 3066 1812 3067
rect 1934 3068 1940 3069
rect 1934 3064 1935 3068
rect 1939 3064 1940 3068
rect 1934 3063 1940 3064
rect 2054 3068 2060 3069
rect 2054 3064 2055 3068
rect 2059 3064 2060 3068
rect 2054 3063 2060 3064
rect 2174 3068 2180 3069
rect 2174 3064 2175 3068
rect 2179 3064 2180 3068
rect 2174 3063 2180 3064
rect 2302 3068 2308 3069
rect 2302 3064 2303 3068
rect 2307 3064 2308 3068
rect 2302 3063 2308 3064
rect 2430 3068 2436 3069
rect 2430 3064 2431 3068
rect 2435 3064 2436 3068
rect 2430 3063 2436 3064
rect 2566 3068 2572 3069
rect 2566 3064 2567 3068
rect 2571 3064 2572 3068
rect 2566 3063 2572 3064
rect 2718 3068 2724 3069
rect 2718 3064 2719 3068
rect 2723 3064 2724 3068
rect 2718 3063 2724 3064
rect 2870 3068 2876 3069
rect 2870 3064 2871 3068
rect 2875 3064 2876 3068
rect 2870 3063 2876 3064
rect 3030 3068 3036 3069
rect 3030 3064 3031 3068
rect 3035 3064 3036 3068
rect 3030 3063 3036 3064
rect 3198 3068 3204 3069
rect 3198 3064 3199 3068
rect 3203 3064 3204 3068
rect 3198 3063 3204 3064
rect 3366 3068 3372 3069
rect 3366 3064 3367 3068
rect 3371 3064 3372 3068
rect 3462 3067 3463 3071
rect 3467 3067 3468 3071
rect 3462 3066 3468 3067
rect 3366 3063 3372 3064
rect 1987 3051 1996 3052
rect 110 3048 116 3049
rect 1766 3048 1772 3049
rect 110 3044 111 3048
rect 115 3044 116 3048
rect 110 3043 116 3044
rect 134 3047 140 3048
rect 134 3043 135 3047
rect 139 3043 140 3047
rect 134 3042 140 3043
rect 262 3047 268 3048
rect 262 3043 263 3047
rect 267 3043 268 3047
rect 262 3042 268 3043
rect 430 3047 436 3048
rect 430 3043 431 3047
rect 435 3043 436 3047
rect 430 3042 436 3043
rect 606 3047 612 3048
rect 606 3043 607 3047
rect 611 3043 612 3047
rect 606 3042 612 3043
rect 790 3047 796 3048
rect 790 3043 791 3047
rect 795 3043 796 3047
rect 790 3042 796 3043
rect 966 3047 972 3048
rect 966 3043 967 3047
rect 971 3043 972 3047
rect 966 3042 972 3043
rect 1142 3047 1148 3048
rect 1142 3043 1143 3047
rect 1147 3043 1148 3047
rect 1142 3042 1148 3043
rect 1326 3047 1332 3048
rect 1326 3043 1327 3047
rect 1331 3043 1332 3047
rect 1326 3042 1332 3043
rect 1510 3047 1516 3048
rect 1510 3043 1511 3047
rect 1515 3043 1516 3047
rect 1766 3044 1767 3048
rect 1771 3044 1772 3048
rect 1987 3047 1988 3051
rect 1995 3047 1996 3051
rect 1987 3046 1996 3047
rect 2006 3051 2012 3052
rect 2006 3047 2007 3051
rect 2011 3050 2012 3051
rect 2107 3051 2113 3052
rect 2107 3050 2108 3051
rect 2011 3048 2108 3050
rect 2011 3047 2012 3048
rect 2006 3046 2012 3047
rect 2107 3047 2108 3048
rect 2112 3047 2113 3051
rect 2107 3046 2113 3047
rect 2126 3051 2132 3052
rect 2126 3047 2127 3051
rect 2131 3050 2132 3051
rect 2227 3051 2233 3052
rect 2227 3050 2228 3051
rect 2131 3048 2228 3050
rect 2131 3047 2132 3048
rect 2126 3046 2132 3047
rect 2227 3047 2228 3048
rect 2232 3047 2233 3051
rect 2227 3046 2233 3047
rect 2355 3051 2361 3052
rect 2355 3047 2356 3051
rect 2360 3050 2361 3051
rect 2414 3051 2420 3052
rect 2414 3050 2415 3051
rect 2360 3048 2415 3050
rect 2360 3047 2361 3048
rect 2355 3046 2361 3047
rect 2414 3047 2415 3048
rect 2419 3047 2420 3051
rect 2414 3046 2420 3047
rect 2478 3051 2489 3052
rect 2478 3047 2479 3051
rect 2483 3047 2484 3051
rect 2488 3047 2489 3051
rect 2478 3046 2489 3047
rect 2619 3051 2625 3052
rect 2619 3047 2620 3051
rect 2624 3050 2625 3051
rect 2638 3051 2644 3052
rect 2624 3048 2634 3050
rect 2624 3047 2625 3048
rect 2619 3046 2625 3047
rect 1766 3043 1772 3044
rect 1510 3042 1516 3043
rect 2632 3042 2634 3048
rect 2638 3047 2639 3051
rect 2643 3050 2644 3051
rect 2771 3051 2777 3052
rect 2771 3050 2772 3051
rect 2643 3048 2772 3050
rect 2643 3047 2644 3048
rect 2638 3046 2644 3047
rect 2771 3047 2772 3048
rect 2776 3047 2777 3051
rect 2771 3046 2777 3047
rect 2790 3051 2796 3052
rect 2790 3047 2791 3051
rect 2795 3050 2796 3051
rect 2923 3051 2929 3052
rect 2923 3050 2924 3051
rect 2795 3048 2924 3050
rect 2795 3047 2796 3048
rect 2790 3046 2796 3047
rect 2923 3047 2924 3048
rect 2928 3047 2929 3051
rect 2923 3046 2929 3047
rect 2942 3051 2948 3052
rect 2942 3047 2943 3051
rect 2947 3050 2948 3051
rect 3083 3051 3089 3052
rect 3083 3050 3084 3051
rect 2947 3048 3084 3050
rect 2947 3047 2948 3048
rect 2942 3046 2948 3047
rect 3083 3047 3084 3048
rect 3088 3047 3089 3051
rect 3083 3046 3089 3047
rect 3206 3051 3212 3052
rect 3206 3047 3207 3051
rect 3211 3050 3212 3051
rect 3251 3051 3257 3052
rect 3251 3050 3252 3051
rect 3211 3048 3252 3050
rect 3211 3047 3212 3048
rect 3206 3046 3212 3047
rect 3251 3047 3252 3048
rect 3256 3047 3257 3051
rect 3251 3046 3257 3047
rect 3270 3051 3276 3052
rect 3270 3047 3271 3051
rect 3275 3050 3276 3051
rect 3419 3051 3425 3052
rect 3419 3050 3420 3051
rect 3275 3048 3420 3050
rect 3275 3047 3276 3048
rect 3270 3046 3276 3047
rect 3419 3047 3420 3048
rect 3424 3047 3425 3051
rect 3419 3046 3425 3047
rect 2822 3043 2828 3044
rect 2822 3042 2823 3043
rect 2632 3040 2823 3042
rect 754 3039 760 3040
rect 206 3035 212 3036
rect 110 3031 116 3032
rect 110 3027 111 3031
rect 115 3027 116 3031
rect 206 3031 207 3035
rect 211 3031 212 3035
rect 206 3030 212 3031
rect 334 3035 340 3036
rect 334 3031 335 3035
rect 339 3031 340 3035
rect 334 3030 340 3031
rect 502 3035 508 3036
rect 502 3031 503 3035
rect 507 3031 508 3035
rect 502 3030 508 3031
rect 678 3035 684 3036
rect 678 3031 679 3035
rect 683 3031 684 3035
rect 754 3035 755 3039
rect 759 3038 760 3039
rect 1582 3039 1588 3040
rect 759 3036 833 3038
rect 759 3035 760 3036
rect 754 3034 760 3035
rect 1038 3035 1044 3036
rect 678 3030 684 3031
rect 1038 3031 1039 3035
rect 1043 3031 1044 3035
rect 1038 3030 1044 3031
rect 1214 3035 1220 3036
rect 1214 3031 1215 3035
rect 1219 3031 1220 3035
rect 1214 3030 1220 3031
rect 1398 3035 1404 3036
rect 1398 3031 1399 3035
rect 1403 3031 1404 3035
rect 1582 3035 1583 3039
rect 1587 3035 1588 3039
rect 2822 3039 2823 3040
rect 2827 3039 2828 3043
rect 2822 3038 2828 3039
rect 1582 3034 1588 3035
rect 1398 3030 1404 3031
rect 1766 3031 1772 3032
rect 110 3026 116 3027
rect 134 3028 140 3029
rect 134 3024 135 3028
rect 139 3024 140 3028
rect 134 3023 140 3024
rect 262 3028 268 3029
rect 262 3024 263 3028
rect 267 3024 268 3028
rect 262 3023 268 3024
rect 430 3028 436 3029
rect 430 3024 431 3028
rect 435 3024 436 3028
rect 430 3023 436 3024
rect 606 3028 612 3029
rect 606 3024 607 3028
rect 611 3024 612 3028
rect 606 3023 612 3024
rect 790 3028 796 3029
rect 790 3024 791 3028
rect 795 3024 796 3028
rect 790 3023 796 3024
rect 966 3028 972 3029
rect 966 3024 967 3028
rect 971 3024 972 3028
rect 966 3023 972 3024
rect 1142 3028 1148 3029
rect 1142 3024 1143 3028
rect 1147 3024 1148 3028
rect 1142 3023 1148 3024
rect 1326 3028 1332 3029
rect 1326 3024 1327 3028
rect 1331 3024 1332 3028
rect 1326 3023 1332 3024
rect 1510 3028 1516 3029
rect 1510 3024 1511 3028
rect 1515 3024 1516 3028
rect 1766 3027 1767 3031
rect 1771 3027 1772 3031
rect 1766 3026 1772 3027
rect 2075 3031 2081 3032
rect 2075 3027 2076 3031
rect 2080 3030 2081 3031
rect 2134 3031 2140 3032
rect 2080 3028 2130 3030
rect 2080 3027 2081 3028
rect 2075 3026 2081 3027
rect 1510 3023 1516 3024
rect 2128 3022 2130 3028
rect 2134 3027 2135 3031
rect 2139 3030 2140 3031
rect 2179 3031 2185 3032
rect 2179 3030 2180 3031
rect 2139 3028 2180 3030
rect 2139 3027 2140 3028
rect 2134 3026 2140 3027
rect 2179 3027 2180 3028
rect 2184 3027 2185 3031
rect 2179 3026 2185 3027
rect 2198 3031 2204 3032
rect 2198 3027 2199 3031
rect 2203 3030 2204 3031
rect 2283 3031 2289 3032
rect 2283 3030 2284 3031
rect 2203 3028 2284 3030
rect 2203 3027 2204 3028
rect 2198 3026 2204 3027
rect 2283 3027 2284 3028
rect 2288 3027 2289 3031
rect 2283 3026 2289 3027
rect 2374 3031 2380 3032
rect 2374 3027 2375 3031
rect 2379 3030 2380 3031
rect 2387 3031 2393 3032
rect 2387 3030 2388 3031
rect 2379 3028 2388 3030
rect 2379 3027 2380 3028
rect 2374 3026 2380 3027
rect 2387 3027 2388 3028
rect 2392 3027 2393 3031
rect 2387 3026 2393 3027
rect 2491 3031 2497 3032
rect 2491 3027 2492 3031
rect 2496 3030 2497 3031
rect 2510 3031 2516 3032
rect 2496 3028 2506 3030
rect 2496 3027 2497 3028
rect 2491 3026 2497 3027
rect 2504 3022 2506 3028
rect 2510 3027 2511 3031
rect 2515 3030 2516 3031
rect 2595 3031 2601 3032
rect 2595 3030 2596 3031
rect 2515 3028 2596 3030
rect 2515 3027 2516 3028
rect 2510 3026 2516 3027
rect 2595 3027 2596 3028
rect 2600 3027 2601 3031
rect 2595 3026 2601 3027
rect 2614 3031 2620 3032
rect 2614 3027 2615 3031
rect 2619 3030 2620 3031
rect 2699 3031 2705 3032
rect 2699 3030 2700 3031
rect 2619 3028 2700 3030
rect 2619 3027 2620 3028
rect 2614 3026 2620 3027
rect 2699 3027 2700 3028
rect 2704 3027 2705 3031
rect 2699 3026 2705 3027
rect 2750 3031 2756 3032
rect 2750 3027 2751 3031
rect 2755 3030 2756 3031
rect 2811 3031 2817 3032
rect 2811 3030 2812 3031
rect 2755 3028 2812 3030
rect 2755 3027 2756 3028
rect 2750 3026 2756 3027
rect 2811 3027 2812 3028
rect 2816 3027 2817 3031
rect 2811 3026 2817 3027
rect 2662 3023 2668 3024
rect 2662 3022 2663 3023
rect 2128 3020 2210 3022
rect 2504 3020 2663 3022
rect 754 3019 760 3020
rect 754 3018 755 3019
rect 188 3016 755 3018
rect 188 3014 190 3016
rect 754 3015 755 3016
rect 759 3015 760 3019
rect 754 3014 760 3015
rect 2022 3016 2028 3017
rect 187 3013 193 3014
rect 187 3009 188 3013
rect 192 3009 193 3013
rect 1806 3013 1812 3014
rect 187 3008 193 3009
rect 206 3011 212 3012
rect 206 3007 207 3011
rect 211 3010 212 3011
rect 315 3011 321 3012
rect 315 3010 316 3011
rect 211 3008 316 3010
rect 211 3007 212 3008
rect 206 3006 212 3007
rect 315 3007 316 3008
rect 320 3007 321 3011
rect 315 3006 321 3007
rect 390 3011 396 3012
rect 390 3007 391 3011
rect 395 3010 396 3011
rect 483 3011 489 3012
rect 483 3010 484 3011
rect 395 3008 484 3010
rect 395 3007 396 3008
rect 390 3006 396 3007
rect 483 3007 484 3008
rect 488 3007 489 3011
rect 483 3006 489 3007
rect 502 3011 508 3012
rect 502 3007 503 3011
rect 507 3010 508 3011
rect 659 3011 665 3012
rect 659 3010 660 3011
rect 507 3008 660 3010
rect 507 3007 508 3008
rect 502 3006 508 3007
rect 659 3007 660 3008
rect 664 3007 665 3011
rect 659 3006 665 3007
rect 678 3011 684 3012
rect 678 3007 679 3011
rect 683 3010 684 3011
rect 843 3011 849 3012
rect 843 3010 844 3011
rect 683 3008 844 3010
rect 683 3007 684 3008
rect 678 3006 684 3007
rect 843 3007 844 3008
rect 848 3007 849 3011
rect 843 3006 849 3007
rect 998 3011 1004 3012
rect 998 3007 999 3011
rect 1003 3010 1004 3011
rect 1019 3011 1025 3012
rect 1019 3010 1020 3011
rect 1003 3008 1020 3010
rect 1003 3007 1004 3008
rect 998 3006 1004 3007
rect 1019 3007 1020 3008
rect 1024 3007 1025 3011
rect 1019 3006 1025 3007
rect 1038 3011 1044 3012
rect 1038 3007 1039 3011
rect 1043 3010 1044 3011
rect 1195 3011 1201 3012
rect 1195 3010 1196 3011
rect 1043 3008 1196 3010
rect 1043 3007 1044 3008
rect 1038 3006 1044 3007
rect 1195 3007 1196 3008
rect 1200 3007 1201 3011
rect 1195 3006 1201 3007
rect 1214 3011 1220 3012
rect 1214 3007 1215 3011
rect 1219 3010 1220 3011
rect 1379 3011 1385 3012
rect 1379 3010 1380 3011
rect 1219 3008 1380 3010
rect 1219 3007 1220 3008
rect 1214 3006 1220 3007
rect 1379 3007 1380 3008
rect 1384 3007 1385 3011
rect 1379 3006 1385 3007
rect 1398 3011 1404 3012
rect 1398 3007 1399 3011
rect 1403 3010 1404 3011
rect 1563 3011 1569 3012
rect 1563 3010 1564 3011
rect 1403 3008 1564 3010
rect 1403 3007 1404 3008
rect 1398 3006 1404 3007
rect 1563 3007 1564 3008
rect 1568 3007 1569 3011
rect 1806 3009 1807 3013
rect 1811 3009 1812 3013
rect 2022 3012 2023 3016
rect 2027 3012 2028 3016
rect 2022 3011 2028 3012
rect 2126 3016 2132 3017
rect 2126 3012 2127 3016
rect 2131 3012 2132 3016
rect 2126 3011 2132 3012
rect 1806 3008 1812 3009
rect 1563 3006 1569 3007
rect 1990 3007 1996 3008
rect 1990 3003 1991 3007
rect 1995 3006 1996 3007
rect 2198 3007 2204 3008
rect 1995 3004 2065 3006
rect 1995 3003 1996 3004
rect 1990 3002 1996 3003
rect 2198 3003 2199 3007
rect 2203 3003 2204 3007
rect 2208 3006 2210 3020
rect 2662 3019 2663 3020
rect 2667 3019 2668 3023
rect 2662 3018 2668 3019
rect 2230 3016 2236 3017
rect 2230 3012 2231 3016
rect 2235 3012 2236 3016
rect 2230 3011 2236 3012
rect 2334 3016 2340 3017
rect 2334 3012 2335 3016
rect 2339 3012 2340 3016
rect 2334 3011 2340 3012
rect 2438 3016 2444 3017
rect 2438 3012 2439 3016
rect 2443 3012 2444 3016
rect 2438 3011 2444 3012
rect 2542 3016 2548 3017
rect 2542 3012 2543 3016
rect 2547 3012 2548 3016
rect 2542 3011 2548 3012
rect 2646 3016 2652 3017
rect 2646 3012 2647 3016
rect 2651 3012 2652 3016
rect 2646 3011 2652 3012
rect 2758 3016 2764 3017
rect 2758 3012 2759 3016
rect 2763 3012 2764 3016
rect 2758 3011 2764 3012
rect 3462 3013 3468 3014
rect 3462 3009 3463 3013
rect 3467 3009 3468 3013
rect 3462 3008 3468 3009
rect 2398 3007 2404 3008
rect 2208 3004 2273 3006
rect 2198 3002 2204 3003
rect 2398 3003 2399 3007
rect 2403 3003 2404 3007
rect 2398 3002 2404 3003
rect 2510 3007 2516 3008
rect 2510 3003 2511 3007
rect 2515 3003 2516 3007
rect 2510 3002 2516 3003
rect 2614 3007 2620 3008
rect 2614 3003 2615 3007
rect 2619 3003 2620 3007
rect 2750 3007 2756 3008
rect 2750 3006 2751 3007
rect 2721 3004 2751 3006
rect 2614 3002 2620 3003
rect 2750 3003 2751 3004
rect 2755 3003 2756 3007
rect 2750 3002 2756 3003
rect 2822 3007 2828 3008
rect 2822 3003 2823 3007
rect 2827 3003 2828 3007
rect 2822 3002 2828 3003
rect 2022 2997 2028 2998
rect 1806 2996 1812 2997
rect 187 2995 193 2996
rect 187 2991 188 2995
rect 192 2994 193 2995
rect 334 2995 340 2996
rect 192 2992 330 2994
rect 192 2991 193 2992
rect 187 2990 193 2991
rect 328 2986 330 2992
rect 334 2991 335 2995
rect 339 2994 340 2995
rect 379 2995 385 2996
rect 379 2994 380 2995
rect 339 2992 380 2994
rect 339 2991 340 2992
rect 334 2990 340 2991
rect 379 2991 380 2992
rect 384 2991 385 2995
rect 379 2990 385 2991
rect 398 2995 404 2996
rect 398 2991 399 2995
rect 403 2994 404 2995
rect 587 2995 593 2996
rect 587 2994 588 2995
rect 403 2992 588 2994
rect 403 2991 404 2992
rect 398 2990 404 2991
rect 587 2991 588 2992
rect 592 2991 593 2995
rect 587 2990 593 2991
rect 710 2995 716 2996
rect 710 2991 711 2995
rect 715 2994 716 2995
rect 787 2995 793 2996
rect 787 2994 788 2995
rect 715 2992 788 2994
rect 715 2991 716 2992
rect 710 2990 716 2991
rect 787 2991 788 2992
rect 792 2991 793 2995
rect 787 2990 793 2991
rect 979 2995 985 2996
rect 979 2991 980 2995
rect 984 2994 985 2995
rect 1006 2995 1012 2996
rect 1006 2994 1007 2995
rect 984 2992 1007 2994
rect 984 2991 985 2992
rect 979 2990 985 2991
rect 1006 2991 1007 2992
rect 1011 2991 1012 2995
rect 1006 2990 1012 2991
rect 1155 2995 1161 2996
rect 1155 2991 1156 2995
rect 1160 2994 1161 2995
rect 1183 2995 1189 2996
rect 1183 2994 1184 2995
rect 1160 2992 1184 2994
rect 1160 2991 1161 2992
rect 1155 2990 1161 2991
rect 1183 2991 1184 2992
rect 1188 2991 1189 2995
rect 1183 2990 1189 2991
rect 1331 2995 1337 2996
rect 1331 2991 1332 2995
rect 1336 2994 1337 2995
rect 1410 2995 1416 2996
rect 1410 2994 1411 2995
rect 1336 2992 1411 2994
rect 1336 2991 1337 2992
rect 1331 2990 1337 2991
rect 1410 2991 1411 2992
rect 1415 2991 1416 2995
rect 1410 2990 1416 2991
rect 1499 2995 1505 2996
rect 1499 2991 1500 2995
rect 1504 2994 1505 2995
rect 1554 2995 1560 2996
rect 1554 2994 1555 2995
rect 1504 2992 1555 2994
rect 1504 2991 1505 2992
rect 1499 2990 1505 2991
rect 1554 2991 1555 2992
rect 1559 2991 1560 2995
rect 1554 2990 1560 2991
rect 1662 2995 1668 2996
rect 1662 2991 1663 2995
rect 1667 2994 1668 2995
rect 1675 2995 1681 2996
rect 1675 2994 1676 2995
rect 1667 2992 1676 2994
rect 1667 2991 1668 2992
rect 1662 2990 1668 2991
rect 1675 2991 1676 2992
rect 1680 2991 1681 2995
rect 1806 2992 1807 2996
rect 1811 2992 1812 2996
rect 2022 2993 2023 2997
rect 2027 2993 2028 2997
rect 2022 2992 2028 2993
rect 2126 2997 2132 2998
rect 2126 2993 2127 2997
rect 2131 2993 2132 2997
rect 2126 2992 2132 2993
rect 2230 2997 2236 2998
rect 2230 2993 2231 2997
rect 2235 2993 2236 2997
rect 2230 2992 2236 2993
rect 2334 2997 2340 2998
rect 2334 2993 2335 2997
rect 2339 2993 2340 2997
rect 2334 2992 2340 2993
rect 2438 2997 2444 2998
rect 2438 2993 2439 2997
rect 2443 2993 2444 2997
rect 2438 2992 2444 2993
rect 2542 2997 2548 2998
rect 2542 2993 2543 2997
rect 2547 2993 2548 2997
rect 2542 2992 2548 2993
rect 2646 2997 2652 2998
rect 2646 2993 2647 2997
rect 2651 2993 2652 2997
rect 2646 2992 2652 2993
rect 2758 2997 2764 2998
rect 2758 2993 2759 2997
rect 2763 2993 2764 2997
rect 2758 2992 2764 2993
rect 3462 2996 3468 2997
rect 3462 2992 3463 2996
rect 3467 2992 3468 2996
rect 1806 2991 1812 2992
rect 3462 2991 3468 2992
rect 1675 2990 1681 2991
rect 328 2984 730 2986
rect 134 2980 140 2981
rect 110 2977 116 2978
rect 110 2973 111 2977
rect 115 2973 116 2977
rect 134 2976 135 2980
rect 139 2976 140 2980
rect 134 2975 140 2976
rect 326 2980 332 2981
rect 326 2976 327 2980
rect 331 2976 332 2980
rect 326 2975 332 2976
rect 534 2980 540 2981
rect 534 2976 535 2980
rect 539 2976 540 2980
rect 534 2975 540 2976
rect 110 2972 116 2973
rect 198 2971 204 2972
rect 198 2967 199 2971
rect 203 2967 204 2971
rect 198 2966 204 2967
rect 398 2971 404 2972
rect 398 2967 399 2971
rect 403 2967 404 2971
rect 710 2971 716 2972
rect 710 2970 711 2971
rect 609 2968 711 2970
rect 398 2966 404 2967
rect 710 2967 711 2968
rect 715 2967 716 2971
rect 728 2970 730 2984
rect 734 2980 740 2981
rect 734 2976 735 2980
rect 739 2976 740 2980
rect 734 2975 740 2976
rect 926 2980 932 2981
rect 926 2976 927 2980
rect 931 2976 932 2980
rect 926 2975 932 2976
rect 1102 2980 1108 2981
rect 1102 2976 1103 2980
rect 1107 2976 1108 2980
rect 1102 2975 1108 2976
rect 1278 2980 1284 2981
rect 1278 2976 1279 2980
rect 1283 2976 1284 2980
rect 1278 2975 1284 2976
rect 1446 2980 1452 2981
rect 1446 2976 1447 2980
rect 1451 2976 1452 2980
rect 1446 2975 1452 2976
rect 1622 2980 1628 2981
rect 1622 2976 1623 2980
rect 1627 2976 1628 2980
rect 1622 2975 1628 2976
rect 1766 2977 1772 2978
rect 1766 2973 1767 2977
rect 1771 2973 1772 2977
rect 1766 2972 1772 2973
rect 998 2971 1004 2972
rect 728 2968 777 2970
rect 710 2966 716 2967
rect 998 2967 999 2971
rect 1003 2967 1004 2971
rect 998 2966 1004 2967
rect 1006 2971 1012 2972
rect 1006 2967 1007 2971
rect 1011 2970 1012 2971
rect 1183 2971 1189 2972
rect 1011 2968 1145 2970
rect 1011 2967 1012 2968
rect 1006 2966 1012 2967
rect 1183 2967 1184 2971
rect 1188 2970 1189 2971
rect 1410 2971 1416 2972
rect 1188 2968 1321 2970
rect 1188 2967 1189 2968
rect 1183 2966 1189 2967
rect 1410 2967 1411 2971
rect 1415 2970 1416 2971
rect 1554 2971 1560 2972
rect 1415 2968 1489 2970
rect 1415 2967 1416 2968
rect 1410 2966 1416 2967
rect 1554 2967 1555 2971
rect 1559 2970 1560 2971
rect 1559 2968 1665 2970
rect 1559 2967 1560 2968
rect 1554 2966 1560 2967
rect 134 2961 140 2962
rect 110 2960 116 2961
rect 110 2956 111 2960
rect 115 2956 116 2960
rect 134 2957 135 2961
rect 139 2957 140 2961
rect 134 2956 140 2957
rect 326 2961 332 2962
rect 326 2957 327 2961
rect 331 2957 332 2961
rect 326 2956 332 2957
rect 534 2961 540 2962
rect 534 2957 535 2961
rect 539 2957 540 2961
rect 534 2956 540 2957
rect 734 2961 740 2962
rect 734 2957 735 2961
rect 739 2957 740 2961
rect 734 2956 740 2957
rect 926 2961 932 2962
rect 926 2957 927 2961
rect 931 2957 932 2961
rect 926 2956 932 2957
rect 1102 2961 1108 2962
rect 1102 2957 1103 2961
rect 1107 2957 1108 2961
rect 1102 2956 1108 2957
rect 1278 2961 1284 2962
rect 1278 2957 1279 2961
rect 1283 2957 1284 2961
rect 1278 2956 1284 2957
rect 1446 2961 1452 2962
rect 1446 2957 1447 2961
rect 1451 2957 1452 2961
rect 1446 2956 1452 2957
rect 1622 2961 1628 2962
rect 1622 2957 1623 2961
rect 1627 2957 1628 2961
rect 1622 2956 1628 2957
rect 1766 2960 1772 2961
rect 1766 2956 1767 2960
rect 1771 2956 1772 2960
rect 110 2955 116 2956
rect 1766 2955 1772 2956
rect 1806 2952 1812 2953
rect 3462 2952 3468 2953
rect 1806 2948 1807 2952
rect 1811 2948 1812 2952
rect 1806 2947 1812 2948
rect 2054 2951 2060 2952
rect 2054 2947 2055 2951
rect 2059 2947 2060 2951
rect 2134 2951 2140 2952
rect 2134 2950 2135 2951
rect 2054 2946 2060 2947
rect 2128 2948 2135 2950
rect 2128 2941 2130 2948
rect 2134 2947 2135 2948
rect 2139 2947 2140 2951
rect 2134 2946 2140 2947
rect 2142 2951 2148 2952
rect 2142 2947 2143 2951
rect 2147 2947 2148 2951
rect 2142 2946 2148 2947
rect 2230 2951 2236 2952
rect 2230 2947 2231 2951
rect 2235 2947 2236 2951
rect 2230 2946 2236 2947
rect 2318 2951 2324 2952
rect 2318 2947 2319 2951
rect 2323 2947 2324 2951
rect 2318 2946 2324 2947
rect 2406 2951 2412 2952
rect 2406 2947 2407 2951
rect 2411 2947 2412 2951
rect 2406 2946 2412 2947
rect 2494 2951 2500 2952
rect 2494 2947 2495 2951
rect 2499 2947 2500 2951
rect 2494 2946 2500 2947
rect 2582 2951 2588 2952
rect 2582 2947 2583 2951
rect 2587 2947 2588 2951
rect 2582 2946 2588 2947
rect 2670 2951 2676 2952
rect 2670 2947 2671 2951
rect 2675 2947 2676 2951
rect 2670 2946 2676 2947
rect 2758 2951 2764 2952
rect 2758 2947 2759 2951
rect 2763 2947 2764 2951
rect 2758 2946 2764 2947
rect 2846 2951 2852 2952
rect 2846 2947 2847 2951
rect 2851 2947 2852 2951
rect 3462 2948 3463 2952
rect 3467 2948 3468 2952
rect 3462 2947 3468 2948
rect 2846 2946 2852 2947
rect 2134 2943 2140 2944
rect 2134 2939 2135 2943
rect 2139 2942 2140 2943
rect 2662 2943 2668 2944
rect 2139 2940 2185 2942
rect 2139 2939 2140 2940
rect 2134 2938 2140 2939
rect 2302 2939 2308 2940
rect 1806 2935 1812 2936
rect 1806 2931 1807 2935
rect 1811 2931 1812 2935
rect 2302 2935 2303 2939
rect 2307 2935 2308 2939
rect 2302 2934 2308 2935
rect 2390 2939 2396 2940
rect 2390 2935 2391 2939
rect 2395 2935 2396 2939
rect 2390 2934 2396 2935
rect 2478 2939 2484 2940
rect 2478 2935 2479 2939
rect 2483 2935 2484 2939
rect 2478 2934 2484 2935
rect 2566 2939 2572 2940
rect 2566 2935 2567 2939
rect 2571 2935 2572 2939
rect 2566 2934 2572 2935
rect 2654 2939 2660 2940
rect 2654 2935 2655 2939
rect 2659 2935 2660 2939
rect 2662 2939 2663 2943
rect 2667 2942 2668 2943
rect 2750 2943 2756 2944
rect 2667 2940 2713 2942
rect 2667 2939 2668 2940
rect 2662 2938 2668 2939
rect 2750 2939 2751 2943
rect 2755 2942 2756 2943
rect 2838 2943 2844 2944
rect 2755 2940 2801 2942
rect 2755 2939 2756 2940
rect 2750 2938 2756 2939
rect 2838 2939 2839 2943
rect 2843 2942 2844 2943
rect 2843 2940 2889 2942
rect 2843 2939 2844 2940
rect 2838 2938 2844 2939
rect 2654 2934 2660 2935
rect 3462 2935 3468 2936
rect 1806 2930 1812 2931
rect 2054 2932 2060 2933
rect 2054 2928 2055 2932
rect 2059 2928 2060 2932
rect 2054 2927 2060 2928
rect 2142 2932 2148 2933
rect 2142 2928 2143 2932
rect 2147 2928 2148 2932
rect 2142 2927 2148 2928
rect 2230 2932 2236 2933
rect 2230 2928 2231 2932
rect 2235 2928 2236 2932
rect 2230 2927 2236 2928
rect 2318 2932 2324 2933
rect 2318 2928 2319 2932
rect 2323 2928 2324 2932
rect 2318 2927 2324 2928
rect 2406 2932 2412 2933
rect 2406 2928 2407 2932
rect 2411 2928 2412 2932
rect 2406 2927 2412 2928
rect 2494 2932 2500 2933
rect 2494 2928 2495 2932
rect 2499 2928 2500 2932
rect 2494 2927 2500 2928
rect 2582 2932 2588 2933
rect 2582 2928 2583 2932
rect 2587 2928 2588 2932
rect 2582 2927 2588 2928
rect 2670 2932 2676 2933
rect 2670 2928 2671 2932
rect 2675 2928 2676 2932
rect 2670 2927 2676 2928
rect 2758 2932 2764 2933
rect 2758 2928 2759 2932
rect 2763 2928 2764 2932
rect 2758 2927 2764 2928
rect 2846 2932 2852 2933
rect 2846 2928 2847 2932
rect 2851 2928 2852 2932
rect 3462 2931 3463 2935
rect 3467 2931 3468 2935
rect 3462 2930 3468 2931
rect 2846 2927 2852 2928
rect 2750 2923 2756 2924
rect 2750 2922 2751 2923
rect 2284 2920 2751 2922
rect 2284 2918 2286 2920
rect 2750 2919 2751 2920
rect 2755 2919 2756 2923
rect 2750 2918 2756 2919
rect 2283 2917 2289 2918
rect 2107 2915 2113 2916
rect 2107 2911 2108 2915
rect 2112 2914 2113 2915
rect 2134 2915 2140 2916
rect 2134 2914 2135 2915
rect 2112 2912 2135 2914
rect 2112 2911 2113 2912
rect 2107 2910 2113 2911
rect 2134 2911 2135 2912
rect 2139 2911 2140 2915
rect 2134 2910 2140 2911
rect 2195 2915 2201 2916
rect 2195 2911 2196 2915
rect 2200 2914 2201 2915
rect 2254 2915 2260 2916
rect 2254 2914 2255 2915
rect 2200 2912 2255 2914
rect 2200 2911 2201 2912
rect 2195 2910 2201 2911
rect 2254 2911 2255 2912
rect 2259 2911 2260 2915
rect 2283 2913 2284 2917
rect 2288 2913 2289 2917
rect 2283 2912 2289 2913
rect 2371 2915 2377 2916
rect 2254 2910 2260 2911
rect 2371 2911 2372 2915
rect 2376 2914 2377 2915
rect 2398 2915 2404 2916
rect 2398 2914 2399 2915
rect 2376 2912 2399 2914
rect 2376 2911 2377 2912
rect 2371 2910 2377 2911
rect 2398 2911 2399 2912
rect 2403 2911 2404 2915
rect 2459 2915 2465 2916
rect 2459 2914 2460 2915
rect 2398 2910 2404 2911
rect 2408 2912 2460 2914
rect 110 2908 116 2909
rect 1766 2908 1772 2909
rect 110 2904 111 2908
rect 115 2904 116 2908
rect 110 2903 116 2904
rect 134 2907 140 2908
rect 134 2903 135 2907
rect 139 2903 140 2907
rect 134 2902 140 2903
rect 262 2907 268 2908
rect 262 2903 263 2907
rect 267 2903 268 2907
rect 262 2902 268 2903
rect 430 2907 436 2908
rect 430 2903 431 2907
rect 435 2903 436 2907
rect 430 2902 436 2903
rect 606 2907 612 2908
rect 606 2903 607 2907
rect 611 2903 612 2907
rect 606 2902 612 2903
rect 782 2907 788 2908
rect 782 2903 783 2907
rect 787 2903 788 2907
rect 782 2902 788 2903
rect 950 2907 956 2908
rect 950 2903 951 2907
rect 955 2903 956 2907
rect 950 2902 956 2903
rect 1110 2907 1116 2908
rect 1110 2903 1111 2907
rect 1115 2903 1116 2907
rect 1110 2902 1116 2903
rect 1270 2907 1276 2908
rect 1270 2903 1271 2907
rect 1275 2903 1276 2907
rect 1270 2902 1276 2903
rect 1430 2907 1436 2908
rect 1430 2903 1431 2907
rect 1435 2903 1436 2907
rect 1430 2902 1436 2903
rect 1590 2907 1596 2908
rect 1590 2903 1591 2907
rect 1595 2903 1596 2907
rect 1766 2904 1767 2908
rect 1771 2904 1772 2908
rect 1766 2903 1772 2904
rect 2302 2907 2308 2908
rect 2302 2903 2303 2907
rect 2307 2906 2308 2907
rect 2408 2906 2410 2912
rect 2459 2911 2460 2912
rect 2464 2911 2465 2915
rect 2459 2910 2465 2911
rect 2478 2915 2484 2916
rect 2478 2911 2479 2915
rect 2483 2914 2484 2915
rect 2547 2915 2553 2916
rect 2547 2914 2548 2915
rect 2483 2912 2548 2914
rect 2483 2911 2484 2912
rect 2478 2910 2484 2911
rect 2547 2911 2548 2912
rect 2552 2911 2553 2915
rect 2547 2910 2553 2911
rect 2566 2915 2572 2916
rect 2566 2911 2567 2915
rect 2571 2914 2572 2915
rect 2635 2915 2641 2916
rect 2635 2914 2636 2915
rect 2571 2912 2636 2914
rect 2571 2911 2572 2912
rect 2566 2910 2572 2911
rect 2635 2911 2636 2912
rect 2640 2911 2641 2915
rect 2635 2910 2641 2911
rect 2654 2915 2660 2916
rect 2654 2911 2655 2915
rect 2659 2914 2660 2915
rect 2723 2915 2729 2916
rect 2723 2914 2724 2915
rect 2659 2912 2724 2914
rect 2659 2911 2660 2912
rect 2654 2910 2660 2911
rect 2723 2911 2724 2912
rect 2728 2911 2729 2915
rect 2723 2910 2729 2911
rect 2811 2915 2817 2916
rect 2811 2911 2812 2915
rect 2816 2914 2817 2915
rect 2838 2915 2844 2916
rect 2838 2914 2839 2915
rect 2816 2912 2839 2914
rect 2816 2911 2817 2912
rect 2811 2910 2817 2911
rect 2838 2911 2839 2912
rect 2843 2911 2844 2915
rect 2838 2910 2844 2911
rect 2854 2915 2860 2916
rect 2854 2911 2855 2915
rect 2859 2914 2860 2915
rect 2899 2915 2905 2916
rect 2899 2914 2900 2915
rect 2859 2912 2900 2914
rect 2859 2911 2860 2912
rect 2854 2910 2860 2911
rect 2899 2911 2900 2912
rect 2904 2911 2905 2915
rect 2899 2910 2905 2911
rect 2307 2904 2410 2906
rect 2307 2903 2308 2904
rect 1590 2902 1596 2903
rect 2302 2902 2308 2903
rect 750 2899 756 2900
rect 206 2895 212 2896
rect 110 2891 116 2892
rect 110 2887 111 2891
rect 115 2887 116 2891
rect 206 2891 207 2895
rect 211 2891 212 2895
rect 206 2890 212 2891
rect 334 2895 340 2896
rect 334 2891 335 2895
rect 339 2891 340 2895
rect 334 2890 340 2891
rect 502 2895 508 2896
rect 502 2891 503 2895
rect 507 2891 508 2895
rect 502 2890 508 2891
rect 678 2895 684 2896
rect 678 2891 679 2895
rect 683 2891 684 2895
rect 750 2895 751 2899
rect 755 2898 756 2899
rect 1662 2899 1668 2900
rect 755 2896 825 2898
rect 755 2895 756 2896
rect 750 2894 756 2895
rect 1022 2895 1028 2896
rect 678 2890 684 2891
rect 1022 2891 1023 2895
rect 1027 2891 1028 2895
rect 1022 2890 1028 2891
rect 1182 2895 1188 2896
rect 1182 2891 1183 2895
rect 1187 2891 1188 2895
rect 1182 2890 1188 2891
rect 1342 2895 1348 2896
rect 1342 2891 1343 2895
rect 1347 2891 1348 2895
rect 1342 2890 1348 2891
rect 1502 2895 1508 2896
rect 1502 2891 1503 2895
rect 1507 2891 1508 2895
rect 1662 2895 1663 2899
rect 1667 2895 1668 2899
rect 1662 2894 1668 2895
rect 2123 2895 2129 2896
rect 2123 2894 2124 2895
rect 2056 2892 2124 2894
rect 1502 2890 1508 2891
rect 1766 2891 1772 2892
rect 110 2886 116 2887
rect 134 2888 140 2889
rect 134 2884 135 2888
rect 139 2884 140 2888
rect 134 2883 140 2884
rect 262 2888 268 2889
rect 262 2884 263 2888
rect 267 2884 268 2888
rect 262 2883 268 2884
rect 430 2888 436 2889
rect 430 2884 431 2888
rect 435 2884 436 2888
rect 430 2883 436 2884
rect 606 2888 612 2889
rect 606 2884 607 2888
rect 611 2884 612 2888
rect 606 2883 612 2884
rect 782 2888 788 2889
rect 782 2884 783 2888
rect 787 2884 788 2888
rect 782 2883 788 2884
rect 950 2888 956 2889
rect 950 2884 951 2888
rect 955 2884 956 2888
rect 950 2883 956 2884
rect 1110 2888 1116 2889
rect 1110 2884 1111 2888
rect 1115 2884 1116 2888
rect 1110 2883 1116 2884
rect 1270 2888 1276 2889
rect 1270 2884 1271 2888
rect 1275 2884 1276 2888
rect 1270 2883 1276 2884
rect 1430 2888 1436 2889
rect 1430 2884 1431 2888
rect 1435 2884 1436 2888
rect 1430 2883 1436 2884
rect 1590 2888 1596 2889
rect 1590 2884 1591 2888
rect 1595 2884 1596 2888
rect 1766 2887 1767 2891
rect 1771 2887 1772 2891
rect 1766 2886 1772 2887
rect 2054 2891 2060 2892
rect 2054 2887 2055 2891
rect 2059 2887 2060 2891
rect 2123 2891 2124 2892
rect 2128 2891 2129 2895
rect 2123 2890 2129 2891
rect 2167 2895 2173 2896
rect 2167 2891 2168 2895
rect 2172 2894 2173 2895
rect 2227 2895 2233 2896
rect 2227 2894 2228 2895
rect 2172 2892 2228 2894
rect 2172 2891 2173 2892
rect 2167 2890 2173 2891
rect 2227 2891 2228 2892
rect 2232 2891 2233 2895
rect 2227 2890 2233 2891
rect 2246 2895 2252 2896
rect 2246 2891 2247 2895
rect 2251 2894 2252 2895
rect 2323 2895 2329 2896
rect 2323 2894 2324 2895
rect 2251 2892 2324 2894
rect 2251 2891 2252 2892
rect 2246 2890 2252 2891
rect 2323 2891 2324 2892
rect 2328 2891 2329 2895
rect 2323 2890 2329 2891
rect 2390 2895 2396 2896
rect 2390 2891 2391 2895
rect 2395 2894 2396 2895
rect 2419 2895 2425 2896
rect 2419 2894 2420 2895
rect 2395 2892 2420 2894
rect 2395 2891 2396 2892
rect 2390 2890 2396 2891
rect 2419 2891 2420 2892
rect 2424 2891 2425 2895
rect 2419 2890 2425 2891
rect 2523 2895 2529 2896
rect 2523 2891 2524 2895
rect 2528 2894 2529 2895
rect 2558 2895 2564 2896
rect 2558 2894 2559 2895
rect 2528 2892 2559 2894
rect 2528 2891 2529 2892
rect 2523 2890 2529 2891
rect 2558 2891 2559 2892
rect 2563 2891 2564 2895
rect 2558 2890 2564 2891
rect 2567 2895 2573 2896
rect 2567 2891 2568 2895
rect 2572 2894 2573 2895
rect 2627 2895 2633 2896
rect 2627 2894 2628 2895
rect 2572 2892 2628 2894
rect 2572 2891 2573 2892
rect 2567 2890 2573 2891
rect 2627 2891 2628 2892
rect 2632 2891 2633 2895
rect 2627 2890 2633 2891
rect 2646 2895 2652 2896
rect 2646 2891 2647 2895
rect 2651 2894 2652 2895
rect 2731 2895 2737 2896
rect 2731 2894 2732 2895
rect 2651 2892 2732 2894
rect 2651 2891 2652 2892
rect 2646 2890 2652 2891
rect 2731 2891 2732 2892
rect 2736 2891 2737 2895
rect 2731 2890 2737 2891
rect 2750 2895 2756 2896
rect 2750 2891 2751 2895
rect 2755 2894 2756 2895
rect 2835 2895 2841 2896
rect 2835 2894 2836 2895
rect 2755 2892 2836 2894
rect 2755 2891 2756 2892
rect 2750 2890 2756 2891
rect 2835 2891 2836 2892
rect 2840 2891 2841 2895
rect 2835 2890 2841 2891
rect 2054 2886 2060 2887
rect 1590 2883 1596 2884
rect 2070 2880 2076 2881
rect 1806 2877 1812 2878
rect 1806 2873 1807 2877
rect 1811 2873 1812 2877
rect 2070 2876 2071 2880
rect 2075 2876 2076 2880
rect 2070 2875 2076 2876
rect 2174 2880 2180 2881
rect 2174 2876 2175 2880
rect 2179 2876 2180 2880
rect 2174 2875 2180 2876
rect 2270 2880 2276 2881
rect 2270 2876 2271 2880
rect 2275 2876 2276 2880
rect 2270 2875 2276 2876
rect 2366 2880 2372 2881
rect 2366 2876 2367 2880
rect 2371 2876 2372 2880
rect 2366 2875 2372 2876
rect 2470 2880 2476 2881
rect 2470 2876 2471 2880
rect 2475 2876 2476 2880
rect 2470 2875 2476 2876
rect 2574 2880 2580 2881
rect 2574 2876 2575 2880
rect 2579 2876 2580 2880
rect 2574 2875 2580 2876
rect 2678 2880 2684 2881
rect 2678 2876 2679 2880
rect 2683 2876 2684 2880
rect 2678 2875 2684 2876
rect 2782 2880 2788 2881
rect 2782 2876 2783 2880
rect 2787 2876 2788 2880
rect 2782 2875 2788 2876
rect 3462 2877 3468 2878
rect 1806 2872 1812 2873
rect 3462 2873 3463 2877
rect 3467 2873 3468 2877
rect 3462 2872 3468 2873
rect 187 2871 193 2872
rect 187 2867 188 2871
rect 192 2870 193 2871
rect 198 2871 204 2872
rect 198 2870 199 2871
rect 192 2868 199 2870
rect 192 2867 193 2868
rect 187 2866 193 2867
rect 198 2867 199 2868
rect 203 2867 204 2871
rect 198 2866 204 2867
rect 206 2871 212 2872
rect 206 2867 207 2871
rect 211 2870 212 2871
rect 315 2871 321 2872
rect 315 2870 316 2871
rect 211 2868 316 2870
rect 211 2867 212 2868
rect 206 2866 212 2867
rect 315 2867 316 2868
rect 320 2867 321 2871
rect 315 2866 321 2867
rect 334 2871 340 2872
rect 334 2867 335 2871
rect 339 2870 340 2871
rect 483 2871 489 2872
rect 483 2870 484 2871
rect 339 2868 484 2870
rect 339 2867 340 2868
rect 334 2866 340 2867
rect 483 2867 484 2868
rect 488 2867 489 2871
rect 483 2866 489 2867
rect 502 2871 508 2872
rect 502 2867 503 2871
rect 507 2870 508 2871
rect 659 2871 665 2872
rect 659 2870 660 2871
rect 507 2868 660 2870
rect 507 2867 508 2868
rect 502 2866 508 2867
rect 659 2867 660 2868
rect 664 2867 665 2871
rect 659 2866 665 2867
rect 678 2871 684 2872
rect 678 2867 679 2871
rect 683 2870 684 2871
rect 835 2871 841 2872
rect 835 2870 836 2871
rect 683 2868 836 2870
rect 683 2867 684 2868
rect 678 2866 684 2867
rect 835 2867 836 2868
rect 840 2867 841 2871
rect 835 2866 841 2867
rect 1003 2871 1009 2872
rect 1003 2867 1004 2871
rect 1008 2870 1009 2871
rect 1022 2871 1028 2872
rect 1008 2868 1018 2870
rect 1008 2867 1009 2868
rect 1003 2866 1009 2867
rect 750 2863 756 2864
rect 750 2862 751 2863
rect 188 2860 751 2862
rect 188 2858 190 2860
rect 750 2859 751 2860
rect 755 2859 756 2863
rect 1016 2862 1018 2868
rect 1022 2867 1023 2871
rect 1027 2870 1028 2871
rect 1163 2871 1169 2872
rect 1163 2870 1164 2871
rect 1027 2868 1164 2870
rect 1027 2867 1028 2868
rect 1022 2866 1028 2867
rect 1163 2867 1164 2868
rect 1168 2867 1169 2871
rect 1163 2866 1169 2867
rect 1182 2871 1188 2872
rect 1182 2867 1183 2871
rect 1187 2870 1188 2871
rect 1323 2871 1329 2872
rect 1323 2870 1324 2871
rect 1187 2868 1324 2870
rect 1187 2867 1188 2868
rect 1182 2866 1188 2867
rect 1323 2867 1324 2868
rect 1328 2867 1329 2871
rect 1323 2866 1329 2867
rect 1342 2871 1348 2872
rect 1342 2867 1343 2871
rect 1347 2870 1348 2871
rect 1483 2871 1489 2872
rect 1483 2870 1484 2871
rect 1347 2868 1484 2870
rect 1347 2867 1348 2868
rect 1342 2866 1348 2867
rect 1483 2867 1484 2868
rect 1488 2867 1489 2871
rect 1483 2866 1489 2867
rect 1502 2871 1508 2872
rect 1502 2867 1503 2871
rect 1507 2870 1508 2871
rect 1643 2871 1649 2872
rect 1643 2870 1644 2871
rect 1507 2868 1644 2870
rect 1507 2867 1508 2868
rect 1502 2866 1508 2867
rect 1643 2867 1644 2868
rect 1648 2867 1649 2871
rect 2167 2871 2173 2872
rect 2167 2870 2168 2871
rect 2145 2868 2168 2870
rect 1643 2866 1649 2867
rect 2167 2867 2168 2868
rect 2172 2867 2173 2871
rect 2167 2866 2173 2867
rect 2246 2871 2252 2872
rect 2246 2867 2247 2871
rect 2251 2867 2252 2871
rect 2246 2866 2252 2867
rect 2254 2871 2260 2872
rect 2254 2867 2255 2871
rect 2259 2870 2260 2871
rect 2430 2871 2436 2872
rect 2259 2868 2313 2870
rect 2259 2867 2260 2868
rect 2254 2866 2260 2867
rect 2430 2867 2431 2871
rect 2435 2867 2436 2871
rect 2567 2871 2573 2872
rect 2567 2870 2568 2871
rect 2545 2868 2568 2870
rect 2430 2866 2436 2867
rect 2567 2867 2568 2868
rect 2572 2867 2573 2871
rect 2567 2866 2573 2867
rect 2646 2871 2652 2872
rect 2646 2867 2647 2871
rect 2651 2867 2652 2871
rect 2646 2866 2652 2867
rect 2750 2871 2756 2872
rect 2750 2867 2751 2871
rect 2755 2867 2756 2871
rect 2750 2866 2756 2867
rect 2854 2871 2860 2872
rect 2854 2867 2855 2871
rect 2859 2867 2860 2871
rect 2854 2866 2860 2867
rect 1398 2863 1404 2864
rect 1398 2862 1399 2863
rect 1016 2860 1399 2862
rect 750 2858 756 2859
rect 1398 2859 1399 2860
rect 1403 2859 1404 2863
rect 2070 2861 2076 2862
rect 1398 2858 1404 2859
rect 1806 2860 1812 2861
rect 187 2857 193 2858
rect 187 2853 188 2857
rect 192 2853 193 2857
rect 1806 2856 1807 2860
rect 1811 2856 1812 2860
rect 2070 2857 2071 2861
rect 2075 2857 2076 2861
rect 2070 2856 2076 2857
rect 2174 2861 2180 2862
rect 2174 2857 2175 2861
rect 2179 2857 2180 2861
rect 2174 2856 2180 2857
rect 2270 2861 2276 2862
rect 2270 2857 2271 2861
rect 2275 2857 2276 2861
rect 2270 2856 2276 2857
rect 2366 2861 2372 2862
rect 2366 2857 2367 2861
rect 2371 2857 2372 2861
rect 2366 2856 2372 2857
rect 2470 2861 2476 2862
rect 2470 2857 2471 2861
rect 2475 2857 2476 2861
rect 2470 2856 2476 2857
rect 2574 2861 2580 2862
rect 2574 2857 2575 2861
rect 2579 2857 2580 2861
rect 2574 2856 2580 2857
rect 2678 2861 2684 2862
rect 2678 2857 2679 2861
rect 2683 2857 2684 2861
rect 2678 2856 2684 2857
rect 2782 2861 2788 2862
rect 2782 2857 2783 2861
rect 2787 2857 2788 2861
rect 2782 2856 2788 2857
rect 3462 2860 3468 2861
rect 3462 2856 3463 2860
rect 3467 2856 3468 2860
rect 187 2852 193 2853
rect 206 2855 212 2856
rect 206 2851 207 2855
rect 211 2854 212 2855
rect 307 2855 313 2856
rect 307 2854 308 2855
rect 211 2852 308 2854
rect 211 2851 212 2852
rect 206 2850 212 2851
rect 307 2851 308 2852
rect 312 2851 313 2855
rect 307 2850 313 2851
rect 326 2855 332 2856
rect 326 2851 327 2855
rect 331 2854 332 2855
rect 459 2855 465 2856
rect 459 2854 460 2855
rect 331 2852 460 2854
rect 331 2851 332 2852
rect 326 2850 332 2851
rect 459 2851 460 2852
rect 464 2851 465 2855
rect 459 2850 465 2851
rect 478 2855 484 2856
rect 478 2851 479 2855
rect 483 2854 484 2855
rect 619 2855 625 2856
rect 619 2854 620 2855
rect 483 2852 620 2854
rect 483 2851 484 2852
rect 478 2850 484 2851
rect 619 2851 620 2852
rect 624 2851 625 2855
rect 619 2850 625 2851
rect 638 2855 644 2856
rect 638 2851 639 2855
rect 643 2854 644 2855
rect 779 2855 785 2856
rect 779 2854 780 2855
rect 643 2852 780 2854
rect 643 2851 644 2852
rect 638 2850 644 2851
rect 779 2851 780 2852
rect 784 2851 785 2855
rect 779 2850 785 2851
rect 931 2855 937 2856
rect 931 2851 932 2855
rect 936 2854 937 2855
rect 998 2855 1004 2856
rect 936 2852 994 2854
rect 936 2851 937 2852
rect 931 2850 937 2851
rect 992 2846 994 2852
rect 998 2851 999 2855
rect 1003 2854 1004 2855
rect 1075 2855 1081 2856
rect 1075 2854 1076 2855
rect 1003 2852 1076 2854
rect 1003 2851 1004 2852
rect 998 2850 1004 2851
rect 1075 2851 1076 2852
rect 1080 2851 1081 2855
rect 1075 2850 1081 2851
rect 1094 2855 1100 2856
rect 1094 2851 1095 2855
rect 1099 2854 1100 2855
rect 1219 2855 1225 2856
rect 1219 2854 1220 2855
rect 1099 2852 1220 2854
rect 1099 2851 1100 2852
rect 1094 2850 1100 2851
rect 1219 2851 1220 2852
rect 1224 2851 1225 2855
rect 1219 2850 1225 2851
rect 1238 2855 1244 2856
rect 1238 2851 1239 2855
rect 1243 2854 1244 2855
rect 1363 2855 1369 2856
rect 1363 2854 1364 2855
rect 1243 2852 1364 2854
rect 1243 2851 1244 2852
rect 1238 2850 1244 2851
rect 1363 2851 1364 2852
rect 1368 2851 1369 2855
rect 1363 2850 1369 2851
rect 1382 2855 1388 2856
rect 1382 2851 1383 2855
rect 1387 2854 1388 2855
rect 1515 2855 1521 2856
rect 1806 2855 1812 2856
rect 3462 2855 3468 2856
rect 1515 2854 1516 2855
rect 1387 2852 1516 2854
rect 1387 2851 1388 2852
rect 1382 2850 1388 2851
rect 1515 2851 1516 2852
rect 1520 2851 1521 2855
rect 1515 2850 1521 2851
rect 1278 2847 1284 2848
rect 1278 2846 1279 2847
rect 992 2844 1279 2846
rect 1278 2843 1279 2844
rect 1283 2843 1284 2847
rect 1278 2842 1284 2843
rect 134 2840 140 2841
rect 110 2837 116 2838
rect 110 2833 111 2837
rect 115 2833 116 2837
rect 134 2836 135 2840
rect 139 2836 140 2840
rect 134 2835 140 2836
rect 254 2840 260 2841
rect 254 2836 255 2840
rect 259 2836 260 2840
rect 254 2835 260 2836
rect 406 2840 412 2841
rect 406 2836 407 2840
rect 411 2836 412 2840
rect 406 2835 412 2836
rect 566 2840 572 2841
rect 566 2836 567 2840
rect 571 2836 572 2840
rect 566 2835 572 2836
rect 726 2840 732 2841
rect 726 2836 727 2840
rect 731 2836 732 2840
rect 726 2835 732 2836
rect 878 2840 884 2841
rect 878 2836 879 2840
rect 883 2836 884 2840
rect 878 2835 884 2836
rect 1022 2840 1028 2841
rect 1022 2836 1023 2840
rect 1027 2836 1028 2840
rect 1022 2835 1028 2836
rect 1166 2840 1172 2841
rect 1166 2836 1167 2840
rect 1171 2836 1172 2840
rect 1166 2835 1172 2836
rect 1310 2840 1316 2841
rect 1310 2836 1311 2840
rect 1315 2836 1316 2840
rect 1310 2835 1316 2836
rect 1462 2840 1468 2841
rect 1462 2836 1463 2840
rect 1467 2836 1468 2840
rect 1462 2835 1468 2836
rect 1766 2837 1772 2838
rect 110 2832 116 2833
rect 1766 2833 1767 2837
rect 1771 2833 1772 2837
rect 1766 2832 1772 2833
rect 206 2831 212 2832
rect 206 2827 207 2831
rect 211 2827 212 2831
rect 206 2826 212 2827
rect 326 2831 332 2832
rect 326 2827 327 2831
rect 331 2827 332 2831
rect 326 2826 332 2827
rect 478 2831 484 2832
rect 478 2827 479 2831
rect 483 2827 484 2831
rect 478 2826 484 2827
rect 638 2831 644 2832
rect 638 2827 639 2831
rect 643 2827 644 2831
rect 638 2826 644 2827
rect 646 2831 652 2832
rect 646 2827 647 2831
rect 651 2830 652 2831
rect 998 2831 1004 2832
rect 998 2830 999 2831
rect 651 2828 769 2830
rect 953 2828 999 2830
rect 651 2827 652 2828
rect 646 2826 652 2827
rect 998 2827 999 2828
rect 1003 2827 1004 2831
rect 998 2826 1004 2827
rect 1094 2831 1100 2832
rect 1094 2827 1095 2831
rect 1099 2827 1100 2831
rect 1094 2826 1100 2827
rect 1238 2831 1244 2832
rect 1238 2827 1239 2831
rect 1243 2827 1244 2831
rect 1238 2826 1244 2827
rect 1382 2831 1388 2832
rect 1382 2827 1383 2831
rect 1387 2827 1388 2831
rect 1382 2826 1388 2827
rect 1398 2831 1404 2832
rect 1398 2827 1399 2831
rect 1403 2830 1404 2831
rect 1403 2828 1505 2830
rect 1403 2827 1404 2828
rect 1398 2826 1404 2827
rect 134 2821 140 2822
rect 110 2820 116 2821
rect 110 2816 111 2820
rect 115 2816 116 2820
rect 134 2817 135 2821
rect 139 2817 140 2821
rect 134 2816 140 2817
rect 254 2821 260 2822
rect 254 2817 255 2821
rect 259 2817 260 2821
rect 254 2816 260 2817
rect 406 2821 412 2822
rect 406 2817 407 2821
rect 411 2817 412 2821
rect 406 2816 412 2817
rect 566 2821 572 2822
rect 566 2817 567 2821
rect 571 2817 572 2821
rect 566 2816 572 2817
rect 726 2821 732 2822
rect 726 2817 727 2821
rect 731 2817 732 2821
rect 726 2816 732 2817
rect 878 2821 884 2822
rect 878 2817 879 2821
rect 883 2817 884 2821
rect 878 2816 884 2817
rect 1022 2821 1028 2822
rect 1022 2817 1023 2821
rect 1027 2817 1028 2821
rect 1022 2816 1028 2817
rect 1166 2821 1172 2822
rect 1166 2817 1167 2821
rect 1171 2817 1172 2821
rect 1166 2816 1172 2817
rect 1310 2821 1316 2822
rect 1310 2817 1311 2821
rect 1315 2817 1316 2821
rect 1310 2816 1316 2817
rect 1462 2821 1468 2822
rect 1462 2817 1463 2821
rect 1467 2817 1468 2821
rect 1462 2816 1468 2817
rect 1766 2820 1772 2821
rect 1766 2816 1767 2820
rect 1771 2816 1772 2820
rect 110 2815 116 2816
rect 1766 2815 1772 2816
rect 1806 2812 1812 2813
rect 3462 2812 3468 2813
rect 1806 2808 1807 2812
rect 1811 2808 1812 2812
rect 1806 2807 1812 2808
rect 1982 2811 1988 2812
rect 1982 2807 1983 2811
rect 1987 2807 1988 2811
rect 1982 2806 1988 2807
rect 2110 2811 2116 2812
rect 2110 2807 2111 2811
rect 2115 2807 2116 2811
rect 2110 2806 2116 2807
rect 2238 2811 2244 2812
rect 2238 2807 2239 2811
rect 2243 2807 2244 2811
rect 2238 2806 2244 2807
rect 2366 2811 2372 2812
rect 2366 2807 2367 2811
rect 2371 2807 2372 2811
rect 2366 2806 2372 2807
rect 2486 2811 2492 2812
rect 2486 2807 2487 2811
rect 2491 2807 2492 2811
rect 2486 2806 2492 2807
rect 2606 2811 2612 2812
rect 2606 2807 2607 2811
rect 2611 2807 2612 2811
rect 2606 2806 2612 2807
rect 2718 2811 2724 2812
rect 2718 2807 2719 2811
rect 2723 2807 2724 2811
rect 2718 2806 2724 2807
rect 2838 2811 2844 2812
rect 2838 2807 2839 2811
rect 2843 2807 2844 2811
rect 2838 2806 2844 2807
rect 2958 2811 2964 2812
rect 2958 2807 2959 2811
rect 2963 2807 2964 2811
rect 3462 2808 3463 2812
rect 3467 2808 3468 2812
rect 3462 2807 3468 2808
rect 2958 2806 2964 2807
rect 2054 2803 2060 2804
rect 2054 2799 2055 2803
rect 2059 2799 2060 2803
rect 2054 2798 2060 2799
rect 2062 2803 2068 2804
rect 2062 2799 2063 2803
rect 2067 2802 2068 2803
rect 2190 2803 2196 2804
rect 2067 2800 2153 2802
rect 2067 2799 2068 2800
rect 2062 2798 2068 2799
rect 2190 2799 2191 2803
rect 2195 2802 2196 2803
rect 2558 2803 2564 2804
rect 2195 2800 2281 2802
rect 2195 2799 2196 2800
rect 2190 2798 2196 2799
rect 2438 2799 2444 2800
rect 1806 2795 1812 2796
rect 1806 2791 1807 2795
rect 1811 2791 1812 2795
rect 2438 2795 2439 2799
rect 2443 2795 2444 2799
rect 2558 2799 2559 2803
rect 2563 2799 2564 2803
rect 2558 2798 2564 2799
rect 2567 2803 2573 2804
rect 2567 2799 2568 2803
rect 2572 2802 2573 2803
rect 2686 2803 2692 2804
rect 2572 2800 2649 2802
rect 2572 2799 2573 2800
rect 2567 2798 2573 2799
rect 2686 2799 2687 2803
rect 2691 2802 2692 2803
rect 2918 2803 2924 2804
rect 2691 2800 2761 2802
rect 2691 2799 2692 2800
rect 2686 2798 2692 2799
rect 2910 2799 2916 2800
rect 2438 2794 2444 2795
rect 2910 2795 2911 2799
rect 2915 2795 2916 2799
rect 2918 2799 2919 2803
rect 2923 2802 2924 2803
rect 2923 2800 3001 2802
rect 2923 2799 2924 2800
rect 2918 2798 2924 2799
rect 2910 2794 2916 2795
rect 3462 2795 3468 2796
rect 1806 2790 1812 2791
rect 1982 2792 1988 2793
rect 1982 2788 1983 2792
rect 1987 2788 1988 2792
rect 1982 2787 1988 2788
rect 2110 2792 2116 2793
rect 2110 2788 2111 2792
rect 2115 2788 2116 2792
rect 2110 2787 2116 2788
rect 2238 2792 2244 2793
rect 2238 2788 2239 2792
rect 2243 2788 2244 2792
rect 2238 2787 2244 2788
rect 2366 2792 2372 2793
rect 2366 2788 2367 2792
rect 2371 2788 2372 2792
rect 2366 2787 2372 2788
rect 2486 2792 2492 2793
rect 2486 2788 2487 2792
rect 2491 2788 2492 2792
rect 2486 2787 2492 2788
rect 2606 2792 2612 2793
rect 2606 2788 2607 2792
rect 2611 2788 2612 2792
rect 2606 2787 2612 2788
rect 2718 2792 2724 2793
rect 2718 2788 2719 2792
rect 2723 2788 2724 2792
rect 2718 2787 2724 2788
rect 2838 2792 2844 2793
rect 2838 2788 2839 2792
rect 2843 2788 2844 2792
rect 2838 2787 2844 2788
rect 2958 2792 2964 2793
rect 2958 2788 2959 2792
rect 2963 2788 2964 2792
rect 3462 2791 3463 2795
rect 3467 2791 3468 2795
rect 3462 2790 3468 2791
rect 2958 2787 2964 2788
rect 2918 2783 2924 2784
rect 2918 2782 2919 2783
rect 2772 2780 2919 2782
rect 2772 2778 2774 2780
rect 2918 2779 2919 2780
rect 2923 2779 2924 2783
rect 2918 2778 2924 2779
rect 2771 2777 2777 2778
rect 2035 2775 2041 2776
rect 2035 2771 2036 2775
rect 2040 2774 2041 2775
rect 2062 2775 2068 2776
rect 2062 2774 2063 2775
rect 2040 2772 2063 2774
rect 2040 2771 2041 2772
rect 2035 2770 2041 2771
rect 2062 2771 2063 2772
rect 2067 2771 2068 2775
rect 2062 2770 2068 2771
rect 2163 2775 2169 2776
rect 2163 2771 2164 2775
rect 2168 2774 2169 2775
rect 2190 2775 2196 2776
rect 2190 2774 2191 2775
rect 2168 2772 2191 2774
rect 2168 2771 2169 2772
rect 2163 2770 2169 2771
rect 2190 2771 2191 2772
rect 2195 2771 2196 2775
rect 2190 2770 2196 2771
rect 2254 2775 2260 2776
rect 2254 2771 2255 2775
rect 2259 2774 2260 2775
rect 2291 2775 2297 2776
rect 2291 2774 2292 2775
rect 2259 2772 2292 2774
rect 2259 2771 2260 2772
rect 2254 2770 2260 2771
rect 2291 2771 2292 2772
rect 2296 2771 2297 2775
rect 2291 2770 2297 2771
rect 2419 2775 2425 2776
rect 2419 2771 2420 2775
rect 2424 2774 2425 2775
rect 2430 2775 2436 2776
rect 2430 2774 2431 2775
rect 2424 2772 2431 2774
rect 2424 2771 2425 2772
rect 2419 2770 2425 2771
rect 2430 2771 2431 2772
rect 2435 2771 2436 2775
rect 2430 2770 2436 2771
rect 2539 2775 2545 2776
rect 2539 2771 2540 2775
rect 2544 2774 2545 2775
rect 2567 2775 2573 2776
rect 2567 2774 2568 2775
rect 2544 2772 2568 2774
rect 2544 2771 2545 2772
rect 2539 2770 2545 2771
rect 2567 2771 2568 2772
rect 2572 2771 2573 2775
rect 2567 2770 2573 2771
rect 2659 2775 2665 2776
rect 2659 2771 2660 2775
rect 2664 2774 2665 2775
rect 2686 2775 2692 2776
rect 2686 2774 2687 2775
rect 2664 2772 2687 2774
rect 2664 2771 2665 2772
rect 2659 2770 2665 2771
rect 2686 2771 2687 2772
rect 2691 2771 2692 2775
rect 2771 2773 2772 2777
rect 2776 2773 2777 2777
rect 2771 2772 2777 2773
rect 2847 2775 2853 2776
rect 2686 2770 2692 2771
rect 2847 2771 2848 2775
rect 2852 2774 2853 2775
rect 2891 2775 2897 2776
rect 2891 2774 2892 2775
rect 2852 2772 2892 2774
rect 2852 2771 2853 2772
rect 2847 2770 2853 2771
rect 2891 2771 2892 2772
rect 2896 2771 2897 2775
rect 2891 2770 2897 2771
rect 2910 2775 2916 2776
rect 2910 2771 2911 2775
rect 2915 2774 2916 2775
rect 3011 2775 3017 2776
rect 3011 2774 3012 2775
rect 2915 2772 3012 2774
rect 2915 2771 2916 2772
rect 2910 2770 2916 2771
rect 3011 2771 3012 2772
rect 3016 2771 3017 2775
rect 3011 2770 3017 2771
rect 110 2768 116 2769
rect 1766 2768 1772 2769
rect 110 2764 111 2768
rect 115 2764 116 2768
rect 110 2763 116 2764
rect 286 2767 292 2768
rect 286 2763 287 2767
rect 291 2763 292 2767
rect 286 2762 292 2763
rect 390 2767 396 2768
rect 390 2763 391 2767
rect 395 2763 396 2767
rect 390 2762 396 2763
rect 502 2767 508 2768
rect 502 2763 503 2767
rect 507 2763 508 2767
rect 502 2762 508 2763
rect 622 2767 628 2768
rect 622 2763 623 2767
rect 627 2763 628 2767
rect 622 2762 628 2763
rect 742 2767 748 2768
rect 742 2763 743 2767
rect 747 2763 748 2767
rect 742 2762 748 2763
rect 854 2767 860 2768
rect 854 2763 855 2767
rect 859 2763 860 2767
rect 854 2762 860 2763
rect 966 2767 972 2768
rect 966 2763 967 2767
rect 971 2763 972 2767
rect 966 2762 972 2763
rect 1078 2767 1084 2768
rect 1078 2763 1079 2767
rect 1083 2763 1084 2767
rect 1078 2762 1084 2763
rect 1198 2767 1204 2768
rect 1198 2763 1199 2767
rect 1203 2763 1204 2767
rect 1198 2762 1204 2763
rect 1318 2767 1324 2768
rect 1318 2763 1319 2767
rect 1323 2763 1324 2767
rect 1766 2764 1767 2768
rect 1771 2764 1772 2768
rect 1766 2763 1772 2764
rect 1318 2762 1324 2763
rect 730 2759 736 2760
rect 358 2755 364 2756
rect 110 2751 116 2752
rect 110 2747 111 2751
rect 115 2747 116 2751
rect 358 2751 359 2755
rect 363 2751 364 2755
rect 358 2750 364 2751
rect 462 2755 468 2756
rect 462 2751 463 2755
rect 467 2751 468 2755
rect 462 2750 468 2751
rect 574 2755 580 2756
rect 574 2751 575 2755
rect 579 2751 580 2755
rect 574 2750 580 2751
rect 694 2755 700 2756
rect 694 2751 695 2755
rect 699 2751 700 2755
rect 730 2755 731 2759
rect 735 2758 736 2759
rect 1278 2759 1284 2760
rect 735 2756 785 2758
rect 735 2755 736 2756
rect 730 2754 736 2755
rect 926 2755 932 2756
rect 694 2750 700 2751
rect 926 2751 927 2755
rect 931 2751 932 2755
rect 926 2750 932 2751
rect 1038 2755 1044 2756
rect 1038 2751 1039 2755
rect 1043 2751 1044 2755
rect 1038 2750 1044 2751
rect 1150 2755 1156 2756
rect 1150 2751 1151 2755
rect 1155 2751 1156 2755
rect 1150 2750 1156 2751
rect 1270 2755 1276 2756
rect 1270 2751 1271 2755
rect 1275 2751 1276 2755
rect 1278 2755 1279 2759
rect 1283 2758 1284 2759
rect 1902 2759 1908 2760
rect 1283 2756 1361 2758
rect 1283 2755 1284 2756
rect 1278 2754 1284 2755
rect 1902 2755 1903 2759
rect 1907 2758 1908 2759
rect 1939 2759 1945 2760
rect 1939 2758 1940 2759
rect 1907 2756 1940 2758
rect 1907 2755 1908 2756
rect 1902 2754 1908 2755
rect 1939 2755 1940 2756
rect 1944 2755 1945 2759
rect 1939 2754 1945 2755
rect 1958 2759 1964 2760
rect 1958 2755 1959 2759
rect 1963 2758 1964 2759
rect 2083 2759 2089 2760
rect 2083 2758 2084 2759
rect 1963 2756 2084 2758
rect 1963 2755 1964 2756
rect 1958 2754 1964 2755
rect 2083 2755 2084 2756
rect 2088 2755 2089 2759
rect 2083 2754 2089 2755
rect 2102 2759 2108 2760
rect 2102 2755 2103 2759
rect 2107 2758 2108 2759
rect 2235 2759 2241 2760
rect 2235 2758 2236 2759
rect 2107 2756 2236 2758
rect 2107 2755 2108 2756
rect 2102 2754 2108 2755
rect 2235 2755 2236 2756
rect 2240 2755 2241 2759
rect 2235 2754 2241 2755
rect 2387 2759 2393 2760
rect 2387 2755 2388 2759
rect 2392 2758 2393 2759
rect 2438 2759 2444 2760
rect 2438 2758 2439 2759
rect 2392 2756 2439 2758
rect 2392 2755 2393 2756
rect 2387 2754 2393 2755
rect 2438 2755 2439 2756
rect 2443 2755 2444 2759
rect 2438 2754 2444 2755
rect 2454 2759 2460 2760
rect 2454 2755 2455 2759
rect 2459 2758 2460 2759
rect 2531 2759 2537 2760
rect 2531 2758 2532 2759
rect 2459 2756 2532 2758
rect 2459 2755 2460 2756
rect 2454 2754 2460 2755
rect 2531 2755 2532 2756
rect 2536 2755 2537 2759
rect 2531 2754 2537 2755
rect 2675 2759 2681 2760
rect 2675 2755 2676 2759
rect 2680 2758 2681 2759
rect 2694 2759 2700 2760
rect 2680 2756 2690 2758
rect 2680 2755 2681 2756
rect 2675 2754 2681 2755
rect 1270 2750 1276 2751
rect 1766 2751 1772 2752
rect 110 2746 116 2747
rect 286 2748 292 2749
rect 286 2744 287 2748
rect 291 2744 292 2748
rect 286 2743 292 2744
rect 390 2748 396 2749
rect 390 2744 391 2748
rect 395 2744 396 2748
rect 390 2743 396 2744
rect 502 2748 508 2749
rect 502 2744 503 2748
rect 507 2744 508 2748
rect 502 2743 508 2744
rect 622 2748 628 2749
rect 622 2744 623 2748
rect 627 2744 628 2748
rect 622 2743 628 2744
rect 742 2748 748 2749
rect 742 2744 743 2748
rect 747 2744 748 2748
rect 742 2743 748 2744
rect 854 2748 860 2749
rect 854 2744 855 2748
rect 859 2744 860 2748
rect 854 2743 860 2744
rect 966 2748 972 2749
rect 966 2744 967 2748
rect 971 2744 972 2748
rect 966 2743 972 2744
rect 1078 2748 1084 2749
rect 1078 2744 1079 2748
rect 1083 2744 1084 2748
rect 1078 2743 1084 2744
rect 1198 2748 1204 2749
rect 1198 2744 1199 2748
rect 1203 2744 1204 2748
rect 1198 2743 1204 2744
rect 1318 2748 1324 2749
rect 1318 2744 1319 2748
rect 1323 2744 1324 2748
rect 1766 2747 1767 2751
rect 1771 2747 1772 2751
rect 2688 2750 2690 2756
rect 2694 2755 2695 2759
rect 2699 2758 2700 2759
rect 2819 2759 2825 2760
rect 2819 2758 2820 2759
rect 2699 2756 2820 2758
rect 2699 2755 2700 2756
rect 2694 2754 2700 2755
rect 2819 2755 2820 2756
rect 2824 2755 2825 2759
rect 2819 2754 2825 2755
rect 2963 2759 2969 2760
rect 2963 2755 2964 2759
rect 2968 2758 2969 2759
rect 2990 2759 2996 2760
rect 2990 2758 2991 2759
rect 2968 2756 2991 2758
rect 2968 2755 2969 2756
rect 2963 2754 2969 2755
rect 2990 2755 2991 2756
rect 2995 2755 2996 2759
rect 2990 2754 2996 2755
rect 3107 2759 3113 2760
rect 3107 2755 3108 2759
rect 3112 2758 3113 2759
rect 3166 2759 3172 2760
rect 3166 2758 3167 2759
rect 3112 2756 3167 2758
rect 3112 2755 3113 2756
rect 3107 2754 3113 2755
rect 3166 2755 3167 2756
rect 3171 2755 3172 2759
rect 3166 2754 3172 2755
rect 2688 2748 2858 2750
rect 1766 2746 1772 2747
rect 1318 2743 1324 2744
rect 1886 2744 1892 2745
rect 1806 2741 1812 2742
rect 646 2739 652 2740
rect 646 2738 647 2739
rect 340 2736 647 2738
rect 340 2734 342 2736
rect 646 2735 647 2736
rect 651 2735 652 2739
rect 1806 2737 1807 2741
rect 1811 2737 1812 2741
rect 1886 2740 1887 2744
rect 1891 2740 1892 2744
rect 1886 2739 1892 2740
rect 2030 2744 2036 2745
rect 2030 2740 2031 2744
rect 2035 2740 2036 2744
rect 2030 2739 2036 2740
rect 2182 2744 2188 2745
rect 2182 2740 2183 2744
rect 2187 2740 2188 2744
rect 2182 2739 2188 2740
rect 2334 2744 2340 2745
rect 2334 2740 2335 2744
rect 2339 2740 2340 2744
rect 2334 2739 2340 2740
rect 2478 2744 2484 2745
rect 2478 2740 2479 2744
rect 2483 2740 2484 2744
rect 2478 2739 2484 2740
rect 2622 2744 2628 2745
rect 2622 2740 2623 2744
rect 2627 2740 2628 2744
rect 2622 2739 2628 2740
rect 2766 2744 2772 2745
rect 2766 2740 2767 2744
rect 2771 2740 2772 2744
rect 2766 2739 2772 2740
rect 1806 2736 1812 2737
rect 646 2734 652 2735
rect 1958 2735 1964 2736
rect 339 2733 345 2734
rect 339 2729 340 2733
rect 344 2729 345 2733
rect 339 2728 345 2729
rect 358 2731 364 2732
rect 358 2727 359 2731
rect 363 2730 364 2731
rect 443 2731 449 2732
rect 443 2730 444 2731
rect 363 2728 444 2730
rect 363 2727 364 2728
rect 358 2726 364 2727
rect 443 2727 444 2728
rect 448 2727 449 2731
rect 443 2726 449 2727
rect 462 2731 468 2732
rect 462 2727 463 2731
rect 467 2730 468 2731
rect 555 2731 561 2732
rect 555 2730 556 2731
rect 467 2728 556 2730
rect 467 2727 468 2728
rect 462 2726 468 2727
rect 555 2727 556 2728
rect 560 2727 561 2731
rect 555 2726 561 2727
rect 574 2731 580 2732
rect 574 2727 575 2731
rect 579 2730 580 2731
rect 675 2731 681 2732
rect 675 2730 676 2731
rect 579 2728 676 2730
rect 579 2727 580 2728
rect 574 2726 580 2727
rect 675 2727 676 2728
rect 680 2727 681 2731
rect 675 2726 681 2727
rect 694 2731 700 2732
rect 694 2727 695 2731
rect 699 2730 700 2731
rect 795 2731 801 2732
rect 795 2730 796 2731
rect 699 2728 796 2730
rect 699 2727 700 2728
rect 694 2726 700 2727
rect 795 2727 796 2728
rect 800 2727 801 2731
rect 795 2726 801 2727
rect 907 2731 913 2732
rect 907 2727 908 2731
rect 912 2730 913 2731
rect 926 2731 932 2732
rect 912 2728 922 2730
rect 912 2727 913 2728
rect 907 2726 913 2727
rect 730 2723 736 2724
rect 730 2722 731 2723
rect 532 2720 731 2722
rect 532 2718 534 2720
rect 730 2719 731 2720
rect 735 2719 736 2723
rect 920 2722 922 2728
rect 926 2727 927 2731
rect 931 2730 932 2731
rect 1019 2731 1025 2732
rect 1019 2730 1020 2731
rect 931 2728 1020 2730
rect 931 2727 932 2728
rect 926 2726 932 2727
rect 1019 2727 1020 2728
rect 1024 2727 1025 2731
rect 1019 2726 1025 2727
rect 1038 2731 1044 2732
rect 1038 2727 1039 2731
rect 1043 2730 1044 2731
rect 1131 2731 1137 2732
rect 1131 2730 1132 2731
rect 1043 2728 1132 2730
rect 1043 2727 1044 2728
rect 1038 2726 1044 2727
rect 1131 2727 1132 2728
rect 1136 2727 1137 2731
rect 1131 2726 1137 2727
rect 1150 2731 1156 2732
rect 1150 2727 1151 2731
rect 1155 2730 1156 2731
rect 1251 2731 1257 2732
rect 1251 2730 1252 2731
rect 1155 2728 1252 2730
rect 1155 2727 1156 2728
rect 1150 2726 1156 2727
rect 1251 2727 1252 2728
rect 1256 2727 1257 2731
rect 1251 2726 1257 2727
rect 1270 2731 1276 2732
rect 1270 2727 1271 2731
rect 1275 2730 1276 2731
rect 1371 2731 1377 2732
rect 1371 2730 1372 2731
rect 1275 2728 1372 2730
rect 1275 2727 1276 2728
rect 1270 2726 1276 2727
rect 1371 2727 1372 2728
rect 1376 2727 1377 2731
rect 1958 2731 1959 2735
rect 1963 2731 1964 2735
rect 1958 2730 1964 2731
rect 2102 2735 2108 2736
rect 2102 2731 2103 2735
rect 2107 2731 2108 2735
rect 2102 2730 2108 2731
rect 2254 2735 2260 2736
rect 2254 2731 2255 2735
rect 2259 2731 2260 2735
rect 2454 2735 2460 2736
rect 2454 2734 2455 2735
rect 2409 2732 2455 2734
rect 2254 2730 2260 2731
rect 2454 2731 2455 2732
rect 2459 2731 2460 2735
rect 2454 2730 2460 2731
rect 2542 2735 2548 2736
rect 2542 2731 2543 2735
rect 2547 2731 2548 2735
rect 2542 2730 2548 2731
rect 2694 2735 2700 2736
rect 2694 2731 2695 2735
rect 2699 2731 2700 2735
rect 2847 2735 2853 2736
rect 2847 2734 2848 2735
rect 2841 2732 2848 2734
rect 2694 2730 2700 2731
rect 2847 2731 2848 2732
rect 2852 2731 2853 2735
rect 2856 2734 2858 2748
rect 2910 2744 2916 2745
rect 2910 2740 2911 2744
rect 2915 2740 2916 2744
rect 2910 2739 2916 2740
rect 3054 2744 3060 2745
rect 3054 2740 3055 2744
rect 3059 2740 3060 2744
rect 3054 2739 3060 2740
rect 3462 2741 3468 2742
rect 3462 2737 3463 2741
rect 3467 2737 3468 2741
rect 3462 2736 3468 2737
rect 2990 2735 2996 2736
rect 2856 2732 2953 2734
rect 2847 2730 2853 2731
rect 2990 2731 2991 2735
rect 2995 2734 2996 2735
rect 2995 2732 3097 2734
rect 2995 2731 2996 2732
rect 2990 2730 2996 2731
rect 1371 2726 1377 2727
rect 1886 2725 1892 2726
rect 1806 2724 1812 2725
rect 1174 2723 1180 2724
rect 1174 2722 1175 2723
rect 920 2720 1175 2722
rect 730 2718 736 2719
rect 1174 2719 1175 2720
rect 1179 2719 1180 2723
rect 1806 2720 1807 2724
rect 1811 2720 1812 2724
rect 1886 2721 1887 2725
rect 1891 2721 1892 2725
rect 1886 2720 1892 2721
rect 2030 2725 2036 2726
rect 2030 2721 2031 2725
rect 2035 2721 2036 2725
rect 2030 2720 2036 2721
rect 2182 2725 2188 2726
rect 2182 2721 2183 2725
rect 2187 2721 2188 2725
rect 2182 2720 2188 2721
rect 2334 2725 2340 2726
rect 2334 2721 2335 2725
rect 2339 2721 2340 2725
rect 2334 2720 2340 2721
rect 2478 2725 2484 2726
rect 2478 2721 2479 2725
rect 2483 2721 2484 2725
rect 2478 2720 2484 2721
rect 2622 2725 2628 2726
rect 2622 2721 2623 2725
rect 2627 2721 2628 2725
rect 2622 2720 2628 2721
rect 2766 2725 2772 2726
rect 2766 2721 2767 2725
rect 2771 2721 2772 2725
rect 2766 2720 2772 2721
rect 2910 2725 2916 2726
rect 2910 2721 2911 2725
rect 2915 2721 2916 2725
rect 2910 2720 2916 2721
rect 3054 2725 3060 2726
rect 3054 2721 3055 2725
rect 3059 2721 3060 2725
rect 3054 2720 3060 2721
rect 3462 2724 3468 2725
rect 3462 2720 3463 2724
rect 3467 2720 3468 2724
rect 1806 2719 1812 2720
rect 3462 2719 3468 2720
rect 1174 2718 1180 2719
rect 531 2717 537 2718
rect 531 2713 532 2717
rect 536 2713 537 2717
rect 531 2712 537 2713
rect 550 2715 556 2716
rect 550 2711 551 2715
rect 555 2714 556 2715
rect 619 2715 625 2716
rect 619 2714 620 2715
rect 555 2712 620 2714
rect 555 2711 556 2712
rect 550 2710 556 2711
rect 619 2711 620 2712
rect 624 2711 625 2715
rect 619 2710 625 2711
rect 638 2715 644 2716
rect 638 2711 639 2715
rect 643 2714 644 2715
rect 707 2715 713 2716
rect 707 2714 708 2715
rect 643 2712 708 2714
rect 643 2711 644 2712
rect 638 2710 644 2711
rect 707 2711 708 2712
rect 712 2711 713 2715
rect 707 2710 713 2711
rect 726 2715 732 2716
rect 726 2711 727 2715
rect 731 2714 732 2715
rect 795 2715 801 2716
rect 795 2714 796 2715
rect 731 2712 796 2714
rect 731 2711 732 2712
rect 726 2710 732 2711
rect 795 2711 796 2712
rect 800 2711 801 2715
rect 795 2710 801 2711
rect 814 2715 820 2716
rect 814 2711 815 2715
rect 819 2714 820 2715
rect 883 2715 889 2716
rect 883 2714 884 2715
rect 819 2712 884 2714
rect 819 2711 820 2712
rect 814 2710 820 2711
rect 883 2711 884 2712
rect 888 2711 889 2715
rect 883 2710 889 2711
rect 971 2715 977 2716
rect 971 2711 972 2715
rect 976 2711 977 2715
rect 971 2710 977 2711
rect 990 2715 996 2716
rect 990 2711 991 2715
rect 995 2714 996 2715
rect 1059 2715 1065 2716
rect 1059 2714 1060 2715
rect 995 2712 1060 2714
rect 995 2711 996 2712
rect 990 2710 996 2711
rect 1059 2711 1060 2712
rect 1064 2711 1065 2715
rect 1059 2710 1065 2711
rect 1087 2715 1093 2716
rect 1087 2711 1088 2715
rect 1092 2714 1093 2715
rect 1147 2715 1153 2716
rect 1147 2714 1148 2715
rect 1092 2712 1148 2714
rect 1092 2711 1093 2712
rect 1087 2710 1093 2711
rect 1147 2711 1148 2712
rect 1152 2711 1153 2715
rect 1147 2710 1153 2711
rect 1166 2715 1172 2716
rect 1166 2711 1167 2715
rect 1171 2714 1172 2715
rect 1235 2715 1241 2716
rect 1235 2714 1236 2715
rect 1171 2712 1236 2714
rect 1171 2711 1172 2712
rect 1166 2710 1172 2711
rect 1235 2711 1236 2712
rect 1240 2711 1241 2715
rect 1235 2710 1241 2711
rect 973 2706 975 2710
rect 1078 2707 1084 2708
rect 1078 2706 1079 2707
rect 973 2704 1079 2706
rect 1078 2703 1079 2704
rect 1083 2703 1084 2707
rect 1078 2702 1084 2703
rect 478 2700 484 2701
rect 110 2697 116 2698
rect 110 2693 111 2697
rect 115 2693 116 2697
rect 478 2696 479 2700
rect 483 2696 484 2700
rect 478 2695 484 2696
rect 566 2700 572 2701
rect 566 2696 567 2700
rect 571 2696 572 2700
rect 566 2695 572 2696
rect 654 2700 660 2701
rect 654 2696 655 2700
rect 659 2696 660 2700
rect 654 2695 660 2696
rect 742 2700 748 2701
rect 742 2696 743 2700
rect 747 2696 748 2700
rect 742 2695 748 2696
rect 830 2700 836 2701
rect 830 2696 831 2700
rect 835 2696 836 2700
rect 830 2695 836 2696
rect 918 2700 924 2701
rect 918 2696 919 2700
rect 923 2696 924 2700
rect 918 2695 924 2696
rect 1006 2700 1012 2701
rect 1006 2696 1007 2700
rect 1011 2696 1012 2700
rect 1006 2695 1012 2696
rect 1094 2700 1100 2701
rect 1094 2696 1095 2700
rect 1099 2696 1100 2700
rect 1094 2695 1100 2696
rect 1182 2700 1188 2701
rect 1182 2696 1183 2700
rect 1187 2696 1188 2700
rect 1182 2695 1188 2696
rect 1766 2697 1772 2698
rect 110 2692 116 2693
rect 1766 2693 1767 2697
rect 1771 2693 1772 2697
rect 1766 2692 1772 2693
rect 550 2691 556 2692
rect 550 2687 551 2691
rect 555 2687 556 2691
rect 550 2686 556 2687
rect 638 2691 644 2692
rect 638 2687 639 2691
rect 643 2687 644 2691
rect 638 2686 644 2687
rect 726 2691 732 2692
rect 726 2687 727 2691
rect 731 2687 732 2691
rect 726 2686 732 2687
rect 814 2691 820 2692
rect 814 2687 815 2691
rect 819 2687 820 2691
rect 814 2686 820 2687
rect 902 2691 908 2692
rect 902 2687 903 2691
rect 907 2687 908 2691
rect 902 2686 908 2687
rect 990 2691 996 2692
rect 990 2687 991 2691
rect 995 2687 996 2691
rect 1087 2691 1093 2692
rect 1087 2690 1088 2691
rect 1081 2688 1088 2690
rect 990 2686 996 2687
rect 1087 2687 1088 2688
rect 1092 2687 1093 2691
rect 1087 2686 1093 2687
rect 1166 2691 1172 2692
rect 1166 2687 1167 2691
rect 1171 2687 1172 2691
rect 1166 2686 1172 2687
rect 1174 2691 1180 2692
rect 1174 2687 1175 2691
rect 1179 2690 1180 2691
rect 1179 2688 1225 2690
rect 1179 2687 1180 2688
rect 1174 2686 1180 2687
rect 478 2681 484 2682
rect 110 2680 116 2681
rect 110 2676 111 2680
rect 115 2676 116 2680
rect 478 2677 479 2681
rect 483 2677 484 2681
rect 478 2676 484 2677
rect 566 2681 572 2682
rect 566 2677 567 2681
rect 571 2677 572 2681
rect 566 2676 572 2677
rect 654 2681 660 2682
rect 654 2677 655 2681
rect 659 2677 660 2681
rect 654 2676 660 2677
rect 742 2681 748 2682
rect 742 2677 743 2681
rect 747 2677 748 2681
rect 742 2676 748 2677
rect 830 2681 836 2682
rect 830 2677 831 2681
rect 835 2677 836 2681
rect 830 2676 836 2677
rect 918 2681 924 2682
rect 918 2677 919 2681
rect 923 2677 924 2681
rect 918 2676 924 2677
rect 1006 2681 1012 2682
rect 1006 2677 1007 2681
rect 1011 2677 1012 2681
rect 1006 2676 1012 2677
rect 1094 2681 1100 2682
rect 1094 2677 1095 2681
rect 1099 2677 1100 2681
rect 1094 2676 1100 2677
rect 1182 2681 1188 2682
rect 1182 2677 1183 2681
rect 1187 2677 1188 2681
rect 1182 2676 1188 2677
rect 1766 2680 1772 2681
rect 1766 2676 1767 2680
rect 1771 2676 1772 2680
rect 110 2675 116 2676
rect 1766 2675 1772 2676
rect 1806 2680 1812 2681
rect 3462 2680 3468 2681
rect 1806 2676 1807 2680
rect 1811 2676 1812 2680
rect 1806 2675 1812 2676
rect 1830 2679 1836 2680
rect 1830 2675 1831 2679
rect 1835 2675 1836 2679
rect 1830 2674 1836 2675
rect 2022 2679 2028 2680
rect 2022 2675 2023 2679
rect 2027 2675 2028 2679
rect 2022 2674 2028 2675
rect 2230 2679 2236 2680
rect 2230 2675 2231 2679
rect 2235 2675 2236 2679
rect 2230 2674 2236 2675
rect 2430 2679 2436 2680
rect 2430 2675 2431 2679
rect 2435 2675 2436 2679
rect 2430 2674 2436 2675
rect 2614 2679 2620 2680
rect 2614 2675 2615 2679
rect 2619 2675 2620 2679
rect 2614 2674 2620 2675
rect 2782 2679 2788 2680
rect 2782 2675 2783 2679
rect 2787 2675 2788 2679
rect 2782 2674 2788 2675
rect 2942 2679 2948 2680
rect 2942 2675 2943 2679
rect 2947 2675 2948 2679
rect 2942 2674 2948 2675
rect 3094 2679 3100 2680
rect 3094 2675 3095 2679
rect 3099 2675 3100 2679
rect 3094 2674 3100 2675
rect 3238 2679 3244 2680
rect 3238 2675 3239 2679
rect 3243 2675 3244 2679
rect 3238 2674 3244 2675
rect 3366 2679 3372 2680
rect 3366 2675 3367 2679
rect 3371 2675 3372 2679
rect 3462 2676 3463 2680
rect 3467 2676 3468 2680
rect 3462 2675 3468 2676
rect 3366 2674 3372 2675
rect 1902 2671 1908 2672
rect 1902 2667 1903 2671
rect 1907 2667 1908 2671
rect 1902 2666 1908 2667
rect 1910 2671 1916 2672
rect 1910 2667 1911 2671
rect 1915 2670 1916 2671
rect 2102 2671 2108 2672
rect 1915 2668 2065 2670
rect 1915 2667 1916 2668
rect 1910 2666 1916 2667
rect 2102 2667 2103 2671
rect 2107 2670 2108 2671
rect 2414 2671 2420 2672
rect 2107 2668 2273 2670
rect 2107 2667 2108 2668
rect 2102 2666 2108 2667
rect 2414 2667 2415 2671
rect 2419 2670 2420 2671
rect 3166 2671 3172 2672
rect 2419 2668 2473 2670
rect 2419 2667 2420 2668
rect 2414 2666 2420 2667
rect 2686 2667 2692 2668
rect 1806 2663 1812 2664
rect 1806 2659 1807 2663
rect 1811 2659 1812 2663
rect 2686 2663 2687 2667
rect 2691 2663 2692 2667
rect 2686 2662 2692 2663
rect 2854 2667 2860 2668
rect 2854 2663 2855 2667
rect 2859 2663 2860 2667
rect 2854 2662 2860 2663
rect 3014 2667 3020 2668
rect 3014 2663 3015 2667
rect 3019 2663 3020 2667
rect 3166 2667 3167 2671
rect 3171 2667 3172 2671
rect 3318 2671 3324 2672
rect 3166 2666 3172 2667
rect 3310 2667 3316 2668
rect 3014 2662 3020 2663
rect 3310 2663 3311 2667
rect 3315 2663 3316 2667
rect 3318 2667 3319 2671
rect 3323 2670 3324 2671
rect 3323 2668 3409 2670
rect 3323 2667 3324 2668
rect 3318 2666 3324 2667
rect 3310 2662 3316 2663
rect 3462 2663 3468 2664
rect 1806 2658 1812 2659
rect 1830 2660 1836 2661
rect 1830 2656 1831 2660
rect 1835 2656 1836 2660
rect 1830 2655 1836 2656
rect 2022 2660 2028 2661
rect 2022 2656 2023 2660
rect 2027 2656 2028 2660
rect 2022 2655 2028 2656
rect 2230 2660 2236 2661
rect 2230 2656 2231 2660
rect 2235 2656 2236 2660
rect 2230 2655 2236 2656
rect 2430 2660 2436 2661
rect 2430 2656 2431 2660
rect 2435 2656 2436 2660
rect 2430 2655 2436 2656
rect 2614 2660 2620 2661
rect 2614 2656 2615 2660
rect 2619 2656 2620 2660
rect 2614 2655 2620 2656
rect 2782 2660 2788 2661
rect 2782 2656 2783 2660
rect 2787 2656 2788 2660
rect 2782 2655 2788 2656
rect 2942 2660 2948 2661
rect 2942 2656 2943 2660
rect 2947 2656 2948 2660
rect 2942 2655 2948 2656
rect 3094 2660 3100 2661
rect 3094 2656 3095 2660
rect 3099 2656 3100 2660
rect 3094 2655 3100 2656
rect 3238 2660 3244 2661
rect 3238 2656 3239 2660
rect 3243 2656 3244 2660
rect 3238 2655 3244 2656
rect 3366 2660 3372 2661
rect 3366 2656 3367 2660
rect 3371 2656 3372 2660
rect 3462 2659 3463 2663
rect 3467 2659 3468 2663
rect 3462 2658 3468 2659
rect 3366 2655 3372 2656
rect 1883 2643 1889 2644
rect 1883 2639 1884 2643
rect 1888 2642 1889 2643
rect 1910 2643 1916 2644
rect 1910 2642 1911 2643
rect 1888 2640 1911 2642
rect 1888 2639 1889 2640
rect 1883 2638 1889 2639
rect 1910 2639 1911 2640
rect 1915 2639 1916 2643
rect 1910 2638 1916 2639
rect 2075 2643 2081 2644
rect 2075 2639 2076 2643
rect 2080 2642 2081 2643
rect 2102 2643 2108 2644
rect 2102 2642 2103 2643
rect 2080 2640 2103 2642
rect 2080 2639 2081 2640
rect 2075 2638 2081 2639
rect 2102 2639 2103 2640
rect 2107 2639 2108 2643
rect 2102 2638 2108 2639
rect 2254 2643 2260 2644
rect 2254 2639 2255 2643
rect 2259 2642 2260 2643
rect 2283 2643 2289 2644
rect 2283 2642 2284 2643
rect 2259 2640 2284 2642
rect 2259 2639 2260 2640
rect 2254 2638 2260 2639
rect 2283 2639 2284 2640
rect 2288 2639 2289 2643
rect 2283 2638 2289 2639
rect 2483 2643 2489 2644
rect 2483 2639 2484 2643
rect 2488 2642 2489 2643
rect 2542 2643 2548 2644
rect 2542 2642 2543 2643
rect 2488 2640 2543 2642
rect 2488 2639 2489 2640
rect 2483 2638 2489 2639
rect 2542 2639 2543 2640
rect 2547 2639 2548 2643
rect 2542 2638 2548 2639
rect 2590 2643 2596 2644
rect 2590 2639 2591 2643
rect 2595 2642 2596 2643
rect 2667 2643 2673 2644
rect 2667 2642 2668 2643
rect 2595 2640 2668 2642
rect 2595 2639 2596 2640
rect 2590 2638 2596 2639
rect 2667 2639 2668 2640
rect 2672 2639 2673 2643
rect 2667 2638 2673 2639
rect 2686 2643 2692 2644
rect 2686 2639 2687 2643
rect 2691 2642 2692 2643
rect 2835 2643 2841 2644
rect 2835 2642 2836 2643
rect 2691 2640 2836 2642
rect 2691 2639 2692 2640
rect 2686 2638 2692 2639
rect 2835 2639 2836 2640
rect 2840 2639 2841 2643
rect 2835 2638 2841 2639
rect 2854 2643 2860 2644
rect 2854 2639 2855 2643
rect 2859 2642 2860 2643
rect 2995 2643 3001 2644
rect 2995 2642 2996 2643
rect 2859 2640 2996 2642
rect 2859 2639 2860 2640
rect 2854 2638 2860 2639
rect 2995 2639 2996 2640
rect 3000 2639 3001 2643
rect 2995 2638 3001 2639
rect 3014 2643 3020 2644
rect 3014 2639 3015 2643
rect 3019 2642 3020 2643
rect 3147 2643 3153 2644
rect 3147 2642 3148 2643
rect 3019 2640 3148 2642
rect 3019 2639 3020 2640
rect 3014 2638 3020 2639
rect 3147 2639 3148 2640
rect 3152 2639 3153 2643
rect 3147 2638 3153 2639
rect 3291 2643 3297 2644
rect 3291 2639 3292 2643
rect 3296 2642 3297 2643
rect 3318 2643 3324 2644
rect 3318 2642 3319 2643
rect 3296 2640 3319 2642
rect 3296 2639 3297 2640
rect 3291 2638 3297 2639
rect 3318 2639 3319 2640
rect 3323 2639 3324 2643
rect 3318 2638 3324 2639
rect 3419 2643 3425 2644
rect 3419 2639 3420 2643
rect 3424 2642 3425 2643
rect 3430 2643 3436 2644
rect 3430 2642 3431 2643
rect 3424 2640 3431 2642
rect 3424 2639 3425 2640
rect 3419 2638 3425 2639
rect 3430 2639 3431 2640
rect 3435 2639 3436 2643
rect 3430 2638 3436 2639
rect 110 2628 116 2629
rect 1766 2628 1772 2629
rect 110 2624 111 2628
rect 115 2624 116 2628
rect 110 2623 116 2624
rect 470 2627 476 2628
rect 470 2623 471 2627
rect 475 2623 476 2627
rect 470 2622 476 2623
rect 558 2627 564 2628
rect 558 2623 559 2627
rect 563 2623 564 2627
rect 558 2622 564 2623
rect 646 2627 652 2628
rect 646 2623 647 2627
rect 651 2623 652 2627
rect 646 2622 652 2623
rect 734 2627 740 2628
rect 734 2623 735 2627
rect 739 2623 740 2627
rect 734 2622 740 2623
rect 822 2627 828 2628
rect 822 2623 823 2627
rect 827 2623 828 2627
rect 822 2622 828 2623
rect 910 2627 916 2628
rect 910 2623 911 2627
rect 915 2623 916 2627
rect 910 2622 916 2623
rect 998 2627 1004 2628
rect 998 2623 999 2627
rect 1003 2623 1004 2627
rect 998 2622 1004 2623
rect 1086 2627 1092 2628
rect 1086 2623 1087 2627
rect 1091 2623 1092 2627
rect 1766 2624 1767 2628
rect 1771 2624 1772 2628
rect 1766 2623 1772 2624
rect 1798 2627 1804 2628
rect 1798 2623 1799 2627
rect 1803 2626 1804 2627
rect 1883 2627 1889 2628
rect 1883 2626 1884 2627
rect 1803 2624 1884 2626
rect 1803 2623 1804 2624
rect 1086 2622 1092 2623
rect 1798 2622 1804 2623
rect 1883 2623 1884 2624
rect 1888 2623 1889 2627
rect 1883 2622 1889 2623
rect 1902 2627 1908 2628
rect 1902 2623 1903 2627
rect 1907 2626 1908 2627
rect 2051 2627 2057 2628
rect 2051 2626 2052 2627
rect 1907 2624 2052 2626
rect 1907 2623 1908 2624
rect 1902 2622 1908 2623
rect 2051 2623 2052 2624
rect 2056 2623 2057 2627
rect 2051 2622 2057 2623
rect 2070 2627 2076 2628
rect 2070 2623 2071 2627
rect 2075 2626 2076 2627
rect 2235 2627 2241 2628
rect 2235 2626 2236 2627
rect 2075 2624 2236 2626
rect 2075 2623 2076 2624
rect 2070 2622 2076 2623
rect 2235 2623 2236 2624
rect 2240 2623 2241 2627
rect 2235 2622 2241 2623
rect 2411 2627 2420 2628
rect 2411 2623 2412 2627
rect 2419 2623 2420 2627
rect 2411 2622 2420 2623
rect 2571 2627 2577 2628
rect 2571 2623 2572 2627
rect 2576 2626 2577 2627
rect 2599 2627 2605 2628
rect 2599 2626 2600 2627
rect 2576 2624 2600 2626
rect 2576 2623 2577 2624
rect 2571 2622 2577 2623
rect 2599 2623 2600 2624
rect 2604 2623 2605 2627
rect 2599 2622 2605 2623
rect 2723 2627 2729 2628
rect 2723 2623 2724 2627
rect 2728 2626 2729 2627
rect 2751 2627 2757 2628
rect 2751 2626 2752 2627
rect 2728 2624 2752 2626
rect 2728 2623 2729 2624
rect 2723 2622 2729 2623
rect 2751 2623 2752 2624
rect 2756 2623 2757 2627
rect 2751 2622 2757 2623
rect 2859 2627 2865 2628
rect 2859 2623 2860 2627
rect 2864 2626 2865 2627
rect 2914 2627 2920 2628
rect 2914 2626 2915 2627
rect 2864 2624 2915 2626
rect 2864 2623 2865 2624
rect 2859 2622 2865 2623
rect 2914 2623 2915 2624
rect 2919 2623 2920 2627
rect 2914 2622 2920 2623
rect 2979 2627 2985 2628
rect 2979 2623 2980 2627
rect 2984 2626 2985 2627
rect 3034 2627 3040 2628
rect 3034 2626 3035 2627
rect 2984 2624 3035 2626
rect 2984 2623 2985 2624
rect 2979 2622 2985 2623
rect 3034 2623 3035 2624
rect 3039 2623 3040 2627
rect 3034 2622 3040 2623
rect 3099 2627 3105 2628
rect 3099 2623 3100 2627
rect 3104 2626 3105 2627
rect 3150 2627 3156 2628
rect 3150 2626 3151 2627
rect 3104 2624 3151 2626
rect 3104 2623 3105 2624
rect 3099 2622 3105 2623
rect 3150 2623 3151 2624
rect 3155 2623 3156 2627
rect 3150 2622 3156 2623
rect 3211 2627 3217 2628
rect 3211 2623 3212 2627
rect 3216 2626 3217 2627
rect 3239 2627 3245 2628
rect 3239 2626 3240 2627
rect 3216 2624 3240 2626
rect 3216 2623 3217 2624
rect 3211 2622 3217 2623
rect 3239 2623 3240 2624
rect 3244 2623 3245 2627
rect 3239 2622 3245 2623
rect 3310 2627 3316 2628
rect 3310 2623 3311 2627
rect 3315 2626 3316 2627
rect 3323 2627 3329 2628
rect 3323 2626 3324 2627
rect 3315 2624 3324 2626
rect 3315 2623 3316 2624
rect 3310 2622 3316 2623
rect 3323 2623 3324 2624
rect 3328 2623 3329 2627
rect 3419 2627 3425 2628
rect 3419 2626 3420 2627
rect 3323 2622 3329 2623
rect 3332 2624 3420 2626
rect 550 2619 556 2620
rect 542 2615 548 2616
rect 110 2611 116 2612
rect 110 2607 111 2611
rect 115 2607 116 2611
rect 542 2611 543 2615
rect 547 2611 548 2615
rect 550 2615 551 2619
rect 555 2618 556 2619
rect 638 2619 644 2620
rect 555 2616 601 2618
rect 555 2615 556 2616
rect 550 2614 556 2615
rect 638 2615 639 2619
rect 643 2618 644 2619
rect 726 2619 732 2620
rect 643 2616 689 2618
rect 643 2615 644 2616
rect 638 2614 644 2615
rect 726 2615 727 2619
rect 731 2618 732 2619
rect 814 2619 820 2620
rect 731 2616 777 2618
rect 731 2615 732 2616
rect 726 2614 732 2615
rect 814 2615 815 2619
rect 819 2618 820 2619
rect 1078 2619 1084 2620
rect 819 2616 865 2618
rect 819 2615 820 2616
rect 814 2614 820 2615
rect 982 2615 988 2616
rect 542 2610 548 2611
rect 982 2611 983 2615
rect 987 2611 988 2615
rect 982 2610 988 2611
rect 1070 2615 1076 2616
rect 1070 2611 1071 2615
rect 1075 2611 1076 2615
rect 1078 2615 1079 2619
rect 1083 2618 1084 2619
rect 2870 2619 2876 2620
rect 1083 2616 1129 2618
rect 1083 2615 1084 2616
rect 1078 2614 1084 2615
rect 2870 2615 2871 2619
rect 2875 2618 2876 2619
rect 3332 2618 3334 2624
rect 3419 2623 3420 2624
rect 3424 2623 3425 2627
rect 3419 2622 3425 2623
rect 2875 2616 3334 2618
rect 2875 2615 2876 2616
rect 2870 2614 2876 2615
rect 1830 2612 1836 2613
rect 1070 2610 1076 2611
rect 1766 2611 1772 2612
rect 110 2606 116 2607
rect 470 2608 476 2609
rect 470 2604 471 2608
rect 475 2604 476 2608
rect 470 2603 476 2604
rect 558 2608 564 2609
rect 558 2604 559 2608
rect 563 2604 564 2608
rect 558 2603 564 2604
rect 646 2608 652 2609
rect 646 2604 647 2608
rect 651 2604 652 2608
rect 646 2603 652 2604
rect 734 2608 740 2609
rect 734 2604 735 2608
rect 739 2604 740 2608
rect 734 2603 740 2604
rect 822 2608 828 2609
rect 822 2604 823 2608
rect 827 2604 828 2608
rect 822 2603 828 2604
rect 910 2608 916 2609
rect 910 2604 911 2608
rect 915 2604 916 2608
rect 910 2603 916 2604
rect 998 2608 1004 2609
rect 998 2604 999 2608
rect 1003 2604 1004 2608
rect 998 2603 1004 2604
rect 1086 2608 1092 2609
rect 1086 2604 1087 2608
rect 1091 2604 1092 2608
rect 1766 2607 1767 2611
rect 1771 2607 1772 2611
rect 1766 2606 1772 2607
rect 1806 2609 1812 2610
rect 1806 2605 1807 2609
rect 1811 2605 1812 2609
rect 1830 2608 1831 2612
rect 1835 2608 1836 2612
rect 1830 2607 1836 2608
rect 1998 2612 2004 2613
rect 1998 2608 1999 2612
rect 2003 2608 2004 2612
rect 1998 2607 2004 2608
rect 2182 2612 2188 2613
rect 2182 2608 2183 2612
rect 2187 2608 2188 2612
rect 2182 2607 2188 2608
rect 2358 2612 2364 2613
rect 2358 2608 2359 2612
rect 2363 2608 2364 2612
rect 2358 2607 2364 2608
rect 2518 2612 2524 2613
rect 2518 2608 2519 2612
rect 2523 2608 2524 2612
rect 2518 2607 2524 2608
rect 2670 2612 2676 2613
rect 2670 2608 2671 2612
rect 2675 2608 2676 2612
rect 2670 2607 2676 2608
rect 2806 2612 2812 2613
rect 2806 2608 2807 2612
rect 2811 2608 2812 2612
rect 2806 2607 2812 2608
rect 2926 2612 2932 2613
rect 2926 2608 2927 2612
rect 2931 2608 2932 2612
rect 2926 2607 2932 2608
rect 3046 2612 3052 2613
rect 3046 2608 3047 2612
rect 3051 2608 3052 2612
rect 3046 2607 3052 2608
rect 3158 2612 3164 2613
rect 3158 2608 3159 2612
rect 3163 2608 3164 2612
rect 3158 2607 3164 2608
rect 3270 2612 3276 2613
rect 3270 2608 3271 2612
rect 3275 2608 3276 2612
rect 3270 2607 3276 2608
rect 3366 2612 3372 2613
rect 3366 2608 3367 2612
rect 3371 2608 3372 2612
rect 3366 2607 3372 2608
rect 3462 2609 3468 2610
rect 1806 2604 1812 2605
rect 3462 2605 3463 2609
rect 3467 2605 3468 2609
rect 3462 2604 3468 2605
rect 1086 2603 1092 2604
rect 1902 2603 1908 2604
rect 1902 2599 1903 2603
rect 1907 2599 1908 2603
rect 1902 2598 1908 2599
rect 2070 2603 2076 2604
rect 2070 2599 2071 2603
rect 2075 2599 2076 2603
rect 2070 2598 2076 2599
rect 2254 2603 2260 2604
rect 2254 2599 2255 2603
rect 2259 2599 2260 2603
rect 2254 2598 2260 2599
rect 2262 2603 2268 2604
rect 2262 2599 2263 2603
rect 2267 2602 2268 2603
rect 2590 2603 2596 2604
rect 2267 2600 2401 2602
rect 2267 2599 2268 2600
rect 2262 2598 2268 2599
rect 2590 2599 2591 2603
rect 2595 2599 2596 2603
rect 2590 2598 2596 2599
rect 2599 2603 2605 2604
rect 2599 2599 2600 2603
rect 2604 2602 2605 2603
rect 2751 2603 2757 2604
rect 2604 2600 2713 2602
rect 2604 2599 2605 2600
rect 2599 2598 2605 2599
rect 2751 2599 2752 2603
rect 2756 2602 2757 2603
rect 2914 2603 2920 2604
rect 2756 2600 2849 2602
rect 2756 2599 2757 2600
rect 2751 2598 2757 2599
rect 2914 2599 2915 2603
rect 2919 2602 2920 2603
rect 3034 2603 3040 2604
rect 2919 2600 2969 2602
rect 2919 2599 2920 2600
rect 2914 2598 2920 2599
rect 3034 2599 3035 2603
rect 3039 2602 3040 2603
rect 3150 2603 3156 2604
rect 3039 2600 3089 2602
rect 3039 2599 3040 2600
rect 3034 2598 3040 2599
rect 3150 2599 3151 2603
rect 3155 2602 3156 2603
rect 3239 2603 3245 2604
rect 3155 2600 3201 2602
rect 3155 2599 3156 2600
rect 3150 2598 3156 2599
rect 3239 2599 3240 2603
rect 3244 2602 3245 2603
rect 3430 2603 3436 2604
rect 3244 2600 3313 2602
rect 3244 2599 3245 2600
rect 3239 2598 3245 2599
rect 3430 2599 3431 2603
rect 3435 2599 3436 2603
rect 3430 2598 3436 2599
rect 1830 2593 1836 2594
rect 1806 2592 1812 2593
rect 523 2591 529 2592
rect 523 2587 524 2591
rect 528 2590 529 2591
rect 550 2591 556 2592
rect 550 2590 551 2591
rect 528 2588 551 2590
rect 528 2587 529 2588
rect 523 2586 529 2587
rect 550 2587 551 2588
rect 555 2587 556 2591
rect 550 2586 556 2587
rect 611 2591 617 2592
rect 611 2587 612 2591
rect 616 2590 617 2591
rect 638 2591 644 2592
rect 638 2590 639 2591
rect 616 2588 639 2590
rect 616 2587 617 2588
rect 611 2586 617 2587
rect 638 2587 639 2588
rect 643 2587 644 2591
rect 638 2586 644 2587
rect 699 2591 705 2592
rect 699 2587 700 2591
rect 704 2590 705 2591
rect 726 2591 732 2592
rect 726 2590 727 2591
rect 704 2588 727 2590
rect 704 2587 705 2588
rect 699 2586 705 2587
rect 726 2587 727 2588
rect 731 2587 732 2591
rect 726 2586 732 2587
rect 787 2591 793 2592
rect 787 2587 788 2591
rect 792 2590 793 2591
rect 814 2591 820 2592
rect 814 2590 815 2591
rect 792 2588 815 2590
rect 792 2587 793 2588
rect 787 2586 793 2587
rect 814 2587 815 2588
rect 819 2587 820 2591
rect 814 2586 820 2587
rect 875 2591 881 2592
rect 875 2587 876 2591
rect 880 2590 881 2591
rect 902 2591 908 2592
rect 902 2590 903 2591
rect 880 2588 903 2590
rect 880 2587 881 2588
rect 875 2586 881 2587
rect 902 2587 903 2588
rect 907 2587 908 2591
rect 963 2591 969 2592
rect 963 2590 964 2591
rect 902 2586 908 2587
rect 912 2588 964 2590
rect 838 2583 844 2584
rect 838 2579 839 2583
rect 843 2582 844 2583
rect 912 2582 914 2588
rect 963 2587 964 2588
rect 968 2587 969 2591
rect 963 2586 969 2587
rect 982 2591 988 2592
rect 982 2587 983 2591
rect 987 2590 988 2591
rect 1051 2591 1057 2592
rect 1051 2590 1052 2591
rect 987 2588 1052 2590
rect 987 2587 988 2588
rect 982 2586 988 2587
rect 1051 2587 1052 2588
rect 1056 2587 1057 2591
rect 1051 2586 1057 2587
rect 1070 2591 1076 2592
rect 1070 2587 1071 2591
rect 1075 2590 1076 2591
rect 1139 2591 1145 2592
rect 1139 2590 1140 2591
rect 1075 2588 1140 2590
rect 1075 2587 1076 2588
rect 1070 2586 1076 2587
rect 1139 2587 1140 2588
rect 1144 2587 1145 2591
rect 1806 2588 1807 2592
rect 1811 2588 1812 2592
rect 1830 2589 1831 2593
rect 1835 2589 1836 2593
rect 1830 2588 1836 2589
rect 1998 2593 2004 2594
rect 1998 2589 1999 2593
rect 2003 2589 2004 2593
rect 1998 2588 2004 2589
rect 2182 2593 2188 2594
rect 2182 2589 2183 2593
rect 2187 2589 2188 2593
rect 2182 2588 2188 2589
rect 2358 2593 2364 2594
rect 2358 2589 2359 2593
rect 2363 2589 2364 2593
rect 2358 2588 2364 2589
rect 2518 2593 2524 2594
rect 2518 2589 2519 2593
rect 2523 2589 2524 2593
rect 2518 2588 2524 2589
rect 2670 2593 2676 2594
rect 2670 2589 2671 2593
rect 2675 2589 2676 2593
rect 2670 2588 2676 2589
rect 2806 2593 2812 2594
rect 2806 2589 2807 2593
rect 2811 2589 2812 2593
rect 2806 2588 2812 2589
rect 2926 2593 2932 2594
rect 2926 2589 2927 2593
rect 2931 2589 2932 2593
rect 2926 2588 2932 2589
rect 3046 2593 3052 2594
rect 3046 2589 3047 2593
rect 3051 2589 3052 2593
rect 3046 2588 3052 2589
rect 3158 2593 3164 2594
rect 3158 2589 3159 2593
rect 3163 2589 3164 2593
rect 3158 2588 3164 2589
rect 3270 2593 3276 2594
rect 3270 2589 3271 2593
rect 3275 2589 3276 2593
rect 3270 2588 3276 2589
rect 3366 2593 3372 2594
rect 3366 2589 3367 2593
rect 3371 2589 3372 2593
rect 3366 2588 3372 2589
rect 3462 2592 3468 2593
rect 3462 2588 3463 2592
rect 3467 2588 3468 2592
rect 1806 2587 1812 2588
rect 3462 2587 3468 2588
rect 1139 2586 1145 2587
rect 843 2580 914 2582
rect 843 2579 844 2580
rect 838 2578 844 2579
rect 275 2567 281 2568
rect 275 2563 276 2567
rect 280 2566 281 2567
rect 294 2567 300 2568
rect 280 2564 290 2566
rect 280 2563 281 2564
rect 275 2562 281 2563
rect 288 2558 290 2564
rect 294 2563 295 2567
rect 299 2566 300 2567
rect 363 2567 369 2568
rect 363 2566 364 2567
rect 299 2564 364 2566
rect 299 2563 300 2564
rect 294 2562 300 2563
rect 363 2563 364 2564
rect 368 2563 369 2567
rect 363 2562 369 2563
rect 459 2567 465 2568
rect 459 2563 460 2567
rect 464 2566 465 2567
rect 542 2567 548 2568
rect 464 2564 538 2566
rect 464 2563 465 2564
rect 459 2562 465 2563
rect 536 2558 538 2564
rect 542 2563 543 2567
rect 547 2566 548 2567
rect 555 2567 561 2568
rect 555 2566 556 2567
rect 547 2564 556 2566
rect 547 2563 548 2564
rect 542 2562 548 2563
rect 555 2563 556 2564
rect 560 2563 561 2567
rect 555 2562 561 2563
rect 574 2567 580 2568
rect 574 2563 575 2567
rect 579 2566 580 2567
rect 643 2567 649 2568
rect 643 2566 644 2567
rect 579 2564 644 2566
rect 579 2563 580 2564
rect 574 2562 580 2563
rect 643 2563 644 2564
rect 648 2563 649 2567
rect 643 2562 649 2563
rect 731 2567 737 2568
rect 731 2563 732 2567
rect 736 2566 737 2567
rect 750 2567 756 2568
rect 736 2564 746 2566
rect 736 2563 737 2564
rect 731 2562 737 2563
rect 744 2558 746 2564
rect 750 2563 751 2567
rect 755 2566 756 2567
rect 819 2567 825 2568
rect 819 2566 820 2567
rect 755 2564 820 2566
rect 755 2563 756 2564
rect 750 2562 756 2563
rect 819 2563 820 2564
rect 824 2563 825 2567
rect 819 2562 825 2563
rect 907 2567 913 2568
rect 907 2563 908 2567
rect 912 2566 913 2567
rect 926 2567 932 2568
rect 912 2564 922 2566
rect 912 2563 913 2564
rect 907 2562 913 2563
rect 806 2559 812 2560
rect 806 2558 807 2559
rect 288 2556 394 2558
rect 536 2556 586 2558
rect 744 2556 807 2558
rect 222 2552 228 2553
rect 110 2549 116 2550
rect 110 2545 111 2549
rect 115 2545 116 2549
rect 222 2548 223 2552
rect 227 2548 228 2552
rect 222 2547 228 2548
rect 310 2552 316 2553
rect 310 2548 311 2552
rect 315 2548 316 2552
rect 310 2547 316 2548
rect 110 2544 116 2545
rect 294 2543 300 2544
rect 294 2539 295 2543
rect 299 2539 300 2543
rect 294 2538 300 2539
rect 382 2543 388 2544
rect 382 2539 383 2543
rect 387 2539 388 2543
rect 392 2542 394 2556
rect 406 2552 412 2553
rect 406 2548 407 2552
rect 411 2548 412 2552
rect 406 2547 412 2548
rect 502 2552 508 2553
rect 502 2548 503 2552
rect 507 2548 508 2552
rect 502 2547 508 2548
rect 574 2543 580 2544
rect 392 2540 449 2542
rect 382 2538 388 2539
rect 574 2539 575 2543
rect 579 2539 580 2543
rect 584 2542 586 2556
rect 806 2555 807 2556
rect 811 2555 812 2559
rect 920 2558 922 2564
rect 926 2563 927 2567
rect 931 2566 932 2567
rect 995 2567 1001 2568
rect 995 2566 996 2567
rect 931 2564 996 2566
rect 931 2563 932 2564
rect 926 2562 932 2563
rect 995 2563 996 2564
rect 1000 2563 1001 2567
rect 995 2562 1001 2563
rect 1014 2567 1020 2568
rect 1014 2563 1015 2567
rect 1019 2566 1020 2567
rect 1083 2567 1089 2568
rect 1083 2566 1084 2567
rect 1019 2564 1084 2566
rect 1019 2563 1020 2564
rect 1014 2562 1020 2563
rect 1083 2563 1084 2564
rect 1088 2563 1089 2567
rect 1083 2562 1089 2563
rect 1102 2567 1108 2568
rect 1102 2563 1103 2567
rect 1107 2566 1108 2567
rect 1171 2567 1177 2568
rect 1171 2566 1172 2567
rect 1107 2564 1172 2566
rect 1107 2563 1108 2564
rect 1102 2562 1108 2563
rect 1171 2563 1172 2564
rect 1176 2563 1177 2567
rect 1171 2562 1177 2563
rect 1190 2567 1196 2568
rect 1190 2563 1191 2567
rect 1195 2566 1196 2567
rect 1267 2567 1273 2568
rect 1267 2566 1268 2567
rect 1195 2564 1268 2566
rect 1195 2563 1196 2564
rect 1190 2562 1196 2563
rect 1267 2563 1268 2564
rect 1272 2563 1273 2567
rect 1267 2562 1273 2563
rect 1286 2567 1292 2568
rect 1286 2563 1287 2567
rect 1291 2566 1292 2567
rect 1363 2567 1369 2568
rect 1363 2566 1364 2567
rect 1291 2564 1364 2566
rect 1291 2563 1292 2564
rect 1286 2562 1292 2563
rect 1363 2563 1364 2564
rect 1368 2563 1369 2567
rect 1363 2562 1369 2563
rect 1459 2567 1465 2568
rect 1459 2563 1460 2567
rect 1464 2566 1465 2567
rect 1495 2567 1501 2568
rect 1464 2564 1490 2566
rect 1464 2563 1465 2564
rect 1459 2562 1465 2563
rect 1054 2559 1060 2560
rect 1054 2558 1055 2559
rect 920 2556 1055 2558
rect 806 2554 812 2555
rect 1054 2555 1055 2556
rect 1059 2555 1060 2559
rect 1488 2558 1490 2564
rect 1495 2563 1496 2567
rect 1500 2566 1501 2567
rect 1547 2567 1553 2568
rect 1547 2566 1548 2567
rect 1500 2564 1548 2566
rect 1500 2563 1501 2564
rect 1495 2562 1501 2563
rect 1547 2563 1548 2564
rect 1552 2563 1553 2567
rect 1547 2562 1553 2563
rect 1566 2567 1572 2568
rect 1566 2563 1567 2567
rect 1571 2566 1572 2567
rect 1635 2567 1641 2568
rect 1635 2566 1636 2567
rect 1571 2564 1636 2566
rect 1571 2563 1572 2564
rect 1566 2562 1572 2563
rect 1635 2563 1636 2564
rect 1640 2563 1641 2567
rect 1635 2562 1641 2563
rect 1654 2567 1660 2568
rect 1654 2563 1655 2567
rect 1659 2566 1660 2567
rect 1723 2567 1729 2568
rect 1723 2566 1724 2567
rect 1659 2564 1724 2566
rect 1659 2563 1660 2564
rect 1654 2562 1660 2563
rect 1723 2563 1724 2564
rect 1728 2563 1729 2567
rect 1723 2562 1729 2563
rect 1662 2559 1668 2560
rect 1662 2558 1663 2559
rect 1488 2556 1663 2558
rect 1054 2554 1060 2555
rect 1662 2555 1663 2556
rect 1667 2555 1668 2559
rect 1662 2554 1668 2555
rect 590 2552 596 2553
rect 590 2548 591 2552
rect 595 2548 596 2552
rect 590 2547 596 2548
rect 678 2552 684 2553
rect 678 2548 679 2552
rect 683 2548 684 2552
rect 678 2547 684 2548
rect 766 2552 772 2553
rect 766 2548 767 2552
rect 771 2548 772 2552
rect 766 2547 772 2548
rect 854 2552 860 2553
rect 854 2548 855 2552
rect 859 2548 860 2552
rect 854 2547 860 2548
rect 942 2552 948 2553
rect 942 2548 943 2552
rect 947 2548 948 2552
rect 942 2547 948 2548
rect 1030 2552 1036 2553
rect 1030 2548 1031 2552
rect 1035 2548 1036 2552
rect 1030 2547 1036 2548
rect 1118 2552 1124 2553
rect 1118 2548 1119 2552
rect 1123 2548 1124 2552
rect 1118 2547 1124 2548
rect 1214 2552 1220 2553
rect 1214 2548 1215 2552
rect 1219 2548 1220 2552
rect 1214 2547 1220 2548
rect 1310 2552 1316 2553
rect 1310 2548 1311 2552
rect 1315 2548 1316 2552
rect 1310 2547 1316 2548
rect 1406 2552 1412 2553
rect 1406 2548 1407 2552
rect 1411 2548 1412 2552
rect 1406 2547 1412 2548
rect 1494 2552 1500 2553
rect 1494 2548 1495 2552
rect 1499 2548 1500 2552
rect 1494 2547 1500 2548
rect 1582 2552 1588 2553
rect 1582 2548 1583 2552
rect 1587 2548 1588 2552
rect 1582 2547 1588 2548
rect 1670 2552 1676 2553
rect 1670 2548 1671 2552
rect 1675 2548 1676 2552
rect 1670 2547 1676 2548
rect 1766 2549 1772 2550
rect 1766 2545 1767 2549
rect 1771 2545 1772 2549
rect 1766 2544 1772 2545
rect 750 2543 756 2544
rect 584 2540 633 2542
rect 574 2538 580 2539
rect 750 2539 751 2543
rect 755 2539 756 2543
rect 750 2538 756 2539
rect 838 2543 844 2544
rect 838 2539 839 2543
rect 843 2539 844 2543
rect 838 2538 844 2539
rect 926 2543 932 2544
rect 926 2539 927 2543
rect 931 2539 932 2543
rect 926 2538 932 2539
rect 1014 2543 1020 2544
rect 1014 2539 1015 2543
rect 1019 2539 1020 2543
rect 1014 2538 1020 2539
rect 1102 2543 1108 2544
rect 1102 2539 1103 2543
rect 1107 2539 1108 2543
rect 1102 2538 1108 2539
rect 1190 2543 1196 2544
rect 1190 2539 1191 2543
rect 1195 2539 1196 2543
rect 1190 2538 1196 2539
rect 1286 2543 1292 2544
rect 1286 2539 1287 2543
rect 1291 2539 1292 2543
rect 1286 2538 1292 2539
rect 1382 2543 1388 2544
rect 1382 2539 1383 2543
rect 1387 2539 1388 2543
rect 1487 2543 1493 2544
rect 1487 2542 1488 2543
rect 1481 2540 1488 2542
rect 1382 2538 1388 2539
rect 1487 2539 1488 2540
rect 1492 2539 1493 2543
rect 1487 2538 1493 2539
rect 1566 2543 1572 2544
rect 1566 2539 1567 2543
rect 1571 2539 1572 2543
rect 1566 2538 1572 2539
rect 1654 2543 1660 2544
rect 1654 2539 1655 2543
rect 1659 2539 1660 2543
rect 1798 2543 1804 2544
rect 1798 2542 1799 2543
rect 1745 2540 1799 2542
rect 1654 2538 1660 2539
rect 1798 2539 1799 2540
rect 1803 2539 1804 2543
rect 1798 2538 1804 2539
rect 1806 2540 1812 2541
rect 3462 2540 3468 2541
rect 1806 2536 1807 2540
rect 1811 2536 1812 2540
rect 1806 2535 1812 2536
rect 2206 2539 2212 2540
rect 2206 2535 2207 2539
rect 2211 2535 2212 2539
rect 2206 2534 2212 2535
rect 2798 2539 2804 2540
rect 2798 2535 2799 2539
rect 2803 2535 2804 2539
rect 2798 2534 2804 2535
rect 3366 2539 3372 2540
rect 3366 2535 3367 2539
rect 3371 2535 3372 2539
rect 3462 2536 3463 2540
rect 3467 2536 3468 2540
rect 3462 2535 3468 2536
rect 3366 2534 3372 2535
rect 222 2533 228 2534
rect 110 2532 116 2533
rect 110 2528 111 2532
rect 115 2528 116 2532
rect 222 2529 223 2533
rect 227 2529 228 2533
rect 222 2528 228 2529
rect 310 2533 316 2534
rect 310 2529 311 2533
rect 315 2529 316 2533
rect 310 2528 316 2529
rect 406 2533 412 2534
rect 406 2529 407 2533
rect 411 2529 412 2533
rect 406 2528 412 2529
rect 502 2533 508 2534
rect 502 2529 503 2533
rect 507 2529 508 2533
rect 502 2528 508 2529
rect 590 2533 596 2534
rect 590 2529 591 2533
rect 595 2529 596 2533
rect 590 2528 596 2529
rect 678 2533 684 2534
rect 678 2529 679 2533
rect 683 2529 684 2533
rect 678 2528 684 2529
rect 766 2533 772 2534
rect 766 2529 767 2533
rect 771 2529 772 2533
rect 766 2528 772 2529
rect 854 2533 860 2534
rect 854 2529 855 2533
rect 859 2529 860 2533
rect 854 2528 860 2529
rect 942 2533 948 2534
rect 942 2529 943 2533
rect 947 2529 948 2533
rect 942 2528 948 2529
rect 1030 2533 1036 2534
rect 1030 2529 1031 2533
rect 1035 2529 1036 2533
rect 1030 2528 1036 2529
rect 1118 2533 1124 2534
rect 1118 2529 1119 2533
rect 1123 2529 1124 2533
rect 1118 2528 1124 2529
rect 1214 2533 1220 2534
rect 1214 2529 1215 2533
rect 1219 2529 1220 2533
rect 1214 2528 1220 2529
rect 1310 2533 1316 2534
rect 1310 2529 1311 2533
rect 1315 2529 1316 2533
rect 1310 2528 1316 2529
rect 1406 2533 1412 2534
rect 1406 2529 1407 2533
rect 1411 2529 1412 2533
rect 1406 2528 1412 2529
rect 1494 2533 1500 2534
rect 1494 2529 1495 2533
rect 1499 2529 1500 2533
rect 1494 2528 1500 2529
rect 1582 2533 1588 2534
rect 1582 2529 1583 2533
rect 1587 2529 1588 2533
rect 1582 2528 1588 2529
rect 1670 2533 1676 2534
rect 1670 2529 1671 2533
rect 1675 2529 1676 2533
rect 1670 2528 1676 2529
rect 1766 2532 1772 2533
rect 1766 2528 1767 2532
rect 1771 2528 1772 2532
rect 110 2527 116 2528
rect 1766 2527 1772 2528
rect 2070 2531 2076 2532
rect 2070 2527 2071 2531
rect 2075 2530 2076 2531
rect 2870 2531 2876 2532
rect 2075 2528 2249 2530
rect 2075 2527 2076 2528
rect 2070 2526 2076 2527
rect 2870 2527 2871 2531
rect 2875 2527 2876 2531
rect 2870 2526 2876 2527
rect 2878 2531 2884 2532
rect 2878 2527 2879 2531
rect 2883 2530 2884 2531
rect 2883 2528 3409 2530
rect 2883 2527 2884 2528
rect 2878 2526 2884 2527
rect 1806 2523 1812 2524
rect 1806 2519 1807 2523
rect 1811 2519 1812 2523
rect 3462 2523 3468 2524
rect 1806 2518 1812 2519
rect 2206 2520 2212 2521
rect 2206 2516 2207 2520
rect 2211 2516 2212 2520
rect 2206 2515 2212 2516
rect 2798 2520 2804 2521
rect 2798 2516 2799 2520
rect 2803 2516 2804 2520
rect 2798 2515 2804 2516
rect 3366 2520 3372 2521
rect 3366 2516 3367 2520
rect 3371 2516 3372 2520
rect 3462 2519 3463 2523
rect 3467 2519 3468 2523
rect 3462 2518 3468 2519
rect 3366 2515 3372 2516
rect 2259 2503 2268 2504
rect 2259 2499 2260 2503
rect 2267 2499 2268 2503
rect 2259 2498 2268 2499
rect 2851 2503 2857 2504
rect 2851 2499 2852 2503
rect 2856 2502 2857 2503
rect 2878 2503 2884 2504
rect 2878 2502 2879 2503
rect 2856 2500 2879 2502
rect 2856 2499 2857 2500
rect 2851 2498 2857 2499
rect 2878 2499 2879 2500
rect 2883 2499 2884 2503
rect 2878 2498 2884 2499
rect 3419 2503 3425 2504
rect 3419 2499 3420 2503
rect 3424 2502 3425 2503
rect 3430 2503 3436 2504
rect 3430 2502 3431 2503
rect 3424 2500 3431 2502
rect 3424 2499 3425 2500
rect 3419 2498 3425 2499
rect 3430 2499 3431 2500
rect 3435 2499 3436 2503
rect 3430 2498 3436 2499
rect 110 2488 116 2489
rect 1766 2488 1772 2489
rect 110 2484 111 2488
rect 115 2484 116 2488
rect 110 2483 116 2484
rect 134 2487 140 2488
rect 134 2483 135 2487
rect 139 2483 140 2487
rect 134 2482 140 2483
rect 246 2487 252 2488
rect 246 2483 247 2487
rect 251 2483 252 2487
rect 246 2482 252 2483
rect 390 2487 396 2488
rect 390 2483 391 2487
rect 395 2483 396 2487
rect 390 2482 396 2483
rect 542 2487 548 2488
rect 542 2483 543 2487
rect 547 2483 548 2487
rect 542 2482 548 2483
rect 694 2487 700 2488
rect 694 2483 695 2487
rect 699 2483 700 2487
rect 694 2482 700 2483
rect 838 2487 844 2488
rect 838 2483 839 2487
rect 843 2483 844 2487
rect 838 2482 844 2483
rect 974 2487 980 2488
rect 974 2483 975 2487
rect 979 2483 980 2487
rect 974 2482 980 2483
rect 1102 2487 1108 2488
rect 1102 2483 1103 2487
rect 1107 2483 1108 2487
rect 1102 2482 1108 2483
rect 1230 2487 1236 2488
rect 1230 2483 1231 2487
rect 1235 2483 1236 2487
rect 1230 2482 1236 2483
rect 1350 2487 1356 2488
rect 1350 2483 1351 2487
rect 1355 2483 1356 2487
rect 1350 2482 1356 2483
rect 1462 2487 1468 2488
rect 1462 2483 1463 2487
rect 1467 2483 1468 2487
rect 1462 2482 1468 2483
rect 1574 2487 1580 2488
rect 1574 2483 1575 2487
rect 1579 2483 1580 2487
rect 1574 2482 1580 2483
rect 1670 2487 1676 2488
rect 1670 2483 1671 2487
rect 1675 2483 1676 2487
rect 1766 2484 1767 2488
rect 1771 2484 1772 2488
rect 1766 2483 1772 2484
rect 1670 2482 1676 2483
rect 214 2479 220 2480
rect 206 2475 212 2476
rect 110 2471 116 2472
rect 110 2467 111 2471
rect 115 2467 116 2471
rect 206 2471 207 2475
rect 211 2471 212 2475
rect 214 2475 215 2479
rect 219 2478 220 2479
rect 622 2479 628 2480
rect 219 2476 289 2478
rect 219 2475 220 2476
rect 214 2474 220 2475
rect 462 2475 468 2476
rect 206 2470 212 2471
rect 462 2471 463 2475
rect 467 2471 468 2475
rect 462 2470 468 2471
rect 614 2475 620 2476
rect 614 2471 615 2475
rect 619 2471 620 2475
rect 622 2475 623 2479
rect 627 2478 628 2479
rect 806 2479 812 2480
rect 627 2476 737 2478
rect 627 2475 628 2476
rect 622 2474 628 2475
rect 806 2475 807 2479
rect 811 2478 812 2479
rect 918 2479 924 2480
rect 811 2476 881 2478
rect 811 2475 812 2476
rect 806 2474 812 2475
rect 918 2475 919 2479
rect 923 2478 924 2479
rect 1054 2479 1060 2480
rect 923 2476 1017 2478
rect 923 2475 924 2476
rect 918 2474 924 2475
rect 1054 2475 1055 2479
rect 1059 2478 1060 2479
rect 1182 2479 1188 2480
rect 1059 2476 1145 2478
rect 1059 2475 1060 2476
rect 1054 2474 1060 2475
rect 1182 2475 1183 2479
rect 1187 2478 1188 2479
rect 1310 2479 1316 2480
rect 1187 2476 1273 2478
rect 1187 2475 1188 2476
rect 1182 2474 1188 2475
rect 1310 2475 1311 2479
rect 1315 2478 1316 2479
rect 1662 2479 1668 2480
rect 1315 2476 1393 2478
rect 1315 2475 1316 2476
rect 1310 2474 1316 2475
rect 1534 2475 1540 2476
rect 614 2470 620 2471
rect 1534 2471 1535 2475
rect 1539 2471 1540 2475
rect 1534 2470 1540 2471
rect 1646 2475 1652 2476
rect 1646 2471 1647 2475
rect 1651 2471 1652 2475
rect 1662 2475 1663 2479
rect 1667 2478 1668 2479
rect 1667 2476 1713 2478
rect 1667 2475 1668 2476
rect 1662 2474 1668 2475
rect 2067 2475 2076 2476
rect 1646 2470 1652 2471
rect 1766 2471 1772 2472
rect 110 2466 116 2467
rect 134 2468 140 2469
rect 134 2464 135 2468
rect 139 2464 140 2468
rect 134 2463 140 2464
rect 246 2468 252 2469
rect 246 2464 247 2468
rect 251 2464 252 2468
rect 246 2463 252 2464
rect 390 2468 396 2469
rect 390 2464 391 2468
rect 395 2464 396 2468
rect 390 2463 396 2464
rect 542 2468 548 2469
rect 542 2464 543 2468
rect 547 2464 548 2468
rect 542 2463 548 2464
rect 694 2468 700 2469
rect 694 2464 695 2468
rect 699 2464 700 2468
rect 694 2463 700 2464
rect 838 2468 844 2469
rect 838 2464 839 2468
rect 843 2464 844 2468
rect 838 2463 844 2464
rect 974 2468 980 2469
rect 974 2464 975 2468
rect 979 2464 980 2468
rect 974 2463 980 2464
rect 1102 2468 1108 2469
rect 1102 2464 1103 2468
rect 1107 2464 1108 2468
rect 1102 2463 1108 2464
rect 1230 2468 1236 2469
rect 1230 2464 1231 2468
rect 1235 2464 1236 2468
rect 1230 2463 1236 2464
rect 1350 2468 1356 2469
rect 1350 2464 1351 2468
rect 1355 2464 1356 2468
rect 1350 2463 1356 2464
rect 1462 2468 1468 2469
rect 1462 2464 1463 2468
rect 1467 2464 1468 2468
rect 1462 2463 1468 2464
rect 1574 2468 1580 2469
rect 1574 2464 1575 2468
rect 1579 2464 1580 2468
rect 1574 2463 1580 2464
rect 1670 2468 1676 2469
rect 1670 2464 1671 2468
rect 1675 2464 1676 2468
rect 1766 2467 1767 2471
rect 1771 2467 1772 2471
rect 2067 2471 2068 2475
rect 2075 2471 2076 2475
rect 2067 2470 2076 2471
rect 2086 2475 2092 2476
rect 2086 2471 2087 2475
rect 2091 2474 2092 2475
rect 2251 2475 2257 2476
rect 2251 2474 2252 2475
rect 2091 2472 2252 2474
rect 2091 2471 2092 2472
rect 2086 2470 2092 2471
rect 2251 2471 2252 2472
rect 2256 2471 2257 2475
rect 2251 2470 2257 2471
rect 2270 2475 2276 2476
rect 2270 2471 2271 2475
rect 2275 2474 2276 2475
rect 2419 2475 2425 2476
rect 2419 2474 2420 2475
rect 2275 2472 2420 2474
rect 2275 2471 2276 2472
rect 2270 2470 2276 2471
rect 2419 2471 2420 2472
rect 2424 2471 2425 2475
rect 2419 2470 2425 2471
rect 2579 2475 2585 2476
rect 2579 2471 2580 2475
rect 2584 2474 2585 2475
rect 2630 2475 2636 2476
rect 2630 2474 2631 2475
rect 2584 2472 2631 2474
rect 2584 2471 2585 2472
rect 2579 2470 2585 2471
rect 2630 2471 2631 2472
rect 2635 2471 2636 2475
rect 2630 2470 2636 2471
rect 2646 2475 2652 2476
rect 2646 2471 2647 2475
rect 2651 2474 2652 2475
rect 2723 2475 2729 2476
rect 2723 2474 2724 2475
rect 2651 2472 2724 2474
rect 2651 2471 2652 2472
rect 2646 2470 2652 2471
rect 2723 2471 2724 2472
rect 2728 2471 2729 2475
rect 2723 2470 2729 2471
rect 2742 2475 2748 2476
rect 2742 2471 2743 2475
rect 2747 2474 2748 2475
rect 2859 2475 2865 2476
rect 2859 2474 2860 2475
rect 2747 2472 2860 2474
rect 2747 2471 2748 2472
rect 2742 2470 2748 2471
rect 2859 2471 2860 2472
rect 2864 2471 2865 2475
rect 2859 2470 2865 2471
rect 2878 2475 2884 2476
rect 2878 2471 2879 2475
rect 2883 2474 2884 2475
rect 2979 2475 2985 2476
rect 2979 2474 2980 2475
rect 2883 2472 2980 2474
rect 2883 2471 2884 2472
rect 2878 2470 2884 2471
rect 2979 2471 2980 2472
rect 2984 2471 2985 2475
rect 2979 2470 2985 2471
rect 2998 2475 3004 2476
rect 2998 2471 2999 2475
rect 3003 2474 3004 2475
rect 3099 2475 3105 2476
rect 3099 2474 3100 2475
rect 3003 2472 3100 2474
rect 3003 2471 3004 2472
rect 2998 2470 3004 2471
rect 3099 2471 3100 2472
rect 3104 2471 3105 2475
rect 3099 2470 3105 2471
rect 3118 2475 3124 2476
rect 3118 2471 3119 2475
rect 3123 2474 3124 2475
rect 3211 2475 3217 2476
rect 3211 2474 3212 2475
rect 3123 2472 3212 2474
rect 3123 2471 3124 2472
rect 3118 2470 3124 2471
rect 3211 2471 3212 2472
rect 3216 2471 3217 2475
rect 3211 2470 3217 2471
rect 3230 2475 3236 2476
rect 3230 2471 3231 2475
rect 3235 2474 3236 2475
rect 3323 2475 3329 2476
rect 3323 2474 3324 2475
rect 3235 2472 3324 2474
rect 3235 2471 3236 2472
rect 3230 2470 3236 2471
rect 3323 2471 3324 2472
rect 3328 2471 3329 2475
rect 3323 2470 3329 2471
rect 3419 2475 3425 2476
rect 3419 2471 3420 2475
rect 3424 2474 3425 2475
rect 3438 2475 3444 2476
rect 3438 2474 3439 2475
rect 3424 2472 3439 2474
rect 3424 2471 3425 2472
rect 3419 2470 3425 2471
rect 3438 2471 3439 2472
rect 3443 2471 3444 2475
rect 3438 2470 3444 2471
rect 1766 2466 1772 2467
rect 1670 2463 1676 2464
rect 2014 2460 2020 2461
rect 622 2459 628 2460
rect 622 2458 623 2459
rect 300 2456 623 2458
rect 300 2454 302 2456
rect 622 2455 623 2456
rect 627 2455 628 2459
rect 622 2454 628 2455
rect 1382 2459 1388 2460
rect 1382 2455 1383 2459
rect 1387 2458 1388 2459
rect 1387 2456 1518 2458
rect 1387 2455 1388 2456
rect 1382 2454 1388 2455
rect 1516 2454 1518 2456
rect 1806 2457 1812 2458
rect 299 2453 305 2454
rect 187 2451 193 2452
rect 187 2447 188 2451
rect 192 2450 193 2451
rect 214 2451 220 2452
rect 214 2450 215 2451
rect 192 2448 215 2450
rect 192 2447 193 2448
rect 187 2446 193 2447
rect 214 2447 215 2448
rect 219 2447 220 2451
rect 299 2449 300 2453
rect 304 2449 305 2453
rect 1515 2453 1521 2454
rect 299 2448 305 2449
rect 382 2451 388 2452
rect 214 2446 220 2447
rect 382 2447 383 2451
rect 387 2450 388 2451
rect 443 2451 449 2452
rect 443 2450 444 2451
rect 387 2448 444 2450
rect 387 2447 388 2448
rect 382 2446 388 2447
rect 443 2447 444 2448
rect 448 2447 449 2451
rect 443 2446 449 2447
rect 462 2451 468 2452
rect 462 2447 463 2451
rect 467 2450 468 2451
rect 595 2451 601 2452
rect 595 2450 596 2451
rect 467 2448 596 2450
rect 467 2447 468 2448
rect 462 2446 468 2447
rect 595 2447 596 2448
rect 600 2447 601 2451
rect 595 2446 601 2447
rect 614 2451 620 2452
rect 614 2447 615 2451
rect 619 2450 620 2451
rect 747 2451 753 2452
rect 747 2450 748 2451
rect 619 2448 748 2450
rect 619 2447 620 2448
rect 614 2446 620 2447
rect 747 2447 748 2448
rect 752 2447 753 2451
rect 747 2446 753 2447
rect 891 2451 897 2452
rect 891 2447 892 2451
rect 896 2450 897 2451
rect 918 2451 924 2452
rect 918 2450 919 2451
rect 896 2448 919 2450
rect 896 2447 897 2448
rect 891 2446 897 2447
rect 918 2447 919 2448
rect 923 2447 924 2451
rect 918 2446 924 2447
rect 1027 2451 1036 2452
rect 1027 2447 1028 2451
rect 1035 2447 1036 2451
rect 1027 2446 1036 2447
rect 1155 2451 1161 2452
rect 1155 2447 1156 2451
rect 1160 2450 1161 2451
rect 1182 2451 1188 2452
rect 1182 2450 1183 2451
rect 1160 2448 1183 2450
rect 1160 2447 1161 2448
rect 1155 2446 1161 2447
rect 1182 2447 1183 2448
rect 1187 2447 1188 2451
rect 1182 2446 1188 2447
rect 1283 2451 1289 2452
rect 1283 2447 1284 2451
rect 1288 2450 1289 2451
rect 1310 2451 1316 2452
rect 1310 2450 1311 2451
rect 1288 2448 1311 2450
rect 1288 2447 1289 2448
rect 1283 2446 1289 2447
rect 1310 2447 1311 2448
rect 1315 2447 1316 2451
rect 1310 2446 1316 2447
rect 1334 2451 1340 2452
rect 1334 2447 1335 2451
rect 1339 2450 1340 2451
rect 1403 2451 1409 2452
rect 1403 2450 1404 2451
rect 1339 2448 1404 2450
rect 1339 2447 1340 2448
rect 1334 2446 1340 2447
rect 1403 2447 1404 2448
rect 1408 2447 1409 2451
rect 1515 2449 1516 2453
rect 1520 2449 1521 2453
rect 1806 2453 1807 2457
rect 1811 2453 1812 2457
rect 2014 2456 2015 2460
rect 2019 2456 2020 2460
rect 2014 2455 2020 2456
rect 2198 2460 2204 2461
rect 2198 2456 2199 2460
rect 2203 2456 2204 2460
rect 2198 2455 2204 2456
rect 2366 2460 2372 2461
rect 2366 2456 2367 2460
rect 2371 2456 2372 2460
rect 2366 2455 2372 2456
rect 2526 2460 2532 2461
rect 2526 2456 2527 2460
rect 2531 2456 2532 2460
rect 2526 2455 2532 2456
rect 2670 2460 2676 2461
rect 2670 2456 2671 2460
rect 2675 2456 2676 2460
rect 2670 2455 2676 2456
rect 2806 2460 2812 2461
rect 2806 2456 2807 2460
rect 2811 2456 2812 2460
rect 2806 2455 2812 2456
rect 2926 2460 2932 2461
rect 2926 2456 2927 2460
rect 2931 2456 2932 2460
rect 2926 2455 2932 2456
rect 3046 2460 3052 2461
rect 3046 2456 3047 2460
rect 3051 2456 3052 2460
rect 3046 2455 3052 2456
rect 3158 2460 3164 2461
rect 3158 2456 3159 2460
rect 3163 2456 3164 2460
rect 3158 2455 3164 2456
rect 3270 2460 3276 2461
rect 3270 2456 3271 2460
rect 3275 2456 3276 2460
rect 3270 2455 3276 2456
rect 3366 2460 3372 2461
rect 3366 2456 3367 2460
rect 3371 2456 3372 2460
rect 3366 2455 3372 2456
rect 3462 2457 3468 2458
rect 1806 2452 1812 2453
rect 3462 2453 3463 2457
rect 3467 2453 3468 2457
rect 3462 2452 3468 2453
rect 1515 2448 1521 2449
rect 1534 2451 1540 2452
rect 1403 2446 1409 2447
rect 1534 2447 1535 2451
rect 1539 2450 1540 2451
rect 1627 2451 1633 2452
rect 1627 2450 1628 2451
rect 1539 2448 1628 2450
rect 1539 2447 1540 2448
rect 1534 2446 1540 2447
rect 1627 2447 1628 2448
rect 1632 2447 1633 2451
rect 1627 2446 1633 2447
rect 1646 2451 1652 2452
rect 1646 2447 1647 2451
rect 1651 2450 1652 2451
rect 1723 2451 1729 2452
rect 1723 2450 1724 2451
rect 1651 2448 1724 2450
rect 1651 2447 1652 2448
rect 1646 2446 1652 2447
rect 1723 2447 1724 2448
rect 1728 2447 1729 2451
rect 1723 2446 1729 2447
rect 2086 2451 2092 2452
rect 2086 2447 2087 2451
rect 2091 2447 2092 2451
rect 2086 2446 2092 2447
rect 2270 2451 2276 2452
rect 2270 2447 2271 2451
rect 2275 2447 2276 2451
rect 2270 2446 2276 2447
rect 2430 2451 2436 2452
rect 2430 2447 2431 2451
rect 2435 2447 2436 2451
rect 2646 2451 2652 2452
rect 2646 2450 2647 2451
rect 2601 2448 2647 2450
rect 2430 2446 2436 2447
rect 2646 2447 2647 2448
rect 2651 2447 2652 2451
rect 2646 2446 2652 2447
rect 2742 2451 2748 2452
rect 2742 2447 2743 2451
rect 2747 2447 2748 2451
rect 2742 2446 2748 2447
rect 2878 2451 2884 2452
rect 2878 2447 2879 2451
rect 2883 2447 2884 2451
rect 2878 2446 2884 2447
rect 2998 2451 3004 2452
rect 2998 2447 2999 2451
rect 3003 2447 3004 2451
rect 2998 2446 3004 2447
rect 3118 2451 3124 2452
rect 3118 2447 3119 2451
rect 3123 2447 3124 2451
rect 3118 2446 3124 2447
rect 3230 2451 3236 2452
rect 3230 2447 3231 2451
rect 3235 2447 3236 2451
rect 3230 2446 3236 2447
rect 3238 2451 3244 2452
rect 3238 2447 3239 2451
rect 3243 2450 3244 2451
rect 3430 2451 3436 2452
rect 3243 2448 3313 2450
rect 3243 2447 3244 2448
rect 3238 2446 3244 2447
rect 3430 2447 3431 2451
rect 3435 2447 3436 2451
rect 3430 2446 3436 2447
rect 2014 2441 2020 2442
rect 1806 2440 1812 2441
rect 1806 2436 1807 2440
rect 1811 2436 1812 2440
rect 2014 2437 2015 2441
rect 2019 2437 2020 2441
rect 2014 2436 2020 2437
rect 2198 2441 2204 2442
rect 2198 2437 2199 2441
rect 2203 2437 2204 2441
rect 2198 2436 2204 2437
rect 2366 2441 2372 2442
rect 2366 2437 2367 2441
rect 2371 2437 2372 2441
rect 2366 2436 2372 2437
rect 2526 2441 2532 2442
rect 2526 2437 2527 2441
rect 2531 2437 2532 2441
rect 2526 2436 2532 2437
rect 2670 2441 2676 2442
rect 2670 2437 2671 2441
rect 2675 2437 2676 2441
rect 2670 2436 2676 2437
rect 2806 2441 2812 2442
rect 2806 2437 2807 2441
rect 2811 2437 2812 2441
rect 2806 2436 2812 2437
rect 2926 2441 2932 2442
rect 2926 2437 2927 2441
rect 2931 2437 2932 2441
rect 2926 2436 2932 2437
rect 3046 2441 3052 2442
rect 3046 2437 3047 2441
rect 3051 2437 3052 2441
rect 3046 2436 3052 2437
rect 3158 2441 3164 2442
rect 3158 2437 3159 2441
rect 3163 2437 3164 2441
rect 3158 2436 3164 2437
rect 3270 2441 3276 2442
rect 3270 2437 3271 2441
rect 3275 2437 3276 2441
rect 3270 2436 3276 2437
rect 3366 2441 3372 2442
rect 3366 2437 3367 2441
rect 3371 2437 3372 2441
rect 3366 2436 3372 2437
rect 3462 2440 3468 2441
rect 3462 2436 3463 2440
rect 3467 2436 3468 2440
rect 1806 2435 1812 2436
rect 3462 2435 3468 2436
rect 187 2423 193 2424
rect 187 2419 188 2423
rect 192 2422 193 2423
rect 206 2423 212 2424
rect 206 2422 207 2423
rect 192 2420 207 2422
rect 192 2419 193 2420
rect 187 2418 193 2419
rect 206 2419 207 2420
rect 211 2419 212 2423
rect 206 2418 212 2419
rect 231 2423 237 2424
rect 231 2419 232 2423
rect 236 2422 237 2423
rect 291 2423 297 2424
rect 291 2422 292 2423
rect 236 2420 292 2422
rect 236 2419 237 2420
rect 231 2418 237 2419
rect 291 2419 292 2420
rect 296 2419 297 2423
rect 291 2418 297 2419
rect 310 2423 316 2424
rect 310 2419 311 2423
rect 315 2422 316 2423
rect 443 2423 449 2424
rect 443 2422 444 2423
rect 315 2420 444 2422
rect 315 2419 316 2420
rect 310 2418 316 2419
rect 443 2419 444 2420
rect 448 2419 449 2423
rect 443 2418 449 2419
rect 462 2423 468 2424
rect 462 2419 463 2423
rect 467 2422 468 2423
rect 603 2423 609 2424
rect 603 2422 604 2423
rect 467 2420 604 2422
rect 467 2419 468 2420
rect 462 2418 468 2419
rect 603 2419 604 2420
rect 608 2419 609 2423
rect 603 2418 609 2419
rect 622 2423 628 2424
rect 622 2419 623 2423
rect 627 2422 628 2423
rect 771 2423 777 2424
rect 771 2422 772 2423
rect 627 2420 772 2422
rect 627 2419 628 2420
rect 622 2418 628 2419
rect 771 2419 772 2420
rect 776 2419 777 2423
rect 771 2418 777 2419
rect 918 2423 924 2424
rect 918 2419 919 2423
rect 923 2422 924 2423
rect 947 2423 953 2424
rect 947 2422 948 2423
rect 923 2420 948 2422
rect 923 2419 924 2420
rect 918 2418 924 2419
rect 947 2419 948 2420
rect 952 2419 953 2423
rect 947 2418 953 2419
rect 966 2423 972 2424
rect 966 2419 967 2423
rect 971 2422 972 2423
rect 1115 2423 1121 2424
rect 1115 2422 1116 2423
rect 971 2420 1116 2422
rect 971 2419 972 2420
rect 966 2418 972 2419
rect 1115 2419 1116 2420
rect 1120 2419 1121 2423
rect 1115 2418 1121 2419
rect 1291 2423 1297 2424
rect 1291 2419 1292 2423
rect 1296 2422 1297 2423
rect 1318 2423 1324 2424
rect 1318 2422 1319 2423
rect 1296 2420 1319 2422
rect 1296 2419 1297 2420
rect 1291 2418 1297 2419
rect 1318 2419 1319 2420
rect 1323 2419 1324 2423
rect 1318 2418 1324 2419
rect 1467 2423 1473 2424
rect 1467 2419 1468 2423
rect 1472 2422 1473 2423
rect 1575 2423 1581 2424
rect 1575 2422 1576 2423
rect 1472 2420 1576 2422
rect 1472 2419 1473 2420
rect 1467 2418 1473 2419
rect 1575 2419 1576 2420
rect 1580 2419 1581 2423
rect 1575 2418 1581 2419
rect 1598 2423 1604 2424
rect 1598 2419 1599 2423
rect 1603 2422 1604 2423
rect 1643 2423 1649 2424
rect 1643 2422 1644 2423
rect 1603 2420 1644 2422
rect 1603 2419 1604 2420
rect 1598 2418 1604 2419
rect 1643 2419 1644 2420
rect 1648 2419 1649 2423
rect 1643 2418 1649 2419
rect 134 2408 140 2409
rect 110 2405 116 2406
rect 110 2401 111 2405
rect 115 2401 116 2405
rect 134 2404 135 2408
rect 139 2404 140 2408
rect 134 2403 140 2404
rect 238 2408 244 2409
rect 238 2404 239 2408
rect 243 2404 244 2408
rect 238 2403 244 2404
rect 390 2408 396 2409
rect 390 2404 391 2408
rect 395 2404 396 2408
rect 390 2403 396 2404
rect 550 2408 556 2409
rect 550 2404 551 2408
rect 555 2404 556 2408
rect 550 2403 556 2404
rect 718 2408 724 2409
rect 718 2404 719 2408
rect 723 2404 724 2408
rect 718 2403 724 2404
rect 894 2408 900 2409
rect 894 2404 895 2408
rect 899 2404 900 2408
rect 894 2403 900 2404
rect 1062 2408 1068 2409
rect 1062 2404 1063 2408
rect 1067 2404 1068 2408
rect 1062 2403 1068 2404
rect 1238 2408 1244 2409
rect 1414 2408 1420 2409
rect 1238 2404 1239 2408
rect 1243 2404 1244 2408
rect 1334 2407 1340 2408
rect 1334 2406 1335 2407
rect 1238 2403 1244 2404
rect 1312 2404 1335 2406
rect 110 2400 116 2401
rect 231 2399 237 2400
rect 231 2398 232 2399
rect 209 2396 232 2398
rect 231 2395 232 2396
rect 236 2395 237 2399
rect 231 2394 237 2395
rect 310 2399 316 2400
rect 310 2395 311 2399
rect 315 2395 316 2399
rect 310 2394 316 2395
rect 462 2399 468 2400
rect 462 2395 463 2399
rect 467 2395 468 2399
rect 462 2394 468 2395
rect 622 2399 628 2400
rect 622 2395 623 2399
rect 627 2395 628 2399
rect 622 2394 628 2395
rect 630 2399 636 2400
rect 630 2395 631 2399
rect 635 2398 636 2399
rect 966 2399 972 2400
rect 635 2396 761 2398
rect 635 2395 636 2396
rect 630 2394 636 2395
rect 966 2395 967 2399
rect 971 2395 972 2399
rect 966 2394 972 2395
rect 1030 2399 1036 2400
rect 1030 2395 1031 2399
rect 1035 2398 1036 2399
rect 1035 2396 1105 2398
rect 1312 2397 1314 2404
rect 1334 2403 1335 2404
rect 1339 2403 1340 2407
rect 1414 2404 1415 2408
rect 1419 2404 1420 2408
rect 1414 2403 1420 2404
rect 1590 2408 1596 2409
rect 1590 2404 1591 2408
rect 1595 2404 1596 2408
rect 1590 2403 1596 2404
rect 1766 2405 1772 2406
rect 1334 2402 1340 2403
rect 1766 2401 1767 2405
rect 1771 2401 1772 2405
rect 1766 2400 1772 2401
rect 1318 2399 1324 2400
rect 1035 2395 1036 2396
rect 1030 2394 1036 2395
rect 1318 2395 1319 2399
rect 1323 2398 1324 2399
rect 1575 2399 1581 2400
rect 1323 2396 1457 2398
rect 1323 2395 1324 2396
rect 1318 2394 1324 2395
rect 1575 2395 1576 2399
rect 1580 2398 1581 2399
rect 1580 2396 1633 2398
rect 1580 2395 1581 2396
rect 1575 2394 1581 2395
rect 1806 2392 1812 2393
rect 3462 2392 3468 2393
rect 134 2389 140 2390
rect 110 2388 116 2389
rect 110 2384 111 2388
rect 115 2384 116 2388
rect 134 2385 135 2389
rect 139 2385 140 2389
rect 134 2384 140 2385
rect 238 2389 244 2390
rect 238 2385 239 2389
rect 243 2385 244 2389
rect 238 2384 244 2385
rect 390 2389 396 2390
rect 390 2385 391 2389
rect 395 2385 396 2389
rect 390 2384 396 2385
rect 550 2389 556 2390
rect 550 2385 551 2389
rect 555 2385 556 2389
rect 550 2384 556 2385
rect 718 2389 724 2390
rect 718 2385 719 2389
rect 723 2385 724 2389
rect 718 2384 724 2385
rect 894 2389 900 2390
rect 894 2385 895 2389
rect 899 2385 900 2389
rect 894 2384 900 2385
rect 1062 2389 1068 2390
rect 1062 2385 1063 2389
rect 1067 2385 1068 2389
rect 1062 2384 1068 2385
rect 1238 2389 1244 2390
rect 1238 2385 1239 2389
rect 1243 2385 1244 2389
rect 1238 2384 1244 2385
rect 1414 2389 1420 2390
rect 1414 2385 1415 2389
rect 1419 2385 1420 2389
rect 1414 2384 1420 2385
rect 1590 2389 1596 2390
rect 1590 2385 1591 2389
rect 1595 2385 1596 2389
rect 1590 2384 1596 2385
rect 1766 2388 1772 2389
rect 1766 2384 1767 2388
rect 1771 2384 1772 2388
rect 1806 2388 1807 2392
rect 1811 2388 1812 2392
rect 1806 2387 1812 2388
rect 1838 2391 1844 2392
rect 1838 2387 1839 2391
rect 1843 2387 1844 2391
rect 1838 2386 1844 2387
rect 2006 2391 2012 2392
rect 2006 2387 2007 2391
rect 2011 2387 2012 2391
rect 2006 2386 2012 2387
rect 2182 2391 2188 2392
rect 2182 2387 2183 2391
rect 2187 2387 2188 2391
rect 2182 2386 2188 2387
rect 2366 2391 2372 2392
rect 2366 2387 2367 2391
rect 2371 2387 2372 2391
rect 2366 2386 2372 2387
rect 2558 2391 2564 2392
rect 2558 2387 2559 2391
rect 2563 2387 2564 2391
rect 2558 2386 2564 2387
rect 2758 2391 2764 2392
rect 2758 2387 2759 2391
rect 2763 2387 2764 2391
rect 2758 2386 2764 2387
rect 2966 2391 2972 2392
rect 2966 2387 2967 2391
rect 2971 2387 2972 2391
rect 2966 2386 2972 2387
rect 3174 2391 3180 2392
rect 3174 2387 3175 2391
rect 3179 2387 3180 2391
rect 3174 2386 3180 2387
rect 3366 2391 3372 2392
rect 3366 2387 3367 2391
rect 3371 2387 3372 2391
rect 3462 2388 3463 2392
rect 3467 2388 3468 2392
rect 3462 2387 3468 2388
rect 3366 2386 3372 2387
rect 110 2383 116 2384
rect 1766 2383 1772 2384
rect 1918 2383 1924 2384
rect 1910 2379 1916 2380
rect 1806 2375 1812 2376
rect 1806 2371 1807 2375
rect 1811 2371 1812 2375
rect 1910 2375 1911 2379
rect 1915 2375 1916 2379
rect 1918 2379 1919 2383
rect 1923 2382 1924 2383
rect 2086 2383 2092 2384
rect 1923 2380 2049 2382
rect 1923 2379 1924 2380
rect 1918 2378 1924 2379
rect 2086 2379 2087 2383
rect 2091 2382 2092 2383
rect 2262 2383 2268 2384
rect 2091 2380 2225 2382
rect 2091 2379 2092 2380
rect 2086 2378 2092 2379
rect 2262 2379 2263 2383
rect 2267 2382 2268 2383
rect 2630 2383 2636 2384
rect 2267 2380 2409 2382
rect 2267 2379 2268 2380
rect 2262 2378 2268 2379
rect 2630 2379 2631 2383
rect 2635 2379 2636 2383
rect 2630 2378 2636 2379
rect 2638 2383 2644 2384
rect 2638 2379 2639 2383
rect 2643 2382 2644 2383
rect 2839 2383 2845 2384
rect 2643 2380 2801 2382
rect 2643 2379 2644 2380
rect 2638 2378 2644 2379
rect 2839 2379 2840 2383
rect 2844 2382 2845 2383
rect 3438 2383 3444 2384
rect 2844 2380 3009 2382
rect 2844 2379 2845 2380
rect 2839 2378 2845 2379
rect 3246 2379 3252 2380
rect 1910 2374 1916 2375
rect 3246 2375 3247 2379
rect 3251 2375 3252 2379
rect 3438 2379 3439 2383
rect 3443 2379 3444 2383
rect 3438 2378 3444 2379
rect 3246 2374 3252 2375
rect 3462 2375 3468 2376
rect 1806 2370 1812 2371
rect 1838 2372 1844 2373
rect 1838 2368 1839 2372
rect 1843 2368 1844 2372
rect 1838 2367 1844 2368
rect 2006 2372 2012 2373
rect 2006 2368 2007 2372
rect 2011 2368 2012 2372
rect 2006 2367 2012 2368
rect 2182 2372 2188 2373
rect 2182 2368 2183 2372
rect 2187 2368 2188 2372
rect 2182 2367 2188 2368
rect 2366 2372 2372 2373
rect 2366 2368 2367 2372
rect 2371 2368 2372 2372
rect 2366 2367 2372 2368
rect 2558 2372 2564 2373
rect 2558 2368 2559 2372
rect 2563 2368 2564 2372
rect 2558 2367 2564 2368
rect 2758 2372 2764 2373
rect 2758 2368 2759 2372
rect 2763 2368 2764 2372
rect 2758 2367 2764 2368
rect 2966 2372 2972 2373
rect 2966 2368 2967 2372
rect 2971 2368 2972 2372
rect 2966 2367 2972 2368
rect 3174 2372 3180 2373
rect 3174 2368 3175 2372
rect 3179 2368 3180 2372
rect 3174 2367 3180 2368
rect 3366 2372 3372 2373
rect 3366 2368 3367 2372
rect 3371 2368 3372 2372
rect 3462 2371 3463 2375
rect 3467 2371 3468 2375
rect 3462 2370 3468 2371
rect 3366 2367 3372 2368
rect 1891 2355 1897 2356
rect 1891 2351 1892 2355
rect 1896 2354 1897 2355
rect 1918 2355 1924 2356
rect 1918 2354 1919 2355
rect 1896 2352 1919 2354
rect 1896 2351 1897 2352
rect 1891 2350 1897 2351
rect 1918 2351 1919 2352
rect 1923 2351 1924 2355
rect 1918 2350 1924 2351
rect 2059 2355 2065 2356
rect 2059 2351 2060 2355
rect 2064 2354 2065 2355
rect 2086 2355 2092 2356
rect 2086 2354 2087 2355
rect 2064 2352 2087 2354
rect 2064 2351 2065 2352
rect 2059 2350 2065 2351
rect 2086 2351 2087 2352
rect 2091 2351 2092 2355
rect 2086 2350 2092 2351
rect 2235 2355 2241 2356
rect 2235 2351 2236 2355
rect 2240 2354 2241 2355
rect 2262 2355 2268 2356
rect 2262 2354 2263 2355
rect 2240 2352 2263 2354
rect 2240 2351 2241 2352
rect 2235 2350 2241 2351
rect 2262 2351 2263 2352
rect 2267 2351 2268 2355
rect 2262 2350 2268 2351
rect 2419 2355 2425 2356
rect 2419 2351 2420 2355
rect 2424 2354 2425 2355
rect 2430 2355 2436 2356
rect 2430 2354 2431 2355
rect 2424 2352 2431 2354
rect 2424 2351 2425 2352
rect 2419 2350 2425 2351
rect 2430 2351 2431 2352
rect 2435 2351 2436 2355
rect 2430 2350 2436 2351
rect 2611 2355 2617 2356
rect 2611 2351 2612 2355
rect 2616 2354 2617 2355
rect 2638 2355 2644 2356
rect 2638 2354 2639 2355
rect 2616 2352 2639 2354
rect 2616 2351 2617 2352
rect 2611 2350 2617 2351
rect 2638 2351 2639 2352
rect 2643 2351 2644 2355
rect 2638 2350 2644 2351
rect 2811 2355 2817 2356
rect 2811 2351 2812 2355
rect 2816 2354 2817 2355
rect 2839 2355 2845 2356
rect 2839 2354 2840 2355
rect 2816 2352 2840 2354
rect 2816 2351 2817 2352
rect 2811 2350 2817 2351
rect 2839 2351 2840 2352
rect 2844 2351 2845 2355
rect 2839 2350 2845 2351
rect 3019 2355 3025 2356
rect 3019 2351 3020 2355
rect 3024 2354 3025 2355
rect 3038 2355 3044 2356
rect 3038 2354 3039 2355
rect 3024 2352 3039 2354
rect 3024 2351 3025 2352
rect 3019 2350 3025 2351
rect 3038 2351 3039 2352
rect 3043 2351 3044 2355
rect 3038 2350 3044 2351
rect 3227 2355 3233 2356
rect 3227 2351 3228 2355
rect 3232 2354 3233 2355
rect 3238 2355 3244 2356
rect 3238 2354 3239 2355
rect 3232 2352 3239 2354
rect 3232 2351 3233 2352
rect 3227 2350 3233 2351
rect 3238 2351 3239 2352
rect 3243 2351 3244 2355
rect 3238 2350 3244 2351
rect 3419 2355 3425 2356
rect 3419 2351 3420 2355
rect 3424 2354 3425 2355
rect 3438 2355 3444 2356
rect 3438 2354 3439 2355
rect 3424 2352 3439 2354
rect 3424 2351 3425 2352
rect 3419 2350 3425 2351
rect 3438 2351 3439 2352
rect 3443 2351 3444 2355
rect 3438 2350 3444 2351
rect 1910 2343 1916 2344
rect 1910 2339 1911 2343
rect 1915 2342 1916 2343
rect 1939 2343 1945 2344
rect 1939 2342 1940 2343
rect 1915 2340 1940 2342
rect 1915 2339 1916 2340
rect 1910 2338 1916 2339
rect 1939 2339 1940 2340
rect 1944 2339 1945 2343
rect 1939 2338 1945 2339
rect 1958 2343 1964 2344
rect 1958 2339 1959 2343
rect 1963 2342 1964 2343
rect 2067 2343 2073 2344
rect 2067 2342 2068 2343
rect 1963 2340 2068 2342
rect 1963 2339 1964 2340
rect 1958 2338 1964 2339
rect 2067 2339 2068 2340
rect 2072 2339 2073 2343
rect 2067 2338 2073 2339
rect 2086 2343 2092 2344
rect 2086 2339 2087 2343
rect 2091 2342 2092 2343
rect 2203 2343 2209 2344
rect 2203 2342 2204 2343
rect 2091 2340 2204 2342
rect 2091 2339 2092 2340
rect 2086 2338 2092 2339
rect 2203 2339 2204 2340
rect 2208 2339 2209 2343
rect 2203 2338 2209 2339
rect 2222 2343 2228 2344
rect 2222 2339 2223 2343
rect 2227 2342 2228 2343
rect 2355 2343 2361 2344
rect 2355 2342 2356 2343
rect 2227 2340 2356 2342
rect 2227 2339 2228 2340
rect 2222 2338 2228 2339
rect 2355 2339 2356 2340
rect 2360 2339 2361 2343
rect 2355 2338 2361 2339
rect 2515 2343 2521 2344
rect 2515 2339 2516 2343
rect 2520 2342 2521 2343
rect 2559 2343 2565 2344
rect 2559 2342 2560 2343
rect 2520 2340 2560 2342
rect 2520 2339 2521 2340
rect 2515 2338 2521 2339
rect 2559 2339 2560 2340
rect 2564 2339 2565 2343
rect 2559 2338 2565 2339
rect 2599 2343 2605 2344
rect 2599 2339 2600 2343
rect 2604 2342 2605 2343
rect 2699 2343 2705 2344
rect 2699 2342 2700 2343
rect 2604 2340 2700 2342
rect 2604 2339 2605 2340
rect 2599 2338 2605 2339
rect 2699 2339 2700 2340
rect 2704 2339 2705 2343
rect 2699 2338 2705 2339
rect 2718 2343 2724 2344
rect 2718 2339 2719 2343
rect 2723 2342 2724 2343
rect 2891 2343 2897 2344
rect 2891 2342 2892 2343
rect 2723 2340 2892 2342
rect 2723 2339 2724 2340
rect 2718 2338 2724 2339
rect 2891 2339 2892 2340
rect 2896 2339 2897 2343
rect 2891 2338 2897 2339
rect 2910 2343 2916 2344
rect 2910 2339 2911 2343
rect 2915 2342 2916 2343
rect 3099 2343 3105 2344
rect 3099 2342 3100 2343
rect 2915 2340 3100 2342
rect 2915 2339 2916 2340
rect 2910 2338 2916 2339
rect 3099 2339 3100 2340
rect 3104 2339 3105 2343
rect 3099 2338 3105 2339
rect 3246 2343 3252 2344
rect 3246 2339 3247 2343
rect 3251 2342 3252 2343
rect 3307 2343 3313 2344
rect 3307 2342 3308 2343
rect 3251 2340 3308 2342
rect 3251 2339 3252 2340
rect 3246 2338 3252 2339
rect 3307 2339 3308 2340
rect 3312 2339 3313 2343
rect 3307 2338 3313 2339
rect 110 2336 116 2337
rect 1766 2336 1772 2337
rect 110 2332 111 2336
rect 115 2332 116 2336
rect 110 2331 116 2332
rect 374 2335 380 2336
rect 374 2331 375 2335
rect 379 2331 380 2335
rect 374 2330 380 2331
rect 478 2335 484 2336
rect 478 2331 479 2335
rect 483 2331 484 2335
rect 478 2330 484 2331
rect 598 2335 604 2336
rect 598 2331 599 2335
rect 603 2331 604 2335
rect 598 2330 604 2331
rect 718 2335 724 2336
rect 718 2331 719 2335
rect 723 2331 724 2335
rect 718 2330 724 2331
rect 846 2335 852 2336
rect 846 2331 847 2335
rect 851 2331 852 2335
rect 846 2330 852 2331
rect 974 2335 980 2336
rect 974 2331 975 2335
rect 979 2331 980 2335
rect 974 2330 980 2331
rect 1102 2335 1108 2336
rect 1102 2331 1103 2335
rect 1107 2331 1108 2335
rect 1102 2330 1108 2331
rect 1238 2335 1244 2336
rect 1238 2331 1239 2335
rect 1243 2331 1244 2335
rect 1238 2330 1244 2331
rect 1374 2335 1380 2336
rect 1374 2331 1375 2335
rect 1379 2331 1380 2335
rect 1374 2330 1380 2331
rect 1510 2335 1516 2336
rect 1510 2331 1511 2335
rect 1515 2331 1516 2335
rect 1766 2332 1767 2336
rect 1771 2332 1772 2336
rect 1766 2331 1772 2332
rect 1510 2330 1516 2331
rect 1886 2328 1892 2329
rect 694 2327 700 2328
rect 446 2323 452 2324
rect 110 2319 116 2320
rect 110 2315 111 2319
rect 115 2315 116 2319
rect 446 2319 447 2323
rect 451 2319 452 2323
rect 446 2318 452 2319
rect 550 2323 556 2324
rect 550 2319 551 2323
rect 555 2319 556 2323
rect 550 2318 556 2319
rect 670 2323 676 2324
rect 670 2319 671 2323
rect 675 2319 676 2323
rect 694 2323 695 2327
rect 699 2326 700 2327
rect 918 2327 924 2328
rect 699 2324 761 2326
rect 699 2323 700 2324
rect 694 2322 700 2323
rect 918 2323 919 2327
rect 923 2323 924 2327
rect 918 2322 924 2323
rect 926 2327 932 2328
rect 926 2323 927 2327
rect 931 2326 932 2327
rect 1054 2327 1060 2328
rect 931 2324 1017 2326
rect 931 2323 932 2324
rect 926 2322 932 2323
rect 1054 2323 1055 2327
rect 1059 2326 1060 2327
rect 1598 2327 1604 2328
rect 1598 2326 1599 2327
rect 1059 2324 1145 2326
rect 1585 2324 1599 2326
rect 1059 2323 1060 2324
rect 1054 2322 1060 2323
rect 1310 2323 1316 2324
rect 670 2318 676 2319
rect 1310 2319 1311 2323
rect 1315 2319 1316 2323
rect 1310 2318 1316 2319
rect 1446 2323 1452 2324
rect 1446 2319 1447 2323
rect 1451 2319 1452 2323
rect 1598 2323 1599 2324
rect 1603 2323 1604 2327
rect 1598 2322 1604 2323
rect 1806 2325 1812 2326
rect 1806 2321 1807 2325
rect 1811 2321 1812 2325
rect 1886 2324 1887 2328
rect 1891 2324 1892 2328
rect 1886 2323 1892 2324
rect 2014 2328 2020 2329
rect 2014 2324 2015 2328
rect 2019 2324 2020 2328
rect 2014 2323 2020 2324
rect 2150 2328 2156 2329
rect 2150 2324 2151 2328
rect 2155 2324 2156 2328
rect 2150 2323 2156 2324
rect 2302 2328 2308 2329
rect 2302 2324 2303 2328
rect 2307 2324 2308 2328
rect 2302 2323 2308 2324
rect 2462 2328 2468 2329
rect 2462 2324 2463 2328
rect 2467 2324 2468 2328
rect 2462 2323 2468 2324
rect 2646 2328 2652 2329
rect 2646 2324 2647 2328
rect 2651 2324 2652 2328
rect 2646 2323 2652 2324
rect 2838 2328 2844 2329
rect 2838 2324 2839 2328
rect 2843 2324 2844 2328
rect 2838 2323 2844 2324
rect 3046 2328 3052 2329
rect 3046 2324 3047 2328
rect 3051 2324 3052 2328
rect 3046 2323 3052 2324
rect 3254 2328 3260 2329
rect 3254 2324 3255 2328
rect 3259 2324 3260 2328
rect 3254 2323 3260 2324
rect 3462 2325 3468 2326
rect 1806 2320 1812 2321
rect 3462 2321 3463 2325
rect 3467 2321 3468 2325
rect 3462 2320 3468 2321
rect 1446 2318 1452 2319
rect 1766 2319 1772 2320
rect 110 2314 116 2315
rect 374 2316 380 2317
rect 374 2312 375 2316
rect 379 2312 380 2316
rect 374 2311 380 2312
rect 478 2316 484 2317
rect 478 2312 479 2316
rect 483 2312 484 2316
rect 478 2311 484 2312
rect 598 2316 604 2317
rect 598 2312 599 2316
rect 603 2312 604 2316
rect 598 2311 604 2312
rect 718 2316 724 2317
rect 718 2312 719 2316
rect 723 2312 724 2316
rect 718 2311 724 2312
rect 846 2316 852 2317
rect 846 2312 847 2316
rect 851 2312 852 2316
rect 846 2311 852 2312
rect 974 2316 980 2317
rect 974 2312 975 2316
rect 979 2312 980 2316
rect 974 2311 980 2312
rect 1102 2316 1108 2317
rect 1102 2312 1103 2316
rect 1107 2312 1108 2316
rect 1102 2311 1108 2312
rect 1238 2316 1244 2317
rect 1238 2312 1239 2316
rect 1243 2312 1244 2316
rect 1238 2311 1244 2312
rect 1374 2316 1380 2317
rect 1374 2312 1375 2316
rect 1379 2312 1380 2316
rect 1374 2311 1380 2312
rect 1510 2316 1516 2317
rect 1510 2312 1511 2316
rect 1515 2312 1516 2316
rect 1766 2315 1767 2319
rect 1771 2315 1772 2319
rect 1766 2314 1772 2315
rect 1958 2319 1964 2320
rect 1958 2315 1959 2319
rect 1963 2315 1964 2319
rect 1958 2314 1964 2315
rect 2086 2319 2092 2320
rect 2086 2315 2087 2319
rect 2091 2315 2092 2319
rect 2086 2314 2092 2315
rect 2222 2319 2228 2320
rect 2222 2315 2223 2319
rect 2227 2315 2228 2319
rect 2222 2314 2228 2315
rect 2230 2319 2236 2320
rect 2230 2315 2231 2319
rect 2235 2318 2236 2319
rect 2599 2319 2605 2320
rect 2599 2318 2600 2319
rect 2235 2316 2345 2318
rect 2537 2316 2600 2318
rect 2235 2315 2236 2316
rect 2230 2314 2236 2315
rect 2599 2315 2600 2316
rect 2604 2315 2605 2319
rect 2599 2314 2605 2315
rect 2718 2319 2724 2320
rect 2718 2315 2719 2319
rect 2723 2315 2724 2319
rect 2718 2314 2724 2315
rect 2910 2319 2916 2320
rect 2910 2315 2911 2319
rect 2915 2315 2916 2319
rect 2910 2314 2916 2315
rect 3038 2319 3044 2320
rect 3038 2315 3039 2319
rect 3043 2318 3044 2319
rect 3318 2319 3324 2320
rect 3043 2316 3089 2318
rect 3043 2315 3044 2316
rect 3038 2314 3044 2315
rect 3318 2315 3319 2319
rect 3323 2315 3324 2319
rect 3318 2314 3324 2315
rect 1510 2311 1516 2312
rect 1886 2309 1892 2310
rect 1806 2308 1812 2309
rect 630 2307 636 2308
rect 630 2306 631 2307
rect 428 2304 631 2306
rect 428 2302 430 2304
rect 630 2303 631 2304
rect 635 2303 636 2307
rect 1806 2304 1807 2308
rect 1811 2304 1812 2308
rect 1886 2305 1887 2309
rect 1891 2305 1892 2309
rect 1886 2304 1892 2305
rect 2014 2309 2020 2310
rect 2014 2305 2015 2309
rect 2019 2305 2020 2309
rect 2014 2304 2020 2305
rect 2150 2309 2156 2310
rect 2150 2305 2151 2309
rect 2155 2305 2156 2309
rect 2150 2304 2156 2305
rect 2302 2309 2308 2310
rect 2302 2305 2303 2309
rect 2307 2305 2308 2309
rect 2302 2304 2308 2305
rect 2462 2309 2468 2310
rect 2462 2305 2463 2309
rect 2467 2305 2468 2309
rect 2462 2304 2468 2305
rect 2646 2309 2652 2310
rect 2646 2305 2647 2309
rect 2651 2305 2652 2309
rect 2646 2304 2652 2305
rect 2838 2309 2844 2310
rect 2838 2305 2839 2309
rect 2843 2305 2844 2309
rect 2838 2304 2844 2305
rect 3046 2309 3052 2310
rect 3046 2305 3047 2309
rect 3051 2305 3052 2309
rect 3046 2304 3052 2305
rect 3254 2309 3260 2310
rect 3254 2305 3255 2309
rect 3259 2305 3260 2309
rect 3254 2304 3260 2305
rect 3462 2308 3468 2309
rect 3462 2304 3463 2308
rect 3467 2304 3468 2308
rect 1806 2303 1812 2304
rect 3462 2303 3468 2304
rect 630 2302 636 2303
rect 427 2301 433 2302
rect 427 2297 428 2301
rect 432 2297 433 2301
rect 427 2296 433 2297
rect 446 2299 452 2300
rect 446 2295 447 2299
rect 451 2298 452 2299
rect 531 2299 537 2300
rect 531 2298 532 2299
rect 451 2296 532 2298
rect 451 2295 452 2296
rect 446 2294 452 2295
rect 531 2295 532 2296
rect 536 2295 537 2299
rect 531 2294 537 2295
rect 550 2299 556 2300
rect 550 2295 551 2299
rect 555 2298 556 2299
rect 651 2299 657 2300
rect 651 2298 652 2299
rect 555 2296 652 2298
rect 555 2295 556 2296
rect 550 2294 556 2295
rect 651 2295 652 2296
rect 656 2295 657 2299
rect 651 2294 657 2295
rect 670 2299 676 2300
rect 670 2295 671 2299
rect 675 2298 676 2299
rect 771 2299 777 2300
rect 771 2298 772 2299
rect 675 2296 772 2298
rect 675 2295 676 2296
rect 670 2294 676 2295
rect 771 2295 772 2296
rect 776 2295 777 2299
rect 771 2294 777 2295
rect 899 2299 905 2300
rect 899 2295 900 2299
rect 904 2298 905 2299
rect 926 2299 932 2300
rect 926 2298 927 2299
rect 904 2296 927 2298
rect 904 2295 905 2296
rect 899 2294 905 2295
rect 926 2295 927 2296
rect 931 2295 932 2299
rect 926 2294 932 2295
rect 1027 2299 1033 2300
rect 1027 2295 1028 2299
rect 1032 2298 1033 2299
rect 1054 2299 1060 2300
rect 1054 2298 1055 2299
rect 1032 2296 1055 2298
rect 1032 2295 1033 2296
rect 1027 2294 1033 2295
rect 1054 2295 1055 2296
rect 1059 2295 1060 2299
rect 1054 2294 1060 2295
rect 1150 2299 1161 2300
rect 1150 2295 1151 2299
rect 1155 2295 1156 2299
rect 1160 2295 1161 2299
rect 1150 2294 1161 2295
rect 1262 2299 1268 2300
rect 1262 2295 1263 2299
rect 1267 2298 1268 2299
rect 1291 2299 1297 2300
rect 1291 2298 1292 2299
rect 1267 2296 1292 2298
rect 1267 2295 1268 2296
rect 1262 2294 1268 2295
rect 1291 2295 1292 2296
rect 1296 2295 1297 2299
rect 1291 2294 1297 2295
rect 1310 2299 1316 2300
rect 1310 2295 1311 2299
rect 1315 2298 1316 2299
rect 1427 2299 1433 2300
rect 1427 2298 1428 2299
rect 1315 2296 1428 2298
rect 1315 2295 1316 2296
rect 1310 2294 1316 2295
rect 1427 2295 1428 2296
rect 1432 2295 1433 2299
rect 1427 2294 1433 2295
rect 1446 2299 1452 2300
rect 1446 2295 1447 2299
rect 1451 2298 1452 2299
rect 1563 2299 1569 2300
rect 1563 2298 1564 2299
rect 1451 2296 1564 2298
rect 1451 2295 1452 2296
rect 1446 2294 1452 2295
rect 1563 2295 1564 2296
rect 1568 2295 1569 2299
rect 1563 2294 1569 2295
rect 694 2287 700 2288
rect 694 2286 695 2287
rect 628 2284 695 2286
rect 628 2282 630 2284
rect 694 2283 695 2284
rect 699 2283 700 2287
rect 694 2282 700 2283
rect 627 2281 633 2282
rect 627 2277 628 2281
rect 632 2277 633 2281
rect 627 2276 633 2277
rect 646 2279 652 2280
rect 646 2275 647 2279
rect 651 2278 652 2279
rect 715 2279 721 2280
rect 715 2278 716 2279
rect 651 2276 716 2278
rect 651 2275 652 2276
rect 646 2274 652 2275
rect 715 2275 716 2276
rect 720 2275 721 2279
rect 715 2274 721 2275
rect 811 2279 817 2280
rect 811 2275 812 2279
rect 816 2278 817 2279
rect 854 2279 860 2280
rect 854 2278 855 2279
rect 816 2276 855 2278
rect 816 2275 817 2276
rect 811 2274 817 2275
rect 854 2275 855 2276
rect 859 2275 860 2279
rect 915 2279 921 2280
rect 915 2278 916 2279
rect 854 2274 860 2275
rect 864 2276 916 2278
rect 864 2270 866 2276
rect 915 2275 916 2276
rect 920 2275 921 2279
rect 915 2274 921 2275
rect 934 2279 940 2280
rect 934 2275 935 2279
rect 939 2278 940 2279
rect 1019 2279 1025 2280
rect 1019 2278 1020 2279
rect 939 2276 1020 2278
rect 939 2275 940 2276
rect 934 2274 940 2275
rect 1019 2275 1020 2276
rect 1024 2275 1025 2279
rect 1019 2274 1025 2275
rect 1038 2279 1044 2280
rect 1038 2275 1039 2279
rect 1043 2278 1044 2279
rect 1131 2279 1137 2280
rect 1131 2278 1132 2279
rect 1043 2276 1132 2278
rect 1043 2275 1044 2276
rect 1038 2274 1044 2275
rect 1131 2275 1132 2276
rect 1136 2275 1137 2279
rect 1131 2274 1137 2275
rect 1243 2279 1249 2280
rect 1243 2275 1244 2279
rect 1248 2278 1249 2279
rect 1271 2279 1277 2280
rect 1271 2278 1272 2279
rect 1248 2276 1272 2278
rect 1248 2275 1249 2276
rect 1243 2274 1249 2275
rect 1271 2275 1272 2276
rect 1276 2275 1277 2279
rect 1271 2274 1277 2275
rect 1355 2279 1361 2280
rect 1355 2275 1356 2279
rect 1360 2278 1361 2279
rect 1383 2279 1389 2280
rect 1383 2278 1384 2279
rect 1360 2276 1384 2278
rect 1360 2275 1361 2276
rect 1355 2274 1361 2275
rect 1383 2275 1384 2276
rect 1388 2275 1389 2279
rect 1383 2274 1389 2275
rect 1407 2279 1413 2280
rect 1407 2275 1408 2279
rect 1412 2278 1413 2279
rect 1467 2279 1473 2280
rect 1467 2278 1468 2279
rect 1412 2276 1468 2278
rect 1412 2275 1413 2276
rect 1407 2274 1413 2275
rect 1467 2275 1468 2276
rect 1472 2275 1473 2279
rect 1467 2274 1473 2275
rect 856 2268 866 2270
rect 574 2264 580 2265
rect 110 2261 116 2262
rect 110 2257 111 2261
rect 115 2257 116 2261
rect 574 2260 575 2264
rect 579 2260 580 2264
rect 574 2259 580 2260
rect 662 2264 668 2265
rect 662 2260 663 2264
rect 667 2260 668 2264
rect 662 2259 668 2260
rect 758 2264 764 2265
rect 758 2260 759 2264
rect 763 2260 764 2264
rect 758 2259 764 2260
rect 110 2256 116 2257
rect 646 2255 652 2256
rect 646 2251 647 2255
rect 651 2251 652 2255
rect 646 2250 652 2251
rect 734 2255 740 2256
rect 734 2251 735 2255
rect 739 2251 740 2255
rect 856 2254 858 2268
rect 862 2264 868 2265
rect 862 2260 863 2264
rect 867 2260 868 2264
rect 862 2259 868 2260
rect 966 2264 972 2265
rect 966 2260 967 2264
rect 971 2260 972 2264
rect 966 2259 972 2260
rect 1078 2264 1084 2265
rect 1078 2260 1079 2264
rect 1083 2260 1084 2264
rect 1078 2259 1084 2260
rect 1190 2264 1196 2265
rect 1190 2260 1191 2264
rect 1195 2260 1196 2264
rect 1190 2259 1196 2260
rect 1302 2264 1308 2265
rect 1302 2260 1303 2264
rect 1307 2260 1308 2264
rect 1302 2259 1308 2260
rect 1414 2264 1420 2265
rect 1414 2260 1415 2264
rect 1419 2260 1420 2264
rect 1414 2259 1420 2260
rect 1766 2261 1772 2262
rect 1766 2257 1767 2261
rect 1771 2257 1772 2261
rect 1766 2256 1772 2257
rect 1806 2260 1812 2261
rect 3462 2260 3468 2261
rect 1806 2256 1807 2260
rect 1811 2256 1812 2260
rect 833 2252 858 2254
rect 934 2255 940 2256
rect 734 2250 740 2251
rect 934 2251 935 2255
rect 939 2251 940 2255
rect 934 2250 940 2251
rect 1038 2255 1044 2256
rect 1038 2251 1039 2255
rect 1043 2251 1044 2255
rect 1038 2250 1044 2251
rect 1150 2255 1156 2256
rect 1150 2251 1151 2255
rect 1155 2251 1156 2255
rect 1150 2250 1156 2251
rect 1262 2255 1268 2256
rect 1262 2251 1263 2255
rect 1267 2251 1268 2255
rect 1262 2250 1268 2251
rect 1271 2255 1277 2256
rect 1271 2251 1272 2255
rect 1276 2254 1277 2255
rect 1383 2255 1389 2256
rect 1806 2255 1812 2256
rect 2038 2259 2044 2260
rect 2038 2255 2039 2259
rect 2043 2255 2044 2259
rect 1276 2252 1345 2254
rect 1276 2251 1277 2252
rect 1271 2250 1277 2251
rect 1383 2251 1384 2255
rect 1388 2254 1389 2255
rect 2038 2254 2044 2255
rect 2134 2259 2140 2260
rect 2134 2255 2135 2259
rect 2139 2255 2140 2259
rect 2134 2254 2140 2255
rect 2238 2259 2244 2260
rect 2238 2255 2239 2259
rect 2243 2255 2244 2259
rect 2238 2254 2244 2255
rect 2342 2259 2348 2260
rect 2342 2255 2343 2259
rect 2347 2255 2348 2259
rect 2342 2254 2348 2255
rect 2462 2259 2468 2260
rect 2462 2255 2463 2259
rect 2467 2255 2468 2259
rect 2462 2254 2468 2255
rect 2590 2259 2596 2260
rect 2590 2255 2591 2259
rect 2595 2255 2596 2259
rect 2590 2254 2596 2255
rect 2734 2259 2740 2260
rect 2734 2255 2735 2259
rect 2739 2255 2740 2259
rect 2734 2254 2740 2255
rect 2886 2259 2892 2260
rect 2886 2255 2887 2259
rect 2891 2255 2892 2259
rect 2886 2254 2892 2255
rect 3046 2259 3052 2260
rect 3046 2255 3047 2259
rect 3051 2255 3052 2259
rect 3046 2254 3052 2255
rect 3214 2259 3220 2260
rect 3214 2255 3215 2259
rect 3219 2255 3220 2259
rect 3214 2254 3220 2255
rect 3366 2259 3372 2260
rect 3366 2255 3367 2259
rect 3371 2255 3372 2259
rect 3462 2256 3463 2260
rect 3467 2256 3468 2260
rect 3462 2255 3468 2256
rect 3366 2254 3372 2255
rect 1388 2252 1457 2254
rect 1388 2251 1389 2252
rect 1383 2250 1389 2251
rect 2430 2251 2436 2252
rect 2110 2247 2116 2248
rect 574 2245 580 2246
rect 110 2244 116 2245
rect 110 2240 111 2244
rect 115 2240 116 2244
rect 574 2241 575 2245
rect 579 2241 580 2245
rect 574 2240 580 2241
rect 662 2245 668 2246
rect 662 2241 663 2245
rect 667 2241 668 2245
rect 662 2240 668 2241
rect 758 2245 764 2246
rect 758 2241 759 2245
rect 763 2241 764 2245
rect 758 2240 764 2241
rect 862 2245 868 2246
rect 862 2241 863 2245
rect 867 2241 868 2245
rect 862 2240 868 2241
rect 966 2245 972 2246
rect 966 2241 967 2245
rect 971 2241 972 2245
rect 966 2240 972 2241
rect 1078 2245 1084 2246
rect 1078 2241 1079 2245
rect 1083 2241 1084 2245
rect 1078 2240 1084 2241
rect 1190 2245 1196 2246
rect 1190 2241 1191 2245
rect 1195 2241 1196 2245
rect 1190 2240 1196 2241
rect 1302 2245 1308 2246
rect 1302 2241 1303 2245
rect 1307 2241 1308 2245
rect 1302 2240 1308 2241
rect 1414 2245 1420 2246
rect 1414 2241 1415 2245
rect 1419 2241 1420 2245
rect 1414 2240 1420 2241
rect 1766 2244 1772 2245
rect 1766 2240 1767 2244
rect 1771 2240 1772 2244
rect 110 2239 116 2240
rect 1766 2239 1772 2240
rect 1806 2243 1812 2244
rect 1806 2239 1807 2243
rect 1811 2239 1812 2243
rect 2110 2243 2111 2247
rect 2115 2243 2116 2247
rect 2110 2242 2116 2243
rect 2206 2247 2212 2248
rect 2206 2243 2207 2247
rect 2211 2243 2212 2247
rect 2206 2242 2212 2243
rect 2310 2247 2316 2248
rect 2310 2243 2311 2247
rect 2315 2243 2316 2247
rect 2310 2242 2316 2243
rect 2414 2247 2420 2248
rect 2414 2243 2415 2247
rect 2419 2243 2420 2247
rect 2430 2247 2431 2251
rect 2435 2250 2436 2251
rect 2559 2251 2565 2252
rect 2435 2248 2505 2250
rect 2435 2247 2436 2248
rect 2430 2246 2436 2247
rect 2559 2247 2560 2251
rect 2564 2250 2565 2251
rect 2670 2251 2676 2252
rect 2564 2248 2633 2250
rect 2564 2247 2565 2248
rect 2559 2246 2565 2247
rect 2670 2247 2671 2251
rect 2675 2250 2676 2251
rect 2814 2251 2820 2252
rect 2675 2248 2777 2250
rect 2675 2247 2676 2248
rect 2670 2246 2676 2247
rect 2814 2247 2815 2251
rect 2819 2250 2820 2251
rect 2966 2251 2972 2252
rect 2819 2248 2929 2250
rect 2819 2247 2820 2248
rect 2814 2246 2820 2247
rect 2966 2247 2967 2251
rect 2971 2250 2972 2251
rect 3438 2251 3444 2252
rect 2971 2248 3089 2250
rect 2971 2247 2972 2248
rect 2966 2246 2972 2247
rect 3338 2247 3344 2248
rect 3338 2246 3339 2247
rect 3289 2244 3339 2246
rect 2414 2242 2420 2243
rect 3338 2243 3339 2244
rect 3343 2243 3344 2247
rect 3438 2247 3439 2251
rect 3443 2247 3444 2251
rect 3438 2246 3444 2247
rect 3338 2242 3344 2243
rect 3462 2243 3468 2244
rect 1806 2238 1812 2239
rect 2038 2240 2044 2241
rect 2038 2236 2039 2240
rect 2043 2236 2044 2240
rect 2038 2235 2044 2236
rect 2134 2240 2140 2241
rect 2134 2236 2135 2240
rect 2139 2236 2140 2240
rect 2134 2235 2140 2236
rect 2238 2240 2244 2241
rect 2238 2236 2239 2240
rect 2243 2236 2244 2240
rect 2238 2235 2244 2236
rect 2342 2240 2348 2241
rect 2342 2236 2343 2240
rect 2347 2236 2348 2240
rect 2342 2235 2348 2236
rect 2462 2240 2468 2241
rect 2462 2236 2463 2240
rect 2467 2236 2468 2240
rect 2462 2235 2468 2236
rect 2590 2240 2596 2241
rect 2590 2236 2591 2240
rect 2595 2236 2596 2240
rect 2590 2235 2596 2236
rect 2734 2240 2740 2241
rect 2734 2236 2735 2240
rect 2739 2236 2740 2240
rect 2734 2235 2740 2236
rect 2886 2240 2892 2241
rect 2886 2236 2887 2240
rect 2891 2236 2892 2240
rect 2886 2235 2892 2236
rect 3046 2240 3052 2241
rect 3046 2236 3047 2240
rect 3051 2236 3052 2240
rect 3046 2235 3052 2236
rect 3214 2240 3220 2241
rect 3214 2236 3215 2240
rect 3219 2236 3220 2240
rect 3214 2235 3220 2236
rect 3366 2240 3372 2241
rect 3366 2236 3367 2240
rect 3371 2236 3372 2240
rect 3462 2239 3463 2243
rect 3467 2239 3468 2243
rect 3462 2238 3468 2239
rect 3366 2235 3372 2236
rect 2230 2231 2236 2232
rect 2230 2230 2231 2231
rect 2092 2228 2231 2230
rect 2092 2226 2094 2228
rect 2230 2227 2231 2228
rect 2235 2227 2236 2231
rect 2230 2226 2236 2227
rect 2091 2225 2097 2226
rect 2091 2221 2092 2225
rect 2096 2221 2097 2225
rect 2091 2220 2097 2221
rect 2110 2223 2116 2224
rect 2110 2219 2111 2223
rect 2115 2222 2116 2223
rect 2187 2223 2193 2224
rect 2187 2222 2188 2223
rect 2115 2220 2188 2222
rect 2115 2219 2116 2220
rect 2110 2218 2116 2219
rect 2187 2219 2188 2220
rect 2192 2219 2193 2223
rect 2187 2218 2193 2219
rect 2206 2223 2212 2224
rect 2206 2219 2207 2223
rect 2211 2222 2212 2223
rect 2291 2223 2297 2224
rect 2291 2222 2292 2223
rect 2211 2220 2292 2222
rect 2211 2219 2212 2220
rect 2206 2218 2212 2219
rect 2291 2219 2292 2220
rect 2296 2219 2297 2223
rect 2291 2218 2297 2219
rect 2310 2223 2316 2224
rect 2310 2219 2311 2223
rect 2315 2222 2316 2223
rect 2395 2223 2401 2224
rect 2395 2222 2396 2223
rect 2315 2220 2396 2222
rect 2315 2219 2316 2220
rect 2310 2218 2316 2219
rect 2395 2219 2396 2220
rect 2400 2219 2401 2223
rect 2395 2218 2401 2219
rect 2414 2223 2420 2224
rect 2414 2219 2415 2223
rect 2419 2222 2420 2223
rect 2515 2223 2521 2224
rect 2515 2222 2516 2223
rect 2419 2220 2516 2222
rect 2419 2219 2420 2220
rect 2414 2218 2420 2219
rect 2515 2219 2516 2220
rect 2520 2219 2521 2223
rect 2515 2218 2521 2219
rect 2643 2223 2649 2224
rect 2643 2219 2644 2223
rect 2648 2222 2649 2223
rect 2670 2223 2676 2224
rect 2670 2222 2671 2223
rect 2648 2220 2671 2222
rect 2648 2219 2649 2220
rect 2643 2218 2649 2219
rect 2670 2219 2671 2220
rect 2675 2219 2676 2223
rect 2670 2218 2676 2219
rect 2787 2223 2793 2224
rect 2787 2219 2788 2223
rect 2792 2222 2793 2223
rect 2814 2223 2820 2224
rect 2814 2222 2815 2223
rect 2792 2220 2815 2222
rect 2792 2219 2793 2220
rect 2787 2218 2793 2219
rect 2814 2219 2815 2220
rect 2819 2219 2820 2223
rect 2814 2218 2820 2219
rect 2939 2223 2945 2224
rect 2939 2219 2940 2223
rect 2944 2222 2945 2223
rect 2966 2223 2972 2224
rect 2966 2222 2967 2223
rect 2944 2220 2967 2222
rect 2944 2219 2945 2220
rect 2939 2218 2945 2219
rect 2966 2219 2967 2220
rect 2971 2219 2972 2223
rect 2966 2218 2972 2219
rect 3038 2223 3044 2224
rect 3038 2219 3039 2223
rect 3043 2222 3044 2223
rect 3099 2223 3105 2224
rect 3099 2222 3100 2223
rect 3043 2220 3100 2222
rect 3043 2219 3044 2220
rect 3038 2218 3044 2219
rect 3099 2219 3100 2220
rect 3104 2219 3105 2223
rect 3099 2218 3105 2219
rect 3267 2223 3273 2224
rect 3267 2219 3268 2223
rect 3272 2222 3273 2223
rect 3318 2223 3324 2224
rect 3318 2222 3319 2223
rect 3272 2220 3319 2222
rect 3272 2219 3273 2220
rect 3267 2218 3273 2219
rect 3318 2219 3319 2220
rect 3323 2219 3324 2223
rect 3318 2218 3324 2219
rect 3419 2223 3425 2224
rect 3419 2219 3420 2223
rect 3424 2222 3425 2223
rect 3430 2223 3436 2224
rect 3430 2222 3431 2223
rect 3424 2220 3431 2222
rect 3424 2219 3425 2220
rect 3419 2218 3425 2219
rect 3430 2219 3431 2220
rect 3435 2219 3436 2223
rect 3430 2218 3436 2219
rect 2430 2207 2436 2208
rect 2430 2206 2431 2207
rect 2236 2204 2431 2206
rect 2236 2202 2238 2204
rect 2430 2203 2431 2204
rect 2435 2203 2436 2207
rect 2430 2202 2436 2203
rect 2235 2201 2241 2202
rect 110 2200 116 2201
rect 1766 2200 1772 2201
rect 110 2196 111 2200
rect 115 2196 116 2200
rect 110 2195 116 2196
rect 438 2199 444 2200
rect 438 2195 439 2199
rect 443 2195 444 2199
rect 438 2194 444 2195
rect 526 2199 532 2200
rect 526 2195 527 2199
rect 531 2195 532 2199
rect 526 2194 532 2195
rect 614 2199 620 2200
rect 614 2195 615 2199
rect 619 2195 620 2199
rect 614 2194 620 2195
rect 702 2199 708 2200
rect 702 2195 703 2199
rect 707 2195 708 2199
rect 702 2194 708 2195
rect 790 2199 796 2200
rect 790 2195 791 2199
rect 795 2195 796 2199
rect 878 2199 884 2200
rect 790 2194 796 2195
rect 854 2195 860 2196
rect 854 2191 855 2195
rect 859 2194 860 2195
rect 878 2195 879 2199
rect 883 2195 884 2199
rect 878 2194 884 2195
rect 966 2199 972 2200
rect 966 2195 967 2199
rect 971 2195 972 2199
rect 966 2194 972 2195
rect 1054 2199 1060 2200
rect 1054 2195 1055 2199
rect 1059 2195 1060 2199
rect 1054 2194 1060 2195
rect 1142 2199 1148 2200
rect 1142 2195 1143 2199
rect 1147 2195 1148 2199
rect 1142 2194 1148 2195
rect 1230 2199 1236 2200
rect 1230 2195 1231 2199
rect 1235 2195 1236 2199
rect 1230 2194 1236 2195
rect 1318 2199 1324 2200
rect 1318 2195 1319 2199
rect 1323 2195 1324 2199
rect 1766 2196 1767 2200
rect 1771 2196 1772 2200
rect 2235 2197 2236 2201
rect 2240 2197 2241 2201
rect 2235 2196 2241 2197
rect 2254 2199 2260 2200
rect 1766 2195 1772 2196
rect 2254 2195 2255 2199
rect 2259 2198 2260 2199
rect 2331 2199 2337 2200
rect 2331 2198 2332 2199
rect 2259 2196 2332 2198
rect 2259 2195 2260 2196
rect 1318 2194 1324 2195
rect 2254 2194 2260 2195
rect 2331 2195 2332 2196
rect 2336 2195 2337 2199
rect 2331 2194 2337 2195
rect 2350 2199 2356 2200
rect 2350 2195 2351 2199
rect 2355 2198 2356 2199
rect 2435 2199 2441 2200
rect 2435 2198 2436 2199
rect 2355 2196 2436 2198
rect 2355 2195 2356 2196
rect 2350 2194 2356 2195
rect 2435 2195 2436 2196
rect 2440 2195 2441 2199
rect 2435 2194 2441 2195
rect 2454 2199 2460 2200
rect 2454 2195 2455 2199
rect 2459 2198 2460 2199
rect 2547 2199 2553 2200
rect 2547 2198 2548 2199
rect 2459 2196 2548 2198
rect 2459 2195 2460 2196
rect 2454 2194 2460 2195
rect 2547 2195 2548 2196
rect 2552 2195 2553 2199
rect 2547 2194 2553 2195
rect 2566 2199 2572 2200
rect 2566 2195 2567 2199
rect 2571 2198 2572 2199
rect 2659 2199 2665 2200
rect 2659 2198 2660 2199
rect 2571 2196 2660 2198
rect 2571 2195 2572 2196
rect 2566 2194 2572 2195
rect 2659 2195 2660 2196
rect 2664 2195 2665 2199
rect 2659 2194 2665 2195
rect 2771 2199 2777 2200
rect 2771 2195 2772 2199
rect 2776 2198 2777 2199
rect 2790 2199 2796 2200
rect 2776 2196 2786 2198
rect 2776 2195 2777 2196
rect 2771 2194 2777 2195
rect 859 2192 866 2194
rect 859 2191 860 2192
rect 854 2190 860 2191
rect 864 2189 866 2192
rect 1407 2191 1413 2192
rect 1407 2190 1408 2191
rect 1393 2188 1408 2190
rect 510 2187 516 2188
rect 110 2183 116 2184
rect 110 2179 111 2183
rect 115 2179 116 2183
rect 510 2183 511 2187
rect 515 2183 516 2187
rect 510 2182 516 2183
rect 598 2187 604 2188
rect 598 2183 599 2187
rect 603 2183 604 2187
rect 598 2182 604 2183
rect 686 2187 692 2188
rect 686 2183 687 2187
rect 691 2183 692 2187
rect 686 2182 692 2183
rect 774 2187 780 2188
rect 774 2183 775 2187
rect 779 2183 780 2187
rect 774 2182 780 2183
rect 950 2187 956 2188
rect 950 2183 951 2187
rect 955 2183 956 2187
rect 950 2182 956 2183
rect 1038 2187 1044 2188
rect 1038 2183 1039 2187
rect 1043 2183 1044 2187
rect 1038 2182 1044 2183
rect 1126 2187 1132 2188
rect 1126 2183 1127 2187
rect 1131 2183 1132 2187
rect 1126 2182 1132 2183
rect 1214 2187 1220 2188
rect 1214 2183 1215 2187
rect 1219 2183 1220 2187
rect 1214 2182 1220 2183
rect 1302 2187 1308 2188
rect 1302 2183 1303 2187
rect 1307 2183 1308 2187
rect 1407 2187 1408 2188
rect 1412 2187 1413 2191
rect 2784 2190 2786 2196
rect 2790 2195 2791 2199
rect 2795 2198 2796 2199
rect 2891 2199 2897 2200
rect 2891 2198 2892 2199
rect 2795 2196 2892 2198
rect 2795 2195 2796 2196
rect 2790 2194 2796 2195
rect 2891 2195 2892 2196
rect 2896 2195 2897 2199
rect 2891 2194 2897 2195
rect 2910 2199 2916 2200
rect 2910 2195 2911 2199
rect 2915 2198 2916 2199
rect 3019 2199 3025 2200
rect 3019 2198 3020 2199
rect 2915 2196 3020 2198
rect 2915 2195 2916 2196
rect 2910 2194 2916 2195
rect 3019 2195 3020 2196
rect 3024 2195 3025 2199
rect 3019 2194 3025 2195
rect 3114 2199 3120 2200
rect 3114 2195 3115 2199
rect 3119 2198 3120 2199
rect 3155 2199 3161 2200
rect 3155 2198 3156 2199
rect 3119 2196 3156 2198
rect 3119 2195 3120 2196
rect 3114 2194 3120 2195
rect 3155 2195 3156 2196
rect 3160 2195 3161 2199
rect 3155 2194 3161 2195
rect 3174 2199 3180 2200
rect 3174 2195 3175 2199
rect 3179 2198 3180 2199
rect 3299 2199 3305 2200
rect 3299 2198 3300 2199
rect 3179 2196 3300 2198
rect 3179 2195 3180 2196
rect 3174 2194 3180 2195
rect 3299 2195 3300 2196
rect 3304 2195 3305 2199
rect 3299 2194 3305 2195
rect 3419 2199 3425 2200
rect 3419 2195 3420 2199
rect 3424 2198 3425 2199
rect 3438 2199 3444 2200
rect 3438 2198 3439 2199
rect 3424 2196 3439 2198
rect 3424 2195 3425 2196
rect 3419 2194 3425 2195
rect 3438 2195 3439 2196
rect 3443 2195 3444 2199
rect 3438 2194 3444 2195
rect 2784 2188 3201 2190
rect 1407 2186 1413 2187
rect 2182 2184 2188 2185
rect 1302 2182 1308 2183
rect 1766 2183 1772 2184
rect 110 2178 116 2179
rect 438 2180 444 2181
rect 438 2176 439 2180
rect 443 2176 444 2180
rect 438 2175 444 2176
rect 526 2180 532 2181
rect 526 2176 527 2180
rect 531 2176 532 2180
rect 526 2175 532 2176
rect 614 2180 620 2181
rect 614 2176 615 2180
rect 619 2176 620 2180
rect 614 2175 620 2176
rect 702 2180 708 2181
rect 702 2176 703 2180
rect 707 2176 708 2180
rect 702 2175 708 2176
rect 790 2180 796 2181
rect 790 2176 791 2180
rect 795 2176 796 2180
rect 790 2175 796 2176
rect 878 2180 884 2181
rect 878 2176 879 2180
rect 883 2176 884 2180
rect 878 2175 884 2176
rect 966 2180 972 2181
rect 966 2176 967 2180
rect 971 2176 972 2180
rect 966 2175 972 2176
rect 1054 2180 1060 2181
rect 1054 2176 1055 2180
rect 1059 2176 1060 2180
rect 1054 2175 1060 2176
rect 1142 2180 1148 2181
rect 1142 2176 1143 2180
rect 1147 2176 1148 2180
rect 1142 2175 1148 2176
rect 1230 2180 1236 2181
rect 1230 2176 1231 2180
rect 1235 2176 1236 2180
rect 1230 2175 1236 2176
rect 1318 2180 1324 2181
rect 1318 2176 1319 2180
rect 1323 2176 1324 2180
rect 1766 2179 1767 2183
rect 1771 2179 1772 2183
rect 1766 2178 1772 2179
rect 1806 2181 1812 2182
rect 1806 2177 1807 2181
rect 1811 2177 1812 2181
rect 2182 2180 2183 2184
rect 2187 2180 2188 2184
rect 2182 2179 2188 2180
rect 2278 2184 2284 2185
rect 2278 2180 2279 2184
rect 2283 2180 2284 2184
rect 2278 2179 2284 2180
rect 2382 2184 2388 2185
rect 2382 2180 2383 2184
rect 2387 2180 2388 2184
rect 2382 2179 2388 2180
rect 2494 2184 2500 2185
rect 2494 2180 2495 2184
rect 2499 2180 2500 2184
rect 2494 2179 2500 2180
rect 2606 2184 2612 2185
rect 2606 2180 2607 2184
rect 2611 2180 2612 2184
rect 2606 2179 2612 2180
rect 2718 2184 2724 2185
rect 2718 2180 2719 2184
rect 2723 2180 2724 2184
rect 2718 2179 2724 2180
rect 2838 2184 2844 2185
rect 2838 2180 2839 2184
rect 2843 2180 2844 2184
rect 2838 2179 2844 2180
rect 2966 2184 2972 2185
rect 2966 2180 2967 2184
rect 2971 2180 2972 2184
rect 2966 2179 2972 2180
rect 3102 2184 3108 2185
rect 3102 2180 3103 2184
rect 3107 2180 3108 2184
rect 3102 2179 3108 2180
rect 1806 2176 1812 2177
rect 1318 2175 1324 2176
rect 2254 2175 2260 2176
rect 734 2171 740 2172
rect 734 2167 735 2171
rect 739 2170 740 2171
rect 2254 2171 2255 2175
rect 2259 2171 2260 2175
rect 2254 2170 2260 2171
rect 2350 2175 2356 2176
rect 2350 2171 2351 2175
rect 2355 2171 2356 2175
rect 2350 2170 2356 2171
rect 2454 2175 2460 2176
rect 2454 2171 2455 2175
rect 2459 2171 2460 2175
rect 2454 2170 2460 2171
rect 2566 2175 2572 2176
rect 2566 2171 2567 2175
rect 2571 2171 2572 2175
rect 2566 2170 2572 2171
rect 2678 2175 2684 2176
rect 2678 2171 2679 2175
rect 2683 2171 2684 2175
rect 2678 2170 2684 2171
rect 2790 2175 2796 2176
rect 2790 2171 2791 2175
rect 2795 2171 2796 2175
rect 2790 2170 2796 2171
rect 2910 2175 2916 2176
rect 2910 2171 2911 2175
rect 2915 2171 2916 2175
rect 2910 2170 2916 2171
rect 3038 2175 3044 2176
rect 3038 2171 3039 2175
rect 3043 2171 3044 2175
rect 3038 2170 3044 2171
rect 3174 2175 3180 2176
rect 3174 2171 3175 2175
rect 3179 2171 3180 2175
rect 3199 2174 3201 2188
rect 3246 2184 3252 2185
rect 3246 2180 3247 2184
rect 3251 2180 3252 2184
rect 3246 2179 3252 2180
rect 3366 2184 3372 2185
rect 3366 2180 3367 2184
rect 3371 2180 3372 2184
rect 3366 2179 3372 2180
rect 3462 2181 3468 2182
rect 3462 2177 3463 2181
rect 3467 2177 3468 2181
rect 3462 2176 3468 2177
rect 3430 2175 3436 2176
rect 3199 2172 3289 2174
rect 3174 2170 3180 2171
rect 3430 2171 3431 2175
rect 3435 2171 3436 2175
rect 3430 2170 3436 2171
rect 739 2168 934 2170
rect 739 2167 740 2168
rect 734 2166 740 2167
rect 932 2166 934 2168
rect 931 2165 937 2166
rect 2182 2165 2188 2166
rect 491 2163 497 2164
rect 491 2159 492 2163
rect 496 2162 497 2163
rect 510 2163 516 2164
rect 496 2160 506 2162
rect 496 2159 497 2160
rect 491 2158 497 2159
rect 504 2154 506 2160
rect 510 2159 511 2163
rect 515 2162 516 2163
rect 579 2163 585 2164
rect 579 2162 580 2163
rect 515 2160 580 2162
rect 515 2159 516 2160
rect 510 2158 516 2159
rect 579 2159 580 2160
rect 584 2159 585 2163
rect 579 2158 585 2159
rect 598 2163 604 2164
rect 598 2159 599 2163
rect 603 2162 604 2163
rect 667 2163 673 2164
rect 667 2162 668 2163
rect 603 2160 668 2162
rect 603 2159 604 2160
rect 598 2158 604 2159
rect 667 2159 668 2160
rect 672 2159 673 2163
rect 667 2158 673 2159
rect 686 2163 692 2164
rect 686 2159 687 2163
rect 691 2162 692 2163
rect 755 2163 761 2164
rect 755 2162 756 2163
rect 691 2160 756 2162
rect 691 2159 692 2160
rect 686 2158 692 2159
rect 755 2159 756 2160
rect 760 2159 761 2163
rect 755 2158 761 2159
rect 774 2163 780 2164
rect 774 2159 775 2163
rect 779 2162 780 2163
rect 843 2163 849 2164
rect 843 2162 844 2163
rect 779 2160 844 2162
rect 779 2159 780 2160
rect 774 2158 780 2159
rect 843 2159 844 2160
rect 848 2159 849 2163
rect 931 2161 932 2165
rect 936 2161 937 2165
rect 1806 2164 1812 2165
rect 931 2160 937 2161
rect 950 2163 956 2164
rect 843 2158 849 2159
rect 950 2159 951 2163
rect 955 2162 956 2163
rect 1019 2163 1025 2164
rect 1019 2162 1020 2163
rect 955 2160 1020 2162
rect 955 2159 956 2160
rect 950 2158 956 2159
rect 1019 2159 1020 2160
rect 1024 2159 1025 2163
rect 1019 2158 1025 2159
rect 1038 2163 1044 2164
rect 1038 2159 1039 2163
rect 1043 2162 1044 2163
rect 1107 2163 1113 2164
rect 1107 2162 1108 2163
rect 1043 2160 1108 2162
rect 1043 2159 1044 2160
rect 1038 2158 1044 2159
rect 1107 2159 1108 2160
rect 1112 2159 1113 2163
rect 1107 2158 1113 2159
rect 1126 2163 1132 2164
rect 1126 2159 1127 2163
rect 1131 2162 1132 2163
rect 1195 2163 1201 2164
rect 1195 2162 1196 2163
rect 1131 2160 1196 2162
rect 1131 2159 1132 2160
rect 1126 2158 1132 2159
rect 1195 2159 1196 2160
rect 1200 2159 1201 2163
rect 1195 2158 1201 2159
rect 1214 2163 1220 2164
rect 1214 2159 1215 2163
rect 1219 2162 1220 2163
rect 1283 2163 1289 2164
rect 1283 2162 1284 2163
rect 1219 2160 1284 2162
rect 1219 2159 1220 2160
rect 1214 2158 1220 2159
rect 1283 2159 1284 2160
rect 1288 2159 1289 2163
rect 1283 2158 1289 2159
rect 1302 2163 1308 2164
rect 1302 2159 1303 2163
rect 1307 2162 1308 2163
rect 1371 2163 1377 2164
rect 1371 2162 1372 2163
rect 1307 2160 1372 2162
rect 1307 2159 1308 2160
rect 1302 2158 1308 2159
rect 1371 2159 1372 2160
rect 1376 2159 1377 2163
rect 1806 2160 1807 2164
rect 1811 2160 1812 2164
rect 2182 2161 2183 2165
rect 2187 2161 2188 2165
rect 2182 2160 2188 2161
rect 2278 2165 2284 2166
rect 2278 2161 2279 2165
rect 2283 2161 2284 2165
rect 2278 2160 2284 2161
rect 2382 2165 2388 2166
rect 2382 2161 2383 2165
rect 2387 2161 2388 2165
rect 2382 2160 2388 2161
rect 2494 2165 2500 2166
rect 2494 2161 2495 2165
rect 2499 2161 2500 2165
rect 2494 2160 2500 2161
rect 2606 2165 2612 2166
rect 2606 2161 2607 2165
rect 2611 2161 2612 2165
rect 2606 2160 2612 2161
rect 2718 2165 2724 2166
rect 2718 2161 2719 2165
rect 2723 2161 2724 2165
rect 2718 2160 2724 2161
rect 2838 2165 2844 2166
rect 2838 2161 2839 2165
rect 2843 2161 2844 2165
rect 2838 2160 2844 2161
rect 2966 2165 2972 2166
rect 2966 2161 2967 2165
rect 2971 2161 2972 2165
rect 2966 2160 2972 2161
rect 3102 2165 3108 2166
rect 3102 2161 3103 2165
rect 3107 2161 3108 2165
rect 3102 2160 3108 2161
rect 3246 2165 3252 2166
rect 3246 2161 3247 2165
rect 3251 2161 3252 2165
rect 3246 2160 3252 2161
rect 3366 2165 3372 2166
rect 3366 2161 3367 2165
rect 3371 2161 3372 2165
rect 3366 2160 3372 2161
rect 3462 2164 3468 2165
rect 3462 2160 3463 2164
rect 3467 2160 3468 2164
rect 1806 2159 1812 2160
rect 3462 2159 3468 2160
rect 1371 2158 1377 2159
rect 598 2155 604 2156
rect 598 2154 599 2155
rect 504 2152 599 2154
rect 598 2151 599 2152
rect 603 2151 604 2155
rect 598 2150 604 2151
rect 326 2135 332 2136
rect 326 2131 327 2135
rect 331 2134 332 2135
rect 355 2135 361 2136
rect 355 2134 356 2135
rect 331 2132 356 2134
rect 331 2131 332 2132
rect 326 2130 332 2131
rect 355 2131 356 2132
rect 360 2131 361 2135
rect 355 2130 361 2131
rect 374 2135 380 2136
rect 374 2131 375 2135
rect 379 2134 380 2135
rect 459 2135 465 2136
rect 459 2134 460 2135
rect 379 2132 460 2134
rect 379 2131 380 2132
rect 374 2130 380 2131
rect 459 2131 460 2132
rect 464 2131 465 2135
rect 459 2130 465 2131
rect 478 2135 484 2136
rect 478 2131 479 2135
rect 483 2134 484 2135
rect 571 2135 577 2136
rect 571 2134 572 2135
rect 483 2132 572 2134
rect 483 2131 484 2132
rect 478 2130 484 2131
rect 571 2131 572 2132
rect 576 2131 577 2135
rect 571 2130 577 2131
rect 590 2135 596 2136
rect 590 2131 591 2135
rect 595 2134 596 2135
rect 683 2135 689 2136
rect 683 2134 684 2135
rect 595 2132 684 2134
rect 595 2131 596 2132
rect 590 2130 596 2131
rect 683 2131 684 2132
rect 688 2131 689 2135
rect 683 2130 689 2131
rect 795 2135 801 2136
rect 795 2131 796 2135
rect 800 2134 801 2135
rect 822 2135 828 2136
rect 822 2134 823 2135
rect 800 2132 823 2134
rect 800 2131 801 2132
rect 795 2130 801 2131
rect 822 2131 823 2132
rect 827 2131 828 2135
rect 822 2130 828 2131
rect 915 2135 921 2136
rect 915 2131 916 2135
rect 920 2134 921 2135
rect 943 2135 949 2136
rect 943 2134 944 2135
rect 920 2132 944 2134
rect 920 2131 921 2132
rect 915 2130 921 2131
rect 943 2131 944 2132
rect 948 2131 949 2135
rect 943 2130 949 2131
rect 1006 2135 1012 2136
rect 1006 2131 1007 2135
rect 1011 2134 1012 2135
rect 1035 2135 1041 2136
rect 1035 2134 1036 2135
rect 1011 2132 1036 2134
rect 1011 2131 1012 2132
rect 1006 2130 1012 2131
rect 1035 2131 1036 2132
rect 1040 2131 1041 2135
rect 1035 2130 1041 2131
rect 302 2120 308 2121
rect 110 2117 116 2118
rect 110 2113 111 2117
rect 115 2113 116 2117
rect 302 2116 303 2120
rect 307 2116 308 2120
rect 302 2115 308 2116
rect 406 2120 412 2121
rect 406 2116 407 2120
rect 411 2116 412 2120
rect 406 2115 412 2116
rect 518 2120 524 2121
rect 518 2116 519 2120
rect 523 2116 524 2120
rect 518 2115 524 2116
rect 630 2120 636 2121
rect 630 2116 631 2120
rect 635 2116 636 2120
rect 630 2115 636 2116
rect 742 2120 748 2121
rect 742 2116 743 2120
rect 747 2116 748 2120
rect 742 2115 748 2116
rect 862 2120 868 2121
rect 862 2116 863 2120
rect 867 2116 868 2120
rect 862 2115 868 2116
rect 982 2120 988 2121
rect 982 2116 983 2120
rect 987 2116 988 2120
rect 982 2115 988 2116
rect 1766 2117 1772 2118
rect 110 2112 116 2113
rect 1766 2113 1767 2117
rect 1771 2113 1772 2117
rect 1766 2112 1772 2113
rect 1806 2112 1812 2113
rect 3462 2112 3468 2113
rect 374 2111 380 2112
rect 374 2107 375 2111
rect 379 2107 380 2111
rect 374 2106 380 2107
rect 478 2111 484 2112
rect 478 2107 479 2111
rect 483 2107 484 2111
rect 478 2106 484 2107
rect 590 2111 596 2112
rect 590 2107 591 2111
rect 595 2107 596 2111
rect 590 2106 596 2107
rect 598 2111 604 2112
rect 598 2107 599 2111
rect 603 2110 604 2111
rect 718 2111 724 2112
rect 603 2108 673 2110
rect 603 2107 604 2108
rect 598 2106 604 2107
rect 718 2107 719 2111
rect 723 2110 724 2111
rect 822 2111 828 2112
rect 723 2108 785 2110
rect 723 2107 724 2108
rect 718 2106 724 2107
rect 822 2107 823 2111
rect 827 2110 828 2111
rect 943 2111 949 2112
rect 827 2108 905 2110
rect 827 2107 828 2108
rect 822 2106 828 2107
rect 943 2107 944 2111
rect 948 2110 949 2111
rect 948 2108 1025 2110
rect 1806 2108 1807 2112
rect 1811 2108 1812 2112
rect 948 2107 949 2108
rect 1806 2107 1812 2108
rect 2134 2111 2140 2112
rect 2134 2107 2135 2111
rect 2139 2107 2140 2111
rect 943 2106 949 2107
rect 2134 2106 2140 2107
rect 2254 2111 2260 2112
rect 2254 2107 2255 2111
rect 2259 2107 2260 2111
rect 2254 2106 2260 2107
rect 2382 2111 2388 2112
rect 2382 2107 2383 2111
rect 2387 2107 2388 2111
rect 2382 2106 2388 2107
rect 2518 2111 2524 2112
rect 2518 2107 2519 2111
rect 2523 2107 2524 2111
rect 2518 2106 2524 2107
rect 2654 2111 2660 2112
rect 2654 2107 2655 2111
rect 2659 2107 2660 2111
rect 2654 2106 2660 2107
rect 2782 2111 2788 2112
rect 2782 2107 2783 2111
rect 2787 2107 2788 2111
rect 2782 2106 2788 2107
rect 2910 2111 2916 2112
rect 2910 2107 2911 2111
rect 2915 2107 2916 2111
rect 2910 2106 2916 2107
rect 3030 2111 3036 2112
rect 3030 2107 3031 2111
rect 3035 2107 3036 2111
rect 3030 2106 3036 2107
rect 3150 2111 3156 2112
rect 3150 2107 3151 2111
rect 3155 2107 3156 2111
rect 3150 2106 3156 2107
rect 3270 2111 3276 2112
rect 3270 2107 3271 2111
rect 3275 2107 3276 2111
rect 3270 2106 3276 2107
rect 3366 2111 3372 2112
rect 3366 2107 3367 2111
rect 3371 2107 3372 2111
rect 3462 2108 3463 2112
rect 3467 2108 3468 2112
rect 3462 2107 3468 2108
rect 3366 2106 3372 2107
rect 2214 2103 2220 2104
rect 302 2101 308 2102
rect 110 2100 116 2101
rect 110 2096 111 2100
rect 115 2096 116 2100
rect 302 2097 303 2101
rect 307 2097 308 2101
rect 302 2096 308 2097
rect 406 2101 412 2102
rect 406 2097 407 2101
rect 411 2097 412 2101
rect 406 2096 412 2097
rect 518 2101 524 2102
rect 518 2097 519 2101
rect 523 2097 524 2101
rect 518 2096 524 2097
rect 630 2101 636 2102
rect 630 2097 631 2101
rect 635 2097 636 2101
rect 630 2096 636 2097
rect 742 2101 748 2102
rect 742 2097 743 2101
rect 747 2097 748 2101
rect 742 2096 748 2097
rect 862 2101 868 2102
rect 862 2097 863 2101
rect 867 2097 868 2101
rect 862 2096 868 2097
rect 982 2101 988 2102
rect 982 2097 983 2101
rect 987 2097 988 2101
rect 982 2096 988 2097
rect 1766 2100 1772 2101
rect 1766 2096 1767 2100
rect 1771 2096 1772 2100
rect 2206 2099 2212 2100
rect 110 2095 116 2096
rect 1766 2095 1772 2096
rect 1806 2095 1812 2096
rect 1806 2091 1807 2095
rect 1811 2091 1812 2095
rect 2206 2095 2207 2099
rect 2211 2095 2212 2099
rect 2214 2099 2215 2103
rect 2219 2102 2220 2103
rect 2334 2103 2340 2104
rect 2219 2100 2297 2102
rect 2219 2099 2220 2100
rect 2214 2098 2220 2099
rect 2334 2099 2335 2103
rect 2339 2102 2340 2103
rect 2462 2103 2468 2104
rect 2339 2100 2425 2102
rect 2339 2099 2340 2100
rect 2334 2098 2340 2099
rect 2462 2099 2463 2103
rect 2467 2102 2468 2103
rect 2598 2103 2604 2104
rect 2467 2100 2561 2102
rect 2467 2099 2468 2100
rect 2462 2098 2468 2099
rect 2598 2099 2599 2103
rect 2603 2102 2604 2103
rect 3114 2103 3120 2104
rect 3114 2102 3115 2103
rect 2603 2100 2697 2102
rect 3105 2100 3115 2102
rect 2603 2099 2604 2100
rect 2598 2098 2604 2099
rect 2854 2099 2860 2100
rect 2206 2094 2212 2095
rect 2854 2095 2855 2099
rect 2859 2095 2860 2099
rect 2854 2094 2860 2095
rect 2982 2099 2988 2100
rect 2982 2095 2983 2099
rect 2987 2095 2988 2099
rect 3114 2099 3115 2100
rect 3119 2099 3120 2103
rect 3114 2098 3120 2099
rect 3122 2103 3128 2104
rect 3122 2099 3123 2103
rect 3127 2102 3128 2103
rect 3230 2103 3236 2104
rect 3127 2100 3193 2102
rect 3127 2099 3128 2100
rect 3122 2098 3128 2099
rect 3230 2099 3231 2103
rect 3235 2102 3236 2103
rect 3358 2103 3364 2104
rect 3235 2100 3313 2102
rect 3235 2099 3236 2100
rect 3230 2098 3236 2099
rect 3358 2099 3359 2103
rect 3363 2102 3364 2103
rect 3363 2100 3409 2102
rect 3363 2099 3364 2100
rect 3358 2098 3364 2099
rect 2982 2094 2988 2095
rect 3462 2095 3468 2096
rect 1806 2090 1812 2091
rect 2134 2092 2140 2093
rect 2134 2088 2135 2092
rect 2139 2088 2140 2092
rect 2134 2087 2140 2088
rect 2254 2092 2260 2093
rect 2254 2088 2255 2092
rect 2259 2088 2260 2092
rect 2254 2087 2260 2088
rect 2382 2092 2388 2093
rect 2382 2088 2383 2092
rect 2387 2088 2388 2092
rect 2382 2087 2388 2088
rect 2518 2092 2524 2093
rect 2518 2088 2519 2092
rect 2523 2088 2524 2092
rect 2518 2087 2524 2088
rect 2654 2092 2660 2093
rect 2654 2088 2655 2092
rect 2659 2088 2660 2092
rect 2654 2087 2660 2088
rect 2782 2092 2788 2093
rect 2782 2088 2783 2092
rect 2787 2088 2788 2092
rect 2782 2087 2788 2088
rect 2910 2092 2916 2093
rect 2910 2088 2911 2092
rect 2915 2088 2916 2092
rect 2910 2087 2916 2088
rect 3030 2092 3036 2093
rect 3030 2088 3031 2092
rect 3035 2088 3036 2092
rect 3030 2087 3036 2088
rect 3150 2092 3156 2093
rect 3150 2088 3151 2092
rect 3155 2088 3156 2092
rect 3150 2087 3156 2088
rect 3270 2092 3276 2093
rect 3270 2088 3271 2092
rect 3275 2088 3276 2092
rect 3270 2087 3276 2088
rect 3366 2092 3372 2093
rect 3366 2088 3367 2092
rect 3371 2088 3372 2092
rect 3462 2091 3463 2095
rect 3467 2091 3468 2095
rect 3462 2090 3468 2091
rect 3366 2087 3372 2088
rect 3122 2083 3128 2084
rect 3122 2082 3123 2083
rect 2836 2080 3123 2082
rect 2836 2078 2838 2080
rect 3122 2079 3123 2080
rect 3127 2079 3128 2083
rect 3122 2078 3128 2079
rect 2835 2077 2841 2078
rect 2187 2075 2193 2076
rect 2187 2071 2188 2075
rect 2192 2074 2193 2075
rect 2214 2075 2220 2076
rect 2214 2074 2215 2075
rect 2192 2072 2215 2074
rect 2192 2071 2193 2072
rect 2187 2070 2193 2071
rect 2214 2071 2215 2072
rect 2219 2071 2220 2075
rect 2214 2070 2220 2071
rect 2307 2075 2313 2076
rect 2307 2071 2308 2075
rect 2312 2074 2313 2075
rect 2334 2075 2340 2076
rect 2334 2074 2335 2075
rect 2312 2072 2335 2074
rect 2312 2071 2313 2072
rect 2307 2070 2313 2071
rect 2334 2071 2335 2072
rect 2339 2071 2340 2075
rect 2334 2070 2340 2071
rect 2435 2075 2441 2076
rect 2435 2071 2436 2075
rect 2440 2074 2441 2075
rect 2462 2075 2468 2076
rect 2462 2074 2463 2075
rect 2440 2072 2463 2074
rect 2440 2071 2441 2072
rect 2435 2070 2441 2071
rect 2462 2071 2463 2072
rect 2467 2071 2468 2075
rect 2462 2070 2468 2071
rect 2571 2075 2577 2076
rect 2571 2071 2572 2075
rect 2576 2074 2577 2075
rect 2598 2075 2604 2076
rect 2598 2074 2599 2075
rect 2576 2072 2599 2074
rect 2576 2071 2577 2072
rect 2571 2070 2577 2071
rect 2598 2071 2599 2072
rect 2603 2071 2604 2075
rect 2598 2070 2604 2071
rect 2678 2075 2684 2076
rect 2678 2071 2679 2075
rect 2683 2074 2684 2075
rect 2707 2075 2713 2076
rect 2707 2074 2708 2075
rect 2683 2072 2708 2074
rect 2683 2071 2684 2072
rect 2678 2070 2684 2071
rect 2707 2071 2708 2072
rect 2712 2071 2713 2075
rect 2835 2073 2836 2077
rect 2840 2073 2841 2077
rect 2835 2072 2841 2073
rect 2854 2075 2860 2076
rect 2707 2070 2713 2071
rect 2854 2071 2855 2075
rect 2859 2074 2860 2075
rect 2963 2075 2969 2076
rect 2963 2074 2964 2075
rect 2859 2072 2964 2074
rect 2859 2071 2860 2072
rect 2854 2070 2860 2071
rect 2963 2071 2964 2072
rect 2968 2071 2969 2075
rect 2963 2070 2969 2071
rect 2982 2075 2988 2076
rect 2982 2071 2983 2075
rect 2987 2074 2988 2075
rect 3083 2075 3089 2076
rect 3083 2074 3084 2075
rect 2987 2072 3084 2074
rect 2987 2071 2988 2072
rect 2982 2070 2988 2071
rect 3083 2071 3084 2072
rect 3088 2071 3089 2075
rect 3083 2070 3089 2071
rect 3203 2075 3209 2076
rect 3203 2071 3204 2075
rect 3208 2074 3209 2075
rect 3230 2075 3236 2076
rect 3230 2074 3231 2075
rect 3208 2072 3231 2074
rect 3208 2071 3209 2072
rect 3203 2070 3209 2071
rect 3230 2071 3231 2072
rect 3235 2071 3236 2075
rect 3230 2070 3236 2071
rect 3323 2075 3332 2076
rect 3323 2071 3324 2075
rect 3331 2071 3332 2075
rect 3323 2070 3332 2071
rect 3338 2075 3344 2076
rect 3338 2071 3339 2075
rect 3343 2074 3344 2075
rect 3419 2075 3425 2076
rect 3419 2074 3420 2075
rect 3343 2072 3420 2074
rect 3343 2071 3344 2072
rect 3338 2070 3344 2071
rect 3419 2071 3420 2072
rect 3424 2071 3425 2075
rect 3419 2070 3425 2071
rect 110 2056 116 2057
rect 1766 2056 1772 2057
rect 110 2052 111 2056
rect 115 2052 116 2056
rect 110 2051 116 2052
rect 254 2055 260 2056
rect 254 2051 255 2055
rect 259 2051 260 2055
rect 254 2050 260 2051
rect 374 2055 380 2056
rect 374 2051 375 2055
rect 379 2051 380 2055
rect 374 2050 380 2051
rect 494 2055 500 2056
rect 494 2051 495 2055
rect 499 2051 500 2055
rect 494 2050 500 2051
rect 614 2055 620 2056
rect 614 2051 615 2055
rect 619 2051 620 2055
rect 614 2050 620 2051
rect 726 2055 732 2056
rect 726 2051 727 2055
rect 731 2051 732 2055
rect 726 2050 732 2051
rect 830 2055 836 2056
rect 830 2051 831 2055
rect 835 2051 836 2055
rect 830 2050 836 2051
rect 934 2055 940 2056
rect 934 2051 935 2055
rect 939 2051 940 2055
rect 934 2050 940 2051
rect 1038 2055 1044 2056
rect 1038 2051 1039 2055
rect 1043 2051 1044 2055
rect 1038 2050 1044 2051
rect 1142 2055 1148 2056
rect 1142 2051 1143 2055
rect 1147 2051 1148 2055
rect 1142 2050 1148 2051
rect 1254 2055 1260 2056
rect 1254 2051 1255 2055
rect 1259 2051 1260 2055
rect 1766 2052 1767 2056
rect 1771 2052 1772 2056
rect 1766 2051 1772 2052
rect 2206 2055 2212 2056
rect 2206 2051 2207 2055
rect 2211 2054 2212 2055
rect 2299 2055 2305 2056
rect 2299 2054 2300 2055
rect 2211 2052 2300 2054
rect 2211 2051 2212 2052
rect 1254 2050 1260 2051
rect 2206 2050 2212 2051
rect 2299 2051 2300 2052
rect 2304 2051 2305 2055
rect 2299 2050 2305 2051
rect 2318 2055 2324 2056
rect 2318 2051 2319 2055
rect 2323 2054 2324 2055
rect 2467 2055 2473 2056
rect 2467 2054 2468 2055
rect 2323 2052 2468 2054
rect 2323 2051 2324 2052
rect 2318 2050 2324 2051
rect 2467 2051 2468 2052
rect 2472 2051 2473 2055
rect 2467 2050 2473 2051
rect 2486 2055 2492 2056
rect 2486 2051 2487 2055
rect 2491 2054 2492 2055
rect 2627 2055 2633 2056
rect 2627 2054 2628 2055
rect 2491 2052 2628 2054
rect 2491 2051 2492 2052
rect 2486 2050 2492 2051
rect 2627 2051 2628 2052
rect 2632 2051 2633 2055
rect 2627 2050 2633 2051
rect 2779 2055 2785 2056
rect 2779 2051 2780 2055
rect 2784 2054 2785 2055
rect 2798 2055 2804 2056
rect 2784 2052 2794 2054
rect 2784 2051 2785 2052
rect 2779 2050 2785 2051
rect 326 2047 332 2048
rect 326 2043 327 2047
rect 331 2043 332 2047
rect 326 2042 332 2043
rect 334 2047 340 2048
rect 334 2043 335 2047
rect 339 2046 340 2047
rect 454 2047 460 2048
rect 339 2044 417 2046
rect 339 2043 340 2044
rect 334 2042 340 2043
rect 454 2043 455 2047
rect 459 2046 460 2047
rect 1006 2047 1012 2048
rect 459 2044 537 2046
rect 459 2043 460 2044
rect 454 2042 460 2043
rect 686 2043 692 2044
rect 110 2039 116 2040
rect 110 2035 111 2039
rect 115 2035 116 2039
rect 686 2039 687 2043
rect 691 2039 692 2043
rect 686 2038 692 2039
rect 798 2043 804 2044
rect 798 2039 799 2043
rect 803 2039 804 2043
rect 798 2038 804 2039
rect 902 2043 908 2044
rect 902 2039 903 2043
rect 907 2039 908 2043
rect 1006 2043 1007 2047
rect 1011 2043 1012 2047
rect 1006 2042 1012 2043
rect 1014 2047 1020 2048
rect 1014 2043 1015 2047
rect 1019 2046 1020 2047
rect 1118 2047 1124 2048
rect 1019 2044 1081 2046
rect 1019 2043 1020 2044
rect 1014 2042 1020 2043
rect 1118 2043 1119 2047
rect 1123 2046 1124 2047
rect 1222 2047 1228 2048
rect 1123 2044 1185 2046
rect 1123 2043 1124 2044
rect 1118 2042 1124 2043
rect 1222 2043 1223 2047
rect 1227 2046 1228 2047
rect 2792 2046 2794 2052
rect 2798 2051 2799 2055
rect 2803 2054 2804 2055
rect 2923 2055 2929 2056
rect 2923 2054 2924 2055
rect 2803 2052 2924 2054
rect 2803 2051 2804 2052
rect 2798 2050 2804 2051
rect 2923 2051 2924 2052
rect 2928 2051 2929 2055
rect 2923 2050 2929 2051
rect 2942 2055 2948 2056
rect 2942 2051 2943 2055
rect 2947 2054 2948 2055
rect 3059 2055 3065 2056
rect 3059 2054 3060 2055
rect 2947 2052 3060 2054
rect 2947 2051 2948 2052
rect 2942 2050 2948 2051
rect 3059 2051 3060 2052
rect 3064 2051 3065 2055
rect 3059 2050 3065 2051
rect 3078 2055 3084 2056
rect 3078 2051 3079 2055
rect 3083 2054 3084 2055
rect 3187 2055 3193 2056
rect 3187 2054 3188 2055
rect 3083 2052 3188 2054
rect 3083 2051 3084 2052
rect 3078 2050 3084 2051
rect 3187 2051 3188 2052
rect 3192 2051 3193 2055
rect 3187 2050 3193 2051
rect 3206 2055 3212 2056
rect 3206 2051 3207 2055
rect 3211 2054 3212 2055
rect 3315 2055 3321 2056
rect 3315 2054 3316 2055
rect 3211 2052 3316 2054
rect 3211 2051 3212 2052
rect 3206 2050 3212 2051
rect 3315 2051 3316 2052
rect 3320 2051 3321 2055
rect 3315 2050 3321 2051
rect 3419 2055 3425 2056
rect 3419 2051 3420 2055
rect 3424 2054 3425 2055
rect 3430 2055 3436 2056
rect 3430 2054 3431 2055
rect 3424 2052 3431 2054
rect 3424 2051 3425 2052
rect 3419 2050 3425 2051
rect 3430 2051 3431 2052
rect 3435 2051 3436 2055
rect 3430 2050 3436 2051
rect 3110 2047 3116 2048
rect 3110 2046 3111 2047
rect 1227 2044 1297 2046
rect 2792 2044 3111 2046
rect 1227 2043 1228 2044
rect 1222 2042 1228 2043
rect 3110 2043 3111 2044
rect 3115 2043 3116 2047
rect 3110 2042 3116 2043
rect 2246 2040 2252 2041
rect 902 2038 908 2039
rect 1766 2039 1772 2040
rect 110 2034 116 2035
rect 254 2036 260 2037
rect 254 2032 255 2036
rect 259 2032 260 2036
rect 254 2031 260 2032
rect 374 2036 380 2037
rect 374 2032 375 2036
rect 379 2032 380 2036
rect 374 2031 380 2032
rect 494 2036 500 2037
rect 494 2032 495 2036
rect 499 2032 500 2036
rect 494 2031 500 2032
rect 614 2036 620 2037
rect 614 2032 615 2036
rect 619 2032 620 2036
rect 614 2031 620 2032
rect 726 2036 732 2037
rect 726 2032 727 2036
rect 731 2032 732 2036
rect 726 2031 732 2032
rect 830 2036 836 2037
rect 830 2032 831 2036
rect 835 2032 836 2036
rect 830 2031 836 2032
rect 934 2036 940 2037
rect 934 2032 935 2036
rect 939 2032 940 2036
rect 934 2031 940 2032
rect 1038 2036 1044 2037
rect 1038 2032 1039 2036
rect 1043 2032 1044 2036
rect 1038 2031 1044 2032
rect 1142 2036 1148 2037
rect 1142 2032 1143 2036
rect 1147 2032 1148 2036
rect 1142 2031 1148 2032
rect 1254 2036 1260 2037
rect 1254 2032 1255 2036
rect 1259 2032 1260 2036
rect 1766 2035 1767 2039
rect 1771 2035 1772 2039
rect 1766 2034 1772 2035
rect 1806 2037 1812 2038
rect 1806 2033 1807 2037
rect 1811 2033 1812 2037
rect 2246 2036 2247 2040
rect 2251 2036 2252 2040
rect 2246 2035 2252 2036
rect 2414 2040 2420 2041
rect 2414 2036 2415 2040
rect 2419 2036 2420 2040
rect 2414 2035 2420 2036
rect 2574 2040 2580 2041
rect 2574 2036 2575 2040
rect 2579 2036 2580 2040
rect 2574 2035 2580 2036
rect 2726 2040 2732 2041
rect 2726 2036 2727 2040
rect 2731 2036 2732 2040
rect 2726 2035 2732 2036
rect 2870 2040 2876 2041
rect 2870 2036 2871 2040
rect 2875 2036 2876 2040
rect 2870 2035 2876 2036
rect 3006 2040 3012 2041
rect 3006 2036 3007 2040
rect 3011 2036 3012 2040
rect 3006 2035 3012 2036
rect 3134 2040 3140 2041
rect 3134 2036 3135 2040
rect 3139 2036 3140 2040
rect 3134 2035 3140 2036
rect 3262 2040 3268 2041
rect 3262 2036 3263 2040
rect 3267 2036 3268 2040
rect 3262 2035 3268 2036
rect 3366 2040 3372 2041
rect 3366 2036 3367 2040
rect 3371 2036 3372 2040
rect 3366 2035 3372 2036
rect 3462 2037 3468 2038
rect 1806 2032 1812 2033
rect 3462 2033 3463 2037
rect 3467 2033 3468 2037
rect 3462 2032 3468 2033
rect 1254 2031 1260 2032
rect 2318 2031 2324 2032
rect 718 2027 724 2028
rect 718 2026 719 2027
rect 668 2024 719 2026
rect 668 2022 670 2024
rect 718 2023 719 2024
rect 723 2023 724 2027
rect 1014 2027 1020 2028
rect 1014 2026 1015 2027
rect 718 2022 724 2023
rect 884 2024 1015 2026
rect 884 2022 886 2024
rect 1014 2023 1015 2024
rect 1019 2023 1020 2027
rect 2318 2027 2319 2031
rect 2323 2027 2324 2031
rect 2318 2026 2324 2027
rect 2486 2031 2492 2032
rect 2486 2027 2487 2031
rect 2491 2027 2492 2031
rect 2486 2026 2492 2027
rect 2526 2031 2532 2032
rect 2526 2027 2527 2031
rect 2531 2030 2532 2031
rect 2798 2031 2804 2032
rect 2531 2028 2617 2030
rect 2531 2027 2532 2028
rect 2526 2026 2532 2027
rect 2798 2027 2799 2031
rect 2803 2027 2804 2031
rect 2798 2026 2804 2027
rect 2942 2031 2948 2032
rect 2942 2027 2943 2031
rect 2947 2027 2948 2031
rect 2942 2026 2948 2027
rect 3078 2031 3084 2032
rect 3078 2027 3079 2031
rect 3083 2027 3084 2031
rect 3078 2026 3084 2027
rect 3206 2031 3212 2032
rect 3206 2027 3207 2031
rect 3211 2027 3212 2031
rect 3206 2026 3212 2027
rect 3326 2031 3332 2032
rect 3326 2027 3327 2031
rect 3331 2027 3332 2031
rect 3326 2026 3332 2027
rect 3438 2031 3444 2032
rect 3438 2027 3439 2031
rect 3443 2027 3444 2031
rect 3438 2026 3444 2027
rect 1014 2022 1020 2023
rect 667 2021 673 2022
rect 307 2019 313 2020
rect 307 2015 308 2019
rect 312 2018 313 2019
rect 334 2019 340 2020
rect 334 2018 335 2019
rect 312 2016 335 2018
rect 312 2015 313 2016
rect 307 2014 313 2015
rect 334 2015 335 2016
rect 339 2015 340 2019
rect 334 2014 340 2015
rect 427 2019 433 2020
rect 427 2015 428 2019
rect 432 2018 433 2019
rect 454 2019 460 2020
rect 454 2018 455 2019
rect 432 2016 455 2018
rect 432 2015 433 2016
rect 427 2014 433 2015
rect 454 2015 455 2016
rect 459 2015 460 2019
rect 454 2014 460 2015
rect 547 2019 556 2020
rect 547 2015 548 2019
rect 555 2015 556 2019
rect 667 2017 668 2021
rect 672 2017 673 2021
rect 883 2021 889 2022
rect 2246 2021 2252 2022
rect 667 2016 673 2017
rect 686 2019 692 2020
rect 547 2014 556 2015
rect 686 2015 687 2019
rect 691 2018 692 2019
rect 779 2019 785 2020
rect 779 2018 780 2019
rect 691 2016 780 2018
rect 691 2015 692 2016
rect 686 2014 692 2015
rect 779 2015 780 2016
rect 784 2015 785 2019
rect 883 2017 884 2021
rect 888 2017 889 2021
rect 1806 2020 1812 2021
rect 883 2016 889 2017
rect 902 2019 908 2020
rect 779 2014 785 2015
rect 902 2015 903 2019
rect 907 2018 908 2019
rect 987 2019 993 2020
rect 987 2018 988 2019
rect 907 2016 988 2018
rect 907 2015 908 2016
rect 902 2014 908 2015
rect 987 2015 988 2016
rect 992 2015 993 2019
rect 987 2014 993 2015
rect 1091 2019 1097 2020
rect 1091 2015 1092 2019
rect 1096 2018 1097 2019
rect 1118 2019 1124 2020
rect 1118 2018 1119 2019
rect 1096 2016 1119 2018
rect 1096 2015 1097 2016
rect 1091 2014 1097 2015
rect 1118 2015 1119 2016
rect 1123 2015 1124 2019
rect 1118 2014 1124 2015
rect 1195 2019 1201 2020
rect 1195 2015 1196 2019
rect 1200 2018 1201 2019
rect 1222 2019 1228 2020
rect 1222 2018 1223 2019
rect 1200 2016 1223 2018
rect 1200 2015 1201 2016
rect 1195 2014 1201 2015
rect 1222 2015 1223 2016
rect 1227 2015 1228 2019
rect 1222 2014 1228 2015
rect 1247 2019 1253 2020
rect 1247 2015 1248 2019
rect 1252 2018 1253 2019
rect 1307 2019 1313 2020
rect 1307 2018 1308 2019
rect 1252 2016 1308 2018
rect 1252 2015 1253 2016
rect 1247 2014 1253 2015
rect 1307 2015 1308 2016
rect 1312 2015 1313 2019
rect 1806 2016 1807 2020
rect 1811 2016 1812 2020
rect 2246 2017 2247 2021
rect 2251 2017 2252 2021
rect 2246 2016 2252 2017
rect 2414 2021 2420 2022
rect 2414 2017 2415 2021
rect 2419 2017 2420 2021
rect 2414 2016 2420 2017
rect 2574 2021 2580 2022
rect 2574 2017 2575 2021
rect 2579 2017 2580 2021
rect 2574 2016 2580 2017
rect 2726 2021 2732 2022
rect 2726 2017 2727 2021
rect 2731 2017 2732 2021
rect 2726 2016 2732 2017
rect 2870 2021 2876 2022
rect 2870 2017 2871 2021
rect 2875 2017 2876 2021
rect 2870 2016 2876 2017
rect 3006 2021 3012 2022
rect 3006 2017 3007 2021
rect 3011 2017 3012 2021
rect 3006 2016 3012 2017
rect 3134 2021 3140 2022
rect 3134 2017 3135 2021
rect 3139 2017 3140 2021
rect 3134 2016 3140 2017
rect 3262 2021 3268 2022
rect 3262 2017 3263 2021
rect 3267 2017 3268 2021
rect 3262 2016 3268 2017
rect 3366 2021 3372 2022
rect 3366 2017 3367 2021
rect 3371 2017 3372 2021
rect 3366 2016 3372 2017
rect 3462 2020 3468 2021
rect 3462 2016 3463 2020
rect 3467 2016 3468 2020
rect 1806 2015 1812 2016
rect 3462 2015 3468 2016
rect 1307 2014 1313 2015
rect 411 2007 417 2008
rect 411 2003 412 2007
rect 416 2006 417 2007
rect 430 2007 436 2008
rect 416 2004 426 2006
rect 416 2003 417 2004
rect 411 2002 417 2003
rect 424 1998 426 2004
rect 430 2003 431 2007
rect 435 2006 436 2007
rect 539 2007 545 2008
rect 539 2006 540 2007
rect 435 2004 540 2006
rect 435 2003 436 2004
rect 430 2002 436 2003
rect 539 2003 540 2004
rect 544 2003 545 2007
rect 539 2002 545 2003
rect 675 2007 681 2008
rect 675 2003 676 2007
rect 680 2006 681 2007
rect 702 2007 708 2008
rect 702 2006 703 2007
rect 680 2004 703 2006
rect 680 2003 681 2004
rect 675 2002 681 2003
rect 702 2003 703 2004
rect 707 2003 708 2007
rect 702 2002 708 2003
rect 798 2007 804 2008
rect 798 2003 799 2007
rect 803 2006 804 2007
rect 811 2007 817 2008
rect 811 2006 812 2007
rect 803 2004 812 2006
rect 803 2003 804 2004
rect 798 2002 804 2003
rect 811 2003 812 2004
rect 816 2003 817 2007
rect 811 2002 817 2003
rect 871 2007 877 2008
rect 871 2003 872 2007
rect 876 2006 877 2007
rect 947 2007 953 2008
rect 947 2006 948 2007
rect 876 2004 948 2006
rect 876 2003 877 2004
rect 871 2002 877 2003
rect 947 2003 948 2004
rect 952 2003 953 2007
rect 947 2002 953 2003
rect 1075 2007 1081 2008
rect 1075 2003 1076 2007
rect 1080 2006 1081 2007
rect 1094 2007 1100 2008
rect 1080 2004 1090 2006
rect 1080 2003 1081 2004
rect 1075 2002 1081 2003
rect 1088 1998 1090 2004
rect 1094 2003 1095 2007
rect 1099 2006 1100 2007
rect 1203 2007 1209 2008
rect 1203 2006 1204 2007
rect 1099 2004 1204 2006
rect 1099 2003 1100 2004
rect 1094 2002 1100 2003
rect 1203 2003 1204 2004
rect 1208 2003 1209 2007
rect 1203 2002 1209 2003
rect 1323 2007 1329 2008
rect 1323 2003 1324 2007
rect 1328 2006 1329 2007
rect 1350 2007 1356 2008
rect 1350 2006 1351 2007
rect 1328 2004 1351 2006
rect 1328 2003 1329 2004
rect 1323 2002 1329 2003
rect 1350 2003 1351 2004
rect 1355 2003 1356 2007
rect 1350 2002 1356 2003
rect 1451 2007 1457 2008
rect 1451 2003 1452 2007
rect 1456 2006 1457 2007
rect 1486 2007 1492 2008
rect 1486 2006 1487 2007
rect 1456 2004 1487 2006
rect 1456 2003 1457 2004
rect 1451 2002 1457 2003
rect 1486 2003 1487 2004
rect 1491 2003 1492 2007
rect 1486 2002 1492 2003
rect 1579 2007 1585 2008
rect 1579 2003 1580 2007
rect 1584 2006 1585 2007
rect 1598 2007 1604 2008
rect 1598 2006 1599 2007
rect 1584 2004 1599 2006
rect 1584 2003 1585 2004
rect 1579 2002 1585 2003
rect 1598 2003 1599 2004
rect 1603 2003 1604 2007
rect 1598 2002 1604 2003
rect 424 1996 618 1998
rect 1088 1996 1258 1998
rect 358 1992 364 1993
rect 110 1989 116 1990
rect 110 1985 111 1989
rect 115 1985 116 1989
rect 358 1988 359 1992
rect 363 1988 364 1992
rect 358 1987 364 1988
rect 486 1992 492 1993
rect 486 1988 487 1992
rect 491 1988 492 1992
rect 486 1987 492 1988
rect 110 1984 116 1985
rect 430 1983 436 1984
rect 430 1979 431 1983
rect 435 1979 436 1983
rect 430 1978 436 1979
rect 550 1983 556 1984
rect 550 1979 551 1983
rect 555 1979 556 1983
rect 616 1982 618 1996
rect 622 1992 628 1993
rect 622 1988 623 1992
rect 627 1988 628 1992
rect 622 1987 628 1988
rect 758 1992 764 1993
rect 758 1988 759 1992
rect 763 1988 764 1992
rect 758 1987 764 1988
rect 894 1992 900 1993
rect 894 1988 895 1992
rect 899 1988 900 1992
rect 894 1987 900 1988
rect 1022 1992 1028 1993
rect 1022 1988 1023 1992
rect 1027 1988 1028 1992
rect 1022 1987 1028 1988
rect 1150 1992 1156 1993
rect 1150 1988 1151 1992
rect 1155 1988 1156 1992
rect 1150 1987 1156 1988
rect 871 1983 877 1984
rect 871 1982 872 1983
rect 616 1980 665 1982
rect 833 1980 872 1982
rect 550 1978 556 1979
rect 871 1979 872 1980
rect 876 1979 877 1983
rect 871 1978 877 1979
rect 966 1983 972 1984
rect 966 1979 967 1983
rect 971 1979 972 1983
rect 966 1978 972 1979
rect 1094 1983 1100 1984
rect 1094 1979 1095 1983
rect 1099 1979 1100 1983
rect 1247 1983 1253 1984
rect 1247 1982 1248 1983
rect 1225 1980 1248 1982
rect 1094 1978 1100 1979
rect 1247 1979 1248 1980
rect 1252 1979 1253 1983
rect 1256 1982 1258 1996
rect 1270 1992 1276 1993
rect 1270 1988 1271 1992
rect 1275 1988 1276 1992
rect 1270 1987 1276 1988
rect 1398 1992 1404 1993
rect 1398 1988 1399 1992
rect 1403 1988 1404 1992
rect 1398 1987 1404 1988
rect 1526 1992 1532 1993
rect 1526 1988 1527 1992
rect 1531 1988 1532 1992
rect 1526 1987 1532 1988
rect 1766 1989 1772 1990
rect 1766 1985 1767 1989
rect 1771 1985 1772 1989
rect 1766 1984 1772 1985
rect 1350 1983 1356 1984
rect 1256 1980 1313 1982
rect 1247 1978 1253 1979
rect 1350 1979 1351 1983
rect 1355 1982 1356 1983
rect 1486 1983 1492 1984
rect 1355 1980 1441 1982
rect 1355 1979 1356 1980
rect 1350 1978 1356 1979
rect 1486 1979 1487 1983
rect 1491 1982 1492 1983
rect 1491 1980 1569 1982
rect 1491 1979 1492 1980
rect 1486 1978 1492 1979
rect 358 1973 364 1974
rect 110 1972 116 1973
rect 110 1968 111 1972
rect 115 1968 116 1972
rect 358 1969 359 1973
rect 363 1969 364 1973
rect 358 1968 364 1969
rect 486 1973 492 1974
rect 486 1969 487 1973
rect 491 1969 492 1973
rect 486 1968 492 1969
rect 622 1973 628 1974
rect 622 1969 623 1973
rect 627 1969 628 1973
rect 622 1968 628 1969
rect 758 1973 764 1974
rect 758 1969 759 1973
rect 763 1969 764 1973
rect 758 1968 764 1969
rect 894 1973 900 1974
rect 894 1969 895 1973
rect 899 1969 900 1973
rect 894 1968 900 1969
rect 1022 1973 1028 1974
rect 1022 1969 1023 1973
rect 1027 1969 1028 1973
rect 1022 1968 1028 1969
rect 1150 1973 1156 1974
rect 1150 1969 1151 1973
rect 1155 1969 1156 1973
rect 1150 1968 1156 1969
rect 1270 1973 1276 1974
rect 1270 1969 1271 1973
rect 1275 1969 1276 1973
rect 1270 1968 1276 1969
rect 1398 1973 1404 1974
rect 1398 1969 1399 1973
rect 1403 1969 1404 1973
rect 1398 1968 1404 1969
rect 1526 1973 1532 1974
rect 1526 1969 1527 1973
rect 1531 1969 1532 1973
rect 1526 1968 1532 1969
rect 1766 1972 1772 1973
rect 1766 1968 1767 1972
rect 1771 1968 1772 1972
rect 110 1967 116 1968
rect 1766 1967 1772 1968
rect 1806 1960 1812 1961
rect 3462 1960 3468 1961
rect 1806 1956 1807 1960
rect 1811 1956 1812 1960
rect 1806 1955 1812 1956
rect 1830 1959 1836 1960
rect 1830 1955 1831 1959
rect 1835 1955 1836 1959
rect 1830 1954 1836 1955
rect 1918 1959 1924 1960
rect 1918 1955 1919 1959
rect 1923 1955 1924 1959
rect 1918 1954 1924 1955
rect 2046 1959 2052 1960
rect 2046 1955 2047 1959
rect 2051 1955 2052 1959
rect 2046 1954 2052 1955
rect 2182 1959 2188 1960
rect 2182 1955 2183 1959
rect 2187 1955 2188 1959
rect 2182 1954 2188 1955
rect 2326 1959 2332 1960
rect 2326 1955 2327 1959
rect 2331 1955 2332 1959
rect 2326 1954 2332 1955
rect 2470 1959 2476 1960
rect 2470 1955 2471 1959
rect 2475 1955 2476 1959
rect 2470 1954 2476 1955
rect 2614 1959 2620 1960
rect 2614 1955 2615 1959
rect 2619 1955 2620 1959
rect 2614 1954 2620 1955
rect 2750 1959 2756 1960
rect 2750 1955 2751 1959
rect 2755 1955 2756 1959
rect 2750 1954 2756 1955
rect 2886 1959 2892 1960
rect 2886 1955 2887 1959
rect 2891 1955 2892 1959
rect 2886 1954 2892 1955
rect 3030 1959 3036 1960
rect 3030 1955 3031 1959
rect 3035 1955 3036 1959
rect 3030 1954 3036 1955
rect 3174 1959 3180 1960
rect 3174 1955 3175 1959
rect 3179 1955 3180 1959
rect 3174 1954 3180 1955
rect 3318 1959 3324 1960
rect 3318 1955 3319 1959
rect 3323 1955 3324 1959
rect 3462 1956 3463 1960
rect 3467 1956 3468 1960
rect 3462 1955 3468 1956
rect 3318 1954 3324 1955
rect 1910 1951 1916 1952
rect 1902 1947 1908 1948
rect 1806 1943 1812 1944
rect 1806 1939 1807 1943
rect 1811 1939 1812 1943
rect 1902 1943 1903 1947
rect 1907 1943 1908 1947
rect 1910 1947 1911 1951
rect 1915 1950 1916 1951
rect 1998 1951 2004 1952
rect 1915 1948 1961 1950
rect 1915 1947 1916 1948
rect 1910 1946 1916 1947
rect 1998 1947 1999 1951
rect 2003 1950 2004 1951
rect 2126 1951 2132 1952
rect 2003 1948 2089 1950
rect 2003 1947 2004 1948
rect 1998 1946 2004 1947
rect 2126 1947 2127 1951
rect 2131 1950 2132 1951
rect 2262 1951 2268 1952
rect 2131 1948 2225 1950
rect 2131 1947 2132 1948
rect 2126 1946 2132 1947
rect 2262 1947 2263 1951
rect 2267 1950 2268 1951
rect 3110 1951 3116 1952
rect 2267 1948 2369 1950
rect 2267 1947 2268 1948
rect 2262 1946 2268 1947
rect 2542 1947 2548 1948
rect 1902 1942 1908 1943
rect 2542 1943 2543 1947
rect 2547 1943 2548 1947
rect 2542 1942 2548 1943
rect 2686 1947 2692 1948
rect 2686 1943 2687 1947
rect 2691 1943 2692 1947
rect 2686 1942 2692 1943
rect 2822 1947 2828 1948
rect 2822 1943 2823 1947
rect 2827 1943 2828 1947
rect 2822 1942 2828 1943
rect 2958 1947 2964 1948
rect 2958 1943 2959 1947
rect 2963 1943 2964 1947
rect 2958 1942 2964 1943
rect 3102 1947 3108 1948
rect 3102 1943 3103 1947
rect 3107 1943 3108 1947
rect 3110 1947 3111 1951
rect 3115 1950 3116 1951
rect 3115 1948 3217 1950
rect 3115 1947 3116 1948
rect 3110 1946 3116 1947
rect 3390 1947 3396 1948
rect 3102 1942 3108 1943
rect 3390 1943 3391 1947
rect 3395 1943 3396 1947
rect 3390 1942 3396 1943
rect 3462 1943 3468 1944
rect 1806 1938 1812 1939
rect 1830 1940 1836 1941
rect 1830 1936 1831 1940
rect 1835 1936 1836 1940
rect 1830 1935 1836 1936
rect 1918 1940 1924 1941
rect 1918 1936 1919 1940
rect 1923 1936 1924 1940
rect 1918 1935 1924 1936
rect 2046 1940 2052 1941
rect 2046 1936 2047 1940
rect 2051 1936 2052 1940
rect 2046 1935 2052 1936
rect 2182 1940 2188 1941
rect 2182 1936 2183 1940
rect 2187 1936 2188 1940
rect 2182 1935 2188 1936
rect 2326 1940 2332 1941
rect 2326 1936 2327 1940
rect 2331 1936 2332 1940
rect 2326 1935 2332 1936
rect 2470 1940 2476 1941
rect 2470 1936 2471 1940
rect 2475 1936 2476 1940
rect 2470 1935 2476 1936
rect 2614 1940 2620 1941
rect 2614 1936 2615 1940
rect 2619 1936 2620 1940
rect 2614 1935 2620 1936
rect 2750 1940 2756 1941
rect 2750 1936 2751 1940
rect 2755 1936 2756 1940
rect 2750 1935 2756 1936
rect 2886 1940 2892 1941
rect 2886 1936 2887 1940
rect 2891 1936 2892 1940
rect 2886 1935 2892 1936
rect 3030 1940 3036 1941
rect 3030 1936 3031 1940
rect 3035 1936 3036 1940
rect 3030 1935 3036 1936
rect 3174 1940 3180 1941
rect 3174 1936 3175 1940
rect 3179 1936 3180 1940
rect 3174 1935 3180 1936
rect 3318 1940 3324 1941
rect 3318 1936 3319 1940
rect 3323 1936 3324 1940
rect 3462 1939 3463 1943
rect 3467 1939 3468 1943
rect 3462 1938 3468 1939
rect 3318 1935 3324 1936
rect 110 1928 116 1929
rect 1766 1928 1772 1929
rect 110 1924 111 1928
rect 115 1924 116 1928
rect 110 1923 116 1924
rect 446 1927 452 1928
rect 446 1923 447 1927
rect 451 1923 452 1927
rect 446 1922 452 1923
rect 574 1927 580 1928
rect 574 1923 575 1927
rect 579 1923 580 1927
rect 574 1922 580 1923
rect 710 1927 716 1928
rect 710 1923 711 1927
rect 715 1923 716 1927
rect 710 1922 716 1923
rect 846 1927 852 1928
rect 846 1923 847 1927
rect 851 1923 852 1927
rect 846 1922 852 1923
rect 982 1927 988 1928
rect 982 1923 983 1927
rect 987 1923 988 1927
rect 982 1922 988 1923
rect 1118 1927 1124 1928
rect 1118 1923 1119 1927
rect 1123 1923 1124 1927
rect 1118 1922 1124 1923
rect 1254 1927 1260 1928
rect 1254 1923 1255 1927
rect 1259 1923 1260 1927
rect 1254 1922 1260 1923
rect 1382 1927 1388 1928
rect 1382 1923 1383 1927
rect 1387 1923 1388 1927
rect 1382 1922 1388 1923
rect 1518 1927 1524 1928
rect 1518 1923 1519 1927
rect 1523 1923 1524 1927
rect 1518 1922 1524 1923
rect 1654 1927 1660 1928
rect 1654 1923 1655 1927
rect 1659 1923 1660 1927
rect 1766 1924 1767 1928
rect 1771 1924 1772 1928
rect 1766 1923 1772 1924
rect 1883 1923 1889 1924
rect 1654 1922 1660 1923
rect 702 1919 708 1920
rect 559 1915 565 1916
rect 559 1914 560 1915
rect 521 1912 560 1914
rect 110 1911 116 1912
rect 110 1907 111 1911
rect 115 1907 116 1911
rect 559 1911 560 1912
rect 564 1911 565 1915
rect 559 1910 565 1911
rect 646 1915 652 1916
rect 646 1911 647 1915
rect 651 1911 652 1915
rect 702 1915 703 1919
rect 707 1918 708 1919
rect 926 1919 932 1920
rect 707 1916 753 1918
rect 707 1915 708 1916
rect 702 1914 708 1915
rect 918 1915 924 1916
rect 646 1910 652 1911
rect 918 1911 919 1915
rect 923 1911 924 1915
rect 926 1915 927 1919
rect 931 1918 932 1919
rect 1598 1919 1604 1920
rect 931 1916 1025 1918
rect 931 1915 932 1916
rect 926 1914 932 1915
rect 1190 1915 1196 1916
rect 918 1910 924 1911
rect 1190 1911 1191 1915
rect 1195 1911 1196 1915
rect 1366 1915 1372 1916
rect 1366 1914 1367 1915
rect 1329 1912 1367 1914
rect 1190 1910 1196 1911
rect 1366 1911 1367 1912
rect 1371 1911 1372 1915
rect 1470 1915 1476 1916
rect 1470 1914 1471 1915
rect 1457 1912 1471 1914
rect 1366 1910 1372 1911
rect 1470 1911 1471 1912
rect 1475 1911 1476 1915
rect 1470 1910 1476 1911
rect 1590 1915 1596 1916
rect 1590 1911 1591 1915
rect 1595 1911 1596 1915
rect 1598 1915 1599 1919
rect 1603 1918 1604 1919
rect 1883 1919 1884 1923
rect 1888 1922 1889 1923
rect 1910 1923 1916 1924
rect 1910 1922 1911 1923
rect 1888 1920 1911 1922
rect 1888 1919 1889 1920
rect 1883 1918 1889 1919
rect 1910 1919 1911 1920
rect 1915 1919 1916 1923
rect 1910 1918 1916 1919
rect 1971 1923 1977 1924
rect 1971 1919 1972 1923
rect 1976 1922 1977 1923
rect 1998 1923 2004 1924
rect 1998 1922 1999 1923
rect 1976 1920 1999 1922
rect 1976 1919 1977 1920
rect 1971 1918 1977 1919
rect 1998 1919 1999 1920
rect 2003 1919 2004 1923
rect 1998 1918 2004 1919
rect 2099 1923 2105 1924
rect 2099 1919 2100 1923
rect 2104 1922 2105 1923
rect 2126 1923 2132 1924
rect 2126 1922 2127 1923
rect 2104 1920 2127 1922
rect 2104 1919 2105 1920
rect 2099 1918 2105 1919
rect 2126 1919 2127 1920
rect 2131 1919 2132 1923
rect 2126 1918 2132 1919
rect 2235 1923 2241 1924
rect 2235 1919 2236 1923
rect 2240 1922 2241 1923
rect 2262 1923 2268 1924
rect 2262 1922 2263 1923
rect 2240 1920 2263 1922
rect 2240 1919 2241 1920
rect 2235 1918 2241 1919
rect 2262 1919 2263 1920
rect 2267 1919 2268 1923
rect 2262 1918 2268 1919
rect 2374 1923 2385 1924
rect 2374 1919 2375 1923
rect 2379 1919 2380 1923
rect 2384 1919 2385 1923
rect 2374 1918 2385 1919
rect 2523 1923 2532 1924
rect 2523 1919 2524 1923
rect 2531 1919 2532 1923
rect 2523 1918 2532 1919
rect 2667 1923 2673 1924
rect 2667 1919 2668 1923
rect 2672 1922 2673 1923
rect 2686 1923 2692 1924
rect 2672 1920 2682 1922
rect 2672 1919 2673 1920
rect 2667 1918 2673 1919
rect 1603 1916 1697 1918
rect 1603 1915 1604 1916
rect 1598 1914 1604 1915
rect 1902 1915 1908 1916
rect 1590 1910 1596 1911
rect 1766 1911 1772 1912
rect 110 1906 116 1907
rect 446 1908 452 1909
rect 446 1904 447 1908
rect 451 1904 452 1908
rect 446 1903 452 1904
rect 574 1908 580 1909
rect 574 1904 575 1908
rect 579 1904 580 1908
rect 574 1903 580 1904
rect 710 1908 716 1909
rect 710 1904 711 1908
rect 715 1904 716 1908
rect 710 1903 716 1904
rect 846 1908 852 1909
rect 846 1904 847 1908
rect 851 1904 852 1908
rect 846 1903 852 1904
rect 982 1908 988 1909
rect 982 1904 983 1908
rect 987 1904 988 1908
rect 982 1903 988 1904
rect 1118 1908 1124 1909
rect 1118 1904 1119 1908
rect 1123 1904 1124 1908
rect 1118 1903 1124 1904
rect 1254 1908 1260 1909
rect 1254 1904 1255 1908
rect 1259 1904 1260 1908
rect 1254 1903 1260 1904
rect 1382 1908 1388 1909
rect 1382 1904 1383 1908
rect 1387 1904 1388 1908
rect 1382 1903 1388 1904
rect 1518 1908 1524 1909
rect 1518 1904 1519 1908
rect 1523 1904 1524 1908
rect 1518 1903 1524 1904
rect 1654 1908 1660 1909
rect 1654 1904 1655 1908
rect 1659 1904 1660 1908
rect 1766 1907 1767 1911
rect 1771 1907 1772 1911
rect 1902 1911 1903 1915
rect 1907 1914 1908 1915
rect 2680 1914 2682 1920
rect 2686 1919 2687 1923
rect 2691 1922 2692 1923
rect 2803 1923 2809 1924
rect 2803 1922 2804 1923
rect 2691 1920 2804 1922
rect 2691 1919 2692 1920
rect 2686 1918 2692 1919
rect 2803 1919 2804 1920
rect 2808 1919 2809 1923
rect 2803 1918 2809 1919
rect 2822 1923 2828 1924
rect 2822 1919 2823 1923
rect 2827 1922 2828 1923
rect 2939 1923 2945 1924
rect 2939 1922 2940 1923
rect 2827 1920 2940 1922
rect 2827 1919 2828 1920
rect 2822 1918 2828 1919
rect 2939 1919 2940 1920
rect 2944 1919 2945 1923
rect 2939 1918 2945 1919
rect 2958 1923 2964 1924
rect 2958 1919 2959 1923
rect 2963 1922 2964 1923
rect 3083 1923 3089 1924
rect 3083 1922 3084 1923
rect 2963 1920 3084 1922
rect 2963 1919 2964 1920
rect 2958 1918 2964 1919
rect 3083 1919 3084 1920
rect 3088 1919 3089 1923
rect 3083 1918 3089 1919
rect 3102 1923 3108 1924
rect 3102 1919 3103 1923
rect 3107 1922 3108 1923
rect 3227 1923 3233 1924
rect 3227 1922 3228 1923
rect 3107 1920 3228 1922
rect 3107 1919 3108 1920
rect 3102 1918 3108 1919
rect 3227 1919 3228 1920
rect 3232 1919 3233 1923
rect 3227 1918 3233 1919
rect 3358 1923 3364 1924
rect 3358 1919 3359 1923
rect 3363 1922 3364 1923
rect 3371 1923 3377 1924
rect 3371 1922 3372 1923
rect 3363 1920 3372 1922
rect 3363 1919 3364 1920
rect 3358 1918 3364 1919
rect 3371 1919 3372 1920
rect 3376 1919 3377 1923
rect 3371 1918 3377 1919
rect 3166 1915 3172 1916
rect 3166 1914 3167 1915
rect 1907 1912 1974 1914
rect 2680 1912 3167 1914
rect 1907 1911 1908 1912
rect 1902 1910 1908 1911
rect 1972 1910 1974 1912
rect 3166 1911 3167 1912
rect 3171 1911 3172 1915
rect 3166 1910 3172 1911
rect 1971 1909 1977 1910
rect 1766 1906 1772 1907
rect 1883 1907 1889 1908
rect 1654 1903 1660 1904
rect 1883 1903 1884 1907
rect 1888 1906 1889 1907
rect 1910 1907 1916 1908
rect 1910 1906 1911 1907
rect 1888 1904 1911 1906
rect 1888 1903 1889 1904
rect 1883 1902 1889 1903
rect 1910 1903 1911 1904
rect 1915 1903 1916 1907
rect 1971 1905 1972 1909
rect 1976 1905 1977 1909
rect 1971 1904 1977 1905
rect 2091 1907 2100 1908
rect 1910 1902 1916 1903
rect 2091 1903 2092 1907
rect 2099 1903 2100 1907
rect 2091 1902 2100 1903
rect 2110 1907 2116 1908
rect 2110 1903 2111 1907
rect 2115 1906 2116 1907
rect 2219 1907 2225 1908
rect 2219 1906 2220 1907
rect 2115 1904 2220 1906
rect 2115 1903 2116 1904
rect 2110 1902 2116 1903
rect 2219 1903 2220 1904
rect 2224 1903 2225 1907
rect 2219 1902 2225 1903
rect 2238 1907 2244 1908
rect 2238 1903 2239 1907
rect 2243 1906 2244 1907
rect 2355 1907 2361 1908
rect 2355 1906 2356 1907
rect 2243 1904 2356 1906
rect 2243 1903 2244 1904
rect 2238 1902 2244 1903
rect 2355 1903 2356 1904
rect 2360 1903 2361 1907
rect 2355 1902 2361 1903
rect 2507 1907 2513 1908
rect 2507 1903 2508 1907
rect 2512 1906 2513 1907
rect 2542 1907 2548 1908
rect 2542 1906 2543 1907
rect 2512 1904 2543 1906
rect 2512 1903 2513 1904
rect 2507 1902 2513 1903
rect 2542 1903 2543 1904
rect 2547 1903 2548 1907
rect 2542 1902 2548 1903
rect 2667 1907 2673 1908
rect 2667 1903 2668 1907
rect 2672 1906 2673 1907
rect 2686 1907 2692 1908
rect 2672 1904 2682 1906
rect 2672 1903 2673 1904
rect 2667 1902 2673 1903
rect 1406 1899 1412 1900
rect 1406 1898 1407 1899
rect 1172 1896 1407 1898
rect 1172 1894 1174 1896
rect 1406 1895 1407 1896
rect 1411 1895 1412 1899
rect 2680 1898 2682 1904
rect 2686 1903 2687 1907
rect 2691 1906 2692 1907
rect 2843 1907 2849 1908
rect 2843 1906 2844 1907
rect 2691 1904 2844 1906
rect 2691 1903 2692 1904
rect 2686 1902 2692 1903
rect 2843 1903 2844 1904
rect 2848 1903 2849 1907
rect 2843 1902 2849 1903
rect 2862 1907 2868 1908
rect 2862 1903 2863 1907
rect 2867 1906 2868 1907
rect 3035 1907 3041 1908
rect 3035 1906 3036 1907
rect 2867 1904 3036 1906
rect 2867 1903 2868 1904
rect 2862 1902 2868 1903
rect 3035 1903 3036 1904
rect 3040 1903 3041 1907
rect 3035 1902 3041 1903
rect 3054 1907 3060 1908
rect 3054 1903 3055 1907
rect 3059 1906 3060 1907
rect 3235 1907 3241 1908
rect 3235 1906 3236 1907
rect 3059 1904 3236 1906
rect 3059 1903 3060 1904
rect 3054 1902 3060 1903
rect 3235 1903 3236 1904
rect 3240 1903 3241 1907
rect 3235 1902 3241 1903
rect 3419 1907 3425 1908
rect 3419 1903 3420 1907
rect 3424 1906 3425 1907
rect 3446 1907 3452 1908
rect 3446 1906 3447 1907
rect 3424 1904 3447 1906
rect 3424 1903 3425 1904
rect 3419 1902 3425 1903
rect 3446 1903 3447 1904
rect 3451 1903 3452 1907
rect 3446 1902 3452 1903
rect 3078 1899 3084 1900
rect 3078 1898 3079 1899
rect 2680 1896 3079 1898
rect 1406 1894 1412 1895
rect 3078 1895 3079 1896
rect 3083 1895 3084 1899
rect 3078 1894 3084 1895
rect 1171 1893 1177 1894
rect 499 1891 505 1892
rect 499 1887 500 1891
rect 504 1890 505 1891
rect 538 1891 544 1892
rect 538 1890 539 1891
rect 504 1888 539 1890
rect 504 1887 505 1888
rect 499 1886 505 1887
rect 538 1887 539 1888
rect 543 1887 544 1891
rect 538 1886 544 1887
rect 559 1891 565 1892
rect 559 1887 560 1891
rect 564 1890 565 1891
rect 627 1891 633 1892
rect 627 1890 628 1891
rect 564 1888 628 1890
rect 564 1887 565 1888
rect 559 1886 565 1887
rect 627 1887 628 1888
rect 632 1887 633 1891
rect 627 1886 633 1887
rect 646 1891 652 1892
rect 646 1887 647 1891
rect 651 1890 652 1891
rect 763 1891 769 1892
rect 763 1890 764 1891
rect 651 1888 764 1890
rect 651 1887 652 1888
rect 646 1886 652 1887
rect 763 1887 764 1888
rect 768 1887 769 1891
rect 763 1886 769 1887
rect 899 1891 905 1892
rect 899 1887 900 1891
rect 904 1890 905 1891
rect 926 1891 932 1892
rect 926 1890 927 1891
rect 904 1888 927 1890
rect 904 1887 905 1888
rect 899 1886 905 1887
rect 926 1887 927 1888
rect 931 1887 932 1891
rect 926 1886 932 1887
rect 966 1891 972 1892
rect 966 1887 967 1891
rect 971 1890 972 1891
rect 1035 1891 1041 1892
rect 1035 1890 1036 1891
rect 971 1888 1036 1890
rect 971 1887 972 1888
rect 966 1886 972 1887
rect 1035 1887 1036 1888
rect 1040 1887 1041 1891
rect 1171 1889 1172 1893
rect 1176 1889 1177 1893
rect 1830 1892 1836 1893
rect 1171 1888 1177 1889
rect 1190 1891 1196 1892
rect 1035 1886 1041 1887
rect 1190 1887 1191 1891
rect 1195 1890 1196 1891
rect 1307 1891 1313 1892
rect 1307 1890 1308 1891
rect 1195 1888 1308 1890
rect 1195 1887 1196 1888
rect 1190 1886 1196 1887
rect 1307 1887 1308 1888
rect 1312 1887 1313 1891
rect 1307 1886 1313 1887
rect 1366 1891 1372 1892
rect 1366 1887 1367 1891
rect 1371 1890 1372 1891
rect 1435 1891 1441 1892
rect 1435 1890 1436 1891
rect 1371 1888 1436 1890
rect 1371 1887 1372 1888
rect 1366 1886 1372 1887
rect 1435 1887 1436 1888
rect 1440 1887 1441 1891
rect 1435 1886 1441 1887
rect 1470 1891 1476 1892
rect 1470 1887 1471 1891
rect 1475 1890 1476 1891
rect 1571 1891 1577 1892
rect 1571 1890 1572 1891
rect 1475 1888 1572 1890
rect 1475 1887 1476 1888
rect 1470 1886 1476 1887
rect 1571 1887 1572 1888
rect 1576 1887 1577 1891
rect 1571 1886 1577 1887
rect 1590 1891 1596 1892
rect 1590 1887 1591 1891
rect 1595 1890 1596 1891
rect 1707 1891 1713 1892
rect 1707 1890 1708 1891
rect 1595 1888 1708 1890
rect 1595 1887 1596 1888
rect 1590 1886 1596 1887
rect 1707 1887 1708 1888
rect 1712 1887 1713 1891
rect 1707 1886 1713 1887
rect 1806 1889 1812 1890
rect 1806 1885 1807 1889
rect 1811 1885 1812 1889
rect 1830 1888 1831 1892
rect 1835 1888 1836 1892
rect 1830 1887 1836 1888
rect 1918 1892 1924 1893
rect 1918 1888 1919 1892
rect 1923 1888 1924 1892
rect 1918 1887 1924 1888
rect 2038 1892 2044 1893
rect 2038 1888 2039 1892
rect 2043 1888 2044 1892
rect 2038 1887 2044 1888
rect 2166 1892 2172 1893
rect 2166 1888 2167 1892
rect 2171 1888 2172 1892
rect 2166 1887 2172 1888
rect 2302 1892 2308 1893
rect 2302 1888 2303 1892
rect 2307 1888 2308 1892
rect 2302 1887 2308 1888
rect 2454 1892 2460 1893
rect 2454 1888 2455 1892
rect 2459 1888 2460 1892
rect 2454 1887 2460 1888
rect 2614 1892 2620 1893
rect 2614 1888 2615 1892
rect 2619 1888 2620 1892
rect 2614 1887 2620 1888
rect 2790 1892 2796 1893
rect 2790 1888 2791 1892
rect 2795 1888 2796 1892
rect 2790 1887 2796 1888
rect 2982 1892 2988 1893
rect 2982 1888 2983 1892
rect 2987 1888 2988 1892
rect 2982 1887 2988 1888
rect 3182 1892 3188 1893
rect 3182 1888 3183 1892
rect 3187 1888 3188 1892
rect 3182 1887 3188 1888
rect 3366 1892 3372 1893
rect 3366 1888 3367 1892
rect 3371 1888 3372 1892
rect 3366 1887 3372 1888
rect 3462 1889 3468 1890
rect 1806 1884 1812 1885
rect 3462 1885 3463 1889
rect 3467 1885 3468 1889
rect 3462 1884 3468 1885
rect 1894 1883 1900 1884
rect 611 1879 617 1880
rect 611 1875 612 1879
rect 616 1878 617 1879
rect 646 1879 652 1880
rect 646 1878 647 1879
rect 616 1876 647 1878
rect 616 1875 617 1876
rect 611 1874 617 1875
rect 646 1875 647 1876
rect 651 1875 652 1879
rect 646 1874 652 1875
rect 747 1879 753 1880
rect 747 1875 748 1879
rect 752 1878 753 1879
rect 774 1879 780 1880
rect 774 1878 775 1879
rect 752 1876 775 1878
rect 752 1875 753 1876
rect 747 1874 753 1875
rect 774 1875 775 1876
rect 779 1875 780 1879
rect 774 1874 780 1875
rect 883 1879 889 1880
rect 883 1875 884 1879
rect 888 1878 889 1879
rect 918 1879 924 1880
rect 918 1878 919 1879
rect 888 1876 919 1878
rect 888 1875 889 1876
rect 883 1874 889 1875
rect 918 1875 919 1876
rect 923 1875 924 1879
rect 918 1874 924 1875
rect 1011 1879 1017 1880
rect 1011 1875 1012 1879
rect 1016 1878 1017 1879
rect 1030 1879 1036 1880
rect 1016 1876 1026 1878
rect 1016 1875 1017 1876
rect 1011 1874 1017 1875
rect 1024 1870 1026 1876
rect 1030 1875 1031 1879
rect 1035 1878 1036 1879
rect 1131 1879 1137 1880
rect 1131 1878 1132 1879
rect 1035 1876 1132 1878
rect 1035 1875 1036 1876
rect 1030 1874 1036 1875
rect 1131 1875 1132 1876
rect 1136 1875 1137 1879
rect 1131 1874 1137 1875
rect 1150 1879 1156 1880
rect 1150 1875 1151 1879
rect 1155 1878 1156 1879
rect 1251 1879 1257 1880
rect 1251 1878 1252 1879
rect 1155 1876 1252 1878
rect 1155 1875 1156 1876
rect 1150 1874 1156 1875
rect 1251 1875 1252 1876
rect 1256 1875 1257 1879
rect 1251 1874 1257 1875
rect 1270 1879 1276 1880
rect 1270 1875 1271 1879
rect 1275 1878 1276 1879
rect 1379 1879 1385 1880
rect 1379 1878 1380 1879
rect 1275 1876 1380 1878
rect 1275 1875 1276 1876
rect 1270 1874 1276 1875
rect 1379 1875 1380 1876
rect 1384 1875 1385 1879
rect 1379 1874 1385 1875
rect 1398 1879 1404 1880
rect 1398 1875 1399 1879
rect 1403 1878 1404 1879
rect 1507 1879 1513 1880
rect 1507 1878 1508 1879
rect 1403 1876 1508 1878
rect 1403 1875 1404 1876
rect 1398 1874 1404 1875
rect 1507 1875 1508 1876
rect 1512 1875 1513 1879
rect 1894 1879 1895 1883
rect 1899 1879 1900 1883
rect 1894 1878 1900 1879
rect 1910 1883 1916 1884
rect 1910 1879 1911 1883
rect 1915 1882 1916 1883
rect 2110 1883 2116 1884
rect 1915 1880 1961 1882
rect 1915 1879 1916 1880
rect 1910 1878 1916 1879
rect 2110 1879 2111 1883
rect 2115 1879 2116 1883
rect 2110 1878 2116 1879
rect 2238 1883 2244 1884
rect 2238 1879 2239 1883
rect 2243 1879 2244 1883
rect 2238 1878 2244 1879
rect 2374 1883 2380 1884
rect 2374 1879 2375 1883
rect 2379 1879 2380 1883
rect 2374 1878 2380 1879
rect 2426 1883 2432 1884
rect 2426 1879 2427 1883
rect 2431 1882 2432 1883
rect 2686 1883 2692 1884
rect 2431 1880 2497 1882
rect 2431 1879 2432 1880
rect 2426 1878 2432 1879
rect 2686 1879 2687 1883
rect 2691 1879 2692 1883
rect 2686 1878 2692 1879
rect 2862 1883 2868 1884
rect 2862 1879 2863 1883
rect 2867 1879 2868 1883
rect 2862 1878 2868 1879
rect 3054 1883 3060 1884
rect 3054 1879 3055 1883
rect 3059 1879 3060 1883
rect 3054 1878 3060 1879
rect 3166 1883 3172 1884
rect 3166 1879 3167 1883
rect 3171 1882 3172 1883
rect 3430 1883 3436 1884
rect 3171 1880 3225 1882
rect 3171 1879 3172 1880
rect 3166 1878 3172 1879
rect 3430 1879 3431 1883
rect 3435 1879 3436 1883
rect 3430 1878 3436 1879
rect 1507 1874 1513 1875
rect 1830 1873 1836 1874
rect 1806 1872 1812 1873
rect 1166 1871 1172 1872
rect 1166 1870 1167 1871
rect 1024 1868 1167 1870
rect 1166 1867 1167 1868
rect 1171 1867 1172 1871
rect 1806 1868 1807 1872
rect 1811 1868 1812 1872
rect 1830 1869 1831 1873
rect 1835 1869 1836 1873
rect 1830 1868 1836 1869
rect 1918 1873 1924 1874
rect 1918 1869 1919 1873
rect 1923 1869 1924 1873
rect 1918 1868 1924 1869
rect 2038 1873 2044 1874
rect 2038 1869 2039 1873
rect 2043 1869 2044 1873
rect 2038 1868 2044 1869
rect 2166 1873 2172 1874
rect 2166 1869 2167 1873
rect 2171 1869 2172 1873
rect 2166 1868 2172 1869
rect 2302 1873 2308 1874
rect 2302 1869 2303 1873
rect 2307 1869 2308 1873
rect 2302 1868 2308 1869
rect 2454 1873 2460 1874
rect 2454 1869 2455 1873
rect 2459 1869 2460 1873
rect 2454 1868 2460 1869
rect 2614 1873 2620 1874
rect 2614 1869 2615 1873
rect 2619 1869 2620 1873
rect 2614 1868 2620 1869
rect 2790 1873 2796 1874
rect 2790 1869 2791 1873
rect 2795 1869 2796 1873
rect 2790 1868 2796 1869
rect 2982 1873 2988 1874
rect 2982 1869 2983 1873
rect 2987 1869 2988 1873
rect 2982 1868 2988 1869
rect 3182 1873 3188 1874
rect 3182 1869 3183 1873
rect 3187 1869 3188 1873
rect 3182 1868 3188 1869
rect 3366 1873 3372 1874
rect 3366 1869 3367 1873
rect 3371 1869 3372 1873
rect 3366 1868 3372 1869
rect 3462 1872 3468 1873
rect 3462 1868 3463 1872
rect 3467 1868 3468 1872
rect 1806 1867 1812 1868
rect 3462 1867 3468 1868
rect 1166 1866 1172 1867
rect 558 1864 564 1865
rect 110 1861 116 1862
rect 110 1857 111 1861
rect 115 1857 116 1861
rect 558 1860 559 1864
rect 563 1860 564 1864
rect 558 1859 564 1860
rect 694 1864 700 1865
rect 694 1860 695 1864
rect 699 1860 700 1864
rect 694 1859 700 1860
rect 830 1864 836 1865
rect 830 1860 831 1864
rect 835 1860 836 1864
rect 830 1859 836 1860
rect 958 1864 964 1865
rect 958 1860 959 1864
rect 963 1860 964 1864
rect 958 1859 964 1860
rect 1078 1864 1084 1865
rect 1078 1860 1079 1864
rect 1083 1860 1084 1864
rect 1078 1859 1084 1860
rect 1198 1864 1204 1865
rect 1198 1860 1199 1864
rect 1203 1860 1204 1864
rect 1198 1859 1204 1860
rect 1326 1864 1332 1865
rect 1326 1860 1327 1864
rect 1331 1860 1332 1864
rect 1326 1859 1332 1860
rect 1454 1864 1460 1865
rect 1454 1860 1455 1864
rect 1459 1860 1460 1864
rect 1454 1859 1460 1860
rect 1766 1861 1772 1862
rect 110 1856 116 1857
rect 1766 1857 1767 1861
rect 1771 1857 1772 1861
rect 1766 1856 1772 1857
rect 538 1855 544 1856
rect 538 1851 539 1855
rect 543 1854 544 1855
rect 646 1855 652 1856
rect 543 1852 601 1854
rect 543 1851 544 1852
rect 538 1850 544 1851
rect 646 1851 647 1855
rect 651 1854 652 1855
rect 774 1855 780 1856
rect 651 1852 737 1854
rect 651 1851 652 1852
rect 646 1850 652 1851
rect 774 1851 775 1855
rect 779 1854 780 1855
rect 1030 1855 1036 1856
rect 779 1852 873 1854
rect 779 1851 780 1852
rect 774 1850 780 1851
rect 1030 1851 1031 1855
rect 1035 1851 1036 1855
rect 1030 1850 1036 1851
rect 1150 1855 1156 1856
rect 1150 1851 1151 1855
rect 1155 1851 1156 1855
rect 1150 1850 1156 1851
rect 1270 1855 1276 1856
rect 1270 1851 1271 1855
rect 1275 1851 1276 1855
rect 1270 1850 1276 1851
rect 1398 1855 1404 1856
rect 1398 1851 1399 1855
rect 1403 1851 1404 1855
rect 1398 1850 1404 1851
rect 1406 1855 1412 1856
rect 1406 1851 1407 1855
rect 1411 1854 1412 1855
rect 1411 1852 1497 1854
rect 1411 1851 1412 1852
rect 1406 1850 1412 1851
rect 558 1845 564 1846
rect 110 1844 116 1845
rect 110 1840 111 1844
rect 115 1840 116 1844
rect 558 1841 559 1845
rect 563 1841 564 1845
rect 558 1840 564 1841
rect 694 1845 700 1846
rect 694 1841 695 1845
rect 699 1841 700 1845
rect 694 1840 700 1841
rect 830 1845 836 1846
rect 830 1841 831 1845
rect 835 1841 836 1845
rect 830 1840 836 1841
rect 958 1845 964 1846
rect 958 1841 959 1845
rect 963 1841 964 1845
rect 958 1840 964 1841
rect 1078 1845 1084 1846
rect 1078 1841 1079 1845
rect 1083 1841 1084 1845
rect 1078 1840 1084 1841
rect 1198 1845 1204 1846
rect 1198 1841 1199 1845
rect 1203 1841 1204 1845
rect 1198 1840 1204 1841
rect 1326 1845 1332 1846
rect 1326 1841 1327 1845
rect 1331 1841 1332 1845
rect 1326 1840 1332 1841
rect 1454 1845 1460 1846
rect 1454 1841 1455 1845
rect 1459 1841 1460 1845
rect 1454 1840 1460 1841
rect 1766 1844 1772 1845
rect 1766 1840 1767 1844
rect 1771 1840 1772 1844
rect 110 1839 116 1840
rect 1766 1839 1772 1840
rect 1806 1824 1812 1825
rect 3462 1824 3468 1825
rect 1806 1820 1807 1824
rect 1811 1820 1812 1824
rect 1806 1819 1812 1820
rect 1830 1823 1836 1824
rect 1830 1819 1831 1823
rect 1835 1819 1836 1823
rect 1830 1818 1836 1819
rect 1958 1823 1964 1824
rect 1958 1819 1959 1823
rect 1963 1819 1964 1823
rect 1958 1818 1964 1819
rect 2110 1823 2116 1824
rect 2110 1819 2111 1823
rect 2115 1819 2116 1823
rect 2110 1818 2116 1819
rect 2254 1823 2260 1824
rect 2254 1819 2255 1823
rect 2259 1819 2260 1823
rect 2254 1818 2260 1819
rect 2406 1823 2412 1824
rect 2406 1819 2407 1823
rect 2411 1819 2412 1823
rect 2406 1818 2412 1819
rect 2566 1823 2572 1824
rect 2566 1819 2567 1823
rect 2571 1819 2572 1823
rect 2566 1818 2572 1819
rect 2742 1823 2748 1824
rect 2742 1819 2743 1823
rect 2747 1819 2748 1823
rect 2742 1818 2748 1819
rect 2934 1823 2940 1824
rect 2934 1819 2935 1823
rect 2939 1819 2940 1823
rect 2934 1818 2940 1819
rect 3134 1823 3140 1824
rect 3134 1819 3135 1823
rect 3139 1819 3140 1823
rect 3134 1818 3140 1819
rect 3342 1823 3348 1824
rect 3342 1819 3343 1823
rect 3347 1819 3348 1823
rect 3462 1820 3463 1824
rect 3467 1820 3468 1824
rect 3462 1819 3468 1820
rect 3342 1818 3348 1819
rect 1726 1815 1732 1816
rect 1726 1811 1727 1815
rect 1731 1814 1732 1815
rect 2094 1815 2100 1816
rect 1731 1812 1873 1814
rect 1731 1811 1732 1812
rect 1726 1810 1732 1811
rect 2030 1811 2036 1812
rect 1806 1807 1812 1808
rect 1806 1803 1807 1807
rect 1811 1803 1812 1807
rect 2030 1807 2031 1811
rect 2035 1807 2036 1811
rect 2094 1811 2095 1815
rect 2099 1814 2100 1815
rect 3078 1815 3084 1816
rect 2099 1812 2153 1814
rect 2099 1811 2100 1812
rect 2094 1810 2100 1811
rect 2326 1811 2332 1812
rect 2030 1806 2036 1807
rect 2326 1807 2327 1811
rect 2331 1807 2332 1811
rect 2326 1806 2332 1807
rect 2478 1811 2484 1812
rect 2478 1807 2479 1811
rect 2483 1807 2484 1811
rect 2478 1806 2484 1807
rect 2638 1811 2644 1812
rect 2638 1807 2639 1811
rect 2643 1807 2644 1811
rect 2638 1806 2644 1807
rect 2814 1811 2820 1812
rect 2814 1807 2815 1811
rect 2819 1807 2820 1811
rect 2814 1806 2820 1807
rect 3006 1811 3012 1812
rect 3006 1807 3007 1811
rect 3011 1807 3012 1811
rect 3078 1811 3079 1815
rect 3083 1814 3084 1815
rect 3270 1815 3276 1816
rect 3083 1812 3177 1814
rect 3083 1811 3084 1812
rect 3078 1810 3084 1811
rect 3270 1811 3271 1815
rect 3275 1814 3276 1815
rect 3275 1812 3385 1814
rect 3275 1811 3276 1812
rect 3270 1810 3276 1811
rect 3006 1806 3012 1807
rect 3462 1807 3468 1808
rect 1806 1802 1812 1803
rect 1830 1804 1836 1805
rect 1830 1800 1831 1804
rect 1835 1800 1836 1804
rect 1830 1799 1836 1800
rect 1958 1804 1964 1805
rect 1958 1800 1959 1804
rect 1963 1800 1964 1804
rect 1958 1799 1964 1800
rect 2110 1804 2116 1805
rect 2110 1800 2111 1804
rect 2115 1800 2116 1804
rect 2110 1799 2116 1800
rect 2254 1804 2260 1805
rect 2254 1800 2255 1804
rect 2259 1800 2260 1804
rect 2254 1799 2260 1800
rect 2406 1804 2412 1805
rect 2406 1800 2407 1804
rect 2411 1800 2412 1804
rect 2406 1799 2412 1800
rect 2566 1804 2572 1805
rect 2566 1800 2567 1804
rect 2571 1800 2572 1804
rect 2566 1799 2572 1800
rect 2742 1804 2748 1805
rect 2742 1800 2743 1804
rect 2747 1800 2748 1804
rect 2742 1799 2748 1800
rect 2934 1804 2940 1805
rect 2934 1800 2935 1804
rect 2939 1800 2940 1804
rect 2934 1799 2940 1800
rect 3134 1804 3140 1805
rect 3134 1800 3135 1804
rect 3139 1800 3140 1804
rect 3134 1799 3140 1800
rect 3342 1804 3348 1805
rect 3342 1800 3343 1804
rect 3347 1800 3348 1804
rect 3462 1803 3463 1807
rect 3467 1803 3468 1807
rect 3462 1802 3468 1803
rect 3342 1799 3348 1800
rect 110 1792 116 1793
rect 1766 1792 1772 1793
rect 110 1788 111 1792
rect 115 1788 116 1792
rect 110 1787 116 1788
rect 134 1791 140 1792
rect 134 1787 135 1791
rect 139 1787 140 1791
rect 134 1786 140 1787
rect 222 1791 228 1792
rect 222 1787 223 1791
rect 227 1787 228 1791
rect 222 1786 228 1787
rect 310 1791 316 1792
rect 310 1787 311 1791
rect 315 1787 316 1791
rect 310 1786 316 1787
rect 406 1791 412 1792
rect 406 1787 407 1791
rect 411 1787 412 1791
rect 406 1786 412 1787
rect 526 1791 532 1792
rect 526 1787 527 1791
rect 531 1787 532 1791
rect 526 1786 532 1787
rect 654 1791 660 1792
rect 654 1787 655 1791
rect 659 1787 660 1791
rect 654 1786 660 1787
rect 798 1791 804 1792
rect 798 1787 799 1791
rect 803 1787 804 1791
rect 798 1786 804 1787
rect 942 1791 948 1792
rect 942 1787 943 1791
rect 947 1787 948 1791
rect 942 1786 948 1787
rect 1086 1791 1092 1792
rect 1086 1787 1087 1791
rect 1091 1787 1092 1791
rect 1086 1786 1092 1787
rect 1238 1791 1244 1792
rect 1238 1787 1239 1791
rect 1243 1787 1244 1791
rect 1238 1786 1244 1787
rect 1390 1791 1396 1792
rect 1390 1787 1391 1791
rect 1395 1787 1396 1791
rect 1390 1786 1396 1787
rect 1542 1791 1548 1792
rect 1542 1787 1543 1791
rect 1547 1787 1548 1791
rect 1542 1786 1548 1787
rect 1670 1791 1676 1792
rect 1670 1787 1671 1791
rect 1675 1787 1676 1791
rect 1766 1788 1767 1792
rect 1771 1788 1772 1792
rect 1766 1787 1772 1788
rect 1883 1787 1889 1788
rect 1670 1786 1676 1787
rect 791 1783 797 1784
rect 206 1779 212 1780
rect 110 1775 116 1776
rect 110 1771 111 1775
rect 115 1771 116 1775
rect 206 1775 207 1779
rect 211 1775 212 1779
rect 206 1774 212 1775
rect 294 1779 300 1780
rect 294 1775 295 1779
rect 299 1775 300 1779
rect 294 1774 300 1775
rect 382 1779 388 1780
rect 382 1775 383 1779
rect 387 1775 388 1779
rect 382 1774 388 1775
rect 478 1779 484 1780
rect 478 1775 479 1779
rect 483 1775 484 1779
rect 478 1774 484 1775
rect 598 1779 604 1780
rect 598 1775 599 1779
rect 603 1775 604 1779
rect 598 1774 604 1775
rect 726 1779 732 1780
rect 726 1775 727 1779
rect 731 1775 732 1779
rect 791 1779 792 1783
rect 796 1782 797 1783
rect 1166 1783 1172 1784
rect 796 1780 841 1782
rect 796 1779 797 1780
rect 791 1778 797 1779
rect 1014 1779 1020 1780
rect 726 1774 732 1775
rect 1014 1775 1015 1779
rect 1019 1775 1020 1779
rect 1014 1774 1020 1775
rect 1158 1779 1164 1780
rect 1158 1775 1159 1779
rect 1163 1775 1164 1779
rect 1166 1779 1167 1783
rect 1171 1782 1172 1783
rect 1366 1783 1372 1784
rect 1171 1780 1281 1782
rect 1171 1779 1172 1780
rect 1166 1778 1172 1779
rect 1366 1779 1367 1783
rect 1371 1782 1372 1783
rect 1471 1783 1477 1784
rect 1371 1780 1433 1782
rect 1371 1779 1372 1780
rect 1366 1778 1372 1779
rect 1471 1779 1472 1783
rect 1476 1782 1477 1783
rect 1622 1783 1628 1784
rect 1476 1780 1585 1782
rect 1476 1779 1477 1780
rect 1471 1778 1477 1779
rect 1622 1779 1623 1783
rect 1627 1782 1628 1783
rect 1883 1783 1884 1787
rect 1888 1786 1889 1787
rect 1894 1787 1900 1788
rect 1894 1786 1895 1787
rect 1888 1784 1895 1786
rect 1888 1783 1889 1784
rect 1883 1782 1889 1783
rect 1894 1783 1895 1784
rect 1899 1783 1900 1787
rect 1894 1782 1900 1783
rect 1950 1787 1956 1788
rect 1950 1783 1951 1787
rect 1955 1786 1956 1787
rect 2011 1787 2017 1788
rect 2011 1786 2012 1787
rect 1955 1784 2012 1786
rect 1955 1783 1956 1784
rect 1950 1782 1956 1783
rect 2011 1783 2012 1784
rect 2016 1783 2017 1787
rect 2011 1782 2017 1783
rect 2030 1787 2036 1788
rect 2030 1783 2031 1787
rect 2035 1786 2036 1787
rect 2163 1787 2169 1788
rect 2163 1786 2164 1787
rect 2035 1784 2164 1786
rect 2035 1783 2036 1784
rect 2030 1782 2036 1783
rect 2163 1783 2164 1784
rect 2168 1783 2169 1787
rect 2163 1782 2169 1783
rect 2307 1787 2313 1788
rect 2307 1783 2308 1787
rect 2312 1786 2313 1787
rect 2426 1787 2432 1788
rect 2426 1786 2427 1787
rect 2312 1784 2427 1786
rect 2312 1783 2313 1784
rect 2307 1782 2313 1783
rect 2426 1783 2427 1784
rect 2431 1783 2432 1787
rect 2426 1782 2432 1783
rect 2459 1787 2468 1788
rect 2459 1783 2460 1787
rect 2467 1783 2468 1787
rect 2459 1782 2468 1783
rect 2478 1787 2484 1788
rect 2478 1783 2479 1787
rect 2483 1786 2484 1787
rect 2619 1787 2625 1788
rect 2619 1786 2620 1787
rect 2483 1784 2620 1786
rect 2483 1783 2484 1784
rect 2478 1782 2484 1783
rect 2619 1783 2620 1784
rect 2624 1783 2625 1787
rect 2619 1782 2625 1783
rect 2638 1787 2644 1788
rect 2638 1783 2639 1787
rect 2643 1786 2644 1787
rect 2795 1787 2801 1788
rect 2795 1786 2796 1787
rect 2643 1784 2796 1786
rect 2643 1783 2644 1784
rect 2638 1782 2644 1783
rect 2795 1783 2796 1784
rect 2800 1783 2801 1787
rect 2795 1782 2801 1783
rect 2814 1787 2820 1788
rect 2814 1783 2815 1787
rect 2819 1786 2820 1787
rect 2987 1787 2993 1788
rect 2987 1786 2988 1787
rect 2819 1784 2988 1786
rect 2819 1783 2820 1784
rect 2814 1782 2820 1783
rect 2987 1783 2988 1784
rect 2992 1783 2993 1787
rect 2987 1782 2993 1783
rect 3006 1787 3012 1788
rect 3006 1783 3007 1787
rect 3011 1786 3012 1787
rect 3187 1787 3193 1788
rect 3187 1786 3188 1787
rect 3011 1784 3188 1786
rect 3011 1783 3012 1784
rect 3006 1782 3012 1783
rect 3187 1783 3188 1784
rect 3192 1783 3193 1787
rect 3187 1782 3193 1783
rect 3390 1787 3401 1788
rect 3390 1783 3391 1787
rect 3395 1783 3396 1787
rect 3400 1783 3401 1787
rect 3390 1782 3401 1783
rect 1627 1780 1713 1782
rect 1627 1779 1628 1780
rect 1622 1778 1628 1779
rect 1158 1774 1164 1775
rect 1766 1775 1772 1776
rect 110 1770 116 1771
rect 134 1772 140 1773
rect 134 1768 135 1772
rect 139 1768 140 1772
rect 134 1767 140 1768
rect 222 1772 228 1773
rect 222 1768 223 1772
rect 227 1768 228 1772
rect 222 1767 228 1768
rect 310 1772 316 1773
rect 310 1768 311 1772
rect 315 1768 316 1772
rect 310 1767 316 1768
rect 406 1772 412 1773
rect 406 1768 407 1772
rect 411 1768 412 1772
rect 406 1767 412 1768
rect 526 1772 532 1773
rect 526 1768 527 1772
rect 531 1768 532 1772
rect 526 1767 532 1768
rect 654 1772 660 1773
rect 654 1768 655 1772
rect 659 1768 660 1772
rect 654 1767 660 1768
rect 798 1772 804 1773
rect 798 1768 799 1772
rect 803 1768 804 1772
rect 798 1767 804 1768
rect 942 1772 948 1773
rect 942 1768 943 1772
rect 947 1768 948 1772
rect 942 1767 948 1768
rect 1086 1772 1092 1773
rect 1086 1768 1087 1772
rect 1091 1768 1092 1772
rect 1086 1767 1092 1768
rect 1238 1772 1244 1773
rect 1238 1768 1239 1772
rect 1243 1768 1244 1772
rect 1238 1767 1244 1768
rect 1390 1772 1396 1773
rect 1390 1768 1391 1772
rect 1395 1768 1396 1772
rect 1390 1767 1396 1768
rect 1542 1772 1548 1773
rect 1542 1768 1543 1772
rect 1547 1768 1548 1772
rect 1542 1767 1548 1768
rect 1670 1772 1676 1773
rect 1670 1768 1671 1772
rect 1675 1768 1676 1772
rect 1766 1771 1767 1775
rect 1771 1771 1772 1775
rect 1766 1770 1772 1771
rect 2798 1771 2804 1772
rect 1670 1767 1676 1768
rect 2798 1767 2799 1771
rect 2803 1770 2804 1771
rect 2803 1768 2966 1770
rect 2803 1767 2804 1768
rect 2798 1766 2804 1767
rect 2964 1766 2966 1768
rect 2963 1765 2969 1766
rect 1931 1763 1937 1764
rect 1931 1759 1932 1763
rect 1936 1762 1937 1763
rect 1959 1763 1965 1764
rect 1959 1762 1960 1763
rect 1936 1760 1960 1762
rect 1936 1759 1937 1760
rect 1931 1758 1937 1759
rect 1959 1759 1960 1760
rect 1964 1759 1965 1763
rect 1959 1758 1965 1759
rect 2067 1763 2073 1764
rect 2067 1759 2068 1763
rect 2072 1762 2073 1763
rect 2094 1763 2100 1764
rect 2094 1762 2095 1763
rect 2072 1760 2095 1762
rect 2072 1759 2073 1760
rect 2067 1758 2073 1759
rect 2094 1759 2095 1760
rect 2099 1759 2100 1763
rect 2094 1758 2100 1759
rect 2203 1763 2209 1764
rect 2203 1759 2204 1763
rect 2208 1762 2209 1763
rect 2326 1763 2332 1764
rect 2208 1760 2258 1762
rect 2208 1759 2209 1760
rect 2203 1758 2209 1759
rect 2254 1759 2260 1760
rect 187 1755 193 1756
rect 187 1751 188 1755
rect 192 1754 193 1755
rect 198 1755 204 1756
rect 198 1754 199 1755
rect 192 1752 199 1754
rect 192 1751 193 1752
rect 187 1750 193 1751
rect 198 1751 199 1752
rect 203 1751 204 1755
rect 198 1750 204 1751
rect 206 1755 212 1756
rect 206 1751 207 1755
rect 211 1754 212 1755
rect 275 1755 281 1756
rect 275 1754 276 1755
rect 211 1752 276 1754
rect 211 1751 212 1752
rect 206 1750 212 1751
rect 275 1751 276 1752
rect 280 1751 281 1755
rect 275 1750 281 1751
rect 294 1755 300 1756
rect 294 1751 295 1755
rect 299 1754 300 1755
rect 363 1755 369 1756
rect 363 1754 364 1755
rect 299 1752 364 1754
rect 299 1751 300 1752
rect 294 1750 300 1751
rect 363 1751 364 1752
rect 368 1751 369 1755
rect 363 1750 369 1751
rect 382 1755 388 1756
rect 382 1751 383 1755
rect 387 1754 388 1755
rect 459 1755 465 1756
rect 459 1754 460 1755
rect 387 1752 460 1754
rect 387 1751 388 1752
rect 382 1750 388 1751
rect 459 1751 460 1752
rect 464 1751 465 1755
rect 459 1750 465 1751
rect 478 1755 484 1756
rect 478 1751 479 1755
rect 483 1754 484 1755
rect 579 1755 585 1756
rect 579 1754 580 1755
rect 483 1752 580 1754
rect 483 1751 484 1752
rect 478 1750 484 1751
rect 579 1751 580 1752
rect 584 1751 585 1755
rect 579 1750 585 1751
rect 598 1755 604 1756
rect 598 1751 599 1755
rect 603 1754 604 1755
rect 707 1755 713 1756
rect 707 1754 708 1755
rect 603 1752 708 1754
rect 603 1751 604 1752
rect 598 1750 604 1751
rect 707 1751 708 1752
rect 712 1751 713 1755
rect 707 1750 713 1751
rect 726 1755 732 1756
rect 726 1751 727 1755
rect 731 1754 732 1755
rect 851 1755 857 1756
rect 851 1754 852 1755
rect 731 1752 852 1754
rect 731 1751 732 1752
rect 726 1750 732 1751
rect 851 1751 852 1752
rect 856 1751 857 1755
rect 851 1750 857 1751
rect 995 1755 1004 1756
rect 995 1751 996 1755
rect 1003 1751 1004 1755
rect 995 1750 1004 1751
rect 1014 1755 1020 1756
rect 1014 1751 1015 1755
rect 1019 1754 1020 1755
rect 1139 1755 1145 1756
rect 1139 1754 1140 1755
rect 1019 1752 1140 1754
rect 1019 1751 1020 1752
rect 1014 1750 1020 1751
rect 1139 1751 1140 1752
rect 1144 1751 1145 1755
rect 1139 1750 1145 1751
rect 1158 1755 1164 1756
rect 1158 1751 1159 1755
rect 1163 1754 1164 1755
rect 1291 1755 1297 1756
rect 1291 1754 1292 1755
rect 1163 1752 1292 1754
rect 1163 1751 1164 1752
rect 1158 1750 1164 1751
rect 1291 1751 1292 1752
rect 1296 1751 1297 1755
rect 1291 1750 1297 1751
rect 1443 1755 1449 1756
rect 1443 1751 1444 1755
rect 1448 1754 1449 1755
rect 1471 1755 1477 1756
rect 1471 1754 1472 1755
rect 1448 1752 1472 1754
rect 1448 1751 1449 1752
rect 1443 1750 1449 1751
rect 1471 1751 1472 1752
rect 1476 1751 1477 1755
rect 1471 1750 1477 1751
rect 1595 1755 1601 1756
rect 1595 1751 1596 1755
rect 1600 1754 1601 1755
rect 1622 1755 1628 1756
rect 1622 1754 1623 1755
rect 1600 1752 1623 1754
rect 1600 1751 1601 1752
rect 1595 1750 1601 1751
rect 1622 1751 1623 1752
rect 1627 1751 1628 1755
rect 1622 1750 1628 1751
rect 1723 1755 1732 1756
rect 1723 1751 1724 1755
rect 1731 1751 1732 1755
rect 2254 1755 2255 1759
rect 2259 1755 2260 1759
rect 2326 1759 2327 1763
rect 2331 1762 2332 1763
rect 2355 1763 2361 1764
rect 2355 1762 2356 1763
rect 2331 1760 2356 1762
rect 2331 1759 2332 1760
rect 2326 1758 2332 1759
rect 2355 1759 2356 1760
rect 2360 1759 2361 1763
rect 2355 1758 2361 1759
rect 2531 1763 2537 1764
rect 2531 1759 2532 1763
rect 2536 1762 2537 1763
rect 2558 1763 2564 1764
rect 2558 1762 2559 1763
rect 2536 1760 2559 1762
rect 2536 1759 2537 1760
rect 2531 1758 2537 1759
rect 2558 1759 2559 1760
rect 2563 1759 2564 1763
rect 2558 1758 2564 1759
rect 2739 1763 2745 1764
rect 2739 1759 2740 1763
rect 2744 1762 2745 1763
rect 2744 1760 2958 1762
rect 2963 1761 2964 1765
rect 2968 1761 2969 1765
rect 2963 1760 2969 1761
rect 2982 1763 2988 1764
rect 2744 1759 2745 1760
rect 2739 1758 2745 1759
rect 2254 1754 2260 1755
rect 2956 1754 2958 1760
rect 2982 1759 2983 1763
rect 2987 1762 2988 1763
rect 3203 1763 3209 1764
rect 3203 1762 3204 1763
rect 2987 1760 3204 1762
rect 2987 1759 2988 1760
rect 2982 1758 2988 1759
rect 3203 1759 3204 1760
rect 3208 1759 3209 1763
rect 3203 1758 3209 1759
rect 3419 1763 3425 1764
rect 3419 1759 3420 1763
rect 3424 1762 3425 1763
rect 3430 1763 3436 1764
rect 3430 1762 3431 1763
rect 3424 1760 3431 1762
rect 3424 1759 3425 1760
rect 3419 1758 3425 1759
rect 3430 1759 3431 1760
rect 3435 1759 3436 1763
rect 3430 1758 3436 1759
rect 2956 1752 3082 1754
rect 1723 1750 1732 1751
rect 1878 1748 1884 1749
rect 1806 1745 1812 1746
rect 1806 1741 1807 1745
rect 1811 1741 1812 1745
rect 1878 1744 1879 1748
rect 1883 1744 1884 1748
rect 1878 1743 1884 1744
rect 2014 1748 2020 1749
rect 2014 1744 2015 1748
rect 2019 1744 2020 1748
rect 2014 1743 2020 1744
rect 2150 1748 2156 1749
rect 2150 1744 2151 1748
rect 2155 1744 2156 1748
rect 2150 1743 2156 1744
rect 2302 1748 2308 1749
rect 2302 1744 2303 1748
rect 2307 1744 2308 1748
rect 2302 1743 2308 1744
rect 2478 1748 2484 1749
rect 2478 1744 2479 1748
rect 2483 1744 2484 1748
rect 2478 1743 2484 1744
rect 2686 1748 2692 1749
rect 2686 1744 2687 1748
rect 2691 1744 2692 1748
rect 2686 1743 2692 1744
rect 2910 1748 2916 1749
rect 2910 1744 2911 1748
rect 2915 1744 2916 1748
rect 2910 1743 2916 1744
rect 1806 1740 1812 1741
rect 1950 1739 1956 1740
rect 1950 1735 1951 1739
rect 1955 1735 1956 1739
rect 1950 1734 1956 1735
rect 1959 1739 1965 1740
rect 1959 1735 1960 1739
rect 1964 1738 1965 1739
rect 2094 1739 2100 1740
rect 1964 1736 2057 1738
rect 1964 1735 1965 1736
rect 1959 1734 1965 1735
rect 2094 1735 2095 1739
rect 2099 1738 2100 1739
rect 2366 1739 2372 1740
rect 2099 1736 2193 1738
rect 2099 1735 2100 1736
rect 2094 1734 2100 1735
rect 2366 1735 2367 1739
rect 2371 1735 2372 1739
rect 2366 1734 2372 1735
rect 2462 1739 2468 1740
rect 2462 1735 2463 1739
rect 2467 1738 2468 1739
rect 2558 1739 2564 1740
rect 2467 1736 2521 1738
rect 2467 1735 2468 1736
rect 2462 1734 2468 1735
rect 2558 1735 2559 1739
rect 2563 1738 2564 1739
rect 2982 1739 2988 1740
rect 2563 1736 2729 1738
rect 2563 1735 2564 1736
rect 2558 1734 2564 1735
rect 2982 1735 2983 1739
rect 2987 1735 2988 1739
rect 3080 1738 3082 1752
rect 3150 1748 3156 1749
rect 3150 1744 3151 1748
rect 3155 1744 3156 1748
rect 3150 1743 3156 1744
rect 3366 1748 3372 1749
rect 3366 1744 3367 1748
rect 3371 1744 3372 1748
rect 3366 1743 3372 1744
rect 3462 1745 3468 1746
rect 3462 1741 3463 1745
rect 3467 1741 3468 1745
rect 3462 1740 3468 1741
rect 3446 1739 3452 1740
rect 3446 1738 3447 1739
rect 3080 1736 3193 1738
rect 3441 1736 3447 1738
rect 2982 1734 2988 1735
rect 3446 1735 3447 1736
rect 3451 1735 3452 1739
rect 3446 1734 3452 1735
rect 187 1731 193 1732
rect 187 1727 188 1731
rect 192 1730 193 1731
rect 214 1731 220 1732
rect 214 1730 215 1731
rect 192 1728 215 1730
rect 192 1727 193 1728
rect 187 1726 193 1727
rect 214 1727 215 1728
rect 219 1727 220 1731
rect 214 1726 220 1727
rect 299 1731 305 1732
rect 299 1727 300 1731
rect 304 1730 305 1731
rect 326 1731 332 1732
rect 326 1730 327 1731
rect 304 1728 327 1730
rect 304 1727 305 1728
rect 299 1726 305 1727
rect 326 1727 327 1728
rect 331 1727 332 1731
rect 326 1726 332 1727
rect 451 1731 457 1732
rect 451 1727 452 1731
rect 456 1730 457 1731
rect 478 1731 484 1732
rect 478 1730 479 1731
rect 456 1728 479 1730
rect 456 1727 457 1728
rect 451 1726 457 1727
rect 478 1727 479 1728
rect 483 1727 484 1731
rect 478 1726 484 1727
rect 619 1731 625 1732
rect 619 1727 620 1731
rect 624 1730 625 1731
rect 734 1731 740 1732
rect 734 1730 735 1731
rect 624 1728 735 1730
rect 624 1727 625 1728
rect 619 1726 625 1727
rect 734 1727 735 1728
rect 739 1727 740 1731
rect 734 1726 740 1727
rect 791 1731 797 1732
rect 791 1727 792 1731
rect 796 1730 797 1731
rect 803 1731 809 1732
rect 803 1730 804 1731
rect 796 1728 804 1730
rect 796 1727 797 1728
rect 791 1726 797 1727
rect 803 1727 804 1728
rect 808 1727 809 1731
rect 803 1726 809 1727
rect 987 1731 993 1732
rect 987 1727 988 1731
rect 992 1730 993 1731
rect 1014 1731 1020 1732
rect 1014 1730 1015 1731
rect 992 1728 1015 1730
rect 992 1727 993 1728
rect 987 1726 993 1727
rect 1014 1727 1015 1728
rect 1019 1727 1020 1731
rect 1014 1726 1020 1727
rect 1171 1731 1180 1732
rect 1171 1727 1172 1731
rect 1179 1727 1180 1731
rect 1171 1726 1180 1727
rect 1363 1731 1372 1732
rect 1363 1727 1364 1731
rect 1371 1727 1372 1731
rect 1363 1726 1372 1727
rect 1382 1731 1388 1732
rect 1382 1727 1383 1731
rect 1387 1730 1388 1731
rect 1555 1731 1561 1732
rect 1555 1730 1556 1731
rect 1387 1728 1556 1730
rect 1387 1727 1388 1728
rect 1382 1726 1388 1727
rect 1555 1727 1556 1728
rect 1560 1727 1561 1731
rect 1555 1726 1561 1727
rect 1574 1731 1580 1732
rect 1574 1727 1575 1731
rect 1579 1730 1580 1731
rect 1723 1731 1729 1732
rect 1723 1730 1724 1731
rect 1579 1728 1724 1730
rect 1579 1727 1580 1728
rect 1574 1726 1580 1727
rect 1723 1727 1724 1728
rect 1728 1727 1729 1731
rect 1878 1729 1884 1730
rect 1723 1726 1729 1727
rect 1806 1728 1812 1729
rect 1806 1724 1807 1728
rect 1811 1724 1812 1728
rect 1878 1725 1879 1729
rect 1883 1725 1884 1729
rect 1878 1724 1884 1725
rect 2014 1729 2020 1730
rect 2014 1725 2015 1729
rect 2019 1725 2020 1729
rect 2014 1724 2020 1725
rect 2150 1729 2156 1730
rect 2150 1725 2151 1729
rect 2155 1725 2156 1729
rect 2150 1724 2156 1725
rect 2302 1729 2308 1730
rect 2302 1725 2303 1729
rect 2307 1725 2308 1729
rect 2302 1724 2308 1725
rect 2478 1729 2484 1730
rect 2478 1725 2479 1729
rect 2483 1725 2484 1729
rect 2478 1724 2484 1725
rect 2686 1729 2692 1730
rect 2686 1725 2687 1729
rect 2691 1725 2692 1729
rect 2686 1724 2692 1725
rect 2910 1729 2916 1730
rect 2910 1725 2911 1729
rect 2915 1725 2916 1729
rect 2910 1724 2916 1725
rect 3150 1729 3156 1730
rect 3150 1725 3151 1729
rect 3155 1725 3156 1729
rect 3150 1724 3156 1725
rect 3366 1729 3372 1730
rect 3366 1725 3367 1729
rect 3371 1725 3372 1729
rect 3366 1724 3372 1725
rect 3462 1728 3468 1729
rect 3462 1724 3463 1728
rect 3467 1724 3468 1728
rect 1806 1723 1812 1724
rect 3462 1723 3468 1724
rect 134 1716 140 1717
rect 110 1713 116 1714
rect 110 1709 111 1713
rect 115 1709 116 1713
rect 134 1712 135 1716
rect 139 1712 140 1716
rect 134 1711 140 1712
rect 246 1716 252 1717
rect 246 1712 247 1716
rect 251 1712 252 1716
rect 246 1711 252 1712
rect 398 1716 404 1717
rect 398 1712 399 1716
rect 403 1712 404 1716
rect 398 1711 404 1712
rect 566 1716 572 1717
rect 566 1712 567 1716
rect 571 1712 572 1716
rect 566 1711 572 1712
rect 750 1716 756 1717
rect 750 1712 751 1716
rect 755 1712 756 1716
rect 750 1711 756 1712
rect 934 1716 940 1717
rect 934 1712 935 1716
rect 939 1712 940 1716
rect 934 1711 940 1712
rect 1118 1716 1124 1717
rect 1118 1712 1119 1716
rect 1123 1712 1124 1716
rect 1118 1711 1124 1712
rect 1310 1716 1316 1717
rect 1310 1712 1311 1716
rect 1315 1712 1316 1716
rect 1310 1711 1316 1712
rect 1502 1716 1508 1717
rect 1502 1712 1503 1716
rect 1507 1712 1508 1716
rect 1502 1711 1508 1712
rect 1670 1716 1676 1717
rect 1670 1712 1671 1716
rect 1675 1712 1676 1716
rect 1670 1711 1676 1712
rect 1766 1713 1772 1714
rect 110 1708 116 1709
rect 1766 1709 1767 1713
rect 1771 1709 1772 1713
rect 1766 1708 1772 1709
rect 198 1707 204 1708
rect 198 1703 199 1707
rect 203 1703 204 1707
rect 198 1702 204 1703
rect 214 1707 220 1708
rect 214 1703 215 1707
rect 219 1706 220 1707
rect 326 1707 332 1708
rect 219 1704 289 1706
rect 219 1703 220 1704
rect 214 1702 220 1703
rect 326 1703 327 1707
rect 331 1706 332 1707
rect 722 1707 728 1708
rect 722 1706 723 1707
rect 331 1704 441 1706
rect 641 1704 723 1706
rect 331 1703 332 1704
rect 326 1702 332 1703
rect 722 1703 723 1704
rect 727 1703 728 1707
rect 722 1702 728 1703
rect 734 1707 740 1708
rect 734 1703 735 1707
rect 739 1706 740 1707
rect 998 1707 1004 1708
rect 739 1704 793 1706
rect 739 1703 740 1704
rect 734 1702 740 1703
rect 998 1703 999 1707
rect 1003 1703 1004 1707
rect 998 1702 1004 1703
rect 1014 1707 1020 1708
rect 1014 1703 1015 1707
rect 1019 1706 1020 1707
rect 1382 1707 1388 1708
rect 1019 1704 1161 1706
rect 1019 1703 1020 1704
rect 1014 1702 1020 1703
rect 1382 1703 1383 1707
rect 1387 1703 1388 1707
rect 1382 1702 1388 1703
rect 1574 1707 1580 1708
rect 1574 1703 1575 1707
rect 1579 1703 1580 1707
rect 1574 1702 1580 1703
rect 1734 1707 1740 1708
rect 1734 1703 1735 1707
rect 1739 1703 1740 1707
rect 1734 1702 1740 1703
rect 134 1697 140 1698
rect 110 1696 116 1697
rect 110 1692 111 1696
rect 115 1692 116 1696
rect 134 1693 135 1697
rect 139 1693 140 1697
rect 134 1692 140 1693
rect 246 1697 252 1698
rect 246 1693 247 1697
rect 251 1693 252 1697
rect 246 1692 252 1693
rect 398 1697 404 1698
rect 398 1693 399 1697
rect 403 1693 404 1697
rect 398 1692 404 1693
rect 566 1697 572 1698
rect 566 1693 567 1697
rect 571 1693 572 1697
rect 566 1692 572 1693
rect 750 1697 756 1698
rect 750 1693 751 1697
rect 755 1693 756 1697
rect 750 1692 756 1693
rect 934 1697 940 1698
rect 934 1693 935 1697
rect 939 1693 940 1697
rect 934 1692 940 1693
rect 1118 1697 1124 1698
rect 1118 1693 1119 1697
rect 1123 1693 1124 1697
rect 1118 1692 1124 1693
rect 1310 1697 1316 1698
rect 1310 1693 1311 1697
rect 1315 1693 1316 1697
rect 1310 1692 1316 1693
rect 1502 1697 1508 1698
rect 1502 1693 1503 1697
rect 1507 1693 1508 1697
rect 1502 1692 1508 1693
rect 1670 1697 1676 1698
rect 1670 1693 1671 1697
rect 1675 1693 1676 1697
rect 1670 1692 1676 1693
rect 1766 1696 1772 1697
rect 1766 1692 1767 1696
rect 1771 1692 1772 1696
rect 110 1691 116 1692
rect 1766 1691 1772 1692
rect 1806 1676 1812 1677
rect 3462 1676 3468 1677
rect 1806 1672 1807 1676
rect 1811 1672 1812 1676
rect 1806 1671 1812 1672
rect 1830 1675 1836 1676
rect 1830 1671 1831 1675
rect 1835 1671 1836 1675
rect 1830 1670 1836 1671
rect 1934 1675 1940 1676
rect 1934 1671 1935 1675
rect 1939 1671 1940 1675
rect 1934 1670 1940 1671
rect 2062 1675 2068 1676
rect 2062 1671 2063 1675
rect 2067 1671 2068 1675
rect 2062 1670 2068 1671
rect 2182 1675 2188 1676
rect 2182 1671 2183 1675
rect 2187 1671 2188 1675
rect 2182 1670 2188 1671
rect 2310 1675 2316 1676
rect 2310 1671 2311 1675
rect 2315 1671 2316 1675
rect 2310 1670 2316 1671
rect 2438 1675 2444 1676
rect 2438 1671 2439 1675
rect 2443 1671 2444 1675
rect 2438 1670 2444 1671
rect 2574 1675 2580 1676
rect 2574 1671 2575 1675
rect 2579 1671 2580 1675
rect 2574 1670 2580 1671
rect 2726 1675 2732 1676
rect 2726 1671 2727 1675
rect 2731 1671 2732 1675
rect 2726 1670 2732 1671
rect 2886 1675 2892 1676
rect 2886 1671 2887 1675
rect 2891 1671 2892 1675
rect 2886 1670 2892 1671
rect 3046 1675 3052 1676
rect 3046 1671 3047 1675
rect 3051 1671 3052 1675
rect 3046 1670 3052 1671
rect 3214 1675 3220 1676
rect 3214 1671 3215 1675
rect 3219 1671 3220 1675
rect 3214 1670 3220 1671
rect 3366 1675 3372 1676
rect 3366 1671 3367 1675
rect 3371 1671 3372 1675
rect 3462 1672 3463 1676
rect 3467 1672 3468 1676
rect 3366 1670 3372 1671
rect 3430 1671 3436 1672
rect 3462 1671 3468 1672
rect 2254 1667 2260 1668
rect 1902 1663 1908 1664
rect 1806 1659 1812 1660
rect 1806 1655 1807 1659
rect 1811 1655 1812 1659
rect 1902 1659 1903 1663
rect 1907 1659 1908 1663
rect 1902 1658 1908 1659
rect 2006 1663 2012 1664
rect 2006 1659 2007 1663
rect 2011 1659 2012 1663
rect 2006 1658 2012 1659
rect 2134 1663 2140 1664
rect 2134 1659 2135 1663
rect 2139 1659 2140 1663
rect 2254 1663 2255 1667
rect 2259 1663 2260 1667
rect 2798 1667 2804 1668
rect 2254 1662 2260 1663
rect 2382 1663 2388 1664
rect 2134 1658 2140 1659
rect 2382 1659 2383 1663
rect 2387 1659 2388 1663
rect 2382 1658 2388 1659
rect 2510 1663 2516 1664
rect 2510 1659 2511 1663
rect 2515 1659 2516 1663
rect 2510 1658 2516 1659
rect 2646 1663 2652 1664
rect 2646 1659 2647 1663
rect 2651 1659 2652 1663
rect 2798 1663 2799 1667
rect 2803 1663 2804 1667
rect 2798 1662 2804 1663
rect 2806 1667 2812 1668
rect 2806 1663 2807 1667
rect 2811 1666 2812 1667
rect 2966 1667 2972 1668
rect 2811 1664 2929 1666
rect 2811 1663 2812 1664
rect 2806 1662 2812 1663
rect 2966 1663 2967 1667
rect 2971 1666 2972 1667
rect 3186 1667 3192 1668
rect 2971 1664 3089 1666
rect 2971 1663 2972 1664
rect 2966 1662 2972 1663
rect 3186 1663 3187 1667
rect 3191 1666 3192 1667
rect 3430 1667 3431 1671
rect 3435 1670 3436 1671
rect 3435 1668 3442 1670
rect 3435 1667 3436 1668
rect 3430 1666 3436 1667
rect 3191 1664 3257 1666
rect 3440 1665 3442 1668
rect 3191 1663 3192 1664
rect 3186 1662 3192 1663
rect 2646 1658 2652 1659
rect 3462 1659 3468 1660
rect 1806 1654 1812 1655
rect 1830 1656 1836 1657
rect 1830 1652 1831 1656
rect 1835 1652 1836 1656
rect 1830 1651 1836 1652
rect 1934 1656 1940 1657
rect 1934 1652 1935 1656
rect 1939 1652 1940 1656
rect 1934 1651 1940 1652
rect 2062 1656 2068 1657
rect 2062 1652 2063 1656
rect 2067 1652 2068 1656
rect 2062 1651 2068 1652
rect 2182 1656 2188 1657
rect 2182 1652 2183 1656
rect 2187 1652 2188 1656
rect 2182 1651 2188 1652
rect 2310 1656 2316 1657
rect 2310 1652 2311 1656
rect 2315 1652 2316 1656
rect 2310 1651 2316 1652
rect 2438 1656 2444 1657
rect 2438 1652 2439 1656
rect 2443 1652 2444 1656
rect 2438 1651 2444 1652
rect 2574 1656 2580 1657
rect 2574 1652 2575 1656
rect 2579 1652 2580 1656
rect 2574 1651 2580 1652
rect 2726 1656 2732 1657
rect 2726 1652 2727 1656
rect 2731 1652 2732 1656
rect 2726 1651 2732 1652
rect 2886 1656 2892 1657
rect 2886 1652 2887 1656
rect 2891 1652 2892 1656
rect 2886 1651 2892 1652
rect 3046 1656 3052 1657
rect 3046 1652 3047 1656
rect 3051 1652 3052 1656
rect 3046 1651 3052 1652
rect 3214 1656 3220 1657
rect 3214 1652 3215 1656
rect 3219 1652 3220 1656
rect 3214 1651 3220 1652
rect 3366 1656 3372 1657
rect 3366 1652 3367 1656
rect 3371 1652 3372 1656
rect 3462 1655 3463 1659
rect 3467 1655 3468 1659
rect 3462 1654 3468 1655
rect 3366 1651 3372 1652
rect 110 1648 116 1649
rect 1766 1648 1772 1649
rect 110 1644 111 1648
rect 115 1644 116 1648
rect 110 1643 116 1644
rect 190 1647 196 1648
rect 190 1643 191 1647
rect 195 1643 196 1647
rect 190 1642 196 1643
rect 294 1647 300 1648
rect 294 1643 295 1647
rect 299 1643 300 1647
rect 294 1642 300 1643
rect 406 1647 412 1648
rect 406 1643 407 1647
rect 411 1643 412 1647
rect 406 1642 412 1643
rect 534 1647 540 1648
rect 534 1643 535 1647
rect 539 1643 540 1647
rect 534 1642 540 1643
rect 686 1647 692 1648
rect 686 1643 687 1647
rect 691 1643 692 1647
rect 686 1642 692 1643
rect 854 1647 860 1648
rect 854 1643 855 1647
rect 859 1643 860 1647
rect 854 1642 860 1643
rect 1038 1647 1044 1648
rect 1038 1643 1039 1647
rect 1043 1643 1044 1647
rect 1038 1642 1044 1643
rect 1230 1647 1236 1648
rect 1230 1643 1231 1647
rect 1235 1643 1236 1647
rect 1230 1642 1236 1643
rect 1430 1647 1436 1648
rect 1430 1643 1431 1647
rect 1435 1643 1436 1647
rect 1430 1642 1436 1643
rect 1638 1647 1644 1648
rect 1638 1643 1639 1647
rect 1643 1643 1644 1647
rect 1766 1644 1767 1648
rect 1771 1644 1772 1648
rect 2806 1647 2812 1648
rect 2806 1646 2807 1647
rect 1766 1643 1772 1644
rect 2492 1644 2807 1646
rect 1638 1642 1644 1643
rect 2492 1642 2494 1644
rect 2806 1643 2807 1644
rect 2811 1643 2812 1647
rect 2806 1642 2812 1643
rect 2491 1641 2497 1642
rect 478 1639 484 1640
rect 262 1635 268 1636
rect 110 1631 116 1632
rect 110 1627 111 1631
rect 115 1627 116 1631
rect 262 1631 263 1635
rect 267 1631 268 1635
rect 262 1630 268 1631
rect 366 1635 372 1636
rect 366 1631 367 1635
rect 371 1631 372 1635
rect 478 1635 479 1639
rect 483 1635 484 1639
rect 614 1639 620 1640
rect 478 1634 484 1635
rect 606 1635 612 1636
rect 366 1630 372 1631
rect 606 1631 607 1635
rect 611 1631 612 1635
rect 614 1635 615 1639
rect 619 1638 620 1639
rect 1174 1639 1180 1640
rect 619 1636 729 1638
rect 619 1635 620 1636
rect 614 1634 620 1635
rect 926 1635 932 1636
rect 606 1630 612 1631
rect 926 1631 927 1635
rect 931 1631 932 1635
rect 926 1630 932 1631
rect 1110 1635 1116 1636
rect 1110 1631 1111 1635
rect 1115 1631 1116 1635
rect 1174 1635 1175 1639
rect 1179 1638 1180 1639
rect 1510 1639 1516 1640
rect 1179 1636 1273 1638
rect 1179 1635 1180 1636
rect 1174 1634 1180 1635
rect 1502 1635 1508 1636
rect 1110 1630 1116 1631
rect 1502 1631 1503 1635
rect 1507 1631 1508 1635
rect 1510 1635 1511 1639
rect 1515 1638 1516 1639
rect 1883 1639 1889 1640
rect 1515 1636 1681 1638
rect 1515 1635 1516 1636
rect 1510 1634 1516 1635
rect 1883 1635 1884 1639
rect 1888 1638 1889 1639
rect 1894 1639 1900 1640
rect 1894 1638 1895 1639
rect 1888 1636 1895 1638
rect 1888 1635 1889 1636
rect 1883 1634 1889 1635
rect 1894 1635 1895 1636
rect 1899 1635 1900 1639
rect 1894 1634 1900 1635
rect 1902 1639 1908 1640
rect 1902 1635 1903 1639
rect 1907 1638 1908 1639
rect 1987 1639 1993 1640
rect 1987 1638 1988 1639
rect 1907 1636 1988 1638
rect 1907 1635 1908 1636
rect 1902 1634 1908 1635
rect 1987 1635 1988 1636
rect 1992 1635 1993 1639
rect 1987 1634 1993 1635
rect 2006 1639 2012 1640
rect 2006 1635 2007 1639
rect 2011 1638 2012 1639
rect 2115 1639 2121 1640
rect 2115 1638 2116 1639
rect 2011 1636 2116 1638
rect 2011 1635 2012 1636
rect 2006 1634 2012 1635
rect 2115 1635 2116 1636
rect 2120 1635 2121 1639
rect 2115 1634 2121 1635
rect 2134 1639 2140 1640
rect 2134 1635 2135 1639
rect 2139 1638 2140 1639
rect 2235 1639 2241 1640
rect 2235 1638 2236 1639
rect 2139 1636 2236 1638
rect 2139 1635 2140 1636
rect 2134 1634 2140 1635
rect 2235 1635 2236 1636
rect 2240 1635 2241 1639
rect 2235 1634 2241 1635
rect 2363 1639 2372 1640
rect 2363 1635 2364 1639
rect 2371 1635 2372 1639
rect 2491 1637 2492 1641
rect 2496 1637 2497 1641
rect 2491 1636 2497 1637
rect 2510 1639 2516 1640
rect 2363 1634 2372 1635
rect 2510 1635 2511 1639
rect 2515 1638 2516 1639
rect 2627 1639 2633 1640
rect 2627 1638 2628 1639
rect 2515 1636 2628 1638
rect 2515 1635 2516 1636
rect 2510 1634 2516 1635
rect 2627 1635 2628 1636
rect 2632 1635 2633 1639
rect 2627 1634 2633 1635
rect 2646 1639 2652 1640
rect 2646 1635 2647 1639
rect 2651 1638 2652 1639
rect 2779 1639 2785 1640
rect 2779 1638 2780 1639
rect 2651 1636 2780 1638
rect 2651 1635 2652 1636
rect 2646 1634 2652 1635
rect 2779 1635 2780 1636
rect 2784 1635 2785 1639
rect 2779 1634 2785 1635
rect 2939 1639 2945 1640
rect 2939 1635 2940 1639
rect 2944 1638 2945 1639
rect 2966 1639 2972 1640
rect 2966 1638 2967 1639
rect 2944 1636 2967 1638
rect 2944 1635 2945 1636
rect 2939 1634 2945 1635
rect 2966 1635 2967 1636
rect 2971 1635 2972 1639
rect 2966 1634 2972 1635
rect 3086 1639 3092 1640
rect 3086 1635 3087 1639
rect 3091 1638 3092 1639
rect 3099 1639 3105 1640
rect 3099 1638 3100 1639
rect 3091 1636 3100 1638
rect 3091 1635 3092 1636
rect 3086 1634 3092 1635
rect 3099 1635 3100 1636
rect 3104 1635 3105 1639
rect 3099 1634 3105 1635
rect 3267 1639 3276 1640
rect 3267 1635 3268 1639
rect 3275 1635 3276 1639
rect 3267 1634 3276 1635
rect 3419 1639 3425 1640
rect 3419 1635 3420 1639
rect 3424 1638 3425 1639
rect 3430 1639 3436 1640
rect 3430 1638 3431 1639
rect 3424 1636 3431 1638
rect 3424 1635 3425 1636
rect 3419 1634 3425 1635
rect 3430 1635 3431 1636
rect 3435 1635 3436 1639
rect 3430 1634 3436 1635
rect 1502 1630 1508 1631
rect 1766 1631 1772 1632
rect 110 1626 116 1627
rect 190 1628 196 1629
rect 190 1624 191 1628
rect 195 1624 196 1628
rect 190 1623 196 1624
rect 294 1628 300 1629
rect 294 1624 295 1628
rect 299 1624 300 1628
rect 294 1623 300 1624
rect 406 1628 412 1629
rect 406 1624 407 1628
rect 411 1624 412 1628
rect 406 1623 412 1624
rect 534 1628 540 1629
rect 534 1624 535 1628
rect 539 1624 540 1628
rect 534 1623 540 1624
rect 686 1628 692 1629
rect 686 1624 687 1628
rect 691 1624 692 1628
rect 686 1623 692 1624
rect 854 1628 860 1629
rect 854 1624 855 1628
rect 859 1624 860 1628
rect 854 1623 860 1624
rect 1038 1628 1044 1629
rect 1038 1624 1039 1628
rect 1043 1624 1044 1628
rect 1038 1623 1044 1624
rect 1230 1628 1236 1629
rect 1230 1624 1231 1628
rect 1235 1624 1236 1628
rect 1230 1623 1236 1624
rect 1430 1628 1436 1629
rect 1430 1624 1431 1628
rect 1435 1624 1436 1628
rect 1430 1623 1436 1624
rect 1638 1628 1644 1629
rect 1638 1624 1639 1628
rect 1643 1624 1644 1628
rect 1766 1627 1767 1631
rect 1771 1627 1772 1631
rect 1766 1626 1772 1627
rect 1638 1623 1644 1624
rect 1883 1619 1889 1620
rect 1883 1615 1884 1619
rect 1888 1618 1889 1619
rect 1910 1619 1916 1620
rect 1910 1618 1911 1619
rect 1888 1616 1911 1618
rect 1888 1615 1889 1616
rect 1883 1614 1889 1615
rect 1910 1615 1911 1616
rect 1915 1615 1916 1619
rect 1910 1614 1916 1615
rect 1995 1619 2001 1620
rect 1995 1615 1996 1619
rect 2000 1618 2001 1619
rect 2022 1619 2028 1620
rect 2022 1618 2023 1619
rect 2000 1616 2023 1618
rect 2000 1615 2001 1616
rect 1995 1614 2001 1615
rect 2022 1615 2023 1616
rect 2027 1615 2028 1619
rect 2022 1614 2028 1615
rect 2139 1619 2145 1620
rect 2139 1615 2140 1619
rect 2144 1618 2145 1619
rect 2166 1619 2172 1620
rect 2166 1618 2167 1619
rect 2144 1616 2167 1618
rect 2144 1615 2145 1616
rect 2139 1614 2145 1615
rect 2166 1615 2167 1616
rect 2171 1615 2172 1619
rect 2166 1614 2172 1615
rect 2283 1619 2292 1620
rect 2283 1615 2284 1619
rect 2291 1615 2292 1619
rect 2283 1614 2292 1615
rect 2382 1619 2388 1620
rect 2382 1615 2383 1619
rect 2387 1618 2388 1619
rect 2419 1619 2425 1620
rect 2419 1618 2420 1619
rect 2387 1616 2420 1618
rect 2387 1615 2388 1616
rect 2382 1614 2388 1615
rect 2419 1615 2420 1616
rect 2424 1615 2425 1619
rect 2419 1614 2425 1615
rect 2555 1619 2564 1620
rect 2555 1615 2556 1619
rect 2563 1615 2564 1619
rect 2555 1614 2564 1615
rect 2615 1619 2621 1620
rect 2615 1615 2616 1619
rect 2620 1618 2621 1619
rect 2691 1619 2697 1620
rect 2691 1618 2692 1619
rect 2620 1616 2692 1618
rect 2620 1615 2621 1616
rect 2615 1614 2621 1615
rect 2691 1615 2692 1616
rect 2696 1615 2697 1619
rect 2691 1614 2697 1615
rect 2710 1619 2716 1620
rect 2710 1615 2711 1619
rect 2715 1618 2716 1619
rect 2819 1619 2825 1620
rect 2819 1618 2820 1619
rect 2715 1616 2820 1618
rect 2715 1615 2716 1616
rect 2710 1614 2716 1615
rect 2819 1615 2820 1616
rect 2824 1615 2825 1619
rect 2819 1614 2825 1615
rect 2838 1619 2844 1620
rect 2838 1615 2839 1619
rect 2843 1618 2844 1619
rect 2947 1619 2953 1620
rect 2947 1618 2948 1619
rect 2843 1616 2948 1618
rect 2843 1615 2844 1616
rect 2838 1614 2844 1615
rect 2947 1615 2948 1616
rect 2952 1615 2953 1619
rect 2947 1614 2953 1615
rect 2966 1619 2972 1620
rect 2966 1615 2967 1619
rect 2971 1618 2972 1619
rect 3067 1619 3073 1620
rect 3067 1618 3068 1619
rect 2971 1616 3068 1618
rect 2971 1615 2972 1616
rect 2966 1614 2972 1615
rect 3067 1615 3068 1616
rect 3072 1615 3073 1619
rect 3067 1614 3073 1615
rect 3186 1619 3193 1620
rect 3186 1615 3187 1619
rect 3192 1615 3193 1619
rect 3186 1614 3193 1615
rect 3206 1619 3212 1620
rect 3206 1615 3207 1619
rect 3211 1618 3212 1619
rect 3315 1619 3321 1620
rect 3315 1618 3316 1619
rect 3211 1616 3316 1618
rect 3211 1615 3212 1616
rect 3206 1614 3212 1615
rect 3315 1615 3316 1616
rect 3320 1615 3321 1619
rect 3315 1614 3321 1615
rect 3334 1619 3340 1620
rect 3334 1615 3335 1619
rect 3339 1618 3340 1619
rect 3419 1619 3425 1620
rect 3419 1618 3420 1619
rect 3339 1616 3420 1618
rect 3339 1615 3340 1616
rect 3334 1614 3340 1615
rect 3419 1615 3420 1616
rect 3424 1615 3425 1619
rect 3419 1614 3425 1615
rect 243 1611 252 1612
rect 243 1607 244 1611
rect 251 1607 252 1611
rect 243 1606 252 1607
rect 262 1611 268 1612
rect 262 1607 263 1611
rect 267 1610 268 1611
rect 347 1611 353 1612
rect 347 1610 348 1611
rect 267 1608 348 1610
rect 267 1607 268 1608
rect 262 1606 268 1607
rect 347 1607 348 1608
rect 352 1607 353 1611
rect 347 1606 353 1607
rect 366 1611 372 1612
rect 366 1607 367 1611
rect 371 1610 372 1611
rect 459 1611 465 1612
rect 459 1610 460 1611
rect 371 1608 460 1610
rect 371 1607 372 1608
rect 366 1606 372 1607
rect 459 1607 460 1608
rect 464 1607 465 1611
rect 459 1606 465 1607
rect 587 1611 593 1612
rect 587 1607 588 1611
rect 592 1610 593 1611
rect 614 1611 620 1612
rect 614 1610 615 1611
rect 592 1608 615 1610
rect 592 1607 593 1608
rect 587 1606 593 1607
rect 614 1607 615 1608
rect 619 1607 620 1611
rect 614 1606 620 1607
rect 722 1611 728 1612
rect 722 1607 723 1611
rect 727 1610 728 1611
rect 739 1611 745 1612
rect 739 1610 740 1611
rect 727 1608 740 1610
rect 727 1607 728 1608
rect 722 1606 728 1607
rect 739 1607 740 1608
rect 744 1607 745 1611
rect 739 1606 745 1607
rect 907 1611 916 1612
rect 907 1607 908 1611
rect 915 1607 916 1611
rect 907 1606 916 1607
rect 926 1611 932 1612
rect 926 1607 927 1611
rect 931 1610 932 1611
rect 1091 1611 1097 1612
rect 1091 1610 1092 1611
rect 931 1608 1092 1610
rect 931 1607 932 1608
rect 926 1606 932 1607
rect 1091 1607 1092 1608
rect 1096 1607 1097 1611
rect 1091 1606 1097 1607
rect 1110 1611 1116 1612
rect 1110 1607 1111 1611
rect 1115 1610 1116 1611
rect 1283 1611 1289 1612
rect 1283 1610 1284 1611
rect 1115 1608 1284 1610
rect 1115 1607 1116 1608
rect 1110 1606 1116 1607
rect 1283 1607 1284 1608
rect 1288 1607 1289 1611
rect 1283 1606 1289 1607
rect 1483 1611 1489 1612
rect 1483 1607 1484 1611
rect 1488 1610 1489 1611
rect 1510 1611 1516 1612
rect 1510 1610 1511 1611
rect 1488 1608 1511 1610
rect 1488 1607 1489 1608
rect 1483 1606 1489 1607
rect 1510 1607 1511 1608
rect 1515 1607 1516 1611
rect 1510 1606 1516 1607
rect 1691 1611 1697 1612
rect 1691 1607 1692 1611
rect 1696 1610 1697 1611
rect 1734 1611 1740 1612
rect 1734 1610 1735 1611
rect 1696 1608 1735 1610
rect 1696 1607 1697 1608
rect 1691 1606 1697 1607
rect 1734 1607 1735 1608
rect 1739 1607 1740 1611
rect 1734 1606 1740 1607
rect 1830 1604 1836 1605
rect 1806 1601 1812 1602
rect 1806 1597 1807 1601
rect 1811 1597 1812 1601
rect 1830 1600 1831 1604
rect 1835 1600 1836 1604
rect 1830 1599 1836 1600
rect 1942 1604 1948 1605
rect 1942 1600 1943 1604
rect 1947 1600 1948 1604
rect 1942 1599 1948 1600
rect 2086 1604 2092 1605
rect 2086 1600 2087 1604
rect 2091 1600 2092 1604
rect 2086 1599 2092 1600
rect 2230 1604 2236 1605
rect 2230 1600 2231 1604
rect 2235 1600 2236 1604
rect 2230 1599 2236 1600
rect 2366 1604 2372 1605
rect 2366 1600 2367 1604
rect 2371 1600 2372 1604
rect 2366 1599 2372 1600
rect 2502 1604 2508 1605
rect 2502 1600 2503 1604
rect 2507 1600 2508 1604
rect 2502 1599 2508 1600
rect 2638 1604 2644 1605
rect 2638 1600 2639 1604
rect 2643 1600 2644 1604
rect 2638 1599 2644 1600
rect 2766 1604 2772 1605
rect 2766 1600 2767 1604
rect 2771 1600 2772 1604
rect 2766 1599 2772 1600
rect 2894 1604 2900 1605
rect 2894 1600 2895 1604
rect 2899 1600 2900 1604
rect 2894 1599 2900 1600
rect 3014 1604 3020 1605
rect 3014 1600 3015 1604
rect 3019 1600 3020 1604
rect 3014 1599 3020 1600
rect 3134 1604 3140 1605
rect 3134 1600 3135 1604
rect 3139 1600 3140 1604
rect 3134 1599 3140 1600
rect 3262 1604 3268 1605
rect 3262 1600 3263 1604
rect 3267 1600 3268 1604
rect 3262 1599 3268 1600
rect 3366 1604 3372 1605
rect 3366 1600 3367 1604
rect 3371 1600 3372 1604
rect 3366 1599 3372 1600
rect 3462 1601 3468 1602
rect 1806 1596 1812 1597
rect 3462 1597 3463 1601
rect 3467 1597 3468 1601
rect 3462 1596 3468 1597
rect 379 1595 385 1596
rect 379 1591 380 1595
rect 384 1594 385 1595
rect 407 1595 413 1596
rect 407 1594 408 1595
rect 384 1592 408 1594
rect 384 1591 385 1592
rect 379 1590 385 1591
rect 407 1591 408 1592
rect 412 1591 413 1595
rect 407 1590 413 1591
rect 462 1595 468 1596
rect 462 1591 463 1595
rect 467 1594 468 1595
rect 483 1595 489 1596
rect 483 1594 484 1595
rect 467 1592 484 1594
rect 467 1591 468 1592
rect 462 1590 468 1591
rect 483 1591 484 1592
rect 488 1591 489 1595
rect 483 1590 489 1591
rect 595 1595 601 1596
rect 595 1591 596 1595
rect 600 1594 601 1595
rect 606 1595 612 1596
rect 606 1594 607 1595
rect 600 1592 607 1594
rect 600 1591 601 1592
rect 595 1590 601 1591
rect 606 1591 607 1592
rect 611 1591 612 1595
rect 606 1590 612 1591
rect 614 1595 620 1596
rect 614 1591 615 1595
rect 619 1594 620 1595
rect 723 1595 729 1596
rect 723 1594 724 1595
rect 619 1592 724 1594
rect 619 1591 620 1592
rect 614 1590 620 1591
rect 723 1591 724 1592
rect 728 1591 729 1595
rect 723 1590 729 1591
rect 742 1595 748 1596
rect 742 1591 743 1595
rect 747 1594 748 1595
rect 867 1595 873 1596
rect 867 1594 868 1595
rect 747 1592 868 1594
rect 747 1591 748 1592
rect 742 1590 748 1591
rect 867 1591 868 1592
rect 872 1591 873 1595
rect 867 1590 873 1591
rect 1019 1595 1025 1596
rect 1019 1591 1020 1595
rect 1024 1594 1025 1595
rect 1047 1595 1053 1596
rect 1047 1594 1048 1595
rect 1024 1592 1048 1594
rect 1024 1591 1025 1592
rect 1019 1590 1025 1591
rect 1047 1591 1048 1592
rect 1052 1591 1053 1595
rect 1047 1590 1053 1591
rect 1171 1595 1177 1596
rect 1171 1591 1172 1595
rect 1176 1594 1177 1595
rect 1190 1595 1196 1596
rect 1190 1594 1191 1595
rect 1176 1592 1191 1594
rect 1176 1591 1177 1592
rect 1171 1590 1177 1591
rect 1190 1591 1191 1592
rect 1195 1591 1196 1595
rect 1190 1590 1196 1591
rect 1331 1595 1337 1596
rect 1331 1591 1332 1595
rect 1336 1594 1337 1595
rect 1491 1595 1497 1596
rect 1336 1592 1430 1594
rect 1336 1591 1337 1592
rect 1331 1590 1337 1591
rect 1428 1586 1430 1592
rect 1491 1591 1492 1595
rect 1496 1594 1497 1595
rect 1502 1595 1508 1596
rect 1502 1594 1503 1595
rect 1496 1592 1503 1594
rect 1496 1591 1497 1592
rect 1491 1590 1497 1591
rect 1502 1591 1503 1592
rect 1507 1591 1508 1595
rect 1502 1590 1508 1591
rect 1510 1595 1516 1596
rect 1510 1591 1511 1595
rect 1515 1594 1516 1595
rect 1659 1595 1665 1596
rect 1659 1594 1660 1595
rect 1515 1592 1660 1594
rect 1515 1591 1516 1592
rect 1510 1590 1516 1591
rect 1659 1591 1660 1592
rect 1664 1591 1665 1595
rect 1659 1590 1665 1591
rect 1894 1595 1900 1596
rect 1894 1591 1895 1595
rect 1899 1591 1900 1595
rect 1894 1590 1900 1591
rect 1910 1595 1916 1596
rect 1910 1591 1911 1595
rect 1915 1594 1916 1595
rect 2022 1595 2028 1596
rect 1915 1592 1985 1594
rect 1915 1591 1916 1592
rect 1910 1590 1916 1591
rect 2022 1591 2023 1595
rect 2027 1594 2028 1595
rect 2166 1595 2172 1596
rect 2027 1592 2129 1594
rect 2027 1591 2028 1592
rect 2022 1590 2028 1591
rect 2166 1591 2167 1595
rect 2171 1594 2172 1595
rect 2438 1595 2444 1596
rect 2171 1592 2273 1594
rect 2171 1591 2172 1592
rect 2166 1590 2172 1591
rect 2438 1591 2439 1595
rect 2443 1591 2444 1595
rect 2615 1595 2621 1596
rect 2615 1594 2616 1595
rect 2577 1592 2616 1594
rect 2438 1590 2444 1591
rect 2615 1591 2616 1592
rect 2620 1591 2621 1595
rect 2615 1590 2621 1591
rect 2710 1595 2716 1596
rect 2710 1591 2711 1595
rect 2715 1591 2716 1595
rect 2710 1590 2716 1591
rect 2838 1595 2844 1596
rect 2838 1591 2839 1595
rect 2843 1591 2844 1595
rect 2838 1590 2844 1591
rect 2966 1595 2972 1596
rect 2966 1591 2967 1595
rect 2971 1591 2972 1595
rect 2966 1590 2972 1591
rect 3086 1595 3092 1596
rect 3086 1591 3087 1595
rect 3091 1591 3092 1595
rect 3086 1590 3092 1591
rect 3206 1595 3212 1596
rect 3206 1591 3207 1595
rect 3211 1591 3212 1595
rect 3206 1590 3212 1591
rect 3334 1595 3340 1596
rect 3334 1591 3335 1595
rect 3339 1591 3340 1595
rect 3334 1590 3340 1591
rect 3430 1595 3436 1596
rect 3430 1591 3431 1595
rect 3435 1591 3436 1595
rect 3430 1590 3436 1591
rect 1428 1584 1586 1586
rect 1830 1585 1836 1586
rect 326 1580 332 1581
rect 110 1577 116 1578
rect 110 1573 111 1577
rect 115 1573 116 1577
rect 326 1576 327 1580
rect 331 1576 332 1580
rect 326 1575 332 1576
rect 430 1580 436 1581
rect 430 1576 431 1580
rect 435 1576 436 1580
rect 430 1575 436 1576
rect 542 1580 548 1581
rect 542 1576 543 1580
rect 547 1576 548 1580
rect 542 1575 548 1576
rect 670 1580 676 1581
rect 670 1576 671 1580
rect 675 1576 676 1580
rect 670 1575 676 1576
rect 814 1580 820 1581
rect 814 1576 815 1580
rect 819 1576 820 1580
rect 814 1575 820 1576
rect 966 1580 972 1581
rect 966 1576 967 1580
rect 971 1576 972 1580
rect 966 1575 972 1576
rect 1118 1580 1124 1581
rect 1118 1576 1119 1580
rect 1123 1576 1124 1580
rect 1118 1575 1124 1576
rect 1278 1580 1284 1581
rect 1278 1576 1279 1580
rect 1283 1576 1284 1580
rect 1278 1575 1284 1576
rect 1438 1580 1444 1581
rect 1438 1576 1439 1580
rect 1443 1576 1444 1580
rect 1438 1575 1444 1576
rect 110 1572 116 1573
rect 246 1571 252 1572
rect 246 1567 247 1571
rect 251 1570 252 1571
rect 407 1571 413 1572
rect 251 1568 369 1570
rect 251 1567 252 1568
rect 246 1566 252 1567
rect 407 1567 408 1571
rect 412 1570 413 1571
rect 614 1571 620 1572
rect 412 1568 473 1570
rect 412 1567 413 1568
rect 407 1566 413 1567
rect 614 1567 615 1571
rect 619 1567 620 1571
rect 614 1566 620 1567
rect 742 1571 748 1572
rect 742 1567 743 1571
rect 747 1567 748 1571
rect 742 1566 748 1567
rect 806 1571 812 1572
rect 806 1567 807 1571
rect 811 1570 812 1571
rect 910 1571 916 1572
rect 811 1568 857 1570
rect 811 1567 812 1568
rect 806 1566 812 1567
rect 910 1567 911 1571
rect 915 1570 916 1571
rect 1047 1571 1053 1572
rect 915 1568 1009 1570
rect 915 1567 916 1568
rect 910 1566 916 1567
rect 1047 1567 1048 1571
rect 1052 1570 1053 1571
rect 1362 1571 1368 1572
rect 1362 1570 1363 1571
rect 1052 1568 1161 1570
rect 1353 1568 1363 1570
rect 1052 1567 1053 1568
rect 1047 1566 1053 1567
rect 1362 1567 1363 1568
rect 1367 1567 1368 1571
rect 1362 1566 1368 1567
rect 1510 1571 1516 1572
rect 1510 1567 1511 1571
rect 1515 1567 1516 1571
rect 1584 1570 1586 1584
rect 1806 1584 1812 1585
rect 1606 1580 1612 1581
rect 1606 1576 1607 1580
rect 1611 1576 1612 1580
rect 1806 1580 1807 1584
rect 1811 1580 1812 1584
rect 1830 1581 1831 1585
rect 1835 1581 1836 1585
rect 1830 1580 1836 1581
rect 1942 1585 1948 1586
rect 1942 1581 1943 1585
rect 1947 1581 1948 1585
rect 1942 1580 1948 1581
rect 2086 1585 2092 1586
rect 2086 1581 2087 1585
rect 2091 1581 2092 1585
rect 2086 1580 2092 1581
rect 2230 1585 2236 1586
rect 2230 1581 2231 1585
rect 2235 1581 2236 1585
rect 2230 1580 2236 1581
rect 2366 1585 2372 1586
rect 2366 1581 2367 1585
rect 2371 1581 2372 1585
rect 2366 1580 2372 1581
rect 2502 1585 2508 1586
rect 2502 1581 2503 1585
rect 2507 1581 2508 1585
rect 2502 1580 2508 1581
rect 2638 1585 2644 1586
rect 2638 1581 2639 1585
rect 2643 1581 2644 1585
rect 2638 1580 2644 1581
rect 2766 1585 2772 1586
rect 2766 1581 2767 1585
rect 2771 1581 2772 1585
rect 2766 1580 2772 1581
rect 2894 1585 2900 1586
rect 2894 1581 2895 1585
rect 2899 1581 2900 1585
rect 2894 1580 2900 1581
rect 3014 1585 3020 1586
rect 3014 1581 3015 1585
rect 3019 1581 3020 1585
rect 3014 1580 3020 1581
rect 3134 1585 3140 1586
rect 3134 1581 3135 1585
rect 3139 1581 3140 1585
rect 3134 1580 3140 1581
rect 3262 1585 3268 1586
rect 3262 1581 3263 1585
rect 3267 1581 3268 1585
rect 3262 1580 3268 1581
rect 3366 1585 3372 1586
rect 3366 1581 3367 1585
rect 3371 1581 3372 1585
rect 3366 1580 3372 1581
rect 3462 1584 3468 1585
rect 3462 1580 3463 1584
rect 3467 1580 3468 1584
rect 1806 1579 1812 1580
rect 3462 1579 3468 1580
rect 1606 1575 1612 1576
rect 1766 1577 1772 1578
rect 1766 1573 1767 1577
rect 1771 1573 1772 1577
rect 1766 1572 1772 1573
rect 1584 1568 1649 1570
rect 1510 1566 1516 1567
rect 326 1561 332 1562
rect 110 1560 116 1561
rect 110 1556 111 1560
rect 115 1556 116 1560
rect 326 1557 327 1561
rect 331 1557 332 1561
rect 326 1556 332 1557
rect 430 1561 436 1562
rect 430 1557 431 1561
rect 435 1557 436 1561
rect 430 1556 436 1557
rect 542 1561 548 1562
rect 542 1557 543 1561
rect 547 1557 548 1561
rect 542 1556 548 1557
rect 670 1561 676 1562
rect 670 1557 671 1561
rect 675 1557 676 1561
rect 670 1556 676 1557
rect 814 1561 820 1562
rect 814 1557 815 1561
rect 819 1557 820 1561
rect 814 1556 820 1557
rect 966 1561 972 1562
rect 966 1557 967 1561
rect 971 1557 972 1561
rect 966 1556 972 1557
rect 1118 1561 1124 1562
rect 1118 1557 1119 1561
rect 1123 1557 1124 1561
rect 1118 1556 1124 1557
rect 1278 1561 1284 1562
rect 1278 1557 1279 1561
rect 1283 1557 1284 1561
rect 1278 1556 1284 1557
rect 1438 1561 1444 1562
rect 1438 1557 1439 1561
rect 1443 1557 1444 1561
rect 1438 1556 1444 1557
rect 1606 1561 1612 1562
rect 1606 1557 1607 1561
rect 1611 1557 1612 1561
rect 1606 1556 1612 1557
rect 1766 1560 1772 1561
rect 1766 1556 1767 1560
rect 1771 1556 1772 1560
rect 110 1555 116 1556
rect 1766 1555 1772 1556
rect 1806 1532 1812 1533
rect 3462 1532 3468 1533
rect 1806 1528 1807 1532
rect 1811 1528 1812 1532
rect 1806 1527 1812 1528
rect 1838 1531 1844 1532
rect 1838 1527 1839 1531
rect 1843 1527 1844 1531
rect 1838 1526 1844 1527
rect 1990 1531 1996 1532
rect 1990 1527 1991 1531
rect 1995 1527 1996 1531
rect 1990 1526 1996 1527
rect 2150 1531 2156 1532
rect 2150 1527 2151 1531
rect 2155 1527 2156 1531
rect 2150 1526 2156 1527
rect 2302 1531 2308 1532
rect 2302 1527 2303 1531
rect 2307 1527 2308 1531
rect 2302 1526 2308 1527
rect 2454 1531 2460 1532
rect 2454 1527 2455 1531
rect 2459 1527 2460 1531
rect 2454 1526 2460 1527
rect 2598 1531 2604 1532
rect 2598 1527 2599 1531
rect 2603 1527 2604 1531
rect 2598 1526 2604 1527
rect 2734 1531 2740 1532
rect 2734 1527 2735 1531
rect 2739 1527 2740 1531
rect 2734 1526 2740 1527
rect 2870 1531 2876 1532
rect 2870 1527 2871 1531
rect 2875 1527 2876 1531
rect 2870 1526 2876 1527
rect 3006 1531 3012 1532
rect 3006 1527 3007 1531
rect 3011 1527 3012 1531
rect 3006 1526 3012 1527
rect 3142 1531 3148 1532
rect 3142 1527 3143 1531
rect 3147 1527 3148 1531
rect 3462 1528 3463 1532
rect 3467 1528 3468 1532
rect 3462 1527 3468 1528
rect 3142 1526 3148 1527
rect 2286 1523 2292 1524
rect 1910 1519 1916 1520
rect 1806 1515 1812 1516
rect 110 1512 116 1513
rect 1766 1512 1772 1513
rect 110 1508 111 1512
rect 115 1508 116 1512
rect 110 1507 116 1508
rect 222 1511 228 1512
rect 222 1507 223 1511
rect 227 1507 228 1511
rect 222 1506 228 1507
rect 342 1511 348 1512
rect 342 1507 343 1511
rect 347 1507 348 1511
rect 342 1506 348 1507
rect 470 1511 476 1512
rect 470 1507 471 1511
rect 475 1507 476 1511
rect 470 1506 476 1507
rect 606 1511 612 1512
rect 606 1507 607 1511
rect 611 1507 612 1511
rect 606 1506 612 1507
rect 750 1511 756 1512
rect 750 1507 751 1511
rect 755 1507 756 1511
rect 750 1506 756 1507
rect 894 1511 900 1512
rect 894 1507 895 1511
rect 899 1507 900 1511
rect 894 1506 900 1507
rect 1046 1511 1052 1512
rect 1046 1507 1047 1511
rect 1051 1507 1052 1511
rect 1046 1506 1052 1507
rect 1198 1511 1204 1512
rect 1198 1507 1199 1511
rect 1203 1507 1204 1511
rect 1198 1506 1204 1507
rect 1350 1511 1356 1512
rect 1350 1507 1351 1511
rect 1355 1507 1356 1511
rect 1350 1506 1356 1507
rect 1502 1511 1508 1512
rect 1502 1507 1503 1511
rect 1507 1507 1508 1511
rect 1766 1508 1767 1512
rect 1771 1508 1772 1512
rect 1806 1511 1807 1515
rect 1811 1511 1812 1515
rect 1910 1515 1911 1519
rect 1915 1515 1916 1519
rect 1910 1514 1916 1515
rect 2062 1519 2068 1520
rect 2062 1515 2063 1519
rect 2067 1515 2068 1519
rect 2062 1514 2068 1515
rect 2222 1519 2228 1520
rect 2222 1515 2223 1519
rect 2227 1515 2228 1519
rect 2286 1519 2287 1523
rect 2291 1522 2292 1523
rect 2558 1523 2564 1524
rect 2291 1520 2345 1522
rect 2291 1519 2292 1520
rect 2286 1518 2292 1519
rect 2550 1519 2556 1520
rect 2550 1518 2551 1519
rect 2529 1516 2551 1518
rect 2222 1514 2228 1515
rect 2550 1515 2551 1516
rect 2555 1515 2556 1519
rect 2558 1519 2559 1523
rect 2563 1522 2564 1523
rect 2678 1523 2684 1524
rect 2563 1520 2641 1522
rect 2563 1519 2564 1520
rect 2558 1518 2564 1519
rect 2678 1519 2679 1523
rect 2683 1522 2684 1523
rect 2814 1523 2820 1524
rect 2683 1520 2777 1522
rect 2683 1519 2684 1520
rect 2678 1518 2684 1519
rect 2814 1519 2815 1523
rect 2819 1522 2820 1523
rect 2950 1523 2956 1524
rect 2819 1520 2913 1522
rect 2819 1519 2820 1520
rect 2814 1518 2820 1519
rect 2950 1519 2951 1523
rect 2955 1522 2956 1523
rect 3086 1523 3092 1524
rect 2955 1520 3049 1522
rect 2955 1519 2956 1520
rect 2950 1518 2956 1519
rect 3086 1519 3087 1523
rect 3091 1522 3092 1523
rect 3091 1520 3185 1522
rect 3091 1519 3092 1520
rect 3086 1518 3092 1519
rect 2550 1514 2556 1515
rect 3462 1515 3468 1516
rect 1806 1510 1812 1511
rect 1838 1512 1844 1513
rect 1766 1507 1772 1508
rect 1838 1508 1839 1512
rect 1843 1508 1844 1512
rect 1838 1507 1844 1508
rect 1990 1512 1996 1513
rect 1990 1508 1991 1512
rect 1995 1508 1996 1512
rect 1990 1507 1996 1508
rect 2150 1512 2156 1513
rect 2150 1508 2151 1512
rect 2155 1508 2156 1512
rect 2150 1507 2156 1508
rect 2302 1512 2308 1513
rect 2302 1508 2303 1512
rect 2307 1508 2308 1512
rect 2302 1507 2308 1508
rect 2454 1512 2460 1513
rect 2454 1508 2455 1512
rect 2459 1508 2460 1512
rect 2454 1507 2460 1508
rect 2598 1512 2604 1513
rect 2598 1508 2599 1512
rect 2603 1508 2604 1512
rect 2598 1507 2604 1508
rect 2734 1512 2740 1513
rect 2734 1508 2735 1512
rect 2739 1508 2740 1512
rect 2734 1507 2740 1508
rect 2870 1512 2876 1513
rect 2870 1508 2871 1512
rect 2875 1508 2876 1512
rect 2870 1507 2876 1508
rect 3006 1512 3012 1513
rect 3006 1508 3007 1512
rect 3011 1508 3012 1512
rect 3006 1507 3012 1508
rect 3142 1512 3148 1513
rect 3142 1508 3143 1512
rect 3147 1508 3148 1512
rect 3462 1511 3463 1515
rect 3467 1511 3468 1515
rect 3462 1510 3468 1511
rect 3142 1507 3148 1508
rect 1502 1506 1508 1507
rect 462 1503 468 1504
rect 294 1499 300 1500
rect 110 1495 116 1496
rect 110 1491 111 1495
rect 115 1491 116 1495
rect 294 1495 295 1499
rect 299 1495 300 1499
rect 294 1494 300 1495
rect 414 1499 420 1500
rect 414 1495 415 1499
rect 419 1495 420 1499
rect 462 1499 463 1503
rect 467 1502 468 1503
rect 550 1503 556 1504
rect 467 1500 513 1502
rect 467 1499 468 1500
rect 462 1498 468 1499
rect 550 1499 551 1503
rect 555 1502 556 1503
rect 735 1503 741 1504
rect 555 1500 649 1502
rect 555 1499 556 1500
rect 550 1498 556 1499
rect 735 1499 736 1503
rect 740 1502 741 1503
rect 1190 1503 1196 1504
rect 740 1500 793 1502
rect 740 1499 741 1500
rect 735 1498 741 1499
rect 966 1499 972 1500
rect 414 1494 420 1495
rect 966 1495 967 1499
rect 971 1495 972 1499
rect 966 1494 972 1495
rect 1118 1499 1124 1500
rect 1118 1495 1119 1499
rect 1123 1495 1124 1499
rect 1190 1499 1191 1503
rect 1195 1502 1196 1503
rect 1195 1500 1241 1502
rect 1195 1499 1196 1500
rect 1190 1498 1196 1499
rect 1422 1499 1428 1500
rect 1118 1494 1124 1495
rect 1422 1495 1423 1499
rect 1427 1495 1428 1499
rect 1422 1494 1428 1495
rect 1574 1499 1580 1500
rect 1574 1495 1575 1499
rect 1579 1495 1580 1499
rect 1574 1494 1580 1495
rect 1766 1495 1772 1496
rect 110 1490 116 1491
rect 222 1492 228 1493
rect 222 1488 223 1492
rect 227 1488 228 1492
rect 222 1487 228 1488
rect 342 1492 348 1493
rect 342 1488 343 1492
rect 347 1488 348 1492
rect 342 1487 348 1488
rect 470 1492 476 1493
rect 470 1488 471 1492
rect 475 1488 476 1492
rect 470 1487 476 1488
rect 606 1492 612 1493
rect 606 1488 607 1492
rect 611 1488 612 1492
rect 606 1487 612 1488
rect 750 1492 756 1493
rect 750 1488 751 1492
rect 755 1488 756 1492
rect 750 1487 756 1488
rect 894 1492 900 1493
rect 894 1488 895 1492
rect 899 1488 900 1492
rect 894 1487 900 1488
rect 1046 1492 1052 1493
rect 1046 1488 1047 1492
rect 1051 1488 1052 1492
rect 1046 1487 1052 1488
rect 1198 1492 1204 1493
rect 1198 1488 1199 1492
rect 1203 1488 1204 1492
rect 1198 1487 1204 1488
rect 1350 1492 1356 1493
rect 1350 1488 1351 1492
rect 1355 1488 1356 1492
rect 1350 1487 1356 1488
rect 1502 1492 1508 1493
rect 1502 1488 1503 1492
rect 1507 1488 1508 1492
rect 1766 1491 1767 1495
rect 1771 1491 1772 1495
rect 1766 1490 1772 1491
rect 1891 1495 1900 1496
rect 1891 1491 1892 1495
rect 1899 1491 1900 1495
rect 1891 1490 1900 1491
rect 1910 1495 1916 1496
rect 1910 1491 1911 1495
rect 1915 1494 1916 1495
rect 2043 1495 2049 1496
rect 2043 1494 2044 1495
rect 1915 1492 2044 1494
rect 1915 1491 1916 1492
rect 1910 1490 1916 1491
rect 2043 1491 2044 1492
rect 2048 1491 2049 1495
rect 2043 1490 2049 1491
rect 2062 1495 2068 1496
rect 2062 1491 2063 1495
rect 2067 1494 2068 1495
rect 2203 1495 2209 1496
rect 2203 1494 2204 1495
rect 2067 1492 2204 1494
rect 2067 1491 2068 1492
rect 2062 1490 2068 1491
rect 2203 1491 2204 1492
rect 2208 1491 2209 1495
rect 2203 1490 2209 1491
rect 2222 1495 2228 1496
rect 2222 1491 2223 1495
rect 2227 1494 2228 1495
rect 2355 1495 2361 1496
rect 2355 1494 2356 1495
rect 2227 1492 2356 1494
rect 2227 1491 2228 1492
rect 2222 1490 2228 1491
rect 2355 1491 2356 1492
rect 2360 1491 2361 1495
rect 2355 1490 2361 1491
rect 2438 1495 2444 1496
rect 2438 1491 2439 1495
rect 2443 1494 2444 1495
rect 2507 1495 2513 1496
rect 2507 1494 2508 1495
rect 2443 1492 2508 1494
rect 2443 1491 2444 1492
rect 2438 1490 2444 1491
rect 2507 1491 2508 1492
rect 2512 1491 2513 1495
rect 2507 1490 2513 1491
rect 2651 1495 2657 1496
rect 2651 1491 2652 1495
rect 2656 1494 2657 1495
rect 2678 1495 2684 1496
rect 2678 1494 2679 1495
rect 2656 1492 2679 1494
rect 2656 1491 2657 1492
rect 2651 1490 2657 1491
rect 2678 1491 2679 1492
rect 2683 1491 2684 1495
rect 2678 1490 2684 1491
rect 2787 1495 2793 1496
rect 2787 1491 2788 1495
rect 2792 1494 2793 1495
rect 2814 1495 2820 1496
rect 2814 1494 2815 1495
rect 2792 1492 2815 1494
rect 2792 1491 2793 1492
rect 2787 1490 2793 1491
rect 2814 1491 2815 1492
rect 2819 1491 2820 1495
rect 2814 1490 2820 1491
rect 2923 1495 2929 1496
rect 2923 1491 2924 1495
rect 2928 1494 2929 1495
rect 2950 1495 2956 1496
rect 2950 1494 2951 1495
rect 2928 1492 2951 1494
rect 2928 1491 2929 1492
rect 2923 1490 2929 1491
rect 2950 1491 2951 1492
rect 2955 1491 2956 1495
rect 2950 1490 2956 1491
rect 3059 1495 3065 1496
rect 3059 1491 3060 1495
rect 3064 1494 3065 1495
rect 3086 1495 3092 1496
rect 3086 1494 3087 1495
rect 3064 1492 3087 1494
rect 3064 1491 3065 1492
rect 3059 1490 3065 1491
rect 3086 1491 3087 1492
rect 3091 1491 3092 1495
rect 3086 1490 3092 1491
rect 3195 1495 3204 1496
rect 3195 1491 3196 1495
rect 3203 1491 3204 1495
rect 3195 1490 3204 1491
rect 1502 1487 1508 1488
rect 206 1475 212 1476
rect 206 1471 207 1475
rect 211 1474 212 1475
rect 275 1475 281 1476
rect 275 1474 276 1475
rect 211 1472 276 1474
rect 211 1471 212 1472
rect 206 1470 212 1471
rect 275 1471 276 1472
rect 280 1471 281 1475
rect 275 1470 281 1471
rect 294 1475 300 1476
rect 294 1471 295 1475
rect 299 1474 300 1475
rect 395 1475 401 1476
rect 395 1474 396 1475
rect 299 1472 396 1474
rect 299 1471 300 1472
rect 294 1470 300 1471
rect 395 1471 396 1472
rect 400 1471 401 1475
rect 395 1470 401 1471
rect 414 1475 420 1476
rect 414 1471 415 1475
rect 419 1474 420 1475
rect 523 1475 529 1476
rect 523 1474 524 1475
rect 419 1472 524 1474
rect 419 1471 420 1472
rect 414 1470 420 1471
rect 523 1471 524 1472
rect 528 1471 529 1475
rect 523 1470 529 1471
rect 659 1475 665 1476
rect 659 1471 660 1475
rect 664 1474 665 1475
rect 735 1475 741 1476
rect 735 1474 736 1475
rect 664 1472 736 1474
rect 664 1471 665 1472
rect 659 1470 665 1471
rect 735 1471 736 1472
rect 740 1471 741 1475
rect 735 1470 741 1471
rect 803 1475 812 1476
rect 803 1471 804 1475
rect 811 1471 812 1475
rect 803 1470 812 1471
rect 947 1475 953 1476
rect 947 1471 948 1475
rect 952 1474 953 1475
rect 966 1475 972 1476
rect 952 1472 962 1474
rect 952 1471 953 1472
rect 947 1470 953 1471
rect 960 1466 962 1472
rect 966 1471 967 1475
rect 971 1474 972 1475
rect 1099 1475 1105 1476
rect 1099 1474 1100 1475
rect 971 1472 1100 1474
rect 971 1471 972 1472
rect 966 1470 972 1471
rect 1099 1471 1100 1472
rect 1104 1471 1105 1475
rect 1099 1470 1105 1471
rect 1118 1475 1124 1476
rect 1118 1471 1119 1475
rect 1123 1474 1124 1475
rect 1251 1475 1257 1476
rect 1251 1474 1252 1475
rect 1123 1472 1252 1474
rect 1123 1471 1124 1472
rect 1118 1470 1124 1471
rect 1251 1471 1252 1472
rect 1256 1471 1257 1475
rect 1251 1470 1257 1471
rect 1362 1475 1368 1476
rect 1362 1471 1363 1475
rect 1367 1474 1368 1475
rect 1403 1475 1409 1476
rect 1403 1474 1404 1475
rect 1367 1472 1404 1474
rect 1367 1471 1368 1472
rect 1362 1470 1368 1471
rect 1403 1471 1404 1472
rect 1408 1471 1409 1475
rect 1403 1470 1409 1471
rect 1422 1475 1428 1476
rect 1422 1471 1423 1475
rect 1427 1474 1428 1475
rect 1555 1475 1561 1476
rect 1555 1474 1556 1475
rect 1427 1472 1556 1474
rect 1427 1471 1428 1472
rect 1422 1470 1428 1471
rect 1555 1471 1556 1472
rect 1560 1471 1561 1475
rect 1555 1470 1561 1471
rect 1995 1475 2001 1476
rect 1995 1471 1996 1475
rect 2000 1474 2001 1475
rect 2023 1475 2029 1476
rect 2023 1474 2024 1475
rect 2000 1472 2024 1474
rect 2000 1471 2001 1472
rect 1995 1470 2001 1471
rect 2023 1471 2024 1472
rect 2028 1471 2029 1475
rect 2023 1470 2029 1471
rect 2107 1475 2113 1476
rect 2107 1471 2108 1475
rect 2112 1474 2113 1475
rect 2134 1475 2140 1476
rect 2134 1474 2135 1475
rect 2112 1472 2135 1474
rect 2112 1471 2113 1472
rect 2107 1470 2113 1471
rect 2134 1471 2135 1472
rect 2139 1471 2140 1475
rect 2134 1470 2140 1471
rect 2243 1475 2249 1476
rect 2243 1471 2244 1475
rect 2248 1474 2249 1475
rect 2387 1475 2396 1476
rect 2248 1472 2361 1474
rect 2248 1471 2249 1472
rect 2243 1470 2249 1471
rect 1010 1467 1016 1468
rect 1010 1466 1011 1467
rect 960 1464 1011 1466
rect 1010 1463 1011 1464
rect 1015 1463 1016 1467
rect 2359 1466 2361 1472
rect 2387 1471 2388 1475
rect 2395 1471 2396 1475
rect 2387 1470 2396 1471
rect 2406 1475 2412 1476
rect 2406 1471 2407 1475
rect 2411 1474 2412 1475
rect 2531 1475 2537 1476
rect 2531 1474 2532 1475
rect 2411 1472 2532 1474
rect 2411 1471 2412 1472
rect 2406 1470 2412 1471
rect 2531 1471 2532 1472
rect 2536 1471 2537 1475
rect 2531 1470 2537 1471
rect 2550 1475 2556 1476
rect 2550 1471 2551 1475
rect 2555 1474 2556 1475
rect 2683 1475 2689 1476
rect 2683 1474 2684 1475
rect 2555 1472 2684 1474
rect 2555 1471 2556 1472
rect 2550 1470 2556 1471
rect 2683 1471 2684 1472
rect 2688 1471 2689 1475
rect 2683 1470 2689 1471
rect 2835 1475 2844 1476
rect 2835 1471 2836 1475
rect 2843 1471 2844 1475
rect 2835 1470 2844 1471
rect 2854 1475 2860 1476
rect 2854 1471 2855 1475
rect 2859 1474 2860 1475
rect 2987 1475 2993 1476
rect 2987 1474 2988 1475
rect 2859 1472 2988 1474
rect 2859 1471 2860 1472
rect 2854 1470 2860 1471
rect 2987 1471 2988 1472
rect 2992 1471 2993 1475
rect 2987 1470 2993 1471
rect 3055 1475 3061 1476
rect 3055 1471 3056 1475
rect 3060 1474 3061 1475
rect 3139 1475 3145 1476
rect 3139 1474 3140 1475
rect 3060 1472 3140 1474
rect 3060 1471 3061 1472
rect 3055 1470 3061 1471
rect 3139 1471 3140 1472
rect 3144 1471 3145 1475
rect 3139 1470 3145 1471
rect 3158 1475 3164 1476
rect 3158 1471 3159 1475
rect 3163 1474 3164 1475
rect 3291 1475 3297 1476
rect 3291 1474 3292 1475
rect 3163 1472 3292 1474
rect 3163 1471 3164 1472
rect 3158 1470 3164 1471
rect 3291 1471 3292 1472
rect 3296 1471 3297 1475
rect 3291 1470 3297 1471
rect 2359 1464 2418 1466
rect 1010 1462 1016 1463
rect 1942 1460 1948 1461
rect 1806 1457 1812 1458
rect 187 1455 193 1456
rect 187 1451 188 1455
rect 192 1454 193 1455
rect 215 1455 221 1456
rect 215 1454 216 1455
rect 192 1452 216 1454
rect 192 1451 193 1452
rect 187 1450 193 1451
rect 215 1451 216 1452
rect 220 1451 221 1455
rect 215 1450 221 1451
rect 355 1455 364 1456
rect 355 1451 356 1455
rect 363 1451 364 1455
rect 355 1450 364 1451
rect 523 1455 529 1456
rect 523 1451 524 1455
rect 528 1454 529 1455
rect 550 1455 556 1456
rect 550 1454 551 1455
rect 528 1452 551 1454
rect 528 1451 529 1452
rect 523 1450 529 1451
rect 550 1451 551 1452
rect 555 1451 556 1455
rect 550 1450 556 1451
rect 598 1455 604 1456
rect 598 1451 599 1455
rect 603 1454 604 1455
rect 683 1455 689 1456
rect 683 1454 684 1455
rect 603 1452 684 1454
rect 603 1451 604 1452
rect 598 1450 604 1451
rect 683 1451 684 1452
rect 688 1451 689 1455
rect 683 1450 689 1451
rect 702 1455 708 1456
rect 702 1451 703 1455
rect 707 1454 708 1455
rect 835 1455 841 1456
rect 835 1454 836 1455
rect 707 1452 836 1454
rect 707 1451 708 1452
rect 702 1450 708 1451
rect 835 1451 836 1452
rect 840 1451 841 1455
rect 835 1450 841 1451
rect 974 1455 985 1456
rect 974 1451 975 1455
rect 979 1451 980 1455
rect 984 1451 985 1455
rect 974 1450 985 1451
rect 998 1455 1004 1456
rect 998 1451 999 1455
rect 1003 1454 1004 1455
rect 1115 1455 1121 1456
rect 1115 1454 1116 1455
rect 1003 1452 1116 1454
rect 1003 1451 1004 1452
rect 998 1450 1004 1451
rect 1115 1451 1116 1452
rect 1120 1451 1121 1455
rect 1115 1450 1121 1451
rect 1251 1455 1257 1456
rect 1251 1451 1252 1455
rect 1256 1454 1257 1455
rect 1278 1455 1284 1456
rect 1278 1454 1279 1455
rect 1256 1452 1279 1454
rect 1256 1451 1257 1452
rect 1251 1450 1257 1451
rect 1278 1451 1279 1452
rect 1283 1451 1284 1455
rect 1278 1450 1284 1451
rect 1387 1455 1393 1456
rect 1387 1451 1388 1455
rect 1392 1454 1393 1455
rect 1414 1455 1420 1456
rect 1414 1454 1415 1455
rect 1392 1452 1415 1454
rect 1392 1451 1393 1452
rect 1387 1450 1393 1451
rect 1414 1451 1415 1452
rect 1419 1451 1420 1455
rect 1414 1450 1420 1451
rect 1523 1455 1529 1456
rect 1523 1451 1524 1455
rect 1528 1454 1529 1455
rect 1574 1455 1580 1456
rect 1574 1454 1575 1455
rect 1528 1452 1575 1454
rect 1528 1451 1529 1452
rect 1523 1450 1529 1451
rect 1574 1451 1575 1452
rect 1579 1451 1580 1455
rect 1806 1453 1807 1457
rect 1811 1453 1812 1457
rect 1942 1456 1943 1460
rect 1947 1456 1948 1460
rect 1942 1455 1948 1456
rect 2054 1460 2060 1461
rect 2054 1456 2055 1460
rect 2059 1456 2060 1460
rect 2054 1455 2060 1456
rect 2190 1460 2196 1461
rect 2190 1456 2191 1460
rect 2195 1456 2196 1460
rect 2190 1455 2196 1456
rect 2334 1460 2340 1461
rect 2334 1456 2335 1460
rect 2339 1456 2340 1460
rect 2334 1455 2340 1456
rect 1806 1452 1812 1453
rect 1574 1450 1580 1451
rect 1894 1451 1900 1452
rect 1894 1447 1895 1451
rect 1899 1450 1900 1451
rect 2023 1451 2029 1452
rect 1899 1448 1985 1450
rect 1899 1447 1900 1448
rect 1894 1446 1900 1447
rect 2023 1447 2024 1451
rect 2028 1450 2029 1451
rect 2134 1451 2140 1452
rect 2028 1448 2097 1450
rect 2028 1447 2029 1448
rect 2023 1446 2029 1447
rect 2134 1447 2135 1451
rect 2139 1450 2140 1451
rect 2406 1451 2412 1452
rect 2139 1448 2233 1450
rect 2139 1447 2140 1448
rect 2134 1446 2140 1447
rect 2406 1447 2407 1451
rect 2411 1447 2412 1451
rect 2416 1450 2418 1464
rect 2478 1460 2484 1461
rect 2478 1456 2479 1460
rect 2483 1456 2484 1460
rect 2478 1455 2484 1456
rect 2630 1460 2636 1461
rect 2630 1456 2631 1460
rect 2635 1456 2636 1460
rect 2630 1455 2636 1456
rect 2782 1460 2788 1461
rect 2782 1456 2783 1460
rect 2787 1456 2788 1460
rect 2782 1455 2788 1456
rect 2934 1460 2940 1461
rect 2934 1456 2935 1460
rect 2939 1456 2940 1460
rect 2934 1455 2940 1456
rect 3086 1460 3092 1461
rect 3086 1456 3087 1460
rect 3091 1456 3092 1460
rect 3086 1455 3092 1456
rect 3238 1460 3244 1461
rect 3238 1456 3239 1460
rect 3243 1456 3244 1460
rect 3238 1455 3244 1456
rect 3462 1457 3468 1458
rect 3462 1453 3463 1457
rect 3467 1453 3468 1457
rect 3462 1452 3468 1453
rect 2702 1451 2708 1452
rect 2416 1448 2521 1450
rect 2406 1446 2412 1447
rect 2702 1447 2703 1451
rect 2707 1447 2708 1451
rect 2702 1446 2708 1447
rect 2854 1451 2860 1452
rect 2854 1447 2855 1451
rect 2859 1447 2860 1451
rect 3055 1451 3061 1452
rect 3055 1450 3056 1451
rect 3009 1448 3056 1450
rect 2854 1446 2860 1447
rect 3055 1447 3056 1448
rect 3060 1447 3061 1451
rect 3055 1446 3061 1447
rect 3158 1451 3164 1452
rect 3158 1447 3159 1451
rect 3163 1447 3164 1451
rect 3158 1446 3164 1447
rect 3198 1451 3204 1452
rect 3198 1447 3199 1451
rect 3203 1450 3204 1451
rect 3203 1448 3281 1450
rect 3203 1447 3204 1448
rect 3198 1446 3204 1447
rect 1942 1441 1948 1442
rect 134 1440 140 1441
rect 110 1437 116 1438
rect 110 1433 111 1437
rect 115 1433 116 1437
rect 134 1436 135 1440
rect 139 1436 140 1440
rect 134 1435 140 1436
rect 302 1440 308 1441
rect 302 1436 303 1440
rect 307 1436 308 1440
rect 302 1435 308 1436
rect 470 1440 476 1441
rect 470 1436 471 1440
rect 475 1436 476 1440
rect 470 1435 476 1436
rect 630 1440 636 1441
rect 630 1436 631 1440
rect 635 1436 636 1440
rect 630 1435 636 1436
rect 782 1440 788 1441
rect 782 1436 783 1440
rect 787 1436 788 1440
rect 782 1435 788 1436
rect 926 1440 932 1441
rect 926 1436 927 1440
rect 931 1436 932 1440
rect 926 1435 932 1436
rect 1062 1440 1068 1441
rect 1062 1436 1063 1440
rect 1067 1436 1068 1440
rect 1062 1435 1068 1436
rect 1198 1440 1204 1441
rect 1198 1436 1199 1440
rect 1203 1436 1204 1440
rect 1198 1435 1204 1436
rect 1334 1440 1340 1441
rect 1334 1436 1335 1440
rect 1339 1436 1340 1440
rect 1334 1435 1340 1436
rect 1470 1440 1476 1441
rect 1470 1436 1471 1440
rect 1475 1436 1476 1440
rect 1806 1440 1812 1441
rect 1470 1435 1476 1436
rect 1766 1437 1772 1438
rect 110 1432 116 1433
rect 1766 1433 1767 1437
rect 1771 1433 1772 1437
rect 1806 1436 1807 1440
rect 1811 1436 1812 1440
rect 1942 1437 1943 1441
rect 1947 1437 1948 1441
rect 1942 1436 1948 1437
rect 2054 1441 2060 1442
rect 2054 1437 2055 1441
rect 2059 1437 2060 1441
rect 2054 1436 2060 1437
rect 2190 1441 2196 1442
rect 2190 1437 2191 1441
rect 2195 1437 2196 1441
rect 2190 1436 2196 1437
rect 2334 1441 2340 1442
rect 2334 1437 2335 1441
rect 2339 1437 2340 1441
rect 2334 1436 2340 1437
rect 2478 1441 2484 1442
rect 2478 1437 2479 1441
rect 2483 1437 2484 1441
rect 2478 1436 2484 1437
rect 2630 1441 2636 1442
rect 2630 1437 2631 1441
rect 2635 1437 2636 1441
rect 2630 1436 2636 1437
rect 2782 1441 2788 1442
rect 2782 1437 2783 1441
rect 2787 1437 2788 1441
rect 2782 1436 2788 1437
rect 2934 1441 2940 1442
rect 2934 1437 2935 1441
rect 2939 1437 2940 1441
rect 2934 1436 2940 1437
rect 3086 1441 3092 1442
rect 3086 1437 3087 1441
rect 3091 1437 3092 1441
rect 3086 1436 3092 1437
rect 3238 1441 3244 1442
rect 3238 1437 3239 1441
rect 3243 1437 3244 1441
rect 3238 1436 3244 1437
rect 3462 1440 3468 1441
rect 3462 1436 3463 1440
rect 3467 1436 3468 1440
rect 1806 1435 1812 1436
rect 3462 1435 3468 1436
rect 1766 1432 1772 1433
rect 206 1431 212 1432
rect 206 1427 207 1431
rect 211 1427 212 1431
rect 206 1426 212 1427
rect 215 1431 221 1432
rect 215 1427 216 1431
rect 220 1430 221 1431
rect 598 1431 604 1432
rect 598 1430 599 1431
rect 220 1428 345 1430
rect 545 1428 599 1430
rect 220 1427 221 1428
rect 215 1426 221 1427
rect 598 1427 599 1428
rect 603 1427 604 1431
rect 598 1426 604 1427
rect 702 1431 708 1432
rect 702 1427 703 1431
rect 707 1427 708 1431
rect 702 1426 708 1427
rect 846 1431 852 1432
rect 846 1427 847 1431
rect 851 1427 852 1431
rect 846 1426 852 1427
rect 998 1431 1004 1432
rect 998 1427 999 1431
rect 1003 1427 1004 1431
rect 998 1426 1004 1427
rect 1010 1431 1016 1432
rect 1010 1427 1011 1431
rect 1015 1430 1016 1431
rect 1270 1431 1276 1432
rect 1015 1428 1105 1430
rect 1015 1427 1016 1428
rect 1010 1426 1016 1427
rect 1270 1427 1271 1431
rect 1275 1427 1276 1431
rect 1270 1426 1276 1427
rect 1278 1431 1284 1432
rect 1278 1427 1279 1431
rect 1283 1430 1284 1431
rect 1414 1431 1420 1432
rect 1283 1428 1377 1430
rect 1283 1427 1284 1428
rect 1278 1426 1284 1427
rect 1414 1427 1415 1431
rect 1419 1430 1420 1431
rect 1419 1428 1513 1430
rect 1419 1427 1420 1428
rect 1414 1426 1420 1427
rect 134 1421 140 1422
rect 110 1420 116 1421
rect 110 1416 111 1420
rect 115 1416 116 1420
rect 134 1417 135 1421
rect 139 1417 140 1421
rect 134 1416 140 1417
rect 302 1421 308 1422
rect 302 1417 303 1421
rect 307 1417 308 1421
rect 302 1416 308 1417
rect 470 1421 476 1422
rect 470 1417 471 1421
rect 475 1417 476 1421
rect 470 1416 476 1417
rect 630 1421 636 1422
rect 630 1417 631 1421
rect 635 1417 636 1421
rect 630 1416 636 1417
rect 782 1421 788 1422
rect 782 1417 783 1421
rect 787 1417 788 1421
rect 782 1416 788 1417
rect 926 1421 932 1422
rect 926 1417 927 1421
rect 931 1417 932 1421
rect 926 1416 932 1417
rect 1062 1421 1068 1422
rect 1062 1417 1063 1421
rect 1067 1417 1068 1421
rect 1062 1416 1068 1417
rect 1198 1421 1204 1422
rect 1198 1417 1199 1421
rect 1203 1417 1204 1421
rect 1198 1416 1204 1417
rect 1334 1421 1340 1422
rect 1334 1417 1335 1421
rect 1339 1417 1340 1421
rect 1334 1416 1340 1417
rect 1470 1421 1476 1422
rect 1470 1417 1471 1421
rect 1475 1417 1476 1421
rect 1470 1416 1476 1417
rect 1766 1420 1772 1421
rect 1766 1416 1767 1420
rect 1771 1416 1772 1420
rect 110 1415 116 1416
rect 1766 1415 1772 1416
rect 1806 1388 1812 1389
rect 3462 1388 3468 1389
rect 1806 1384 1807 1388
rect 1811 1384 1812 1388
rect 1806 1383 1812 1384
rect 2094 1387 2100 1388
rect 2094 1383 2095 1387
rect 2099 1383 2100 1387
rect 2094 1382 2100 1383
rect 2198 1387 2204 1388
rect 2198 1383 2199 1387
rect 2203 1383 2204 1387
rect 2198 1382 2204 1383
rect 2318 1387 2324 1388
rect 2318 1383 2319 1387
rect 2323 1383 2324 1387
rect 2318 1382 2324 1383
rect 2454 1387 2460 1388
rect 2454 1383 2455 1387
rect 2459 1383 2460 1387
rect 2454 1382 2460 1383
rect 2598 1387 2604 1388
rect 2598 1383 2599 1387
rect 2603 1383 2604 1387
rect 2598 1382 2604 1383
rect 2742 1387 2748 1388
rect 2742 1383 2743 1387
rect 2747 1383 2748 1387
rect 2742 1382 2748 1383
rect 2886 1387 2892 1388
rect 2886 1383 2887 1387
rect 2891 1383 2892 1387
rect 2886 1382 2892 1383
rect 3030 1387 3036 1388
rect 3030 1383 3031 1387
rect 3035 1383 3036 1387
rect 3030 1382 3036 1383
rect 3174 1387 3180 1388
rect 3174 1383 3175 1387
rect 3179 1383 3180 1387
rect 3174 1382 3180 1383
rect 3326 1387 3332 1388
rect 3326 1383 3327 1387
rect 3331 1383 3332 1387
rect 3462 1384 3463 1388
rect 3467 1384 3468 1388
rect 3462 1383 3468 1384
rect 3326 1382 3332 1383
rect 2390 1379 2396 1380
rect 2166 1375 2172 1376
rect 110 1372 116 1373
rect 1766 1372 1772 1373
rect 110 1368 111 1372
rect 115 1368 116 1372
rect 110 1367 116 1368
rect 134 1371 140 1372
rect 134 1367 135 1371
rect 139 1367 140 1371
rect 134 1366 140 1367
rect 278 1371 284 1372
rect 278 1367 279 1371
rect 283 1367 284 1371
rect 278 1366 284 1367
rect 446 1371 452 1372
rect 446 1367 447 1371
rect 451 1367 452 1371
rect 446 1366 452 1367
rect 606 1371 612 1372
rect 606 1367 607 1371
rect 611 1367 612 1371
rect 606 1366 612 1367
rect 758 1371 764 1372
rect 758 1367 759 1371
rect 763 1367 764 1371
rect 758 1366 764 1367
rect 902 1371 908 1372
rect 902 1367 903 1371
rect 907 1367 908 1371
rect 902 1366 908 1367
rect 1030 1371 1036 1372
rect 1030 1367 1031 1371
rect 1035 1367 1036 1371
rect 1030 1366 1036 1367
rect 1158 1371 1164 1372
rect 1158 1367 1159 1371
rect 1163 1367 1164 1371
rect 1158 1366 1164 1367
rect 1286 1371 1292 1372
rect 1286 1367 1287 1371
rect 1291 1367 1292 1371
rect 1286 1366 1292 1367
rect 1414 1371 1420 1372
rect 1414 1367 1415 1371
rect 1419 1367 1420 1371
rect 1766 1368 1767 1372
rect 1771 1368 1772 1372
rect 1766 1367 1772 1368
rect 1806 1371 1812 1372
rect 1806 1367 1807 1371
rect 1811 1367 1812 1371
rect 2166 1371 2167 1375
rect 2171 1371 2172 1375
rect 2166 1370 2172 1371
rect 2270 1375 2276 1376
rect 2270 1371 2271 1375
rect 2275 1371 2276 1375
rect 2390 1375 2391 1379
rect 2395 1375 2396 1379
rect 2390 1374 2396 1375
rect 2426 1379 2432 1380
rect 2426 1375 2427 1379
rect 2431 1378 2432 1379
rect 2534 1379 2540 1380
rect 2431 1376 2497 1378
rect 2431 1375 2432 1376
rect 2426 1374 2432 1375
rect 2534 1375 2535 1379
rect 2539 1378 2540 1379
rect 2734 1379 2740 1380
rect 2539 1376 2641 1378
rect 2539 1375 2540 1376
rect 2534 1374 2540 1375
rect 2734 1375 2735 1379
rect 2739 1378 2740 1379
rect 2838 1379 2844 1380
rect 2739 1376 2785 1378
rect 2739 1375 2740 1376
rect 2734 1374 2740 1375
rect 2838 1375 2839 1379
rect 2843 1378 2844 1379
rect 2966 1379 2972 1380
rect 2843 1376 2929 1378
rect 2843 1375 2844 1376
rect 2838 1374 2844 1375
rect 2966 1375 2967 1379
rect 2971 1378 2972 1379
rect 3111 1379 3117 1380
rect 2971 1376 3073 1378
rect 2971 1375 2972 1376
rect 2966 1374 2972 1375
rect 3111 1375 3112 1379
rect 3116 1378 3117 1379
rect 3254 1379 3260 1380
rect 3116 1376 3217 1378
rect 3116 1375 3117 1376
rect 3111 1374 3117 1375
rect 3254 1375 3255 1379
rect 3259 1378 3260 1379
rect 3259 1376 3369 1378
rect 3259 1375 3260 1376
rect 3254 1374 3260 1375
rect 2270 1370 2276 1371
rect 3462 1371 3468 1372
rect 1414 1366 1420 1367
rect 1806 1366 1812 1367
rect 2094 1368 2100 1369
rect 2094 1364 2095 1368
rect 2099 1364 2100 1368
rect 358 1363 364 1364
rect 206 1359 212 1360
rect 110 1355 116 1356
rect 110 1351 111 1355
rect 115 1351 116 1355
rect 206 1355 207 1359
rect 211 1355 212 1359
rect 206 1354 212 1355
rect 350 1359 356 1360
rect 350 1355 351 1359
rect 355 1355 356 1359
rect 358 1359 359 1363
rect 363 1362 364 1363
rect 558 1363 564 1364
rect 363 1360 489 1362
rect 363 1359 364 1360
rect 358 1358 364 1359
rect 558 1359 559 1363
rect 563 1362 564 1363
rect 738 1363 744 1364
rect 563 1360 649 1362
rect 563 1359 564 1360
rect 558 1358 564 1359
rect 738 1359 739 1363
rect 743 1362 744 1363
rect 974 1363 980 1364
rect 743 1360 801 1362
rect 743 1359 744 1360
rect 738 1358 744 1359
rect 974 1359 975 1363
rect 979 1359 980 1363
rect 974 1358 980 1359
rect 982 1363 988 1364
rect 982 1359 983 1363
rect 987 1362 988 1363
rect 1110 1363 1116 1364
rect 987 1360 1073 1362
rect 987 1359 988 1360
rect 982 1358 988 1359
rect 1110 1359 1111 1363
rect 1115 1362 1116 1363
rect 1366 1363 1372 1364
rect 2094 1363 2100 1364
rect 2198 1368 2204 1369
rect 2198 1364 2199 1368
rect 2203 1364 2204 1368
rect 2198 1363 2204 1364
rect 2318 1368 2324 1369
rect 2318 1364 2319 1368
rect 2323 1364 2324 1368
rect 2318 1363 2324 1364
rect 2454 1368 2460 1369
rect 2454 1364 2455 1368
rect 2459 1364 2460 1368
rect 2454 1363 2460 1364
rect 2598 1368 2604 1369
rect 2598 1364 2599 1368
rect 2603 1364 2604 1368
rect 2598 1363 2604 1364
rect 2742 1368 2748 1369
rect 2742 1364 2743 1368
rect 2747 1364 2748 1368
rect 2742 1363 2748 1364
rect 2886 1368 2892 1369
rect 2886 1364 2887 1368
rect 2891 1364 2892 1368
rect 2886 1363 2892 1364
rect 3030 1368 3036 1369
rect 3030 1364 3031 1368
rect 3035 1364 3036 1368
rect 3030 1363 3036 1364
rect 3174 1368 3180 1369
rect 3174 1364 3175 1368
rect 3179 1364 3180 1368
rect 3174 1363 3180 1364
rect 3326 1368 3332 1369
rect 3326 1364 3327 1368
rect 3331 1364 3332 1368
rect 3462 1367 3463 1371
rect 3467 1367 3468 1371
rect 3462 1366 3468 1367
rect 3326 1363 3332 1364
rect 1115 1360 1201 1362
rect 1115 1359 1116 1360
rect 1110 1358 1116 1359
rect 1358 1359 1364 1360
rect 350 1354 356 1355
rect 1358 1355 1359 1359
rect 1363 1355 1364 1359
rect 1366 1359 1367 1363
rect 1371 1362 1372 1363
rect 1371 1360 1457 1362
rect 1371 1359 1372 1360
rect 1366 1358 1372 1359
rect 2426 1359 2432 1360
rect 2426 1358 2427 1359
rect 2148 1356 2427 1358
rect 1358 1354 1364 1355
rect 1766 1355 1772 1356
rect 110 1350 116 1351
rect 134 1352 140 1353
rect 134 1348 135 1352
rect 139 1348 140 1352
rect 134 1347 140 1348
rect 278 1352 284 1353
rect 278 1348 279 1352
rect 283 1348 284 1352
rect 278 1347 284 1348
rect 446 1352 452 1353
rect 446 1348 447 1352
rect 451 1348 452 1352
rect 446 1347 452 1348
rect 606 1352 612 1353
rect 606 1348 607 1352
rect 611 1348 612 1352
rect 606 1347 612 1348
rect 758 1352 764 1353
rect 758 1348 759 1352
rect 763 1348 764 1352
rect 758 1347 764 1348
rect 902 1352 908 1353
rect 902 1348 903 1352
rect 907 1348 908 1352
rect 902 1347 908 1348
rect 1030 1352 1036 1353
rect 1030 1348 1031 1352
rect 1035 1348 1036 1352
rect 1030 1347 1036 1348
rect 1158 1352 1164 1353
rect 1158 1348 1159 1352
rect 1163 1348 1164 1352
rect 1158 1347 1164 1348
rect 1286 1352 1292 1353
rect 1286 1348 1287 1352
rect 1291 1348 1292 1352
rect 1286 1347 1292 1348
rect 1414 1352 1420 1353
rect 1414 1348 1415 1352
rect 1419 1348 1420 1352
rect 1766 1351 1767 1355
rect 1771 1351 1772 1355
rect 2148 1354 2150 1356
rect 2426 1355 2427 1356
rect 2431 1355 2432 1359
rect 2426 1354 2432 1355
rect 1766 1350 1772 1351
rect 2147 1353 2153 1354
rect 2147 1349 2148 1353
rect 2152 1349 2153 1353
rect 2147 1348 2153 1349
rect 2166 1351 2172 1352
rect 1414 1347 1420 1348
rect 2166 1347 2167 1351
rect 2171 1350 2172 1351
rect 2251 1351 2257 1352
rect 2251 1350 2252 1351
rect 2171 1348 2252 1350
rect 2171 1347 2172 1348
rect 2166 1346 2172 1347
rect 2251 1347 2252 1348
rect 2256 1347 2257 1351
rect 2251 1346 2257 1347
rect 2270 1351 2276 1352
rect 2270 1347 2271 1351
rect 2275 1350 2276 1351
rect 2371 1351 2377 1352
rect 2371 1350 2372 1351
rect 2275 1348 2372 1350
rect 2275 1347 2276 1348
rect 2270 1346 2276 1347
rect 2371 1347 2372 1348
rect 2376 1347 2377 1351
rect 2371 1346 2377 1347
rect 2507 1351 2513 1352
rect 2507 1347 2508 1351
rect 2512 1350 2513 1351
rect 2534 1351 2540 1352
rect 2534 1350 2535 1351
rect 2512 1348 2535 1350
rect 2512 1347 2513 1348
rect 2507 1346 2513 1347
rect 2534 1347 2535 1348
rect 2539 1347 2540 1351
rect 2534 1346 2540 1347
rect 2606 1351 2612 1352
rect 2606 1347 2607 1351
rect 2611 1350 2612 1351
rect 2651 1351 2657 1352
rect 2651 1350 2652 1351
rect 2611 1348 2652 1350
rect 2611 1347 2612 1348
rect 2606 1346 2612 1347
rect 2651 1347 2652 1348
rect 2656 1347 2657 1351
rect 2651 1346 2657 1347
rect 2702 1351 2708 1352
rect 2702 1347 2703 1351
rect 2707 1350 2708 1351
rect 2795 1351 2801 1352
rect 2795 1350 2796 1351
rect 2707 1348 2796 1350
rect 2707 1347 2708 1348
rect 2702 1346 2708 1347
rect 2795 1347 2796 1348
rect 2800 1347 2801 1351
rect 2795 1346 2801 1347
rect 2939 1351 2945 1352
rect 2939 1347 2940 1351
rect 2944 1350 2945 1351
rect 2966 1351 2972 1352
rect 2966 1350 2967 1351
rect 2944 1348 2967 1350
rect 2944 1347 2945 1348
rect 2939 1346 2945 1347
rect 2966 1347 2967 1348
rect 2971 1347 2972 1351
rect 2966 1346 2972 1347
rect 3083 1351 3089 1352
rect 3083 1347 3084 1351
rect 3088 1350 3089 1351
rect 3111 1351 3117 1352
rect 3111 1350 3112 1351
rect 3088 1348 3112 1350
rect 3088 1347 3089 1348
rect 3083 1346 3089 1347
rect 3111 1347 3112 1348
rect 3116 1347 3117 1351
rect 3111 1346 3117 1347
rect 3227 1351 3233 1352
rect 3227 1347 3228 1351
rect 3232 1350 3233 1351
rect 3254 1351 3260 1352
rect 3254 1350 3255 1351
rect 3232 1348 3255 1350
rect 3232 1347 3233 1348
rect 3227 1346 3233 1347
rect 3254 1347 3255 1348
rect 3259 1347 3260 1351
rect 3254 1346 3260 1347
rect 3374 1351 3385 1352
rect 3374 1347 3375 1351
rect 3379 1347 3380 1351
rect 3384 1347 3385 1351
rect 3374 1346 3385 1347
rect 187 1335 193 1336
rect 187 1331 188 1335
rect 192 1334 193 1335
rect 198 1335 204 1336
rect 198 1334 199 1335
rect 192 1332 199 1334
rect 192 1331 193 1332
rect 187 1330 193 1331
rect 198 1331 199 1332
rect 203 1331 204 1335
rect 198 1330 204 1331
rect 206 1335 212 1336
rect 206 1331 207 1335
rect 211 1334 212 1335
rect 331 1335 337 1336
rect 331 1334 332 1335
rect 211 1332 332 1334
rect 211 1331 212 1332
rect 206 1330 212 1331
rect 331 1331 332 1332
rect 336 1331 337 1335
rect 331 1330 337 1331
rect 350 1335 356 1336
rect 350 1331 351 1335
rect 355 1334 356 1335
rect 499 1335 505 1336
rect 499 1334 500 1335
rect 355 1332 500 1334
rect 355 1331 356 1332
rect 350 1330 356 1331
rect 499 1331 500 1332
rect 504 1331 505 1335
rect 499 1330 505 1331
rect 659 1335 665 1336
rect 659 1331 660 1335
rect 664 1334 665 1335
rect 738 1335 744 1336
rect 738 1334 739 1335
rect 664 1332 739 1334
rect 664 1331 665 1332
rect 659 1330 665 1331
rect 738 1331 739 1332
rect 743 1331 744 1335
rect 738 1330 744 1331
rect 811 1335 817 1336
rect 811 1331 812 1335
rect 816 1334 817 1335
rect 846 1335 852 1336
rect 846 1334 847 1335
rect 816 1332 847 1334
rect 816 1331 817 1332
rect 811 1330 817 1331
rect 846 1331 847 1332
rect 851 1331 852 1335
rect 846 1330 852 1331
rect 955 1335 961 1336
rect 955 1331 956 1335
rect 960 1334 961 1335
rect 982 1335 988 1336
rect 982 1334 983 1335
rect 960 1332 983 1334
rect 960 1331 961 1332
rect 955 1330 961 1331
rect 982 1331 983 1332
rect 987 1331 988 1335
rect 982 1330 988 1331
rect 1083 1335 1089 1336
rect 1083 1331 1084 1335
rect 1088 1334 1089 1335
rect 1110 1335 1116 1336
rect 1110 1334 1111 1335
rect 1088 1332 1111 1334
rect 1088 1331 1089 1332
rect 1083 1330 1089 1331
rect 1110 1331 1111 1332
rect 1115 1331 1116 1335
rect 1110 1330 1116 1331
rect 1211 1335 1217 1336
rect 1211 1331 1212 1335
rect 1216 1334 1217 1335
rect 1254 1335 1260 1336
rect 1254 1334 1255 1335
rect 1216 1332 1255 1334
rect 1216 1331 1217 1332
rect 1211 1330 1217 1331
rect 1254 1331 1255 1332
rect 1259 1331 1260 1335
rect 1254 1330 1260 1331
rect 1270 1335 1276 1336
rect 1270 1331 1271 1335
rect 1275 1334 1276 1335
rect 1339 1335 1345 1336
rect 1339 1334 1340 1335
rect 1275 1332 1340 1334
rect 1275 1331 1276 1332
rect 1270 1330 1276 1331
rect 1339 1331 1340 1332
rect 1344 1331 1345 1335
rect 1339 1330 1345 1331
rect 1358 1335 1364 1336
rect 1358 1331 1359 1335
rect 1363 1334 1364 1335
rect 1467 1335 1473 1336
rect 1467 1334 1468 1335
rect 1363 1332 1468 1334
rect 1363 1331 1364 1332
rect 1358 1330 1364 1331
rect 1467 1331 1468 1332
rect 1472 1331 1473 1335
rect 1467 1330 1473 1331
rect 2155 1335 2161 1336
rect 2155 1331 2156 1335
rect 2160 1334 2161 1335
rect 2174 1335 2180 1336
rect 2160 1332 2170 1334
rect 2160 1331 2161 1332
rect 2155 1330 2161 1331
rect 558 1327 564 1328
rect 558 1326 559 1327
rect 332 1324 559 1326
rect 332 1322 334 1324
rect 558 1323 559 1324
rect 563 1323 564 1327
rect 2168 1326 2170 1332
rect 2174 1331 2175 1335
rect 2179 1334 2180 1335
rect 2291 1335 2297 1336
rect 2291 1334 2292 1335
rect 2179 1332 2292 1334
rect 2179 1331 2180 1332
rect 2174 1330 2180 1331
rect 2291 1331 2292 1332
rect 2296 1331 2297 1335
rect 2291 1330 2297 1331
rect 2310 1335 2316 1336
rect 2310 1331 2311 1335
rect 2315 1334 2316 1335
rect 2435 1335 2441 1336
rect 2435 1334 2436 1335
rect 2315 1332 2436 1334
rect 2315 1331 2316 1332
rect 2310 1330 2316 1331
rect 2435 1331 2436 1332
rect 2440 1331 2441 1335
rect 2435 1330 2441 1331
rect 2503 1335 2509 1336
rect 2503 1331 2504 1335
rect 2508 1334 2509 1335
rect 2587 1335 2593 1336
rect 2587 1334 2588 1335
rect 2508 1332 2588 1334
rect 2508 1331 2509 1332
rect 2503 1330 2509 1331
rect 2587 1331 2588 1332
rect 2592 1331 2593 1335
rect 2587 1330 2593 1331
rect 2734 1335 2745 1336
rect 2734 1331 2735 1335
rect 2739 1331 2740 1335
rect 2744 1331 2745 1335
rect 2734 1330 2745 1331
rect 2891 1335 2897 1336
rect 2891 1331 2892 1335
rect 2896 1334 2897 1335
rect 2910 1335 2916 1336
rect 2896 1332 2906 1334
rect 2896 1331 2897 1332
rect 2891 1330 2897 1331
rect 2322 1327 2328 1328
rect 2322 1326 2323 1327
rect 2168 1324 2323 1326
rect 558 1322 564 1323
rect 2322 1323 2323 1324
rect 2327 1323 2328 1327
rect 2904 1326 2906 1332
rect 2910 1331 2911 1335
rect 2915 1334 2916 1335
rect 3043 1335 3049 1336
rect 3043 1334 3044 1335
rect 2915 1332 3044 1334
rect 2915 1331 2916 1332
rect 2910 1330 2916 1331
rect 3043 1331 3044 1332
rect 3048 1331 3049 1335
rect 3043 1330 3049 1331
rect 3062 1335 3068 1336
rect 3062 1331 3063 1335
rect 3067 1334 3068 1335
rect 3195 1335 3201 1336
rect 3195 1334 3196 1335
rect 3067 1332 3196 1334
rect 3067 1331 3068 1332
rect 3062 1330 3068 1331
rect 3195 1331 3196 1332
rect 3200 1331 3201 1335
rect 3195 1330 3201 1331
rect 3214 1335 3220 1336
rect 3214 1331 3215 1335
rect 3219 1334 3220 1335
rect 3355 1335 3361 1336
rect 3355 1334 3356 1335
rect 3219 1332 3356 1334
rect 3219 1331 3220 1332
rect 3214 1330 3220 1331
rect 3355 1331 3356 1332
rect 3360 1331 3361 1335
rect 3355 1330 3361 1331
rect 3054 1327 3060 1328
rect 3054 1326 3055 1327
rect 2904 1324 3055 1326
rect 2322 1322 2328 1323
rect 3054 1323 3055 1324
rect 3059 1323 3060 1327
rect 3054 1322 3060 1323
rect 331 1321 337 1322
rect 187 1319 193 1320
rect 187 1315 188 1319
rect 192 1318 193 1319
rect 206 1319 212 1320
rect 206 1318 207 1319
rect 192 1316 207 1318
rect 192 1315 193 1316
rect 187 1314 193 1315
rect 206 1315 207 1316
rect 211 1315 212 1319
rect 331 1317 332 1321
rect 336 1317 337 1321
rect 2102 1320 2108 1321
rect 331 1316 337 1317
rect 350 1319 356 1320
rect 206 1314 212 1315
rect 350 1315 351 1319
rect 355 1318 356 1319
rect 491 1319 497 1320
rect 491 1318 492 1319
rect 355 1316 492 1318
rect 355 1315 356 1316
rect 350 1314 356 1315
rect 491 1315 492 1316
rect 496 1315 497 1319
rect 491 1314 497 1315
rect 510 1319 516 1320
rect 510 1315 511 1319
rect 515 1318 516 1319
rect 635 1319 641 1320
rect 635 1318 636 1319
rect 515 1316 636 1318
rect 515 1315 516 1316
rect 510 1314 516 1315
rect 635 1315 636 1316
rect 640 1315 641 1319
rect 635 1314 641 1315
rect 686 1319 692 1320
rect 686 1315 687 1319
rect 691 1318 692 1319
rect 771 1319 777 1320
rect 771 1318 772 1319
rect 691 1316 772 1318
rect 691 1315 692 1316
rect 686 1314 692 1315
rect 771 1315 772 1316
rect 776 1315 777 1319
rect 771 1314 777 1315
rect 790 1319 796 1320
rect 790 1315 791 1319
rect 795 1318 796 1319
rect 899 1319 905 1320
rect 899 1318 900 1319
rect 795 1316 900 1318
rect 795 1315 796 1316
rect 790 1314 796 1315
rect 899 1315 900 1316
rect 904 1315 905 1319
rect 899 1314 905 1315
rect 918 1319 924 1320
rect 918 1315 919 1319
rect 923 1318 924 1319
rect 1019 1319 1025 1320
rect 1019 1318 1020 1319
rect 923 1316 1020 1318
rect 923 1315 924 1316
rect 918 1314 924 1315
rect 1019 1315 1020 1316
rect 1024 1315 1025 1319
rect 1019 1314 1025 1315
rect 1038 1319 1044 1320
rect 1038 1315 1039 1319
rect 1043 1318 1044 1319
rect 1131 1319 1137 1320
rect 1131 1318 1132 1319
rect 1043 1316 1132 1318
rect 1043 1315 1044 1316
rect 1038 1314 1044 1315
rect 1131 1315 1132 1316
rect 1136 1315 1137 1319
rect 1131 1314 1137 1315
rect 1243 1319 1249 1320
rect 1243 1315 1244 1319
rect 1248 1318 1249 1319
rect 1298 1319 1304 1320
rect 1298 1318 1299 1319
rect 1248 1316 1299 1318
rect 1248 1315 1249 1316
rect 1243 1314 1249 1315
rect 1298 1315 1299 1316
rect 1303 1315 1304 1319
rect 1298 1314 1304 1315
rect 1363 1319 1372 1320
rect 1363 1315 1364 1319
rect 1371 1315 1372 1319
rect 1363 1314 1372 1315
rect 1806 1317 1812 1318
rect 1806 1313 1807 1317
rect 1811 1313 1812 1317
rect 2102 1316 2103 1320
rect 2107 1316 2108 1320
rect 2102 1315 2108 1316
rect 2238 1320 2244 1321
rect 2238 1316 2239 1320
rect 2243 1316 2244 1320
rect 2238 1315 2244 1316
rect 2382 1320 2388 1321
rect 2382 1316 2383 1320
rect 2387 1316 2388 1320
rect 2382 1315 2388 1316
rect 2534 1320 2540 1321
rect 2534 1316 2535 1320
rect 2539 1316 2540 1320
rect 2534 1315 2540 1316
rect 2686 1320 2692 1321
rect 2686 1316 2687 1320
rect 2691 1316 2692 1320
rect 2686 1315 2692 1316
rect 2838 1320 2844 1321
rect 2838 1316 2839 1320
rect 2843 1316 2844 1320
rect 2838 1315 2844 1316
rect 2990 1320 2996 1321
rect 2990 1316 2991 1320
rect 2995 1316 2996 1320
rect 2990 1315 2996 1316
rect 3142 1320 3148 1321
rect 3142 1316 3143 1320
rect 3147 1316 3148 1320
rect 3142 1315 3148 1316
rect 3302 1320 3308 1321
rect 3302 1316 3303 1320
rect 3307 1316 3308 1320
rect 3302 1315 3308 1316
rect 3462 1317 3468 1318
rect 1806 1312 1812 1313
rect 3462 1313 3463 1317
rect 3467 1313 3468 1317
rect 3462 1312 3468 1313
rect 2174 1311 2180 1312
rect 2174 1307 2175 1311
rect 2179 1307 2180 1311
rect 2174 1306 2180 1307
rect 2310 1311 2316 1312
rect 2310 1307 2311 1311
rect 2315 1307 2316 1311
rect 2503 1311 2509 1312
rect 2503 1310 2504 1311
rect 2457 1308 2504 1310
rect 2310 1306 2316 1307
rect 2503 1307 2504 1308
rect 2508 1307 2509 1311
rect 2503 1306 2509 1307
rect 2606 1311 2612 1312
rect 2606 1307 2607 1311
rect 2611 1307 2612 1311
rect 2606 1306 2612 1307
rect 2750 1311 2756 1312
rect 2750 1307 2751 1311
rect 2755 1307 2756 1311
rect 2750 1306 2756 1307
rect 2910 1311 2916 1312
rect 2910 1307 2911 1311
rect 2915 1307 2916 1311
rect 2910 1306 2916 1307
rect 3062 1311 3068 1312
rect 3062 1307 3063 1311
rect 3067 1307 3068 1311
rect 3062 1306 3068 1307
rect 3214 1311 3220 1312
rect 3214 1307 3215 1311
rect 3219 1307 3220 1311
rect 3214 1306 3220 1307
rect 3374 1311 3380 1312
rect 3374 1307 3375 1311
rect 3379 1307 3380 1311
rect 3374 1306 3380 1307
rect 134 1304 140 1305
rect 110 1301 116 1302
rect 110 1297 111 1301
rect 115 1297 116 1301
rect 134 1300 135 1304
rect 139 1300 140 1304
rect 134 1299 140 1300
rect 278 1304 284 1305
rect 278 1300 279 1304
rect 283 1300 284 1304
rect 278 1299 284 1300
rect 438 1304 444 1305
rect 438 1300 439 1304
rect 443 1300 444 1304
rect 438 1299 444 1300
rect 582 1304 588 1305
rect 582 1300 583 1304
rect 587 1300 588 1304
rect 582 1299 588 1300
rect 718 1304 724 1305
rect 718 1300 719 1304
rect 723 1300 724 1304
rect 718 1299 724 1300
rect 846 1304 852 1305
rect 846 1300 847 1304
rect 851 1300 852 1304
rect 846 1299 852 1300
rect 966 1304 972 1305
rect 966 1300 967 1304
rect 971 1300 972 1304
rect 966 1299 972 1300
rect 1078 1304 1084 1305
rect 1078 1300 1079 1304
rect 1083 1300 1084 1304
rect 1078 1299 1084 1300
rect 1190 1304 1196 1305
rect 1190 1300 1191 1304
rect 1195 1300 1196 1304
rect 1190 1299 1196 1300
rect 1310 1304 1316 1305
rect 1310 1300 1311 1304
rect 1315 1300 1316 1304
rect 1310 1299 1316 1300
rect 1766 1301 1772 1302
rect 2102 1301 2108 1302
rect 110 1296 116 1297
rect 1766 1297 1767 1301
rect 1771 1297 1772 1301
rect 1766 1296 1772 1297
rect 1806 1300 1812 1301
rect 1806 1296 1807 1300
rect 1811 1296 1812 1300
rect 2102 1297 2103 1301
rect 2107 1297 2108 1301
rect 2102 1296 2108 1297
rect 2238 1301 2244 1302
rect 2238 1297 2239 1301
rect 2243 1297 2244 1301
rect 2238 1296 2244 1297
rect 2382 1301 2388 1302
rect 2382 1297 2383 1301
rect 2387 1297 2388 1301
rect 2382 1296 2388 1297
rect 2534 1301 2540 1302
rect 2534 1297 2535 1301
rect 2539 1297 2540 1301
rect 2534 1296 2540 1297
rect 2686 1301 2692 1302
rect 2686 1297 2687 1301
rect 2691 1297 2692 1301
rect 2686 1296 2692 1297
rect 2838 1301 2844 1302
rect 2838 1297 2839 1301
rect 2843 1297 2844 1301
rect 2838 1296 2844 1297
rect 2990 1301 2996 1302
rect 2990 1297 2991 1301
rect 2995 1297 2996 1301
rect 2990 1296 2996 1297
rect 3142 1301 3148 1302
rect 3142 1297 3143 1301
rect 3147 1297 3148 1301
rect 3142 1296 3148 1297
rect 3302 1301 3308 1302
rect 3302 1297 3303 1301
rect 3307 1297 3308 1301
rect 3302 1296 3308 1297
rect 3462 1300 3468 1301
rect 3462 1296 3463 1300
rect 3467 1296 3468 1300
rect 198 1295 204 1296
rect 198 1291 199 1295
rect 203 1291 204 1295
rect 198 1290 204 1291
rect 350 1295 356 1296
rect 350 1291 351 1295
rect 355 1291 356 1295
rect 350 1290 356 1291
rect 510 1295 516 1296
rect 510 1291 511 1295
rect 515 1291 516 1295
rect 510 1290 516 1291
rect 654 1295 660 1296
rect 654 1291 655 1295
rect 659 1291 660 1295
rect 654 1290 660 1291
rect 790 1295 796 1296
rect 790 1291 791 1295
rect 795 1291 796 1295
rect 790 1290 796 1291
rect 918 1295 924 1296
rect 918 1291 919 1295
rect 923 1291 924 1295
rect 918 1290 924 1291
rect 1038 1295 1044 1296
rect 1038 1291 1039 1295
rect 1043 1291 1044 1295
rect 1038 1290 1044 1291
rect 1046 1295 1052 1296
rect 1046 1291 1047 1295
rect 1051 1294 1052 1295
rect 1254 1295 1260 1296
rect 1051 1292 1121 1294
rect 1051 1291 1052 1292
rect 1046 1290 1052 1291
rect 1254 1291 1255 1295
rect 1259 1291 1260 1295
rect 1254 1290 1260 1291
rect 1298 1295 1304 1296
rect 1806 1295 1812 1296
rect 3462 1295 3468 1296
rect 1298 1291 1299 1295
rect 1303 1294 1304 1295
rect 1303 1292 1353 1294
rect 1303 1291 1304 1292
rect 1298 1290 1304 1291
rect 134 1285 140 1286
rect 110 1284 116 1285
rect 110 1280 111 1284
rect 115 1280 116 1284
rect 134 1281 135 1285
rect 139 1281 140 1285
rect 134 1280 140 1281
rect 278 1285 284 1286
rect 278 1281 279 1285
rect 283 1281 284 1285
rect 278 1280 284 1281
rect 438 1285 444 1286
rect 438 1281 439 1285
rect 443 1281 444 1285
rect 438 1280 444 1281
rect 582 1285 588 1286
rect 582 1281 583 1285
rect 587 1281 588 1285
rect 582 1280 588 1281
rect 718 1285 724 1286
rect 718 1281 719 1285
rect 723 1281 724 1285
rect 718 1280 724 1281
rect 846 1285 852 1286
rect 846 1281 847 1285
rect 851 1281 852 1285
rect 846 1280 852 1281
rect 966 1285 972 1286
rect 966 1281 967 1285
rect 971 1281 972 1285
rect 966 1280 972 1281
rect 1078 1285 1084 1286
rect 1078 1281 1079 1285
rect 1083 1281 1084 1285
rect 1078 1280 1084 1281
rect 1190 1285 1196 1286
rect 1190 1281 1191 1285
rect 1195 1281 1196 1285
rect 1190 1280 1196 1281
rect 1310 1285 1316 1286
rect 1310 1281 1311 1285
rect 1315 1281 1316 1285
rect 1310 1280 1316 1281
rect 1766 1284 1772 1285
rect 1766 1280 1767 1284
rect 1771 1280 1772 1284
rect 110 1279 116 1280
rect 1766 1279 1772 1280
rect 1806 1256 1812 1257
rect 3462 1256 3468 1257
rect 1806 1252 1807 1256
rect 1811 1252 1812 1256
rect 1806 1251 1812 1252
rect 1934 1255 1940 1256
rect 1934 1251 1935 1255
rect 1939 1251 1940 1255
rect 1934 1250 1940 1251
rect 2062 1255 2068 1256
rect 2062 1251 2063 1255
rect 2067 1251 2068 1255
rect 2062 1250 2068 1251
rect 2198 1255 2204 1256
rect 2198 1251 2199 1255
rect 2203 1251 2204 1255
rect 2198 1250 2204 1251
rect 2342 1255 2348 1256
rect 2342 1251 2343 1255
rect 2347 1251 2348 1255
rect 2342 1250 2348 1251
rect 2494 1255 2500 1256
rect 2494 1251 2495 1255
rect 2499 1251 2500 1255
rect 2494 1250 2500 1251
rect 2654 1255 2660 1256
rect 2654 1251 2655 1255
rect 2659 1251 2660 1255
rect 2654 1250 2660 1251
rect 2814 1255 2820 1256
rect 2814 1251 2815 1255
rect 2819 1251 2820 1255
rect 2814 1250 2820 1251
rect 2974 1255 2980 1256
rect 2974 1251 2975 1255
rect 2979 1251 2980 1255
rect 2974 1250 2980 1251
rect 3142 1255 3148 1256
rect 3142 1251 3143 1255
rect 3147 1251 3148 1255
rect 3462 1252 3463 1256
rect 3467 1252 3468 1256
rect 3462 1251 3468 1252
rect 3142 1250 3148 1251
rect 2322 1247 2328 1248
rect 2006 1243 2012 1244
rect 1806 1239 1812 1240
rect 110 1236 116 1237
rect 1766 1236 1772 1237
rect 110 1232 111 1236
rect 115 1232 116 1236
rect 110 1231 116 1232
rect 134 1235 140 1236
rect 134 1231 135 1235
rect 139 1231 140 1235
rect 134 1230 140 1231
rect 238 1235 244 1236
rect 238 1231 239 1235
rect 243 1231 244 1235
rect 238 1230 244 1231
rect 366 1235 372 1236
rect 366 1231 367 1235
rect 371 1231 372 1235
rect 366 1230 372 1231
rect 494 1235 500 1236
rect 494 1231 495 1235
rect 499 1231 500 1235
rect 494 1230 500 1231
rect 614 1235 620 1236
rect 614 1231 615 1235
rect 619 1231 620 1235
rect 614 1230 620 1231
rect 734 1235 740 1236
rect 734 1231 735 1235
rect 739 1231 740 1235
rect 734 1230 740 1231
rect 846 1235 852 1236
rect 846 1231 847 1235
rect 851 1231 852 1235
rect 846 1230 852 1231
rect 958 1235 964 1236
rect 958 1231 959 1235
rect 963 1231 964 1235
rect 958 1230 964 1231
rect 1070 1235 1076 1236
rect 1070 1231 1071 1235
rect 1075 1231 1076 1235
rect 1070 1230 1076 1231
rect 1190 1235 1196 1236
rect 1190 1231 1191 1235
rect 1195 1231 1196 1235
rect 1766 1232 1767 1236
rect 1771 1232 1772 1236
rect 1806 1235 1807 1239
rect 1811 1235 1812 1239
rect 2006 1239 2007 1243
rect 2011 1239 2012 1243
rect 2006 1238 2012 1239
rect 2134 1243 2140 1244
rect 2134 1239 2135 1243
rect 2139 1239 2140 1243
rect 2134 1238 2140 1239
rect 2270 1243 2276 1244
rect 2270 1239 2271 1243
rect 2275 1239 2276 1243
rect 2322 1243 2323 1247
rect 2327 1246 2328 1247
rect 2574 1247 2580 1248
rect 2327 1244 2385 1246
rect 2327 1243 2328 1244
rect 2322 1242 2328 1243
rect 2566 1243 2572 1244
rect 2270 1238 2276 1239
rect 2566 1239 2567 1243
rect 2571 1239 2572 1243
rect 2574 1243 2575 1247
rect 2579 1246 2580 1247
rect 3054 1247 3060 1248
rect 2579 1244 2697 1246
rect 2579 1243 2580 1244
rect 2574 1242 2580 1243
rect 2886 1243 2892 1244
rect 2566 1238 2572 1239
rect 2886 1239 2887 1243
rect 2891 1239 2892 1243
rect 2886 1238 2892 1239
rect 3046 1243 3052 1244
rect 3046 1239 3047 1243
rect 3051 1239 3052 1243
rect 3054 1243 3055 1247
rect 3059 1246 3060 1247
rect 3059 1244 3185 1246
rect 3059 1243 3060 1244
rect 3054 1242 3060 1243
rect 3046 1238 3052 1239
rect 3462 1239 3468 1240
rect 1806 1234 1812 1235
rect 1934 1236 1940 1237
rect 1766 1231 1772 1232
rect 1934 1232 1935 1236
rect 1939 1232 1940 1236
rect 1934 1231 1940 1232
rect 2062 1236 2068 1237
rect 2062 1232 2063 1236
rect 2067 1232 2068 1236
rect 2062 1231 2068 1232
rect 2198 1236 2204 1237
rect 2198 1232 2199 1236
rect 2203 1232 2204 1236
rect 2198 1231 2204 1232
rect 2342 1236 2348 1237
rect 2342 1232 2343 1236
rect 2347 1232 2348 1236
rect 2342 1231 2348 1232
rect 2494 1236 2500 1237
rect 2494 1232 2495 1236
rect 2499 1232 2500 1236
rect 2494 1231 2500 1232
rect 2654 1236 2660 1237
rect 2654 1232 2655 1236
rect 2659 1232 2660 1236
rect 2654 1231 2660 1232
rect 2814 1236 2820 1237
rect 2814 1232 2815 1236
rect 2819 1232 2820 1236
rect 2814 1231 2820 1232
rect 2974 1236 2980 1237
rect 2974 1232 2975 1236
rect 2979 1232 2980 1236
rect 2974 1231 2980 1232
rect 3142 1236 3148 1237
rect 3142 1232 3143 1236
rect 3147 1232 3148 1236
rect 3462 1235 3463 1239
rect 3467 1235 3468 1239
rect 3462 1234 3468 1235
rect 3142 1231 3148 1232
rect 1190 1230 1196 1231
rect 206 1227 212 1228
rect 206 1223 207 1227
rect 211 1223 212 1227
rect 206 1222 212 1223
rect 214 1227 220 1228
rect 214 1223 215 1227
rect 219 1226 220 1227
rect 318 1227 324 1228
rect 219 1224 281 1226
rect 219 1223 220 1224
rect 214 1222 220 1223
rect 318 1223 319 1227
rect 323 1226 324 1227
rect 446 1227 452 1228
rect 323 1224 409 1226
rect 323 1223 324 1224
rect 318 1222 324 1223
rect 446 1223 447 1227
rect 451 1226 452 1227
rect 686 1227 692 1228
rect 451 1224 537 1226
rect 451 1223 452 1224
rect 446 1222 452 1223
rect 686 1223 687 1227
rect 691 1223 692 1227
rect 1150 1227 1156 1228
rect 686 1222 692 1223
rect 806 1223 812 1224
rect 110 1219 116 1220
rect 110 1215 111 1219
rect 115 1215 116 1219
rect 806 1219 807 1223
rect 811 1219 812 1223
rect 806 1218 812 1219
rect 918 1223 924 1224
rect 918 1219 919 1223
rect 923 1219 924 1223
rect 918 1218 924 1219
rect 1030 1223 1036 1224
rect 1030 1219 1031 1223
rect 1035 1219 1036 1223
rect 1030 1218 1036 1219
rect 1142 1223 1148 1224
rect 1142 1219 1143 1223
rect 1147 1219 1148 1223
rect 1150 1223 1151 1227
rect 1155 1226 1156 1227
rect 2310 1227 2316 1228
rect 2310 1226 2311 1227
rect 1155 1224 1233 1226
rect 1988 1224 2311 1226
rect 1155 1223 1156 1224
rect 1150 1222 1156 1223
rect 1988 1222 1990 1224
rect 2310 1223 2311 1224
rect 2315 1223 2316 1227
rect 2310 1222 2316 1223
rect 1987 1221 1993 1222
rect 1142 1218 1148 1219
rect 1766 1219 1772 1220
rect 110 1214 116 1215
rect 134 1216 140 1217
rect 134 1212 135 1216
rect 139 1212 140 1216
rect 134 1211 140 1212
rect 238 1216 244 1217
rect 238 1212 239 1216
rect 243 1212 244 1216
rect 238 1211 244 1212
rect 366 1216 372 1217
rect 366 1212 367 1216
rect 371 1212 372 1216
rect 366 1211 372 1212
rect 494 1216 500 1217
rect 494 1212 495 1216
rect 499 1212 500 1216
rect 494 1211 500 1212
rect 614 1216 620 1217
rect 614 1212 615 1216
rect 619 1212 620 1216
rect 614 1211 620 1212
rect 734 1216 740 1217
rect 734 1212 735 1216
rect 739 1212 740 1216
rect 734 1211 740 1212
rect 846 1216 852 1217
rect 846 1212 847 1216
rect 851 1212 852 1216
rect 846 1211 852 1212
rect 958 1216 964 1217
rect 958 1212 959 1216
rect 963 1212 964 1216
rect 958 1211 964 1212
rect 1070 1216 1076 1217
rect 1070 1212 1071 1216
rect 1075 1212 1076 1216
rect 1070 1211 1076 1212
rect 1190 1216 1196 1217
rect 1190 1212 1191 1216
rect 1195 1212 1196 1216
rect 1766 1215 1767 1219
rect 1771 1215 1772 1219
rect 1987 1217 1988 1221
rect 1992 1217 1993 1221
rect 1987 1216 1993 1217
rect 2006 1219 2012 1220
rect 1766 1214 1772 1215
rect 2006 1215 2007 1219
rect 2011 1218 2012 1219
rect 2115 1219 2121 1220
rect 2115 1218 2116 1219
rect 2011 1216 2116 1218
rect 2011 1215 2012 1216
rect 2006 1214 2012 1215
rect 2115 1215 2116 1216
rect 2120 1215 2121 1219
rect 2115 1214 2121 1215
rect 2134 1219 2140 1220
rect 2134 1215 2135 1219
rect 2139 1218 2140 1219
rect 2251 1219 2257 1220
rect 2251 1218 2252 1219
rect 2139 1216 2252 1218
rect 2139 1215 2140 1216
rect 2134 1214 2140 1215
rect 2251 1215 2252 1216
rect 2256 1215 2257 1219
rect 2251 1214 2257 1215
rect 2270 1219 2276 1220
rect 2270 1215 2271 1219
rect 2275 1218 2276 1219
rect 2395 1219 2401 1220
rect 2395 1218 2396 1219
rect 2275 1216 2396 1218
rect 2275 1215 2276 1216
rect 2270 1214 2276 1215
rect 2395 1215 2396 1216
rect 2400 1215 2401 1219
rect 2395 1214 2401 1215
rect 2547 1219 2553 1220
rect 2547 1215 2548 1219
rect 2552 1218 2553 1219
rect 2574 1219 2580 1220
rect 2574 1218 2575 1219
rect 2552 1216 2575 1218
rect 2552 1215 2553 1216
rect 2547 1214 2553 1215
rect 2574 1215 2575 1216
rect 2579 1215 2580 1219
rect 2574 1214 2580 1215
rect 2707 1219 2713 1220
rect 2707 1215 2708 1219
rect 2712 1218 2713 1219
rect 2750 1219 2756 1220
rect 2750 1218 2751 1219
rect 2712 1216 2751 1218
rect 2712 1215 2713 1216
rect 2707 1214 2713 1215
rect 2750 1215 2751 1216
rect 2755 1215 2756 1219
rect 2750 1214 2756 1215
rect 2766 1219 2772 1220
rect 2766 1215 2767 1219
rect 2771 1218 2772 1219
rect 2867 1219 2873 1220
rect 2867 1218 2868 1219
rect 2771 1216 2868 1218
rect 2771 1215 2772 1216
rect 2766 1214 2772 1215
rect 2867 1215 2868 1216
rect 2872 1215 2873 1219
rect 2867 1214 2873 1215
rect 2886 1219 2892 1220
rect 2886 1215 2887 1219
rect 2891 1218 2892 1219
rect 3027 1219 3033 1220
rect 3027 1218 3028 1219
rect 2891 1216 3028 1218
rect 2891 1215 2892 1216
rect 2886 1214 2892 1215
rect 3027 1215 3028 1216
rect 3032 1215 3033 1219
rect 3027 1214 3033 1215
rect 3046 1219 3052 1220
rect 3046 1215 3047 1219
rect 3051 1218 3052 1219
rect 3195 1219 3201 1220
rect 3195 1218 3196 1219
rect 3051 1216 3196 1218
rect 3051 1215 3052 1216
rect 3046 1214 3052 1215
rect 3195 1215 3196 1216
rect 3200 1215 3201 1219
rect 3195 1214 3201 1215
rect 1190 1211 1196 1212
rect 1046 1207 1052 1208
rect 1046 1206 1047 1207
rect 788 1204 1047 1206
rect 788 1202 790 1204
rect 1046 1203 1047 1204
rect 1051 1203 1052 1207
rect 1046 1202 1052 1203
rect 1883 1207 1889 1208
rect 1883 1203 1884 1207
rect 1888 1206 1889 1207
rect 1926 1207 1932 1208
rect 1926 1206 1927 1207
rect 1888 1204 1927 1206
rect 1888 1203 1889 1204
rect 1883 1202 1889 1203
rect 1926 1203 1927 1204
rect 1931 1203 1932 1207
rect 1987 1207 1993 1208
rect 1987 1206 1988 1207
rect 1926 1202 1932 1203
rect 1936 1204 1988 1206
rect 787 1201 793 1202
rect 187 1199 193 1200
rect 187 1195 188 1199
rect 192 1198 193 1199
rect 214 1199 220 1200
rect 214 1198 215 1199
rect 192 1196 215 1198
rect 192 1195 193 1196
rect 187 1194 193 1195
rect 214 1195 215 1196
rect 219 1195 220 1199
rect 214 1194 220 1195
rect 291 1199 297 1200
rect 291 1195 292 1199
rect 296 1198 297 1199
rect 318 1199 324 1200
rect 318 1198 319 1199
rect 296 1196 319 1198
rect 296 1195 297 1196
rect 291 1194 297 1195
rect 318 1195 319 1196
rect 323 1195 324 1199
rect 318 1194 324 1195
rect 419 1199 425 1200
rect 419 1195 420 1199
rect 424 1198 425 1199
rect 446 1199 452 1200
rect 446 1198 447 1199
rect 424 1196 447 1198
rect 424 1195 425 1196
rect 419 1194 425 1195
rect 446 1195 447 1196
rect 451 1195 452 1199
rect 446 1194 452 1195
rect 547 1199 553 1200
rect 547 1195 548 1199
rect 552 1198 553 1199
rect 622 1199 628 1200
rect 622 1198 623 1199
rect 552 1196 623 1198
rect 552 1195 553 1196
rect 547 1194 553 1195
rect 622 1195 623 1196
rect 627 1195 628 1199
rect 622 1194 628 1195
rect 654 1199 660 1200
rect 654 1195 655 1199
rect 659 1198 660 1199
rect 667 1199 673 1200
rect 667 1198 668 1199
rect 659 1196 668 1198
rect 659 1195 660 1196
rect 654 1194 660 1195
rect 667 1195 668 1196
rect 672 1195 673 1199
rect 787 1197 788 1201
rect 792 1197 793 1201
rect 787 1196 793 1197
rect 806 1199 812 1200
rect 667 1194 673 1195
rect 806 1195 807 1199
rect 811 1198 812 1199
rect 899 1199 905 1200
rect 899 1198 900 1199
rect 811 1196 900 1198
rect 811 1195 812 1196
rect 806 1194 812 1195
rect 899 1195 900 1196
rect 904 1195 905 1199
rect 899 1194 905 1195
rect 918 1199 924 1200
rect 918 1195 919 1199
rect 923 1198 924 1199
rect 1011 1199 1017 1200
rect 1011 1198 1012 1199
rect 923 1196 1012 1198
rect 923 1195 924 1196
rect 918 1194 924 1195
rect 1011 1195 1012 1196
rect 1016 1195 1017 1199
rect 1011 1194 1017 1195
rect 1030 1199 1036 1200
rect 1030 1195 1031 1199
rect 1035 1198 1036 1199
rect 1123 1199 1129 1200
rect 1123 1198 1124 1199
rect 1035 1196 1124 1198
rect 1035 1195 1036 1196
rect 1030 1194 1036 1195
rect 1123 1195 1124 1196
rect 1128 1195 1129 1199
rect 1123 1194 1129 1195
rect 1142 1199 1148 1200
rect 1142 1195 1143 1199
rect 1147 1198 1148 1199
rect 1243 1199 1249 1200
rect 1243 1198 1244 1199
rect 1147 1196 1244 1198
rect 1147 1195 1148 1196
rect 1142 1194 1148 1195
rect 1243 1195 1244 1196
rect 1248 1195 1249 1199
rect 1936 1198 1938 1204
rect 1987 1203 1988 1204
rect 1992 1203 1993 1207
rect 1987 1202 1993 1203
rect 2006 1207 2012 1208
rect 2006 1203 2007 1207
rect 2011 1206 2012 1207
rect 2131 1207 2137 1208
rect 2131 1206 2132 1207
rect 2011 1204 2132 1206
rect 2011 1203 2012 1204
rect 2006 1202 2012 1203
rect 2131 1203 2132 1204
rect 2136 1203 2137 1207
rect 2131 1202 2137 1203
rect 2150 1207 2156 1208
rect 2150 1203 2151 1207
rect 2155 1206 2156 1207
rect 2283 1207 2289 1208
rect 2283 1206 2284 1207
rect 2155 1204 2284 1206
rect 2155 1203 2156 1204
rect 2150 1202 2156 1203
rect 2283 1203 2284 1204
rect 2288 1203 2289 1207
rect 2283 1202 2289 1203
rect 2302 1207 2308 1208
rect 2302 1203 2303 1207
rect 2307 1206 2308 1207
rect 2443 1207 2449 1208
rect 2443 1206 2444 1207
rect 2307 1204 2444 1206
rect 2307 1203 2308 1204
rect 2302 1202 2308 1203
rect 2443 1203 2444 1204
rect 2448 1203 2449 1207
rect 2443 1202 2449 1203
rect 2566 1207 2572 1208
rect 2566 1203 2567 1207
rect 2571 1206 2572 1207
rect 2595 1207 2601 1208
rect 2595 1206 2596 1207
rect 2571 1204 2596 1206
rect 2571 1203 2572 1204
rect 2566 1202 2572 1203
rect 2595 1203 2596 1204
rect 2600 1203 2601 1207
rect 2595 1202 2601 1203
rect 2747 1207 2753 1208
rect 2747 1203 2748 1207
rect 2752 1206 2753 1207
rect 2774 1207 2780 1208
rect 2774 1206 2775 1207
rect 2752 1204 2775 1206
rect 2752 1203 2753 1204
rect 2747 1202 2753 1203
rect 2774 1203 2775 1204
rect 2779 1203 2780 1207
rect 2774 1202 2780 1203
rect 2899 1207 2905 1208
rect 2899 1203 2900 1207
rect 2904 1206 2905 1207
rect 2942 1207 2948 1208
rect 2904 1204 2938 1206
rect 2904 1203 2905 1204
rect 2899 1202 2905 1203
rect 1243 1194 1249 1195
rect 1904 1196 1938 1198
rect 2936 1198 2938 1204
rect 2942 1203 2943 1207
rect 2947 1206 2948 1207
rect 3051 1207 3057 1208
rect 3051 1206 3052 1207
rect 2947 1204 3052 1206
rect 2947 1203 2948 1204
rect 2942 1202 2948 1203
rect 3051 1203 3052 1204
rect 3056 1203 3057 1207
rect 3051 1202 3057 1203
rect 3070 1207 3076 1208
rect 3070 1203 3071 1207
rect 3075 1206 3076 1207
rect 3211 1207 3217 1208
rect 3211 1206 3212 1207
rect 3075 1204 3212 1206
rect 3075 1203 3076 1204
rect 3070 1202 3076 1203
rect 3211 1203 3212 1204
rect 3216 1203 3217 1207
rect 3211 1202 3217 1203
rect 2936 1196 3082 1198
rect 1830 1192 1836 1193
rect 1150 1191 1156 1192
rect 1150 1190 1151 1191
rect 844 1188 1151 1190
rect 844 1186 846 1188
rect 1150 1187 1151 1188
rect 1155 1187 1156 1191
rect 1150 1186 1156 1187
rect 1806 1189 1812 1190
rect 843 1185 849 1186
rect 182 1183 193 1184
rect 182 1179 183 1183
rect 187 1179 188 1183
rect 192 1179 193 1183
rect 182 1178 193 1179
rect 206 1183 212 1184
rect 206 1179 207 1183
rect 211 1182 212 1183
rect 291 1183 297 1184
rect 291 1182 292 1183
rect 211 1180 292 1182
rect 211 1179 212 1180
rect 206 1178 212 1179
rect 291 1179 292 1180
rect 296 1179 297 1183
rect 291 1178 297 1179
rect 310 1183 316 1184
rect 310 1179 311 1183
rect 315 1182 316 1183
rect 427 1183 433 1184
rect 427 1182 428 1183
rect 315 1180 428 1182
rect 315 1179 316 1180
rect 310 1178 316 1179
rect 427 1179 428 1180
rect 432 1179 433 1183
rect 427 1178 433 1179
rect 446 1183 452 1184
rect 446 1179 447 1183
rect 451 1182 452 1183
rect 563 1183 569 1184
rect 563 1182 564 1183
rect 451 1180 564 1182
rect 451 1179 452 1180
rect 446 1178 452 1179
rect 563 1179 564 1180
rect 568 1179 569 1183
rect 563 1178 569 1179
rect 582 1183 588 1184
rect 582 1179 583 1183
rect 587 1182 588 1183
rect 707 1183 713 1184
rect 707 1182 708 1183
rect 587 1180 708 1182
rect 587 1179 588 1180
rect 582 1178 588 1179
rect 707 1179 708 1180
rect 712 1179 713 1183
rect 843 1181 844 1185
rect 848 1181 849 1185
rect 1806 1185 1807 1189
rect 1811 1185 1812 1189
rect 1830 1188 1831 1192
rect 1835 1188 1836 1192
rect 1830 1187 1836 1188
rect 1806 1184 1812 1185
rect 843 1180 849 1181
rect 862 1183 868 1184
rect 707 1178 713 1179
rect 862 1179 863 1183
rect 867 1182 868 1183
rect 979 1183 985 1184
rect 979 1182 980 1183
rect 867 1180 980 1182
rect 867 1179 868 1180
rect 862 1178 868 1179
rect 979 1179 980 1180
rect 984 1179 985 1183
rect 979 1178 985 1179
rect 998 1183 1004 1184
rect 998 1179 999 1183
rect 1003 1182 1004 1183
rect 1115 1183 1121 1184
rect 1115 1182 1116 1183
rect 1003 1180 1116 1182
rect 1003 1179 1004 1180
rect 998 1178 1004 1179
rect 1115 1179 1116 1180
rect 1120 1179 1121 1183
rect 1115 1178 1121 1179
rect 1134 1183 1140 1184
rect 1134 1179 1135 1183
rect 1139 1182 1140 1183
rect 1251 1183 1257 1184
rect 1251 1182 1252 1183
rect 1139 1180 1252 1182
rect 1139 1179 1140 1180
rect 1134 1178 1140 1179
rect 1251 1179 1252 1180
rect 1256 1179 1257 1183
rect 1251 1178 1257 1179
rect 1270 1183 1276 1184
rect 1270 1179 1271 1183
rect 1275 1182 1276 1183
rect 1387 1183 1393 1184
rect 1387 1182 1388 1183
rect 1275 1180 1388 1182
rect 1275 1179 1276 1180
rect 1270 1178 1276 1179
rect 1387 1179 1388 1180
rect 1392 1179 1393 1183
rect 1904 1181 1906 1196
rect 1934 1192 1940 1193
rect 1934 1188 1935 1192
rect 1939 1188 1940 1192
rect 1934 1187 1940 1188
rect 2078 1192 2084 1193
rect 2078 1188 2079 1192
rect 2083 1188 2084 1192
rect 2078 1187 2084 1188
rect 2230 1192 2236 1193
rect 2230 1188 2231 1192
rect 2235 1188 2236 1192
rect 2230 1187 2236 1188
rect 2390 1192 2396 1193
rect 2390 1188 2391 1192
rect 2395 1188 2396 1192
rect 2390 1187 2396 1188
rect 2542 1192 2548 1193
rect 2542 1188 2543 1192
rect 2547 1188 2548 1192
rect 2542 1187 2548 1188
rect 2694 1192 2700 1193
rect 2694 1188 2695 1192
rect 2699 1188 2700 1192
rect 2694 1187 2700 1188
rect 2846 1192 2852 1193
rect 2846 1188 2847 1192
rect 2851 1188 2852 1192
rect 2846 1187 2852 1188
rect 2998 1192 3004 1193
rect 2998 1188 2999 1192
rect 3003 1188 3004 1192
rect 2998 1187 3004 1188
rect 2006 1183 2012 1184
rect 1387 1178 1393 1179
rect 2006 1179 2007 1183
rect 2011 1179 2012 1183
rect 2006 1178 2012 1179
rect 2150 1183 2156 1184
rect 2150 1179 2151 1183
rect 2155 1179 2156 1183
rect 2150 1178 2156 1179
rect 2302 1183 2308 1184
rect 2302 1179 2303 1183
rect 2307 1179 2308 1183
rect 2302 1178 2308 1179
rect 2310 1183 2316 1184
rect 2310 1179 2311 1183
rect 2315 1182 2316 1183
rect 2606 1183 2612 1184
rect 2315 1180 2433 1182
rect 2315 1179 2316 1180
rect 2310 1178 2316 1179
rect 2606 1179 2607 1183
rect 2611 1179 2612 1183
rect 2606 1178 2612 1179
rect 2766 1183 2772 1184
rect 2766 1179 2767 1183
rect 2771 1179 2772 1183
rect 2766 1178 2772 1179
rect 2774 1183 2780 1184
rect 2774 1179 2775 1183
rect 2779 1182 2780 1183
rect 3070 1183 3076 1184
rect 2779 1180 2889 1182
rect 2779 1179 2780 1180
rect 2774 1178 2780 1179
rect 3070 1179 3071 1183
rect 3075 1179 3076 1183
rect 3080 1182 3082 1196
rect 3158 1192 3164 1193
rect 3158 1188 3159 1192
rect 3163 1188 3164 1192
rect 3158 1187 3164 1188
rect 3462 1189 3468 1190
rect 3462 1185 3463 1189
rect 3467 1185 3468 1189
rect 3462 1184 3468 1185
rect 3080 1180 3201 1182
rect 3070 1178 3076 1179
rect 1830 1173 1836 1174
rect 1806 1172 1812 1173
rect 134 1168 140 1169
rect 110 1165 116 1166
rect 110 1161 111 1165
rect 115 1161 116 1165
rect 134 1164 135 1168
rect 139 1164 140 1168
rect 134 1163 140 1164
rect 238 1168 244 1169
rect 238 1164 239 1168
rect 243 1164 244 1168
rect 238 1163 244 1164
rect 374 1168 380 1169
rect 374 1164 375 1168
rect 379 1164 380 1168
rect 374 1163 380 1164
rect 510 1168 516 1169
rect 510 1164 511 1168
rect 515 1164 516 1168
rect 510 1163 516 1164
rect 654 1168 660 1169
rect 654 1164 655 1168
rect 659 1164 660 1168
rect 654 1163 660 1164
rect 790 1168 796 1169
rect 790 1164 791 1168
rect 795 1164 796 1168
rect 790 1163 796 1164
rect 926 1168 932 1169
rect 926 1164 927 1168
rect 931 1164 932 1168
rect 926 1163 932 1164
rect 1062 1168 1068 1169
rect 1062 1164 1063 1168
rect 1067 1164 1068 1168
rect 1062 1163 1068 1164
rect 1198 1168 1204 1169
rect 1198 1164 1199 1168
rect 1203 1164 1204 1168
rect 1198 1163 1204 1164
rect 1334 1168 1340 1169
rect 1334 1164 1335 1168
rect 1339 1164 1340 1168
rect 1806 1168 1807 1172
rect 1811 1168 1812 1172
rect 1830 1169 1831 1173
rect 1835 1169 1836 1173
rect 1830 1168 1836 1169
rect 1934 1173 1940 1174
rect 1934 1169 1935 1173
rect 1939 1169 1940 1173
rect 1934 1168 1940 1169
rect 2078 1173 2084 1174
rect 2078 1169 2079 1173
rect 2083 1169 2084 1173
rect 2078 1168 2084 1169
rect 2230 1173 2236 1174
rect 2230 1169 2231 1173
rect 2235 1169 2236 1173
rect 2230 1168 2236 1169
rect 2390 1173 2396 1174
rect 2390 1169 2391 1173
rect 2395 1169 2396 1173
rect 2390 1168 2396 1169
rect 2542 1173 2548 1174
rect 2542 1169 2543 1173
rect 2547 1169 2548 1173
rect 2542 1168 2548 1169
rect 2694 1173 2700 1174
rect 2694 1169 2695 1173
rect 2699 1169 2700 1173
rect 2694 1168 2700 1169
rect 2846 1173 2852 1174
rect 2846 1169 2847 1173
rect 2851 1169 2852 1173
rect 2846 1168 2852 1169
rect 2998 1173 3004 1174
rect 2998 1169 2999 1173
rect 3003 1169 3004 1173
rect 2998 1168 3004 1169
rect 3158 1173 3164 1174
rect 3158 1169 3159 1173
rect 3163 1169 3164 1173
rect 3158 1168 3164 1169
rect 3462 1172 3468 1173
rect 3462 1168 3463 1172
rect 3467 1168 3468 1172
rect 1806 1167 1812 1168
rect 3462 1167 3468 1168
rect 1334 1163 1340 1164
rect 1766 1165 1772 1166
rect 110 1160 116 1161
rect 1766 1161 1767 1165
rect 1771 1161 1772 1165
rect 1766 1160 1772 1161
rect 206 1159 212 1160
rect 206 1155 207 1159
rect 211 1155 212 1159
rect 206 1154 212 1155
rect 310 1159 316 1160
rect 310 1155 311 1159
rect 315 1155 316 1159
rect 310 1154 316 1155
rect 446 1159 452 1160
rect 446 1155 447 1159
rect 451 1155 452 1159
rect 446 1154 452 1155
rect 582 1159 588 1160
rect 582 1155 583 1159
rect 587 1155 588 1159
rect 582 1154 588 1155
rect 622 1159 628 1160
rect 622 1155 623 1159
rect 627 1158 628 1159
rect 862 1159 868 1160
rect 627 1156 697 1158
rect 627 1155 628 1156
rect 622 1154 628 1155
rect 862 1155 863 1159
rect 867 1155 868 1159
rect 862 1154 868 1155
rect 998 1159 1004 1160
rect 998 1155 999 1159
rect 1003 1155 1004 1159
rect 998 1154 1004 1155
rect 1134 1159 1140 1160
rect 1134 1155 1135 1159
rect 1139 1155 1140 1159
rect 1134 1154 1140 1155
rect 1270 1159 1276 1160
rect 1270 1155 1271 1159
rect 1275 1155 1276 1159
rect 1270 1154 1276 1155
rect 1278 1159 1284 1160
rect 1278 1155 1279 1159
rect 1283 1158 1284 1159
rect 1283 1156 1377 1158
rect 1283 1155 1284 1156
rect 1278 1154 1284 1155
rect 134 1149 140 1150
rect 110 1148 116 1149
rect 110 1144 111 1148
rect 115 1144 116 1148
rect 134 1145 135 1149
rect 139 1145 140 1149
rect 134 1144 140 1145
rect 238 1149 244 1150
rect 238 1145 239 1149
rect 243 1145 244 1149
rect 238 1144 244 1145
rect 374 1149 380 1150
rect 374 1145 375 1149
rect 379 1145 380 1149
rect 374 1144 380 1145
rect 510 1149 516 1150
rect 510 1145 511 1149
rect 515 1145 516 1149
rect 510 1144 516 1145
rect 654 1149 660 1150
rect 654 1145 655 1149
rect 659 1145 660 1149
rect 654 1144 660 1145
rect 790 1149 796 1150
rect 790 1145 791 1149
rect 795 1145 796 1149
rect 790 1144 796 1145
rect 926 1149 932 1150
rect 926 1145 927 1149
rect 931 1145 932 1149
rect 926 1144 932 1145
rect 1062 1149 1068 1150
rect 1062 1145 1063 1149
rect 1067 1145 1068 1149
rect 1062 1144 1068 1145
rect 1198 1149 1204 1150
rect 1198 1145 1199 1149
rect 1203 1145 1204 1149
rect 1198 1144 1204 1145
rect 1334 1149 1340 1150
rect 1334 1145 1335 1149
rect 1339 1145 1340 1149
rect 1334 1144 1340 1145
rect 1766 1148 1772 1149
rect 1766 1144 1767 1148
rect 1771 1144 1772 1148
rect 110 1143 116 1144
rect 1766 1143 1772 1144
rect 1806 1116 1812 1117
rect 3462 1116 3468 1117
rect 1806 1112 1807 1116
rect 1811 1112 1812 1116
rect 1806 1111 1812 1112
rect 1862 1115 1868 1116
rect 1862 1111 1863 1115
rect 1867 1111 1868 1115
rect 1982 1115 1988 1116
rect 1862 1110 1868 1111
rect 1926 1111 1932 1112
rect 1926 1107 1927 1111
rect 1931 1110 1932 1111
rect 1982 1111 1983 1115
rect 1987 1111 1988 1115
rect 1982 1110 1988 1111
rect 2110 1115 2116 1116
rect 2110 1111 2111 1115
rect 2115 1111 2116 1115
rect 2110 1110 2116 1111
rect 2246 1115 2252 1116
rect 2246 1111 2247 1115
rect 2251 1111 2252 1115
rect 2246 1110 2252 1111
rect 2382 1115 2388 1116
rect 2382 1111 2383 1115
rect 2387 1111 2388 1115
rect 2382 1110 2388 1111
rect 2510 1115 2516 1116
rect 2510 1111 2511 1115
rect 2515 1111 2516 1115
rect 2510 1110 2516 1111
rect 2638 1115 2644 1116
rect 2638 1111 2639 1115
rect 2643 1111 2644 1115
rect 2638 1110 2644 1111
rect 2758 1115 2764 1116
rect 2758 1111 2759 1115
rect 2763 1111 2764 1115
rect 2758 1110 2764 1111
rect 2870 1115 2876 1116
rect 2870 1111 2871 1115
rect 2875 1111 2876 1115
rect 2870 1110 2876 1111
rect 2974 1115 2980 1116
rect 2974 1111 2975 1115
rect 2979 1111 2980 1115
rect 2974 1110 2980 1111
rect 3078 1115 3084 1116
rect 3078 1111 3079 1115
rect 3083 1111 3084 1115
rect 3078 1110 3084 1111
rect 3182 1115 3188 1116
rect 3182 1111 3183 1115
rect 3187 1111 3188 1115
rect 3182 1110 3188 1111
rect 3278 1115 3284 1116
rect 3278 1111 3279 1115
rect 3283 1111 3284 1115
rect 3278 1110 3284 1111
rect 3366 1115 3372 1116
rect 3366 1111 3367 1115
rect 3371 1111 3372 1115
rect 3462 1112 3463 1116
rect 3467 1112 3468 1116
rect 3462 1111 3468 1112
rect 3366 1110 3372 1111
rect 1931 1108 1938 1110
rect 1931 1107 1932 1108
rect 1926 1106 1932 1107
rect 1936 1105 1938 1108
rect 1942 1107 1948 1108
rect 1942 1103 1943 1107
rect 1947 1106 1948 1107
rect 2062 1107 2068 1108
rect 1947 1104 2025 1106
rect 1947 1103 1948 1104
rect 1942 1102 1948 1103
rect 2062 1103 2063 1107
rect 2067 1106 2068 1107
rect 2190 1107 2196 1108
rect 2067 1104 2153 1106
rect 2067 1103 2068 1104
rect 2062 1102 2068 1103
rect 2190 1103 2191 1107
rect 2195 1106 2196 1107
rect 2327 1107 2333 1108
rect 2195 1104 2289 1106
rect 2195 1103 2196 1104
rect 2190 1102 2196 1103
rect 2327 1103 2328 1107
rect 2332 1106 2333 1107
rect 2942 1107 2948 1108
rect 2332 1104 2425 1106
rect 2332 1103 2333 1104
rect 2327 1102 2333 1103
rect 2582 1103 2588 1104
rect 110 1100 116 1101
rect 1766 1100 1772 1101
rect 110 1096 111 1100
rect 115 1096 116 1100
rect 110 1095 116 1096
rect 190 1099 196 1100
rect 190 1095 191 1099
rect 195 1095 196 1099
rect 190 1094 196 1095
rect 334 1099 340 1100
rect 334 1095 335 1099
rect 339 1095 340 1099
rect 334 1094 340 1095
rect 494 1099 500 1100
rect 494 1095 495 1099
rect 499 1095 500 1099
rect 494 1094 500 1095
rect 654 1099 660 1100
rect 654 1095 655 1099
rect 659 1095 660 1099
rect 654 1094 660 1095
rect 814 1099 820 1100
rect 814 1095 815 1099
rect 819 1095 820 1099
rect 814 1094 820 1095
rect 966 1099 972 1100
rect 966 1095 967 1099
rect 971 1095 972 1099
rect 966 1094 972 1095
rect 1118 1099 1124 1100
rect 1118 1095 1119 1099
rect 1123 1095 1124 1099
rect 1118 1094 1124 1095
rect 1262 1099 1268 1100
rect 1262 1095 1263 1099
rect 1267 1095 1268 1099
rect 1262 1094 1268 1095
rect 1406 1099 1412 1100
rect 1406 1095 1407 1099
rect 1411 1095 1412 1099
rect 1406 1094 1412 1095
rect 1558 1099 1564 1100
rect 1558 1095 1559 1099
rect 1563 1095 1564 1099
rect 1766 1096 1767 1100
rect 1771 1096 1772 1100
rect 1766 1095 1772 1096
rect 1806 1099 1812 1100
rect 1806 1095 1807 1099
rect 1811 1095 1812 1099
rect 2582 1099 2583 1103
rect 2587 1099 2588 1103
rect 2582 1098 2588 1099
rect 2710 1103 2716 1104
rect 2710 1099 2711 1103
rect 2715 1099 2716 1103
rect 2710 1098 2716 1099
rect 2830 1103 2836 1104
rect 2830 1099 2831 1103
rect 2835 1099 2836 1103
rect 2942 1103 2943 1107
rect 2947 1103 2948 1107
rect 2942 1102 2948 1103
rect 2950 1107 2956 1108
rect 2950 1103 2951 1107
rect 2955 1106 2956 1107
rect 3054 1107 3060 1108
rect 2955 1104 3017 1106
rect 2955 1103 2956 1104
rect 2950 1102 2956 1103
rect 3054 1103 3055 1107
rect 3059 1106 3060 1107
rect 3158 1107 3164 1108
rect 3059 1104 3121 1106
rect 3059 1103 3060 1104
rect 3054 1102 3060 1103
rect 3158 1103 3159 1107
rect 3163 1106 3164 1107
rect 3262 1107 3268 1108
rect 3163 1104 3225 1106
rect 3163 1103 3164 1104
rect 3158 1102 3164 1103
rect 3262 1103 3263 1107
rect 3267 1106 3268 1107
rect 3359 1107 3365 1108
rect 3267 1104 3321 1106
rect 3267 1103 3268 1104
rect 3262 1102 3268 1103
rect 3359 1103 3360 1107
rect 3364 1106 3365 1107
rect 3364 1104 3409 1106
rect 3364 1103 3365 1104
rect 3359 1102 3365 1103
rect 2830 1098 2836 1099
rect 3462 1099 3468 1100
rect 1558 1094 1564 1095
rect 1806 1094 1812 1095
rect 1862 1096 1868 1097
rect 1862 1092 1863 1096
rect 1867 1092 1868 1096
rect 182 1091 188 1092
rect 182 1087 183 1091
rect 187 1090 188 1091
rect 270 1091 276 1092
rect 187 1088 233 1090
rect 187 1087 188 1088
rect 182 1086 188 1087
rect 270 1087 271 1091
rect 275 1090 276 1091
rect 414 1091 420 1092
rect 275 1088 377 1090
rect 275 1087 276 1088
rect 270 1086 276 1087
rect 414 1087 415 1091
rect 419 1090 420 1091
rect 766 1091 772 1092
rect 419 1088 537 1090
rect 419 1087 420 1088
rect 414 1086 420 1087
rect 726 1087 732 1088
rect 110 1083 116 1084
rect 110 1079 111 1083
rect 115 1079 116 1083
rect 726 1083 727 1087
rect 731 1083 732 1087
rect 766 1087 767 1091
rect 771 1090 772 1091
rect 1527 1091 1533 1092
rect 1862 1091 1868 1092
rect 1982 1096 1988 1097
rect 1982 1092 1983 1096
rect 1987 1092 1988 1096
rect 1982 1091 1988 1092
rect 2110 1096 2116 1097
rect 2110 1092 2111 1096
rect 2115 1092 2116 1096
rect 2110 1091 2116 1092
rect 2246 1096 2252 1097
rect 2246 1092 2247 1096
rect 2251 1092 2252 1096
rect 2246 1091 2252 1092
rect 2382 1096 2388 1097
rect 2382 1092 2383 1096
rect 2387 1092 2388 1096
rect 2382 1091 2388 1092
rect 2510 1096 2516 1097
rect 2510 1092 2511 1096
rect 2515 1092 2516 1096
rect 2510 1091 2516 1092
rect 2638 1096 2644 1097
rect 2638 1092 2639 1096
rect 2643 1092 2644 1096
rect 2638 1091 2644 1092
rect 2758 1096 2764 1097
rect 2758 1092 2759 1096
rect 2763 1092 2764 1096
rect 2758 1091 2764 1092
rect 2870 1096 2876 1097
rect 2870 1092 2871 1096
rect 2875 1092 2876 1096
rect 2870 1091 2876 1092
rect 2974 1096 2980 1097
rect 2974 1092 2975 1096
rect 2979 1092 2980 1096
rect 2974 1091 2980 1092
rect 3078 1096 3084 1097
rect 3078 1092 3079 1096
rect 3083 1092 3084 1096
rect 3078 1091 3084 1092
rect 3182 1096 3188 1097
rect 3182 1092 3183 1096
rect 3187 1092 3188 1096
rect 3182 1091 3188 1092
rect 3278 1096 3284 1097
rect 3278 1092 3279 1096
rect 3283 1092 3284 1096
rect 3278 1091 3284 1092
rect 3366 1096 3372 1097
rect 3366 1092 3367 1096
rect 3371 1092 3372 1096
rect 3462 1095 3463 1099
rect 3467 1095 3468 1099
rect 3462 1094 3468 1095
rect 3366 1091 3372 1092
rect 771 1088 857 1090
rect 771 1087 772 1088
rect 766 1086 772 1087
rect 1038 1087 1044 1088
rect 726 1082 732 1083
rect 1038 1083 1039 1087
rect 1043 1083 1044 1087
rect 1038 1082 1044 1083
rect 1190 1087 1196 1088
rect 1190 1083 1191 1087
rect 1195 1083 1196 1087
rect 1190 1082 1196 1083
rect 1334 1087 1340 1088
rect 1334 1083 1335 1087
rect 1339 1083 1340 1087
rect 1334 1082 1340 1083
rect 1478 1087 1484 1088
rect 1478 1083 1479 1087
rect 1483 1083 1484 1087
rect 1527 1087 1528 1091
rect 1532 1090 1533 1091
rect 1532 1088 1601 1090
rect 1532 1087 1533 1088
rect 1527 1086 1533 1087
rect 2950 1087 2956 1088
rect 2950 1086 2951 1087
rect 2692 1084 2951 1086
rect 1478 1082 1484 1083
rect 1766 1083 1772 1084
rect 110 1078 116 1079
rect 190 1080 196 1081
rect 190 1076 191 1080
rect 195 1076 196 1080
rect 190 1075 196 1076
rect 334 1080 340 1081
rect 334 1076 335 1080
rect 339 1076 340 1080
rect 334 1075 340 1076
rect 494 1080 500 1081
rect 494 1076 495 1080
rect 499 1076 500 1080
rect 494 1075 500 1076
rect 654 1080 660 1081
rect 654 1076 655 1080
rect 659 1076 660 1080
rect 654 1075 660 1076
rect 814 1080 820 1081
rect 814 1076 815 1080
rect 819 1076 820 1080
rect 814 1075 820 1076
rect 966 1080 972 1081
rect 966 1076 967 1080
rect 971 1076 972 1080
rect 966 1075 972 1076
rect 1118 1080 1124 1081
rect 1118 1076 1119 1080
rect 1123 1076 1124 1080
rect 1118 1075 1124 1076
rect 1262 1080 1268 1081
rect 1262 1076 1263 1080
rect 1267 1076 1268 1080
rect 1262 1075 1268 1076
rect 1406 1080 1412 1081
rect 1406 1076 1407 1080
rect 1411 1076 1412 1080
rect 1406 1075 1412 1076
rect 1558 1080 1564 1081
rect 1558 1076 1559 1080
rect 1563 1076 1564 1080
rect 1766 1079 1767 1083
rect 1771 1079 1772 1083
rect 2692 1082 2694 1084
rect 2950 1083 2951 1084
rect 2955 1083 2956 1087
rect 2950 1082 2956 1083
rect 2691 1081 2697 1082
rect 1766 1078 1772 1079
rect 1915 1079 1921 1080
rect 1558 1075 1564 1076
rect 1915 1075 1916 1079
rect 1920 1078 1921 1079
rect 1942 1079 1948 1080
rect 1942 1078 1943 1079
rect 1920 1076 1943 1078
rect 1920 1075 1921 1076
rect 1915 1074 1921 1075
rect 1942 1075 1943 1076
rect 1947 1075 1948 1079
rect 1942 1074 1948 1075
rect 2035 1079 2041 1080
rect 2035 1075 2036 1079
rect 2040 1078 2041 1079
rect 2062 1079 2068 1080
rect 2062 1078 2063 1079
rect 2040 1076 2063 1078
rect 2040 1075 2041 1076
rect 2035 1074 2041 1075
rect 2062 1075 2063 1076
rect 2067 1075 2068 1079
rect 2062 1074 2068 1075
rect 2163 1079 2169 1080
rect 2163 1075 2164 1079
rect 2168 1078 2169 1079
rect 2190 1079 2196 1080
rect 2190 1078 2191 1079
rect 2168 1076 2191 1078
rect 2168 1075 2169 1076
rect 2163 1074 2169 1075
rect 2190 1075 2191 1076
rect 2195 1075 2196 1079
rect 2190 1074 2196 1075
rect 2299 1079 2305 1080
rect 2299 1075 2300 1079
rect 2304 1078 2305 1079
rect 2327 1079 2333 1080
rect 2327 1078 2328 1079
rect 2304 1076 2328 1078
rect 2304 1075 2305 1076
rect 2299 1074 2305 1075
rect 2327 1075 2328 1076
rect 2332 1075 2333 1079
rect 2327 1074 2333 1075
rect 2350 1079 2356 1080
rect 2350 1075 2351 1079
rect 2355 1078 2356 1079
rect 2435 1079 2441 1080
rect 2435 1078 2436 1079
rect 2355 1076 2436 1078
rect 2355 1075 2356 1076
rect 2350 1074 2356 1075
rect 2435 1075 2436 1076
rect 2440 1075 2441 1079
rect 2435 1074 2441 1075
rect 2563 1079 2569 1080
rect 2563 1075 2564 1079
rect 2568 1078 2569 1079
rect 2606 1079 2612 1080
rect 2606 1078 2607 1079
rect 2568 1076 2607 1078
rect 2568 1075 2569 1076
rect 2563 1074 2569 1075
rect 2606 1075 2607 1076
rect 2611 1075 2612 1079
rect 2691 1077 2692 1081
rect 2696 1077 2697 1081
rect 2691 1076 2697 1077
rect 2710 1079 2716 1080
rect 2606 1074 2612 1075
rect 2710 1075 2711 1079
rect 2715 1078 2716 1079
rect 2811 1079 2817 1080
rect 2811 1078 2812 1079
rect 2715 1076 2812 1078
rect 2715 1075 2716 1076
rect 2710 1074 2716 1075
rect 2811 1075 2812 1076
rect 2816 1075 2817 1079
rect 2811 1074 2817 1075
rect 2830 1079 2836 1080
rect 2830 1075 2831 1079
rect 2835 1078 2836 1079
rect 2923 1079 2929 1080
rect 2923 1078 2924 1079
rect 2835 1076 2924 1078
rect 2835 1075 2836 1076
rect 2830 1074 2836 1075
rect 2923 1075 2924 1076
rect 2928 1075 2929 1079
rect 2923 1074 2929 1075
rect 3027 1079 3033 1080
rect 3027 1075 3028 1079
rect 3032 1078 3033 1079
rect 3054 1079 3060 1080
rect 3054 1078 3055 1079
rect 3032 1076 3055 1078
rect 3032 1075 3033 1076
rect 3027 1074 3033 1075
rect 3054 1075 3055 1076
rect 3059 1075 3060 1079
rect 3054 1074 3060 1075
rect 3131 1079 3137 1080
rect 3131 1075 3132 1079
rect 3136 1078 3137 1079
rect 3158 1079 3164 1080
rect 3158 1078 3159 1079
rect 3136 1076 3159 1078
rect 3136 1075 3137 1076
rect 3131 1074 3137 1075
rect 3158 1075 3159 1076
rect 3163 1075 3164 1079
rect 3158 1074 3164 1075
rect 3235 1079 3241 1080
rect 3235 1075 3236 1079
rect 3240 1078 3241 1079
rect 3262 1079 3268 1080
rect 3262 1078 3263 1079
rect 3240 1076 3263 1078
rect 3240 1075 3241 1076
rect 3235 1074 3241 1075
rect 3262 1075 3263 1076
rect 3267 1075 3268 1079
rect 3262 1074 3268 1075
rect 3331 1079 3337 1080
rect 3331 1075 3332 1079
rect 3336 1078 3337 1079
rect 3359 1079 3365 1080
rect 3359 1078 3360 1079
rect 3336 1076 3360 1078
rect 3336 1075 3337 1076
rect 3331 1074 3337 1075
rect 3359 1075 3360 1076
rect 3364 1075 3365 1079
rect 3359 1074 3365 1075
rect 3419 1079 3425 1080
rect 3419 1075 3420 1079
rect 3424 1078 3425 1079
rect 3438 1079 3444 1080
rect 3438 1078 3439 1079
rect 3424 1076 3439 1078
rect 3424 1075 3425 1076
rect 3419 1074 3425 1075
rect 3438 1075 3439 1076
rect 3443 1075 3444 1079
rect 3438 1074 3444 1075
rect 766 1071 772 1072
rect 766 1070 767 1071
rect 548 1068 767 1070
rect 548 1066 550 1068
rect 766 1067 767 1068
rect 771 1067 772 1071
rect 1278 1071 1284 1072
rect 1278 1070 1279 1071
rect 766 1066 772 1067
rect 1020 1068 1279 1070
rect 1020 1066 1022 1068
rect 1278 1067 1279 1068
rect 1283 1067 1284 1071
rect 1278 1066 1284 1067
rect 2174 1067 2180 1068
rect 547 1065 553 1066
rect 243 1063 249 1064
rect 243 1059 244 1063
rect 248 1062 249 1063
rect 270 1063 276 1064
rect 270 1062 271 1063
rect 248 1060 271 1062
rect 248 1059 249 1060
rect 243 1058 249 1059
rect 270 1059 271 1060
rect 275 1059 276 1063
rect 270 1058 276 1059
rect 387 1063 393 1064
rect 387 1059 388 1063
rect 392 1062 393 1063
rect 414 1063 420 1064
rect 414 1062 415 1063
rect 392 1060 415 1062
rect 392 1059 393 1060
rect 387 1058 393 1059
rect 414 1059 415 1060
rect 419 1059 420 1063
rect 547 1061 548 1065
rect 552 1061 553 1065
rect 1019 1065 1025 1066
rect 547 1060 553 1061
rect 678 1063 684 1064
rect 414 1058 420 1059
rect 678 1059 679 1063
rect 683 1062 684 1063
rect 707 1063 713 1064
rect 707 1062 708 1063
rect 683 1060 708 1062
rect 683 1059 684 1060
rect 678 1058 684 1059
rect 707 1059 708 1060
rect 712 1059 713 1063
rect 707 1058 713 1059
rect 726 1063 732 1064
rect 726 1059 727 1063
rect 731 1062 732 1063
rect 867 1063 873 1064
rect 867 1062 868 1063
rect 731 1060 868 1062
rect 731 1059 732 1060
rect 726 1058 732 1059
rect 867 1059 868 1060
rect 872 1059 873 1063
rect 1019 1061 1020 1065
rect 1024 1061 1025 1065
rect 1019 1060 1025 1061
rect 1038 1063 1044 1064
rect 867 1058 873 1059
rect 1038 1059 1039 1063
rect 1043 1062 1044 1063
rect 1171 1063 1177 1064
rect 1171 1062 1172 1063
rect 1043 1060 1172 1062
rect 1043 1059 1044 1060
rect 1038 1058 1044 1059
rect 1171 1059 1172 1060
rect 1176 1059 1177 1063
rect 1171 1058 1177 1059
rect 1190 1063 1196 1064
rect 1190 1059 1191 1063
rect 1195 1062 1196 1063
rect 1315 1063 1321 1064
rect 1315 1062 1316 1063
rect 1195 1060 1316 1062
rect 1195 1059 1196 1060
rect 1190 1058 1196 1059
rect 1315 1059 1316 1060
rect 1320 1059 1321 1063
rect 1315 1058 1321 1059
rect 1334 1063 1340 1064
rect 1334 1059 1335 1063
rect 1339 1062 1340 1063
rect 1459 1063 1465 1064
rect 1459 1062 1460 1063
rect 1339 1060 1460 1062
rect 1339 1059 1340 1060
rect 1334 1058 1340 1059
rect 1459 1059 1460 1060
rect 1464 1059 1465 1063
rect 1459 1058 1465 1059
rect 1478 1063 1484 1064
rect 1478 1059 1479 1063
rect 1483 1062 1484 1063
rect 1611 1063 1617 1064
rect 1611 1062 1612 1063
rect 1483 1060 1612 1062
rect 1483 1059 1484 1060
rect 1478 1058 1484 1059
rect 1611 1059 1612 1060
rect 1616 1059 1617 1063
rect 2174 1063 2175 1067
rect 2179 1066 2180 1067
rect 2179 1064 2247 1066
rect 2179 1063 2180 1064
rect 2174 1062 2180 1063
rect 2245 1062 2247 1064
rect 2243 1061 2249 1062
rect 1611 1058 1617 1059
rect 2155 1059 2161 1060
rect 2155 1055 2156 1059
rect 2160 1058 2161 1059
rect 2160 1056 2238 1058
rect 2243 1057 2244 1061
rect 2248 1057 2249 1061
rect 2243 1056 2249 1057
rect 2262 1059 2268 1060
rect 2160 1055 2161 1056
rect 2155 1054 2161 1055
rect 398 1051 404 1052
rect 398 1047 399 1051
rect 403 1050 404 1051
rect 1527 1051 1533 1052
rect 1527 1050 1528 1051
rect 403 1048 518 1050
rect 403 1047 404 1048
rect 398 1046 404 1047
rect 516 1046 518 1048
rect 1284 1048 1528 1050
rect 1284 1046 1286 1048
rect 1527 1047 1528 1048
rect 1532 1047 1533 1051
rect 2236 1050 2238 1056
rect 2262 1055 2263 1059
rect 2267 1058 2268 1059
rect 2331 1059 2337 1060
rect 2331 1058 2332 1059
rect 2267 1056 2332 1058
rect 2267 1055 2268 1056
rect 2262 1054 2268 1055
rect 2331 1055 2332 1056
rect 2336 1055 2337 1059
rect 2331 1054 2337 1055
rect 2419 1059 2425 1060
rect 2419 1055 2420 1059
rect 2424 1058 2425 1059
rect 2446 1059 2452 1060
rect 2446 1058 2447 1059
rect 2424 1056 2447 1058
rect 2424 1055 2425 1056
rect 2419 1054 2425 1055
rect 2446 1055 2447 1056
rect 2451 1055 2452 1059
rect 2446 1054 2452 1055
rect 2502 1059 2513 1060
rect 2502 1055 2503 1059
rect 2507 1055 2508 1059
rect 2512 1055 2513 1059
rect 2502 1054 2513 1055
rect 2582 1059 2588 1060
rect 2582 1055 2583 1059
rect 2587 1058 2588 1059
rect 2595 1059 2601 1060
rect 2595 1058 2596 1059
rect 2587 1056 2596 1058
rect 2587 1055 2588 1056
rect 2582 1054 2588 1055
rect 2595 1055 2596 1056
rect 2600 1055 2601 1059
rect 2595 1054 2601 1055
rect 2614 1059 2620 1060
rect 2614 1055 2615 1059
rect 2619 1058 2620 1059
rect 2683 1059 2689 1060
rect 2683 1058 2684 1059
rect 2619 1056 2684 1058
rect 2619 1055 2620 1056
rect 2614 1054 2620 1055
rect 2683 1055 2684 1056
rect 2688 1055 2689 1059
rect 2683 1054 2689 1055
rect 2702 1059 2708 1060
rect 2702 1055 2703 1059
rect 2707 1058 2708 1059
rect 2771 1059 2777 1060
rect 2771 1058 2772 1059
rect 2707 1056 2772 1058
rect 2707 1055 2708 1056
rect 2702 1054 2708 1055
rect 2771 1055 2772 1056
rect 2776 1055 2777 1059
rect 2771 1054 2777 1055
rect 2790 1059 2796 1060
rect 2790 1055 2791 1059
rect 2795 1058 2796 1059
rect 2859 1059 2865 1060
rect 2859 1058 2860 1059
rect 2795 1056 2860 1058
rect 2795 1055 2796 1056
rect 2790 1054 2796 1055
rect 2859 1055 2860 1056
rect 2864 1055 2865 1059
rect 2859 1054 2865 1055
rect 2236 1048 2361 1050
rect 1527 1046 1533 1047
rect 515 1045 521 1046
rect 379 1043 385 1044
rect 379 1039 380 1043
rect 384 1042 385 1043
rect 384 1040 510 1042
rect 515 1041 516 1045
rect 520 1041 521 1045
rect 1283 1045 1289 1046
rect 515 1040 521 1041
rect 534 1043 540 1044
rect 384 1039 385 1040
rect 379 1038 385 1039
rect 508 1034 510 1040
rect 534 1039 535 1043
rect 539 1042 540 1043
rect 659 1043 665 1044
rect 659 1042 660 1043
rect 539 1040 660 1042
rect 539 1039 540 1040
rect 534 1038 540 1039
rect 659 1039 660 1040
rect 664 1039 665 1043
rect 659 1038 665 1039
rect 819 1043 825 1044
rect 819 1039 820 1043
rect 824 1042 825 1043
rect 846 1043 852 1044
rect 846 1042 847 1043
rect 824 1040 847 1042
rect 824 1039 825 1040
rect 819 1038 825 1039
rect 846 1039 847 1040
rect 851 1039 852 1043
rect 846 1038 852 1039
rect 958 1043 964 1044
rect 958 1039 959 1043
rect 963 1042 964 1043
rect 979 1043 985 1044
rect 979 1042 980 1043
rect 963 1040 980 1042
rect 963 1039 964 1040
rect 958 1038 964 1039
rect 979 1039 980 1040
rect 984 1039 985 1043
rect 979 1038 985 1039
rect 1131 1043 1137 1044
rect 1131 1039 1132 1043
rect 1136 1042 1137 1043
rect 1158 1043 1164 1044
rect 1158 1042 1159 1043
rect 1136 1040 1159 1042
rect 1136 1039 1137 1040
rect 1131 1038 1137 1039
rect 1158 1039 1159 1040
rect 1163 1039 1164 1043
rect 1283 1041 1284 1045
rect 1288 1041 1289 1045
rect 2102 1044 2108 1045
rect 1283 1040 1289 1041
rect 1435 1043 1441 1044
rect 1158 1038 1164 1039
rect 1435 1039 1436 1043
rect 1440 1042 1441 1043
rect 1462 1043 1468 1044
rect 1462 1042 1463 1043
rect 1440 1040 1463 1042
rect 1440 1039 1441 1040
rect 1435 1038 1441 1039
rect 1462 1039 1463 1040
rect 1467 1039 1468 1043
rect 1462 1038 1468 1039
rect 1470 1043 1476 1044
rect 1470 1039 1471 1043
rect 1475 1042 1476 1043
rect 1587 1043 1593 1044
rect 1587 1042 1588 1043
rect 1475 1040 1588 1042
rect 1475 1039 1476 1040
rect 1470 1038 1476 1039
rect 1587 1039 1588 1040
rect 1592 1039 1593 1043
rect 1587 1038 1593 1039
rect 1606 1043 1612 1044
rect 1606 1039 1607 1043
rect 1611 1042 1612 1043
rect 1723 1043 1729 1044
rect 1723 1042 1724 1043
rect 1611 1040 1724 1042
rect 1611 1039 1612 1040
rect 1606 1038 1612 1039
rect 1723 1039 1724 1040
rect 1728 1039 1729 1043
rect 1723 1038 1729 1039
rect 1806 1041 1812 1042
rect 1806 1037 1807 1041
rect 1811 1037 1812 1041
rect 2102 1040 2103 1044
rect 2107 1040 2108 1044
rect 2102 1039 2108 1040
rect 2190 1044 2196 1045
rect 2190 1040 2191 1044
rect 2195 1040 2196 1044
rect 2190 1039 2196 1040
rect 2278 1044 2284 1045
rect 2278 1040 2279 1044
rect 2283 1040 2284 1044
rect 2278 1039 2284 1040
rect 1806 1036 1812 1037
rect 2174 1035 2180 1036
rect 508 1032 746 1034
rect 326 1028 332 1029
rect 110 1025 116 1026
rect 110 1021 111 1025
rect 115 1021 116 1025
rect 326 1024 327 1028
rect 331 1024 332 1028
rect 326 1023 332 1024
rect 462 1028 468 1029
rect 462 1024 463 1028
rect 467 1024 468 1028
rect 462 1023 468 1024
rect 606 1028 612 1029
rect 606 1024 607 1028
rect 611 1024 612 1028
rect 606 1023 612 1024
rect 110 1020 116 1021
rect 398 1019 404 1020
rect 398 1015 399 1019
rect 403 1015 404 1019
rect 398 1014 404 1015
rect 534 1019 540 1020
rect 534 1015 535 1019
rect 539 1015 540 1019
rect 534 1014 540 1015
rect 678 1019 684 1020
rect 678 1015 679 1019
rect 683 1015 684 1019
rect 744 1018 746 1032
rect 2174 1031 2175 1035
rect 2179 1031 2180 1035
rect 2174 1030 2180 1031
rect 2262 1035 2268 1036
rect 2262 1031 2263 1035
rect 2267 1031 2268 1035
rect 2262 1030 2268 1031
rect 2350 1035 2356 1036
rect 2350 1031 2351 1035
rect 2355 1031 2356 1035
rect 2359 1034 2361 1048
rect 2366 1044 2372 1045
rect 2366 1040 2367 1044
rect 2371 1040 2372 1044
rect 2366 1039 2372 1040
rect 2454 1044 2460 1045
rect 2454 1040 2455 1044
rect 2459 1040 2460 1044
rect 2454 1039 2460 1040
rect 2542 1044 2548 1045
rect 2542 1040 2543 1044
rect 2547 1040 2548 1044
rect 2542 1039 2548 1040
rect 2630 1044 2636 1045
rect 2630 1040 2631 1044
rect 2635 1040 2636 1044
rect 2630 1039 2636 1040
rect 2718 1044 2724 1045
rect 2718 1040 2719 1044
rect 2723 1040 2724 1044
rect 2718 1039 2724 1040
rect 2806 1044 2812 1045
rect 2806 1040 2807 1044
rect 2811 1040 2812 1044
rect 2806 1039 2812 1040
rect 3462 1041 3468 1042
rect 3462 1037 3463 1041
rect 3467 1037 3468 1041
rect 3462 1036 3468 1037
rect 2446 1035 2452 1036
rect 2359 1032 2409 1034
rect 2350 1030 2356 1031
rect 2446 1031 2447 1035
rect 2451 1034 2452 1035
rect 2614 1035 2620 1036
rect 2451 1032 2497 1034
rect 2451 1031 2452 1032
rect 2446 1030 2452 1031
rect 2614 1031 2615 1035
rect 2619 1031 2620 1035
rect 2614 1030 2620 1031
rect 2702 1035 2708 1036
rect 2702 1031 2703 1035
rect 2707 1031 2708 1035
rect 2702 1030 2708 1031
rect 2790 1035 2796 1036
rect 2790 1031 2791 1035
rect 2795 1031 2796 1035
rect 2790 1030 2796 1031
rect 2878 1035 2884 1036
rect 2878 1031 2879 1035
rect 2883 1031 2884 1035
rect 2878 1030 2884 1031
rect 766 1028 772 1029
rect 766 1024 767 1028
rect 771 1024 772 1028
rect 766 1023 772 1024
rect 926 1028 932 1029
rect 926 1024 927 1028
rect 931 1024 932 1028
rect 926 1023 932 1024
rect 1078 1028 1084 1029
rect 1078 1024 1079 1028
rect 1083 1024 1084 1028
rect 1078 1023 1084 1024
rect 1230 1028 1236 1029
rect 1230 1024 1231 1028
rect 1235 1024 1236 1028
rect 1230 1023 1236 1024
rect 1382 1028 1388 1029
rect 1382 1024 1383 1028
rect 1387 1024 1388 1028
rect 1382 1023 1388 1024
rect 1534 1028 1540 1029
rect 1534 1024 1535 1028
rect 1539 1024 1540 1028
rect 1534 1023 1540 1024
rect 1670 1028 1676 1029
rect 1670 1024 1671 1028
rect 1675 1024 1676 1028
rect 1670 1023 1676 1024
rect 1766 1025 1772 1026
rect 2102 1025 2108 1026
rect 1766 1021 1767 1025
rect 1771 1021 1772 1025
rect 1766 1020 1772 1021
rect 1806 1024 1812 1025
rect 1806 1020 1807 1024
rect 1811 1020 1812 1024
rect 2102 1021 2103 1025
rect 2107 1021 2108 1025
rect 2102 1020 2108 1021
rect 2190 1025 2196 1026
rect 2190 1021 2191 1025
rect 2195 1021 2196 1025
rect 2190 1020 2196 1021
rect 2278 1025 2284 1026
rect 2278 1021 2279 1025
rect 2283 1021 2284 1025
rect 2278 1020 2284 1021
rect 2366 1025 2372 1026
rect 2366 1021 2367 1025
rect 2371 1021 2372 1025
rect 2366 1020 2372 1021
rect 2454 1025 2460 1026
rect 2454 1021 2455 1025
rect 2459 1021 2460 1025
rect 2454 1020 2460 1021
rect 2542 1025 2548 1026
rect 2542 1021 2543 1025
rect 2547 1021 2548 1025
rect 2542 1020 2548 1021
rect 2630 1025 2636 1026
rect 2630 1021 2631 1025
rect 2635 1021 2636 1025
rect 2630 1020 2636 1021
rect 2718 1025 2724 1026
rect 2718 1021 2719 1025
rect 2723 1021 2724 1025
rect 2718 1020 2724 1021
rect 2806 1025 2812 1026
rect 2806 1021 2807 1025
rect 2811 1021 2812 1025
rect 2806 1020 2812 1021
rect 3462 1024 3468 1025
rect 3462 1020 3463 1024
rect 3467 1020 3468 1024
rect 846 1019 852 1020
rect 744 1016 809 1018
rect 678 1014 684 1015
rect 846 1015 847 1019
rect 851 1018 852 1019
rect 1046 1019 1052 1020
rect 851 1016 969 1018
rect 851 1015 852 1016
rect 846 1014 852 1015
rect 1046 1015 1047 1019
rect 1051 1018 1052 1019
rect 1158 1019 1164 1020
rect 1051 1016 1121 1018
rect 1051 1015 1052 1016
rect 1046 1014 1052 1015
rect 1158 1015 1159 1019
rect 1163 1018 1164 1019
rect 1470 1019 1476 1020
rect 1470 1018 1471 1019
rect 1163 1016 1273 1018
rect 1457 1016 1471 1018
rect 1163 1015 1164 1016
rect 1158 1014 1164 1015
rect 1470 1015 1471 1016
rect 1475 1015 1476 1019
rect 1470 1014 1476 1015
rect 1606 1019 1612 1020
rect 1606 1015 1607 1019
rect 1611 1015 1612 1019
rect 1606 1014 1612 1015
rect 1614 1019 1620 1020
rect 1806 1019 1812 1020
rect 3462 1019 3468 1020
rect 1614 1015 1615 1019
rect 1619 1018 1620 1019
rect 1619 1016 1713 1018
rect 1619 1015 1620 1016
rect 1614 1014 1620 1015
rect 326 1009 332 1010
rect 110 1008 116 1009
rect 110 1004 111 1008
rect 115 1004 116 1008
rect 326 1005 327 1009
rect 331 1005 332 1009
rect 326 1004 332 1005
rect 462 1009 468 1010
rect 462 1005 463 1009
rect 467 1005 468 1009
rect 462 1004 468 1005
rect 606 1009 612 1010
rect 606 1005 607 1009
rect 611 1005 612 1009
rect 606 1004 612 1005
rect 766 1009 772 1010
rect 766 1005 767 1009
rect 771 1005 772 1009
rect 766 1004 772 1005
rect 926 1009 932 1010
rect 926 1005 927 1009
rect 931 1005 932 1009
rect 926 1004 932 1005
rect 1078 1009 1084 1010
rect 1078 1005 1079 1009
rect 1083 1005 1084 1009
rect 1078 1004 1084 1005
rect 1230 1009 1236 1010
rect 1230 1005 1231 1009
rect 1235 1005 1236 1009
rect 1230 1004 1236 1005
rect 1382 1009 1388 1010
rect 1382 1005 1383 1009
rect 1387 1005 1388 1009
rect 1382 1004 1388 1005
rect 1534 1009 1540 1010
rect 1534 1005 1535 1009
rect 1539 1005 1540 1009
rect 1534 1004 1540 1005
rect 1670 1009 1676 1010
rect 1670 1005 1671 1009
rect 1675 1005 1676 1009
rect 1670 1004 1676 1005
rect 1766 1008 1772 1009
rect 1766 1004 1767 1008
rect 1771 1004 1772 1008
rect 110 1003 116 1004
rect 1766 1003 1772 1004
rect 1806 980 1812 981
rect 3462 980 3468 981
rect 1806 976 1807 980
rect 1811 976 1812 980
rect 1806 975 1812 976
rect 2310 979 2316 980
rect 2310 975 2311 979
rect 2315 975 2316 979
rect 2310 974 2316 975
rect 2406 979 2412 980
rect 2406 975 2407 979
rect 2411 975 2412 979
rect 2406 974 2412 975
rect 2510 979 2516 980
rect 2510 975 2511 979
rect 2515 975 2516 979
rect 2510 974 2516 975
rect 2622 979 2628 980
rect 2622 975 2623 979
rect 2627 975 2628 979
rect 2622 974 2628 975
rect 2750 979 2756 980
rect 2750 975 2751 979
rect 2755 975 2756 979
rect 2750 974 2756 975
rect 2894 979 2900 980
rect 2894 975 2895 979
rect 2899 975 2900 979
rect 2894 974 2900 975
rect 3054 979 3060 980
rect 3054 975 3055 979
rect 3059 975 3060 979
rect 3054 974 3060 975
rect 3222 979 3228 980
rect 3222 975 3223 979
rect 3227 975 3228 979
rect 3222 974 3228 975
rect 3366 979 3372 980
rect 3366 975 3367 979
rect 3371 975 3372 979
rect 3462 976 3463 980
rect 3467 976 3468 980
rect 3462 975 3468 976
rect 3366 974 3372 975
rect 2502 971 2508 972
rect 2382 967 2388 968
rect 1806 963 1812 964
rect 110 960 116 961
rect 1766 960 1772 961
rect 110 956 111 960
rect 115 956 116 960
rect 110 955 116 956
rect 470 959 476 960
rect 470 955 471 959
rect 475 955 476 959
rect 470 954 476 955
rect 566 959 572 960
rect 566 955 567 959
rect 571 955 572 959
rect 566 954 572 955
rect 670 959 676 960
rect 670 955 671 959
rect 675 955 676 959
rect 670 954 676 955
rect 782 959 788 960
rect 782 955 783 959
rect 787 955 788 959
rect 782 954 788 955
rect 886 959 892 960
rect 886 955 887 959
rect 891 955 892 959
rect 886 954 892 955
rect 990 959 996 960
rect 990 955 991 959
rect 995 955 996 959
rect 990 954 996 955
rect 1094 959 1100 960
rect 1094 955 1095 959
rect 1099 955 1100 959
rect 1094 954 1100 955
rect 1198 959 1204 960
rect 1198 955 1199 959
rect 1203 955 1204 959
rect 1198 954 1204 955
rect 1294 959 1300 960
rect 1294 955 1295 959
rect 1299 955 1300 959
rect 1294 954 1300 955
rect 1390 959 1396 960
rect 1390 955 1391 959
rect 1395 955 1396 959
rect 1390 954 1396 955
rect 1486 959 1492 960
rect 1486 955 1487 959
rect 1491 955 1492 959
rect 1486 954 1492 955
rect 1582 959 1588 960
rect 1582 955 1583 959
rect 1587 955 1588 959
rect 1582 954 1588 955
rect 1670 959 1676 960
rect 1670 955 1671 959
rect 1675 955 1676 959
rect 1766 956 1767 960
rect 1771 956 1772 960
rect 1806 959 1807 963
rect 1811 959 1812 963
rect 2382 963 2383 967
rect 2387 963 2388 967
rect 2382 962 2388 963
rect 2478 967 2484 968
rect 2478 963 2479 967
rect 2483 963 2484 967
rect 2502 967 2503 971
rect 2507 970 2508 971
rect 3138 971 3144 972
rect 2507 968 2553 970
rect 2507 967 2508 968
rect 2502 966 2508 967
rect 2694 967 2700 968
rect 2478 962 2484 963
rect 2694 963 2695 967
rect 2699 963 2700 967
rect 2694 962 2700 963
rect 2822 967 2828 968
rect 2822 963 2823 967
rect 2827 963 2828 967
rect 2822 962 2828 963
rect 2966 967 2972 968
rect 2966 963 2967 967
rect 2971 963 2972 967
rect 2966 962 2972 963
rect 3126 967 3132 968
rect 3126 963 3127 967
rect 3131 963 3132 967
rect 3138 967 3139 971
rect 3143 970 3144 971
rect 3438 971 3444 972
rect 3143 968 3265 970
rect 3143 967 3144 968
rect 3138 966 3144 967
rect 3438 967 3439 971
rect 3443 967 3444 971
rect 3438 966 3444 967
rect 3126 962 3132 963
rect 3462 963 3468 964
rect 1806 958 1812 959
rect 2310 960 2316 961
rect 1766 955 1772 956
rect 2310 956 2311 960
rect 2315 956 2316 960
rect 2310 955 2316 956
rect 2406 960 2412 961
rect 2406 956 2407 960
rect 2411 956 2412 960
rect 2406 955 2412 956
rect 2510 960 2516 961
rect 2510 956 2511 960
rect 2515 956 2516 960
rect 2510 955 2516 956
rect 2622 960 2628 961
rect 2622 956 2623 960
rect 2627 956 2628 960
rect 2622 955 2628 956
rect 2750 960 2756 961
rect 2750 956 2751 960
rect 2755 956 2756 960
rect 2750 955 2756 956
rect 2894 960 2900 961
rect 2894 956 2895 960
rect 2899 956 2900 960
rect 2894 955 2900 956
rect 3054 960 3060 961
rect 3054 956 3055 960
rect 3059 956 3060 960
rect 3054 955 3060 956
rect 3222 960 3228 961
rect 3222 956 3223 960
rect 3227 956 3228 960
rect 3222 955 3228 956
rect 3366 960 3372 961
rect 3366 956 3367 960
rect 3371 956 3372 960
rect 3462 959 3463 963
rect 3467 959 3468 963
rect 3462 958 3468 959
rect 3366 955 3372 956
rect 1670 954 1676 955
rect 958 951 964 952
rect 542 947 548 948
rect 110 943 116 944
rect 110 939 111 943
rect 115 939 116 943
rect 542 943 543 947
rect 547 943 548 947
rect 542 942 548 943
rect 638 947 644 948
rect 638 943 639 947
rect 643 943 644 947
rect 638 942 644 943
rect 742 947 748 948
rect 742 943 743 947
rect 747 943 748 947
rect 742 942 748 943
rect 854 947 860 948
rect 854 943 855 947
rect 859 943 860 947
rect 958 947 959 951
rect 963 947 964 951
rect 1462 951 1468 952
rect 958 946 964 947
rect 1062 947 1068 948
rect 854 942 860 943
rect 1062 943 1063 947
rect 1067 943 1068 947
rect 1062 942 1068 943
rect 1166 947 1172 948
rect 1166 943 1167 947
rect 1171 943 1172 947
rect 1166 942 1172 943
rect 1270 947 1276 948
rect 1270 943 1271 947
rect 1275 943 1276 947
rect 1270 942 1276 943
rect 1366 947 1372 948
rect 1366 943 1367 947
rect 1371 943 1372 947
rect 1462 947 1463 951
rect 1467 947 1468 951
rect 3138 951 3144 952
rect 3138 950 3139 951
rect 2676 948 3139 950
rect 1462 946 1468 947
rect 1558 947 1564 948
rect 1366 942 1372 943
rect 1558 943 1559 947
rect 1563 943 1564 947
rect 1558 942 1564 943
rect 1654 947 1660 948
rect 1654 943 1655 947
rect 1659 943 1660 947
rect 1654 942 1660 943
rect 1742 947 1748 948
rect 1742 943 1743 947
rect 1747 943 1748 947
rect 2676 946 2678 948
rect 3138 947 3139 948
rect 3143 947 3144 951
rect 3138 946 3144 947
rect 2675 945 2681 946
rect 1742 942 1748 943
rect 1766 943 1772 944
rect 110 938 116 939
rect 470 940 476 941
rect 470 936 471 940
rect 475 936 476 940
rect 470 935 476 936
rect 566 940 572 941
rect 566 936 567 940
rect 571 936 572 940
rect 566 935 572 936
rect 670 940 676 941
rect 670 936 671 940
rect 675 936 676 940
rect 670 935 676 936
rect 782 940 788 941
rect 782 936 783 940
rect 787 936 788 940
rect 782 935 788 936
rect 886 940 892 941
rect 886 936 887 940
rect 891 936 892 940
rect 886 935 892 936
rect 990 940 996 941
rect 990 936 991 940
rect 995 936 996 940
rect 990 935 996 936
rect 1094 940 1100 941
rect 1094 936 1095 940
rect 1099 936 1100 940
rect 1094 935 1100 936
rect 1198 940 1204 941
rect 1198 936 1199 940
rect 1203 936 1204 940
rect 1198 935 1204 936
rect 1294 940 1300 941
rect 1294 936 1295 940
rect 1299 936 1300 940
rect 1294 935 1300 936
rect 1390 940 1396 941
rect 1390 936 1391 940
rect 1395 936 1396 940
rect 1390 935 1396 936
rect 1486 940 1492 941
rect 1486 936 1487 940
rect 1491 936 1492 940
rect 1486 935 1492 936
rect 1582 940 1588 941
rect 1582 936 1583 940
rect 1587 936 1588 940
rect 1582 935 1588 936
rect 1670 940 1676 941
rect 1670 936 1671 940
rect 1675 936 1676 940
rect 1766 939 1767 943
rect 1771 939 1772 943
rect 1766 938 1772 939
rect 2222 943 2228 944
rect 2222 939 2223 943
rect 2227 942 2228 943
rect 2363 943 2369 944
rect 2363 942 2364 943
rect 2227 940 2364 942
rect 2227 939 2228 940
rect 2222 938 2228 939
rect 2363 939 2364 940
rect 2368 939 2369 943
rect 2363 938 2369 939
rect 2382 943 2388 944
rect 2382 939 2383 943
rect 2387 942 2388 943
rect 2459 943 2465 944
rect 2459 942 2460 943
rect 2387 940 2460 942
rect 2387 939 2388 940
rect 2382 938 2388 939
rect 2459 939 2460 940
rect 2464 939 2465 943
rect 2459 938 2465 939
rect 2478 943 2484 944
rect 2478 939 2479 943
rect 2483 942 2484 943
rect 2563 943 2569 944
rect 2563 942 2564 943
rect 2483 940 2564 942
rect 2483 939 2484 940
rect 2478 938 2484 939
rect 2563 939 2564 940
rect 2568 939 2569 943
rect 2675 941 2676 945
rect 2680 941 2681 945
rect 2675 940 2681 941
rect 2694 943 2700 944
rect 2563 938 2569 939
rect 2694 939 2695 943
rect 2699 942 2700 943
rect 2803 943 2809 944
rect 2803 942 2804 943
rect 2699 940 2804 942
rect 2699 939 2700 940
rect 2694 938 2700 939
rect 2803 939 2804 940
rect 2808 939 2809 943
rect 2803 938 2809 939
rect 2878 943 2884 944
rect 2878 939 2879 943
rect 2883 942 2884 943
rect 2947 943 2953 944
rect 2947 942 2948 943
rect 2883 940 2948 942
rect 2883 939 2884 940
rect 2878 938 2884 939
rect 2947 939 2948 940
rect 2952 939 2953 943
rect 2947 938 2953 939
rect 2966 943 2972 944
rect 2966 939 2967 943
rect 2971 942 2972 943
rect 3107 943 3113 944
rect 3107 942 3108 943
rect 2971 940 3108 942
rect 2971 939 2972 940
rect 2966 938 2972 939
rect 3107 939 3108 940
rect 3112 939 3113 943
rect 3107 938 3113 939
rect 3126 943 3132 944
rect 3126 939 3127 943
rect 3131 942 3132 943
rect 3275 943 3281 944
rect 3275 942 3276 943
rect 3131 940 3276 942
rect 3131 939 3132 940
rect 3126 938 3132 939
rect 3275 939 3276 940
rect 3280 939 3281 943
rect 3275 938 3281 939
rect 3419 943 3425 944
rect 3419 939 3420 943
rect 3424 942 3425 943
rect 3430 943 3436 944
rect 3430 942 3431 943
rect 3424 940 3431 942
rect 3424 939 3425 940
rect 3419 938 3425 939
rect 3430 939 3431 940
rect 3435 939 3436 943
rect 3430 938 3436 939
rect 1670 935 1676 936
rect 1614 931 1620 932
rect 1614 930 1615 931
rect 1540 928 1615 930
rect 1540 926 1542 928
rect 1614 927 1615 928
rect 1619 927 1620 931
rect 1614 926 1620 927
rect 2822 927 2828 928
rect 1539 925 1545 926
rect 523 923 532 924
rect 523 919 524 923
rect 531 919 532 923
rect 523 918 532 919
rect 542 923 548 924
rect 542 919 543 923
rect 547 922 548 923
rect 619 923 625 924
rect 619 922 620 923
rect 547 920 620 922
rect 547 919 548 920
rect 542 918 548 919
rect 619 919 620 920
rect 624 919 625 923
rect 619 918 625 919
rect 638 923 644 924
rect 638 919 639 923
rect 643 922 644 923
rect 723 923 729 924
rect 723 922 724 923
rect 643 920 724 922
rect 643 919 644 920
rect 638 918 644 919
rect 723 919 724 920
rect 728 919 729 923
rect 723 918 729 919
rect 742 923 748 924
rect 742 919 743 923
rect 747 922 748 923
rect 835 923 841 924
rect 835 922 836 923
rect 747 920 836 922
rect 747 919 748 920
rect 742 918 748 919
rect 835 919 836 920
rect 840 919 841 923
rect 835 918 841 919
rect 854 923 860 924
rect 854 919 855 923
rect 859 922 860 923
rect 939 923 945 924
rect 939 922 940 923
rect 859 920 940 922
rect 859 919 860 920
rect 854 918 860 919
rect 939 919 940 920
rect 944 919 945 923
rect 939 918 945 919
rect 1043 923 1052 924
rect 1043 919 1044 923
rect 1051 919 1052 923
rect 1043 918 1052 919
rect 1147 923 1153 924
rect 1147 919 1148 923
rect 1152 922 1153 923
rect 1166 923 1172 924
rect 1152 920 1162 922
rect 1152 919 1153 920
rect 1147 918 1153 919
rect 1160 914 1162 920
rect 1166 919 1167 923
rect 1171 922 1172 923
rect 1251 923 1257 924
rect 1251 922 1252 923
rect 1171 920 1252 922
rect 1171 919 1172 920
rect 1166 918 1172 919
rect 1251 919 1252 920
rect 1256 919 1257 923
rect 1251 918 1257 919
rect 1270 923 1276 924
rect 1270 919 1271 923
rect 1275 922 1276 923
rect 1347 923 1353 924
rect 1347 922 1348 923
rect 1275 920 1348 922
rect 1275 919 1276 920
rect 1270 918 1276 919
rect 1347 919 1348 920
rect 1352 919 1353 923
rect 1347 918 1353 919
rect 1366 923 1372 924
rect 1366 919 1367 923
rect 1371 922 1372 923
rect 1443 923 1449 924
rect 1443 922 1444 923
rect 1371 920 1444 922
rect 1371 919 1372 920
rect 1366 918 1372 919
rect 1443 919 1444 920
rect 1448 919 1449 923
rect 1539 921 1540 925
rect 1544 921 1545 925
rect 1539 920 1545 921
rect 1558 923 1564 924
rect 1443 918 1449 919
rect 1558 919 1559 923
rect 1563 922 1564 923
rect 1635 923 1641 924
rect 1635 922 1636 923
rect 1563 920 1636 922
rect 1563 919 1564 920
rect 1558 918 1564 919
rect 1635 919 1636 920
rect 1640 919 1641 923
rect 1635 918 1641 919
rect 1654 923 1660 924
rect 1654 919 1655 923
rect 1659 922 1660 923
rect 1723 923 1729 924
rect 1723 922 1724 923
rect 1659 920 1724 922
rect 1659 919 1660 920
rect 1654 918 1660 919
rect 1723 919 1724 920
rect 1728 919 1729 923
rect 2822 923 2823 927
rect 2827 926 2828 927
rect 2827 924 2991 926
rect 2827 923 2828 924
rect 2822 922 2828 923
rect 2989 922 2991 924
rect 2987 921 2993 922
rect 1723 918 1729 919
rect 1742 919 1748 920
rect 1302 915 1308 916
rect 1302 914 1303 915
rect 1160 912 1303 914
rect 1302 911 1303 912
rect 1307 911 1308 915
rect 1742 915 1743 919
rect 1747 918 1748 919
rect 1883 919 1889 920
rect 1883 918 1884 919
rect 1747 916 1884 918
rect 1747 915 1748 916
rect 1742 914 1748 915
rect 1883 915 1884 916
rect 1888 915 1889 919
rect 1883 914 1889 915
rect 2035 919 2044 920
rect 2035 915 2036 919
rect 2043 915 2044 919
rect 2035 914 2044 915
rect 2054 919 2060 920
rect 2054 915 2055 919
rect 2059 918 2060 919
rect 2203 919 2209 920
rect 2203 918 2204 919
rect 2059 916 2204 918
rect 2059 915 2060 916
rect 2054 914 2060 915
rect 2203 915 2204 916
rect 2208 915 2209 919
rect 2203 914 2209 915
rect 2379 919 2385 920
rect 2379 915 2380 919
rect 2384 918 2385 919
rect 2407 919 2413 920
rect 2407 918 2408 919
rect 2384 916 2408 918
rect 2384 915 2385 916
rect 2379 914 2385 915
rect 2407 915 2408 916
rect 2412 915 2413 919
rect 2407 914 2413 915
rect 2571 919 2577 920
rect 2571 915 2572 919
rect 2576 918 2577 919
rect 2598 919 2604 920
rect 2598 918 2599 919
rect 2576 916 2599 918
rect 2576 915 2577 916
rect 2571 914 2577 915
rect 2598 915 2599 916
rect 2603 915 2604 919
rect 2598 914 2604 915
rect 2771 919 2777 920
rect 2771 915 2772 919
rect 2776 918 2777 919
rect 2776 916 2982 918
rect 2987 917 2988 921
rect 2992 917 2993 921
rect 2987 916 2993 917
rect 3006 919 3012 920
rect 2776 915 2777 916
rect 2771 914 2777 915
rect 1302 910 1308 911
rect 659 907 665 908
rect 659 903 660 907
rect 664 906 665 907
rect 687 907 693 908
rect 687 906 688 907
rect 664 904 688 906
rect 664 903 665 904
rect 659 902 665 903
rect 687 903 688 904
rect 692 903 693 907
rect 687 902 693 903
rect 747 907 753 908
rect 747 903 748 907
rect 752 906 753 907
rect 774 907 780 908
rect 774 906 775 907
rect 752 904 775 906
rect 752 903 753 904
rect 747 902 753 903
rect 774 903 775 904
rect 779 903 780 907
rect 774 902 780 903
rect 843 907 849 908
rect 843 903 844 907
rect 848 906 849 907
rect 870 907 876 908
rect 870 906 871 907
rect 848 904 871 906
rect 848 903 849 904
rect 843 902 849 903
rect 870 903 871 904
rect 875 903 876 907
rect 870 902 876 903
rect 947 907 953 908
rect 947 903 948 907
rect 952 906 953 907
rect 975 907 981 908
rect 975 906 976 907
rect 952 904 976 906
rect 952 903 953 904
rect 947 902 953 903
rect 975 903 976 904
rect 980 903 981 907
rect 975 902 981 903
rect 1022 907 1028 908
rect 1022 903 1023 907
rect 1027 906 1028 907
rect 1051 907 1057 908
rect 1051 906 1052 907
rect 1027 904 1052 906
rect 1027 903 1028 904
rect 1022 902 1028 903
rect 1051 903 1052 904
rect 1056 903 1057 907
rect 1051 902 1057 903
rect 1062 907 1068 908
rect 1062 903 1063 907
rect 1067 906 1068 907
rect 1163 907 1169 908
rect 1163 906 1164 907
rect 1067 904 1164 906
rect 1067 903 1068 904
rect 1062 902 1068 903
rect 1163 903 1164 904
rect 1168 903 1169 907
rect 1163 902 1169 903
rect 1182 907 1188 908
rect 1182 903 1183 907
rect 1187 906 1188 907
rect 1275 907 1281 908
rect 1275 906 1276 907
rect 1187 904 1276 906
rect 1187 903 1188 904
rect 1182 902 1188 903
rect 1275 903 1276 904
rect 1280 903 1281 907
rect 1275 902 1281 903
rect 1395 907 1401 908
rect 1395 903 1396 907
rect 1400 906 1401 907
rect 1447 907 1453 908
rect 1447 906 1448 907
rect 1400 904 1448 906
rect 1400 903 1401 904
rect 1395 902 1401 903
rect 1447 903 1448 904
rect 1452 903 1453 907
rect 1447 902 1453 903
rect 1515 907 1521 908
rect 1515 903 1516 907
rect 1520 906 1521 907
rect 1566 907 1572 908
rect 1566 906 1567 907
rect 1520 904 1567 906
rect 1520 903 1521 904
rect 1515 902 1521 903
rect 1566 903 1567 904
rect 1571 903 1572 907
rect 1566 902 1572 903
rect 1630 907 1641 908
rect 1630 903 1631 907
rect 1635 903 1636 907
rect 1640 903 1641 907
rect 2980 906 2982 916
rect 3006 915 3007 919
rect 3011 918 3012 919
rect 3211 919 3217 920
rect 3211 918 3212 919
rect 3011 916 3212 918
rect 3011 915 3012 916
rect 3006 914 3012 915
rect 3211 915 3212 916
rect 3216 915 3217 919
rect 3211 914 3217 915
rect 3419 919 3425 920
rect 3419 915 3420 919
rect 3424 918 3425 919
rect 3438 919 3444 920
rect 3438 918 3439 919
rect 3424 916 3439 918
rect 3424 915 3425 916
rect 3419 914 3425 915
rect 3438 915 3439 916
rect 3443 915 3444 919
rect 3438 914 3444 915
rect 1630 902 1641 903
rect 1830 904 1836 905
rect 1806 901 1812 902
rect 1806 897 1807 901
rect 1811 897 1812 901
rect 1830 900 1831 904
rect 1835 900 1836 904
rect 1830 899 1836 900
rect 1982 904 1988 905
rect 1982 900 1983 904
rect 1987 900 1988 904
rect 1982 899 1988 900
rect 2150 904 2156 905
rect 2150 900 2151 904
rect 2155 900 2156 904
rect 2150 899 2156 900
rect 2326 904 2332 905
rect 2326 900 2327 904
rect 2331 900 2332 904
rect 2326 899 2332 900
rect 2518 904 2524 905
rect 2518 900 2519 904
rect 2523 900 2524 904
rect 2518 899 2524 900
rect 2718 904 2724 905
rect 2718 900 2719 904
rect 2723 900 2724 904
rect 2718 899 2724 900
rect 2934 904 2940 905
rect 2980 904 3014 906
rect 2934 900 2935 904
rect 2939 900 2940 904
rect 3012 902 3014 904
rect 3158 904 3164 905
rect 3012 900 3138 902
rect 2934 899 2940 900
rect 1806 896 1812 897
rect 1894 895 1900 896
rect 606 892 612 893
rect 110 889 116 890
rect 110 885 111 889
rect 115 885 116 889
rect 606 888 607 892
rect 611 888 612 892
rect 606 887 612 888
rect 694 892 700 893
rect 694 888 695 892
rect 699 888 700 892
rect 694 887 700 888
rect 790 892 796 893
rect 790 888 791 892
rect 795 888 796 892
rect 790 887 796 888
rect 894 892 900 893
rect 894 888 895 892
rect 899 888 900 892
rect 894 887 900 888
rect 998 892 1004 893
rect 998 888 999 892
rect 1003 888 1004 892
rect 998 887 1004 888
rect 1110 892 1116 893
rect 1110 888 1111 892
rect 1115 888 1116 892
rect 1110 887 1116 888
rect 1222 892 1228 893
rect 1222 888 1223 892
rect 1227 888 1228 892
rect 1222 887 1228 888
rect 1342 892 1348 893
rect 1342 888 1343 892
rect 1347 888 1348 892
rect 1342 887 1348 888
rect 1462 892 1468 893
rect 1462 888 1463 892
rect 1467 888 1468 892
rect 1462 887 1468 888
rect 1582 892 1588 893
rect 1582 888 1583 892
rect 1587 888 1588 892
rect 1894 891 1895 895
rect 1899 891 1900 895
rect 1894 890 1900 891
rect 2054 895 2060 896
rect 2054 891 2055 895
rect 2059 891 2060 895
rect 2054 890 2060 891
rect 2222 895 2228 896
rect 2222 891 2223 895
rect 2227 891 2228 895
rect 2222 890 2228 891
rect 2398 895 2404 896
rect 2398 891 2399 895
rect 2403 891 2404 895
rect 2398 890 2404 891
rect 2407 895 2413 896
rect 2407 891 2408 895
rect 2412 894 2413 895
rect 2598 895 2604 896
rect 2412 892 2561 894
rect 2412 891 2413 892
rect 2407 890 2413 891
rect 2598 891 2599 895
rect 2603 894 2604 895
rect 3006 895 3012 896
rect 2603 892 2761 894
rect 2603 891 2604 892
rect 2598 890 2604 891
rect 3006 891 3007 895
rect 3011 891 3012 895
rect 3136 894 3138 900
rect 3158 900 3159 904
rect 3163 900 3164 904
rect 3158 899 3164 900
rect 3366 904 3372 905
rect 3366 900 3367 904
rect 3371 900 3372 904
rect 3366 899 3372 900
rect 3462 901 3468 902
rect 3462 897 3463 901
rect 3467 897 3468 901
rect 3462 896 3468 897
rect 3430 895 3436 896
rect 3136 892 3201 894
rect 3006 890 3012 891
rect 3430 891 3431 895
rect 3435 891 3436 895
rect 3430 890 3436 891
rect 1582 887 1588 888
rect 1766 889 1772 890
rect 110 884 116 885
rect 1766 885 1767 889
rect 1771 885 1772 889
rect 1830 885 1836 886
rect 1766 884 1772 885
rect 1806 884 1812 885
rect 526 883 532 884
rect 526 879 527 883
rect 531 882 532 883
rect 687 883 693 884
rect 531 880 649 882
rect 531 879 532 880
rect 526 878 532 879
rect 687 879 688 883
rect 692 882 693 883
rect 774 883 780 884
rect 692 880 737 882
rect 692 879 693 880
rect 687 878 693 879
rect 774 879 775 883
rect 779 882 780 883
rect 870 883 876 884
rect 779 880 833 882
rect 779 879 780 880
rect 774 878 780 879
rect 870 879 871 883
rect 875 882 876 883
rect 975 883 981 884
rect 875 880 937 882
rect 875 879 876 880
rect 870 878 876 879
rect 975 879 976 883
rect 980 882 981 883
rect 1182 883 1188 884
rect 980 880 1041 882
rect 980 879 981 880
rect 975 878 981 879
rect 1182 879 1183 883
rect 1187 879 1188 883
rect 1182 878 1188 879
rect 1198 883 1204 884
rect 1198 879 1199 883
rect 1203 882 1204 883
rect 1302 883 1308 884
rect 1203 880 1265 882
rect 1203 879 1204 880
rect 1198 878 1204 879
rect 1302 879 1303 883
rect 1307 882 1308 883
rect 1447 883 1453 884
rect 1307 880 1385 882
rect 1307 879 1308 880
rect 1302 878 1308 879
rect 1447 879 1448 883
rect 1452 882 1453 883
rect 1566 883 1572 884
rect 1452 880 1505 882
rect 1452 879 1453 880
rect 1447 878 1453 879
rect 1566 879 1567 883
rect 1571 882 1572 883
rect 1571 880 1625 882
rect 1806 880 1807 884
rect 1811 880 1812 884
rect 1830 881 1831 885
rect 1835 881 1836 885
rect 1830 880 1836 881
rect 1982 885 1988 886
rect 1982 881 1983 885
rect 1987 881 1988 885
rect 1982 880 1988 881
rect 2150 885 2156 886
rect 2150 881 2151 885
rect 2155 881 2156 885
rect 2150 880 2156 881
rect 2326 885 2332 886
rect 2326 881 2327 885
rect 2331 881 2332 885
rect 2326 880 2332 881
rect 2518 885 2524 886
rect 2518 881 2519 885
rect 2523 881 2524 885
rect 2518 880 2524 881
rect 2718 885 2724 886
rect 2718 881 2719 885
rect 2723 881 2724 885
rect 2718 880 2724 881
rect 2934 885 2940 886
rect 2934 881 2935 885
rect 2939 881 2940 885
rect 2934 880 2940 881
rect 3158 885 3164 886
rect 3158 881 3159 885
rect 3163 881 3164 885
rect 3158 880 3164 881
rect 3366 885 3372 886
rect 3366 881 3367 885
rect 3371 881 3372 885
rect 3366 880 3372 881
rect 3462 884 3468 885
rect 3462 880 3463 884
rect 3467 880 3468 884
rect 1571 879 1572 880
rect 1806 879 1812 880
rect 3462 879 3468 880
rect 1566 878 1572 879
rect 606 873 612 874
rect 110 872 116 873
rect 110 868 111 872
rect 115 868 116 872
rect 606 869 607 873
rect 611 869 612 873
rect 606 868 612 869
rect 694 873 700 874
rect 694 869 695 873
rect 699 869 700 873
rect 694 868 700 869
rect 790 873 796 874
rect 790 869 791 873
rect 795 869 796 873
rect 790 868 796 869
rect 894 873 900 874
rect 894 869 895 873
rect 899 869 900 873
rect 894 868 900 869
rect 998 873 1004 874
rect 998 869 999 873
rect 1003 869 1004 873
rect 998 868 1004 869
rect 1110 873 1116 874
rect 1110 869 1111 873
rect 1115 869 1116 873
rect 1110 868 1116 869
rect 1222 873 1228 874
rect 1222 869 1223 873
rect 1227 869 1228 873
rect 1222 868 1228 869
rect 1342 873 1348 874
rect 1342 869 1343 873
rect 1347 869 1348 873
rect 1342 868 1348 869
rect 1462 873 1468 874
rect 1462 869 1463 873
rect 1467 869 1468 873
rect 1462 868 1468 869
rect 1582 873 1588 874
rect 1582 869 1583 873
rect 1587 869 1588 873
rect 1582 868 1588 869
rect 1766 872 1772 873
rect 1766 868 1767 872
rect 1771 868 1772 872
rect 110 867 116 868
rect 1766 867 1772 868
rect 1806 836 1812 837
rect 3462 836 3468 837
rect 1806 832 1807 836
rect 1811 832 1812 836
rect 1806 831 1812 832
rect 1830 835 1836 836
rect 1830 831 1831 835
rect 1835 831 1836 835
rect 1830 830 1836 831
rect 1958 835 1964 836
rect 1958 831 1959 835
rect 1963 831 1964 835
rect 1958 830 1964 831
rect 2086 835 2092 836
rect 2086 831 2087 835
rect 2091 831 2092 835
rect 2086 830 2092 831
rect 2206 835 2212 836
rect 2206 831 2207 835
rect 2211 831 2212 835
rect 2206 830 2212 831
rect 2326 835 2332 836
rect 2326 831 2327 835
rect 2331 831 2332 835
rect 2326 830 2332 831
rect 2462 835 2468 836
rect 2462 831 2463 835
rect 2467 831 2468 835
rect 2462 830 2468 831
rect 2614 835 2620 836
rect 2614 831 2615 835
rect 2619 831 2620 835
rect 2614 830 2620 831
rect 2790 835 2796 836
rect 2790 831 2791 835
rect 2795 831 2796 835
rect 2790 830 2796 831
rect 2982 835 2988 836
rect 2982 831 2983 835
rect 2987 831 2988 835
rect 2982 830 2988 831
rect 3182 835 3188 836
rect 3182 831 3183 835
rect 3187 831 3188 835
rect 3182 830 3188 831
rect 3366 835 3372 836
rect 3366 831 3367 835
rect 3371 831 3372 835
rect 3462 832 3463 836
rect 3467 832 3468 836
rect 3462 831 3468 832
rect 3366 830 3372 831
rect 2038 827 2044 828
rect 110 824 116 825
rect 1766 824 1772 825
rect 110 820 111 824
rect 115 820 116 824
rect 110 819 116 820
rect 518 823 524 824
rect 518 819 519 823
rect 523 819 524 823
rect 518 818 524 819
rect 614 823 620 824
rect 614 819 615 823
rect 619 819 620 823
rect 614 818 620 819
rect 718 823 724 824
rect 718 819 719 823
rect 723 819 724 823
rect 718 818 724 819
rect 830 823 836 824
rect 830 819 831 823
rect 835 819 836 823
rect 830 818 836 819
rect 950 823 956 824
rect 950 819 951 823
rect 955 819 956 823
rect 950 818 956 819
rect 1070 823 1076 824
rect 1070 819 1071 823
rect 1075 819 1076 823
rect 1070 818 1076 819
rect 1190 823 1196 824
rect 1190 819 1191 823
rect 1195 819 1196 823
rect 1190 818 1196 819
rect 1310 823 1316 824
rect 1310 819 1311 823
rect 1315 819 1316 823
rect 1310 818 1316 819
rect 1430 823 1436 824
rect 1430 819 1431 823
rect 1435 819 1436 823
rect 1430 818 1436 819
rect 1558 823 1564 824
rect 1558 819 1559 823
rect 1563 819 1564 823
rect 1766 820 1767 824
rect 1771 820 1772 824
rect 1902 823 1908 824
rect 1766 819 1772 820
rect 1806 819 1812 820
rect 1558 818 1564 819
rect 1022 815 1028 816
rect 686 811 692 812
rect 593 808 610 810
rect 110 807 116 808
rect 110 803 111 807
rect 115 803 116 807
rect 110 802 116 803
rect 518 804 524 805
rect 518 800 519 804
rect 523 800 524 804
rect 518 799 524 800
rect 608 794 610 808
rect 686 807 687 811
rect 691 807 692 811
rect 686 806 692 807
rect 790 811 796 812
rect 790 807 791 811
rect 795 807 796 811
rect 790 806 796 807
rect 902 811 908 812
rect 902 807 903 811
rect 907 807 908 811
rect 1022 811 1023 815
rect 1027 811 1028 815
rect 1630 815 1636 816
rect 1022 810 1028 811
rect 1142 811 1148 812
rect 902 806 908 807
rect 1142 807 1143 811
rect 1147 807 1148 811
rect 1142 806 1148 807
rect 1262 811 1268 812
rect 1262 807 1263 811
rect 1267 807 1268 811
rect 1262 806 1268 807
rect 1382 811 1388 812
rect 1382 807 1383 811
rect 1387 807 1388 811
rect 1382 806 1388 807
rect 1502 811 1508 812
rect 1502 807 1503 811
rect 1507 807 1508 811
rect 1630 811 1631 815
rect 1635 811 1636 815
rect 1806 815 1807 819
rect 1811 815 1812 819
rect 1902 819 1903 823
rect 1907 819 1908 823
rect 1902 818 1908 819
rect 2030 823 2036 824
rect 2030 819 2031 823
rect 2035 819 2036 823
rect 2038 823 2039 827
rect 2043 826 2044 827
rect 2286 827 2292 828
rect 2043 824 2129 826
rect 2043 823 2044 824
rect 2038 822 2044 823
rect 2278 823 2284 824
rect 2030 818 2036 819
rect 2278 819 2279 823
rect 2283 819 2284 823
rect 2286 823 2287 827
rect 2291 826 2292 827
rect 3138 827 3144 828
rect 2291 824 2369 826
rect 2291 823 2292 824
rect 2286 822 2292 823
rect 2534 823 2540 824
rect 2278 818 2284 819
rect 2534 819 2535 823
rect 2539 819 2540 823
rect 2534 818 2540 819
rect 2686 823 2692 824
rect 2686 819 2687 823
rect 2691 819 2692 823
rect 2686 818 2692 819
rect 2862 823 2868 824
rect 2862 819 2863 823
rect 2867 819 2868 823
rect 2862 818 2868 819
rect 3054 823 3060 824
rect 3054 819 3055 823
rect 3059 819 3060 823
rect 3138 823 3139 827
rect 3143 826 3144 827
rect 3438 827 3444 828
rect 3143 824 3225 826
rect 3143 823 3144 824
rect 3138 822 3144 823
rect 3438 823 3439 827
rect 3443 823 3444 827
rect 3438 822 3444 823
rect 3054 818 3060 819
rect 3462 819 3468 820
rect 1806 814 1812 815
rect 1830 816 1836 817
rect 1830 812 1831 816
rect 1835 812 1836 816
rect 1830 811 1836 812
rect 1958 816 1964 817
rect 1958 812 1959 816
rect 1963 812 1964 816
rect 1958 811 1964 812
rect 2086 816 2092 817
rect 2086 812 2087 816
rect 2091 812 2092 816
rect 2086 811 2092 812
rect 2206 816 2212 817
rect 2206 812 2207 816
rect 2211 812 2212 816
rect 2206 811 2212 812
rect 2326 816 2332 817
rect 2326 812 2327 816
rect 2331 812 2332 816
rect 2326 811 2332 812
rect 2462 816 2468 817
rect 2462 812 2463 816
rect 2467 812 2468 816
rect 2462 811 2468 812
rect 2614 816 2620 817
rect 2614 812 2615 816
rect 2619 812 2620 816
rect 2614 811 2620 812
rect 2790 816 2796 817
rect 2790 812 2791 816
rect 2795 812 2796 816
rect 2790 811 2796 812
rect 2982 816 2988 817
rect 2982 812 2983 816
rect 2987 812 2988 816
rect 2982 811 2988 812
rect 3182 816 3188 817
rect 3182 812 3183 816
rect 3187 812 3188 816
rect 3182 811 3188 812
rect 3366 816 3372 817
rect 3366 812 3367 816
rect 3371 812 3372 816
rect 3462 815 3463 819
rect 3467 815 3468 819
rect 3462 814 3468 815
rect 3366 811 3372 812
rect 1630 810 1636 811
rect 1502 806 1508 807
rect 1766 807 1772 808
rect 614 804 620 805
rect 614 800 615 804
rect 619 800 620 804
rect 614 799 620 800
rect 718 804 724 805
rect 718 800 719 804
rect 723 800 724 804
rect 718 799 724 800
rect 830 804 836 805
rect 830 800 831 804
rect 835 800 836 804
rect 830 799 836 800
rect 950 804 956 805
rect 950 800 951 804
rect 955 800 956 804
rect 950 799 956 800
rect 1070 804 1076 805
rect 1070 800 1071 804
rect 1075 800 1076 804
rect 1070 799 1076 800
rect 1190 804 1196 805
rect 1190 800 1191 804
rect 1195 800 1196 804
rect 1190 799 1196 800
rect 1310 804 1316 805
rect 1310 800 1311 804
rect 1315 800 1316 804
rect 1310 799 1316 800
rect 1430 804 1436 805
rect 1430 800 1431 804
rect 1435 800 1436 804
rect 1430 799 1436 800
rect 1558 804 1564 805
rect 1558 800 1559 804
rect 1563 800 1564 804
rect 1766 803 1767 807
rect 1771 803 1772 807
rect 2286 807 2292 808
rect 2286 806 2287 807
rect 1766 802 1772 803
rect 2140 804 2287 806
rect 2140 802 2142 804
rect 2286 803 2287 804
rect 2291 803 2292 807
rect 2286 802 2292 803
rect 2139 801 2145 802
rect 1558 799 1564 800
rect 1883 799 1889 800
rect 1883 795 1884 799
rect 1888 798 1889 799
rect 1894 799 1900 800
rect 1894 798 1895 799
rect 1888 796 1895 798
rect 1888 795 1889 796
rect 1883 794 1889 795
rect 1894 795 1895 796
rect 1899 795 1900 799
rect 1894 794 1900 795
rect 1902 799 1908 800
rect 1902 795 1903 799
rect 1907 798 1908 799
rect 2011 799 2017 800
rect 2011 798 2012 799
rect 1907 796 2012 798
rect 1907 795 1908 796
rect 1902 794 1908 795
rect 2011 795 2012 796
rect 2016 795 2017 799
rect 2139 797 2140 801
rect 2144 797 2145 801
rect 2139 796 2145 797
rect 2222 799 2228 800
rect 2011 794 2017 795
rect 2222 795 2223 799
rect 2227 798 2228 799
rect 2259 799 2265 800
rect 2259 798 2260 799
rect 2227 796 2260 798
rect 2227 795 2228 796
rect 2222 794 2228 795
rect 2259 795 2260 796
rect 2264 795 2265 799
rect 2259 794 2265 795
rect 2278 799 2284 800
rect 2278 795 2279 799
rect 2283 798 2284 799
rect 2379 799 2385 800
rect 2379 798 2380 799
rect 2283 796 2380 798
rect 2283 795 2284 796
rect 2278 794 2284 795
rect 2379 795 2380 796
rect 2384 795 2385 799
rect 2379 794 2385 795
rect 2398 799 2404 800
rect 2398 795 2399 799
rect 2403 798 2404 799
rect 2515 799 2521 800
rect 2515 798 2516 799
rect 2403 796 2516 798
rect 2403 795 2404 796
rect 2398 794 2404 795
rect 2515 795 2516 796
rect 2520 795 2521 799
rect 2515 794 2521 795
rect 2534 799 2540 800
rect 2534 795 2535 799
rect 2539 798 2540 799
rect 2667 799 2673 800
rect 2667 798 2668 799
rect 2539 796 2668 798
rect 2539 795 2540 796
rect 2534 794 2540 795
rect 2667 795 2668 796
rect 2672 795 2673 799
rect 2667 794 2673 795
rect 2686 799 2692 800
rect 2686 795 2687 799
rect 2691 798 2692 799
rect 2843 799 2849 800
rect 2843 798 2844 799
rect 2691 796 2844 798
rect 2691 795 2692 796
rect 2686 794 2692 795
rect 2843 795 2844 796
rect 2848 795 2849 799
rect 2843 794 2849 795
rect 2862 799 2868 800
rect 2862 795 2863 799
rect 2867 798 2868 799
rect 3035 799 3041 800
rect 3035 798 3036 799
rect 2867 796 3036 798
rect 2867 795 2868 796
rect 2862 794 2868 795
rect 3035 795 3036 796
rect 3040 795 3041 799
rect 3035 794 3041 795
rect 3054 799 3060 800
rect 3054 795 3055 799
rect 3059 798 3060 799
rect 3235 799 3241 800
rect 3235 798 3236 799
rect 3059 796 3236 798
rect 3059 795 3060 796
rect 3054 794 3060 795
rect 3235 795 3236 796
rect 3240 795 3241 799
rect 3235 794 3241 795
rect 3419 799 3425 800
rect 3419 795 3420 799
rect 3424 798 3425 799
rect 3430 799 3436 800
rect 3430 798 3431 799
rect 3424 796 3431 798
rect 3424 795 3425 796
rect 3419 794 3425 795
rect 3430 795 3431 796
rect 3435 795 3436 799
rect 3430 794 3436 795
rect 608 792 670 794
rect 668 790 670 792
rect 3138 791 3144 792
rect 3138 790 3139 791
rect 667 789 673 790
rect 571 787 577 788
rect 571 783 572 787
rect 576 786 577 787
rect 576 784 630 786
rect 667 785 668 789
rect 672 785 673 789
rect 2612 788 3139 790
rect 667 784 673 785
rect 686 787 692 788
rect 576 783 577 784
rect 571 782 577 783
rect 628 778 630 784
rect 686 783 687 787
rect 691 786 692 787
rect 771 787 777 788
rect 771 786 772 787
rect 691 784 772 786
rect 691 783 692 784
rect 686 782 692 783
rect 771 783 772 784
rect 776 783 777 787
rect 771 782 777 783
rect 790 787 796 788
rect 790 783 791 787
rect 795 786 796 787
rect 883 787 889 788
rect 883 786 884 787
rect 795 784 884 786
rect 795 783 796 784
rect 790 782 796 783
rect 883 783 884 784
rect 888 783 889 787
rect 883 782 889 783
rect 902 787 908 788
rect 902 783 903 787
rect 907 786 908 787
rect 1003 787 1009 788
rect 1003 786 1004 787
rect 907 784 1004 786
rect 907 783 908 784
rect 902 782 908 783
rect 1003 783 1004 784
rect 1008 783 1009 787
rect 1003 782 1009 783
rect 1123 787 1129 788
rect 1123 783 1124 787
rect 1128 786 1129 787
rect 1198 787 1204 788
rect 1198 786 1199 787
rect 1128 784 1199 786
rect 1128 783 1129 784
rect 1123 782 1129 783
rect 1198 783 1199 784
rect 1203 783 1204 787
rect 1198 782 1204 783
rect 1230 787 1236 788
rect 1230 783 1231 787
rect 1235 786 1236 787
rect 1243 787 1249 788
rect 1243 786 1244 787
rect 1235 784 1244 786
rect 1235 783 1236 784
rect 1230 782 1236 783
rect 1243 783 1244 784
rect 1248 783 1249 787
rect 1243 782 1249 783
rect 1262 787 1268 788
rect 1262 783 1263 787
rect 1267 786 1268 787
rect 1363 787 1369 788
rect 1363 786 1364 787
rect 1267 784 1364 786
rect 1267 783 1268 784
rect 1262 782 1268 783
rect 1363 783 1364 784
rect 1368 783 1369 787
rect 1363 782 1369 783
rect 1382 787 1388 788
rect 1382 783 1383 787
rect 1387 786 1388 787
rect 1483 787 1489 788
rect 1483 786 1484 787
rect 1387 784 1484 786
rect 1387 783 1388 784
rect 1382 782 1388 783
rect 1483 783 1484 784
rect 1488 783 1489 787
rect 1483 782 1489 783
rect 1502 787 1508 788
rect 1502 783 1503 787
rect 1507 786 1508 787
rect 1611 787 1617 788
rect 1611 786 1612 787
rect 1507 784 1612 786
rect 1507 783 1508 784
rect 1502 782 1508 783
rect 1611 783 1612 784
rect 1616 783 1617 787
rect 2612 786 2614 788
rect 3138 787 3139 788
rect 3143 787 3144 791
rect 3138 786 3144 787
rect 2611 785 2617 786
rect 1611 782 1617 783
rect 1931 783 1937 784
rect 758 779 764 780
rect 758 778 759 779
rect 628 776 759 778
rect 758 775 759 776
rect 763 775 764 779
rect 1931 779 1932 783
rect 1936 782 1937 783
rect 1959 783 1965 784
rect 1959 782 1960 783
rect 1936 780 1960 782
rect 1936 779 1937 780
rect 1931 778 1937 779
rect 1959 779 1960 780
rect 1964 779 1965 783
rect 1959 778 1965 779
rect 2030 783 2036 784
rect 2030 779 2031 783
rect 2035 782 2036 783
rect 2067 783 2073 784
rect 2067 782 2068 783
rect 2035 780 2068 782
rect 2035 779 2036 780
rect 2030 778 2036 779
rect 2067 779 2068 780
rect 2072 779 2073 783
rect 2067 778 2073 779
rect 2203 783 2209 784
rect 2203 779 2204 783
rect 2208 782 2209 783
rect 2230 783 2236 784
rect 2230 782 2231 783
rect 2208 780 2231 782
rect 2208 779 2209 780
rect 2203 778 2209 779
rect 2230 779 2231 780
rect 2235 779 2236 783
rect 2230 778 2236 779
rect 2339 783 2345 784
rect 2339 779 2340 783
rect 2344 782 2345 783
rect 2366 783 2372 784
rect 2366 782 2367 783
rect 2344 780 2367 782
rect 2344 779 2345 780
rect 2339 778 2345 779
rect 2366 779 2367 780
rect 2371 779 2372 783
rect 2366 778 2372 779
rect 2475 783 2481 784
rect 2475 779 2476 783
rect 2480 782 2481 783
rect 2486 783 2492 784
rect 2486 782 2487 783
rect 2480 780 2487 782
rect 2480 779 2481 780
rect 2475 778 2481 779
rect 2486 779 2487 780
rect 2491 779 2492 783
rect 2611 781 2612 785
rect 2616 781 2617 785
rect 2611 780 2617 781
rect 2630 783 2636 784
rect 2486 778 2492 779
rect 2630 779 2631 783
rect 2635 782 2636 783
rect 2763 783 2769 784
rect 2763 782 2764 783
rect 2635 780 2764 782
rect 2635 779 2636 780
rect 2630 778 2636 779
rect 2763 779 2764 780
rect 2768 779 2769 783
rect 2763 778 2769 779
rect 2782 783 2788 784
rect 2782 779 2783 783
rect 2787 782 2788 783
rect 2923 783 2929 784
rect 2923 782 2924 783
rect 2787 780 2924 782
rect 2787 779 2788 780
rect 2782 778 2788 779
rect 2923 779 2924 780
rect 2928 779 2929 783
rect 2923 778 2929 779
rect 2942 783 2948 784
rect 2942 779 2943 783
rect 2947 782 2948 783
rect 3091 783 3097 784
rect 3091 782 3092 783
rect 2947 780 3092 782
rect 2947 779 2948 780
rect 2942 778 2948 779
rect 3091 779 3092 780
rect 3096 779 3097 783
rect 3091 778 3097 779
rect 3110 783 3116 784
rect 3110 779 3111 783
rect 3115 782 3116 783
rect 3267 783 3273 784
rect 3267 782 3268 783
rect 3115 780 3268 782
rect 3115 779 3116 780
rect 3110 778 3116 779
rect 3267 779 3268 780
rect 3272 779 3273 783
rect 3267 778 3273 779
rect 3419 783 3425 784
rect 3419 779 3420 783
rect 3424 782 3425 783
rect 3438 783 3444 784
rect 3438 782 3439 783
rect 3424 780 3439 782
rect 3424 779 3425 780
rect 3419 778 3425 779
rect 3438 779 3439 780
rect 3443 779 3444 783
rect 3438 778 3444 779
rect 758 774 764 775
rect 435 771 441 772
rect 435 767 436 771
rect 440 770 441 771
rect 454 771 460 772
rect 440 768 450 770
rect 440 767 441 768
rect 435 766 441 767
rect 448 762 450 768
rect 454 767 455 771
rect 459 770 460 771
rect 523 771 529 772
rect 523 770 524 771
rect 459 768 524 770
rect 459 767 460 768
rect 454 766 460 767
rect 523 767 524 768
rect 528 767 529 771
rect 523 766 529 767
rect 542 771 548 772
rect 542 767 543 771
rect 547 770 548 771
rect 627 771 633 772
rect 627 770 628 771
rect 547 768 628 770
rect 547 767 548 768
rect 542 766 548 767
rect 627 767 628 768
rect 632 767 633 771
rect 627 766 633 767
rect 646 771 652 772
rect 646 767 647 771
rect 651 770 652 771
rect 731 771 737 772
rect 731 770 732 771
rect 651 768 732 770
rect 651 767 652 768
rect 646 766 652 767
rect 731 767 732 768
rect 736 767 737 771
rect 731 766 737 767
rect 750 771 756 772
rect 750 767 751 771
rect 755 770 756 771
rect 843 771 849 772
rect 843 770 844 771
rect 755 768 844 770
rect 755 767 756 768
rect 750 766 756 767
rect 843 767 844 768
rect 848 767 849 771
rect 843 766 849 767
rect 963 771 969 772
rect 963 767 964 771
rect 968 770 969 771
rect 990 771 996 772
rect 990 770 991 771
rect 968 768 991 770
rect 968 767 969 768
rect 963 766 969 767
rect 990 767 991 768
rect 995 767 996 771
rect 990 766 996 767
rect 1083 771 1089 772
rect 1083 767 1084 771
rect 1088 770 1089 771
rect 1142 771 1148 772
rect 1142 770 1143 771
rect 1088 768 1143 770
rect 1088 767 1089 768
rect 1083 766 1089 767
rect 1142 767 1143 768
rect 1147 767 1148 771
rect 1142 766 1148 767
rect 1211 771 1217 772
rect 1211 767 1212 771
rect 1216 770 1217 771
rect 1238 771 1244 772
rect 1238 770 1239 771
rect 1216 768 1239 770
rect 1216 767 1217 768
rect 1211 766 1217 767
rect 1238 767 1239 768
rect 1243 767 1244 771
rect 1238 766 1244 767
rect 1339 771 1345 772
rect 1339 767 1340 771
rect 1344 770 1345 771
rect 1366 771 1372 772
rect 1366 770 1367 771
rect 1344 768 1367 770
rect 1344 767 1345 768
rect 1339 766 1345 767
rect 1366 767 1367 768
rect 1371 767 1372 771
rect 1366 766 1372 767
rect 1467 771 1473 772
rect 1467 767 1468 771
rect 1472 770 1473 771
rect 1503 771 1509 772
rect 1503 770 1504 771
rect 1472 768 1504 770
rect 1472 767 1473 768
rect 1467 766 1473 767
rect 1503 767 1504 768
rect 1508 767 1509 771
rect 1503 766 1509 767
rect 1878 768 1884 769
rect 1806 765 1812 766
rect 654 763 660 764
rect 654 762 655 763
rect 448 760 655 762
rect 654 759 655 760
rect 659 759 660 763
rect 1806 761 1807 765
rect 1811 761 1812 765
rect 1878 764 1879 768
rect 1883 764 1884 768
rect 1878 763 1884 764
rect 2014 768 2020 769
rect 2014 764 2015 768
rect 2019 764 2020 768
rect 2014 763 2020 764
rect 2150 768 2156 769
rect 2150 764 2151 768
rect 2155 764 2156 768
rect 2150 763 2156 764
rect 2286 768 2292 769
rect 2286 764 2287 768
rect 2291 764 2292 768
rect 2286 763 2292 764
rect 2422 768 2428 769
rect 2422 764 2423 768
rect 2427 764 2428 768
rect 2422 763 2428 764
rect 2558 768 2564 769
rect 2558 764 2559 768
rect 2563 764 2564 768
rect 2558 763 2564 764
rect 2710 768 2716 769
rect 2710 764 2711 768
rect 2715 764 2716 768
rect 2710 763 2716 764
rect 2870 768 2876 769
rect 2870 764 2871 768
rect 2875 764 2876 768
rect 2870 763 2876 764
rect 3038 768 3044 769
rect 3038 764 3039 768
rect 3043 764 3044 768
rect 3038 763 3044 764
rect 3214 768 3220 769
rect 3214 764 3215 768
rect 3219 764 3220 768
rect 3214 763 3220 764
rect 3366 768 3372 769
rect 3366 764 3367 768
rect 3371 764 3372 768
rect 3366 763 3372 764
rect 3462 765 3468 766
rect 1806 760 1812 761
rect 3462 761 3463 765
rect 3467 761 3468 765
rect 3462 760 3468 761
rect 654 758 660 759
rect 1959 759 1965 760
rect 382 756 388 757
rect 110 753 116 754
rect 110 749 111 753
rect 115 749 116 753
rect 382 752 383 756
rect 387 752 388 756
rect 382 751 388 752
rect 470 756 476 757
rect 470 752 471 756
rect 475 752 476 756
rect 470 751 476 752
rect 574 756 580 757
rect 574 752 575 756
rect 579 752 580 756
rect 574 751 580 752
rect 678 756 684 757
rect 678 752 679 756
rect 683 752 684 756
rect 678 751 684 752
rect 790 756 796 757
rect 790 752 791 756
rect 795 752 796 756
rect 790 751 796 752
rect 910 756 916 757
rect 910 752 911 756
rect 915 752 916 756
rect 910 751 916 752
rect 1030 756 1036 757
rect 1030 752 1031 756
rect 1035 752 1036 756
rect 1030 751 1036 752
rect 1158 756 1164 757
rect 1158 752 1159 756
rect 1163 752 1164 756
rect 1158 751 1164 752
rect 1286 756 1292 757
rect 1286 752 1287 756
rect 1291 752 1292 756
rect 1286 751 1292 752
rect 1414 756 1420 757
rect 1414 752 1415 756
rect 1419 752 1420 756
rect 1959 755 1960 759
rect 1964 758 1965 759
rect 2222 759 2228 760
rect 1964 756 2057 758
rect 1964 755 1965 756
rect 1959 754 1965 755
rect 2222 755 2223 759
rect 2227 755 2228 759
rect 2222 754 2228 755
rect 2230 759 2236 760
rect 2230 755 2231 759
rect 2235 758 2236 759
rect 2366 759 2372 760
rect 2235 756 2329 758
rect 2235 755 2236 756
rect 2230 754 2236 755
rect 2366 755 2367 759
rect 2371 758 2372 759
rect 2630 759 2636 760
rect 2371 756 2465 758
rect 2371 755 2372 756
rect 2366 754 2372 755
rect 2630 755 2631 759
rect 2635 755 2636 759
rect 2630 754 2636 755
rect 2782 759 2788 760
rect 2782 755 2783 759
rect 2787 755 2788 759
rect 2782 754 2788 755
rect 2942 759 2948 760
rect 2942 755 2943 759
rect 2947 755 2948 759
rect 2942 754 2948 755
rect 3110 759 3116 760
rect 3110 755 3111 759
rect 3115 755 3116 759
rect 3110 754 3116 755
rect 3278 759 3284 760
rect 3278 755 3279 759
rect 3283 755 3284 759
rect 3278 754 3284 755
rect 3430 759 3436 760
rect 3430 755 3431 759
rect 3435 755 3436 759
rect 3430 754 3436 755
rect 1414 751 1420 752
rect 1766 753 1772 754
rect 110 748 116 749
rect 1766 749 1767 753
rect 1771 749 1772 753
rect 1951 751 1957 752
rect 1878 749 1884 750
rect 1766 748 1772 749
rect 1806 748 1812 749
rect 454 747 460 748
rect 454 743 455 747
rect 459 743 460 747
rect 454 742 460 743
rect 542 747 548 748
rect 542 743 543 747
rect 547 743 548 747
rect 542 742 548 743
rect 646 747 652 748
rect 646 743 647 747
rect 651 743 652 747
rect 646 742 652 743
rect 750 747 756 748
rect 750 743 751 747
rect 755 743 756 747
rect 750 742 756 743
rect 758 747 764 748
rect 758 743 759 747
rect 763 746 764 747
rect 990 747 996 748
rect 763 744 833 746
rect 763 743 764 744
rect 758 742 764 743
rect 990 743 991 747
rect 995 746 996 747
rect 1230 747 1236 748
rect 995 744 1073 746
rect 995 743 996 744
rect 990 742 996 743
rect 1230 743 1231 747
rect 1235 743 1236 747
rect 1230 742 1236 743
rect 1238 747 1244 748
rect 1238 743 1239 747
rect 1243 746 1244 747
rect 1366 747 1372 748
rect 1243 744 1329 746
rect 1243 743 1244 744
rect 1238 742 1244 743
rect 1366 743 1367 747
rect 1371 746 1372 747
rect 1371 744 1457 746
rect 1806 744 1807 748
rect 1811 744 1812 748
rect 1878 745 1879 749
rect 1883 745 1884 749
rect 1951 747 1952 751
rect 1956 750 1957 751
rect 1962 751 1968 752
rect 1962 750 1963 751
rect 1956 748 1963 750
rect 1956 747 1957 748
rect 1951 746 1957 747
rect 1962 747 1963 748
rect 1967 747 1968 751
rect 1962 746 1968 747
rect 2014 749 2020 750
rect 1878 744 1884 745
rect 2014 745 2015 749
rect 2019 745 2020 749
rect 2014 744 2020 745
rect 2150 749 2156 750
rect 2150 745 2151 749
rect 2155 745 2156 749
rect 2150 744 2156 745
rect 2286 749 2292 750
rect 2286 745 2287 749
rect 2291 745 2292 749
rect 2286 744 2292 745
rect 2422 749 2428 750
rect 2422 745 2423 749
rect 2427 745 2428 749
rect 2422 744 2428 745
rect 2558 749 2564 750
rect 2558 745 2559 749
rect 2563 745 2564 749
rect 2558 744 2564 745
rect 2710 749 2716 750
rect 2710 745 2711 749
rect 2715 745 2716 749
rect 2710 744 2716 745
rect 2870 749 2876 750
rect 2870 745 2871 749
rect 2875 745 2876 749
rect 2870 744 2876 745
rect 3038 749 3044 750
rect 3038 745 3039 749
rect 3043 745 3044 749
rect 3038 744 3044 745
rect 3214 749 3220 750
rect 3214 745 3215 749
rect 3219 745 3220 749
rect 3214 744 3220 745
rect 3366 749 3372 750
rect 3366 745 3367 749
rect 3371 745 3372 749
rect 3366 744 3372 745
rect 3462 748 3468 749
rect 3462 744 3463 748
rect 3467 744 3468 748
rect 1371 743 1372 744
rect 1806 743 1812 744
rect 3462 743 3468 744
rect 1366 742 1372 743
rect 983 739 989 740
rect 382 737 388 738
rect 110 736 116 737
rect 110 732 111 736
rect 115 732 116 736
rect 382 733 383 737
rect 387 733 388 737
rect 382 732 388 733
rect 470 737 476 738
rect 470 733 471 737
rect 475 733 476 737
rect 470 732 476 733
rect 574 737 580 738
rect 574 733 575 737
rect 579 733 580 737
rect 574 732 580 733
rect 678 737 684 738
rect 678 733 679 737
rect 683 733 684 737
rect 678 732 684 733
rect 790 737 796 738
rect 790 733 791 737
rect 795 733 796 737
rect 790 732 796 733
rect 910 737 916 738
rect 910 733 911 737
rect 915 733 916 737
rect 983 735 984 739
rect 988 738 989 739
rect 994 739 1000 740
rect 994 738 995 739
rect 988 736 995 738
rect 988 735 989 736
rect 983 734 989 735
rect 994 735 995 736
rect 999 735 1000 739
rect 994 734 1000 735
rect 1030 737 1036 738
rect 910 732 916 733
rect 1030 733 1031 737
rect 1035 733 1036 737
rect 1030 732 1036 733
rect 1158 737 1164 738
rect 1158 733 1159 737
rect 1163 733 1164 737
rect 1158 732 1164 733
rect 1286 737 1292 738
rect 1286 733 1287 737
rect 1291 733 1292 737
rect 1286 732 1292 733
rect 1414 737 1420 738
rect 1414 733 1415 737
rect 1419 733 1420 737
rect 1414 732 1420 733
rect 1766 736 1772 737
rect 1766 732 1767 736
rect 1771 732 1772 736
rect 110 731 116 732
rect 1766 731 1772 732
rect 1806 700 1812 701
rect 3462 700 3468 701
rect 1806 696 1807 700
rect 1811 696 1812 700
rect 1806 695 1812 696
rect 1830 699 1836 700
rect 1830 695 1831 699
rect 1835 695 1836 699
rect 1830 694 1836 695
rect 1950 699 1956 700
rect 1950 695 1951 699
rect 1955 695 1956 699
rect 1950 694 1956 695
rect 2102 699 2108 700
rect 2102 695 2103 699
rect 2107 695 2108 699
rect 2102 694 2108 695
rect 2262 699 2268 700
rect 2262 695 2263 699
rect 2267 695 2268 699
rect 2262 694 2268 695
rect 2414 699 2420 700
rect 2414 695 2415 699
rect 2419 695 2420 699
rect 2414 694 2420 695
rect 2566 699 2572 700
rect 2566 695 2567 699
rect 2571 695 2572 699
rect 2566 694 2572 695
rect 2718 699 2724 700
rect 2718 695 2719 699
rect 2723 695 2724 699
rect 2718 694 2724 695
rect 2878 699 2884 700
rect 2878 695 2879 699
rect 2883 695 2884 699
rect 2878 694 2884 695
rect 3038 699 3044 700
rect 3038 695 3039 699
rect 3043 695 3044 699
rect 3038 694 3044 695
rect 3198 699 3204 700
rect 3198 695 3199 699
rect 3203 695 3204 699
rect 3462 696 3463 700
rect 3467 696 3468 700
rect 3462 695 3468 696
rect 3198 694 3204 695
rect 1750 691 1756 692
rect 1750 687 1751 691
rect 1755 690 1756 691
rect 1910 691 1916 692
rect 1755 688 1873 690
rect 1755 687 1756 688
rect 1750 686 1756 687
rect 1910 687 1911 691
rect 1915 690 1916 691
rect 2486 691 2492 692
rect 1915 688 1993 690
rect 1915 687 1916 688
rect 1910 686 1916 687
rect 2174 687 2180 688
rect 110 684 116 685
rect 1766 684 1772 685
rect 110 680 111 684
rect 115 680 116 684
rect 110 679 116 680
rect 246 683 252 684
rect 246 679 247 683
rect 251 679 252 683
rect 246 678 252 679
rect 342 683 348 684
rect 342 679 343 683
rect 347 679 348 683
rect 342 678 348 679
rect 454 683 460 684
rect 454 679 455 683
rect 459 679 460 683
rect 454 678 460 679
rect 566 683 572 684
rect 566 679 567 683
rect 571 679 572 683
rect 566 678 572 679
rect 694 683 700 684
rect 694 679 695 683
rect 699 679 700 683
rect 694 678 700 679
rect 830 683 836 684
rect 830 679 831 683
rect 835 679 836 683
rect 830 678 836 679
rect 982 683 988 684
rect 982 679 983 683
rect 987 679 988 683
rect 982 678 988 679
rect 1150 683 1156 684
rect 1150 679 1151 683
rect 1155 679 1156 683
rect 1150 678 1156 679
rect 1326 683 1332 684
rect 1326 679 1327 683
rect 1331 679 1332 683
rect 1326 678 1332 679
rect 1510 683 1516 684
rect 1510 679 1511 683
rect 1515 679 1516 683
rect 1510 678 1516 679
rect 1670 683 1676 684
rect 1670 679 1671 683
rect 1675 679 1676 683
rect 1766 680 1767 684
rect 1771 680 1772 684
rect 1766 679 1772 680
rect 1806 683 1812 684
rect 1806 679 1807 683
rect 1811 679 1812 683
rect 2174 683 2175 687
rect 2179 683 2180 687
rect 2174 682 2180 683
rect 2334 687 2340 688
rect 2334 683 2335 687
rect 2339 683 2340 687
rect 2486 687 2487 691
rect 2491 687 2492 691
rect 2486 686 2492 687
rect 2646 691 2652 692
rect 2646 687 2647 691
rect 2651 690 2652 691
rect 2798 691 2804 692
rect 2651 688 2761 690
rect 2651 687 2652 688
rect 2646 686 2652 687
rect 2798 687 2799 691
rect 2803 690 2804 691
rect 3138 691 3144 692
rect 2803 688 2921 690
rect 2803 687 2804 688
rect 2798 686 2804 687
rect 3110 687 3116 688
rect 2632 684 2641 686
rect 2334 682 2340 683
rect 2630 683 2636 684
rect 1670 678 1676 679
rect 1806 678 1812 679
rect 1830 680 1836 681
rect 1830 676 1831 680
rect 1835 676 1836 680
rect 654 675 660 676
rect 318 671 324 672
rect 110 667 116 668
rect 110 663 111 667
rect 115 663 116 667
rect 318 667 319 671
rect 323 667 324 671
rect 318 666 324 667
rect 414 671 420 672
rect 414 667 415 671
rect 419 667 420 671
rect 414 666 420 667
rect 526 671 532 672
rect 526 667 527 671
rect 531 667 532 671
rect 526 666 532 667
rect 638 671 644 672
rect 638 667 639 671
rect 643 667 644 671
rect 654 671 655 675
rect 659 674 660 675
rect 822 675 828 676
rect 659 672 737 674
rect 659 671 660 672
rect 654 670 660 671
rect 822 671 823 675
rect 827 674 828 675
rect 910 675 916 676
rect 827 672 873 674
rect 827 671 828 672
rect 822 670 828 671
rect 910 671 911 675
rect 915 674 916 675
rect 1503 675 1509 676
rect 1830 675 1836 676
rect 1950 680 1956 681
rect 1950 676 1951 680
rect 1955 676 1956 680
rect 1950 675 1956 676
rect 2102 680 2108 681
rect 2102 676 2103 680
rect 2107 676 2108 680
rect 2102 675 2108 676
rect 2262 680 2268 681
rect 2262 676 2263 680
rect 2267 676 2268 680
rect 2262 675 2268 676
rect 2414 680 2420 681
rect 2414 676 2415 680
rect 2419 676 2420 680
rect 2414 675 2420 676
rect 2566 680 2572 681
rect 2566 676 2567 680
rect 2571 676 2572 680
rect 2630 679 2631 683
rect 2635 679 2636 683
rect 3110 683 3111 687
rect 3115 683 3116 687
rect 3138 687 3139 691
rect 3143 690 3144 691
rect 3143 688 3241 690
rect 3143 687 3144 688
rect 3138 686 3144 687
rect 3110 682 3116 683
rect 3462 683 3468 684
rect 2630 678 2636 679
rect 2718 680 2724 681
rect 2566 675 2572 676
rect 2718 676 2719 680
rect 2723 676 2724 680
rect 2718 675 2724 676
rect 2878 680 2884 681
rect 2878 676 2879 680
rect 2883 676 2884 680
rect 2878 675 2884 676
rect 3038 680 3044 681
rect 3038 676 3039 680
rect 3043 676 3044 680
rect 3038 675 3044 676
rect 3198 680 3204 681
rect 3198 676 3199 680
rect 3203 676 3204 680
rect 3462 679 3463 683
rect 3467 679 3468 683
rect 3462 678 3468 679
rect 3198 675 3204 676
rect 915 672 1025 674
rect 915 671 916 672
rect 910 670 916 671
rect 1294 671 1300 672
rect 1294 670 1295 671
rect 1225 668 1295 670
rect 638 666 644 667
rect 1294 667 1295 668
rect 1299 667 1300 671
rect 1294 666 1300 667
rect 1398 671 1404 672
rect 1398 667 1399 671
rect 1403 667 1404 671
rect 1503 671 1504 675
rect 1508 674 1509 675
rect 1508 672 1553 674
rect 1508 671 1509 672
rect 1503 670 1509 671
rect 1742 671 1748 672
rect 1398 666 1404 667
rect 1742 667 1743 671
rect 1747 667 1748 671
rect 3138 671 3144 672
rect 3138 670 3139 671
rect 2932 668 3139 670
rect 1742 666 1748 667
rect 1766 667 1772 668
rect 110 662 116 663
rect 246 664 252 665
rect 246 660 247 664
rect 251 660 252 664
rect 246 659 252 660
rect 342 664 348 665
rect 342 660 343 664
rect 347 660 348 664
rect 342 659 348 660
rect 454 664 460 665
rect 454 660 455 664
rect 459 660 460 664
rect 454 659 460 660
rect 566 664 572 665
rect 566 660 567 664
rect 571 660 572 664
rect 566 659 572 660
rect 694 664 700 665
rect 694 660 695 664
rect 699 660 700 664
rect 694 659 700 660
rect 830 664 836 665
rect 830 660 831 664
rect 835 660 836 664
rect 830 659 836 660
rect 982 664 988 665
rect 982 660 983 664
rect 987 660 988 664
rect 982 659 988 660
rect 1150 664 1156 665
rect 1150 660 1151 664
rect 1155 660 1156 664
rect 1150 659 1156 660
rect 1326 664 1332 665
rect 1326 660 1327 664
rect 1331 660 1332 664
rect 1326 659 1332 660
rect 1510 664 1516 665
rect 1510 660 1511 664
rect 1515 660 1516 664
rect 1510 659 1516 660
rect 1670 664 1676 665
rect 1670 660 1671 664
rect 1675 660 1676 664
rect 1766 663 1767 667
rect 1771 663 1772 667
rect 2932 666 2934 668
rect 3138 667 3139 668
rect 3143 667 3144 671
rect 3138 666 3144 667
rect 2931 665 2937 666
rect 1766 662 1772 663
rect 1883 663 1889 664
rect 1670 659 1676 660
rect 1883 659 1884 663
rect 1888 662 1889 663
rect 1910 663 1916 664
rect 1910 662 1911 663
rect 1888 660 1911 662
rect 1888 659 1889 660
rect 1883 658 1889 659
rect 1910 659 1911 660
rect 1915 659 1916 663
rect 1910 658 1916 659
rect 1962 663 1968 664
rect 1962 659 1963 663
rect 1967 662 1968 663
rect 2003 663 2009 664
rect 2003 662 2004 663
rect 1967 660 2004 662
rect 1967 659 1968 660
rect 1962 658 1968 659
rect 2003 659 2004 660
rect 2008 659 2009 663
rect 2003 658 2009 659
rect 2155 663 2164 664
rect 2155 659 2156 663
rect 2163 659 2164 663
rect 2155 658 2164 659
rect 2174 663 2180 664
rect 2174 659 2175 663
rect 2179 662 2180 663
rect 2315 663 2321 664
rect 2315 662 2316 663
rect 2179 660 2316 662
rect 2179 659 2180 660
rect 2174 658 2180 659
rect 2315 659 2316 660
rect 2320 659 2321 663
rect 2315 658 2321 659
rect 2334 663 2340 664
rect 2334 659 2335 663
rect 2339 662 2340 663
rect 2467 663 2473 664
rect 2467 662 2468 663
rect 2339 660 2468 662
rect 2339 659 2340 660
rect 2334 658 2340 659
rect 2467 659 2468 660
rect 2472 659 2473 663
rect 2467 658 2473 659
rect 2619 663 2625 664
rect 2619 659 2620 663
rect 2624 662 2625 663
rect 2646 663 2652 664
rect 2646 662 2647 663
rect 2624 660 2647 662
rect 2624 659 2625 660
rect 2619 658 2625 659
rect 2646 659 2647 660
rect 2651 659 2652 663
rect 2646 658 2652 659
rect 2771 663 2777 664
rect 2771 659 2772 663
rect 2776 662 2777 663
rect 2798 663 2804 664
rect 2798 662 2799 663
rect 2776 660 2799 662
rect 2776 659 2777 660
rect 2771 658 2777 659
rect 2798 659 2799 660
rect 2803 659 2804 663
rect 2931 661 2932 665
rect 2936 661 2937 665
rect 2931 660 2937 661
rect 2950 663 2956 664
rect 2798 658 2804 659
rect 2950 659 2951 663
rect 2955 662 2956 663
rect 3091 663 3097 664
rect 3091 662 3092 663
rect 2955 660 3092 662
rect 2955 659 2956 660
rect 2950 658 2956 659
rect 3091 659 3092 660
rect 3096 659 3097 663
rect 3091 658 3097 659
rect 3251 663 3257 664
rect 3251 659 3252 663
rect 3256 662 3257 663
rect 3278 663 3284 664
rect 3278 662 3279 663
rect 3256 660 3279 662
rect 3256 659 3257 660
rect 3251 658 3257 659
rect 3278 659 3279 660
rect 3283 659 3284 663
rect 3278 658 3284 659
rect 1966 651 1972 652
rect 299 647 305 648
rect 299 643 300 647
rect 304 646 305 647
rect 318 647 324 648
rect 304 644 314 646
rect 304 643 305 644
rect 299 642 305 643
rect 312 638 314 644
rect 318 643 319 647
rect 323 646 324 647
rect 395 647 401 648
rect 395 646 396 647
rect 323 644 396 646
rect 323 643 324 644
rect 318 642 324 643
rect 395 643 396 644
rect 400 643 401 647
rect 395 642 401 643
rect 414 647 420 648
rect 414 643 415 647
rect 419 646 420 647
rect 507 647 513 648
rect 507 646 508 647
rect 419 644 508 646
rect 419 643 420 644
rect 414 642 420 643
rect 507 643 508 644
rect 512 643 513 647
rect 507 642 513 643
rect 526 647 532 648
rect 526 643 527 647
rect 531 646 532 647
rect 619 647 625 648
rect 619 646 620 647
rect 531 644 620 646
rect 531 643 532 644
rect 526 642 532 643
rect 619 643 620 644
rect 624 643 625 647
rect 619 642 625 643
rect 638 647 644 648
rect 638 643 639 647
rect 643 646 644 647
rect 747 647 753 648
rect 747 646 748 647
rect 643 644 748 646
rect 643 643 644 644
rect 638 642 644 643
rect 747 643 748 644
rect 752 643 753 647
rect 747 642 753 643
rect 883 647 889 648
rect 883 643 884 647
rect 888 646 889 647
rect 910 647 916 648
rect 910 646 911 647
rect 888 644 911 646
rect 888 643 889 644
rect 883 642 889 643
rect 910 643 911 644
rect 915 643 916 647
rect 910 642 916 643
rect 994 647 1000 648
rect 994 643 995 647
rect 999 646 1000 647
rect 1035 647 1041 648
rect 1035 646 1036 647
rect 999 644 1036 646
rect 999 643 1000 644
rect 994 642 1000 643
rect 1035 643 1036 644
rect 1040 643 1041 647
rect 1035 642 1041 643
rect 1203 647 1209 648
rect 1203 643 1204 647
rect 1208 646 1209 647
rect 1286 647 1292 648
rect 1286 646 1287 647
rect 1208 644 1287 646
rect 1208 643 1209 644
rect 1203 642 1209 643
rect 1286 643 1287 644
rect 1291 643 1292 647
rect 1286 642 1292 643
rect 1294 647 1300 648
rect 1294 643 1295 647
rect 1299 646 1300 647
rect 1379 647 1385 648
rect 1379 646 1380 647
rect 1299 644 1380 646
rect 1299 643 1300 644
rect 1294 642 1300 643
rect 1379 643 1380 644
rect 1384 643 1385 647
rect 1379 642 1385 643
rect 1398 647 1404 648
rect 1398 643 1399 647
rect 1403 646 1404 647
rect 1563 647 1569 648
rect 1563 646 1564 647
rect 1403 644 1564 646
rect 1403 643 1404 644
rect 1398 642 1404 643
rect 1563 643 1564 644
rect 1568 643 1569 647
rect 1563 642 1569 643
rect 1723 647 1729 648
rect 1723 643 1724 647
rect 1728 646 1729 647
rect 1750 647 1756 648
rect 1750 646 1751 647
rect 1728 644 1751 646
rect 1728 643 1729 644
rect 1723 642 1729 643
rect 1750 643 1751 644
rect 1755 643 1756 647
rect 1966 647 1967 651
rect 1971 650 1972 651
rect 2027 651 2033 652
rect 2027 650 2028 651
rect 1971 648 2028 650
rect 1971 647 1972 648
rect 1966 646 1972 647
rect 2027 647 2028 648
rect 2032 647 2033 651
rect 2027 646 2033 647
rect 2046 651 2052 652
rect 2046 647 2047 651
rect 2051 650 2052 651
rect 2291 651 2297 652
rect 2291 650 2292 651
rect 2051 648 2292 650
rect 2051 647 2052 648
rect 2046 646 2052 647
rect 2291 647 2292 648
rect 2296 647 2297 651
rect 2291 646 2297 647
rect 2531 651 2537 652
rect 2531 647 2532 651
rect 2536 647 2537 651
rect 2531 646 2537 647
rect 2550 651 2556 652
rect 2550 647 2551 651
rect 2555 650 2556 651
rect 2739 651 2745 652
rect 2739 650 2740 651
rect 2555 648 2740 650
rect 2555 647 2556 648
rect 2550 646 2556 647
rect 2739 647 2740 648
rect 2744 647 2745 651
rect 2739 646 2745 647
rect 2758 651 2764 652
rect 2758 647 2759 651
rect 2763 650 2764 651
rect 2931 651 2937 652
rect 2931 650 2932 651
rect 2763 648 2932 650
rect 2763 647 2764 648
rect 2758 646 2764 647
rect 2931 647 2932 648
rect 2936 647 2937 651
rect 2931 646 2937 647
rect 3107 651 3116 652
rect 3107 647 3108 651
rect 3115 647 3116 651
rect 3107 646 3116 647
rect 3126 651 3132 652
rect 3126 647 3127 651
rect 3131 650 3132 651
rect 3275 651 3281 652
rect 3275 650 3276 651
rect 3131 648 3276 650
rect 3131 647 3132 648
rect 3126 646 3132 647
rect 3275 647 3276 648
rect 3280 647 3281 651
rect 3275 646 3281 647
rect 3419 651 3425 652
rect 3419 647 3420 651
rect 3424 650 3425 651
rect 3430 651 3436 652
rect 3430 650 3431 651
rect 3424 648 3431 650
rect 3424 647 3425 648
rect 3419 646 3425 647
rect 3430 647 3431 648
rect 3435 647 3436 651
rect 3430 646 3436 647
rect 1750 642 1756 643
rect 2533 642 2535 646
rect 2838 643 2844 644
rect 2838 642 2839 643
rect 2533 640 2839 642
rect 567 639 573 640
rect 567 638 568 639
rect 312 636 568 638
rect 567 635 568 636
rect 572 635 573 639
rect 2838 639 2839 640
rect 2843 639 2844 643
rect 2838 638 2844 639
rect 567 634 573 635
rect 1974 636 1980 637
rect 1806 633 1812 634
rect 187 631 193 632
rect 187 627 188 631
rect 192 630 193 631
rect 198 631 204 632
rect 198 630 199 631
rect 192 628 199 630
rect 192 627 193 628
rect 187 626 193 627
rect 198 627 199 628
rect 203 627 204 631
rect 198 626 204 627
rect 206 631 212 632
rect 206 627 207 631
rect 211 630 212 631
rect 283 631 289 632
rect 283 630 284 631
rect 211 628 284 630
rect 211 627 212 628
rect 206 626 212 627
rect 283 627 284 628
rect 288 627 289 631
rect 283 626 289 627
rect 302 631 308 632
rect 302 627 303 631
rect 307 630 308 631
rect 411 631 417 632
rect 411 630 412 631
rect 307 628 412 630
rect 307 627 308 628
rect 302 626 308 627
rect 411 627 412 628
rect 416 627 417 631
rect 411 626 417 627
rect 430 631 436 632
rect 430 627 431 631
rect 435 630 436 631
rect 539 631 545 632
rect 539 630 540 631
rect 435 628 540 630
rect 435 627 436 628
rect 430 626 436 627
rect 539 627 540 628
rect 544 627 545 631
rect 539 626 545 627
rect 558 631 564 632
rect 558 627 559 631
rect 563 630 564 631
rect 675 631 681 632
rect 675 630 676 631
rect 563 628 676 630
rect 563 627 564 628
rect 558 626 564 627
rect 675 627 676 628
rect 680 627 681 631
rect 675 626 681 627
rect 819 631 828 632
rect 819 627 820 631
rect 827 627 828 631
rect 963 631 969 632
rect 963 630 964 631
rect 819 626 828 627
rect 864 628 964 630
rect 134 616 140 617
rect 110 613 116 614
rect 110 609 111 613
rect 115 609 116 613
rect 134 612 135 616
rect 139 612 140 616
rect 134 611 140 612
rect 230 616 236 617
rect 230 612 231 616
rect 235 612 236 616
rect 230 611 236 612
rect 358 616 364 617
rect 358 612 359 616
rect 363 612 364 616
rect 358 611 364 612
rect 486 616 492 617
rect 486 612 487 616
rect 491 612 492 616
rect 486 611 492 612
rect 622 616 628 617
rect 622 612 623 616
rect 627 612 628 616
rect 622 611 628 612
rect 766 616 772 617
rect 766 612 767 616
rect 771 612 772 616
rect 766 611 772 612
rect 110 608 116 609
rect 206 607 212 608
rect 206 603 207 607
rect 211 603 212 607
rect 206 602 212 603
rect 302 607 308 608
rect 302 603 303 607
rect 307 603 308 607
rect 302 602 308 603
rect 430 607 436 608
rect 430 603 431 607
rect 435 603 436 607
rect 430 602 436 603
rect 558 607 564 608
rect 558 603 559 607
rect 563 603 564 607
rect 558 602 564 603
rect 567 607 573 608
rect 567 603 568 607
rect 572 606 573 607
rect 864 606 866 628
rect 963 627 964 628
rect 968 627 969 631
rect 963 626 969 627
rect 1107 631 1116 632
rect 1107 627 1108 631
rect 1115 627 1116 631
rect 1107 626 1116 627
rect 1126 631 1132 632
rect 1126 627 1127 631
rect 1131 630 1132 631
rect 1259 631 1265 632
rect 1259 630 1260 631
rect 1131 628 1260 630
rect 1131 627 1132 628
rect 1126 626 1132 627
rect 1259 627 1260 628
rect 1264 627 1265 631
rect 1259 626 1265 627
rect 1278 631 1284 632
rect 1278 627 1279 631
rect 1283 630 1284 631
rect 1419 631 1425 632
rect 1419 630 1420 631
rect 1283 628 1420 630
rect 1283 627 1284 628
rect 1278 626 1284 627
rect 1419 627 1420 628
rect 1424 627 1425 631
rect 1419 626 1425 627
rect 1579 631 1585 632
rect 1579 627 1580 631
rect 1584 630 1585 631
rect 1606 631 1612 632
rect 1606 630 1607 631
rect 1584 628 1607 630
rect 1584 627 1585 628
rect 1579 626 1585 627
rect 1606 627 1607 628
rect 1611 627 1612 631
rect 1606 626 1612 627
rect 1723 631 1729 632
rect 1723 627 1724 631
rect 1728 630 1729 631
rect 1742 631 1748 632
rect 1742 630 1743 631
rect 1728 628 1743 630
rect 1728 627 1729 628
rect 1723 626 1729 627
rect 1742 627 1743 628
rect 1747 627 1748 631
rect 1806 629 1807 633
rect 1811 629 1812 633
rect 1974 632 1975 636
rect 1979 632 1980 636
rect 1974 631 1980 632
rect 2238 636 2244 637
rect 2238 632 2239 636
rect 2243 632 2244 636
rect 2238 631 2244 632
rect 2478 636 2484 637
rect 2478 632 2479 636
rect 2483 632 2484 636
rect 2478 631 2484 632
rect 2686 636 2692 637
rect 2686 632 2687 636
rect 2691 632 2692 636
rect 2686 631 2692 632
rect 2878 636 2884 637
rect 2878 632 2879 636
rect 2883 632 2884 636
rect 2878 631 2884 632
rect 3054 636 3060 637
rect 3054 632 3055 636
rect 3059 632 3060 636
rect 3054 631 3060 632
rect 3222 636 3228 637
rect 3222 632 3223 636
rect 3227 632 3228 636
rect 3222 631 3228 632
rect 3366 636 3372 637
rect 3366 632 3367 636
rect 3371 632 3372 636
rect 3366 631 3372 632
rect 3462 633 3468 634
rect 1806 628 1812 629
rect 3462 629 3463 633
rect 3467 629 3468 633
rect 3462 628 3468 629
rect 1742 626 1748 627
rect 2046 627 2052 628
rect 2046 623 2047 627
rect 2051 623 2052 627
rect 2046 622 2052 623
rect 2158 627 2164 628
rect 2158 623 2159 627
rect 2163 626 2164 627
rect 2550 627 2556 628
rect 2163 624 2281 626
rect 2163 623 2164 624
rect 2158 622 2164 623
rect 2550 623 2551 627
rect 2555 623 2556 627
rect 2550 622 2556 623
rect 2758 627 2764 628
rect 2758 623 2759 627
rect 2763 623 2764 627
rect 2758 622 2764 623
rect 2950 627 2956 628
rect 2950 623 2951 627
rect 2955 623 2956 627
rect 2950 622 2956 623
rect 3126 627 3132 628
rect 3126 623 3127 627
rect 3131 623 3132 627
rect 3126 622 3132 623
rect 3190 627 3196 628
rect 3190 623 3191 627
rect 3195 626 3196 627
rect 3438 627 3444 628
rect 3195 624 3265 626
rect 3195 623 3196 624
rect 3190 622 3196 623
rect 3438 623 3439 627
rect 3443 623 3444 627
rect 3438 622 3444 623
rect 1974 617 1980 618
rect 910 616 916 617
rect 910 612 911 616
rect 915 612 916 616
rect 910 611 916 612
rect 1054 616 1060 617
rect 1054 612 1055 616
rect 1059 612 1060 616
rect 1054 611 1060 612
rect 1206 616 1212 617
rect 1206 612 1207 616
rect 1211 612 1212 616
rect 1206 611 1212 612
rect 1366 616 1372 617
rect 1366 612 1367 616
rect 1371 612 1372 616
rect 1366 611 1372 612
rect 1526 616 1532 617
rect 1526 612 1527 616
rect 1531 612 1532 616
rect 1526 611 1532 612
rect 1670 616 1676 617
rect 1670 612 1671 616
rect 1675 612 1676 616
rect 1806 616 1812 617
rect 1670 611 1676 612
rect 1766 613 1772 614
rect 1766 609 1767 613
rect 1771 609 1772 613
rect 1806 612 1807 616
rect 1811 612 1812 616
rect 1974 613 1975 617
rect 1979 613 1980 617
rect 1974 612 1980 613
rect 2238 617 2244 618
rect 2238 613 2239 617
rect 2243 613 2244 617
rect 2238 612 2244 613
rect 2478 617 2484 618
rect 2478 613 2479 617
rect 2483 613 2484 617
rect 2478 612 2484 613
rect 2686 617 2692 618
rect 2686 613 2687 617
rect 2691 613 2692 617
rect 2686 612 2692 613
rect 2878 617 2884 618
rect 2878 613 2879 617
rect 2883 613 2884 617
rect 2878 612 2884 613
rect 3054 617 3060 618
rect 3054 613 3055 617
rect 3059 613 3060 617
rect 3054 612 3060 613
rect 3222 617 3228 618
rect 3222 613 3223 617
rect 3227 613 3228 617
rect 3222 612 3228 613
rect 3366 617 3372 618
rect 3366 613 3367 617
rect 3371 613 3372 617
rect 3366 612 3372 613
rect 3462 616 3468 617
rect 3462 612 3463 616
rect 3467 612 3468 616
rect 1806 611 1812 612
rect 3462 611 3468 612
rect 1766 608 1772 609
rect 572 604 665 606
rect 841 604 866 606
rect 982 607 988 608
rect 572 603 573 604
rect 567 602 573 603
rect 982 603 983 607
rect 987 603 988 607
rect 982 602 988 603
rect 1126 607 1132 608
rect 1126 603 1127 607
rect 1131 603 1132 607
rect 1126 602 1132 603
rect 1278 607 1284 608
rect 1278 603 1279 607
rect 1283 603 1284 607
rect 1278 602 1284 603
rect 1286 607 1292 608
rect 1286 603 1287 607
rect 1291 606 1292 607
rect 1446 607 1452 608
rect 1291 604 1409 606
rect 1291 603 1292 604
rect 1286 602 1292 603
rect 1446 603 1447 607
rect 1451 606 1452 607
rect 1606 607 1612 608
rect 1451 604 1569 606
rect 1451 603 1452 604
rect 1446 602 1452 603
rect 1606 603 1607 607
rect 1611 606 1612 607
rect 1611 604 1713 606
rect 1611 603 1612 604
rect 1606 602 1612 603
rect 134 597 140 598
rect 110 596 116 597
rect 110 592 111 596
rect 115 592 116 596
rect 134 593 135 597
rect 139 593 140 597
rect 134 592 140 593
rect 230 597 236 598
rect 230 593 231 597
rect 235 593 236 597
rect 230 592 236 593
rect 358 597 364 598
rect 358 593 359 597
rect 363 593 364 597
rect 358 592 364 593
rect 486 597 492 598
rect 486 593 487 597
rect 491 593 492 597
rect 486 592 492 593
rect 622 597 628 598
rect 622 593 623 597
rect 627 593 628 597
rect 622 592 628 593
rect 766 597 772 598
rect 766 593 767 597
rect 771 593 772 597
rect 766 592 772 593
rect 910 597 916 598
rect 910 593 911 597
rect 915 593 916 597
rect 910 592 916 593
rect 1054 597 1060 598
rect 1054 593 1055 597
rect 1059 593 1060 597
rect 1054 592 1060 593
rect 1206 597 1212 598
rect 1206 593 1207 597
rect 1211 593 1212 597
rect 1206 592 1212 593
rect 1366 597 1372 598
rect 1366 593 1367 597
rect 1371 593 1372 597
rect 1366 592 1372 593
rect 1526 597 1532 598
rect 1526 593 1527 597
rect 1531 593 1532 597
rect 1526 592 1532 593
rect 1670 597 1676 598
rect 1670 593 1671 597
rect 1675 593 1676 597
rect 1670 592 1676 593
rect 1766 596 1772 597
rect 1766 592 1767 596
rect 1771 592 1772 596
rect 110 591 116 592
rect 1766 591 1772 592
rect 1806 564 1812 565
rect 3462 564 3468 565
rect 1806 560 1807 564
rect 1811 560 1812 564
rect 1806 559 1812 560
rect 1894 563 1900 564
rect 1894 559 1895 563
rect 1899 559 1900 563
rect 1894 558 1900 559
rect 2014 563 2020 564
rect 2014 559 2015 563
rect 2019 559 2020 563
rect 2014 558 2020 559
rect 2142 563 2148 564
rect 2142 559 2143 563
rect 2147 559 2148 563
rect 2142 558 2148 559
rect 2278 563 2284 564
rect 2278 559 2279 563
rect 2283 559 2284 563
rect 2278 558 2284 559
rect 2422 563 2428 564
rect 2422 559 2423 563
rect 2427 559 2428 563
rect 2422 558 2428 559
rect 2566 563 2572 564
rect 2566 559 2567 563
rect 2571 559 2572 563
rect 2566 558 2572 559
rect 2718 563 2724 564
rect 2718 559 2719 563
rect 2723 559 2724 563
rect 2718 558 2724 559
rect 2870 563 2876 564
rect 2870 559 2871 563
rect 2875 559 2876 563
rect 2870 558 2876 559
rect 3030 563 3036 564
rect 3030 559 3031 563
rect 3035 559 3036 563
rect 3030 558 3036 559
rect 3198 563 3204 564
rect 3198 559 3199 563
rect 3203 559 3204 563
rect 3198 558 3204 559
rect 3366 563 3372 564
rect 3366 559 3367 563
rect 3371 559 3372 563
rect 3462 560 3463 564
rect 3467 560 3468 564
rect 3366 558 3372 559
rect 3430 559 3436 560
rect 3462 559 3468 560
rect 1966 555 1972 556
rect 1966 551 1967 555
rect 1971 551 1972 555
rect 1966 550 1972 551
rect 1974 555 1980 556
rect 1974 551 1975 555
rect 1979 554 1980 555
rect 2094 555 2100 556
rect 1979 552 2057 554
rect 1979 551 1980 552
rect 1974 550 1980 551
rect 2094 551 2095 555
rect 2099 554 2100 555
rect 2222 555 2228 556
rect 2099 552 2185 554
rect 2099 551 2100 552
rect 2094 550 2100 551
rect 2222 551 2223 555
rect 2227 554 2228 555
rect 2410 555 2416 556
rect 2227 552 2321 554
rect 2227 551 2228 552
rect 2222 550 2228 551
rect 2410 551 2411 555
rect 2415 554 2416 555
rect 2838 555 2844 556
rect 2415 552 2465 554
rect 2415 551 2416 552
rect 2410 550 2416 551
rect 2638 551 2644 552
rect 110 548 116 549
rect 1766 548 1772 549
rect 110 544 111 548
rect 115 544 116 548
rect 110 543 116 544
rect 134 547 140 548
rect 134 543 135 547
rect 139 543 140 547
rect 246 547 252 548
rect 134 542 140 543
rect 198 543 204 544
rect 198 539 199 543
rect 203 539 204 543
rect 246 543 247 547
rect 251 543 252 547
rect 246 542 252 543
rect 406 547 412 548
rect 406 543 407 547
rect 411 543 412 547
rect 406 542 412 543
rect 582 547 588 548
rect 582 543 583 547
rect 587 543 588 547
rect 582 542 588 543
rect 766 547 772 548
rect 766 543 767 547
rect 771 543 772 547
rect 766 542 772 543
rect 950 547 956 548
rect 950 543 951 547
rect 955 543 956 547
rect 950 542 956 543
rect 1134 547 1140 548
rect 1134 543 1135 547
rect 1139 543 1140 547
rect 1134 542 1140 543
rect 1318 547 1324 548
rect 1318 543 1319 547
rect 1323 543 1324 547
rect 1318 542 1324 543
rect 1502 547 1508 548
rect 1502 543 1503 547
rect 1507 543 1508 547
rect 1502 542 1508 543
rect 1670 547 1676 548
rect 1670 543 1671 547
rect 1675 543 1676 547
rect 1766 544 1767 548
rect 1771 544 1772 548
rect 1766 543 1772 544
rect 1806 547 1812 548
rect 1806 543 1807 547
rect 1811 543 1812 547
rect 2638 547 2639 551
rect 2643 547 2644 551
rect 2638 546 2644 547
rect 2790 551 2796 552
rect 2790 547 2791 551
rect 2795 547 2796 551
rect 2838 551 2839 555
rect 2843 554 2844 555
rect 3138 555 3144 556
rect 2843 552 2913 554
rect 2843 551 2844 552
rect 2838 550 2844 551
rect 3102 551 3108 552
rect 2790 546 2796 547
rect 3102 547 3103 551
rect 3107 547 3108 551
rect 3138 551 3139 555
rect 3143 554 3144 555
rect 3430 555 3431 559
rect 3435 555 3436 559
rect 3430 554 3436 555
rect 3143 552 3241 554
rect 3432 552 3441 554
rect 3143 551 3144 552
rect 3138 550 3144 551
rect 3102 546 3108 547
rect 3462 547 3468 548
rect 1670 542 1676 543
rect 1806 542 1812 543
rect 1894 544 1900 545
rect 1894 540 1895 544
rect 1899 540 1900 544
rect 198 538 204 539
rect 214 539 220 540
rect 200 536 209 538
rect 214 535 215 539
rect 219 538 220 539
rect 326 539 332 540
rect 219 536 289 538
rect 219 535 220 536
rect 214 534 220 535
rect 326 535 327 539
rect 331 538 332 539
rect 742 539 748 540
rect 331 536 449 538
rect 331 535 332 536
rect 326 534 332 535
rect 654 535 660 536
rect 110 531 116 532
rect 110 527 111 531
rect 115 527 116 531
rect 654 531 655 535
rect 659 531 660 535
rect 742 535 743 539
rect 747 538 748 539
rect 1110 539 1116 540
rect 1894 539 1900 540
rect 2014 544 2020 545
rect 2014 540 2015 544
rect 2019 540 2020 544
rect 2014 539 2020 540
rect 2142 544 2148 545
rect 2142 540 2143 544
rect 2147 540 2148 544
rect 2142 539 2148 540
rect 2278 544 2284 545
rect 2278 540 2279 544
rect 2283 540 2284 544
rect 2278 539 2284 540
rect 2422 544 2428 545
rect 2422 540 2423 544
rect 2427 540 2428 544
rect 2422 539 2428 540
rect 2566 544 2572 545
rect 2566 540 2567 544
rect 2571 540 2572 544
rect 2566 539 2572 540
rect 2718 544 2724 545
rect 2718 540 2719 544
rect 2723 540 2724 544
rect 2718 539 2724 540
rect 2870 544 2876 545
rect 2870 540 2871 544
rect 2875 540 2876 544
rect 2870 539 2876 540
rect 3030 544 3036 545
rect 3030 540 3031 544
rect 3035 540 3036 544
rect 3030 539 3036 540
rect 3198 544 3204 545
rect 3198 540 3199 544
rect 3203 540 3204 544
rect 3198 539 3204 540
rect 3366 544 3372 545
rect 3366 540 3367 544
rect 3371 540 3372 544
rect 3462 543 3463 547
rect 3467 543 3468 547
rect 3462 542 3468 543
rect 3366 539 3372 540
rect 747 536 809 538
rect 747 535 748 536
rect 742 534 748 535
rect 1022 535 1028 536
rect 654 530 660 531
rect 1022 531 1023 535
rect 1027 531 1028 535
rect 1110 535 1111 539
rect 1115 538 1116 539
rect 1115 536 1177 538
rect 1115 535 1116 536
rect 1110 534 1116 535
rect 1390 535 1396 536
rect 1022 530 1028 531
rect 1390 531 1391 535
rect 1395 531 1396 535
rect 1390 530 1396 531
rect 1574 535 1580 536
rect 1574 531 1575 535
rect 1579 531 1580 535
rect 1574 530 1580 531
rect 1742 535 1748 536
rect 1742 531 1743 535
rect 1747 531 1748 535
rect 3138 535 3144 536
rect 3138 534 3139 535
rect 2924 532 3139 534
rect 1742 530 1748 531
rect 1766 531 1772 532
rect 110 526 116 527
rect 134 528 140 529
rect 134 524 135 528
rect 139 524 140 528
rect 134 523 140 524
rect 246 528 252 529
rect 246 524 247 528
rect 251 524 252 528
rect 246 523 252 524
rect 406 528 412 529
rect 406 524 407 528
rect 411 524 412 528
rect 406 523 412 524
rect 582 528 588 529
rect 582 524 583 528
rect 587 524 588 528
rect 582 523 588 524
rect 766 528 772 529
rect 766 524 767 528
rect 771 524 772 528
rect 766 523 772 524
rect 950 528 956 529
rect 950 524 951 528
rect 955 524 956 528
rect 950 523 956 524
rect 1134 528 1140 529
rect 1134 524 1135 528
rect 1139 524 1140 528
rect 1134 523 1140 524
rect 1318 528 1324 529
rect 1318 524 1319 528
rect 1323 524 1324 528
rect 1318 523 1324 524
rect 1502 528 1508 529
rect 1502 524 1503 528
rect 1507 524 1508 528
rect 1502 523 1508 524
rect 1670 528 1676 529
rect 1670 524 1671 528
rect 1675 524 1676 528
rect 1766 527 1767 531
rect 1771 527 1772 531
rect 2924 530 2926 532
rect 3138 531 3139 532
rect 3143 531 3144 535
rect 3138 530 3144 531
rect 2923 529 2929 530
rect 1766 526 1772 527
rect 1947 527 1953 528
rect 1670 523 1676 524
rect 1947 523 1948 527
rect 1952 526 1953 527
rect 1974 527 1980 528
rect 1974 526 1975 527
rect 1952 524 1975 526
rect 1952 523 1953 524
rect 1947 522 1953 523
rect 1974 523 1975 524
rect 1979 523 1980 527
rect 1974 522 1980 523
rect 2067 527 2073 528
rect 2067 523 2068 527
rect 2072 526 2073 527
rect 2094 527 2100 528
rect 2094 526 2095 527
rect 2072 524 2095 526
rect 2072 523 2073 524
rect 2067 522 2073 523
rect 2094 523 2095 524
rect 2099 523 2100 527
rect 2094 522 2100 523
rect 2195 527 2201 528
rect 2195 523 2196 527
rect 2200 526 2201 527
rect 2222 527 2228 528
rect 2222 526 2223 527
rect 2200 524 2223 526
rect 2200 523 2201 524
rect 2195 522 2201 523
rect 2222 523 2223 524
rect 2227 523 2228 527
rect 2222 522 2228 523
rect 2331 527 2337 528
rect 2331 523 2332 527
rect 2336 526 2337 527
rect 2410 527 2416 528
rect 2410 526 2411 527
rect 2336 524 2411 526
rect 2336 523 2337 524
rect 2331 522 2337 523
rect 2410 523 2411 524
rect 2415 523 2416 527
rect 2410 522 2416 523
rect 2430 527 2436 528
rect 2430 523 2431 527
rect 2435 526 2436 527
rect 2475 527 2481 528
rect 2475 526 2476 527
rect 2435 524 2476 526
rect 2435 523 2436 524
rect 2430 522 2436 523
rect 2475 523 2476 524
rect 2480 523 2481 527
rect 2475 522 2481 523
rect 2619 527 2625 528
rect 2619 523 2620 527
rect 2624 526 2625 527
rect 2630 527 2636 528
rect 2630 526 2631 527
rect 2624 524 2631 526
rect 2624 523 2625 524
rect 2619 522 2625 523
rect 2630 523 2631 524
rect 2635 523 2636 527
rect 2630 522 2636 523
rect 2638 527 2644 528
rect 2638 523 2639 527
rect 2643 526 2644 527
rect 2771 527 2777 528
rect 2771 526 2772 527
rect 2643 524 2772 526
rect 2643 523 2644 524
rect 2638 522 2644 523
rect 2771 523 2772 524
rect 2776 523 2777 527
rect 2923 525 2924 529
rect 2928 525 2929 529
rect 2923 524 2929 525
rect 3078 527 3089 528
rect 2771 522 2777 523
rect 3078 523 3079 527
rect 3083 523 3084 527
rect 3088 523 3089 527
rect 3078 522 3089 523
rect 3102 527 3108 528
rect 3102 523 3103 527
rect 3107 526 3108 527
rect 3251 527 3257 528
rect 3251 526 3252 527
rect 3107 524 3252 526
rect 3107 523 3108 524
rect 3102 522 3108 523
rect 3251 523 3252 524
rect 3256 523 3257 527
rect 3251 522 3257 523
rect 3419 527 3425 528
rect 3419 523 3420 527
rect 3424 526 3425 527
rect 3430 527 3436 528
rect 3430 526 3431 527
rect 3424 524 3431 526
rect 3424 523 3425 524
rect 3419 522 3425 523
rect 3430 523 3431 524
rect 3435 523 3436 527
rect 3430 522 3436 523
rect 742 519 748 520
rect 742 518 743 519
rect 460 516 743 518
rect 460 514 462 516
rect 742 515 743 516
rect 747 515 748 519
rect 1446 519 1452 520
rect 1446 518 1447 519
rect 742 514 748 515
rect 1372 516 1447 518
rect 1372 514 1374 516
rect 1446 515 1447 516
rect 1451 515 1452 519
rect 1446 514 1452 515
rect 2206 519 2212 520
rect 2206 515 2207 519
rect 2211 518 2212 519
rect 2211 516 2294 518
rect 2211 515 2212 516
rect 2206 514 2212 515
rect 2292 514 2294 516
rect 459 513 465 514
rect 187 511 193 512
rect 187 507 188 511
rect 192 510 193 511
rect 214 511 220 512
rect 214 510 215 511
rect 192 508 215 510
rect 192 507 193 508
rect 187 506 193 507
rect 214 507 215 508
rect 219 507 220 511
rect 214 506 220 507
rect 299 511 305 512
rect 299 507 300 511
rect 304 510 305 511
rect 326 511 332 512
rect 326 510 327 511
rect 304 508 327 510
rect 304 507 305 508
rect 299 506 305 507
rect 326 507 327 508
rect 331 507 332 511
rect 459 509 460 513
rect 464 509 465 513
rect 1371 513 1377 514
rect 459 508 465 509
rect 634 511 641 512
rect 326 506 332 507
rect 634 507 635 511
rect 640 507 641 511
rect 634 506 641 507
rect 654 511 660 512
rect 654 507 655 511
rect 659 510 660 511
rect 819 511 825 512
rect 819 510 820 511
rect 659 508 820 510
rect 659 507 660 508
rect 654 506 660 507
rect 819 507 820 508
rect 824 507 825 511
rect 819 506 825 507
rect 982 511 988 512
rect 982 507 983 511
rect 987 510 988 511
rect 1003 511 1009 512
rect 1003 510 1004 511
rect 987 508 1004 510
rect 987 507 988 508
rect 982 506 988 507
rect 1003 507 1004 508
rect 1008 507 1009 511
rect 1003 506 1009 507
rect 1022 511 1028 512
rect 1022 507 1023 511
rect 1027 510 1028 511
rect 1187 511 1193 512
rect 1187 510 1188 511
rect 1027 508 1188 510
rect 1027 507 1028 508
rect 1022 506 1028 507
rect 1187 507 1188 508
rect 1192 507 1193 511
rect 1371 509 1372 513
rect 1376 509 1377 513
rect 2291 513 2297 514
rect 1371 508 1377 509
rect 1390 511 1396 512
rect 1187 506 1193 507
rect 1390 507 1391 511
rect 1395 510 1396 511
rect 1555 511 1561 512
rect 1555 510 1556 511
rect 1395 508 1556 510
rect 1395 507 1396 508
rect 1390 506 1396 507
rect 1555 507 1556 508
rect 1560 507 1561 511
rect 1555 506 1561 507
rect 1574 511 1580 512
rect 1574 507 1575 511
rect 1579 510 1580 511
rect 1723 511 1729 512
rect 1723 510 1724 511
rect 1579 508 1724 510
rect 1579 507 1580 508
rect 1574 506 1580 507
rect 1723 507 1724 508
rect 1728 507 1729 511
rect 1723 506 1729 507
rect 2187 511 2193 512
rect 2187 507 2188 511
rect 2192 510 2193 511
rect 2192 508 2278 510
rect 2291 509 2292 513
rect 2296 509 2297 513
rect 2291 508 2297 509
rect 2310 511 2316 512
rect 2192 507 2193 508
rect 2187 506 2193 507
rect 2276 502 2278 508
rect 2310 507 2311 511
rect 2315 510 2316 511
rect 2411 511 2417 512
rect 2411 510 2412 511
rect 2315 508 2412 510
rect 2315 507 2316 508
rect 2310 506 2316 507
rect 2411 507 2412 508
rect 2416 507 2417 511
rect 2411 506 2417 507
rect 2539 511 2545 512
rect 2539 507 2540 511
rect 2544 510 2545 511
rect 2567 511 2573 512
rect 2567 510 2568 511
rect 2544 508 2568 510
rect 2544 507 2545 508
rect 2539 506 2545 507
rect 2567 507 2568 508
rect 2572 507 2573 511
rect 2567 506 2573 507
rect 2667 511 2676 512
rect 2667 507 2668 511
rect 2675 507 2676 511
rect 2667 506 2676 507
rect 2790 511 2796 512
rect 2790 507 2791 511
rect 2795 510 2796 511
rect 2803 511 2809 512
rect 2803 510 2804 511
rect 2795 508 2804 510
rect 2795 507 2796 508
rect 2790 506 2796 507
rect 2803 507 2804 508
rect 2808 507 2809 511
rect 2803 506 2809 507
rect 2931 511 2937 512
rect 2931 507 2932 511
rect 2936 510 2937 511
rect 2950 511 2956 512
rect 2936 508 2946 510
rect 2936 507 2937 508
rect 2931 506 2937 507
rect 2944 502 2946 508
rect 2950 507 2951 511
rect 2955 510 2956 511
rect 3059 511 3065 512
rect 3059 510 3060 511
rect 2955 508 3060 510
rect 2955 507 2956 508
rect 2950 506 2956 507
rect 3059 507 3060 508
rect 3064 507 3065 511
rect 3059 506 3065 507
rect 3187 511 3196 512
rect 3187 507 3188 511
rect 3195 507 3196 511
rect 3187 506 3196 507
rect 3206 511 3212 512
rect 3206 507 3207 511
rect 3211 510 3212 511
rect 3315 511 3321 512
rect 3315 510 3316 511
rect 3211 508 3316 510
rect 3211 507 3212 508
rect 3206 506 3212 507
rect 3315 507 3316 508
rect 3320 507 3321 511
rect 3315 506 3321 507
rect 3419 511 3425 512
rect 3419 507 3420 511
rect 3424 510 3425 511
rect 3438 511 3444 512
rect 3438 510 3439 511
rect 3424 508 3439 510
rect 3424 507 3425 508
rect 3419 506 3425 507
rect 3438 507 3439 508
rect 3443 507 3444 511
rect 3438 506 3444 507
rect 3102 503 3108 504
rect 3102 502 3103 503
rect 2276 500 2446 502
rect 2944 500 3103 502
rect 2134 496 2140 497
rect 299 495 305 496
rect 299 491 300 495
rect 304 494 305 495
rect 318 495 324 496
rect 304 492 314 494
rect 304 491 305 492
rect 299 490 305 491
rect 312 486 314 492
rect 318 491 319 495
rect 323 494 324 495
rect 451 495 457 496
rect 451 494 452 495
rect 323 492 452 494
rect 323 491 324 492
rect 318 490 324 491
rect 451 491 452 492
rect 456 491 457 495
rect 451 490 457 491
rect 470 495 476 496
rect 470 491 471 495
rect 475 494 476 495
rect 619 495 625 496
rect 619 494 620 495
rect 475 492 620 494
rect 475 491 476 492
rect 470 490 476 491
rect 619 491 620 492
rect 624 491 625 495
rect 619 490 625 491
rect 787 495 793 496
rect 787 491 788 495
rect 792 494 793 495
rect 814 495 820 496
rect 814 494 815 495
rect 792 492 815 494
rect 792 491 793 492
rect 787 490 793 491
rect 814 491 815 492
rect 819 491 820 495
rect 814 490 820 491
rect 955 495 961 496
rect 955 491 956 495
rect 960 494 961 495
rect 998 495 1004 496
rect 998 494 999 495
rect 960 492 999 494
rect 960 491 961 492
rect 955 490 961 491
rect 998 491 999 492
rect 1003 491 1004 495
rect 998 490 1004 491
rect 1115 495 1121 496
rect 1115 491 1116 495
rect 1120 494 1121 495
rect 1186 495 1192 496
rect 1120 492 1182 494
rect 1120 491 1121 492
rect 1115 490 1121 491
rect 1180 486 1182 492
rect 1186 491 1187 495
rect 1191 494 1192 495
rect 1275 495 1281 496
rect 1275 494 1276 495
rect 1191 492 1276 494
rect 1191 491 1192 492
rect 1186 490 1192 491
rect 1275 491 1276 492
rect 1280 491 1281 495
rect 1275 490 1281 491
rect 1427 495 1433 496
rect 1427 491 1428 495
rect 1432 494 1433 495
rect 1471 495 1477 496
rect 1471 494 1472 495
rect 1432 492 1472 494
rect 1432 491 1433 492
rect 1427 490 1433 491
rect 1471 491 1472 492
rect 1476 491 1477 495
rect 1471 490 1477 491
rect 1579 495 1585 496
rect 1579 491 1580 495
rect 1584 494 1585 495
rect 1606 495 1612 496
rect 1606 494 1607 495
rect 1584 492 1607 494
rect 1584 491 1585 492
rect 1579 490 1585 491
rect 1606 491 1607 492
rect 1611 491 1612 495
rect 1606 490 1612 491
rect 1723 495 1729 496
rect 1723 491 1724 495
rect 1728 494 1729 495
rect 1742 495 1748 496
rect 1742 494 1743 495
rect 1728 492 1743 494
rect 1728 491 1729 492
rect 1723 490 1729 491
rect 1742 491 1743 492
rect 1747 491 1748 495
rect 1742 490 1748 491
rect 1806 493 1812 494
rect 1806 489 1807 493
rect 1811 489 1812 493
rect 2134 492 2135 496
rect 2139 492 2140 496
rect 2134 491 2140 492
rect 2238 496 2244 497
rect 2238 492 2239 496
rect 2243 492 2244 496
rect 2238 491 2244 492
rect 2358 496 2364 497
rect 2358 492 2359 496
rect 2363 492 2364 496
rect 2358 491 2364 492
rect 1806 488 1812 489
rect 2206 487 2212 488
rect 312 484 681 486
rect 1180 484 1306 486
rect 246 480 252 481
rect 110 477 116 478
rect 110 473 111 477
rect 115 473 116 477
rect 246 476 247 480
rect 251 476 252 480
rect 246 475 252 476
rect 398 480 404 481
rect 398 476 399 480
rect 403 476 404 480
rect 398 475 404 476
rect 566 480 572 481
rect 566 476 567 480
rect 571 476 572 480
rect 566 475 572 476
rect 110 472 116 473
rect 318 471 324 472
rect 318 467 319 471
rect 323 467 324 471
rect 318 466 324 467
rect 470 471 476 472
rect 470 467 471 471
rect 475 467 476 471
rect 470 466 476 467
rect 634 471 640 472
rect 634 467 635 471
rect 639 467 640 471
rect 679 470 681 484
rect 734 480 740 481
rect 734 476 735 480
rect 739 476 740 480
rect 734 475 740 476
rect 902 480 908 481
rect 902 476 903 480
rect 907 476 908 480
rect 902 475 908 476
rect 1062 480 1068 481
rect 1062 476 1063 480
rect 1067 476 1068 480
rect 1062 475 1068 476
rect 1222 480 1228 481
rect 1222 476 1223 480
rect 1227 476 1228 480
rect 1222 475 1228 476
rect 814 471 820 472
rect 679 468 777 470
rect 634 466 640 467
rect 814 467 815 471
rect 819 470 820 471
rect 1186 471 1192 472
rect 1186 470 1187 471
rect 819 468 945 470
rect 1137 468 1187 470
rect 819 467 820 468
rect 814 466 820 467
rect 1186 467 1187 468
rect 1191 467 1192 471
rect 1186 466 1192 467
rect 1294 471 1300 472
rect 1294 467 1295 471
rect 1299 467 1300 471
rect 1304 470 1306 484
rect 2206 483 2207 487
rect 2211 483 2212 487
rect 2206 482 2212 483
rect 2310 487 2316 488
rect 2310 483 2311 487
rect 2315 483 2316 487
rect 2310 482 2316 483
rect 2430 487 2436 488
rect 2430 483 2431 487
rect 2435 483 2436 487
rect 2444 486 2446 500
rect 3102 499 3103 500
rect 3107 499 3108 503
rect 3102 498 3108 499
rect 2486 496 2492 497
rect 2486 492 2487 496
rect 2491 492 2492 496
rect 2486 491 2492 492
rect 2614 496 2620 497
rect 2614 492 2615 496
rect 2619 492 2620 496
rect 2614 491 2620 492
rect 2750 496 2756 497
rect 2750 492 2751 496
rect 2755 492 2756 496
rect 2750 491 2756 492
rect 2878 496 2884 497
rect 2878 492 2879 496
rect 2883 492 2884 496
rect 2878 491 2884 492
rect 3006 496 3012 497
rect 3006 492 3007 496
rect 3011 492 3012 496
rect 3006 491 3012 492
rect 3134 496 3140 497
rect 3134 492 3135 496
rect 3139 492 3140 496
rect 3134 491 3140 492
rect 3262 496 3268 497
rect 3262 492 3263 496
rect 3267 492 3268 496
rect 3262 491 3268 492
rect 3366 496 3372 497
rect 3366 492 3367 496
rect 3371 492 3372 496
rect 3366 491 3372 492
rect 3462 493 3468 494
rect 3462 489 3463 493
rect 3467 489 3468 493
rect 3462 488 3468 489
rect 2567 487 2573 488
rect 2444 484 2529 486
rect 2430 482 2436 483
rect 2567 483 2568 487
rect 2572 486 2573 487
rect 2822 487 2828 488
rect 2572 484 2657 486
rect 2572 483 2573 484
rect 2567 482 2573 483
rect 2822 483 2823 487
rect 2827 483 2828 487
rect 2822 482 2828 483
rect 2950 487 2956 488
rect 2950 483 2951 487
rect 2955 483 2956 487
rect 2950 482 2956 483
rect 3078 487 3084 488
rect 3078 483 3079 487
rect 3083 483 3084 487
rect 3078 482 3084 483
rect 3206 487 3212 488
rect 3206 483 3207 487
rect 3211 483 3212 487
rect 3206 482 3212 483
rect 3326 487 3332 488
rect 3326 483 3327 487
rect 3331 483 3332 487
rect 3326 482 3332 483
rect 3430 487 3436 488
rect 3430 483 3431 487
rect 3435 483 3436 487
rect 3430 482 3436 483
rect 1374 480 1380 481
rect 1374 476 1375 480
rect 1379 476 1380 480
rect 1374 475 1380 476
rect 1526 480 1532 481
rect 1526 476 1527 480
rect 1531 476 1532 480
rect 1526 475 1532 476
rect 1670 480 1676 481
rect 1670 476 1671 480
rect 1675 476 1676 480
rect 1670 475 1676 476
rect 1766 477 1772 478
rect 2134 477 2140 478
rect 1766 473 1767 477
rect 1771 473 1772 477
rect 1766 472 1772 473
rect 1806 476 1812 477
rect 1806 472 1807 476
rect 1811 472 1812 476
rect 2134 473 2135 477
rect 2139 473 2140 477
rect 2134 472 2140 473
rect 2238 477 2244 478
rect 2238 473 2239 477
rect 2243 473 2244 477
rect 2238 472 2244 473
rect 2358 477 2364 478
rect 2358 473 2359 477
rect 2363 473 2364 477
rect 2358 472 2364 473
rect 2486 477 2492 478
rect 2486 473 2487 477
rect 2491 473 2492 477
rect 2486 472 2492 473
rect 2614 477 2620 478
rect 2614 473 2615 477
rect 2619 473 2620 477
rect 2614 472 2620 473
rect 2750 477 2756 478
rect 2750 473 2751 477
rect 2755 473 2756 477
rect 2750 472 2756 473
rect 2878 477 2884 478
rect 2878 473 2879 477
rect 2883 473 2884 477
rect 2878 472 2884 473
rect 3006 477 3012 478
rect 3006 473 3007 477
rect 3011 473 3012 477
rect 3006 472 3012 473
rect 3134 477 3140 478
rect 3134 473 3135 477
rect 3139 473 3140 477
rect 3134 472 3140 473
rect 3262 477 3268 478
rect 3262 473 3263 477
rect 3267 473 3268 477
rect 3262 472 3268 473
rect 3366 477 3372 478
rect 3366 473 3367 477
rect 3371 473 3372 477
rect 3366 472 3372 473
rect 3462 476 3468 477
rect 3462 472 3463 476
rect 3467 472 3468 476
rect 1471 471 1477 472
rect 1304 468 1417 470
rect 1294 466 1300 467
rect 1471 467 1472 471
rect 1476 470 1477 471
rect 1606 471 1612 472
rect 1806 471 1812 472
rect 3462 471 3468 472
rect 1476 468 1569 470
rect 1476 467 1477 468
rect 1471 466 1477 467
rect 1606 467 1607 471
rect 1611 470 1612 471
rect 1611 468 1713 470
rect 1611 467 1612 468
rect 1606 466 1612 467
rect 246 461 252 462
rect 110 460 116 461
rect 110 456 111 460
rect 115 456 116 460
rect 246 457 247 461
rect 251 457 252 461
rect 246 456 252 457
rect 398 461 404 462
rect 398 457 399 461
rect 403 457 404 461
rect 398 456 404 457
rect 566 461 572 462
rect 566 457 567 461
rect 571 457 572 461
rect 566 456 572 457
rect 734 461 740 462
rect 734 457 735 461
rect 739 457 740 461
rect 734 456 740 457
rect 902 461 908 462
rect 902 457 903 461
rect 907 457 908 461
rect 902 456 908 457
rect 1062 461 1068 462
rect 1062 457 1063 461
rect 1067 457 1068 461
rect 1062 456 1068 457
rect 1222 461 1228 462
rect 1222 457 1223 461
rect 1227 457 1228 461
rect 1222 456 1228 457
rect 1374 461 1380 462
rect 1374 457 1375 461
rect 1379 457 1380 461
rect 1374 456 1380 457
rect 1526 461 1532 462
rect 1526 457 1527 461
rect 1531 457 1532 461
rect 1526 456 1532 457
rect 1670 461 1676 462
rect 1670 457 1671 461
rect 1675 457 1676 461
rect 1670 456 1676 457
rect 1766 460 1772 461
rect 1766 456 1767 460
rect 1771 456 1772 460
rect 110 455 116 456
rect 1766 455 1772 456
rect 1806 424 1812 425
rect 3462 424 3468 425
rect 1806 420 1807 424
rect 1811 420 1812 424
rect 1806 419 1812 420
rect 2238 423 2244 424
rect 2238 419 2239 423
rect 2243 419 2244 423
rect 2238 418 2244 419
rect 2334 423 2340 424
rect 2334 419 2335 423
rect 2339 419 2340 423
rect 2334 418 2340 419
rect 2446 423 2452 424
rect 2446 419 2447 423
rect 2451 419 2452 423
rect 2446 418 2452 419
rect 2558 423 2564 424
rect 2558 419 2559 423
rect 2563 419 2564 423
rect 2558 418 2564 419
rect 2678 423 2684 424
rect 2678 419 2679 423
rect 2683 419 2684 423
rect 2678 418 2684 419
rect 2798 423 2804 424
rect 2798 419 2799 423
rect 2803 419 2804 423
rect 2798 418 2804 419
rect 2910 423 2916 424
rect 2910 419 2911 423
rect 2915 419 2916 423
rect 2910 418 2916 419
rect 3022 423 3028 424
rect 3022 419 3023 423
rect 3027 419 3028 423
rect 3022 418 3028 419
rect 3142 423 3148 424
rect 3142 419 3143 423
rect 3147 419 3148 423
rect 3142 418 3148 419
rect 3262 423 3268 424
rect 3262 419 3263 423
rect 3267 419 3268 423
rect 3262 418 3268 419
rect 3366 423 3372 424
rect 3366 419 3367 423
rect 3371 419 3372 423
rect 3462 420 3463 424
rect 3467 420 3468 424
rect 3462 419 3468 420
rect 3366 418 3372 419
rect 2670 415 2676 416
rect 110 412 116 413
rect 1766 412 1772 413
rect 110 408 111 412
rect 115 408 116 412
rect 110 407 116 408
rect 518 411 524 412
rect 518 407 519 411
rect 523 407 524 411
rect 518 406 524 407
rect 614 411 620 412
rect 614 407 615 411
rect 619 407 620 411
rect 614 406 620 407
rect 718 411 724 412
rect 718 407 719 411
rect 723 407 724 411
rect 718 406 724 407
rect 822 411 828 412
rect 822 407 823 411
rect 827 407 828 411
rect 822 406 828 407
rect 926 411 932 412
rect 926 407 927 411
rect 931 407 932 411
rect 926 406 932 407
rect 1022 411 1028 412
rect 1022 407 1023 411
rect 1027 407 1028 411
rect 1022 406 1028 407
rect 1126 411 1132 412
rect 1126 407 1127 411
rect 1131 407 1132 411
rect 1126 406 1132 407
rect 1230 411 1236 412
rect 1230 407 1231 411
rect 1235 407 1236 411
rect 1230 406 1236 407
rect 1334 411 1340 412
rect 1334 407 1335 411
rect 1339 407 1340 411
rect 1334 406 1340 407
rect 1438 411 1444 412
rect 1438 407 1439 411
rect 1443 407 1444 411
rect 1766 408 1767 412
rect 1771 408 1772 412
rect 2406 411 2412 412
rect 2313 408 2322 410
rect 1766 407 1772 408
rect 1806 407 1812 408
rect 1438 406 1444 407
rect 798 403 804 404
rect 590 399 596 400
rect 110 395 116 396
rect 110 391 111 395
rect 115 391 116 395
rect 590 395 591 399
rect 595 395 596 399
rect 590 394 596 395
rect 686 399 692 400
rect 686 395 687 399
rect 691 395 692 399
rect 798 399 799 403
rect 803 402 804 403
rect 998 403 1004 404
rect 803 400 865 402
rect 803 399 804 400
rect 798 398 804 399
rect 998 399 999 403
rect 1003 399 1004 403
rect 1206 403 1212 404
rect 998 398 1004 399
rect 1094 399 1100 400
rect 686 394 692 395
rect 110 390 116 391
rect 518 392 524 393
rect 518 388 519 392
rect 523 388 524 392
rect 518 387 524 388
rect 614 392 620 393
rect 614 388 615 392
rect 619 388 620 392
rect 614 387 620 388
rect 718 392 724 393
rect 718 388 719 392
rect 723 388 724 392
rect 792 390 794 397
rect 1094 395 1095 399
rect 1099 395 1100 399
rect 1094 394 1100 395
rect 1198 399 1204 400
rect 1198 395 1199 399
rect 1203 395 1204 399
rect 1206 399 1207 403
rect 1211 402 1212 403
rect 1414 403 1420 404
rect 1211 400 1273 402
rect 1211 399 1212 400
rect 1206 398 1212 399
rect 1406 399 1412 400
rect 1198 394 1204 395
rect 1406 395 1407 399
rect 1411 395 1412 399
rect 1414 399 1415 403
rect 1419 402 1420 403
rect 1806 403 1807 407
rect 1811 403 1812 407
rect 1806 402 1812 403
rect 2238 404 2244 405
rect 1419 400 1481 402
rect 2238 400 2239 404
rect 2243 400 2244 404
rect 1419 399 1420 400
rect 2238 399 2244 400
rect 1414 398 1420 399
rect 1406 394 1412 395
rect 1766 395 1772 396
rect 822 392 828 393
rect 792 388 810 390
rect 718 387 724 388
rect 798 383 804 384
rect 798 382 799 383
rect 572 380 799 382
rect 572 378 574 380
rect 798 379 799 380
rect 803 379 804 383
rect 808 382 810 388
rect 822 388 823 392
rect 827 388 828 392
rect 822 387 828 388
rect 926 392 932 393
rect 926 388 927 392
rect 931 388 932 392
rect 926 387 932 388
rect 1022 392 1028 393
rect 1022 388 1023 392
rect 1027 388 1028 392
rect 1022 387 1028 388
rect 1126 392 1132 393
rect 1126 388 1127 392
rect 1131 388 1132 392
rect 1126 387 1132 388
rect 1230 392 1236 393
rect 1230 388 1231 392
rect 1235 388 1236 392
rect 1230 387 1236 388
rect 1334 392 1340 393
rect 1334 388 1335 392
rect 1339 388 1340 392
rect 1334 387 1340 388
rect 1438 392 1444 393
rect 1438 388 1439 392
rect 1443 388 1444 392
rect 1766 391 1767 395
rect 1771 391 1772 395
rect 2320 394 2322 408
rect 2406 407 2407 411
rect 2411 407 2412 411
rect 2406 406 2412 407
rect 2518 411 2524 412
rect 2518 407 2519 411
rect 2523 407 2524 411
rect 2518 406 2524 407
rect 2630 411 2636 412
rect 2630 407 2631 411
rect 2635 407 2636 411
rect 2670 411 2671 415
rect 2675 414 2676 415
rect 3102 415 3108 416
rect 2675 412 2721 414
rect 2675 411 2676 412
rect 2670 410 2676 411
rect 2870 411 2876 412
rect 2630 406 2636 407
rect 2870 407 2871 411
rect 2875 407 2876 411
rect 2870 406 2876 407
rect 2982 411 2988 412
rect 2982 407 2983 411
rect 2987 407 2988 411
rect 2982 406 2988 407
rect 3094 411 3100 412
rect 3094 407 3095 411
rect 3099 407 3100 411
rect 3102 411 3103 415
rect 3107 414 3108 415
rect 3438 415 3444 416
rect 3107 412 3185 414
rect 3107 411 3108 412
rect 3102 410 3108 411
rect 3334 411 3340 412
rect 3094 406 3100 407
rect 3334 407 3335 411
rect 3339 407 3340 411
rect 3438 411 3439 415
rect 3443 411 3444 415
rect 3438 410 3444 411
rect 3334 406 3340 407
rect 3462 407 3468 408
rect 2334 404 2340 405
rect 2334 400 2335 404
rect 2339 400 2340 404
rect 2334 399 2340 400
rect 2446 404 2452 405
rect 2446 400 2447 404
rect 2451 400 2452 404
rect 2446 399 2452 400
rect 2558 404 2564 405
rect 2558 400 2559 404
rect 2563 400 2564 404
rect 2558 399 2564 400
rect 2678 404 2684 405
rect 2678 400 2679 404
rect 2683 400 2684 404
rect 2678 399 2684 400
rect 2798 404 2804 405
rect 2798 400 2799 404
rect 2803 400 2804 404
rect 2798 399 2804 400
rect 2910 404 2916 405
rect 2910 400 2911 404
rect 2915 400 2916 404
rect 2910 399 2916 400
rect 3022 404 3028 405
rect 3022 400 3023 404
rect 3027 400 3028 404
rect 3022 399 3028 400
rect 3142 404 3148 405
rect 3142 400 3143 404
rect 3147 400 3148 404
rect 3142 399 3148 400
rect 3262 404 3268 405
rect 3262 400 3263 404
rect 3267 400 3268 404
rect 3262 399 3268 400
rect 3366 404 3372 405
rect 3366 400 3367 404
rect 3371 400 3372 404
rect 3462 403 3463 407
rect 3467 403 3468 407
rect 3462 402 3468 403
rect 3366 399 3372 400
rect 2320 392 2361 394
rect 1766 390 1772 391
rect 2359 390 2361 392
rect 2359 389 2393 390
rect 2359 388 2388 389
rect 1438 387 1444 388
rect 2291 387 2297 388
rect 1206 383 1212 384
rect 1206 382 1207 383
rect 808 380 982 382
rect 798 378 804 379
rect 980 378 982 380
rect 1076 380 1207 382
rect 1076 378 1078 380
rect 1206 379 1207 380
rect 1211 379 1212 383
rect 1414 383 1420 384
rect 1414 382 1415 383
rect 1206 378 1212 379
rect 1284 380 1415 382
rect 1284 378 1286 380
rect 1414 379 1415 380
rect 1419 379 1420 383
rect 2291 383 2292 387
rect 2296 386 2297 387
rect 2296 384 2330 386
rect 2387 385 2388 388
rect 2392 385 2393 389
rect 2387 384 2393 385
rect 2406 387 2412 388
rect 2296 383 2297 384
rect 2291 382 2297 383
rect 1414 378 1420 379
rect 2328 378 2330 384
rect 2406 383 2407 387
rect 2411 386 2412 387
rect 2499 387 2505 388
rect 2499 386 2500 387
rect 2411 384 2500 386
rect 2411 383 2412 384
rect 2406 382 2412 383
rect 2499 383 2500 384
rect 2504 383 2505 387
rect 2499 382 2505 383
rect 2518 387 2524 388
rect 2518 383 2519 387
rect 2523 386 2524 387
rect 2611 387 2617 388
rect 2611 386 2612 387
rect 2523 384 2612 386
rect 2523 383 2524 384
rect 2518 382 2524 383
rect 2611 383 2612 384
rect 2616 383 2617 387
rect 2611 382 2617 383
rect 2630 387 2636 388
rect 2630 383 2631 387
rect 2635 386 2636 387
rect 2731 387 2737 388
rect 2731 386 2732 387
rect 2635 384 2732 386
rect 2635 383 2636 384
rect 2630 382 2636 383
rect 2731 383 2732 384
rect 2736 383 2737 387
rect 2731 382 2737 383
rect 2822 387 2828 388
rect 2822 383 2823 387
rect 2827 386 2828 387
rect 2851 387 2857 388
rect 2851 386 2852 387
rect 2827 384 2852 386
rect 2827 383 2828 384
rect 2822 382 2828 383
rect 2851 383 2852 384
rect 2856 383 2857 387
rect 2851 382 2857 383
rect 2963 387 2969 388
rect 2963 383 2964 387
rect 2968 386 2969 387
rect 2974 387 2980 388
rect 2974 386 2975 387
rect 2968 384 2975 386
rect 2968 383 2969 384
rect 2963 382 2969 383
rect 2974 383 2975 384
rect 2979 383 2980 387
rect 2974 382 2980 383
rect 2982 387 2988 388
rect 2982 383 2983 387
rect 2987 386 2988 387
rect 3075 387 3081 388
rect 3075 386 3076 387
rect 2987 384 3076 386
rect 2987 383 2988 384
rect 2982 382 2988 383
rect 3075 383 3076 384
rect 3080 383 3081 387
rect 3075 382 3081 383
rect 3094 387 3100 388
rect 3094 383 3095 387
rect 3099 386 3100 387
rect 3195 387 3201 388
rect 3195 386 3196 387
rect 3099 384 3196 386
rect 3099 383 3100 384
rect 3094 382 3100 383
rect 3195 383 3196 384
rect 3200 383 3201 387
rect 3195 382 3201 383
rect 3315 387 3321 388
rect 3315 383 3316 387
rect 3320 386 3321 387
rect 3326 387 3332 388
rect 3326 386 3327 387
rect 3320 384 3327 386
rect 3320 383 3321 384
rect 3315 382 3321 383
rect 3326 383 3327 384
rect 3331 383 3332 387
rect 3326 382 3332 383
rect 3419 387 3425 388
rect 3419 383 3420 387
rect 3424 386 3425 387
rect 3430 387 3436 388
rect 3430 386 3431 387
rect 3424 384 3431 386
rect 3424 383 3425 384
rect 3419 382 3425 383
rect 3430 383 3431 384
rect 3435 383 3436 387
rect 3430 382 3436 383
rect 2438 379 2444 380
rect 2438 378 2439 379
rect 571 377 577 378
rect 571 373 572 377
rect 576 373 577 377
rect 979 377 985 378
rect 571 372 577 373
rect 590 375 596 376
rect 590 371 591 375
rect 595 374 596 375
rect 667 375 673 376
rect 667 374 668 375
rect 595 372 668 374
rect 595 371 596 372
rect 590 370 596 371
rect 667 371 668 372
rect 672 371 673 375
rect 667 370 673 371
rect 686 375 692 376
rect 686 371 687 375
rect 691 374 692 375
rect 771 375 777 376
rect 771 374 772 375
rect 691 372 772 374
rect 691 371 692 372
rect 686 370 692 371
rect 771 371 772 372
rect 776 371 777 375
rect 771 370 777 371
rect 875 375 881 376
rect 875 371 876 375
rect 880 374 881 375
rect 886 375 892 376
rect 886 374 887 375
rect 880 372 887 374
rect 880 371 881 372
rect 875 370 881 371
rect 886 371 887 372
rect 891 371 892 375
rect 979 373 980 377
rect 984 373 985 377
rect 979 372 985 373
rect 1075 377 1081 378
rect 1075 373 1076 377
rect 1080 373 1081 377
rect 1283 377 1289 378
rect 1075 372 1081 373
rect 1094 375 1100 376
rect 886 370 892 371
rect 1094 371 1095 375
rect 1099 374 1100 375
rect 1179 375 1185 376
rect 1179 374 1180 375
rect 1099 372 1180 374
rect 1099 371 1100 372
rect 1094 370 1100 371
rect 1179 371 1180 372
rect 1184 371 1185 375
rect 1283 373 1284 377
rect 1288 373 1289 377
rect 2328 376 2439 378
rect 1283 372 1289 373
rect 1294 375 1300 376
rect 1179 370 1185 371
rect 1294 371 1295 375
rect 1299 374 1300 375
rect 1387 375 1393 376
rect 1387 374 1388 375
rect 1299 372 1388 374
rect 1299 371 1300 372
rect 1294 370 1300 371
rect 1387 371 1388 372
rect 1392 371 1393 375
rect 1387 370 1393 371
rect 1406 375 1412 376
rect 1406 371 1407 375
rect 1411 374 1412 375
rect 1491 375 1497 376
rect 1491 374 1492 375
rect 1411 372 1492 374
rect 1411 371 1412 372
rect 1406 370 1412 371
rect 1491 371 1492 372
rect 1496 371 1497 375
rect 2438 375 2439 376
rect 2443 375 2444 379
rect 2438 374 2444 375
rect 1491 370 1497 371
rect 2115 371 2121 372
rect 2115 367 2116 371
rect 2120 370 2121 371
rect 2134 371 2140 372
rect 2120 368 2130 370
rect 2120 367 2121 368
rect 2115 366 2121 367
rect 2128 362 2130 368
rect 2134 367 2135 371
rect 2139 370 2140 371
rect 2203 371 2209 372
rect 2203 370 2204 371
rect 2139 368 2204 370
rect 2139 367 2140 368
rect 2134 366 2140 367
rect 2203 367 2204 368
rect 2208 367 2209 371
rect 2203 366 2209 367
rect 2222 371 2228 372
rect 2222 367 2223 371
rect 2227 370 2228 371
rect 2299 371 2305 372
rect 2299 370 2300 371
rect 2227 368 2300 370
rect 2227 367 2228 368
rect 2222 366 2228 367
rect 2299 367 2300 368
rect 2304 367 2305 371
rect 2299 366 2305 367
rect 2318 371 2324 372
rect 2318 367 2319 371
rect 2323 370 2324 371
rect 2411 371 2417 372
rect 2411 370 2412 371
rect 2323 368 2412 370
rect 2323 367 2324 368
rect 2318 366 2324 367
rect 2411 367 2412 368
rect 2416 367 2417 371
rect 2411 366 2417 367
rect 2430 371 2436 372
rect 2430 367 2431 371
rect 2435 370 2436 371
rect 2531 371 2537 372
rect 2531 370 2532 371
rect 2435 368 2532 370
rect 2435 367 2436 368
rect 2430 366 2436 367
rect 2531 367 2532 368
rect 2536 367 2537 371
rect 2531 366 2537 367
rect 2667 371 2673 372
rect 2667 367 2668 371
rect 2672 370 2673 371
rect 2694 371 2700 372
rect 2694 370 2695 371
rect 2672 368 2695 370
rect 2672 367 2673 368
rect 2667 366 2673 367
rect 2694 367 2695 368
rect 2699 367 2700 371
rect 2694 366 2700 367
rect 2811 371 2817 372
rect 2811 367 2812 371
rect 2816 370 2817 371
rect 2870 371 2876 372
rect 2870 370 2871 371
rect 2816 368 2871 370
rect 2816 367 2817 368
rect 2811 366 2817 367
rect 2870 367 2871 368
rect 2875 367 2876 371
rect 2870 366 2876 367
rect 2963 371 2969 372
rect 2963 367 2964 371
rect 2968 370 2969 371
rect 2990 371 2996 372
rect 2990 370 2991 371
rect 2968 368 2991 370
rect 2968 367 2969 368
rect 2963 366 2969 367
rect 2990 367 2991 368
rect 2995 367 2996 371
rect 2990 366 2996 367
rect 3115 371 3121 372
rect 3115 367 3116 371
rect 3120 370 3121 371
rect 3158 371 3164 372
rect 3158 370 3159 371
rect 3120 368 3159 370
rect 3120 367 3121 368
rect 3115 366 3121 367
rect 3158 367 3159 368
rect 3163 367 3164 371
rect 3158 366 3164 367
rect 3166 371 3172 372
rect 3166 367 3167 371
rect 3171 370 3172 371
rect 3275 371 3281 372
rect 3275 370 3276 371
rect 3171 368 3276 370
rect 3171 367 3172 368
rect 3166 366 3172 367
rect 3275 367 3276 368
rect 3280 367 3281 371
rect 3275 366 3281 367
rect 3419 371 3425 372
rect 3419 367 3420 371
rect 3424 370 3425 371
rect 3438 371 3444 372
rect 3438 370 3439 371
rect 3424 368 3439 370
rect 3424 367 3425 368
rect 3419 366 3425 367
rect 3438 367 3439 368
rect 3443 367 3444 371
rect 3438 366 3444 367
rect 2422 363 2428 364
rect 2422 362 2423 363
rect 2128 360 2423 362
rect 523 359 529 360
rect 523 355 524 359
rect 528 358 529 359
rect 542 359 548 360
rect 528 356 538 358
rect 528 355 529 356
rect 523 354 529 355
rect 536 350 538 356
rect 542 355 543 359
rect 547 358 548 359
rect 611 359 617 360
rect 611 358 612 359
rect 547 356 612 358
rect 547 355 548 356
rect 542 354 548 355
rect 611 355 612 356
rect 616 355 617 359
rect 611 354 617 355
rect 630 359 636 360
rect 630 355 631 359
rect 635 358 636 359
rect 699 359 705 360
rect 699 358 700 359
rect 635 356 700 358
rect 635 355 636 356
rect 630 354 636 355
rect 699 355 700 356
rect 704 355 705 359
rect 699 354 705 355
rect 727 359 733 360
rect 727 355 728 359
rect 732 358 733 359
rect 787 359 793 360
rect 787 358 788 359
rect 732 356 788 358
rect 732 355 733 356
rect 727 354 733 355
rect 787 355 788 356
rect 792 355 793 359
rect 787 354 793 355
rect 806 359 812 360
rect 806 355 807 359
rect 811 358 812 359
rect 875 359 881 360
rect 875 358 876 359
rect 811 356 876 358
rect 811 355 812 356
rect 806 354 812 355
rect 875 355 876 356
rect 880 355 881 359
rect 875 354 881 355
rect 963 359 969 360
rect 963 355 964 359
rect 968 358 969 359
rect 990 359 996 360
rect 990 358 991 359
rect 968 356 991 358
rect 968 355 969 356
rect 963 354 969 355
rect 990 355 991 356
rect 995 355 996 359
rect 990 354 996 355
rect 1051 359 1057 360
rect 1051 355 1052 359
rect 1056 358 1057 359
rect 1078 359 1084 360
rect 1078 358 1079 359
rect 1056 356 1079 358
rect 1056 355 1057 356
rect 1051 354 1057 355
rect 1078 355 1079 356
rect 1083 355 1084 359
rect 1078 354 1084 355
rect 1139 359 1145 360
rect 1139 355 1140 359
rect 1144 358 1145 359
rect 1198 359 1204 360
rect 1144 356 1194 358
rect 1144 355 1145 356
rect 1139 354 1145 355
rect 638 351 644 352
rect 638 350 639 351
rect 536 348 639 350
rect 638 347 639 348
rect 643 347 644 351
rect 1192 350 1194 356
rect 1198 355 1199 359
rect 1203 358 1204 359
rect 1227 359 1233 360
rect 1227 358 1228 359
rect 1203 356 1228 358
rect 1203 355 1204 356
rect 1198 354 1204 355
rect 1227 355 1228 356
rect 1232 355 1233 359
rect 1227 354 1233 355
rect 1246 359 1252 360
rect 1246 355 1247 359
rect 1251 358 1252 359
rect 1315 359 1321 360
rect 1315 358 1316 359
rect 1251 356 1316 358
rect 1251 355 1252 356
rect 1246 354 1252 355
rect 1315 355 1316 356
rect 1320 355 1321 359
rect 2422 359 2423 360
rect 2427 359 2428 363
rect 2422 358 2428 359
rect 1315 354 1321 355
rect 2062 356 2068 357
rect 1806 353 1812 354
rect 1192 348 1258 350
rect 1806 349 1807 353
rect 1811 349 1812 353
rect 2062 352 2063 356
rect 2067 352 2068 356
rect 2062 351 2068 352
rect 2150 356 2156 357
rect 2150 352 2151 356
rect 2155 352 2156 356
rect 2150 351 2156 352
rect 2246 356 2252 357
rect 2246 352 2247 356
rect 2251 352 2252 356
rect 2246 351 2252 352
rect 2358 356 2364 357
rect 2358 352 2359 356
rect 2363 352 2364 356
rect 2358 351 2364 352
rect 2478 356 2484 357
rect 2478 352 2479 356
rect 2483 352 2484 356
rect 2478 351 2484 352
rect 2614 356 2620 357
rect 2614 352 2615 356
rect 2619 352 2620 356
rect 2614 351 2620 352
rect 2758 356 2764 357
rect 2758 352 2759 356
rect 2763 352 2764 356
rect 2758 351 2764 352
rect 2910 356 2916 357
rect 2910 352 2911 356
rect 2915 352 2916 356
rect 2910 351 2916 352
rect 3062 356 3068 357
rect 3062 352 3063 356
rect 3067 352 3068 356
rect 3062 351 3068 352
rect 3222 356 3228 357
rect 3222 352 3223 356
rect 3227 352 3228 356
rect 3222 351 3228 352
rect 3366 356 3372 357
rect 3366 352 3367 356
rect 3371 352 3372 356
rect 3366 351 3372 352
rect 3462 353 3468 354
rect 1806 348 1812 349
rect 3462 349 3463 353
rect 3467 349 3468 353
rect 3462 348 3468 349
rect 638 346 644 347
rect 470 344 476 345
rect 110 341 116 342
rect 110 337 111 341
rect 115 337 116 341
rect 470 340 471 344
rect 475 340 476 344
rect 470 339 476 340
rect 558 344 564 345
rect 558 340 559 344
rect 563 340 564 344
rect 558 339 564 340
rect 646 344 652 345
rect 646 340 647 344
rect 651 340 652 344
rect 646 339 652 340
rect 734 344 740 345
rect 734 340 735 344
rect 739 340 740 344
rect 734 339 740 340
rect 822 344 828 345
rect 822 340 823 344
rect 827 340 828 344
rect 822 339 828 340
rect 910 344 916 345
rect 910 340 911 344
rect 915 340 916 344
rect 910 339 916 340
rect 998 344 1004 345
rect 998 340 999 344
rect 1003 340 1004 344
rect 998 339 1004 340
rect 1086 344 1092 345
rect 1086 340 1087 344
rect 1091 340 1092 344
rect 1086 339 1092 340
rect 1174 344 1180 345
rect 1174 340 1175 344
rect 1179 340 1180 344
rect 1174 339 1180 340
rect 110 336 116 337
rect 542 335 548 336
rect 542 331 543 335
rect 547 331 548 335
rect 542 330 548 331
rect 630 335 636 336
rect 630 331 631 335
rect 635 331 636 335
rect 727 335 733 336
rect 727 334 728 335
rect 721 332 728 334
rect 630 330 636 331
rect 727 331 728 332
rect 732 331 733 335
rect 727 330 733 331
rect 806 335 812 336
rect 806 331 807 335
rect 811 331 812 335
rect 806 330 812 331
rect 886 335 892 336
rect 886 331 887 335
rect 891 331 892 335
rect 886 330 892 331
rect 902 335 908 336
rect 902 331 903 335
rect 907 334 908 335
rect 990 335 996 336
rect 907 332 953 334
rect 907 331 908 332
rect 902 330 908 331
rect 990 331 991 335
rect 995 334 996 335
rect 1078 335 1084 336
rect 995 332 1041 334
rect 995 331 996 332
rect 990 330 996 331
rect 1078 331 1079 335
rect 1083 334 1084 335
rect 1246 335 1252 336
rect 1083 332 1129 334
rect 1083 331 1084 332
rect 1078 330 1084 331
rect 1246 331 1247 335
rect 1251 331 1252 335
rect 1256 334 1258 348
rect 2134 347 2140 348
rect 1262 344 1268 345
rect 1262 340 1263 344
rect 1267 340 1268 344
rect 2134 343 2135 347
rect 2139 343 2140 347
rect 2134 342 2140 343
rect 2222 347 2228 348
rect 2222 343 2223 347
rect 2227 343 2228 347
rect 2222 342 2228 343
rect 2318 347 2324 348
rect 2318 343 2319 347
rect 2323 343 2324 347
rect 2318 342 2324 343
rect 2430 347 2436 348
rect 2430 343 2431 347
rect 2435 343 2436 347
rect 2430 342 2436 343
rect 2438 347 2444 348
rect 2438 343 2439 347
rect 2443 346 2444 347
rect 2678 347 2684 348
rect 2443 344 2521 346
rect 2443 343 2444 344
rect 2438 342 2444 343
rect 2678 343 2679 347
rect 2683 343 2684 347
rect 2678 342 2684 343
rect 2694 347 2700 348
rect 2694 343 2695 347
rect 2699 346 2700 347
rect 2974 347 2980 348
rect 2699 344 2801 346
rect 2699 343 2700 344
rect 2694 342 2700 343
rect 2974 343 2975 347
rect 2979 343 2980 347
rect 2974 342 2980 343
rect 2990 347 2996 348
rect 2990 343 2991 347
rect 2995 346 2996 347
rect 3158 347 3164 348
rect 2995 344 3105 346
rect 2995 343 2996 344
rect 2990 342 2996 343
rect 3158 343 3159 347
rect 3163 346 3164 347
rect 3430 347 3436 348
rect 3163 344 3265 346
rect 3163 343 3164 344
rect 3158 342 3164 343
rect 3430 343 3431 347
rect 3435 343 3436 347
rect 3430 342 3436 343
rect 1262 339 1268 340
rect 1766 341 1772 342
rect 1766 337 1767 341
rect 1771 337 1772 341
rect 2062 337 2068 338
rect 1766 336 1772 337
rect 1806 336 1812 337
rect 1256 332 1305 334
rect 1806 332 1807 336
rect 1811 332 1812 336
rect 2062 333 2063 337
rect 2067 333 2068 337
rect 2062 332 2068 333
rect 2150 337 2156 338
rect 2150 333 2151 337
rect 2155 333 2156 337
rect 2150 332 2156 333
rect 2246 337 2252 338
rect 2246 333 2247 337
rect 2251 333 2252 337
rect 2246 332 2252 333
rect 2358 337 2364 338
rect 2358 333 2359 337
rect 2363 333 2364 337
rect 2358 332 2364 333
rect 2478 337 2484 338
rect 2478 333 2479 337
rect 2483 333 2484 337
rect 2478 332 2484 333
rect 2614 337 2620 338
rect 2614 333 2615 337
rect 2619 333 2620 337
rect 2614 332 2620 333
rect 2758 337 2764 338
rect 2758 333 2759 337
rect 2763 333 2764 337
rect 2758 332 2764 333
rect 2910 337 2916 338
rect 2910 333 2911 337
rect 2915 333 2916 337
rect 2910 332 2916 333
rect 3062 337 3068 338
rect 3062 333 3063 337
rect 3067 333 3068 337
rect 3062 332 3068 333
rect 3222 337 3228 338
rect 3222 333 3223 337
rect 3227 333 3228 337
rect 3222 332 3228 333
rect 3366 337 3372 338
rect 3366 333 3367 337
rect 3371 333 3372 337
rect 3366 332 3372 333
rect 3462 336 3468 337
rect 3462 332 3463 336
rect 3467 332 3468 336
rect 1806 331 1812 332
rect 3462 331 3468 332
rect 1246 330 1252 331
rect 470 325 476 326
rect 110 324 116 325
rect 110 320 111 324
rect 115 320 116 324
rect 470 321 471 325
rect 475 321 476 325
rect 470 320 476 321
rect 558 325 564 326
rect 558 321 559 325
rect 563 321 564 325
rect 558 320 564 321
rect 646 325 652 326
rect 646 321 647 325
rect 651 321 652 325
rect 646 320 652 321
rect 734 325 740 326
rect 734 321 735 325
rect 739 321 740 325
rect 734 320 740 321
rect 822 325 828 326
rect 822 321 823 325
rect 827 321 828 325
rect 822 320 828 321
rect 910 325 916 326
rect 910 321 911 325
rect 915 321 916 325
rect 910 320 916 321
rect 998 325 1004 326
rect 998 321 999 325
rect 1003 321 1004 325
rect 998 320 1004 321
rect 1086 325 1092 326
rect 1086 321 1087 325
rect 1091 321 1092 325
rect 1086 320 1092 321
rect 1174 325 1180 326
rect 1174 321 1175 325
rect 1179 321 1180 325
rect 1174 320 1180 321
rect 1262 325 1268 326
rect 1262 321 1263 325
rect 1267 321 1268 325
rect 1262 320 1268 321
rect 1766 324 1772 325
rect 1766 320 1767 324
rect 1771 320 1772 324
rect 110 319 116 320
rect 1766 319 1772 320
rect 1806 288 1812 289
rect 3462 288 3468 289
rect 1806 284 1807 288
rect 1811 284 1812 288
rect 1806 283 1812 284
rect 1926 287 1932 288
rect 1926 283 1927 287
rect 1931 283 1932 287
rect 1926 282 1932 283
rect 2038 287 2044 288
rect 2038 283 2039 287
rect 2043 283 2044 287
rect 2038 282 2044 283
rect 2166 287 2172 288
rect 2166 283 2167 287
rect 2171 283 2172 287
rect 2166 282 2172 283
rect 2302 287 2308 288
rect 2302 283 2303 287
rect 2307 283 2308 287
rect 2302 282 2308 283
rect 2446 287 2452 288
rect 2446 283 2447 287
rect 2451 283 2452 287
rect 2446 282 2452 283
rect 2598 287 2604 288
rect 2598 283 2599 287
rect 2603 283 2604 287
rect 2598 282 2604 283
rect 2758 287 2764 288
rect 2758 283 2759 287
rect 2763 283 2764 287
rect 2758 282 2764 283
rect 2918 287 2924 288
rect 2918 283 2919 287
rect 2923 283 2924 287
rect 2918 282 2924 283
rect 3086 287 3092 288
rect 3086 283 3087 287
rect 3091 283 3092 287
rect 3086 282 3092 283
rect 3254 287 3260 288
rect 3254 283 3255 287
rect 3259 283 3260 287
rect 3462 284 3463 288
rect 3467 284 3468 288
rect 3462 283 3468 284
rect 3254 282 3260 283
rect 2422 279 2428 280
rect 110 276 116 277
rect 1766 276 1772 277
rect 110 272 111 276
rect 115 272 116 276
rect 110 271 116 272
rect 278 275 284 276
rect 278 271 279 275
rect 283 271 284 275
rect 278 270 284 271
rect 366 275 372 276
rect 366 271 367 275
rect 371 271 372 275
rect 366 270 372 271
rect 462 275 468 276
rect 462 271 463 275
rect 467 271 468 275
rect 462 270 468 271
rect 558 275 564 276
rect 558 271 559 275
rect 563 271 564 275
rect 558 270 564 271
rect 654 275 660 276
rect 654 271 655 275
rect 659 271 660 275
rect 654 270 660 271
rect 750 275 756 276
rect 750 271 751 275
rect 755 271 756 275
rect 750 270 756 271
rect 846 275 852 276
rect 846 271 847 275
rect 851 271 852 275
rect 846 270 852 271
rect 942 275 948 276
rect 942 271 943 275
rect 947 271 948 275
rect 942 270 948 271
rect 1046 275 1052 276
rect 1046 271 1047 275
rect 1051 271 1052 275
rect 1046 270 1052 271
rect 1150 275 1156 276
rect 1150 271 1151 275
rect 1155 271 1156 275
rect 1766 272 1767 276
rect 1771 272 1772 276
rect 1998 275 2004 276
rect 1766 271 1772 272
rect 1806 271 1812 272
rect 1150 270 1156 271
rect 638 267 644 268
rect 350 263 356 264
rect 110 259 116 260
rect 110 255 111 259
rect 115 255 116 259
rect 350 259 351 263
rect 355 259 356 263
rect 350 258 356 259
rect 438 263 444 264
rect 438 259 439 263
rect 443 259 444 263
rect 438 258 444 259
rect 534 263 540 264
rect 534 259 535 263
rect 539 259 540 263
rect 534 258 540 259
rect 630 263 636 264
rect 630 259 631 263
rect 635 259 636 263
rect 638 263 639 267
rect 643 266 644 267
rect 1126 267 1132 268
rect 643 264 697 266
rect 643 263 644 264
rect 638 262 644 263
rect 822 263 828 264
rect 630 258 636 259
rect 822 259 823 263
rect 827 259 828 263
rect 822 258 828 259
rect 918 263 924 264
rect 918 259 919 263
rect 923 259 924 263
rect 918 258 924 259
rect 1014 263 1020 264
rect 1014 259 1015 263
rect 1019 259 1020 263
rect 1014 258 1020 259
rect 1118 263 1124 264
rect 1118 259 1119 263
rect 1123 259 1124 263
rect 1126 263 1127 267
rect 1131 266 1132 267
rect 1806 267 1807 271
rect 1811 267 1812 271
rect 1998 271 1999 275
rect 2003 271 2004 275
rect 1998 270 2004 271
rect 2110 275 2116 276
rect 2110 271 2111 275
rect 2115 271 2116 275
rect 2110 270 2116 271
rect 2238 275 2244 276
rect 2238 271 2239 275
rect 2243 271 2244 275
rect 2238 270 2244 271
rect 2374 275 2380 276
rect 2374 271 2375 275
rect 2379 271 2380 275
rect 2422 275 2423 279
rect 2427 278 2428 279
rect 3166 279 3172 280
rect 3166 278 3167 279
rect 2427 276 2489 278
rect 3161 276 3167 278
rect 2427 275 2428 276
rect 2422 274 2428 275
rect 2670 275 2676 276
rect 2374 270 2380 271
rect 2670 271 2671 275
rect 2675 271 2676 275
rect 2670 270 2676 271
rect 2830 275 2836 276
rect 2830 271 2831 275
rect 2835 271 2836 275
rect 2830 270 2836 271
rect 2990 275 2996 276
rect 2990 271 2991 275
rect 2995 271 2996 275
rect 3166 275 3167 276
rect 3171 275 3172 279
rect 3166 274 3172 275
rect 3247 279 3253 280
rect 3247 275 3248 279
rect 3252 278 3253 279
rect 3252 276 3297 278
rect 3252 275 3253 276
rect 3247 274 3253 275
rect 2990 270 2996 271
rect 3462 271 3468 272
rect 1806 266 1812 267
rect 1926 268 1932 269
rect 1131 264 1193 266
rect 1926 264 1927 268
rect 1931 264 1932 268
rect 1131 263 1132 264
rect 1926 263 1932 264
rect 2038 268 2044 269
rect 2038 264 2039 268
rect 2043 264 2044 268
rect 2038 263 2044 264
rect 2166 268 2172 269
rect 2166 264 2167 268
rect 2171 264 2172 268
rect 2166 263 2172 264
rect 2302 268 2308 269
rect 2302 264 2303 268
rect 2307 264 2308 268
rect 2302 263 2308 264
rect 2446 268 2452 269
rect 2446 264 2447 268
rect 2451 264 2452 268
rect 2446 263 2452 264
rect 2598 268 2604 269
rect 2598 264 2599 268
rect 2603 264 2604 268
rect 2598 263 2604 264
rect 2758 268 2764 269
rect 2758 264 2759 268
rect 2763 264 2764 268
rect 2758 263 2764 264
rect 2918 268 2924 269
rect 2918 264 2919 268
rect 2923 264 2924 268
rect 2918 263 2924 264
rect 3086 268 3092 269
rect 3086 264 3087 268
rect 3091 264 3092 268
rect 3086 263 3092 264
rect 3254 268 3260 269
rect 3254 264 3255 268
rect 3259 264 3260 268
rect 3462 267 3463 271
rect 3467 267 3468 271
rect 3462 266 3468 267
rect 3254 263 3260 264
rect 1126 262 1132 263
rect 1118 258 1124 259
rect 1766 259 1772 260
rect 110 254 116 255
rect 278 256 284 257
rect 278 252 279 256
rect 283 252 284 256
rect 278 251 284 252
rect 366 256 372 257
rect 366 252 367 256
rect 371 252 372 256
rect 366 251 372 252
rect 462 256 468 257
rect 462 252 463 256
rect 467 252 468 256
rect 462 251 468 252
rect 558 256 564 257
rect 558 252 559 256
rect 563 252 564 256
rect 558 251 564 252
rect 654 256 660 257
rect 654 252 655 256
rect 659 252 660 256
rect 654 251 660 252
rect 750 256 756 257
rect 750 252 751 256
rect 755 252 756 256
rect 750 251 756 252
rect 846 256 852 257
rect 846 252 847 256
rect 851 252 852 256
rect 846 251 852 252
rect 942 256 948 257
rect 942 252 943 256
rect 947 252 948 256
rect 942 251 948 252
rect 1046 256 1052 257
rect 1046 252 1047 256
rect 1051 252 1052 256
rect 1046 251 1052 252
rect 1150 256 1156 257
rect 1150 252 1151 256
rect 1155 252 1156 256
rect 1766 255 1767 259
rect 1771 255 1772 259
rect 1766 254 1772 255
rect 1150 251 1156 252
rect 1979 251 1985 252
rect 902 247 908 248
rect 902 246 903 247
rect 804 244 903 246
rect 804 242 806 244
rect 902 243 903 244
rect 907 243 908 247
rect 1979 247 1980 251
rect 1984 250 1985 251
rect 1998 251 2004 252
rect 1984 248 1994 250
rect 1984 247 1985 248
rect 1979 246 1985 247
rect 902 242 908 243
rect 1992 242 1994 248
rect 1998 247 1999 251
rect 2003 250 2004 251
rect 2091 251 2097 252
rect 2091 250 2092 251
rect 2003 248 2092 250
rect 2003 247 2004 248
rect 1998 246 2004 247
rect 2091 247 2092 248
rect 2096 247 2097 251
rect 2091 246 2097 247
rect 2110 251 2116 252
rect 2110 247 2111 251
rect 2115 250 2116 251
rect 2219 251 2225 252
rect 2219 250 2220 251
rect 2115 248 2220 250
rect 2115 247 2116 248
rect 2110 246 2116 247
rect 2219 247 2220 248
rect 2224 247 2225 251
rect 2219 246 2225 247
rect 2238 251 2244 252
rect 2238 247 2239 251
rect 2243 250 2244 251
rect 2355 251 2361 252
rect 2355 250 2356 251
rect 2243 248 2356 250
rect 2243 247 2244 248
rect 2238 246 2244 247
rect 2355 247 2356 248
rect 2360 247 2361 251
rect 2355 246 2361 247
rect 2374 251 2380 252
rect 2374 247 2375 251
rect 2379 250 2380 251
rect 2499 251 2505 252
rect 2499 250 2500 251
rect 2379 248 2500 250
rect 2379 247 2380 248
rect 2374 246 2380 247
rect 2499 247 2500 248
rect 2504 247 2505 251
rect 2499 246 2505 247
rect 2651 251 2657 252
rect 2651 247 2652 251
rect 2656 250 2657 251
rect 2678 251 2684 252
rect 2678 250 2679 251
rect 2656 248 2679 250
rect 2656 247 2657 248
rect 2651 246 2657 247
rect 2678 247 2679 248
rect 2683 247 2684 251
rect 2678 246 2684 247
rect 2811 251 2820 252
rect 2811 247 2812 251
rect 2819 247 2820 251
rect 2811 246 2820 247
rect 2830 251 2836 252
rect 2830 247 2831 251
rect 2835 250 2836 251
rect 2971 251 2977 252
rect 2971 250 2972 251
rect 2835 248 2972 250
rect 2835 247 2836 248
rect 2830 246 2836 247
rect 2971 247 2972 248
rect 2976 247 2977 251
rect 2971 246 2977 247
rect 2990 251 2996 252
rect 2990 247 2991 251
rect 2995 250 2996 251
rect 3139 251 3145 252
rect 3139 250 3140 251
rect 2995 248 3140 250
rect 2995 247 2996 248
rect 2990 246 2996 247
rect 3139 247 3140 248
rect 3144 247 3145 251
rect 3139 246 3145 247
rect 3307 251 3313 252
rect 3307 247 3308 251
rect 3312 250 3313 251
rect 3334 251 3340 252
rect 3334 250 3335 251
rect 3312 248 3335 250
rect 3312 247 3313 248
rect 3307 246 3313 247
rect 3334 247 3335 248
rect 3339 247 3340 251
rect 3334 246 3340 247
rect 2322 243 2328 244
rect 2322 242 2323 243
rect 803 241 809 242
rect 331 239 337 240
rect 331 235 332 239
rect 336 238 337 239
rect 350 239 356 240
rect 336 236 346 238
rect 336 235 337 236
rect 331 234 337 235
rect 344 230 346 236
rect 350 235 351 239
rect 355 238 356 239
rect 419 239 425 240
rect 419 238 420 239
rect 355 236 420 238
rect 355 235 356 236
rect 350 234 356 235
rect 419 235 420 236
rect 424 235 425 239
rect 419 234 425 235
rect 438 239 444 240
rect 438 235 439 239
rect 443 238 444 239
rect 515 239 521 240
rect 515 238 516 239
rect 443 236 516 238
rect 443 235 444 236
rect 438 234 444 235
rect 515 235 516 236
rect 520 235 521 239
rect 515 234 521 235
rect 534 239 540 240
rect 534 235 535 239
rect 539 238 540 239
rect 611 239 617 240
rect 611 238 612 239
rect 539 236 612 238
rect 539 235 540 236
rect 534 234 540 235
rect 611 235 612 236
rect 616 235 617 239
rect 611 234 617 235
rect 630 239 636 240
rect 630 235 631 239
rect 635 238 636 239
rect 707 239 713 240
rect 707 238 708 239
rect 635 236 708 238
rect 635 235 636 236
rect 630 234 636 235
rect 707 235 708 236
rect 712 235 713 239
rect 803 237 804 241
rect 808 237 809 241
rect 1992 240 2323 242
rect 803 236 809 237
rect 822 239 828 240
rect 707 234 713 235
rect 822 235 823 239
rect 827 238 828 239
rect 899 239 905 240
rect 899 238 900 239
rect 827 236 900 238
rect 827 235 828 236
rect 822 234 828 235
rect 899 235 900 236
rect 904 235 905 239
rect 899 234 905 235
rect 918 239 924 240
rect 918 235 919 239
rect 923 238 924 239
rect 995 239 1001 240
rect 995 238 996 239
rect 923 236 996 238
rect 923 235 924 236
rect 918 234 924 235
rect 995 235 996 236
rect 1000 235 1001 239
rect 995 234 1001 235
rect 1014 239 1020 240
rect 1014 235 1015 239
rect 1019 238 1020 239
rect 1099 239 1105 240
rect 1099 238 1100 239
rect 1019 236 1100 238
rect 1019 235 1020 236
rect 1014 234 1020 235
rect 1099 235 1100 236
rect 1104 235 1105 239
rect 1099 234 1105 235
rect 1118 239 1124 240
rect 1118 235 1119 239
rect 1123 238 1124 239
rect 1203 239 1209 240
rect 1203 238 1204 239
rect 1123 236 1204 238
rect 1123 235 1124 236
rect 1118 234 1124 235
rect 1203 235 1204 236
rect 1208 235 1209 239
rect 2322 239 2323 240
rect 2327 239 2328 243
rect 2322 238 2328 239
rect 1203 234 1209 235
rect 1883 235 1889 236
rect 590 231 596 232
rect 590 230 591 231
rect 344 228 591 230
rect 590 227 591 228
rect 595 227 596 231
rect 1126 231 1132 232
rect 1126 230 1127 231
rect 590 226 596 227
rect 892 228 1127 230
rect 892 226 894 228
rect 1126 227 1127 228
rect 1131 227 1132 231
rect 1883 231 1884 235
rect 1888 234 1889 235
rect 1902 235 1908 236
rect 1888 232 1898 234
rect 1888 231 1889 232
rect 1883 230 1889 231
rect 1126 226 1132 227
rect 1896 226 1898 232
rect 1902 231 1903 235
rect 1907 234 1908 235
rect 1979 235 1985 236
rect 1979 234 1980 235
rect 1907 232 1980 234
rect 1907 231 1908 232
rect 1902 230 1908 231
rect 1979 231 1980 232
rect 1984 231 1985 235
rect 1979 230 1985 231
rect 1998 235 2004 236
rect 1998 231 1999 235
rect 2003 234 2004 235
rect 2107 235 2113 236
rect 2107 234 2108 235
rect 2003 232 2108 234
rect 2003 231 2004 232
rect 1998 230 2004 231
rect 2107 231 2108 232
rect 2112 231 2113 235
rect 2107 230 2113 231
rect 2126 235 2132 236
rect 2126 231 2127 235
rect 2131 234 2132 235
rect 2251 235 2257 236
rect 2251 234 2252 235
rect 2131 232 2252 234
rect 2131 231 2132 232
rect 2126 230 2132 231
rect 2251 231 2252 232
rect 2256 231 2257 235
rect 2251 230 2257 231
rect 2270 235 2276 236
rect 2270 231 2271 235
rect 2275 234 2276 235
rect 2403 235 2409 236
rect 2403 234 2404 235
rect 2275 232 2404 234
rect 2275 231 2276 232
rect 2270 230 2276 231
rect 2403 231 2404 232
rect 2408 231 2409 235
rect 2403 230 2409 231
rect 2563 235 2569 236
rect 2563 231 2564 235
rect 2568 234 2569 235
rect 2590 235 2596 236
rect 2590 234 2591 235
rect 2568 232 2591 234
rect 2568 231 2569 232
rect 2563 230 2569 231
rect 2590 231 2591 232
rect 2595 231 2596 235
rect 2590 230 2596 231
rect 2670 235 2676 236
rect 2670 231 2671 235
rect 2675 234 2676 235
rect 2731 235 2737 236
rect 2731 234 2732 235
rect 2675 232 2732 234
rect 2675 231 2676 232
rect 2670 230 2676 231
rect 2731 231 2732 232
rect 2736 231 2737 235
rect 2731 230 2737 231
rect 2899 235 2905 236
rect 2899 231 2900 235
rect 2904 234 2905 235
rect 2926 235 2932 236
rect 2926 234 2927 235
rect 2904 232 2927 234
rect 2904 231 2905 232
rect 2899 230 2905 231
rect 2926 231 2927 232
rect 2931 231 2932 235
rect 2926 230 2932 231
rect 3075 235 3081 236
rect 3075 231 3076 235
rect 3080 234 3081 235
rect 3126 235 3132 236
rect 3126 234 3127 235
rect 3080 232 3127 234
rect 3080 231 3081 232
rect 3075 230 3081 231
rect 3126 231 3127 232
rect 3131 231 3132 235
rect 3126 230 3132 231
rect 3247 235 3253 236
rect 3247 231 3248 235
rect 3252 234 3253 235
rect 3259 235 3265 236
rect 3259 234 3260 235
rect 3252 232 3260 234
rect 3252 231 3253 232
rect 3247 230 3253 231
rect 3259 231 3260 232
rect 3264 231 3265 235
rect 3259 230 3265 231
rect 3419 235 3425 236
rect 3419 231 3420 235
rect 3424 234 3425 235
rect 3430 235 3436 236
rect 3430 234 3431 235
rect 3424 232 3431 234
rect 3424 231 3425 232
rect 3419 230 3425 231
rect 3430 231 3431 232
rect 3435 231 3436 235
rect 3430 230 3436 231
rect 2238 227 2244 228
rect 2238 226 2239 227
rect 891 225 897 226
rect 219 223 225 224
rect 219 219 220 223
rect 224 222 225 223
rect 230 223 236 224
rect 230 222 231 223
rect 224 220 231 222
rect 224 219 225 220
rect 219 218 225 219
rect 230 219 231 220
rect 235 219 236 223
rect 230 218 236 219
rect 238 223 244 224
rect 238 219 239 223
rect 243 222 244 223
rect 395 223 401 224
rect 395 222 396 223
rect 243 220 396 222
rect 243 219 244 220
rect 238 218 244 219
rect 395 219 396 220
rect 400 219 401 223
rect 395 218 401 219
rect 414 223 420 224
rect 414 219 415 223
rect 419 222 420 223
rect 563 223 569 224
rect 563 222 564 223
rect 419 220 564 222
rect 419 219 420 220
rect 414 218 420 219
rect 563 219 564 220
rect 568 219 569 223
rect 563 218 569 219
rect 582 223 588 224
rect 582 219 583 223
rect 587 222 588 223
rect 731 223 737 224
rect 731 222 732 223
rect 587 220 732 222
rect 587 219 588 220
rect 582 218 588 219
rect 731 219 732 220
rect 736 219 737 223
rect 891 221 892 225
rect 896 221 897 225
rect 1896 224 2239 226
rect 891 220 897 221
rect 910 223 916 224
rect 731 218 737 219
rect 910 219 911 223
rect 915 222 916 223
rect 1043 223 1049 224
rect 1043 222 1044 223
rect 915 220 1044 222
rect 915 219 916 220
rect 910 218 916 219
rect 1043 219 1044 220
rect 1048 219 1049 223
rect 1043 218 1049 219
rect 1062 223 1068 224
rect 1062 219 1063 223
rect 1067 222 1068 223
rect 1187 223 1193 224
rect 1187 222 1188 223
rect 1067 220 1188 222
rect 1067 219 1068 220
rect 1062 218 1068 219
rect 1187 219 1188 220
rect 1192 219 1193 223
rect 1187 218 1193 219
rect 1206 223 1212 224
rect 1206 219 1207 223
rect 1211 222 1212 223
rect 1331 223 1337 224
rect 1331 222 1332 223
rect 1211 220 1332 222
rect 1211 219 1212 220
rect 1206 218 1212 219
rect 1331 219 1332 220
rect 1336 219 1337 223
rect 1331 218 1337 219
rect 1350 223 1356 224
rect 1350 219 1351 223
rect 1355 222 1356 223
rect 1483 223 1489 224
rect 1483 222 1484 223
rect 1355 220 1484 222
rect 1355 219 1356 220
rect 1350 218 1356 219
rect 1483 219 1484 220
rect 1488 219 1489 223
rect 2238 223 2239 224
rect 2243 223 2244 227
rect 2238 222 2244 223
rect 1483 218 1489 219
rect 1830 220 1836 221
rect 1806 217 1812 218
rect 1806 213 1807 217
rect 1811 213 1812 217
rect 1830 216 1831 220
rect 1835 216 1836 220
rect 1830 215 1836 216
rect 1926 220 1932 221
rect 1926 216 1927 220
rect 1931 216 1932 220
rect 1926 215 1932 216
rect 2054 220 2060 221
rect 2054 216 2055 220
rect 2059 216 2060 220
rect 2054 215 2060 216
rect 2198 220 2204 221
rect 2198 216 2199 220
rect 2203 216 2204 220
rect 2198 215 2204 216
rect 2350 220 2356 221
rect 2350 216 2351 220
rect 2355 216 2356 220
rect 2350 215 2356 216
rect 2510 220 2516 221
rect 2510 216 2511 220
rect 2515 216 2516 220
rect 2510 215 2516 216
rect 2678 220 2684 221
rect 2678 216 2679 220
rect 2683 216 2684 220
rect 2678 215 2684 216
rect 2846 220 2852 221
rect 2846 216 2847 220
rect 2851 216 2852 220
rect 2846 215 2852 216
rect 3022 220 3028 221
rect 3022 216 3023 220
rect 3027 216 3028 220
rect 3022 215 3028 216
rect 3206 220 3212 221
rect 3206 216 3207 220
rect 3211 216 3212 220
rect 3206 215 3212 216
rect 3366 220 3372 221
rect 3366 216 3367 220
rect 3371 216 3372 220
rect 3366 215 3372 216
rect 3462 217 3468 218
rect 1806 212 1812 213
rect 3462 213 3463 217
rect 3467 213 3468 217
rect 3462 212 3468 213
rect 1902 211 1908 212
rect 166 208 172 209
rect 110 205 116 206
rect 110 201 111 205
rect 115 201 116 205
rect 166 204 167 208
rect 171 204 172 208
rect 166 203 172 204
rect 342 208 348 209
rect 342 204 343 208
rect 347 204 348 208
rect 342 203 348 204
rect 510 208 516 209
rect 510 204 511 208
rect 515 204 516 208
rect 510 203 516 204
rect 678 208 684 209
rect 678 204 679 208
rect 683 204 684 208
rect 678 203 684 204
rect 838 208 844 209
rect 838 204 839 208
rect 843 204 844 208
rect 838 203 844 204
rect 990 208 996 209
rect 990 204 991 208
rect 995 204 996 208
rect 990 203 996 204
rect 1134 208 1140 209
rect 1134 204 1135 208
rect 1139 204 1140 208
rect 1134 203 1140 204
rect 1278 208 1284 209
rect 1278 204 1279 208
rect 1283 204 1284 208
rect 1278 203 1284 204
rect 1430 208 1436 209
rect 1430 204 1431 208
rect 1435 204 1436 208
rect 1902 207 1903 211
rect 1907 207 1908 211
rect 1902 206 1908 207
rect 1998 211 2004 212
rect 1998 207 1999 211
rect 2003 207 2004 211
rect 1998 206 2004 207
rect 2126 211 2132 212
rect 2126 207 2127 211
rect 2131 207 2132 211
rect 2126 206 2132 207
rect 2270 211 2276 212
rect 2270 207 2271 211
rect 2275 207 2276 211
rect 2270 206 2276 207
rect 2322 211 2328 212
rect 2322 207 2323 211
rect 2327 210 2328 211
rect 2454 211 2460 212
rect 2327 208 2393 210
rect 2327 207 2328 208
rect 2322 206 2328 207
rect 2454 207 2455 211
rect 2459 210 2460 211
rect 2590 211 2596 212
rect 2459 208 2553 210
rect 2459 207 2460 208
rect 2454 206 2460 207
rect 2590 207 2591 211
rect 2595 210 2596 211
rect 2814 211 2820 212
rect 2595 208 2721 210
rect 2595 207 2596 208
rect 2590 206 2596 207
rect 2814 207 2815 211
rect 2819 210 2820 211
rect 2926 211 2932 212
rect 2819 208 2889 210
rect 2819 207 2820 208
rect 2814 206 2820 207
rect 2926 207 2927 211
rect 2931 210 2932 211
rect 3270 211 3276 212
rect 2931 208 3065 210
rect 2931 207 2932 208
rect 2926 206 2932 207
rect 3270 207 3271 211
rect 3275 207 3276 211
rect 3270 206 3276 207
rect 3438 211 3444 212
rect 3438 207 3439 211
rect 3443 207 3444 211
rect 3438 206 3444 207
rect 1430 203 1436 204
rect 1766 205 1772 206
rect 110 200 116 201
rect 1766 201 1767 205
rect 1771 201 1772 205
rect 1830 201 1836 202
rect 1766 200 1772 201
rect 1806 200 1812 201
rect 238 199 244 200
rect 238 195 239 199
rect 243 195 244 199
rect 238 194 244 195
rect 414 199 420 200
rect 414 195 415 199
rect 419 195 420 199
rect 414 194 420 195
rect 582 199 588 200
rect 582 195 583 199
rect 587 195 588 199
rect 582 194 588 195
rect 590 199 596 200
rect 590 195 591 199
rect 595 198 596 199
rect 910 199 916 200
rect 595 196 721 198
rect 595 195 596 196
rect 590 194 596 195
rect 910 195 911 199
rect 915 195 916 199
rect 910 194 916 195
rect 1062 199 1068 200
rect 1062 195 1063 199
rect 1067 195 1068 199
rect 1062 194 1068 195
rect 1206 199 1212 200
rect 1206 195 1207 199
rect 1211 195 1212 199
rect 1206 194 1212 195
rect 1350 199 1356 200
rect 1350 195 1351 199
rect 1355 195 1356 199
rect 1350 194 1356 195
rect 1398 199 1404 200
rect 1398 195 1399 199
rect 1403 198 1404 199
rect 1403 196 1473 198
rect 1806 196 1807 200
rect 1811 196 1812 200
rect 1830 197 1831 201
rect 1835 197 1836 201
rect 1830 196 1836 197
rect 1926 201 1932 202
rect 1926 197 1927 201
rect 1931 197 1932 201
rect 1926 196 1932 197
rect 2054 201 2060 202
rect 2054 197 2055 201
rect 2059 197 2060 201
rect 2054 196 2060 197
rect 2198 201 2204 202
rect 2198 197 2199 201
rect 2203 197 2204 201
rect 2198 196 2204 197
rect 2350 201 2356 202
rect 2350 197 2351 201
rect 2355 197 2356 201
rect 2350 196 2356 197
rect 2510 201 2516 202
rect 2510 197 2511 201
rect 2515 197 2516 201
rect 2510 196 2516 197
rect 2678 201 2684 202
rect 2678 197 2679 201
rect 2683 197 2684 201
rect 2678 196 2684 197
rect 2846 201 2852 202
rect 2846 197 2847 201
rect 2851 197 2852 201
rect 2846 196 2852 197
rect 3022 201 3028 202
rect 3022 197 3023 201
rect 3027 197 3028 201
rect 3022 196 3028 197
rect 3206 201 3212 202
rect 3206 197 3207 201
rect 3211 197 3212 201
rect 3206 196 3212 197
rect 3366 201 3372 202
rect 3366 197 3367 201
rect 3371 197 3372 201
rect 3366 196 3372 197
rect 3462 200 3468 201
rect 3462 196 3463 200
rect 3467 196 3468 200
rect 1403 195 1404 196
rect 1806 195 1812 196
rect 3462 195 3468 196
rect 1398 194 1404 195
rect 166 189 172 190
rect 110 188 116 189
rect 110 184 111 188
rect 115 184 116 188
rect 166 185 167 189
rect 171 185 172 189
rect 166 184 172 185
rect 342 189 348 190
rect 342 185 343 189
rect 347 185 348 189
rect 342 184 348 185
rect 510 189 516 190
rect 510 185 511 189
rect 515 185 516 189
rect 510 184 516 185
rect 678 189 684 190
rect 678 185 679 189
rect 683 185 684 189
rect 678 184 684 185
rect 838 189 844 190
rect 838 185 839 189
rect 843 185 844 189
rect 838 184 844 185
rect 990 189 996 190
rect 990 185 991 189
rect 995 185 996 189
rect 990 184 996 185
rect 1134 189 1140 190
rect 1134 185 1135 189
rect 1139 185 1140 189
rect 1134 184 1140 185
rect 1278 189 1284 190
rect 1278 185 1279 189
rect 1283 185 1284 189
rect 1278 184 1284 185
rect 1430 189 1436 190
rect 1430 185 1431 189
rect 1435 185 1436 189
rect 1430 184 1436 185
rect 1766 188 1772 189
rect 1766 184 1767 188
rect 1771 184 1772 188
rect 110 183 116 184
rect 1766 183 1772 184
rect 1806 136 1812 137
rect 3462 136 3468 137
rect 1806 132 1807 136
rect 1811 132 1812 136
rect 1806 131 1812 132
rect 1830 135 1836 136
rect 1830 131 1831 135
rect 1835 131 1836 135
rect 1830 130 1836 131
rect 1918 135 1924 136
rect 1918 131 1919 135
rect 1923 131 1924 135
rect 1918 130 1924 131
rect 2038 135 2044 136
rect 2038 131 2039 135
rect 2043 131 2044 135
rect 2038 130 2044 131
rect 2158 135 2164 136
rect 2158 131 2159 135
rect 2163 131 2164 135
rect 2158 130 2164 131
rect 2278 135 2284 136
rect 2278 131 2279 135
rect 2283 131 2284 135
rect 2278 130 2284 131
rect 2398 135 2404 136
rect 2398 131 2399 135
rect 2403 131 2404 135
rect 2398 130 2404 131
rect 2510 135 2516 136
rect 2510 131 2511 135
rect 2515 131 2516 135
rect 2510 130 2516 131
rect 2622 135 2628 136
rect 2622 131 2623 135
rect 2627 131 2628 135
rect 2622 130 2628 131
rect 2734 135 2740 136
rect 2734 131 2735 135
rect 2739 131 2740 135
rect 2734 130 2740 131
rect 2838 135 2844 136
rect 2838 131 2839 135
rect 2843 131 2844 135
rect 2838 130 2844 131
rect 2942 135 2948 136
rect 2942 131 2943 135
rect 2947 131 2948 135
rect 2942 130 2948 131
rect 3054 135 3060 136
rect 3054 131 3055 135
rect 3059 131 3060 135
rect 3054 130 3060 131
rect 3166 135 3172 136
rect 3166 131 3167 135
rect 3171 131 3172 135
rect 3166 130 3172 131
rect 3278 135 3284 136
rect 3278 131 3279 135
rect 3283 131 3284 135
rect 3278 130 3284 131
rect 3366 135 3372 136
rect 3366 131 3367 135
rect 3371 131 3372 135
rect 3462 132 3463 136
rect 3467 132 3468 136
rect 3366 130 3372 131
rect 3430 131 3436 132
rect 3462 131 3468 132
rect 2238 127 2244 128
rect 1902 123 1908 124
rect 110 120 116 121
rect 1766 120 1772 121
rect 110 116 111 120
rect 115 116 116 120
rect 110 115 116 116
rect 134 119 140 120
rect 134 115 135 119
rect 139 115 140 119
rect 134 114 140 115
rect 222 119 228 120
rect 222 115 223 119
rect 227 115 228 119
rect 222 114 228 115
rect 310 119 316 120
rect 310 115 311 119
rect 315 115 316 119
rect 310 114 316 115
rect 398 119 404 120
rect 398 115 399 119
rect 403 115 404 119
rect 398 114 404 115
rect 486 119 492 120
rect 486 115 487 119
rect 491 115 492 119
rect 486 114 492 115
rect 574 119 580 120
rect 574 115 575 119
rect 579 115 580 119
rect 574 114 580 115
rect 662 119 668 120
rect 662 115 663 119
rect 667 115 668 119
rect 662 114 668 115
rect 750 119 756 120
rect 750 115 751 119
rect 755 115 756 119
rect 750 114 756 115
rect 846 119 852 120
rect 846 115 847 119
rect 851 115 852 119
rect 846 114 852 115
rect 942 119 948 120
rect 942 115 943 119
rect 947 115 948 119
rect 942 114 948 115
rect 1030 119 1036 120
rect 1030 115 1031 119
rect 1035 115 1036 119
rect 1030 114 1036 115
rect 1118 119 1124 120
rect 1118 115 1119 119
rect 1123 115 1124 119
rect 1118 114 1124 115
rect 1214 119 1220 120
rect 1214 115 1215 119
rect 1219 115 1220 119
rect 1214 114 1220 115
rect 1310 119 1316 120
rect 1310 115 1311 119
rect 1315 115 1316 119
rect 1310 114 1316 115
rect 1406 119 1412 120
rect 1406 115 1407 119
rect 1411 115 1412 119
rect 1406 114 1412 115
rect 1494 119 1500 120
rect 1494 115 1495 119
rect 1499 115 1500 119
rect 1494 114 1500 115
rect 1582 119 1588 120
rect 1582 115 1583 119
rect 1587 115 1588 119
rect 1582 114 1588 115
rect 1670 119 1676 120
rect 1670 115 1671 119
rect 1675 115 1676 119
rect 1766 116 1767 120
rect 1771 116 1772 120
rect 1766 115 1772 116
rect 1806 119 1812 120
rect 1806 115 1807 119
rect 1811 115 1812 119
rect 1902 119 1903 123
rect 1907 119 1908 123
rect 1902 118 1908 119
rect 1990 123 1996 124
rect 1990 119 1991 123
rect 1995 119 1996 123
rect 1990 118 1996 119
rect 2110 123 2116 124
rect 2110 119 2111 123
rect 2115 119 2116 123
rect 2110 118 2116 119
rect 2230 123 2236 124
rect 2230 119 2231 123
rect 2235 119 2236 123
rect 2238 123 2239 127
rect 2243 126 2244 127
rect 3126 127 3132 128
rect 2243 124 2321 126
rect 2243 123 2244 124
rect 2238 122 2244 123
rect 2470 123 2476 124
rect 2230 118 2236 119
rect 2470 119 2471 123
rect 2475 119 2476 123
rect 2470 118 2476 119
rect 2582 123 2588 124
rect 2582 119 2583 123
rect 2587 119 2588 123
rect 2582 118 2588 119
rect 2694 123 2700 124
rect 2694 119 2695 123
rect 2699 119 2700 123
rect 2694 118 2700 119
rect 2806 123 2812 124
rect 2806 119 2807 123
rect 2811 119 2812 123
rect 2806 118 2812 119
rect 2910 123 2916 124
rect 2910 119 2911 123
rect 2915 119 2916 123
rect 2910 118 2916 119
rect 3014 123 3020 124
rect 3014 119 3015 123
rect 3019 119 3020 123
rect 3126 123 3127 127
rect 3131 123 3132 127
rect 3430 127 3431 131
rect 3435 130 3436 131
rect 3435 128 3442 130
rect 3435 127 3436 128
rect 3430 126 3436 127
rect 3440 125 3442 128
rect 3126 122 3132 123
rect 3350 123 3356 124
rect 3241 120 3274 122
rect 3014 118 3020 119
rect 1670 114 1676 115
rect 1806 114 1812 115
rect 1830 116 1836 117
rect 1830 112 1831 116
rect 1835 112 1836 116
rect 742 111 748 112
rect 1830 111 1836 112
rect 1918 116 1924 117
rect 1918 112 1919 116
rect 1923 112 1924 116
rect 1918 111 1924 112
rect 2038 116 2044 117
rect 2038 112 2039 116
rect 2043 112 2044 116
rect 2038 111 2044 112
rect 2158 116 2164 117
rect 2158 112 2159 116
rect 2163 112 2164 116
rect 2158 111 2164 112
rect 2278 116 2284 117
rect 2278 112 2279 116
rect 2283 112 2284 116
rect 2278 111 2284 112
rect 2398 116 2404 117
rect 2398 112 2399 116
rect 2403 112 2404 116
rect 2398 111 2404 112
rect 2510 116 2516 117
rect 2510 112 2511 116
rect 2515 112 2516 116
rect 2510 111 2516 112
rect 2622 116 2628 117
rect 2622 112 2623 116
rect 2627 112 2628 116
rect 2622 111 2628 112
rect 2734 116 2740 117
rect 2734 112 2735 116
rect 2739 112 2740 116
rect 2734 111 2740 112
rect 2838 116 2844 117
rect 2838 112 2839 116
rect 2843 112 2844 116
rect 2838 111 2844 112
rect 2942 116 2948 117
rect 2942 112 2943 116
rect 2947 112 2948 116
rect 2942 111 2948 112
rect 3054 116 3060 117
rect 3054 112 3055 116
rect 3059 112 3060 116
rect 3054 111 3060 112
rect 3166 116 3172 117
rect 3166 112 3167 116
rect 3171 112 3172 116
rect 3166 111 3172 112
rect 206 107 212 108
rect 110 103 116 104
rect 110 99 111 103
rect 115 99 116 103
rect 206 103 207 107
rect 211 103 212 107
rect 206 102 212 103
rect 294 107 300 108
rect 294 103 295 107
rect 299 103 300 107
rect 294 102 300 103
rect 382 107 388 108
rect 382 103 383 107
rect 387 103 388 107
rect 382 102 388 103
rect 470 107 476 108
rect 470 103 471 107
rect 475 103 476 107
rect 470 102 476 103
rect 558 107 564 108
rect 558 103 559 107
rect 563 103 564 107
rect 558 102 564 103
rect 646 107 652 108
rect 646 103 647 107
rect 651 103 652 107
rect 646 102 652 103
rect 734 107 740 108
rect 734 103 735 107
rect 739 103 740 107
rect 742 107 743 111
rect 747 110 748 111
rect 747 108 793 110
rect 1745 108 1802 110
rect 747 107 748 108
rect 742 106 748 107
rect 918 107 924 108
rect 734 102 740 103
rect 918 103 919 107
rect 923 103 924 107
rect 918 102 924 103
rect 1014 107 1020 108
rect 1014 103 1015 107
rect 1019 103 1020 107
rect 1014 102 1020 103
rect 1102 107 1108 108
rect 1102 103 1103 107
rect 1107 103 1108 107
rect 1102 102 1108 103
rect 1190 107 1196 108
rect 1190 103 1191 107
rect 1195 103 1196 107
rect 1190 102 1196 103
rect 1286 107 1292 108
rect 1286 103 1287 107
rect 1291 103 1292 107
rect 1286 102 1292 103
rect 1382 107 1388 108
rect 1382 103 1383 107
rect 1387 103 1388 107
rect 1382 102 1388 103
rect 1478 107 1484 108
rect 1478 103 1479 107
rect 1483 103 1484 107
rect 1478 102 1484 103
rect 1566 107 1572 108
rect 1566 103 1567 107
rect 1571 103 1572 107
rect 1566 102 1572 103
rect 1654 107 1660 108
rect 1654 103 1655 107
rect 1659 103 1660 107
rect 1800 106 1802 108
rect 3272 106 3274 120
rect 3350 119 3351 123
rect 3355 119 3356 123
rect 3350 118 3356 119
rect 3462 119 3468 120
rect 3278 116 3284 117
rect 3278 112 3279 116
rect 3283 112 3284 116
rect 3278 111 3284 112
rect 3366 116 3372 117
rect 3366 112 3367 116
rect 3371 112 3372 116
rect 3462 115 3463 119
rect 3467 115 3468 119
rect 3462 114 3468 115
rect 3366 111 3372 112
rect 1800 104 1886 106
rect 3272 104 3334 106
rect 1654 102 1660 103
rect 1766 103 1772 104
rect 110 98 116 99
rect 134 100 140 101
rect 134 96 135 100
rect 139 96 140 100
rect 134 95 140 96
rect 222 100 228 101
rect 222 96 223 100
rect 227 96 228 100
rect 222 95 228 96
rect 310 100 316 101
rect 310 96 311 100
rect 315 96 316 100
rect 310 95 316 96
rect 398 100 404 101
rect 398 96 399 100
rect 403 96 404 100
rect 398 95 404 96
rect 486 100 492 101
rect 486 96 487 100
rect 491 96 492 100
rect 486 95 492 96
rect 574 100 580 101
rect 574 96 575 100
rect 579 96 580 100
rect 574 95 580 96
rect 662 100 668 101
rect 662 96 663 100
rect 667 96 668 100
rect 662 95 668 96
rect 750 100 756 101
rect 750 96 751 100
rect 755 96 756 100
rect 750 95 756 96
rect 846 100 852 101
rect 846 96 847 100
rect 851 96 852 100
rect 846 95 852 96
rect 942 100 948 101
rect 942 96 943 100
rect 947 96 948 100
rect 942 95 948 96
rect 1030 100 1036 101
rect 1030 96 1031 100
rect 1035 96 1036 100
rect 1030 95 1036 96
rect 1118 100 1124 101
rect 1118 96 1119 100
rect 1123 96 1124 100
rect 1118 95 1124 96
rect 1214 100 1220 101
rect 1214 96 1215 100
rect 1219 96 1220 100
rect 1214 95 1220 96
rect 1310 100 1316 101
rect 1310 96 1311 100
rect 1315 96 1316 100
rect 1310 95 1316 96
rect 1406 100 1412 101
rect 1406 96 1407 100
rect 1411 96 1412 100
rect 1406 95 1412 96
rect 1494 100 1500 101
rect 1494 96 1495 100
rect 1499 96 1500 100
rect 1494 95 1500 96
rect 1582 100 1588 101
rect 1582 96 1583 100
rect 1587 96 1588 100
rect 1582 95 1588 96
rect 1670 100 1676 101
rect 1670 96 1671 100
rect 1675 96 1676 100
rect 1766 99 1767 103
rect 1771 99 1772 103
rect 1884 102 1886 104
rect 3332 102 3334 104
rect 1766 98 1772 99
rect 1883 101 1889 102
rect 1883 97 1884 101
rect 1888 97 1889 101
rect 3331 101 3337 102
rect 1883 96 1889 97
rect 1902 99 1908 100
rect 1670 95 1676 96
rect 1902 95 1903 99
rect 1907 98 1908 99
rect 1971 99 1977 100
rect 1971 98 1972 99
rect 1907 96 1972 98
rect 1907 95 1908 96
rect 1902 94 1908 95
rect 1971 95 1972 96
rect 1976 95 1977 99
rect 1971 94 1977 95
rect 1990 99 1996 100
rect 1990 95 1991 99
rect 1995 98 1996 99
rect 2091 99 2097 100
rect 2091 98 2092 99
rect 1995 96 2092 98
rect 1995 95 1996 96
rect 1990 94 1996 95
rect 2091 95 2092 96
rect 2096 95 2097 99
rect 2091 94 2097 95
rect 2110 99 2116 100
rect 2110 95 2111 99
rect 2115 98 2116 99
rect 2211 99 2217 100
rect 2211 98 2212 99
rect 2115 96 2212 98
rect 2115 95 2116 96
rect 2110 94 2116 95
rect 2211 95 2212 96
rect 2216 95 2217 99
rect 2211 94 2217 95
rect 2230 99 2236 100
rect 2230 95 2231 99
rect 2235 98 2236 99
rect 2331 99 2337 100
rect 2331 98 2332 99
rect 2235 96 2332 98
rect 2235 95 2236 96
rect 2230 94 2236 95
rect 2331 95 2332 96
rect 2336 95 2337 99
rect 2331 94 2337 95
rect 2451 99 2460 100
rect 2451 95 2452 99
rect 2459 95 2460 99
rect 2451 94 2460 95
rect 2470 99 2476 100
rect 2470 95 2471 99
rect 2475 98 2476 99
rect 2563 99 2569 100
rect 2563 98 2564 99
rect 2475 96 2564 98
rect 2475 95 2476 96
rect 2470 94 2476 95
rect 2563 95 2564 96
rect 2568 95 2569 99
rect 2563 94 2569 95
rect 2582 99 2588 100
rect 2582 95 2583 99
rect 2587 98 2588 99
rect 2675 99 2681 100
rect 2675 98 2676 99
rect 2587 96 2676 98
rect 2587 95 2588 96
rect 2582 94 2588 95
rect 2675 95 2676 96
rect 2680 95 2681 99
rect 2675 94 2681 95
rect 2694 99 2700 100
rect 2694 95 2695 99
rect 2699 98 2700 99
rect 2787 99 2793 100
rect 2787 98 2788 99
rect 2699 96 2788 98
rect 2699 95 2700 96
rect 2694 94 2700 95
rect 2787 95 2788 96
rect 2792 95 2793 99
rect 2787 94 2793 95
rect 2806 99 2812 100
rect 2806 95 2807 99
rect 2811 98 2812 99
rect 2891 99 2897 100
rect 2891 98 2892 99
rect 2811 96 2892 98
rect 2811 95 2812 96
rect 2806 94 2812 95
rect 2891 95 2892 96
rect 2896 95 2897 99
rect 2891 94 2897 95
rect 2910 99 2916 100
rect 2910 95 2911 99
rect 2915 98 2916 99
rect 2995 99 3001 100
rect 2995 98 2996 99
rect 2915 96 2996 98
rect 2915 95 2916 96
rect 2910 94 2916 95
rect 2995 95 2996 96
rect 3000 95 3001 99
rect 2995 94 3001 95
rect 3014 99 3020 100
rect 3014 95 3015 99
rect 3019 98 3020 99
rect 3107 99 3113 100
rect 3107 98 3108 99
rect 3019 96 3108 98
rect 3019 95 3020 96
rect 3014 94 3020 95
rect 3107 95 3108 96
rect 3112 95 3113 99
rect 3107 94 3113 95
rect 3219 99 3225 100
rect 3219 95 3220 99
rect 3224 98 3225 99
rect 3270 99 3276 100
rect 3270 98 3271 99
rect 3224 96 3271 98
rect 3224 95 3225 96
rect 3219 94 3225 95
rect 3270 95 3271 96
rect 3275 95 3276 99
rect 3331 97 3332 101
rect 3336 97 3337 101
rect 3331 96 3337 97
rect 3350 99 3356 100
rect 3270 94 3276 95
rect 3350 95 3351 99
rect 3355 98 3356 99
rect 3419 99 3425 100
rect 3419 98 3420 99
rect 3355 96 3420 98
rect 3355 95 3356 96
rect 3350 94 3356 95
rect 3419 95 3420 96
rect 3424 95 3425 99
rect 3419 94 3425 95
rect 206 83 212 84
rect 206 79 207 83
rect 211 82 212 83
rect 275 83 281 84
rect 275 82 276 83
rect 211 80 276 82
rect 211 79 212 80
rect 206 78 212 79
rect 275 79 276 80
rect 280 79 281 83
rect 275 78 281 79
rect 294 83 300 84
rect 294 79 295 83
rect 299 82 300 83
rect 363 83 369 84
rect 363 82 364 83
rect 299 80 364 82
rect 299 79 300 80
rect 294 78 300 79
rect 363 79 364 80
rect 368 79 369 83
rect 363 78 369 79
rect 382 83 388 84
rect 382 79 383 83
rect 387 82 388 83
rect 451 83 457 84
rect 451 82 452 83
rect 387 80 452 82
rect 387 79 388 80
rect 382 78 388 79
rect 451 79 452 80
rect 456 79 457 83
rect 451 78 457 79
rect 470 83 476 84
rect 470 79 471 83
rect 475 82 476 83
rect 539 83 545 84
rect 539 82 540 83
rect 475 80 540 82
rect 475 79 476 80
rect 470 78 476 79
rect 539 79 540 80
rect 544 79 545 83
rect 539 78 545 79
rect 558 83 564 84
rect 558 79 559 83
rect 563 82 564 83
rect 627 83 633 84
rect 627 82 628 83
rect 563 80 628 82
rect 563 79 564 80
rect 558 78 564 79
rect 627 79 628 80
rect 632 79 633 83
rect 627 78 633 79
rect 646 83 652 84
rect 646 79 647 83
rect 651 82 652 83
rect 715 83 721 84
rect 715 82 716 83
rect 651 80 716 82
rect 651 79 652 80
rect 646 78 652 79
rect 715 79 716 80
rect 720 79 721 83
rect 715 78 721 79
rect 734 83 740 84
rect 734 79 735 83
rect 739 82 740 83
rect 803 83 809 84
rect 803 82 804 83
rect 739 80 804 82
rect 739 79 740 80
rect 734 78 740 79
rect 803 79 804 80
rect 808 79 809 83
rect 803 78 809 79
rect 899 83 908 84
rect 899 79 900 83
rect 907 79 908 83
rect 899 78 908 79
rect 918 83 924 84
rect 918 79 919 83
rect 923 82 924 83
rect 995 83 1001 84
rect 995 82 996 83
rect 923 80 996 82
rect 923 79 924 80
rect 918 78 924 79
rect 995 79 996 80
rect 1000 79 1001 83
rect 995 78 1001 79
rect 1014 83 1020 84
rect 1014 79 1015 83
rect 1019 82 1020 83
rect 1083 83 1089 84
rect 1083 82 1084 83
rect 1019 80 1084 82
rect 1019 79 1020 80
rect 1014 78 1020 79
rect 1083 79 1084 80
rect 1088 79 1089 83
rect 1083 78 1089 79
rect 1102 83 1108 84
rect 1102 79 1103 83
rect 1107 82 1108 83
rect 1171 83 1177 84
rect 1171 82 1172 83
rect 1107 80 1172 82
rect 1107 79 1108 80
rect 1102 78 1108 79
rect 1171 79 1172 80
rect 1176 79 1177 83
rect 1171 78 1177 79
rect 1190 83 1196 84
rect 1190 79 1191 83
rect 1195 82 1196 83
rect 1267 83 1273 84
rect 1267 82 1268 83
rect 1195 80 1268 82
rect 1195 79 1196 80
rect 1190 78 1196 79
rect 1267 79 1268 80
rect 1272 79 1273 83
rect 1267 78 1273 79
rect 1286 83 1292 84
rect 1286 79 1287 83
rect 1291 82 1292 83
rect 1363 83 1369 84
rect 1363 82 1364 83
rect 1291 80 1364 82
rect 1291 79 1292 80
rect 1286 78 1292 79
rect 1363 79 1364 80
rect 1368 79 1369 83
rect 1363 78 1369 79
rect 1382 83 1388 84
rect 1382 79 1383 83
rect 1387 82 1388 83
rect 1459 83 1465 84
rect 1459 82 1460 83
rect 1387 80 1460 82
rect 1387 79 1388 80
rect 1382 78 1388 79
rect 1459 79 1460 80
rect 1464 79 1465 83
rect 1459 78 1465 79
rect 1478 83 1484 84
rect 1478 79 1479 83
rect 1483 82 1484 83
rect 1547 83 1553 84
rect 1547 82 1548 83
rect 1483 80 1548 82
rect 1483 79 1484 80
rect 1478 78 1484 79
rect 1547 79 1548 80
rect 1552 79 1553 83
rect 1547 78 1553 79
rect 1566 83 1572 84
rect 1566 79 1567 83
rect 1571 82 1572 83
rect 1635 83 1641 84
rect 1635 82 1636 83
rect 1571 80 1636 82
rect 1571 79 1572 80
rect 1566 78 1572 79
rect 1635 79 1636 80
rect 1640 79 1641 83
rect 1635 78 1641 79
rect 1654 83 1660 84
rect 1654 79 1655 83
rect 1659 82 1660 83
rect 1723 83 1729 84
rect 1723 82 1724 83
rect 1659 80 1724 82
rect 1659 79 1660 80
rect 1654 78 1660 79
rect 1723 79 1724 80
rect 1728 79 1729 83
rect 1723 78 1729 79
<< m3c >>
rect 1807 3496 1811 3500
rect 2007 3495 2011 3499
rect 2239 3495 2243 3499
rect 2455 3495 2459 3499
rect 2655 3495 2659 3499
rect 2855 3495 2859 3499
rect 3047 3495 3051 3499
rect 3247 3495 3251 3499
rect 3463 3496 3467 3500
rect 1807 3479 1811 3483
rect 2311 3483 2315 3487
rect 2407 3487 2411 3491
rect 2727 3483 2731 3487
rect 2927 3483 2931 3487
rect 3119 3483 3123 3487
rect 2007 3476 2011 3480
rect 2239 3476 2243 3480
rect 2455 3476 2459 3480
rect 2655 3476 2659 3480
rect 2855 3476 2859 3480
rect 3047 3476 3051 3480
rect 3247 3476 3251 3480
rect 3463 3479 3467 3483
rect 111 3460 115 3464
rect 455 3459 459 3463
rect 543 3459 547 3463
rect 631 3459 635 3463
rect 719 3459 723 3463
rect 807 3459 811 3463
rect 895 3459 899 3463
rect 983 3459 987 3463
rect 1071 3459 1075 3463
rect 1159 3459 1163 3463
rect 1767 3460 1771 3464
rect 2015 3459 2019 3463
rect 2311 3459 2315 3463
rect 2727 3459 2731 3463
rect 2927 3459 2931 3463
rect 3119 3459 3123 3463
rect 111 3443 115 3447
rect 527 3447 531 3451
rect 615 3447 619 3451
rect 623 3451 627 3455
rect 711 3451 715 3455
rect 799 3451 803 3455
rect 887 3451 891 3455
rect 975 3451 979 3455
rect 1143 3447 1147 3451
rect 1151 3451 1155 3455
rect 455 3440 459 3444
rect 543 3440 547 3444
rect 631 3440 635 3444
rect 719 3440 723 3444
rect 807 3440 811 3444
rect 895 3440 899 3444
rect 983 3440 987 3444
rect 1071 3440 1075 3444
rect 1159 3440 1163 3444
rect 1767 3443 1771 3447
rect 1903 3447 1907 3451
rect 2167 3447 2171 3451
rect 2407 3447 2408 3451
rect 2408 3447 2411 3451
rect 2591 3447 2595 3451
rect 2671 3447 2675 3451
rect 2791 3447 2795 3451
rect 2919 3447 2923 3451
rect 623 3431 627 3435
rect 1151 3431 1155 3435
rect 527 3423 531 3427
rect 711 3423 715 3427
rect 799 3423 803 3427
rect 887 3423 891 3427
rect 975 3423 979 3427
rect 1807 3429 1811 3433
rect 1831 3432 1835 3436
rect 1943 3432 1947 3436
rect 1103 3423 1107 3427
rect 1143 3423 1147 3427
rect 1903 3423 1907 3427
rect 2015 3423 2019 3427
rect 2079 3432 2083 3436
rect 2215 3432 2219 3436
rect 2351 3432 2355 3436
rect 2479 3432 2483 3436
rect 2287 3423 2291 3427
rect 2599 3432 2603 3436
rect 2719 3432 2723 3436
rect 2847 3432 2851 3436
rect 2975 3432 2979 3436
rect 3463 3429 3467 3433
rect 2671 3423 2675 3427
rect 2791 3423 2795 3427
rect 2919 3423 2923 3427
rect 495 3411 499 3415
rect 615 3411 619 3415
rect 663 3411 667 3415
rect 751 3411 755 3415
rect 927 3411 931 3415
rect 1015 3411 1019 3415
rect 1259 3411 1260 3415
rect 1260 3411 1263 3415
rect 1279 3411 1283 3415
rect 1807 3412 1811 3416
rect 1831 3413 1835 3417
rect 1943 3413 1947 3417
rect 2079 3413 2083 3417
rect 2215 3413 2219 3417
rect 2351 3413 2355 3417
rect 2479 3413 2483 3417
rect 2599 3413 2603 3417
rect 2719 3413 2723 3417
rect 2847 3413 2851 3417
rect 2975 3413 2979 3417
rect 3463 3412 3467 3416
rect 111 3393 115 3397
rect 415 3396 419 3400
rect 503 3396 507 3400
rect 591 3396 595 3400
rect 679 3396 683 3400
rect 479 3387 483 3391
rect 495 3387 499 3391
rect 663 3387 667 3391
rect 751 3387 755 3391
rect 767 3396 771 3400
rect 855 3396 859 3400
rect 943 3396 947 3400
rect 1031 3396 1035 3400
rect 927 3387 931 3391
rect 1015 3387 1019 3391
rect 1103 3387 1107 3391
rect 1119 3396 1123 3400
rect 1207 3396 1211 3400
rect 1279 3387 1283 3391
rect 1303 3396 1307 3400
rect 1767 3393 1771 3397
rect 111 3376 115 3380
rect 415 3377 419 3381
rect 503 3377 507 3381
rect 591 3377 595 3381
rect 679 3377 683 3381
rect 767 3377 771 3381
rect 855 3377 859 3381
rect 943 3377 947 3381
rect 1031 3377 1035 3381
rect 1119 3377 1123 3381
rect 1207 3377 1211 3381
rect 1303 3377 1307 3381
rect 1767 3376 1771 3380
rect 1807 3360 1811 3364
rect 1831 3359 1835 3363
rect 1951 3359 1955 3363
rect 2095 3359 2099 3363
rect 2239 3359 2243 3363
rect 2383 3359 2387 3363
rect 2519 3359 2523 3363
rect 2647 3359 2651 3363
rect 2775 3359 2779 3363
rect 2903 3359 2907 3363
rect 3039 3359 3043 3363
rect 3463 3360 3467 3364
rect 1191 3343 1195 3347
rect 1259 3343 1263 3347
rect 1807 3343 1811 3347
rect 1903 3347 1907 3351
rect 2023 3347 2027 3351
rect 2167 3351 2171 3355
rect 2311 3347 2315 3351
rect 2455 3347 2459 3351
rect 2591 3351 2595 3355
rect 2599 3351 2603 3355
rect 2727 3351 2731 3355
rect 2975 3347 2979 3351
rect 2983 3351 2987 3355
rect 1831 3340 1835 3344
rect 1951 3340 1955 3344
rect 2095 3340 2099 3344
rect 2239 3340 2243 3344
rect 2383 3340 2387 3344
rect 2519 3340 2523 3344
rect 2647 3340 2651 3344
rect 2775 3340 2779 3344
rect 2903 3340 2907 3344
rect 3039 3340 3043 3344
rect 3463 3343 3467 3347
rect 111 3328 115 3332
rect 399 3327 403 3331
rect 495 3327 499 3331
rect 599 3327 603 3331
rect 703 3327 707 3331
rect 807 3327 811 3331
rect 911 3327 915 3331
rect 1015 3327 1019 3331
rect 1119 3327 1123 3331
rect 1223 3327 1227 3331
rect 1327 3327 1331 3331
rect 1767 3328 1771 3332
rect 2983 3331 2987 3335
rect 111 3311 115 3315
rect 487 3315 491 3319
rect 567 3315 571 3319
rect 671 3315 675 3319
rect 775 3315 779 3319
rect 879 3315 883 3319
rect 983 3315 987 3319
rect 1087 3315 1091 3319
rect 1191 3319 1195 3323
rect 1199 3319 1203 3323
rect 1303 3319 1307 3323
rect 1895 3323 1899 3327
rect 1903 3323 1907 3327
rect 2023 3323 2027 3327
rect 2287 3323 2291 3327
rect 2311 3323 2315 3327
rect 2599 3323 2603 3327
rect 2727 3323 2731 3327
rect 2975 3323 2979 3327
rect 399 3308 403 3312
rect 495 3308 499 3312
rect 599 3308 603 3312
rect 703 3308 707 3312
rect 807 3308 811 3312
rect 911 3308 915 3312
rect 1015 3308 1019 3312
rect 1119 3308 1123 3312
rect 1223 3308 1227 3312
rect 1327 3308 1331 3312
rect 1767 3311 1771 3315
rect 1199 3299 1203 3303
rect 1911 3303 1915 3307
rect 2055 3303 2059 3307
rect 2103 3303 2107 3307
rect 2415 3303 2419 3307
rect 2455 3303 2459 3307
rect 2751 3303 2755 3307
rect 3055 3303 3059 3307
rect 3327 3303 3331 3307
rect 3439 3303 3443 3307
rect 479 3291 483 3295
rect 487 3291 491 3295
rect 567 3291 571 3295
rect 671 3291 675 3295
rect 775 3291 779 3295
rect 983 3291 987 3295
rect 1087 3291 1091 3295
rect 1303 3291 1307 3295
rect 1399 3291 1403 3295
rect 1807 3285 1811 3289
rect 1831 3288 1835 3292
rect 1975 3288 1979 3292
rect 2151 3288 2155 3292
rect 2335 3288 2339 3292
rect 2511 3288 2515 3292
rect 2679 3288 2683 3292
rect 2831 3288 2835 3292
rect 455 3275 459 3279
rect 695 3275 699 3279
rect 879 3275 883 3279
rect 999 3275 1003 3279
rect 1039 3275 1043 3279
rect 1159 3275 1163 3279
rect 1279 3275 1283 3279
rect 1895 3279 1899 3283
rect 1911 3279 1915 3283
rect 2055 3279 2059 3283
rect 2303 3279 2307 3283
rect 2415 3279 2419 3283
rect 2751 3279 2755 3283
rect 2975 3288 2979 3292
rect 3111 3288 3115 3292
rect 3247 3288 3251 3292
rect 3367 3288 3371 3292
rect 3463 3285 3467 3289
rect 3055 3279 3059 3283
rect 3327 3279 3331 3283
rect 111 3257 115 3261
rect 383 3260 387 3264
rect 495 3260 499 3264
rect 455 3251 459 3255
rect 567 3251 571 3255
rect 1807 3268 1811 3272
rect 1831 3269 1835 3273
rect 1975 3269 1979 3273
rect 2151 3269 2155 3273
rect 2335 3269 2339 3273
rect 2511 3269 2515 3273
rect 2679 3269 2683 3273
rect 2831 3269 2835 3273
rect 2975 3269 2979 3273
rect 3111 3269 3115 3273
rect 3247 3269 3251 3273
rect 3367 3269 3371 3273
rect 3463 3268 3467 3272
rect 607 3260 611 3264
rect 727 3260 731 3264
rect 847 3260 851 3264
rect 967 3260 971 3264
rect 1087 3260 1091 3264
rect 1207 3260 1211 3264
rect 1335 3260 1339 3264
rect 1767 3257 1771 3261
rect 695 3251 699 3255
rect 1039 3251 1043 3255
rect 1159 3251 1163 3255
rect 1279 3251 1283 3255
rect 1399 3251 1403 3255
rect 111 3240 115 3244
rect 383 3241 387 3245
rect 495 3241 499 3245
rect 607 3241 611 3245
rect 727 3241 731 3245
rect 847 3241 851 3245
rect 967 3241 971 3245
rect 1087 3241 1091 3245
rect 1207 3241 1211 3245
rect 1335 3241 1339 3245
rect 1767 3240 1771 3244
rect 1807 3216 1811 3220
rect 1831 3215 1835 3219
rect 2031 3215 2035 3219
rect 2247 3215 2251 3219
rect 2455 3215 2459 3219
rect 2655 3215 2659 3219
rect 2839 3215 2843 3219
rect 3023 3215 3027 3219
rect 3207 3215 3211 3219
rect 3367 3215 3371 3219
rect 3463 3216 3467 3220
rect 1807 3199 1811 3203
rect 2103 3207 2107 3211
rect 2319 3203 2323 3207
rect 2727 3203 2731 3207
rect 2911 3203 2915 3207
rect 3095 3203 3099 3207
rect 111 3192 115 3196
rect 303 3191 307 3195
rect 423 3191 427 3195
rect 543 3191 547 3195
rect 671 3191 675 3195
rect 799 3191 803 3195
rect 927 3191 931 3195
rect 1055 3191 1059 3195
rect 1175 3191 1179 3195
rect 1303 3191 1307 3195
rect 1431 3191 1435 3195
rect 1767 3192 1771 3196
rect 1831 3196 1835 3200
rect 2031 3196 2035 3200
rect 2247 3196 2251 3200
rect 2455 3196 2459 3200
rect 2655 3196 2659 3200
rect 2839 3196 2843 3200
rect 3023 3196 3027 3200
rect 3063 3191 3067 3195
rect 3439 3207 3443 3211
rect 3207 3196 3211 3200
rect 3367 3196 3371 3200
rect 3463 3199 3467 3203
rect 111 3175 115 3179
rect 375 3179 379 3183
rect 495 3179 499 3183
rect 615 3179 619 3183
rect 743 3179 747 3183
rect 759 3183 763 3187
rect 999 3183 1003 3187
rect 1007 3183 1011 3187
rect 1135 3183 1139 3187
rect 1375 3179 1379 3183
rect 1383 3183 1387 3187
rect 303 3172 307 3176
rect 423 3172 427 3176
rect 543 3172 547 3176
rect 671 3172 675 3176
rect 799 3172 803 3176
rect 927 3172 931 3176
rect 1055 3172 1059 3176
rect 1175 3172 1179 3176
rect 1303 3172 1307 3176
rect 1431 3172 1435 3176
rect 1767 3175 1771 3179
rect 1903 3179 1907 3183
rect 2303 3179 2304 3183
rect 2304 3179 2307 3183
rect 2319 3179 2323 3183
rect 2647 3179 2651 3183
rect 2727 3179 2731 3183
rect 2911 3179 2915 3183
rect 3095 3179 3099 3183
rect 3431 3179 3435 3183
rect 759 3163 763 3167
rect 1383 3163 1387 3167
rect 1919 3167 1923 3171
rect 2111 3167 2115 3171
rect 2255 3167 2259 3171
rect 2815 3167 2819 3171
rect 2975 3167 2979 3171
rect 3063 3167 3064 3171
rect 3064 3167 3067 3171
rect 3079 3167 3083 3171
rect 3351 3167 3355 3171
rect 375 3155 379 3159
rect 567 3155 571 3159
rect 615 3155 619 3159
rect 743 3155 747 3159
rect 1007 3155 1011 3159
rect 1135 3155 1139 3159
rect 1271 3155 1275 3159
rect 1375 3155 1379 3159
rect 1807 3149 1811 3153
rect 1839 3152 1843 3156
rect 2031 3152 2035 3156
rect 2223 3152 2227 3156
rect 2407 3152 2411 3156
rect 2575 3152 2579 3156
rect 2735 3152 2739 3156
rect 2879 3152 2883 3156
rect 3007 3152 3011 3156
rect 3135 3152 3139 3156
rect 3263 3152 3267 3156
rect 3367 3152 3371 3156
rect 3463 3149 3467 3153
rect 1903 3143 1907 3147
rect 1919 3143 1923 3147
rect 2111 3143 2115 3147
rect 2479 3143 2483 3147
rect 2647 3143 2651 3147
rect 2815 3143 2819 3147
rect 3079 3143 3083 3147
rect 3207 3143 3211 3147
rect 3431 3143 3435 3147
rect 247 3131 251 3135
rect 495 3131 499 3135
rect 695 3131 699 3135
rect 991 3131 995 3135
rect 1135 3131 1139 3135
rect 1423 3131 1427 3135
rect 1583 3131 1587 3135
rect 1807 3132 1811 3136
rect 1839 3133 1843 3137
rect 2031 3133 2035 3137
rect 2223 3133 2227 3137
rect 2407 3133 2411 3137
rect 2575 3133 2579 3137
rect 2735 3133 2739 3137
rect 2879 3133 2883 3137
rect 3007 3133 3011 3137
rect 3135 3133 3139 3137
rect 3263 3133 3267 3137
rect 3367 3133 3371 3137
rect 3463 3132 3467 3136
rect 111 3113 115 3117
rect 175 3116 179 3120
rect 319 3116 323 3120
rect 471 3116 475 3120
rect 623 3116 627 3120
rect 247 3107 251 3111
rect 391 3107 395 3111
rect 695 3107 699 3111
rect 775 3116 779 3120
rect 919 3116 923 3120
rect 1063 3116 1067 3120
rect 1199 3116 1203 3120
rect 991 3107 995 3111
rect 1135 3107 1139 3111
rect 1271 3107 1275 3111
rect 1343 3116 1347 3120
rect 1487 3116 1491 3120
rect 1767 3113 1771 3117
rect 1423 3107 1427 3111
rect 111 3096 115 3100
rect 175 3097 179 3101
rect 319 3097 323 3101
rect 471 3097 475 3101
rect 623 3097 627 3101
rect 775 3097 779 3101
rect 919 3097 923 3101
rect 1063 3097 1067 3101
rect 1199 3097 1203 3101
rect 1343 3097 1347 3101
rect 1487 3097 1491 3101
rect 1767 3096 1771 3100
rect 1807 3084 1811 3088
rect 1935 3083 1939 3087
rect 2055 3083 2059 3087
rect 2175 3083 2179 3087
rect 2303 3083 2307 3087
rect 2431 3083 2435 3087
rect 2567 3083 2571 3087
rect 2719 3083 2723 3087
rect 2871 3083 2875 3087
rect 3031 3083 3035 3087
rect 3199 3083 3203 3087
rect 3367 3083 3371 3087
rect 3463 3084 3467 3088
rect 1807 3067 1811 3071
rect 2007 3071 2011 3075
rect 2127 3071 2131 3075
rect 2255 3075 2259 3079
rect 2375 3071 2379 3075
rect 2415 3075 2419 3079
rect 2639 3071 2643 3075
rect 2791 3071 2795 3075
rect 2943 3071 2947 3075
rect 2975 3075 2979 3079
rect 3271 3071 3275 3075
rect 3351 3075 3355 3079
rect 1935 3064 1939 3068
rect 2055 3064 2059 3068
rect 2175 3064 2179 3068
rect 2303 3064 2307 3068
rect 2431 3064 2435 3068
rect 2567 3064 2571 3068
rect 2719 3064 2723 3068
rect 2871 3064 2875 3068
rect 3031 3064 3035 3068
rect 3199 3064 3203 3068
rect 3367 3064 3371 3068
rect 3463 3067 3467 3071
rect 111 3044 115 3048
rect 135 3043 139 3047
rect 263 3043 267 3047
rect 431 3043 435 3047
rect 607 3043 611 3047
rect 791 3043 795 3047
rect 967 3043 971 3047
rect 1143 3043 1147 3047
rect 1327 3043 1331 3047
rect 1511 3043 1515 3047
rect 1767 3044 1771 3048
rect 1991 3047 1992 3051
rect 1992 3047 1995 3051
rect 2007 3047 2011 3051
rect 2127 3047 2131 3051
rect 2415 3047 2419 3051
rect 2479 3047 2483 3051
rect 2639 3047 2643 3051
rect 2791 3047 2795 3051
rect 2943 3047 2947 3051
rect 3207 3047 3211 3051
rect 3271 3047 3275 3051
rect 111 3027 115 3031
rect 207 3031 211 3035
rect 335 3031 339 3035
rect 503 3031 507 3035
rect 679 3031 683 3035
rect 755 3035 759 3039
rect 1039 3031 1043 3035
rect 1215 3031 1219 3035
rect 1399 3031 1403 3035
rect 1583 3035 1587 3039
rect 2823 3039 2827 3043
rect 135 3024 139 3028
rect 263 3024 267 3028
rect 431 3024 435 3028
rect 607 3024 611 3028
rect 791 3024 795 3028
rect 967 3024 971 3028
rect 1143 3024 1147 3028
rect 1327 3024 1331 3028
rect 1511 3024 1515 3028
rect 1767 3027 1771 3031
rect 2135 3027 2139 3031
rect 2199 3027 2203 3031
rect 2375 3027 2379 3031
rect 2511 3027 2515 3031
rect 2615 3027 2619 3031
rect 2751 3027 2755 3031
rect 755 3015 759 3019
rect 207 3007 211 3011
rect 391 3007 395 3011
rect 503 3007 507 3011
rect 679 3007 683 3011
rect 999 3007 1003 3011
rect 1039 3007 1043 3011
rect 1215 3007 1219 3011
rect 1399 3007 1403 3011
rect 1807 3009 1811 3013
rect 2023 3012 2027 3016
rect 2127 3012 2131 3016
rect 1991 3003 1995 3007
rect 2199 3003 2203 3007
rect 2663 3019 2667 3023
rect 2231 3012 2235 3016
rect 2335 3012 2339 3016
rect 2439 3012 2443 3016
rect 2543 3012 2547 3016
rect 2647 3012 2651 3016
rect 2759 3012 2763 3016
rect 3463 3009 3467 3013
rect 2399 3003 2403 3007
rect 2511 3003 2515 3007
rect 2615 3003 2619 3007
rect 2751 3003 2755 3007
rect 2823 3003 2827 3007
rect 335 2991 339 2995
rect 399 2991 403 2995
rect 711 2991 715 2995
rect 1007 2991 1011 2995
rect 1411 2991 1415 2995
rect 1555 2991 1559 2995
rect 1663 2991 1667 2995
rect 1807 2992 1811 2996
rect 2023 2993 2027 2997
rect 2127 2993 2131 2997
rect 2231 2993 2235 2997
rect 2335 2993 2339 2997
rect 2439 2993 2443 2997
rect 2543 2993 2547 2997
rect 2647 2993 2651 2997
rect 2759 2993 2763 2997
rect 3463 2992 3467 2996
rect 111 2973 115 2977
rect 135 2976 139 2980
rect 327 2976 331 2980
rect 535 2976 539 2980
rect 199 2967 203 2971
rect 399 2967 403 2971
rect 711 2967 715 2971
rect 735 2976 739 2980
rect 927 2976 931 2980
rect 1103 2976 1107 2980
rect 1279 2976 1283 2980
rect 1447 2976 1451 2980
rect 1623 2976 1627 2980
rect 1767 2973 1771 2977
rect 999 2967 1003 2971
rect 1007 2967 1011 2971
rect 1411 2967 1415 2971
rect 1555 2967 1559 2971
rect 111 2956 115 2960
rect 135 2957 139 2961
rect 327 2957 331 2961
rect 535 2957 539 2961
rect 735 2957 739 2961
rect 927 2957 931 2961
rect 1103 2957 1107 2961
rect 1279 2957 1283 2961
rect 1447 2957 1451 2961
rect 1623 2957 1627 2961
rect 1767 2956 1771 2960
rect 1807 2948 1811 2952
rect 2055 2947 2059 2951
rect 2135 2947 2139 2951
rect 2143 2947 2147 2951
rect 2231 2947 2235 2951
rect 2319 2947 2323 2951
rect 2407 2947 2411 2951
rect 2495 2947 2499 2951
rect 2583 2947 2587 2951
rect 2671 2947 2675 2951
rect 2759 2947 2763 2951
rect 2847 2947 2851 2951
rect 3463 2948 3467 2952
rect 2135 2939 2139 2943
rect 1807 2931 1811 2935
rect 2303 2935 2307 2939
rect 2391 2935 2395 2939
rect 2479 2935 2483 2939
rect 2567 2935 2571 2939
rect 2655 2935 2659 2939
rect 2663 2939 2667 2943
rect 2751 2939 2755 2943
rect 2839 2939 2843 2943
rect 2055 2928 2059 2932
rect 2143 2928 2147 2932
rect 2231 2928 2235 2932
rect 2319 2928 2323 2932
rect 2407 2928 2411 2932
rect 2495 2928 2499 2932
rect 2583 2928 2587 2932
rect 2671 2928 2675 2932
rect 2759 2928 2763 2932
rect 2847 2928 2851 2932
rect 3463 2931 3467 2935
rect 2751 2919 2755 2923
rect 2135 2911 2139 2915
rect 2255 2911 2259 2915
rect 2399 2911 2403 2915
rect 111 2904 115 2908
rect 135 2903 139 2907
rect 263 2903 267 2907
rect 431 2903 435 2907
rect 607 2903 611 2907
rect 783 2903 787 2907
rect 951 2903 955 2907
rect 1111 2903 1115 2907
rect 1271 2903 1275 2907
rect 1431 2903 1435 2907
rect 1591 2903 1595 2907
rect 1767 2904 1771 2908
rect 2303 2903 2307 2907
rect 2479 2911 2483 2915
rect 2567 2911 2571 2915
rect 2655 2911 2659 2915
rect 2839 2911 2843 2915
rect 2855 2911 2859 2915
rect 111 2887 115 2891
rect 207 2891 211 2895
rect 335 2891 339 2895
rect 503 2891 507 2895
rect 679 2891 683 2895
rect 751 2895 755 2899
rect 1023 2891 1027 2895
rect 1183 2891 1187 2895
rect 1343 2891 1347 2895
rect 1503 2891 1507 2895
rect 1663 2895 1667 2899
rect 135 2884 139 2888
rect 263 2884 267 2888
rect 431 2884 435 2888
rect 607 2884 611 2888
rect 783 2884 787 2888
rect 951 2884 955 2888
rect 1111 2884 1115 2888
rect 1271 2884 1275 2888
rect 1431 2884 1435 2888
rect 1591 2884 1595 2888
rect 1767 2887 1771 2891
rect 2055 2887 2059 2891
rect 2247 2891 2251 2895
rect 2391 2891 2395 2895
rect 2559 2891 2563 2895
rect 2647 2891 2651 2895
rect 2751 2891 2755 2895
rect 1807 2873 1811 2877
rect 2071 2876 2075 2880
rect 2175 2876 2179 2880
rect 2271 2876 2275 2880
rect 2367 2876 2371 2880
rect 2471 2876 2475 2880
rect 2575 2876 2579 2880
rect 2679 2876 2683 2880
rect 2783 2876 2787 2880
rect 3463 2873 3467 2877
rect 199 2867 203 2871
rect 207 2867 211 2871
rect 335 2867 339 2871
rect 503 2867 507 2871
rect 679 2867 683 2871
rect 751 2859 755 2863
rect 1023 2867 1027 2871
rect 1183 2867 1187 2871
rect 1343 2867 1347 2871
rect 1503 2867 1507 2871
rect 2247 2867 2251 2871
rect 2255 2867 2259 2871
rect 2431 2867 2435 2871
rect 2647 2867 2651 2871
rect 2751 2867 2755 2871
rect 2855 2867 2859 2871
rect 1399 2859 1403 2863
rect 1807 2856 1811 2860
rect 2071 2857 2075 2861
rect 2175 2857 2179 2861
rect 2271 2857 2275 2861
rect 2367 2857 2371 2861
rect 2471 2857 2475 2861
rect 2575 2857 2579 2861
rect 2679 2857 2683 2861
rect 2783 2857 2787 2861
rect 3463 2856 3467 2860
rect 207 2851 211 2855
rect 327 2851 331 2855
rect 479 2851 483 2855
rect 639 2851 643 2855
rect 999 2851 1003 2855
rect 1095 2851 1099 2855
rect 1239 2851 1243 2855
rect 1383 2851 1387 2855
rect 1279 2843 1283 2847
rect 111 2833 115 2837
rect 135 2836 139 2840
rect 255 2836 259 2840
rect 407 2836 411 2840
rect 567 2836 571 2840
rect 727 2836 731 2840
rect 879 2836 883 2840
rect 1023 2836 1027 2840
rect 1167 2836 1171 2840
rect 1311 2836 1315 2840
rect 1463 2836 1467 2840
rect 1767 2833 1771 2837
rect 207 2827 211 2831
rect 327 2827 331 2831
rect 479 2827 483 2831
rect 639 2827 643 2831
rect 647 2827 651 2831
rect 999 2827 1003 2831
rect 1095 2827 1099 2831
rect 1239 2827 1243 2831
rect 1383 2827 1387 2831
rect 1399 2827 1403 2831
rect 111 2816 115 2820
rect 135 2817 139 2821
rect 255 2817 259 2821
rect 407 2817 411 2821
rect 567 2817 571 2821
rect 727 2817 731 2821
rect 879 2817 883 2821
rect 1023 2817 1027 2821
rect 1167 2817 1171 2821
rect 1311 2817 1315 2821
rect 1463 2817 1467 2821
rect 1767 2816 1771 2820
rect 1807 2808 1811 2812
rect 1983 2807 1987 2811
rect 2111 2807 2115 2811
rect 2239 2807 2243 2811
rect 2367 2807 2371 2811
rect 2487 2807 2491 2811
rect 2607 2807 2611 2811
rect 2719 2807 2723 2811
rect 2839 2807 2843 2811
rect 2959 2807 2963 2811
rect 3463 2808 3467 2812
rect 2055 2799 2059 2803
rect 2063 2799 2067 2803
rect 2191 2799 2195 2803
rect 1807 2791 1811 2795
rect 2439 2795 2443 2799
rect 2559 2799 2563 2803
rect 2687 2799 2691 2803
rect 2911 2795 2915 2799
rect 2919 2799 2923 2803
rect 1983 2788 1987 2792
rect 2111 2788 2115 2792
rect 2239 2788 2243 2792
rect 2367 2788 2371 2792
rect 2487 2788 2491 2792
rect 2607 2788 2611 2792
rect 2719 2788 2723 2792
rect 2839 2788 2843 2792
rect 2959 2788 2963 2792
rect 3463 2791 3467 2795
rect 2919 2779 2923 2783
rect 2063 2771 2067 2775
rect 2191 2771 2195 2775
rect 2255 2771 2259 2775
rect 2431 2771 2435 2775
rect 2687 2771 2691 2775
rect 2911 2771 2915 2775
rect 111 2764 115 2768
rect 287 2763 291 2767
rect 391 2763 395 2767
rect 503 2763 507 2767
rect 623 2763 627 2767
rect 743 2763 747 2767
rect 855 2763 859 2767
rect 967 2763 971 2767
rect 1079 2763 1083 2767
rect 1199 2763 1203 2767
rect 1319 2763 1323 2767
rect 1767 2764 1771 2768
rect 111 2747 115 2751
rect 359 2751 363 2755
rect 463 2751 467 2755
rect 575 2751 579 2755
rect 695 2751 699 2755
rect 731 2755 735 2759
rect 927 2751 931 2755
rect 1039 2751 1043 2755
rect 1151 2751 1155 2755
rect 1271 2751 1275 2755
rect 1279 2755 1283 2759
rect 1903 2755 1907 2759
rect 1959 2755 1963 2759
rect 2103 2755 2107 2759
rect 2439 2755 2443 2759
rect 2455 2755 2459 2759
rect 287 2744 291 2748
rect 391 2744 395 2748
rect 503 2744 507 2748
rect 623 2744 627 2748
rect 743 2744 747 2748
rect 855 2744 859 2748
rect 967 2744 971 2748
rect 1079 2744 1083 2748
rect 1199 2744 1203 2748
rect 1319 2744 1323 2748
rect 1767 2747 1771 2751
rect 2695 2755 2699 2759
rect 2991 2755 2995 2759
rect 3167 2755 3171 2759
rect 647 2735 651 2739
rect 1807 2737 1811 2741
rect 1887 2740 1891 2744
rect 2031 2740 2035 2744
rect 2183 2740 2187 2744
rect 2335 2740 2339 2744
rect 2479 2740 2483 2744
rect 2623 2740 2627 2744
rect 2767 2740 2771 2744
rect 359 2727 363 2731
rect 463 2727 467 2731
rect 575 2727 579 2731
rect 695 2727 699 2731
rect 731 2719 735 2723
rect 927 2727 931 2731
rect 1039 2727 1043 2731
rect 1151 2727 1155 2731
rect 1271 2727 1275 2731
rect 1959 2731 1963 2735
rect 2103 2731 2107 2735
rect 2255 2731 2259 2735
rect 2455 2731 2459 2735
rect 2543 2731 2547 2735
rect 2695 2731 2699 2735
rect 2911 2740 2915 2744
rect 3055 2740 3059 2744
rect 3463 2737 3467 2741
rect 2991 2731 2995 2735
rect 1175 2719 1179 2723
rect 1807 2720 1811 2724
rect 1887 2721 1891 2725
rect 2031 2721 2035 2725
rect 2183 2721 2187 2725
rect 2335 2721 2339 2725
rect 2479 2721 2483 2725
rect 2623 2721 2627 2725
rect 2767 2721 2771 2725
rect 2911 2721 2915 2725
rect 3055 2721 3059 2725
rect 3463 2720 3467 2724
rect 551 2711 555 2715
rect 639 2711 643 2715
rect 727 2711 731 2715
rect 815 2711 819 2715
rect 991 2711 995 2715
rect 1167 2711 1171 2715
rect 1079 2703 1083 2707
rect 111 2693 115 2697
rect 479 2696 483 2700
rect 567 2696 571 2700
rect 655 2696 659 2700
rect 743 2696 747 2700
rect 831 2696 835 2700
rect 919 2696 923 2700
rect 1007 2696 1011 2700
rect 1095 2696 1099 2700
rect 1183 2696 1187 2700
rect 1767 2693 1771 2697
rect 551 2687 555 2691
rect 639 2687 643 2691
rect 727 2687 731 2691
rect 815 2687 819 2691
rect 903 2687 907 2691
rect 991 2687 995 2691
rect 1167 2687 1171 2691
rect 1175 2687 1179 2691
rect 111 2676 115 2680
rect 479 2677 483 2681
rect 567 2677 571 2681
rect 655 2677 659 2681
rect 743 2677 747 2681
rect 831 2677 835 2681
rect 919 2677 923 2681
rect 1007 2677 1011 2681
rect 1095 2677 1099 2681
rect 1183 2677 1187 2681
rect 1767 2676 1771 2680
rect 1807 2676 1811 2680
rect 1831 2675 1835 2679
rect 2023 2675 2027 2679
rect 2231 2675 2235 2679
rect 2431 2675 2435 2679
rect 2615 2675 2619 2679
rect 2783 2675 2787 2679
rect 2943 2675 2947 2679
rect 3095 2675 3099 2679
rect 3239 2675 3243 2679
rect 3367 2675 3371 2679
rect 3463 2676 3467 2680
rect 1903 2667 1907 2671
rect 1911 2667 1915 2671
rect 2103 2667 2107 2671
rect 2415 2667 2419 2671
rect 1807 2659 1811 2663
rect 2687 2663 2691 2667
rect 2855 2663 2859 2667
rect 3015 2663 3019 2667
rect 3167 2667 3171 2671
rect 3311 2663 3315 2667
rect 3319 2667 3323 2671
rect 1831 2656 1835 2660
rect 2023 2656 2027 2660
rect 2231 2656 2235 2660
rect 2431 2656 2435 2660
rect 2615 2656 2619 2660
rect 2783 2656 2787 2660
rect 2943 2656 2947 2660
rect 3095 2656 3099 2660
rect 3239 2656 3243 2660
rect 3367 2656 3371 2660
rect 3463 2659 3467 2663
rect 1911 2639 1915 2643
rect 2103 2639 2107 2643
rect 2255 2639 2259 2643
rect 2543 2639 2547 2643
rect 2591 2639 2595 2643
rect 2687 2639 2691 2643
rect 2855 2639 2859 2643
rect 3015 2639 3019 2643
rect 3319 2639 3323 2643
rect 3431 2639 3435 2643
rect 111 2624 115 2628
rect 471 2623 475 2627
rect 559 2623 563 2627
rect 647 2623 651 2627
rect 735 2623 739 2627
rect 823 2623 827 2627
rect 911 2623 915 2627
rect 999 2623 1003 2627
rect 1087 2623 1091 2627
rect 1767 2624 1771 2628
rect 1799 2623 1803 2627
rect 1903 2623 1907 2627
rect 2071 2623 2075 2627
rect 2415 2623 2416 2627
rect 2416 2623 2419 2627
rect 2915 2623 2919 2627
rect 3035 2623 3039 2627
rect 3151 2623 3155 2627
rect 3311 2623 3315 2627
rect 111 2607 115 2611
rect 543 2611 547 2615
rect 551 2615 555 2619
rect 639 2615 643 2619
rect 727 2615 731 2619
rect 815 2615 819 2619
rect 983 2611 987 2615
rect 1071 2611 1075 2615
rect 1079 2615 1083 2619
rect 2871 2615 2875 2619
rect 471 2604 475 2608
rect 559 2604 563 2608
rect 647 2604 651 2608
rect 735 2604 739 2608
rect 823 2604 827 2608
rect 911 2604 915 2608
rect 999 2604 1003 2608
rect 1087 2604 1091 2608
rect 1767 2607 1771 2611
rect 1807 2605 1811 2609
rect 1831 2608 1835 2612
rect 1999 2608 2003 2612
rect 2183 2608 2187 2612
rect 2359 2608 2363 2612
rect 2519 2608 2523 2612
rect 2671 2608 2675 2612
rect 2807 2608 2811 2612
rect 2927 2608 2931 2612
rect 3047 2608 3051 2612
rect 3159 2608 3163 2612
rect 3271 2608 3275 2612
rect 3367 2608 3371 2612
rect 3463 2605 3467 2609
rect 1903 2599 1907 2603
rect 2071 2599 2075 2603
rect 2255 2599 2259 2603
rect 2263 2599 2267 2603
rect 2591 2599 2595 2603
rect 2915 2599 2919 2603
rect 3035 2599 3039 2603
rect 3151 2599 3155 2603
rect 3431 2599 3435 2603
rect 551 2587 555 2591
rect 639 2587 643 2591
rect 727 2587 731 2591
rect 815 2587 819 2591
rect 903 2587 907 2591
rect 839 2579 843 2583
rect 983 2587 987 2591
rect 1071 2587 1075 2591
rect 1807 2588 1811 2592
rect 1831 2589 1835 2593
rect 1999 2589 2003 2593
rect 2183 2589 2187 2593
rect 2359 2589 2363 2593
rect 2519 2589 2523 2593
rect 2671 2589 2675 2593
rect 2807 2589 2811 2593
rect 2927 2589 2931 2593
rect 3047 2589 3051 2593
rect 3159 2589 3163 2593
rect 3271 2589 3275 2593
rect 3367 2589 3371 2593
rect 3463 2588 3467 2592
rect 295 2563 299 2567
rect 543 2563 547 2567
rect 575 2563 579 2567
rect 751 2563 755 2567
rect 111 2545 115 2549
rect 223 2548 227 2552
rect 311 2548 315 2552
rect 295 2539 299 2543
rect 383 2539 387 2543
rect 407 2548 411 2552
rect 503 2548 507 2552
rect 575 2539 579 2543
rect 807 2555 811 2559
rect 927 2563 931 2567
rect 1015 2563 1019 2567
rect 1103 2563 1107 2567
rect 1191 2563 1195 2567
rect 1287 2563 1291 2567
rect 1055 2555 1059 2559
rect 1567 2563 1571 2567
rect 1655 2563 1659 2567
rect 1663 2555 1667 2559
rect 591 2548 595 2552
rect 679 2548 683 2552
rect 767 2548 771 2552
rect 855 2548 859 2552
rect 943 2548 947 2552
rect 1031 2548 1035 2552
rect 1119 2548 1123 2552
rect 1215 2548 1219 2552
rect 1311 2548 1315 2552
rect 1407 2548 1411 2552
rect 1495 2548 1499 2552
rect 1583 2548 1587 2552
rect 1671 2548 1675 2552
rect 1767 2545 1771 2549
rect 751 2539 755 2543
rect 839 2539 843 2543
rect 927 2539 931 2543
rect 1015 2539 1019 2543
rect 1103 2539 1107 2543
rect 1191 2539 1195 2543
rect 1287 2539 1291 2543
rect 1383 2539 1387 2543
rect 1567 2539 1571 2543
rect 1655 2539 1659 2543
rect 1799 2539 1803 2543
rect 1807 2536 1811 2540
rect 2207 2535 2211 2539
rect 2799 2535 2803 2539
rect 3367 2535 3371 2539
rect 3463 2536 3467 2540
rect 111 2528 115 2532
rect 223 2529 227 2533
rect 311 2529 315 2533
rect 407 2529 411 2533
rect 503 2529 507 2533
rect 591 2529 595 2533
rect 679 2529 683 2533
rect 767 2529 771 2533
rect 855 2529 859 2533
rect 943 2529 947 2533
rect 1031 2529 1035 2533
rect 1119 2529 1123 2533
rect 1215 2529 1219 2533
rect 1311 2529 1315 2533
rect 1407 2529 1411 2533
rect 1495 2529 1499 2533
rect 1583 2529 1587 2533
rect 1671 2529 1675 2533
rect 1767 2528 1771 2532
rect 2071 2527 2075 2531
rect 2871 2527 2875 2531
rect 2879 2527 2883 2531
rect 1807 2519 1811 2523
rect 2207 2516 2211 2520
rect 2799 2516 2803 2520
rect 3367 2516 3371 2520
rect 3463 2519 3467 2523
rect 2263 2499 2264 2503
rect 2264 2499 2267 2503
rect 2879 2499 2883 2503
rect 3431 2499 3435 2503
rect 111 2484 115 2488
rect 135 2483 139 2487
rect 247 2483 251 2487
rect 391 2483 395 2487
rect 543 2483 547 2487
rect 695 2483 699 2487
rect 839 2483 843 2487
rect 975 2483 979 2487
rect 1103 2483 1107 2487
rect 1231 2483 1235 2487
rect 1351 2483 1355 2487
rect 1463 2483 1467 2487
rect 1575 2483 1579 2487
rect 1671 2483 1675 2487
rect 1767 2484 1771 2488
rect 111 2467 115 2471
rect 207 2471 211 2475
rect 215 2475 219 2479
rect 463 2471 467 2475
rect 615 2471 619 2475
rect 623 2475 627 2479
rect 807 2475 811 2479
rect 919 2475 923 2479
rect 1055 2475 1059 2479
rect 1183 2475 1187 2479
rect 1311 2475 1315 2479
rect 1535 2471 1539 2475
rect 1647 2471 1651 2475
rect 1663 2475 1667 2479
rect 135 2464 139 2468
rect 247 2464 251 2468
rect 391 2464 395 2468
rect 543 2464 547 2468
rect 695 2464 699 2468
rect 839 2464 843 2468
rect 975 2464 979 2468
rect 1103 2464 1107 2468
rect 1231 2464 1235 2468
rect 1351 2464 1355 2468
rect 1463 2464 1467 2468
rect 1575 2464 1579 2468
rect 1671 2464 1675 2468
rect 1767 2467 1771 2471
rect 2071 2471 2072 2475
rect 2072 2471 2075 2475
rect 2087 2471 2091 2475
rect 2271 2471 2275 2475
rect 2631 2471 2635 2475
rect 2647 2471 2651 2475
rect 2743 2471 2747 2475
rect 2879 2471 2883 2475
rect 2999 2471 3003 2475
rect 3119 2471 3123 2475
rect 3231 2471 3235 2475
rect 3439 2471 3443 2475
rect 623 2455 627 2459
rect 1383 2455 1387 2459
rect 215 2447 219 2451
rect 383 2447 387 2451
rect 463 2447 467 2451
rect 615 2447 619 2451
rect 919 2447 923 2451
rect 1031 2447 1032 2451
rect 1032 2447 1035 2451
rect 1183 2447 1187 2451
rect 1311 2447 1315 2451
rect 1335 2447 1339 2451
rect 1807 2453 1811 2457
rect 2015 2456 2019 2460
rect 2199 2456 2203 2460
rect 2367 2456 2371 2460
rect 2527 2456 2531 2460
rect 2671 2456 2675 2460
rect 2807 2456 2811 2460
rect 2927 2456 2931 2460
rect 3047 2456 3051 2460
rect 3159 2456 3163 2460
rect 3271 2456 3275 2460
rect 3367 2456 3371 2460
rect 3463 2453 3467 2457
rect 1535 2447 1539 2451
rect 1647 2447 1651 2451
rect 2087 2447 2091 2451
rect 2271 2447 2275 2451
rect 2431 2447 2435 2451
rect 2647 2447 2651 2451
rect 2743 2447 2747 2451
rect 2879 2447 2883 2451
rect 2999 2447 3003 2451
rect 3119 2447 3123 2451
rect 3231 2447 3235 2451
rect 3239 2447 3243 2451
rect 3431 2447 3435 2451
rect 1807 2436 1811 2440
rect 2015 2437 2019 2441
rect 2199 2437 2203 2441
rect 2367 2437 2371 2441
rect 2527 2437 2531 2441
rect 2671 2437 2675 2441
rect 2807 2437 2811 2441
rect 2927 2437 2931 2441
rect 3047 2437 3051 2441
rect 3159 2437 3163 2441
rect 3271 2437 3275 2441
rect 3367 2437 3371 2441
rect 3463 2436 3467 2440
rect 207 2419 211 2423
rect 311 2419 315 2423
rect 463 2419 467 2423
rect 623 2419 627 2423
rect 919 2419 923 2423
rect 967 2419 971 2423
rect 1319 2419 1323 2423
rect 1599 2419 1603 2423
rect 111 2401 115 2405
rect 135 2404 139 2408
rect 239 2404 243 2408
rect 391 2404 395 2408
rect 551 2404 555 2408
rect 719 2404 723 2408
rect 895 2404 899 2408
rect 1063 2404 1067 2408
rect 1239 2404 1243 2408
rect 311 2395 315 2399
rect 463 2395 467 2399
rect 623 2395 627 2399
rect 631 2395 635 2399
rect 967 2395 971 2399
rect 1031 2395 1035 2399
rect 1335 2403 1339 2407
rect 1415 2404 1419 2408
rect 1591 2404 1595 2408
rect 1767 2401 1771 2405
rect 1319 2395 1323 2399
rect 111 2384 115 2388
rect 135 2385 139 2389
rect 239 2385 243 2389
rect 391 2385 395 2389
rect 551 2385 555 2389
rect 719 2385 723 2389
rect 895 2385 899 2389
rect 1063 2385 1067 2389
rect 1239 2385 1243 2389
rect 1415 2385 1419 2389
rect 1591 2385 1595 2389
rect 1767 2384 1771 2388
rect 1807 2388 1811 2392
rect 1839 2387 1843 2391
rect 2007 2387 2011 2391
rect 2183 2387 2187 2391
rect 2367 2387 2371 2391
rect 2559 2387 2563 2391
rect 2759 2387 2763 2391
rect 2967 2387 2971 2391
rect 3175 2387 3179 2391
rect 3367 2387 3371 2391
rect 3463 2388 3467 2392
rect 1807 2371 1811 2375
rect 1911 2375 1915 2379
rect 1919 2379 1923 2383
rect 2087 2379 2091 2383
rect 2263 2379 2267 2383
rect 2631 2379 2635 2383
rect 2639 2379 2643 2383
rect 3247 2375 3251 2379
rect 3439 2379 3443 2383
rect 1839 2368 1843 2372
rect 2007 2368 2011 2372
rect 2183 2368 2187 2372
rect 2367 2368 2371 2372
rect 2559 2368 2563 2372
rect 2759 2368 2763 2372
rect 2967 2368 2971 2372
rect 3175 2368 3179 2372
rect 3367 2368 3371 2372
rect 3463 2371 3467 2375
rect 1919 2351 1923 2355
rect 2087 2351 2091 2355
rect 2263 2351 2267 2355
rect 2431 2351 2435 2355
rect 2639 2351 2643 2355
rect 3039 2351 3043 2355
rect 3239 2351 3243 2355
rect 3439 2351 3443 2355
rect 1911 2339 1915 2343
rect 1959 2339 1963 2343
rect 2087 2339 2091 2343
rect 2223 2339 2227 2343
rect 2719 2339 2723 2343
rect 2911 2339 2915 2343
rect 3247 2339 3251 2343
rect 111 2332 115 2336
rect 375 2331 379 2335
rect 479 2331 483 2335
rect 599 2331 603 2335
rect 719 2331 723 2335
rect 847 2331 851 2335
rect 975 2331 979 2335
rect 1103 2331 1107 2335
rect 1239 2331 1243 2335
rect 1375 2331 1379 2335
rect 1511 2331 1515 2335
rect 1767 2332 1771 2336
rect 111 2315 115 2319
rect 447 2319 451 2323
rect 551 2319 555 2323
rect 671 2319 675 2323
rect 695 2323 699 2327
rect 919 2323 923 2327
rect 927 2323 931 2327
rect 1055 2323 1059 2327
rect 1311 2319 1315 2323
rect 1447 2319 1451 2323
rect 1599 2323 1603 2327
rect 1807 2321 1811 2325
rect 1887 2324 1891 2328
rect 2015 2324 2019 2328
rect 2151 2324 2155 2328
rect 2303 2324 2307 2328
rect 2463 2324 2467 2328
rect 2647 2324 2651 2328
rect 2839 2324 2843 2328
rect 3047 2324 3051 2328
rect 3255 2324 3259 2328
rect 3463 2321 3467 2325
rect 375 2312 379 2316
rect 479 2312 483 2316
rect 599 2312 603 2316
rect 719 2312 723 2316
rect 847 2312 851 2316
rect 975 2312 979 2316
rect 1103 2312 1107 2316
rect 1239 2312 1243 2316
rect 1375 2312 1379 2316
rect 1511 2312 1515 2316
rect 1767 2315 1771 2319
rect 1959 2315 1963 2319
rect 2087 2315 2091 2319
rect 2223 2315 2227 2319
rect 2231 2315 2235 2319
rect 2719 2315 2723 2319
rect 2911 2315 2915 2319
rect 3039 2315 3043 2319
rect 3319 2315 3323 2319
rect 631 2303 635 2307
rect 1807 2304 1811 2308
rect 1887 2305 1891 2309
rect 2015 2305 2019 2309
rect 2151 2305 2155 2309
rect 2303 2305 2307 2309
rect 2463 2305 2467 2309
rect 2647 2305 2651 2309
rect 2839 2305 2843 2309
rect 3047 2305 3051 2309
rect 3255 2305 3259 2309
rect 3463 2304 3467 2308
rect 447 2295 451 2299
rect 551 2295 555 2299
rect 671 2295 675 2299
rect 927 2295 931 2299
rect 1055 2295 1059 2299
rect 1151 2295 1155 2299
rect 1263 2295 1267 2299
rect 1311 2295 1315 2299
rect 1447 2295 1451 2299
rect 695 2283 699 2287
rect 647 2275 651 2279
rect 855 2275 859 2279
rect 935 2275 939 2279
rect 1039 2275 1043 2279
rect 111 2257 115 2261
rect 575 2260 579 2264
rect 663 2260 667 2264
rect 759 2260 763 2264
rect 647 2251 651 2255
rect 735 2251 739 2255
rect 863 2260 867 2264
rect 967 2260 971 2264
rect 1079 2260 1083 2264
rect 1191 2260 1195 2264
rect 1303 2260 1307 2264
rect 1415 2260 1419 2264
rect 1767 2257 1771 2261
rect 1807 2256 1811 2260
rect 935 2251 939 2255
rect 1039 2251 1043 2255
rect 1151 2251 1155 2255
rect 1263 2251 1267 2255
rect 2039 2255 2043 2259
rect 2135 2255 2139 2259
rect 2239 2255 2243 2259
rect 2343 2255 2347 2259
rect 2463 2255 2467 2259
rect 2591 2255 2595 2259
rect 2735 2255 2739 2259
rect 2887 2255 2891 2259
rect 3047 2255 3051 2259
rect 3215 2255 3219 2259
rect 3367 2255 3371 2259
rect 3463 2256 3467 2260
rect 111 2240 115 2244
rect 575 2241 579 2245
rect 663 2241 667 2245
rect 759 2241 763 2245
rect 863 2241 867 2245
rect 967 2241 971 2245
rect 1079 2241 1083 2245
rect 1191 2241 1195 2245
rect 1303 2241 1307 2245
rect 1415 2241 1419 2245
rect 1767 2240 1771 2244
rect 1807 2239 1811 2243
rect 2111 2243 2115 2247
rect 2207 2243 2211 2247
rect 2311 2243 2315 2247
rect 2415 2243 2419 2247
rect 2431 2247 2435 2251
rect 2671 2247 2675 2251
rect 2815 2247 2819 2251
rect 2967 2247 2971 2251
rect 3339 2243 3343 2247
rect 3439 2247 3443 2251
rect 2039 2236 2043 2240
rect 2135 2236 2139 2240
rect 2239 2236 2243 2240
rect 2343 2236 2347 2240
rect 2463 2236 2467 2240
rect 2591 2236 2595 2240
rect 2735 2236 2739 2240
rect 2887 2236 2891 2240
rect 3047 2236 3051 2240
rect 3215 2236 3219 2240
rect 3367 2236 3371 2240
rect 3463 2239 3467 2243
rect 2231 2227 2235 2231
rect 2111 2219 2115 2223
rect 2207 2219 2211 2223
rect 2311 2219 2315 2223
rect 2415 2219 2419 2223
rect 2671 2219 2675 2223
rect 2815 2219 2819 2223
rect 2967 2219 2971 2223
rect 3039 2219 3043 2223
rect 3319 2219 3323 2223
rect 3431 2219 3435 2223
rect 2431 2203 2435 2207
rect 111 2196 115 2200
rect 439 2195 443 2199
rect 527 2195 531 2199
rect 615 2195 619 2199
rect 703 2195 707 2199
rect 791 2195 795 2199
rect 855 2191 859 2195
rect 879 2195 883 2199
rect 967 2195 971 2199
rect 1055 2195 1059 2199
rect 1143 2195 1147 2199
rect 1231 2195 1235 2199
rect 1319 2195 1323 2199
rect 1767 2196 1771 2200
rect 2255 2195 2259 2199
rect 2351 2195 2355 2199
rect 2455 2195 2459 2199
rect 2567 2195 2571 2199
rect 111 2179 115 2183
rect 511 2183 515 2187
rect 599 2183 603 2187
rect 687 2183 691 2187
rect 775 2183 779 2187
rect 951 2183 955 2187
rect 1039 2183 1043 2187
rect 1127 2183 1131 2187
rect 1215 2183 1219 2187
rect 1303 2183 1307 2187
rect 2791 2195 2795 2199
rect 2911 2195 2915 2199
rect 3115 2195 3119 2199
rect 3175 2195 3179 2199
rect 3439 2195 3443 2199
rect 439 2176 443 2180
rect 527 2176 531 2180
rect 615 2176 619 2180
rect 703 2176 707 2180
rect 791 2176 795 2180
rect 879 2176 883 2180
rect 967 2176 971 2180
rect 1055 2176 1059 2180
rect 1143 2176 1147 2180
rect 1231 2176 1235 2180
rect 1319 2176 1323 2180
rect 1767 2179 1771 2183
rect 1807 2177 1811 2181
rect 2183 2180 2187 2184
rect 2279 2180 2283 2184
rect 2383 2180 2387 2184
rect 2495 2180 2499 2184
rect 2607 2180 2611 2184
rect 2719 2180 2723 2184
rect 2839 2180 2843 2184
rect 2967 2180 2971 2184
rect 3103 2180 3107 2184
rect 735 2167 739 2171
rect 2255 2171 2259 2175
rect 2351 2171 2355 2175
rect 2455 2171 2459 2175
rect 2567 2171 2571 2175
rect 2679 2171 2683 2175
rect 2791 2171 2795 2175
rect 2911 2171 2915 2175
rect 3039 2171 3043 2175
rect 3175 2171 3179 2175
rect 3247 2180 3251 2184
rect 3367 2180 3371 2184
rect 3463 2177 3467 2181
rect 3431 2171 3435 2175
rect 511 2159 515 2163
rect 599 2159 603 2163
rect 687 2159 691 2163
rect 775 2159 779 2163
rect 951 2159 955 2163
rect 1039 2159 1043 2163
rect 1127 2159 1131 2163
rect 1215 2159 1219 2163
rect 1303 2159 1307 2163
rect 1807 2160 1811 2164
rect 2183 2161 2187 2165
rect 2279 2161 2283 2165
rect 2383 2161 2387 2165
rect 2495 2161 2499 2165
rect 2607 2161 2611 2165
rect 2719 2161 2723 2165
rect 2839 2161 2843 2165
rect 2967 2161 2971 2165
rect 3103 2161 3107 2165
rect 3247 2161 3251 2165
rect 3367 2161 3371 2165
rect 3463 2160 3467 2164
rect 599 2151 603 2155
rect 327 2131 331 2135
rect 375 2131 379 2135
rect 479 2131 483 2135
rect 591 2131 595 2135
rect 823 2131 827 2135
rect 1007 2131 1011 2135
rect 111 2113 115 2117
rect 303 2116 307 2120
rect 407 2116 411 2120
rect 519 2116 523 2120
rect 631 2116 635 2120
rect 743 2116 747 2120
rect 863 2116 867 2120
rect 983 2116 987 2120
rect 1767 2113 1771 2117
rect 375 2107 379 2111
rect 479 2107 483 2111
rect 591 2107 595 2111
rect 599 2107 603 2111
rect 719 2107 723 2111
rect 823 2107 827 2111
rect 1807 2108 1811 2112
rect 2135 2107 2139 2111
rect 2255 2107 2259 2111
rect 2383 2107 2387 2111
rect 2519 2107 2523 2111
rect 2655 2107 2659 2111
rect 2783 2107 2787 2111
rect 2911 2107 2915 2111
rect 3031 2107 3035 2111
rect 3151 2107 3155 2111
rect 3271 2107 3275 2111
rect 3367 2107 3371 2111
rect 3463 2108 3467 2112
rect 111 2096 115 2100
rect 303 2097 307 2101
rect 407 2097 411 2101
rect 519 2097 523 2101
rect 631 2097 635 2101
rect 743 2097 747 2101
rect 863 2097 867 2101
rect 983 2097 987 2101
rect 1767 2096 1771 2100
rect 1807 2091 1811 2095
rect 2207 2095 2211 2099
rect 2215 2099 2219 2103
rect 2335 2099 2339 2103
rect 2463 2099 2467 2103
rect 2599 2099 2603 2103
rect 2855 2095 2859 2099
rect 2983 2095 2987 2099
rect 3115 2099 3119 2103
rect 3123 2099 3127 2103
rect 3231 2099 3235 2103
rect 3359 2099 3363 2103
rect 2135 2088 2139 2092
rect 2255 2088 2259 2092
rect 2383 2088 2387 2092
rect 2519 2088 2523 2092
rect 2655 2088 2659 2092
rect 2783 2088 2787 2092
rect 2911 2088 2915 2092
rect 3031 2088 3035 2092
rect 3151 2088 3155 2092
rect 3271 2088 3275 2092
rect 3367 2088 3371 2092
rect 3463 2091 3467 2095
rect 3123 2079 3127 2083
rect 2215 2071 2219 2075
rect 2335 2071 2339 2075
rect 2463 2071 2467 2075
rect 2599 2071 2603 2075
rect 2679 2071 2683 2075
rect 2855 2071 2859 2075
rect 2983 2071 2987 2075
rect 3231 2071 3235 2075
rect 3327 2071 3328 2075
rect 3328 2071 3331 2075
rect 3339 2071 3343 2075
rect 111 2052 115 2056
rect 255 2051 259 2055
rect 375 2051 379 2055
rect 495 2051 499 2055
rect 615 2051 619 2055
rect 727 2051 731 2055
rect 831 2051 835 2055
rect 935 2051 939 2055
rect 1039 2051 1043 2055
rect 1143 2051 1147 2055
rect 1255 2051 1259 2055
rect 1767 2052 1771 2056
rect 2207 2051 2211 2055
rect 2319 2051 2323 2055
rect 2487 2051 2491 2055
rect 327 2043 331 2047
rect 335 2043 339 2047
rect 455 2043 459 2047
rect 111 2035 115 2039
rect 687 2039 691 2043
rect 799 2039 803 2043
rect 903 2039 907 2043
rect 1007 2043 1011 2047
rect 1015 2043 1019 2047
rect 1119 2043 1123 2047
rect 1223 2043 1227 2047
rect 2799 2051 2803 2055
rect 2943 2051 2947 2055
rect 3079 2051 3083 2055
rect 3207 2051 3211 2055
rect 3431 2051 3435 2055
rect 3111 2043 3115 2047
rect 255 2032 259 2036
rect 375 2032 379 2036
rect 495 2032 499 2036
rect 615 2032 619 2036
rect 727 2032 731 2036
rect 831 2032 835 2036
rect 935 2032 939 2036
rect 1039 2032 1043 2036
rect 1143 2032 1147 2036
rect 1255 2032 1259 2036
rect 1767 2035 1771 2039
rect 1807 2033 1811 2037
rect 2247 2036 2251 2040
rect 2415 2036 2419 2040
rect 2575 2036 2579 2040
rect 2727 2036 2731 2040
rect 2871 2036 2875 2040
rect 3007 2036 3011 2040
rect 3135 2036 3139 2040
rect 3263 2036 3267 2040
rect 3367 2036 3371 2040
rect 3463 2033 3467 2037
rect 719 2023 723 2027
rect 1015 2023 1019 2027
rect 2319 2027 2323 2031
rect 2487 2027 2491 2031
rect 2527 2027 2531 2031
rect 2799 2027 2803 2031
rect 2943 2027 2947 2031
rect 3079 2027 3083 2031
rect 3207 2027 3211 2031
rect 3327 2027 3331 2031
rect 3439 2027 3443 2031
rect 335 2015 339 2019
rect 455 2015 459 2019
rect 551 2015 552 2019
rect 552 2015 555 2019
rect 687 2015 691 2019
rect 903 2015 907 2019
rect 1119 2015 1123 2019
rect 1223 2015 1227 2019
rect 1807 2016 1811 2020
rect 2247 2017 2251 2021
rect 2415 2017 2419 2021
rect 2575 2017 2579 2021
rect 2727 2017 2731 2021
rect 2871 2017 2875 2021
rect 3007 2017 3011 2021
rect 3135 2017 3139 2021
rect 3263 2017 3267 2021
rect 3367 2017 3371 2021
rect 3463 2016 3467 2020
rect 431 2003 435 2007
rect 703 2003 707 2007
rect 799 2003 803 2007
rect 1095 2003 1099 2007
rect 1351 2003 1355 2007
rect 1487 2003 1491 2007
rect 1599 2003 1603 2007
rect 111 1985 115 1989
rect 359 1988 363 1992
rect 487 1988 491 1992
rect 431 1979 435 1983
rect 551 1979 555 1983
rect 623 1988 627 1992
rect 759 1988 763 1992
rect 895 1988 899 1992
rect 1023 1988 1027 1992
rect 1151 1988 1155 1992
rect 967 1979 971 1983
rect 1095 1979 1099 1983
rect 1271 1988 1275 1992
rect 1399 1988 1403 1992
rect 1527 1988 1531 1992
rect 1767 1985 1771 1989
rect 1351 1979 1355 1983
rect 1487 1979 1491 1983
rect 111 1968 115 1972
rect 359 1969 363 1973
rect 487 1969 491 1973
rect 623 1969 627 1973
rect 759 1969 763 1973
rect 895 1969 899 1973
rect 1023 1969 1027 1973
rect 1151 1969 1155 1973
rect 1271 1969 1275 1973
rect 1399 1969 1403 1973
rect 1527 1969 1531 1973
rect 1767 1968 1771 1972
rect 1807 1956 1811 1960
rect 1831 1955 1835 1959
rect 1919 1955 1923 1959
rect 2047 1955 2051 1959
rect 2183 1955 2187 1959
rect 2327 1955 2331 1959
rect 2471 1955 2475 1959
rect 2615 1955 2619 1959
rect 2751 1955 2755 1959
rect 2887 1955 2891 1959
rect 3031 1955 3035 1959
rect 3175 1955 3179 1959
rect 3319 1955 3323 1959
rect 3463 1956 3467 1960
rect 1807 1939 1811 1943
rect 1903 1943 1907 1947
rect 1911 1947 1915 1951
rect 1999 1947 2003 1951
rect 2127 1947 2131 1951
rect 2263 1947 2267 1951
rect 2543 1943 2547 1947
rect 2687 1943 2691 1947
rect 2823 1943 2827 1947
rect 2959 1943 2963 1947
rect 3103 1943 3107 1947
rect 3111 1947 3115 1951
rect 3391 1943 3395 1947
rect 1831 1936 1835 1940
rect 1919 1936 1923 1940
rect 2047 1936 2051 1940
rect 2183 1936 2187 1940
rect 2327 1936 2331 1940
rect 2471 1936 2475 1940
rect 2615 1936 2619 1940
rect 2751 1936 2755 1940
rect 2887 1936 2891 1940
rect 3031 1936 3035 1940
rect 3175 1936 3179 1940
rect 3319 1936 3323 1940
rect 3463 1939 3467 1943
rect 111 1924 115 1928
rect 447 1923 451 1927
rect 575 1923 579 1927
rect 711 1923 715 1927
rect 847 1923 851 1927
rect 983 1923 987 1927
rect 1119 1923 1123 1927
rect 1255 1923 1259 1927
rect 1383 1923 1387 1927
rect 1519 1923 1523 1927
rect 1655 1923 1659 1927
rect 1767 1924 1771 1928
rect 111 1907 115 1911
rect 647 1911 651 1915
rect 703 1915 707 1919
rect 919 1911 923 1915
rect 927 1915 931 1919
rect 1191 1911 1195 1915
rect 1367 1911 1371 1915
rect 1471 1911 1475 1915
rect 1591 1911 1595 1915
rect 1599 1915 1603 1919
rect 1911 1919 1915 1923
rect 1999 1919 2003 1923
rect 2127 1919 2131 1923
rect 2263 1919 2267 1923
rect 2375 1919 2379 1923
rect 2527 1919 2528 1923
rect 2528 1919 2531 1923
rect 447 1904 451 1908
rect 575 1904 579 1908
rect 711 1904 715 1908
rect 847 1904 851 1908
rect 983 1904 987 1908
rect 1119 1904 1123 1908
rect 1255 1904 1259 1908
rect 1383 1904 1387 1908
rect 1519 1904 1523 1908
rect 1655 1904 1659 1908
rect 1767 1907 1771 1911
rect 1903 1911 1907 1915
rect 2687 1919 2691 1923
rect 2823 1919 2827 1923
rect 2959 1919 2963 1923
rect 3103 1919 3107 1923
rect 3359 1919 3363 1923
rect 3167 1911 3171 1915
rect 1911 1903 1915 1907
rect 2095 1903 2096 1907
rect 2096 1903 2099 1907
rect 2111 1903 2115 1907
rect 2239 1903 2243 1907
rect 2543 1903 2547 1907
rect 1407 1895 1411 1899
rect 2687 1903 2691 1907
rect 2863 1903 2867 1907
rect 3055 1903 3059 1907
rect 3447 1903 3451 1907
rect 3079 1895 3083 1899
rect 539 1887 543 1891
rect 647 1887 651 1891
rect 927 1887 931 1891
rect 967 1887 971 1891
rect 1191 1887 1195 1891
rect 1367 1887 1371 1891
rect 1471 1887 1475 1891
rect 1591 1887 1595 1891
rect 1807 1885 1811 1889
rect 1831 1888 1835 1892
rect 1919 1888 1923 1892
rect 2039 1888 2043 1892
rect 2167 1888 2171 1892
rect 2303 1888 2307 1892
rect 2455 1888 2459 1892
rect 2615 1888 2619 1892
rect 2791 1888 2795 1892
rect 2983 1888 2987 1892
rect 3183 1888 3187 1892
rect 3367 1888 3371 1892
rect 3463 1885 3467 1889
rect 647 1875 651 1879
rect 775 1875 779 1879
rect 919 1875 923 1879
rect 1031 1875 1035 1879
rect 1151 1875 1155 1879
rect 1271 1875 1275 1879
rect 1399 1875 1403 1879
rect 1895 1879 1899 1883
rect 1911 1879 1915 1883
rect 2111 1879 2115 1883
rect 2239 1879 2243 1883
rect 2375 1879 2379 1883
rect 2427 1879 2431 1883
rect 2687 1879 2691 1883
rect 2863 1879 2867 1883
rect 3055 1879 3059 1883
rect 3167 1879 3171 1883
rect 3431 1879 3435 1883
rect 1167 1867 1171 1871
rect 1807 1868 1811 1872
rect 1831 1869 1835 1873
rect 1919 1869 1923 1873
rect 2039 1869 2043 1873
rect 2167 1869 2171 1873
rect 2303 1869 2307 1873
rect 2455 1869 2459 1873
rect 2615 1869 2619 1873
rect 2791 1869 2795 1873
rect 2983 1869 2987 1873
rect 3183 1869 3187 1873
rect 3367 1869 3371 1873
rect 3463 1868 3467 1872
rect 111 1857 115 1861
rect 559 1860 563 1864
rect 695 1860 699 1864
rect 831 1860 835 1864
rect 959 1860 963 1864
rect 1079 1860 1083 1864
rect 1199 1860 1203 1864
rect 1327 1860 1331 1864
rect 1455 1860 1459 1864
rect 1767 1857 1771 1861
rect 539 1851 543 1855
rect 647 1851 651 1855
rect 775 1851 779 1855
rect 1031 1851 1035 1855
rect 1151 1851 1155 1855
rect 1271 1851 1275 1855
rect 1399 1851 1403 1855
rect 1407 1851 1411 1855
rect 111 1840 115 1844
rect 559 1841 563 1845
rect 695 1841 699 1845
rect 831 1841 835 1845
rect 959 1841 963 1845
rect 1079 1841 1083 1845
rect 1199 1841 1203 1845
rect 1327 1841 1331 1845
rect 1455 1841 1459 1845
rect 1767 1840 1771 1844
rect 1807 1820 1811 1824
rect 1831 1819 1835 1823
rect 1959 1819 1963 1823
rect 2111 1819 2115 1823
rect 2255 1819 2259 1823
rect 2407 1819 2411 1823
rect 2567 1819 2571 1823
rect 2743 1819 2747 1823
rect 2935 1819 2939 1823
rect 3135 1819 3139 1823
rect 3343 1819 3347 1823
rect 3463 1820 3467 1824
rect 1727 1811 1731 1815
rect 1807 1803 1811 1807
rect 2031 1807 2035 1811
rect 2095 1811 2099 1815
rect 2327 1807 2331 1811
rect 2479 1807 2483 1811
rect 2639 1807 2643 1811
rect 2815 1807 2819 1811
rect 3007 1807 3011 1811
rect 3079 1811 3083 1815
rect 3271 1811 3275 1815
rect 1831 1800 1835 1804
rect 1959 1800 1963 1804
rect 2111 1800 2115 1804
rect 2255 1800 2259 1804
rect 2407 1800 2411 1804
rect 2567 1800 2571 1804
rect 2743 1800 2747 1804
rect 2935 1800 2939 1804
rect 3135 1800 3139 1804
rect 3343 1800 3347 1804
rect 3463 1803 3467 1807
rect 111 1788 115 1792
rect 135 1787 139 1791
rect 223 1787 227 1791
rect 311 1787 315 1791
rect 407 1787 411 1791
rect 527 1787 531 1791
rect 655 1787 659 1791
rect 799 1787 803 1791
rect 943 1787 947 1791
rect 1087 1787 1091 1791
rect 1239 1787 1243 1791
rect 1391 1787 1395 1791
rect 1543 1787 1547 1791
rect 1671 1787 1675 1791
rect 1767 1788 1771 1792
rect 111 1771 115 1775
rect 207 1775 211 1779
rect 295 1775 299 1779
rect 383 1775 387 1779
rect 479 1775 483 1779
rect 599 1775 603 1779
rect 727 1775 731 1779
rect 1015 1775 1019 1779
rect 1159 1775 1163 1779
rect 1167 1779 1171 1783
rect 1367 1779 1371 1783
rect 1623 1779 1627 1783
rect 1895 1783 1899 1787
rect 1951 1783 1955 1787
rect 2031 1783 2035 1787
rect 2427 1783 2431 1787
rect 2463 1783 2464 1787
rect 2464 1783 2467 1787
rect 2479 1783 2483 1787
rect 2639 1783 2643 1787
rect 2815 1783 2819 1787
rect 3007 1783 3011 1787
rect 3391 1783 3395 1787
rect 135 1768 139 1772
rect 223 1768 227 1772
rect 311 1768 315 1772
rect 407 1768 411 1772
rect 527 1768 531 1772
rect 655 1768 659 1772
rect 799 1768 803 1772
rect 943 1768 947 1772
rect 1087 1768 1091 1772
rect 1239 1768 1243 1772
rect 1391 1768 1395 1772
rect 1543 1768 1547 1772
rect 1671 1768 1675 1772
rect 1767 1771 1771 1775
rect 2799 1767 2803 1771
rect 2095 1759 2099 1763
rect 199 1751 203 1755
rect 207 1751 211 1755
rect 295 1751 299 1755
rect 383 1751 387 1755
rect 479 1751 483 1755
rect 599 1751 603 1755
rect 727 1751 731 1755
rect 999 1751 1000 1755
rect 1000 1751 1003 1755
rect 1015 1751 1019 1755
rect 1159 1751 1163 1755
rect 1623 1751 1627 1755
rect 1727 1751 1728 1755
rect 1728 1751 1731 1755
rect 2255 1755 2259 1759
rect 2327 1759 2331 1763
rect 2559 1759 2563 1763
rect 2983 1759 2987 1763
rect 3431 1759 3435 1763
rect 1807 1741 1811 1745
rect 1879 1744 1883 1748
rect 2015 1744 2019 1748
rect 2151 1744 2155 1748
rect 2303 1744 2307 1748
rect 2479 1744 2483 1748
rect 2687 1744 2691 1748
rect 2911 1744 2915 1748
rect 1951 1735 1955 1739
rect 2095 1735 2099 1739
rect 2367 1735 2371 1739
rect 2463 1735 2467 1739
rect 2559 1735 2563 1739
rect 2983 1735 2987 1739
rect 3151 1744 3155 1748
rect 3367 1744 3371 1748
rect 3463 1741 3467 1745
rect 3447 1735 3451 1739
rect 215 1727 219 1731
rect 327 1727 331 1731
rect 479 1727 483 1731
rect 735 1727 739 1731
rect 1015 1727 1019 1731
rect 1175 1727 1176 1731
rect 1176 1727 1179 1731
rect 1367 1727 1368 1731
rect 1368 1727 1371 1731
rect 1383 1727 1387 1731
rect 1575 1727 1579 1731
rect 1807 1724 1811 1728
rect 1879 1725 1883 1729
rect 2015 1725 2019 1729
rect 2151 1725 2155 1729
rect 2303 1725 2307 1729
rect 2479 1725 2483 1729
rect 2687 1725 2691 1729
rect 2911 1725 2915 1729
rect 3151 1725 3155 1729
rect 3367 1725 3371 1729
rect 3463 1724 3467 1728
rect 111 1709 115 1713
rect 135 1712 139 1716
rect 247 1712 251 1716
rect 399 1712 403 1716
rect 567 1712 571 1716
rect 751 1712 755 1716
rect 935 1712 939 1716
rect 1119 1712 1123 1716
rect 1311 1712 1315 1716
rect 1503 1712 1507 1716
rect 1671 1712 1675 1716
rect 1767 1709 1771 1713
rect 199 1703 203 1707
rect 215 1703 219 1707
rect 327 1703 331 1707
rect 723 1703 727 1707
rect 735 1703 739 1707
rect 999 1703 1003 1707
rect 1015 1703 1019 1707
rect 1383 1703 1387 1707
rect 1575 1703 1579 1707
rect 1735 1703 1739 1707
rect 111 1692 115 1696
rect 135 1693 139 1697
rect 247 1693 251 1697
rect 399 1693 403 1697
rect 567 1693 571 1697
rect 751 1693 755 1697
rect 935 1693 939 1697
rect 1119 1693 1123 1697
rect 1311 1693 1315 1697
rect 1503 1693 1507 1697
rect 1671 1693 1675 1697
rect 1767 1692 1771 1696
rect 1807 1672 1811 1676
rect 1831 1671 1835 1675
rect 1935 1671 1939 1675
rect 2063 1671 2067 1675
rect 2183 1671 2187 1675
rect 2311 1671 2315 1675
rect 2439 1671 2443 1675
rect 2575 1671 2579 1675
rect 2727 1671 2731 1675
rect 2887 1671 2891 1675
rect 3047 1671 3051 1675
rect 3215 1671 3219 1675
rect 3367 1671 3371 1675
rect 3463 1672 3467 1676
rect 1807 1655 1811 1659
rect 1903 1659 1907 1663
rect 2007 1659 2011 1663
rect 2135 1659 2139 1663
rect 2255 1663 2259 1667
rect 2383 1659 2387 1663
rect 2511 1659 2515 1663
rect 2647 1659 2651 1663
rect 2799 1663 2803 1667
rect 2807 1663 2811 1667
rect 2967 1663 2971 1667
rect 3187 1663 3191 1667
rect 3431 1667 3435 1671
rect 1831 1652 1835 1656
rect 1935 1652 1939 1656
rect 2063 1652 2067 1656
rect 2183 1652 2187 1656
rect 2311 1652 2315 1656
rect 2439 1652 2443 1656
rect 2575 1652 2579 1656
rect 2727 1652 2731 1656
rect 2887 1652 2891 1656
rect 3047 1652 3051 1656
rect 3215 1652 3219 1656
rect 3367 1652 3371 1656
rect 3463 1655 3467 1659
rect 111 1644 115 1648
rect 191 1643 195 1647
rect 295 1643 299 1647
rect 407 1643 411 1647
rect 535 1643 539 1647
rect 687 1643 691 1647
rect 855 1643 859 1647
rect 1039 1643 1043 1647
rect 1231 1643 1235 1647
rect 1431 1643 1435 1647
rect 1639 1643 1643 1647
rect 1767 1644 1771 1648
rect 2807 1643 2811 1647
rect 111 1627 115 1631
rect 263 1631 267 1635
rect 367 1631 371 1635
rect 479 1635 483 1639
rect 607 1631 611 1635
rect 615 1635 619 1639
rect 927 1631 931 1635
rect 1111 1631 1115 1635
rect 1175 1635 1179 1639
rect 1503 1631 1507 1635
rect 1511 1635 1515 1639
rect 1895 1635 1899 1639
rect 1903 1635 1907 1639
rect 2007 1635 2011 1639
rect 2135 1635 2139 1639
rect 2367 1635 2368 1639
rect 2368 1635 2371 1639
rect 2511 1635 2515 1639
rect 2647 1635 2651 1639
rect 2967 1635 2971 1639
rect 3087 1635 3091 1639
rect 3271 1635 3272 1639
rect 3272 1635 3275 1639
rect 3431 1635 3435 1639
rect 191 1624 195 1628
rect 295 1624 299 1628
rect 407 1624 411 1628
rect 535 1624 539 1628
rect 687 1624 691 1628
rect 855 1624 859 1628
rect 1039 1624 1043 1628
rect 1231 1624 1235 1628
rect 1431 1624 1435 1628
rect 1639 1624 1643 1628
rect 1767 1627 1771 1631
rect 1911 1615 1915 1619
rect 2023 1615 2027 1619
rect 2167 1615 2171 1619
rect 2287 1615 2288 1619
rect 2288 1615 2291 1619
rect 2383 1615 2387 1619
rect 2559 1615 2560 1619
rect 2560 1615 2563 1619
rect 2711 1615 2715 1619
rect 2839 1615 2843 1619
rect 2967 1615 2971 1619
rect 3187 1615 3188 1619
rect 3188 1615 3191 1619
rect 3207 1615 3211 1619
rect 3335 1615 3339 1619
rect 247 1607 248 1611
rect 248 1607 251 1611
rect 263 1607 267 1611
rect 367 1607 371 1611
rect 615 1607 619 1611
rect 723 1607 727 1611
rect 911 1607 912 1611
rect 912 1607 915 1611
rect 927 1607 931 1611
rect 1111 1607 1115 1611
rect 1511 1607 1515 1611
rect 1735 1607 1739 1611
rect 1807 1597 1811 1601
rect 1831 1600 1835 1604
rect 1943 1600 1947 1604
rect 2087 1600 2091 1604
rect 2231 1600 2235 1604
rect 2367 1600 2371 1604
rect 2503 1600 2507 1604
rect 2639 1600 2643 1604
rect 2767 1600 2771 1604
rect 2895 1600 2899 1604
rect 3015 1600 3019 1604
rect 3135 1600 3139 1604
rect 3263 1600 3267 1604
rect 3367 1600 3371 1604
rect 3463 1597 3467 1601
rect 463 1591 467 1595
rect 607 1591 611 1595
rect 615 1591 619 1595
rect 743 1591 747 1595
rect 1191 1591 1195 1595
rect 1503 1591 1507 1595
rect 1511 1591 1515 1595
rect 1895 1591 1899 1595
rect 1911 1591 1915 1595
rect 2023 1591 2027 1595
rect 2167 1591 2171 1595
rect 2439 1591 2443 1595
rect 2711 1591 2715 1595
rect 2839 1591 2843 1595
rect 2967 1591 2971 1595
rect 3087 1591 3091 1595
rect 3207 1591 3211 1595
rect 3335 1591 3339 1595
rect 3431 1591 3435 1595
rect 111 1573 115 1577
rect 327 1576 331 1580
rect 431 1576 435 1580
rect 543 1576 547 1580
rect 671 1576 675 1580
rect 815 1576 819 1580
rect 967 1576 971 1580
rect 1119 1576 1123 1580
rect 1279 1576 1283 1580
rect 1439 1576 1443 1580
rect 247 1567 251 1571
rect 615 1567 619 1571
rect 743 1567 747 1571
rect 807 1567 811 1571
rect 911 1567 915 1571
rect 1363 1567 1367 1571
rect 1511 1567 1515 1571
rect 1607 1576 1611 1580
rect 1807 1580 1811 1584
rect 1831 1581 1835 1585
rect 1943 1581 1947 1585
rect 2087 1581 2091 1585
rect 2231 1581 2235 1585
rect 2367 1581 2371 1585
rect 2503 1581 2507 1585
rect 2639 1581 2643 1585
rect 2767 1581 2771 1585
rect 2895 1581 2899 1585
rect 3015 1581 3019 1585
rect 3135 1581 3139 1585
rect 3263 1581 3267 1585
rect 3367 1581 3371 1585
rect 3463 1580 3467 1584
rect 1767 1573 1771 1577
rect 111 1556 115 1560
rect 327 1557 331 1561
rect 431 1557 435 1561
rect 543 1557 547 1561
rect 671 1557 675 1561
rect 815 1557 819 1561
rect 967 1557 971 1561
rect 1119 1557 1123 1561
rect 1279 1557 1283 1561
rect 1439 1557 1443 1561
rect 1607 1557 1611 1561
rect 1767 1556 1771 1560
rect 1807 1528 1811 1532
rect 1839 1527 1843 1531
rect 1991 1527 1995 1531
rect 2151 1527 2155 1531
rect 2303 1527 2307 1531
rect 2455 1527 2459 1531
rect 2599 1527 2603 1531
rect 2735 1527 2739 1531
rect 2871 1527 2875 1531
rect 3007 1527 3011 1531
rect 3143 1527 3147 1531
rect 3463 1528 3467 1532
rect 111 1508 115 1512
rect 223 1507 227 1511
rect 343 1507 347 1511
rect 471 1507 475 1511
rect 607 1507 611 1511
rect 751 1507 755 1511
rect 895 1507 899 1511
rect 1047 1507 1051 1511
rect 1199 1507 1203 1511
rect 1351 1507 1355 1511
rect 1503 1507 1507 1511
rect 1767 1508 1771 1512
rect 1807 1511 1811 1515
rect 1911 1515 1915 1519
rect 2063 1515 2067 1519
rect 2223 1515 2227 1519
rect 2287 1519 2291 1523
rect 2551 1515 2555 1519
rect 2559 1519 2563 1523
rect 2679 1519 2683 1523
rect 2815 1519 2819 1523
rect 2951 1519 2955 1523
rect 3087 1519 3091 1523
rect 1839 1508 1843 1512
rect 1991 1508 1995 1512
rect 2151 1508 2155 1512
rect 2303 1508 2307 1512
rect 2455 1508 2459 1512
rect 2599 1508 2603 1512
rect 2735 1508 2739 1512
rect 2871 1508 2875 1512
rect 3007 1508 3011 1512
rect 3143 1508 3147 1512
rect 3463 1511 3467 1515
rect 111 1491 115 1495
rect 295 1495 299 1499
rect 415 1495 419 1499
rect 463 1499 467 1503
rect 551 1499 555 1503
rect 967 1495 971 1499
rect 1119 1495 1123 1499
rect 1191 1499 1195 1503
rect 1423 1495 1427 1499
rect 1575 1495 1579 1499
rect 223 1488 227 1492
rect 343 1488 347 1492
rect 471 1488 475 1492
rect 607 1488 611 1492
rect 751 1488 755 1492
rect 895 1488 899 1492
rect 1047 1488 1051 1492
rect 1199 1488 1203 1492
rect 1351 1488 1355 1492
rect 1503 1488 1507 1492
rect 1767 1491 1771 1495
rect 1895 1491 1896 1495
rect 1896 1491 1899 1495
rect 1911 1491 1915 1495
rect 2063 1491 2067 1495
rect 2223 1491 2227 1495
rect 2439 1491 2443 1495
rect 2679 1491 2683 1495
rect 2815 1491 2819 1495
rect 2951 1491 2955 1495
rect 3087 1491 3091 1495
rect 3199 1491 3200 1495
rect 3200 1491 3203 1495
rect 207 1471 211 1475
rect 295 1471 299 1475
rect 415 1471 419 1475
rect 807 1471 808 1475
rect 808 1471 811 1475
rect 967 1471 971 1475
rect 1119 1471 1123 1475
rect 1363 1471 1367 1475
rect 1423 1471 1427 1475
rect 2135 1471 2139 1475
rect 1011 1463 1015 1467
rect 2391 1471 2392 1475
rect 2392 1471 2395 1475
rect 2407 1471 2411 1475
rect 2551 1471 2555 1475
rect 2839 1471 2840 1475
rect 2840 1471 2843 1475
rect 2855 1471 2859 1475
rect 3159 1471 3163 1475
rect 359 1451 360 1455
rect 360 1451 363 1455
rect 551 1451 555 1455
rect 599 1451 603 1455
rect 703 1451 707 1455
rect 975 1451 979 1455
rect 999 1451 1003 1455
rect 1279 1451 1283 1455
rect 1415 1451 1419 1455
rect 1575 1451 1579 1455
rect 1807 1453 1811 1457
rect 1943 1456 1947 1460
rect 2055 1456 2059 1460
rect 2191 1456 2195 1460
rect 2335 1456 2339 1460
rect 1895 1447 1899 1451
rect 2135 1447 2139 1451
rect 2407 1447 2411 1451
rect 2479 1456 2483 1460
rect 2631 1456 2635 1460
rect 2783 1456 2787 1460
rect 2935 1456 2939 1460
rect 3087 1456 3091 1460
rect 3239 1456 3243 1460
rect 3463 1453 3467 1457
rect 2703 1447 2707 1451
rect 2855 1447 2859 1451
rect 3159 1447 3163 1451
rect 3199 1447 3203 1451
rect 111 1433 115 1437
rect 135 1436 139 1440
rect 303 1436 307 1440
rect 471 1436 475 1440
rect 631 1436 635 1440
rect 783 1436 787 1440
rect 927 1436 931 1440
rect 1063 1436 1067 1440
rect 1199 1436 1203 1440
rect 1335 1436 1339 1440
rect 1471 1436 1475 1440
rect 1767 1433 1771 1437
rect 1807 1436 1811 1440
rect 1943 1437 1947 1441
rect 2055 1437 2059 1441
rect 2191 1437 2195 1441
rect 2335 1437 2339 1441
rect 2479 1437 2483 1441
rect 2631 1437 2635 1441
rect 2783 1437 2787 1441
rect 2935 1437 2939 1441
rect 3087 1437 3091 1441
rect 3239 1437 3243 1441
rect 3463 1436 3467 1440
rect 207 1427 211 1431
rect 599 1427 603 1431
rect 703 1427 707 1431
rect 847 1427 851 1431
rect 999 1427 1003 1431
rect 1011 1427 1015 1431
rect 1271 1427 1275 1431
rect 1279 1427 1283 1431
rect 1415 1427 1419 1431
rect 111 1416 115 1420
rect 135 1417 139 1421
rect 303 1417 307 1421
rect 471 1417 475 1421
rect 631 1417 635 1421
rect 783 1417 787 1421
rect 927 1417 931 1421
rect 1063 1417 1067 1421
rect 1199 1417 1203 1421
rect 1335 1417 1339 1421
rect 1471 1417 1475 1421
rect 1767 1416 1771 1420
rect 1807 1384 1811 1388
rect 2095 1383 2099 1387
rect 2199 1383 2203 1387
rect 2319 1383 2323 1387
rect 2455 1383 2459 1387
rect 2599 1383 2603 1387
rect 2743 1383 2747 1387
rect 2887 1383 2891 1387
rect 3031 1383 3035 1387
rect 3175 1383 3179 1387
rect 3327 1383 3331 1387
rect 3463 1384 3467 1388
rect 111 1368 115 1372
rect 135 1367 139 1371
rect 279 1367 283 1371
rect 447 1367 451 1371
rect 607 1367 611 1371
rect 759 1367 763 1371
rect 903 1367 907 1371
rect 1031 1367 1035 1371
rect 1159 1367 1163 1371
rect 1287 1367 1291 1371
rect 1415 1367 1419 1371
rect 1767 1368 1771 1372
rect 1807 1367 1811 1371
rect 2167 1371 2171 1375
rect 2271 1371 2275 1375
rect 2391 1375 2395 1379
rect 2427 1375 2431 1379
rect 2535 1375 2539 1379
rect 2735 1375 2739 1379
rect 2839 1375 2843 1379
rect 2967 1375 2971 1379
rect 3255 1375 3259 1379
rect 2095 1364 2099 1368
rect 111 1351 115 1355
rect 207 1355 211 1359
rect 351 1355 355 1359
rect 359 1359 363 1363
rect 559 1359 563 1363
rect 739 1359 743 1363
rect 975 1359 979 1363
rect 983 1359 987 1363
rect 1111 1359 1115 1363
rect 2199 1364 2203 1368
rect 2319 1364 2323 1368
rect 2455 1364 2459 1368
rect 2599 1364 2603 1368
rect 2743 1364 2747 1368
rect 2887 1364 2891 1368
rect 3031 1364 3035 1368
rect 3175 1364 3179 1368
rect 3327 1364 3331 1368
rect 3463 1367 3467 1371
rect 1359 1355 1363 1359
rect 1367 1359 1371 1363
rect 135 1348 139 1352
rect 279 1348 283 1352
rect 447 1348 451 1352
rect 607 1348 611 1352
rect 759 1348 763 1352
rect 903 1348 907 1352
rect 1031 1348 1035 1352
rect 1159 1348 1163 1352
rect 1287 1348 1291 1352
rect 1415 1348 1419 1352
rect 1767 1351 1771 1355
rect 2427 1355 2431 1359
rect 2167 1347 2171 1351
rect 2271 1347 2275 1351
rect 2535 1347 2539 1351
rect 2607 1347 2611 1351
rect 2703 1347 2707 1351
rect 2967 1347 2971 1351
rect 3255 1347 3259 1351
rect 3375 1347 3379 1351
rect 199 1331 203 1335
rect 207 1331 211 1335
rect 351 1331 355 1335
rect 739 1331 743 1335
rect 847 1331 851 1335
rect 983 1331 987 1335
rect 1111 1331 1115 1335
rect 1255 1331 1259 1335
rect 1271 1331 1275 1335
rect 1359 1331 1363 1335
rect 559 1323 563 1327
rect 2175 1331 2179 1335
rect 2311 1331 2315 1335
rect 2735 1331 2739 1335
rect 2323 1323 2327 1327
rect 2911 1331 2915 1335
rect 3063 1331 3067 1335
rect 3215 1331 3219 1335
rect 3055 1323 3059 1327
rect 207 1315 211 1319
rect 351 1315 355 1319
rect 511 1315 515 1319
rect 687 1315 691 1319
rect 791 1315 795 1319
rect 919 1315 923 1319
rect 1039 1315 1043 1319
rect 1299 1315 1303 1319
rect 1367 1315 1368 1319
rect 1368 1315 1371 1319
rect 1807 1313 1811 1317
rect 2103 1316 2107 1320
rect 2239 1316 2243 1320
rect 2383 1316 2387 1320
rect 2535 1316 2539 1320
rect 2687 1316 2691 1320
rect 2839 1316 2843 1320
rect 2991 1316 2995 1320
rect 3143 1316 3147 1320
rect 3303 1316 3307 1320
rect 3463 1313 3467 1317
rect 2175 1307 2179 1311
rect 2311 1307 2315 1311
rect 2607 1307 2611 1311
rect 2751 1307 2755 1311
rect 2911 1307 2915 1311
rect 3063 1307 3067 1311
rect 3215 1307 3219 1311
rect 3375 1307 3379 1311
rect 111 1297 115 1301
rect 135 1300 139 1304
rect 279 1300 283 1304
rect 439 1300 443 1304
rect 583 1300 587 1304
rect 719 1300 723 1304
rect 847 1300 851 1304
rect 967 1300 971 1304
rect 1079 1300 1083 1304
rect 1191 1300 1195 1304
rect 1311 1300 1315 1304
rect 1767 1297 1771 1301
rect 1807 1296 1811 1300
rect 2103 1297 2107 1301
rect 2239 1297 2243 1301
rect 2383 1297 2387 1301
rect 2535 1297 2539 1301
rect 2687 1297 2691 1301
rect 2839 1297 2843 1301
rect 2991 1297 2995 1301
rect 3143 1297 3147 1301
rect 3303 1297 3307 1301
rect 3463 1296 3467 1300
rect 199 1291 203 1295
rect 351 1291 355 1295
rect 511 1291 515 1295
rect 655 1291 659 1295
rect 791 1291 795 1295
rect 919 1291 923 1295
rect 1039 1291 1043 1295
rect 1047 1291 1051 1295
rect 1255 1291 1259 1295
rect 1299 1291 1303 1295
rect 111 1280 115 1284
rect 135 1281 139 1285
rect 279 1281 283 1285
rect 439 1281 443 1285
rect 583 1281 587 1285
rect 719 1281 723 1285
rect 847 1281 851 1285
rect 967 1281 971 1285
rect 1079 1281 1083 1285
rect 1191 1281 1195 1285
rect 1311 1281 1315 1285
rect 1767 1280 1771 1284
rect 1807 1252 1811 1256
rect 1935 1251 1939 1255
rect 2063 1251 2067 1255
rect 2199 1251 2203 1255
rect 2343 1251 2347 1255
rect 2495 1251 2499 1255
rect 2655 1251 2659 1255
rect 2815 1251 2819 1255
rect 2975 1251 2979 1255
rect 3143 1251 3147 1255
rect 3463 1252 3467 1256
rect 111 1232 115 1236
rect 135 1231 139 1235
rect 239 1231 243 1235
rect 367 1231 371 1235
rect 495 1231 499 1235
rect 615 1231 619 1235
rect 735 1231 739 1235
rect 847 1231 851 1235
rect 959 1231 963 1235
rect 1071 1231 1075 1235
rect 1191 1231 1195 1235
rect 1767 1232 1771 1236
rect 1807 1235 1811 1239
rect 2007 1239 2011 1243
rect 2135 1239 2139 1243
rect 2271 1239 2275 1243
rect 2323 1243 2327 1247
rect 2567 1239 2571 1243
rect 2575 1243 2579 1247
rect 2887 1239 2891 1243
rect 3047 1239 3051 1243
rect 3055 1243 3059 1247
rect 1935 1232 1939 1236
rect 2063 1232 2067 1236
rect 2199 1232 2203 1236
rect 2343 1232 2347 1236
rect 2495 1232 2499 1236
rect 2655 1232 2659 1236
rect 2815 1232 2819 1236
rect 2975 1232 2979 1236
rect 3143 1232 3147 1236
rect 3463 1235 3467 1239
rect 207 1223 211 1227
rect 215 1223 219 1227
rect 319 1223 323 1227
rect 447 1223 451 1227
rect 687 1223 691 1227
rect 111 1215 115 1219
rect 807 1219 811 1223
rect 919 1219 923 1223
rect 1031 1219 1035 1223
rect 1143 1219 1147 1223
rect 1151 1223 1155 1227
rect 2311 1223 2315 1227
rect 135 1212 139 1216
rect 239 1212 243 1216
rect 367 1212 371 1216
rect 495 1212 499 1216
rect 615 1212 619 1216
rect 735 1212 739 1216
rect 847 1212 851 1216
rect 959 1212 963 1216
rect 1071 1212 1075 1216
rect 1191 1212 1195 1216
rect 1767 1215 1771 1219
rect 2007 1215 2011 1219
rect 2135 1215 2139 1219
rect 2271 1215 2275 1219
rect 2575 1215 2579 1219
rect 2751 1215 2755 1219
rect 2767 1215 2771 1219
rect 2887 1215 2891 1219
rect 3047 1215 3051 1219
rect 1047 1203 1051 1207
rect 1927 1203 1931 1207
rect 215 1195 219 1199
rect 319 1195 323 1199
rect 447 1195 451 1199
rect 623 1195 627 1199
rect 655 1195 659 1199
rect 807 1195 811 1199
rect 919 1195 923 1199
rect 1031 1195 1035 1199
rect 1143 1195 1147 1199
rect 2007 1203 2011 1207
rect 2151 1203 2155 1207
rect 2303 1203 2307 1207
rect 2567 1203 2571 1207
rect 2775 1203 2779 1207
rect 2943 1203 2947 1207
rect 3071 1203 3075 1207
rect 1151 1187 1155 1191
rect 183 1179 187 1183
rect 207 1179 211 1183
rect 311 1179 315 1183
rect 447 1179 451 1183
rect 583 1179 587 1183
rect 1807 1185 1811 1189
rect 1831 1188 1835 1192
rect 863 1179 867 1183
rect 999 1179 1003 1183
rect 1135 1179 1139 1183
rect 1271 1179 1275 1183
rect 1935 1188 1939 1192
rect 2079 1188 2083 1192
rect 2231 1188 2235 1192
rect 2391 1188 2395 1192
rect 2543 1188 2547 1192
rect 2695 1188 2699 1192
rect 2847 1188 2851 1192
rect 2999 1188 3003 1192
rect 2007 1179 2011 1183
rect 2151 1179 2155 1183
rect 2303 1179 2307 1183
rect 2311 1179 2315 1183
rect 2607 1179 2611 1183
rect 2767 1179 2771 1183
rect 2775 1179 2779 1183
rect 3071 1179 3075 1183
rect 3159 1188 3163 1192
rect 3463 1185 3467 1189
rect 111 1161 115 1165
rect 135 1164 139 1168
rect 239 1164 243 1168
rect 375 1164 379 1168
rect 511 1164 515 1168
rect 655 1164 659 1168
rect 791 1164 795 1168
rect 927 1164 931 1168
rect 1063 1164 1067 1168
rect 1199 1164 1203 1168
rect 1335 1164 1339 1168
rect 1807 1168 1811 1172
rect 1831 1169 1835 1173
rect 1935 1169 1939 1173
rect 2079 1169 2083 1173
rect 2231 1169 2235 1173
rect 2391 1169 2395 1173
rect 2543 1169 2547 1173
rect 2695 1169 2699 1173
rect 2847 1169 2851 1173
rect 2999 1169 3003 1173
rect 3159 1169 3163 1173
rect 3463 1168 3467 1172
rect 1767 1161 1771 1165
rect 207 1155 211 1159
rect 311 1155 315 1159
rect 447 1155 451 1159
rect 583 1155 587 1159
rect 623 1155 627 1159
rect 863 1155 867 1159
rect 999 1155 1003 1159
rect 1135 1155 1139 1159
rect 1271 1155 1275 1159
rect 1279 1155 1283 1159
rect 111 1144 115 1148
rect 135 1145 139 1149
rect 239 1145 243 1149
rect 375 1145 379 1149
rect 511 1145 515 1149
rect 655 1145 659 1149
rect 791 1145 795 1149
rect 927 1145 931 1149
rect 1063 1145 1067 1149
rect 1199 1145 1203 1149
rect 1335 1145 1339 1149
rect 1767 1144 1771 1148
rect 1807 1112 1811 1116
rect 1863 1111 1867 1115
rect 1927 1107 1931 1111
rect 1983 1111 1987 1115
rect 2111 1111 2115 1115
rect 2247 1111 2251 1115
rect 2383 1111 2387 1115
rect 2511 1111 2515 1115
rect 2639 1111 2643 1115
rect 2759 1111 2763 1115
rect 2871 1111 2875 1115
rect 2975 1111 2979 1115
rect 3079 1111 3083 1115
rect 3183 1111 3187 1115
rect 3279 1111 3283 1115
rect 3367 1111 3371 1115
rect 3463 1112 3467 1116
rect 1943 1103 1947 1107
rect 2063 1103 2067 1107
rect 2191 1103 2195 1107
rect 111 1096 115 1100
rect 191 1095 195 1099
rect 335 1095 339 1099
rect 495 1095 499 1099
rect 655 1095 659 1099
rect 815 1095 819 1099
rect 967 1095 971 1099
rect 1119 1095 1123 1099
rect 1263 1095 1267 1099
rect 1407 1095 1411 1099
rect 1559 1095 1563 1099
rect 1767 1096 1771 1100
rect 1807 1095 1811 1099
rect 2583 1099 2587 1103
rect 2711 1099 2715 1103
rect 2831 1099 2835 1103
rect 2943 1103 2947 1107
rect 2951 1103 2955 1107
rect 3055 1103 3059 1107
rect 3159 1103 3163 1107
rect 3263 1103 3267 1107
rect 1863 1092 1867 1096
rect 183 1087 187 1091
rect 271 1087 275 1091
rect 415 1087 419 1091
rect 111 1079 115 1083
rect 727 1083 731 1087
rect 767 1087 771 1091
rect 1983 1092 1987 1096
rect 2111 1092 2115 1096
rect 2247 1092 2251 1096
rect 2383 1092 2387 1096
rect 2511 1092 2515 1096
rect 2639 1092 2643 1096
rect 2759 1092 2763 1096
rect 2871 1092 2875 1096
rect 2975 1092 2979 1096
rect 3079 1092 3083 1096
rect 3183 1092 3187 1096
rect 3279 1092 3283 1096
rect 3367 1092 3371 1096
rect 3463 1095 3467 1099
rect 1039 1083 1043 1087
rect 1191 1083 1195 1087
rect 1335 1083 1339 1087
rect 1479 1083 1483 1087
rect 191 1076 195 1080
rect 335 1076 339 1080
rect 495 1076 499 1080
rect 655 1076 659 1080
rect 815 1076 819 1080
rect 967 1076 971 1080
rect 1119 1076 1123 1080
rect 1263 1076 1267 1080
rect 1407 1076 1411 1080
rect 1559 1076 1563 1080
rect 1767 1079 1771 1083
rect 2951 1083 2955 1087
rect 1943 1075 1947 1079
rect 2063 1075 2067 1079
rect 2191 1075 2195 1079
rect 2351 1075 2355 1079
rect 2607 1075 2611 1079
rect 2711 1075 2715 1079
rect 2831 1075 2835 1079
rect 3055 1075 3059 1079
rect 3159 1075 3163 1079
rect 3263 1075 3267 1079
rect 3439 1075 3443 1079
rect 767 1067 771 1071
rect 1279 1067 1283 1071
rect 271 1059 275 1063
rect 415 1059 419 1063
rect 679 1059 683 1063
rect 727 1059 731 1063
rect 1039 1059 1043 1063
rect 1191 1059 1195 1063
rect 1335 1059 1339 1063
rect 1479 1059 1483 1063
rect 2175 1063 2179 1067
rect 399 1047 403 1051
rect 2263 1055 2267 1059
rect 2447 1055 2451 1059
rect 2503 1055 2507 1059
rect 2583 1055 2587 1059
rect 2615 1055 2619 1059
rect 2703 1055 2707 1059
rect 2791 1055 2795 1059
rect 535 1039 539 1043
rect 847 1039 851 1043
rect 959 1039 963 1043
rect 1159 1039 1163 1043
rect 1463 1039 1467 1043
rect 1471 1039 1475 1043
rect 1607 1039 1611 1043
rect 1807 1037 1811 1041
rect 2103 1040 2107 1044
rect 2191 1040 2195 1044
rect 2279 1040 2283 1044
rect 111 1021 115 1025
rect 327 1024 331 1028
rect 463 1024 467 1028
rect 607 1024 611 1028
rect 399 1015 403 1019
rect 535 1015 539 1019
rect 679 1015 683 1019
rect 2175 1031 2179 1035
rect 2263 1031 2267 1035
rect 2351 1031 2355 1035
rect 2367 1040 2371 1044
rect 2455 1040 2459 1044
rect 2543 1040 2547 1044
rect 2631 1040 2635 1044
rect 2719 1040 2723 1044
rect 2807 1040 2811 1044
rect 3463 1037 3467 1041
rect 2447 1031 2451 1035
rect 2615 1031 2619 1035
rect 2703 1031 2707 1035
rect 2791 1031 2795 1035
rect 2879 1031 2883 1035
rect 767 1024 771 1028
rect 927 1024 931 1028
rect 1079 1024 1083 1028
rect 1231 1024 1235 1028
rect 1383 1024 1387 1028
rect 1535 1024 1539 1028
rect 1671 1024 1675 1028
rect 1767 1021 1771 1025
rect 1807 1020 1811 1024
rect 2103 1021 2107 1025
rect 2191 1021 2195 1025
rect 2279 1021 2283 1025
rect 2367 1021 2371 1025
rect 2455 1021 2459 1025
rect 2543 1021 2547 1025
rect 2631 1021 2635 1025
rect 2719 1021 2723 1025
rect 2807 1021 2811 1025
rect 3463 1020 3467 1024
rect 847 1015 851 1019
rect 1047 1015 1051 1019
rect 1159 1015 1163 1019
rect 1471 1015 1475 1019
rect 1607 1015 1611 1019
rect 1615 1015 1619 1019
rect 111 1004 115 1008
rect 327 1005 331 1009
rect 463 1005 467 1009
rect 607 1005 611 1009
rect 767 1005 771 1009
rect 927 1005 931 1009
rect 1079 1005 1083 1009
rect 1231 1005 1235 1009
rect 1383 1005 1387 1009
rect 1535 1005 1539 1009
rect 1671 1005 1675 1009
rect 1767 1004 1771 1008
rect 1807 976 1811 980
rect 2311 975 2315 979
rect 2407 975 2411 979
rect 2511 975 2515 979
rect 2623 975 2627 979
rect 2751 975 2755 979
rect 2895 975 2899 979
rect 3055 975 3059 979
rect 3223 975 3227 979
rect 3367 975 3371 979
rect 3463 976 3467 980
rect 111 956 115 960
rect 471 955 475 959
rect 567 955 571 959
rect 671 955 675 959
rect 783 955 787 959
rect 887 955 891 959
rect 991 955 995 959
rect 1095 955 1099 959
rect 1199 955 1203 959
rect 1295 955 1299 959
rect 1391 955 1395 959
rect 1487 955 1491 959
rect 1583 955 1587 959
rect 1671 955 1675 959
rect 1767 956 1771 960
rect 1807 959 1811 963
rect 2383 963 2387 967
rect 2479 963 2483 967
rect 2503 967 2507 971
rect 2695 963 2699 967
rect 2823 963 2827 967
rect 2967 963 2971 967
rect 3127 963 3131 967
rect 3139 967 3143 971
rect 3439 967 3443 971
rect 2311 956 2315 960
rect 2407 956 2411 960
rect 2511 956 2515 960
rect 2623 956 2627 960
rect 2751 956 2755 960
rect 2895 956 2899 960
rect 3055 956 3059 960
rect 3223 956 3227 960
rect 3367 956 3371 960
rect 3463 959 3467 963
rect 111 939 115 943
rect 543 943 547 947
rect 639 943 643 947
rect 743 943 747 947
rect 855 943 859 947
rect 959 947 963 951
rect 1063 943 1067 947
rect 1167 943 1171 947
rect 1271 943 1275 947
rect 1367 943 1371 947
rect 1463 947 1467 951
rect 1559 943 1563 947
rect 1655 943 1659 947
rect 1743 943 1747 947
rect 3139 947 3143 951
rect 471 936 475 940
rect 567 936 571 940
rect 671 936 675 940
rect 783 936 787 940
rect 887 936 891 940
rect 991 936 995 940
rect 1095 936 1099 940
rect 1199 936 1203 940
rect 1295 936 1299 940
rect 1391 936 1395 940
rect 1487 936 1491 940
rect 1583 936 1587 940
rect 1671 936 1675 940
rect 1767 939 1771 943
rect 2223 939 2227 943
rect 2383 939 2387 943
rect 2479 939 2483 943
rect 2695 939 2699 943
rect 2879 939 2883 943
rect 2967 939 2971 943
rect 3127 939 3131 943
rect 3431 939 3435 943
rect 1615 927 1619 931
rect 527 919 528 923
rect 528 919 531 923
rect 543 919 547 923
rect 639 919 643 923
rect 743 919 747 923
rect 855 919 859 923
rect 1047 919 1048 923
rect 1048 919 1051 923
rect 1167 919 1171 923
rect 1271 919 1275 923
rect 1367 919 1371 923
rect 1559 919 1563 923
rect 1655 919 1659 923
rect 2823 923 2827 927
rect 1303 911 1307 915
rect 1743 915 1747 919
rect 2039 915 2040 919
rect 2040 915 2043 919
rect 2055 915 2059 919
rect 2599 915 2603 919
rect 775 903 779 907
rect 871 903 875 907
rect 1023 903 1027 907
rect 1063 903 1067 907
rect 1183 903 1187 907
rect 1567 903 1571 907
rect 1631 903 1635 907
rect 3007 915 3011 919
rect 3439 915 3443 919
rect 1807 897 1811 901
rect 1831 900 1835 904
rect 1983 900 1987 904
rect 2151 900 2155 904
rect 2327 900 2331 904
rect 2519 900 2523 904
rect 2719 900 2723 904
rect 2935 900 2939 904
rect 111 885 115 889
rect 607 888 611 892
rect 695 888 699 892
rect 791 888 795 892
rect 895 888 899 892
rect 999 888 1003 892
rect 1111 888 1115 892
rect 1223 888 1227 892
rect 1343 888 1347 892
rect 1463 888 1467 892
rect 1583 888 1587 892
rect 1895 891 1899 895
rect 2055 891 2059 895
rect 2223 891 2227 895
rect 2399 891 2403 895
rect 2599 891 2603 895
rect 3007 891 3011 895
rect 3159 900 3163 904
rect 3367 900 3371 904
rect 3463 897 3467 901
rect 3431 891 3435 895
rect 1767 885 1771 889
rect 527 879 531 883
rect 775 879 779 883
rect 871 879 875 883
rect 1183 879 1187 883
rect 1199 879 1203 883
rect 1303 879 1307 883
rect 1567 879 1571 883
rect 1807 880 1811 884
rect 1831 881 1835 885
rect 1983 881 1987 885
rect 2151 881 2155 885
rect 2327 881 2331 885
rect 2519 881 2523 885
rect 2719 881 2723 885
rect 2935 881 2939 885
rect 3159 881 3163 885
rect 3367 881 3371 885
rect 3463 880 3467 884
rect 111 868 115 872
rect 607 869 611 873
rect 695 869 699 873
rect 791 869 795 873
rect 895 869 899 873
rect 999 869 1003 873
rect 1111 869 1115 873
rect 1223 869 1227 873
rect 1343 869 1347 873
rect 1463 869 1467 873
rect 1583 869 1587 873
rect 1767 868 1771 872
rect 1807 832 1811 836
rect 1831 831 1835 835
rect 1959 831 1963 835
rect 2087 831 2091 835
rect 2207 831 2211 835
rect 2327 831 2331 835
rect 2463 831 2467 835
rect 2615 831 2619 835
rect 2791 831 2795 835
rect 2983 831 2987 835
rect 3183 831 3187 835
rect 3367 831 3371 835
rect 3463 832 3467 836
rect 111 820 115 824
rect 519 819 523 823
rect 615 819 619 823
rect 719 819 723 823
rect 831 819 835 823
rect 951 819 955 823
rect 1071 819 1075 823
rect 1191 819 1195 823
rect 1311 819 1315 823
rect 1431 819 1435 823
rect 1559 819 1563 823
rect 1767 820 1771 824
rect 111 803 115 807
rect 519 800 523 804
rect 687 807 691 811
rect 791 807 795 811
rect 903 807 907 811
rect 1023 811 1027 815
rect 1143 807 1147 811
rect 1263 807 1267 811
rect 1383 807 1387 811
rect 1503 807 1507 811
rect 1631 811 1635 815
rect 1807 815 1811 819
rect 1903 819 1907 823
rect 2031 819 2035 823
rect 2039 823 2043 827
rect 2279 819 2283 823
rect 2287 823 2291 827
rect 2535 819 2539 823
rect 2687 819 2691 823
rect 2863 819 2867 823
rect 3055 819 3059 823
rect 3139 823 3143 827
rect 3439 823 3443 827
rect 1831 812 1835 816
rect 1959 812 1963 816
rect 2087 812 2091 816
rect 2207 812 2211 816
rect 2327 812 2331 816
rect 2463 812 2467 816
rect 2615 812 2619 816
rect 2791 812 2795 816
rect 2983 812 2987 816
rect 3183 812 3187 816
rect 3367 812 3371 816
rect 3463 815 3467 819
rect 615 800 619 804
rect 719 800 723 804
rect 831 800 835 804
rect 951 800 955 804
rect 1071 800 1075 804
rect 1191 800 1195 804
rect 1311 800 1315 804
rect 1431 800 1435 804
rect 1559 800 1563 804
rect 1767 803 1771 807
rect 2287 803 2291 807
rect 1895 795 1899 799
rect 1903 795 1907 799
rect 2223 795 2227 799
rect 2279 795 2283 799
rect 2399 795 2403 799
rect 2535 795 2539 799
rect 2687 795 2691 799
rect 2863 795 2867 799
rect 3055 795 3059 799
rect 3431 795 3435 799
rect 687 783 691 787
rect 791 783 795 787
rect 903 783 907 787
rect 1199 783 1203 787
rect 1231 783 1235 787
rect 1263 783 1267 787
rect 1383 783 1387 787
rect 1503 783 1507 787
rect 3139 787 3143 791
rect 759 775 763 779
rect 2031 779 2035 783
rect 2231 779 2235 783
rect 2367 779 2371 783
rect 2487 779 2491 783
rect 2631 779 2635 783
rect 2783 779 2787 783
rect 2943 779 2947 783
rect 3111 779 3115 783
rect 3439 779 3443 783
rect 455 767 459 771
rect 543 767 547 771
rect 647 767 651 771
rect 751 767 755 771
rect 991 767 995 771
rect 1143 767 1147 771
rect 1239 767 1243 771
rect 1367 767 1371 771
rect 655 759 659 763
rect 1807 761 1811 765
rect 1879 764 1883 768
rect 2015 764 2019 768
rect 2151 764 2155 768
rect 2287 764 2291 768
rect 2423 764 2427 768
rect 2559 764 2563 768
rect 2711 764 2715 768
rect 2871 764 2875 768
rect 3039 764 3043 768
rect 3215 764 3219 768
rect 3367 764 3371 768
rect 3463 761 3467 765
rect 111 749 115 753
rect 383 752 387 756
rect 471 752 475 756
rect 575 752 579 756
rect 679 752 683 756
rect 791 752 795 756
rect 911 752 915 756
rect 1031 752 1035 756
rect 1159 752 1163 756
rect 1287 752 1291 756
rect 1415 752 1419 756
rect 2223 755 2227 759
rect 2231 755 2235 759
rect 2367 755 2371 759
rect 2631 755 2635 759
rect 2783 755 2787 759
rect 2943 755 2947 759
rect 3111 755 3115 759
rect 3279 755 3283 759
rect 3431 755 3435 759
rect 1767 749 1771 753
rect 455 743 459 747
rect 543 743 547 747
rect 647 743 651 747
rect 751 743 755 747
rect 759 743 763 747
rect 991 743 995 747
rect 1231 743 1235 747
rect 1239 743 1243 747
rect 1367 743 1371 747
rect 1807 744 1811 748
rect 1879 745 1883 749
rect 1963 747 1967 751
rect 2015 745 2019 749
rect 2151 745 2155 749
rect 2287 745 2291 749
rect 2423 745 2427 749
rect 2559 745 2563 749
rect 2711 745 2715 749
rect 2871 745 2875 749
rect 3039 745 3043 749
rect 3215 745 3219 749
rect 3367 745 3371 749
rect 3463 744 3467 748
rect 111 732 115 736
rect 383 733 387 737
rect 471 733 475 737
rect 575 733 579 737
rect 679 733 683 737
rect 791 733 795 737
rect 911 733 915 737
rect 995 735 999 739
rect 1031 733 1035 737
rect 1159 733 1163 737
rect 1287 733 1291 737
rect 1415 733 1419 737
rect 1767 732 1771 736
rect 1807 696 1811 700
rect 1831 695 1835 699
rect 1951 695 1955 699
rect 2103 695 2107 699
rect 2263 695 2267 699
rect 2415 695 2419 699
rect 2567 695 2571 699
rect 2719 695 2723 699
rect 2879 695 2883 699
rect 3039 695 3043 699
rect 3199 695 3203 699
rect 3463 696 3467 700
rect 1751 687 1755 691
rect 1911 687 1915 691
rect 111 680 115 684
rect 247 679 251 683
rect 343 679 347 683
rect 455 679 459 683
rect 567 679 571 683
rect 695 679 699 683
rect 831 679 835 683
rect 983 679 987 683
rect 1151 679 1155 683
rect 1327 679 1331 683
rect 1511 679 1515 683
rect 1671 679 1675 683
rect 1767 680 1771 684
rect 1807 679 1811 683
rect 2175 683 2179 687
rect 2335 683 2339 687
rect 2487 687 2491 691
rect 2647 687 2651 691
rect 2799 687 2803 691
rect 1831 676 1835 680
rect 111 663 115 667
rect 319 667 323 671
rect 415 667 419 671
rect 527 667 531 671
rect 639 667 643 671
rect 655 671 659 675
rect 823 671 827 675
rect 911 671 915 675
rect 1951 676 1955 680
rect 2103 676 2107 680
rect 2263 676 2267 680
rect 2415 676 2419 680
rect 2567 676 2571 680
rect 2631 679 2635 683
rect 3111 683 3115 687
rect 3139 687 3143 691
rect 2719 676 2723 680
rect 2879 676 2883 680
rect 3039 676 3043 680
rect 3199 676 3203 680
rect 3463 679 3467 683
rect 1295 667 1299 671
rect 1399 667 1403 671
rect 1743 667 1747 671
rect 247 660 251 664
rect 343 660 347 664
rect 455 660 459 664
rect 567 660 571 664
rect 695 660 699 664
rect 831 660 835 664
rect 983 660 987 664
rect 1151 660 1155 664
rect 1327 660 1331 664
rect 1511 660 1515 664
rect 1671 660 1675 664
rect 1767 663 1771 667
rect 3139 667 3143 671
rect 1911 659 1915 663
rect 1963 659 1967 663
rect 2159 659 2160 663
rect 2160 659 2163 663
rect 2175 659 2179 663
rect 2335 659 2339 663
rect 2647 659 2651 663
rect 2799 659 2803 663
rect 2951 659 2955 663
rect 3279 659 3283 663
rect 319 643 323 647
rect 415 643 419 647
rect 527 643 531 647
rect 639 643 643 647
rect 911 643 915 647
rect 995 643 999 647
rect 1287 643 1291 647
rect 1295 643 1299 647
rect 1399 643 1403 647
rect 1751 643 1755 647
rect 1967 647 1971 651
rect 2047 647 2051 651
rect 2551 647 2555 651
rect 2759 647 2763 651
rect 3111 647 3112 651
rect 3112 647 3115 651
rect 3127 647 3131 651
rect 3431 647 3435 651
rect 2839 639 2843 643
rect 199 627 203 631
rect 207 627 211 631
rect 303 627 307 631
rect 431 627 435 631
rect 559 627 563 631
rect 823 627 824 631
rect 824 627 827 631
rect 111 609 115 613
rect 135 612 139 616
rect 231 612 235 616
rect 359 612 363 616
rect 487 612 491 616
rect 623 612 627 616
rect 767 612 771 616
rect 207 603 211 607
rect 303 603 307 607
rect 431 603 435 607
rect 559 603 563 607
rect 1111 627 1112 631
rect 1112 627 1115 631
rect 1127 627 1131 631
rect 1279 627 1283 631
rect 1607 627 1611 631
rect 1743 627 1747 631
rect 1807 629 1811 633
rect 1975 632 1979 636
rect 2239 632 2243 636
rect 2479 632 2483 636
rect 2687 632 2691 636
rect 2879 632 2883 636
rect 3055 632 3059 636
rect 3223 632 3227 636
rect 3367 632 3371 636
rect 3463 629 3467 633
rect 2047 623 2051 627
rect 2159 623 2163 627
rect 2551 623 2555 627
rect 2759 623 2763 627
rect 2951 623 2955 627
rect 3127 623 3131 627
rect 3191 623 3195 627
rect 3439 623 3443 627
rect 911 612 915 616
rect 1055 612 1059 616
rect 1207 612 1211 616
rect 1367 612 1371 616
rect 1527 612 1531 616
rect 1671 612 1675 616
rect 1767 609 1771 613
rect 1807 612 1811 616
rect 1975 613 1979 617
rect 2239 613 2243 617
rect 2479 613 2483 617
rect 2687 613 2691 617
rect 2879 613 2883 617
rect 3055 613 3059 617
rect 3223 613 3227 617
rect 3367 613 3371 617
rect 3463 612 3467 616
rect 983 603 987 607
rect 1127 603 1131 607
rect 1279 603 1283 607
rect 1287 603 1291 607
rect 1447 603 1451 607
rect 1607 603 1611 607
rect 111 592 115 596
rect 135 593 139 597
rect 231 593 235 597
rect 359 593 363 597
rect 487 593 491 597
rect 623 593 627 597
rect 767 593 771 597
rect 911 593 915 597
rect 1055 593 1059 597
rect 1207 593 1211 597
rect 1367 593 1371 597
rect 1527 593 1531 597
rect 1671 593 1675 597
rect 1767 592 1771 596
rect 1807 560 1811 564
rect 1895 559 1899 563
rect 2015 559 2019 563
rect 2143 559 2147 563
rect 2279 559 2283 563
rect 2423 559 2427 563
rect 2567 559 2571 563
rect 2719 559 2723 563
rect 2871 559 2875 563
rect 3031 559 3035 563
rect 3199 559 3203 563
rect 3367 559 3371 563
rect 3463 560 3467 564
rect 1967 551 1971 555
rect 1975 551 1979 555
rect 2095 551 2099 555
rect 2223 551 2227 555
rect 2411 551 2415 555
rect 111 544 115 548
rect 135 543 139 547
rect 199 539 203 543
rect 247 543 251 547
rect 407 543 411 547
rect 583 543 587 547
rect 767 543 771 547
rect 951 543 955 547
rect 1135 543 1139 547
rect 1319 543 1323 547
rect 1503 543 1507 547
rect 1671 543 1675 547
rect 1767 544 1771 548
rect 1807 543 1811 547
rect 2639 547 2643 551
rect 2791 547 2795 551
rect 2839 551 2843 555
rect 3103 547 3107 551
rect 3139 551 3143 555
rect 3431 555 3435 559
rect 1895 540 1899 544
rect 215 535 219 539
rect 327 535 331 539
rect 111 527 115 531
rect 655 531 659 535
rect 743 535 747 539
rect 2015 540 2019 544
rect 2143 540 2147 544
rect 2279 540 2283 544
rect 2423 540 2427 544
rect 2567 540 2571 544
rect 2719 540 2723 544
rect 2871 540 2875 544
rect 3031 540 3035 544
rect 3199 540 3203 544
rect 3367 540 3371 544
rect 3463 543 3467 547
rect 1023 531 1027 535
rect 1111 535 1115 539
rect 1391 531 1395 535
rect 1575 531 1579 535
rect 1743 531 1747 535
rect 135 524 139 528
rect 247 524 251 528
rect 407 524 411 528
rect 583 524 587 528
rect 767 524 771 528
rect 951 524 955 528
rect 1135 524 1139 528
rect 1319 524 1323 528
rect 1503 524 1507 528
rect 1671 524 1675 528
rect 1767 527 1771 531
rect 3139 531 3143 535
rect 1975 523 1979 527
rect 2095 523 2099 527
rect 2223 523 2227 527
rect 2411 523 2415 527
rect 2431 523 2435 527
rect 2631 523 2635 527
rect 2639 523 2643 527
rect 3079 523 3083 527
rect 3103 523 3107 527
rect 3431 523 3435 527
rect 743 515 747 519
rect 1447 515 1451 519
rect 2207 515 2211 519
rect 215 507 219 511
rect 327 507 331 511
rect 635 507 636 511
rect 636 507 639 511
rect 655 507 659 511
rect 983 507 987 511
rect 1023 507 1027 511
rect 1391 507 1395 511
rect 1575 507 1579 511
rect 2311 507 2315 511
rect 2671 507 2672 511
rect 2672 507 2675 511
rect 2791 507 2795 511
rect 2951 507 2955 511
rect 3191 507 3192 511
rect 3192 507 3195 511
rect 3207 507 3211 511
rect 3439 507 3443 511
rect 319 491 323 495
rect 471 491 475 495
rect 815 491 819 495
rect 999 491 1003 495
rect 1187 491 1191 495
rect 1607 491 1611 495
rect 1743 491 1747 495
rect 1807 489 1811 493
rect 2135 492 2139 496
rect 2239 492 2243 496
rect 2359 492 2363 496
rect 111 473 115 477
rect 247 476 251 480
rect 399 476 403 480
rect 567 476 571 480
rect 319 467 323 471
rect 471 467 475 471
rect 635 467 639 471
rect 735 476 739 480
rect 903 476 907 480
rect 1063 476 1067 480
rect 1223 476 1227 480
rect 815 467 819 471
rect 1187 467 1191 471
rect 1295 467 1299 471
rect 2207 483 2211 487
rect 2311 483 2315 487
rect 2431 483 2435 487
rect 3103 499 3107 503
rect 2487 492 2491 496
rect 2615 492 2619 496
rect 2751 492 2755 496
rect 2879 492 2883 496
rect 3007 492 3011 496
rect 3135 492 3139 496
rect 3263 492 3267 496
rect 3367 492 3371 496
rect 3463 489 3467 493
rect 2823 483 2827 487
rect 2951 483 2955 487
rect 3079 483 3083 487
rect 3207 483 3211 487
rect 3327 483 3331 487
rect 3431 483 3435 487
rect 1375 476 1379 480
rect 1527 476 1531 480
rect 1671 476 1675 480
rect 1767 473 1771 477
rect 1807 472 1811 476
rect 2135 473 2139 477
rect 2239 473 2243 477
rect 2359 473 2363 477
rect 2487 473 2491 477
rect 2615 473 2619 477
rect 2751 473 2755 477
rect 2879 473 2883 477
rect 3007 473 3011 477
rect 3135 473 3139 477
rect 3263 473 3267 477
rect 3367 473 3371 477
rect 3463 472 3467 476
rect 1607 467 1611 471
rect 111 456 115 460
rect 247 457 251 461
rect 399 457 403 461
rect 567 457 571 461
rect 735 457 739 461
rect 903 457 907 461
rect 1063 457 1067 461
rect 1223 457 1227 461
rect 1375 457 1379 461
rect 1527 457 1531 461
rect 1671 457 1675 461
rect 1767 456 1771 460
rect 1807 420 1811 424
rect 2239 419 2243 423
rect 2335 419 2339 423
rect 2447 419 2451 423
rect 2559 419 2563 423
rect 2679 419 2683 423
rect 2799 419 2803 423
rect 2911 419 2915 423
rect 3023 419 3027 423
rect 3143 419 3147 423
rect 3263 419 3267 423
rect 3367 419 3371 423
rect 3463 420 3467 424
rect 111 408 115 412
rect 519 407 523 411
rect 615 407 619 411
rect 719 407 723 411
rect 823 407 827 411
rect 927 407 931 411
rect 1023 407 1027 411
rect 1127 407 1131 411
rect 1231 407 1235 411
rect 1335 407 1339 411
rect 1439 407 1443 411
rect 1767 408 1771 412
rect 111 391 115 395
rect 591 395 595 399
rect 687 395 691 399
rect 799 399 803 403
rect 999 399 1003 403
rect 519 388 523 392
rect 615 388 619 392
rect 719 388 723 392
rect 1095 395 1099 399
rect 1199 395 1203 399
rect 1207 399 1211 403
rect 1407 395 1411 399
rect 1415 399 1419 403
rect 1807 403 1811 407
rect 2239 400 2243 404
rect 799 379 803 383
rect 823 388 827 392
rect 927 388 931 392
rect 1023 388 1027 392
rect 1127 388 1131 392
rect 1231 388 1235 392
rect 1335 388 1339 392
rect 1439 388 1443 392
rect 1767 391 1771 395
rect 2407 407 2411 411
rect 2519 407 2523 411
rect 2631 407 2635 411
rect 2671 411 2675 415
rect 2871 407 2875 411
rect 2983 407 2987 411
rect 3095 407 3099 411
rect 3103 411 3107 415
rect 3335 407 3339 411
rect 3439 411 3443 415
rect 2335 400 2339 404
rect 2447 400 2451 404
rect 2559 400 2563 404
rect 2679 400 2683 404
rect 2799 400 2803 404
rect 2911 400 2915 404
rect 3023 400 3027 404
rect 3143 400 3147 404
rect 3263 400 3267 404
rect 3367 400 3371 404
rect 3463 403 3467 407
rect 1207 379 1211 383
rect 1415 379 1419 383
rect 2407 383 2411 387
rect 2519 383 2523 387
rect 2631 383 2635 387
rect 2823 383 2827 387
rect 2975 383 2979 387
rect 2983 383 2987 387
rect 3095 383 3099 387
rect 3327 383 3331 387
rect 3431 383 3435 387
rect 591 371 595 375
rect 687 371 691 375
rect 887 371 891 375
rect 1095 371 1099 375
rect 1295 371 1299 375
rect 1407 371 1411 375
rect 2439 375 2443 379
rect 2135 367 2139 371
rect 2223 367 2227 371
rect 2319 367 2323 371
rect 2431 367 2435 371
rect 2695 367 2699 371
rect 2871 367 2875 371
rect 2991 367 2995 371
rect 3159 367 3163 371
rect 3167 367 3171 371
rect 3439 367 3443 371
rect 543 355 547 359
rect 631 355 635 359
rect 807 355 811 359
rect 991 355 995 359
rect 1079 355 1083 359
rect 639 347 643 351
rect 1199 355 1203 359
rect 1247 355 1251 359
rect 2423 359 2427 363
rect 1807 349 1811 353
rect 2063 352 2067 356
rect 2151 352 2155 356
rect 2247 352 2251 356
rect 2359 352 2363 356
rect 2479 352 2483 356
rect 2615 352 2619 356
rect 2759 352 2763 356
rect 2911 352 2915 356
rect 3063 352 3067 356
rect 3223 352 3227 356
rect 3367 352 3371 356
rect 3463 349 3467 353
rect 111 337 115 341
rect 471 340 475 344
rect 559 340 563 344
rect 647 340 651 344
rect 735 340 739 344
rect 823 340 827 344
rect 911 340 915 344
rect 999 340 1003 344
rect 1087 340 1091 344
rect 1175 340 1179 344
rect 543 331 547 335
rect 631 331 635 335
rect 807 331 811 335
rect 887 331 891 335
rect 903 331 907 335
rect 991 331 995 335
rect 1079 331 1083 335
rect 1247 331 1251 335
rect 1263 340 1267 344
rect 2135 343 2139 347
rect 2223 343 2227 347
rect 2319 343 2323 347
rect 2431 343 2435 347
rect 2439 343 2443 347
rect 2679 343 2683 347
rect 2695 343 2699 347
rect 2975 343 2979 347
rect 2991 343 2995 347
rect 3159 343 3163 347
rect 3431 343 3435 347
rect 1767 337 1771 341
rect 1807 332 1811 336
rect 2063 333 2067 337
rect 2151 333 2155 337
rect 2247 333 2251 337
rect 2359 333 2363 337
rect 2479 333 2483 337
rect 2615 333 2619 337
rect 2759 333 2763 337
rect 2911 333 2915 337
rect 3063 333 3067 337
rect 3223 333 3227 337
rect 3367 333 3371 337
rect 3463 332 3467 336
rect 111 320 115 324
rect 471 321 475 325
rect 559 321 563 325
rect 647 321 651 325
rect 735 321 739 325
rect 823 321 827 325
rect 911 321 915 325
rect 999 321 1003 325
rect 1087 321 1091 325
rect 1175 321 1179 325
rect 1263 321 1267 325
rect 1767 320 1771 324
rect 1807 284 1811 288
rect 1927 283 1931 287
rect 2039 283 2043 287
rect 2167 283 2171 287
rect 2303 283 2307 287
rect 2447 283 2451 287
rect 2599 283 2603 287
rect 2759 283 2763 287
rect 2919 283 2923 287
rect 3087 283 3091 287
rect 3255 283 3259 287
rect 3463 284 3467 288
rect 111 272 115 276
rect 279 271 283 275
rect 367 271 371 275
rect 463 271 467 275
rect 559 271 563 275
rect 655 271 659 275
rect 751 271 755 275
rect 847 271 851 275
rect 943 271 947 275
rect 1047 271 1051 275
rect 1151 271 1155 275
rect 1767 272 1771 276
rect 111 255 115 259
rect 351 259 355 263
rect 439 259 443 263
rect 535 259 539 263
rect 631 259 635 263
rect 639 263 643 267
rect 823 259 827 263
rect 919 259 923 263
rect 1015 259 1019 263
rect 1119 259 1123 263
rect 1127 263 1131 267
rect 1807 267 1811 271
rect 1999 271 2003 275
rect 2111 271 2115 275
rect 2239 271 2243 275
rect 2375 271 2379 275
rect 2423 275 2427 279
rect 2671 271 2675 275
rect 2831 271 2835 275
rect 2991 271 2995 275
rect 3167 275 3171 279
rect 1927 264 1931 268
rect 2039 264 2043 268
rect 2167 264 2171 268
rect 2303 264 2307 268
rect 2447 264 2451 268
rect 2599 264 2603 268
rect 2759 264 2763 268
rect 2919 264 2923 268
rect 3087 264 3091 268
rect 3255 264 3259 268
rect 3463 267 3467 271
rect 279 252 283 256
rect 367 252 371 256
rect 463 252 467 256
rect 559 252 563 256
rect 655 252 659 256
rect 751 252 755 256
rect 847 252 851 256
rect 943 252 947 256
rect 1047 252 1051 256
rect 1151 252 1155 256
rect 1767 255 1771 259
rect 903 243 907 247
rect 1999 247 2003 251
rect 2111 247 2115 251
rect 2239 247 2243 251
rect 2375 247 2379 251
rect 2679 247 2683 251
rect 2815 247 2816 251
rect 2816 247 2819 251
rect 2831 247 2835 251
rect 2991 247 2995 251
rect 3335 247 3339 251
rect 351 235 355 239
rect 439 235 443 239
rect 535 235 539 239
rect 631 235 635 239
rect 823 235 827 239
rect 919 235 923 239
rect 1015 235 1019 239
rect 1119 235 1123 239
rect 2323 239 2327 243
rect 591 227 595 231
rect 1127 227 1131 231
rect 1903 231 1907 235
rect 1999 231 2003 235
rect 2127 231 2131 235
rect 2271 231 2275 235
rect 2591 231 2595 235
rect 2671 231 2675 235
rect 2927 231 2931 235
rect 3127 231 3131 235
rect 3431 231 3435 235
rect 231 219 235 223
rect 239 219 243 223
rect 415 219 419 223
rect 583 219 587 223
rect 911 219 915 223
rect 1063 219 1067 223
rect 1207 219 1211 223
rect 1351 219 1355 223
rect 2239 223 2243 227
rect 1807 213 1811 217
rect 1831 216 1835 220
rect 1927 216 1931 220
rect 2055 216 2059 220
rect 2199 216 2203 220
rect 2351 216 2355 220
rect 2511 216 2515 220
rect 2679 216 2683 220
rect 2847 216 2851 220
rect 3023 216 3027 220
rect 3207 216 3211 220
rect 3367 216 3371 220
rect 3463 213 3467 217
rect 111 201 115 205
rect 167 204 171 208
rect 343 204 347 208
rect 511 204 515 208
rect 679 204 683 208
rect 839 204 843 208
rect 991 204 995 208
rect 1135 204 1139 208
rect 1279 204 1283 208
rect 1431 204 1435 208
rect 1903 207 1907 211
rect 1999 207 2003 211
rect 2127 207 2131 211
rect 2271 207 2275 211
rect 2323 207 2327 211
rect 2455 207 2459 211
rect 2591 207 2595 211
rect 2815 207 2819 211
rect 2927 207 2931 211
rect 3271 207 3275 211
rect 3439 207 3443 211
rect 1767 201 1771 205
rect 239 195 243 199
rect 415 195 419 199
rect 583 195 587 199
rect 591 195 595 199
rect 911 195 915 199
rect 1063 195 1067 199
rect 1207 195 1211 199
rect 1351 195 1355 199
rect 1399 195 1403 199
rect 1807 196 1811 200
rect 1831 197 1835 201
rect 1927 197 1931 201
rect 2055 197 2059 201
rect 2199 197 2203 201
rect 2351 197 2355 201
rect 2511 197 2515 201
rect 2679 197 2683 201
rect 2847 197 2851 201
rect 3023 197 3027 201
rect 3207 197 3211 201
rect 3367 197 3371 201
rect 3463 196 3467 200
rect 111 184 115 188
rect 167 185 171 189
rect 343 185 347 189
rect 511 185 515 189
rect 679 185 683 189
rect 839 185 843 189
rect 991 185 995 189
rect 1135 185 1139 189
rect 1279 185 1283 189
rect 1431 185 1435 189
rect 1767 184 1771 188
rect 1807 132 1811 136
rect 1831 131 1835 135
rect 1919 131 1923 135
rect 2039 131 2043 135
rect 2159 131 2163 135
rect 2279 131 2283 135
rect 2399 131 2403 135
rect 2511 131 2515 135
rect 2623 131 2627 135
rect 2735 131 2739 135
rect 2839 131 2843 135
rect 2943 131 2947 135
rect 3055 131 3059 135
rect 3167 131 3171 135
rect 3279 131 3283 135
rect 3367 131 3371 135
rect 3463 132 3467 136
rect 111 116 115 120
rect 135 115 139 119
rect 223 115 227 119
rect 311 115 315 119
rect 399 115 403 119
rect 487 115 491 119
rect 575 115 579 119
rect 663 115 667 119
rect 751 115 755 119
rect 847 115 851 119
rect 943 115 947 119
rect 1031 115 1035 119
rect 1119 115 1123 119
rect 1215 115 1219 119
rect 1311 115 1315 119
rect 1407 115 1411 119
rect 1495 115 1499 119
rect 1583 115 1587 119
rect 1671 115 1675 119
rect 1767 116 1771 120
rect 1807 115 1811 119
rect 1903 119 1907 123
rect 1991 119 1995 123
rect 2111 119 2115 123
rect 2231 119 2235 123
rect 2239 123 2243 127
rect 2471 119 2475 123
rect 2583 119 2587 123
rect 2695 119 2699 123
rect 2807 119 2811 123
rect 2911 119 2915 123
rect 3015 119 3019 123
rect 3127 123 3131 127
rect 3431 127 3435 131
rect 1831 112 1835 116
rect 1919 112 1923 116
rect 2039 112 2043 116
rect 2159 112 2163 116
rect 2279 112 2283 116
rect 2399 112 2403 116
rect 2511 112 2515 116
rect 2623 112 2627 116
rect 2735 112 2739 116
rect 2839 112 2843 116
rect 2943 112 2947 116
rect 3055 112 3059 116
rect 3167 112 3171 116
rect 111 99 115 103
rect 207 103 211 107
rect 295 103 299 107
rect 383 103 387 107
rect 471 103 475 107
rect 559 103 563 107
rect 647 103 651 107
rect 735 103 739 107
rect 743 107 747 111
rect 919 103 923 107
rect 1015 103 1019 107
rect 1103 103 1107 107
rect 1191 103 1195 107
rect 1287 103 1291 107
rect 1383 103 1387 107
rect 1479 103 1483 107
rect 1567 103 1571 107
rect 1655 103 1659 107
rect 3351 119 3355 123
rect 3279 112 3283 116
rect 3367 112 3371 116
rect 3463 115 3467 119
rect 135 96 139 100
rect 223 96 227 100
rect 311 96 315 100
rect 399 96 403 100
rect 487 96 491 100
rect 575 96 579 100
rect 663 96 667 100
rect 751 96 755 100
rect 847 96 851 100
rect 943 96 947 100
rect 1031 96 1035 100
rect 1119 96 1123 100
rect 1215 96 1219 100
rect 1311 96 1315 100
rect 1407 96 1411 100
rect 1495 96 1499 100
rect 1583 96 1587 100
rect 1671 96 1675 100
rect 1767 99 1771 103
rect 1903 95 1907 99
rect 1991 95 1995 99
rect 2111 95 2115 99
rect 2231 95 2235 99
rect 2455 95 2456 99
rect 2456 95 2459 99
rect 2471 95 2475 99
rect 2583 95 2587 99
rect 2695 95 2699 99
rect 2807 95 2811 99
rect 2911 95 2915 99
rect 3015 95 3019 99
rect 3271 95 3275 99
rect 3351 95 3355 99
rect 207 79 211 83
rect 295 79 299 83
rect 383 79 387 83
rect 471 79 475 83
rect 559 79 563 83
rect 647 79 651 83
rect 735 79 739 83
rect 903 79 904 83
rect 904 79 907 83
rect 919 79 923 83
rect 1015 79 1019 83
rect 1103 79 1107 83
rect 1191 79 1195 83
rect 1287 79 1291 83
rect 1383 79 1387 83
rect 1479 79 1483 83
rect 1567 79 1571 83
rect 1655 79 1659 83
<< m3 >>
rect 1807 3522 1811 3523
rect 1807 3517 1811 3518
rect 2007 3522 2011 3523
rect 2007 3517 2011 3518
rect 2239 3522 2243 3523
rect 2239 3517 2243 3518
rect 2455 3522 2459 3523
rect 2455 3517 2459 3518
rect 2655 3522 2659 3523
rect 2655 3517 2659 3518
rect 2855 3522 2859 3523
rect 2855 3517 2859 3518
rect 3047 3522 3051 3523
rect 3047 3517 3051 3518
rect 3247 3522 3251 3523
rect 3247 3517 3251 3518
rect 3463 3522 3467 3523
rect 3463 3517 3467 3518
rect 1808 3501 1810 3517
rect 1806 3500 1812 3501
rect 2008 3500 2010 3517
rect 2240 3500 2242 3517
rect 2456 3500 2458 3517
rect 2656 3500 2658 3517
rect 2856 3500 2858 3517
rect 3048 3500 3050 3517
rect 3248 3500 3250 3517
rect 3464 3501 3466 3517
rect 3462 3500 3468 3501
rect 1806 3496 1807 3500
rect 1811 3496 1812 3500
rect 1806 3495 1812 3496
rect 2006 3499 2012 3500
rect 2006 3495 2007 3499
rect 2011 3495 2012 3499
rect 2006 3494 2012 3495
rect 2238 3499 2244 3500
rect 2238 3495 2239 3499
rect 2243 3495 2244 3499
rect 2238 3494 2244 3495
rect 2454 3499 2460 3500
rect 2454 3495 2455 3499
rect 2459 3495 2460 3499
rect 2454 3494 2460 3495
rect 2654 3499 2660 3500
rect 2654 3495 2655 3499
rect 2659 3495 2660 3499
rect 2654 3494 2660 3495
rect 2854 3499 2860 3500
rect 2854 3495 2855 3499
rect 2859 3495 2860 3499
rect 2854 3494 2860 3495
rect 3046 3499 3052 3500
rect 3046 3495 3047 3499
rect 3051 3495 3052 3499
rect 3046 3494 3052 3495
rect 3246 3499 3252 3500
rect 3246 3495 3247 3499
rect 3251 3495 3252 3499
rect 3462 3496 3463 3500
rect 3467 3496 3468 3500
rect 3462 3495 3468 3496
rect 3246 3494 3252 3495
rect 2406 3491 2412 3492
rect 2310 3487 2316 3488
rect 111 3486 115 3487
rect 111 3481 115 3482
rect 455 3486 459 3487
rect 455 3481 459 3482
rect 543 3486 547 3487
rect 543 3481 547 3482
rect 631 3486 635 3487
rect 631 3481 635 3482
rect 719 3486 723 3487
rect 719 3481 723 3482
rect 807 3486 811 3487
rect 807 3481 811 3482
rect 895 3486 899 3487
rect 895 3481 899 3482
rect 983 3486 987 3487
rect 983 3481 987 3482
rect 1071 3486 1075 3487
rect 1071 3481 1075 3482
rect 1159 3486 1163 3487
rect 1159 3481 1163 3482
rect 1767 3486 1771 3487
rect 1767 3481 1771 3482
rect 1806 3483 1812 3484
rect 112 3465 114 3481
rect 110 3464 116 3465
rect 456 3464 458 3481
rect 544 3464 546 3481
rect 632 3464 634 3481
rect 720 3464 722 3481
rect 808 3464 810 3481
rect 896 3464 898 3481
rect 984 3464 986 3481
rect 1072 3464 1074 3481
rect 1160 3464 1162 3481
rect 1768 3465 1770 3481
rect 1806 3479 1807 3483
rect 1811 3479 1812 3483
rect 2310 3483 2311 3487
rect 2315 3483 2316 3487
rect 2406 3487 2407 3491
rect 2411 3487 2412 3491
rect 2406 3486 2412 3487
rect 2726 3487 2732 3488
rect 2310 3482 2316 3483
rect 1806 3478 1812 3479
rect 2006 3480 2012 3481
rect 1766 3464 1772 3465
rect 110 3460 111 3464
rect 115 3460 116 3464
rect 110 3459 116 3460
rect 454 3463 460 3464
rect 454 3459 455 3463
rect 459 3459 460 3463
rect 454 3458 460 3459
rect 542 3463 548 3464
rect 542 3459 543 3463
rect 547 3459 548 3463
rect 542 3458 548 3459
rect 630 3463 636 3464
rect 630 3459 631 3463
rect 635 3459 636 3463
rect 630 3458 636 3459
rect 718 3463 724 3464
rect 718 3459 719 3463
rect 723 3459 724 3463
rect 718 3458 724 3459
rect 806 3463 812 3464
rect 806 3459 807 3463
rect 811 3459 812 3463
rect 806 3458 812 3459
rect 894 3463 900 3464
rect 894 3459 895 3463
rect 899 3459 900 3463
rect 894 3458 900 3459
rect 982 3463 988 3464
rect 982 3459 983 3463
rect 987 3459 988 3463
rect 982 3458 988 3459
rect 1070 3463 1076 3464
rect 1070 3459 1071 3463
rect 1075 3459 1076 3463
rect 1070 3458 1076 3459
rect 1158 3463 1164 3464
rect 1158 3459 1159 3463
rect 1163 3459 1164 3463
rect 1766 3460 1767 3464
rect 1771 3460 1772 3464
rect 1766 3459 1772 3460
rect 1808 3459 1810 3478
rect 2006 3476 2007 3480
rect 2011 3476 2012 3480
rect 2006 3475 2012 3476
rect 2238 3480 2244 3481
rect 2238 3476 2239 3480
rect 2243 3476 2244 3480
rect 2238 3475 2244 3476
rect 2008 3459 2010 3475
rect 2014 3463 2020 3464
rect 2014 3459 2015 3463
rect 2019 3459 2020 3463
rect 2240 3459 2242 3475
rect 2312 3464 2314 3482
rect 2310 3463 2316 3464
rect 2310 3459 2311 3463
rect 2315 3459 2316 3463
rect 1158 3458 1164 3459
rect 1807 3458 1811 3459
rect 622 3455 628 3456
rect 526 3451 532 3452
rect 110 3447 116 3448
rect 110 3443 111 3447
rect 115 3443 116 3447
rect 526 3447 527 3451
rect 531 3447 532 3451
rect 526 3446 532 3447
rect 614 3451 620 3452
rect 614 3447 615 3451
rect 619 3447 620 3451
rect 622 3451 623 3455
rect 627 3451 628 3455
rect 622 3450 628 3451
rect 710 3455 716 3456
rect 710 3451 711 3455
rect 715 3451 716 3455
rect 710 3450 716 3451
rect 798 3455 804 3456
rect 798 3451 799 3455
rect 803 3451 804 3455
rect 798 3450 804 3451
rect 886 3455 892 3456
rect 886 3451 887 3455
rect 891 3451 892 3455
rect 886 3450 892 3451
rect 974 3455 980 3456
rect 974 3451 975 3455
rect 979 3451 980 3455
rect 1150 3455 1156 3456
rect 974 3450 980 3451
rect 1142 3451 1148 3452
rect 614 3446 620 3447
rect 110 3442 116 3443
rect 454 3444 460 3445
rect 112 3423 114 3442
rect 454 3440 455 3444
rect 459 3440 460 3444
rect 454 3439 460 3440
rect 456 3423 458 3439
rect 528 3428 530 3446
rect 542 3444 548 3445
rect 542 3440 543 3444
rect 547 3440 548 3444
rect 542 3439 548 3440
rect 526 3427 532 3428
rect 526 3423 527 3427
rect 531 3423 532 3427
rect 544 3423 546 3439
rect 111 3422 115 3423
rect 111 3417 115 3418
rect 415 3422 419 3423
rect 415 3417 419 3418
rect 455 3422 459 3423
rect 455 3417 459 3418
rect 503 3422 507 3423
rect 526 3422 532 3423
rect 543 3422 547 3423
rect 503 3417 507 3418
rect 543 3417 547 3418
rect 591 3422 595 3423
rect 591 3417 595 3418
rect 112 3398 114 3417
rect 416 3401 418 3417
rect 494 3415 500 3416
rect 494 3411 495 3415
rect 499 3411 500 3415
rect 494 3410 500 3411
rect 414 3400 420 3401
rect 110 3397 116 3398
rect 110 3393 111 3397
rect 115 3393 116 3397
rect 414 3396 415 3400
rect 419 3396 420 3400
rect 414 3395 420 3396
rect 110 3392 116 3393
rect 496 3392 498 3410
rect 504 3401 506 3417
rect 592 3401 594 3417
rect 616 3416 618 3446
rect 624 3436 626 3450
rect 630 3444 636 3445
rect 630 3440 631 3444
rect 635 3440 636 3444
rect 630 3439 636 3440
rect 622 3435 628 3436
rect 622 3431 623 3435
rect 627 3431 628 3435
rect 622 3430 628 3431
rect 632 3423 634 3439
rect 712 3428 714 3450
rect 718 3444 724 3445
rect 718 3440 719 3444
rect 723 3440 724 3444
rect 718 3439 724 3440
rect 710 3427 716 3428
rect 710 3423 711 3427
rect 715 3423 716 3427
rect 720 3423 722 3439
rect 800 3428 802 3450
rect 806 3444 812 3445
rect 806 3440 807 3444
rect 811 3440 812 3444
rect 806 3439 812 3440
rect 798 3427 804 3428
rect 798 3423 799 3427
rect 803 3423 804 3427
rect 808 3423 810 3439
rect 888 3428 890 3450
rect 894 3444 900 3445
rect 894 3440 895 3444
rect 899 3440 900 3444
rect 894 3439 900 3440
rect 886 3427 892 3428
rect 886 3423 887 3427
rect 891 3423 892 3427
rect 896 3423 898 3439
rect 976 3428 978 3450
rect 1142 3447 1143 3451
rect 1147 3447 1148 3451
rect 1150 3451 1151 3455
rect 1155 3451 1156 3455
rect 1807 3453 1811 3454
rect 1831 3458 1835 3459
rect 1831 3453 1835 3454
rect 1943 3458 1947 3459
rect 1943 3453 1947 3454
rect 2007 3458 2011 3459
rect 2014 3458 2020 3459
rect 2079 3458 2083 3459
rect 2007 3453 2011 3454
rect 1150 3450 1156 3451
rect 1142 3446 1148 3447
rect 982 3444 988 3445
rect 982 3440 983 3444
rect 987 3440 988 3444
rect 982 3439 988 3440
rect 1070 3444 1076 3445
rect 1070 3440 1071 3444
rect 1075 3440 1076 3444
rect 1070 3439 1076 3440
rect 974 3427 980 3428
rect 974 3423 975 3427
rect 979 3423 980 3427
rect 984 3423 986 3439
rect 1072 3423 1074 3439
rect 1144 3428 1146 3446
rect 1152 3436 1154 3450
rect 1766 3447 1772 3448
rect 1158 3444 1164 3445
rect 1158 3440 1159 3444
rect 1163 3440 1164 3444
rect 1766 3443 1767 3447
rect 1771 3443 1772 3447
rect 1766 3442 1772 3443
rect 1158 3439 1164 3440
rect 1150 3435 1156 3436
rect 1150 3431 1151 3435
rect 1155 3431 1156 3435
rect 1150 3430 1156 3431
rect 1102 3427 1108 3428
rect 1102 3423 1103 3427
rect 1107 3423 1108 3427
rect 1142 3427 1148 3428
rect 1142 3423 1143 3427
rect 1147 3423 1148 3427
rect 1160 3423 1162 3439
rect 1768 3423 1770 3442
rect 1808 3434 1810 3453
rect 1832 3437 1834 3453
rect 1902 3451 1908 3452
rect 1902 3447 1903 3451
rect 1907 3447 1908 3451
rect 1902 3446 1908 3447
rect 1830 3436 1836 3437
rect 1806 3433 1812 3434
rect 1806 3429 1807 3433
rect 1811 3429 1812 3433
rect 1830 3432 1831 3436
rect 1835 3432 1836 3436
rect 1830 3431 1836 3432
rect 1806 3428 1812 3429
rect 1904 3428 1906 3446
rect 1944 3437 1946 3453
rect 1942 3436 1948 3437
rect 1942 3432 1943 3436
rect 1947 3432 1948 3436
rect 1942 3431 1948 3432
rect 2016 3428 2018 3458
rect 2079 3453 2083 3454
rect 2215 3458 2219 3459
rect 2215 3453 2219 3454
rect 2239 3458 2243 3459
rect 2310 3458 2316 3459
rect 2351 3458 2355 3459
rect 2239 3453 2243 3454
rect 2351 3453 2355 3454
rect 2080 3437 2082 3453
rect 2166 3451 2172 3452
rect 2166 3447 2167 3451
rect 2171 3447 2172 3451
rect 2166 3446 2172 3447
rect 2078 3436 2084 3437
rect 2078 3432 2079 3436
rect 2083 3432 2084 3436
rect 2078 3431 2084 3432
rect 1902 3427 1908 3428
rect 1902 3423 1903 3427
rect 1907 3423 1908 3427
rect 631 3422 635 3423
rect 631 3417 635 3418
rect 679 3422 683 3423
rect 710 3422 716 3423
rect 719 3422 723 3423
rect 679 3417 683 3418
rect 719 3417 723 3418
rect 767 3422 771 3423
rect 798 3422 804 3423
rect 807 3422 811 3423
rect 767 3417 771 3418
rect 807 3417 811 3418
rect 855 3422 859 3423
rect 886 3422 892 3423
rect 895 3422 899 3423
rect 855 3417 859 3418
rect 895 3417 899 3418
rect 943 3422 947 3423
rect 974 3422 980 3423
rect 983 3422 987 3423
rect 943 3417 947 3418
rect 983 3417 987 3418
rect 1031 3422 1035 3423
rect 1031 3417 1035 3418
rect 1071 3422 1075 3423
rect 1102 3422 1108 3423
rect 1119 3422 1123 3423
rect 1142 3422 1148 3423
rect 1159 3422 1163 3423
rect 1071 3417 1075 3418
rect 614 3415 620 3416
rect 614 3411 615 3415
rect 619 3411 620 3415
rect 614 3410 620 3411
rect 662 3415 668 3416
rect 662 3411 663 3415
rect 667 3411 668 3415
rect 662 3410 668 3411
rect 502 3400 508 3401
rect 502 3396 503 3400
rect 507 3396 508 3400
rect 502 3395 508 3396
rect 590 3400 596 3401
rect 590 3396 591 3400
rect 595 3396 596 3400
rect 590 3395 596 3396
rect 664 3392 666 3410
rect 680 3401 682 3417
rect 750 3415 756 3416
rect 750 3411 751 3415
rect 755 3411 756 3415
rect 750 3410 756 3411
rect 678 3400 684 3401
rect 678 3396 679 3400
rect 683 3396 684 3400
rect 678 3395 684 3396
rect 752 3392 754 3410
rect 768 3401 770 3417
rect 856 3401 858 3417
rect 926 3415 932 3416
rect 926 3411 927 3415
rect 931 3411 932 3415
rect 926 3410 932 3411
rect 766 3400 772 3401
rect 766 3396 767 3400
rect 771 3396 772 3400
rect 766 3395 772 3396
rect 854 3400 860 3401
rect 854 3396 855 3400
rect 859 3396 860 3400
rect 854 3395 860 3396
rect 928 3392 930 3410
rect 944 3401 946 3417
rect 1014 3415 1020 3416
rect 1014 3411 1015 3415
rect 1019 3411 1020 3415
rect 1014 3410 1020 3411
rect 942 3400 948 3401
rect 942 3396 943 3400
rect 947 3396 948 3400
rect 942 3395 948 3396
rect 1016 3392 1018 3410
rect 1032 3401 1034 3417
rect 1030 3400 1036 3401
rect 1030 3396 1031 3400
rect 1035 3396 1036 3400
rect 1030 3395 1036 3396
rect 1104 3392 1106 3422
rect 1119 3417 1123 3418
rect 1159 3417 1163 3418
rect 1207 3422 1211 3423
rect 1207 3417 1211 3418
rect 1303 3422 1307 3423
rect 1303 3417 1307 3418
rect 1767 3422 1771 3423
rect 1902 3422 1908 3423
rect 2014 3427 2020 3428
rect 2014 3423 2015 3427
rect 2019 3423 2020 3427
rect 2014 3422 2020 3423
rect 1767 3417 1771 3418
rect 1830 3417 1836 3418
rect 1120 3401 1122 3417
rect 1208 3401 1210 3417
rect 1258 3415 1264 3416
rect 1258 3411 1259 3415
rect 1263 3411 1264 3415
rect 1258 3410 1264 3411
rect 1278 3415 1284 3416
rect 1278 3411 1279 3415
rect 1283 3411 1284 3415
rect 1278 3410 1284 3411
rect 1118 3400 1124 3401
rect 1118 3396 1119 3400
rect 1123 3396 1124 3400
rect 1118 3395 1124 3396
rect 1206 3400 1212 3401
rect 1206 3396 1207 3400
rect 1211 3396 1212 3400
rect 1206 3395 1212 3396
rect 478 3391 484 3392
rect 478 3387 479 3391
rect 483 3387 484 3391
rect 478 3386 484 3387
rect 494 3391 500 3392
rect 494 3387 495 3391
rect 499 3387 500 3391
rect 494 3386 500 3387
rect 662 3391 668 3392
rect 662 3387 663 3391
rect 667 3387 668 3391
rect 662 3386 668 3387
rect 750 3391 756 3392
rect 750 3387 751 3391
rect 755 3387 756 3391
rect 750 3386 756 3387
rect 926 3391 932 3392
rect 926 3387 927 3391
rect 931 3387 932 3391
rect 926 3386 932 3387
rect 1014 3391 1020 3392
rect 1014 3387 1015 3391
rect 1019 3387 1020 3391
rect 1014 3386 1020 3387
rect 1102 3391 1108 3392
rect 1102 3387 1103 3391
rect 1107 3387 1108 3391
rect 1102 3386 1108 3387
rect 414 3381 420 3382
rect 110 3380 116 3381
rect 110 3376 111 3380
rect 115 3376 116 3380
rect 414 3377 415 3381
rect 419 3377 420 3381
rect 414 3376 420 3377
rect 110 3375 116 3376
rect 112 3355 114 3375
rect 416 3355 418 3376
rect 111 3354 115 3355
rect 111 3349 115 3350
rect 399 3354 403 3355
rect 399 3349 403 3350
rect 415 3354 419 3355
rect 415 3349 419 3350
rect 112 3333 114 3349
rect 110 3332 116 3333
rect 400 3332 402 3349
rect 110 3328 111 3332
rect 115 3328 116 3332
rect 110 3327 116 3328
rect 398 3331 404 3332
rect 398 3327 399 3331
rect 403 3327 404 3331
rect 398 3326 404 3327
rect 110 3315 116 3316
rect 110 3311 111 3315
rect 115 3311 116 3315
rect 110 3310 116 3311
rect 398 3312 404 3313
rect 112 3287 114 3310
rect 398 3308 399 3312
rect 403 3308 404 3312
rect 398 3307 404 3308
rect 400 3287 402 3307
rect 480 3296 482 3386
rect 502 3381 508 3382
rect 502 3377 503 3381
rect 507 3377 508 3381
rect 502 3376 508 3377
rect 590 3381 596 3382
rect 590 3377 591 3381
rect 595 3377 596 3381
rect 590 3376 596 3377
rect 678 3381 684 3382
rect 678 3377 679 3381
rect 683 3377 684 3381
rect 678 3376 684 3377
rect 766 3381 772 3382
rect 766 3377 767 3381
rect 771 3377 772 3381
rect 766 3376 772 3377
rect 854 3381 860 3382
rect 854 3377 855 3381
rect 859 3377 860 3381
rect 854 3376 860 3377
rect 942 3381 948 3382
rect 942 3377 943 3381
rect 947 3377 948 3381
rect 942 3376 948 3377
rect 1030 3381 1036 3382
rect 1030 3377 1031 3381
rect 1035 3377 1036 3381
rect 1030 3376 1036 3377
rect 1118 3381 1124 3382
rect 1118 3377 1119 3381
rect 1123 3377 1124 3381
rect 1118 3376 1124 3377
rect 1206 3381 1212 3382
rect 1206 3377 1207 3381
rect 1211 3377 1212 3381
rect 1206 3376 1212 3377
rect 504 3355 506 3376
rect 592 3355 594 3376
rect 680 3355 682 3376
rect 768 3355 770 3376
rect 856 3355 858 3376
rect 944 3355 946 3376
rect 1032 3355 1034 3376
rect 1120 3355 1122 3376
rect 1208 3355 1210 3376
rect 495 3354 499 3355
rect 495 3349 499 3350
rect 503 3354 507 3355
rect 503 3349 507 3350
rect 591 3354 595 3355
rect 591 3349 595 3350
rect 599 3354 603 3355
rect 599 3349 603 3350
rect 679 3354 683 3355
rect 679 3349 683 3350
rect 703 3354 707 3355
rect 703 3349 707 3350
rect 767 3354 771 3355
rect 767 3349 771 3350
rect 807 3354 811 3355
rect 807 3349 811 3350
rect 855 3354 859 3355
rect 855 3349 859 3350
rect 911 3354 915 3355
rect 911 3349 915 3350
rect 943 3354 947 3355
rect 943 3349 947 3350
rect 1015 3354 1019 3355
rect 1015 3349 1019 3350
rect 1031 3354 1035 3355
rect 1031 3349 1035 3350
rect 1119 3354 1123 3355
rect 1119 3349 1123 3350
rect 1207 3354 1211 3355
rect 1207 3349 1211 3350
rect 1223 3354 1227 3355
rect 1223 3349 1227 3350
rect 496 3332 498 3349
rect 600 3332 602 3349
rect 704 3332 706 3349
rect 808 3332 810 3349
rect 912 3332 914 3349
rect 1016 3332 1018 3349
rect 1120 3332 1122 3349
rect 1190 3347 1196 3348
rect 1190 3343 1191 3347
rect 1195 3343 1196 3347
rect 1190 3342 1196 3343
rect 494 3331 500 3332
rect 494 3327 495 3331
rect 499 3327 500 3331
rect 494 3326 500 3327
rect 598 3331 604 3332
rect 598 3327 599 3331
rect 603 3327 604 3331
rect 598 3326 604 3327
rect 702 3331 708 3332
rect 702 3327 703 3331
rect 707 3327 708 3331
rect 702 3326 708 3327
rect 806 3331 812 3332
rect 806 3327 807 3331
rect 811 3327 812 3331
rect 806 3326 812 3327
rect 910 3331 916 3332
rect 910 3327 911 3331
rect 915 3327 916 3331
rect 910 3326 916 3327
rect 1014 3331 1020 3332
rect 1014 3327 1015 3331
rect 1019 3327 1020 3331
rect 1014 3326 1020 3327
rect 1118 3331 1124 3332
rect 1118 3327 1119 3331
rect 1123 3327 1124 3331
rect 1118 3326 1124 3327
rect 1192 3324 1194 3342
rect 1224 3332 1226 3349
rect 1260 3348 1262 3410
rect 1280 3392 1282 3410
rect 1304 3401 1306 3417
rect 1302 3400 1308 3401
rect 1302 3396 1303 3400
rect 1307 3396 1308 3400
rect 1768 3398 1770 3417
rect 1806 3416 1812 3417
rect 1806 3412 1807 3416
rect 1811 3412 1812 3416
rect 1830 3413 1831 3417
rect 1835 3413 1836 3417
rect 1830 3412 1836 3413
rect 1942 3417 1948 3418
rect 1942 3413 1943 3417
rect 1947 3413 1948 3417
rect 1942 3412 1948 3413
rect 2078 3417 2084 3418
rect 2078 3413 2079 3417
rect 2083 3413 2084 3417
rect 2078 3412 2084 3413
rect 1806 3411 1812 3412
rect 1302 3395 1308 3396
rect 1766 3397 1772 3398
rect 1766 3393 1767 3397
rect 1771 3393 1772 3397
rect 1766 3392 1772 3393
rect 1278 3391 1284 3392
rect 1278 3387 1279 3391
rect 1283 3387 1284 3391
rect 1808 3387 1810 3411
rect 1832 3387 1834 3412
rect 1944 3387 1946 3412
rect 2080 3387 2082 3412
rect 1278 3386 1284 3387
rect 1807 3386 1811 3387
rect 1302 3381 1308 3382
rect 1807 3381 1811 3382
rect 1831 3386 1835 3387
rect 1831 3381 1835 3382
rect 1943 3386 1947 3387
rect 1943 3381 1947 3382
rect 1951 3386 1955 3387
rect 1951 3381 1955 3382
rect 2079 3386 2083 3387
rect 2079 3381 2083 3382
rect 2095 3386 2099 3387
rect 2095 3381 2099 3382
rect 1302 3377 1303 3381
rect 1307 3377 1308 3381
rect 1302 3376 1308 3377
rect 1766 3380 1772 3381
rect 1766 3376 1767 3380
rect 1771 3376 1772 3380
rect 1304 3355 1306 3376
rect 1766 3375 1772 3376
rect 1768 3355 1770 3375
rect 1808 3365 1810 3381
rect 1806 3364 1812 3365
rect 1832 3364 1834 3381
rect 1952 3364 1954 3381
rect 2096 3364 2098 3381
rect 1806 3360 1807 3364
rect 1811 3360 1812 3364
rect 1806 3359 1812 3360
rect 1830 3363 1836 3364
rect 1830 3359 1831 3363
rect 1835 3359 1836 3363
rect 1830 3358 1836 3359
rect 1950 3363 1956 3364
rect 1950 3359 1951 3363
rect 1955 3359 1956 3363
rect 1950 3358 1956 3359
rect 2094 3363 2100 3364
rect 2094 3359 2095 3363
rect 2099 3359 2100 3363
rect 2094 3358 2100 3359
rect 2168 3356 2170 3446
rect 2216 3437 2218 3453
rect 2352 3437 2354 3453
rect 2408 3452 2410 3486
rect 2726 3483 2727 3487
rect 2731 3483 2732 3487
rect 2726 3482 2732 3483
rect 2926 3487 2932 3488
rect 2926 3483 2927 3487
rect 2931 3483 2932 3487
rect 2926 3482 2932 3483
rect 3118 3487 3124 3488
rect 3118 3483 3119 3487
rect 3123 3483 3124 3487
rect 3118 3482 3124 3483
rect 3462 3483 3468 3484
rect 2454 3480 2460 3481
rect 2454 3476 2455 3480
rect 2459 3476 2460 3480
rect 2454 3475 2460 3476
rect 2654 3480 2660 3481
rect 2654 3476 2655 3480
rect 2659 3476 2660 3480
rect 2654 3475 2660 3476
rect 2456 3459 2458 3475
rect 2656 3459 2658 3475
rect 2728 3464 2730 3482
rect 2854 3480 2860 3481
rect 2854 3476 2855 3480
rect 2859 3476 2860 3480
rect 2854 3475 2860 3476
rect 2726 3463 2732 3464
rect 2726 3459 2727 3463
rect 2731 3459 2732 3463
rect 2856 3459 2858 3475
rect 2928 3464 2930 3482
rect 3046 3480 3052 3481
rect 3046 3476 3047 3480
rect 3051 3476 3052 3480
rect 3046 3475 3052 3476
rect 2926 3463 2932 3464
rect 2926 3459 2927 3463
rect 2931 3459 2932 3463
rect 3048 3459 3050 3475
rect 3120 3464 3122 3482
rect 3246 3480 3252 3481
rect 3246 3476 3247 3480
rect 3251 3476 3252 3480
rect 3462 3479 3463 3483
rect 3467 3479 3468 3483
rect 3462 3478 3468 3479
rect 3246 3475 3252 3476
rect 3118 3463 3124 3464
rect 3118 3459 3119 3463
rect 3123 3459 3124 3463
rect 3248 3459 3250 3475
rect 3464 3459 3466 3478
rect 2455 3458 2459 3459
rect 2455 3453 2459 3454
rect 2479 3458 2483 3459
rect 2479 3453 2483 3454
rect 2599 3458 2603 3459
rect 2599 3453 2603 3454
rect 2655 3458 2659 3459
rect 2655 3453 2659 3454
rect 2719 3458 2723 3459
rect 2726 3458 2732 3459
rect 2847 3458 2851 3459
rect 2719 3453 2723 3454
rect 2847 3453 2851 3454
rect 2855 3458 2859 3459
rect 2926 3458 2932 3459
rect 2975 3458 2979 3459
rect 2855 3453 2859 3454
rect 2975 3453 2979 3454
rect 3047 3458 3051 3459
rect 3118 3458 3124 3459
rect 3247 3458 3251 3459
rect 3047 3453 3051 3454
rect 3247 3453 3251 3454
rect 3463 3458 3467 3459
rect 3463 3453 3467 3454
rect 2406 3451 2412 3452
rect 2406 3447 2407 3451
rect 2411 3447 2412 3451
rect 2406 3446 2412 3447
rect 2480 3437 2482 3453
rect 2590 3451 2596 3452
rect 2590 3447 2591 3451
rect 2595 3447 2596 3451
rect 2590 3446 2596 3447
rect 2214 3436 2220 3437
rect 2214 3432 2215 3436
rect 2219 3432 2220 3436
rect 2214 3431 2220 3432
rect 2350 3436 2356 3437
rect 2350 3432 2351 3436
rect 2355 3432 2356 3436
rect 2350 3431 2356 3432
rect 2478 3436 2484 3437
rect 2478 3432 2479 3436
rect 2483 3432 2484 3436
rect 2478 3431 2484 3432
rect 2286 3427 2292 3428
rect 2286 3423 2287 3427
rect 2291 3423 2292 3427
rect 2286 3422 2292 3423
rect 2214 3417 2220 3418
rect 2214 3413 2215 3417
rect 2219 3413 2220 3417
rect 2214 3412 2220 3413
rect 2216 3387 2218 3412
rect 2215 3386 2219 3387
rect 2215 3381 2219 3382
rect 2239 3386 2243 3387
rect 2239 3381 2243 3382
rect 2240 3364 2242 3381
rect 2238 3363 2244 3364
rect 2238 3359 2239 3363
rect 2243 3359 2244 3363
rect 2238 3358 2244 3359
rect 2166 3355 2172 3356
rect 1303 3354 1307 3355
rect 1303 3349 1307 3350
rect 1327 3354 1331 3355
rect 1327 3349 1331 3350
rect 1767 3354 1771 3355
rect 1767 3349 1771 3350
rect 1902 3351 1908 3352
rect 1258 3347 1264 3348
rect 1258 3343 1259 3347
rect 1263 3343 1264 3347
rect 1258 3342 1264 3343
rect 1328 3332 1330 3349
rect 1768 3333 1770 3349
rect 1806 3347 1812 3348
rect 1806 3343 1807 3347
rect 1811 3343 1812 3347
rect 1902 3347 1903 3351
rect 1907 3347 1908 3351
rect 1902 3346 1908 3347
rect 2022 3351 2028 3352
rect 2022 3347 2023 3351
rect 2027 3347 2028 3351
rect 2166 3351 2167 3355
rect 2171 3351 2172 3355
rect 2166 3350 2172 3351
rect 2022 3346 2028 3347
rect 1806 3342 1812 3343
rect 1830 3344 1836 3345
rect 1766 3332 1772 3333
rect 1222 3331 1228 3332
rect 1222 3327 1223 3331
rect 1227 3327 1228 3331
rect 1222 3326 1228 3327
rect 1326 3331 1332 3332
rect 1326 3327 1327 3331
rect 1331 3327 1332 3331
rect 1766 3328 1767 3332
rect 1771 3328 1772 3332
rect 1766 3327 1772 3328
rect 1326 3326 1332 3327
rect 1190 3323 1196 3324
rect 486 3319 492 3320
rect 486 3315 487 3319
rect 491 3315 492 3319
rect 486 3314 492 3315
rect 566 3319 572 3320
rect 566 3315 567 3319
rect 571 3315 572 3319
rect 566 3314 572 3315
rect 670 3319 676 3320
rect 670 3315 671 3319
rect 675 3315 676 3319
rect 670 3314 676 3315
rect 774 3319 780 3320
rect 774 3315 775 3319
rect 779 3315 780 3319
rect 774 3314 780 3315
rect 878 3319 884 3320
rect 878 3315 879 3319
rect 883 3315 884 3319
rect 878 3314 884 3315
rect 982 3319 988 3320
rect 982 3315 983 3319
rect 987 3315 988 3319
rect 982 3314 988 3315
rect 1086 3319 1092 3320
rect 1086 3315 1087 3319
rect 1091 3315 1092 3319
rect 1190 3319 1191 3323
rect 1195 3319 1196 3323
rect 1190 3318 1196 3319
rect 1198 3323 1204 3324
rect 1198 3319 1199 3323
rect 1203 3319 1204 3323
rect 1198 3318 1204 3319
rect 1302 3323 1308 3324
rect 1302 3319 1303 3323
rect 1307 3319 1308 3323
rect 1302 3318 1308 3319
rect 1086 3314 1092 3315
rect 488 3296 490 3314
rect 494 3312 500 3313
rect 494 3308 495 3312
rect 499 3308 500 3312
rect 494 3307 500 3308
rect 478 3295 484 3296
rect 478 3291 479 3295
rect 483 3291 484 3295
rect 478 3290 484 3291
rect 486 3295 492 3296
rect 486 3291 487 3295
rect 491 3291 492 3295
rect 486 3290 492 3291
rect 496 3287 498 3307
rect 568 3296 570 3314
rect 598 3312 604 3313
rect 598 3308 599 3312
rect 603 3308 604 3312
rect 598 3307 604 3308
rect 566 3295 572 3296
rect 566 3291 567 3295
rect 571 3291 572 3295
rect 566 3290 572 3291
rect 600 3287 602 3307
rect 672 3296 674 3314
rect 702 3312 708 3313
rect 702 3308 703 3312
rect 707 3308 708 3312
rect 702 3307 708 3308
rect 670 3295 676 3296
rect 670 3291 671 3295
rect 675 3291 676 3295
rect 670 3290 676 3291
rect 704 3287 706 3307
rect 776 3296 778 3314
rect 806 3312 812 3313
rect 806 3308 807 3312
rect 811 3308 812 3312
rect 806 3307 812 3308
rect 774 3295 780 3296
rect 774 3291 775 3295
rect 779 3291 780 3295
rect 774 3290 780 3291
rect 808 3287 810 3307
rect 111 3286 115 3287
rect 111 3281 115 3282
rect 383 3286 387 3287
rect 383 3281 387 3282
rect 399 3286 403 3287
rect 399 3281 403 3282
rect 495 3286 499 3287
rect 495 3281 499 3282
rect 599 3286 603 3287
rect 599 3281 603 3282
rect 607 3286 611 3287
rect 607 3281 611 3282
rect 703 3286 707 3287
rect 703 3281 707 3282
rect 727 3286 731 3287
rect 727 3281 731 3282
rect 807 3286 811 3287
rect 807 3281 811 3282
rect 847 3286 851 3287
rect 847 3281 851 3282
rect 112 3262 114 3281
rect 384 3265 386 3281
rect 454 3279 460 3280
rect 454 3275 455 3279
rect 459 3275 460 3279
rect 454 3274 460 3275
rect 382 3264 388 3265
rect 110 3261 116 3262
rect 110 3257 111 3261
rect 115 3257 116 3261
rect 382 3260 383 3264
rect 387 3260 388 3264
rect 382 3259 388 3260
rect 110 3256 116 3257
rect 456 3256 458 3274
rect 496 3265 498 3281
rect 608 3265 610 3281
rect 694 3279 700 3280
rect 694 3275 695 3279
rect 699 3275 700 3279
rect 694 3274 700 3275
rect 494 3264 500 3265
rect 494 3260 495 3264
rect 499 3260 500 3264
rect 494 3259 500 3260
rect 606 3264 612 3265
rect 606 3260 607 3264
rect 611 3260 612 3264
rect 606 3259 612 3260
rect 696 3256 698 3274
rect 728 3265 730 3281
rect 848 3265 850 3281
rect 880 3280 882 3314
rect 910 3312 916 3313
rect 910 3308 911 3312
rect 915 3308 916 3312
rect 910 3307 916 3308
rect 912 3287 914 3307
rect 984 3296 986 3314
rect 1014 3312 1020 3313
rect 1014 3308 1015 3312
rect 1019 3308 1020 3312
rect 1014 3307 1020 3308
rect 982 3295 988 3296
rect 982 3291 983 3295
rect 987 3291 988 3295
rect 982 3290 988 3291
rect 1016 3287 1018 3307
rect 1088 3296 1090 3314
rect 1118 3312 1124 3313
rect 1118 3308 1119 3312
rect 1123 3308 1124 3312
rect 1118 3307 1124 3308
rect 1086 3295 1092 3296
rect 1086 3291 1087 3295
rect 1091 3291 1092 3295
rect 1086 3290 1092 3291
rect 1120 3287 1122 3307
rect 1200 3304 1202 3318
rect 1222 3312 1228 3313
rect 1222 3308 1223 3312
rect 1227 3308 1228 3312
rect 1222 3307 1228 3308
rect 1198 3303 1204 3304
rect 1198 3299 1199 3303
rect 1203 3299 1204 3303
rect 1198 3298 1204 3299
rect 1224 3287 1226 3307
rect 1304 3296 1306 3318
rect 1766 3315 1772 3316
rect 1808 3315 1810 3342
rect 1830 3340 1831 3344
rect 1835 3340 1836 3344
rect 1830 3339 1836 3340
rect 1832 3315 1834 3339
rect 1904 3328 1906 3346
rect 1950 3344 1956 3345
rect 1950 3340 1951 3344
rect 1955 3340 1956 3344
rect 1950 3339 1956 3340
rect 1894 3327 1900 3328
rect 1894 3323 1895 3327
rect 1899 3323 1900 3327
rect 1894 3322 1900 3323
rect 1902 3327 1908 3328
rect 1902 3323 1903 3327
rect 1907 3323 1908 3327
rect 1902 3322 1908 3323
rect 1326 3312 1332 3313
rect 1326 3308 1327 3312
rect 1331 3308 1332 3312
rect 1766 3311 1767 3315
rect 1771 3311 1772 3315
rect 1766 3310 1772 3311
rect 1807 3314 1811 3315
rect 1326 3307 1332 3308
rect 1302 3295 1308 3296
rect 1302 3291 1303 3295
rect 1307 3291 1308 3295
rect 1302 3290 1308 3291
rect 1328 3287 1330 3307
rect 1398 3295 1404 3296
rect 1398 3291 1399 3295
rect 1403 3291 1404 3295
rect 1398 3290 1404 3291
rect 911 3286 915 3287
rect 911 3281 915 3282
rect 967 3286 971 3287
rect 967 3281 971 3282
rect 1015 3286 1019 3287
rect 1015 3281 1019 3282
rect 1087 3286 1091 3287
rect 1087 3281 1091 3282
rect 1119 3286 1123 3287
rect 1119 3281 1123 3282
rect 1207 3286 1211 3287
rect 1207 3281 1211 3282
rect 1223 3286 1227 3287
rect 1223 3281 1227 3282
rect 1327 3286 1331 3287
rect 1327 3281 1331 3282
rect 1335 3286 1339 3287
rect 1335 3281 1339 3282
rect 878 3279 884 3280
rect 878 3275 879 3279
rect 883 3275 884 3279
rect 878 3274 884 3275
rect 968 3265 970 3281
rect 998 3279 1004 3280
rect 998 3275 999 3279
rect 1003 3275 1004 3279
rect 998 3274 1004 3275
rect 1038 3279 1044 3280
rect 1038 3275 1039 3279
rect 1043 3275 1044 3279
rect 1038 3274 1044 3275
rect 726 3264 732 3265
rect 726 3260 727 3264
rect 731 3260 732 3264
rect 726 3259 732 3260
rect 846 3264 852 3265
rect 846 3260 847 3264
rect 851 3260 852 3264
rect 846 3259 852 3260
rect 966 3264 972 3265
rect 966 3260 967 3264
rect 971 3260 972 3264
rect 966 3259 972 3260
rect 454 3255 460 3256
rect 454 3251 455 3255
rect 459 3251 460 3255
rect 454 3250 460 3251
rect 566 3255 572 3256
rect 566 3251 567 3255
rect 571 3251 572 3255
rect 566 3250 572 3251
rect 694 3255 700 3256
rect 694 3251 695 3255
rect 699 3251 700 3255
rect 694 3250 700 3251
rect 382 3245 388 3246
rect 110 3244 116 3245
rect 110 3240 111 3244
rect 115 3240 116 3244
rect 382 3241 383 3245
rect 387 3241 388 3245
rect 382 3240 388 3241
rect 494 3245 500 3246
rect 494 3241 495 3245
rect 499 3241 500 3245
rect 494 3240 500 3241
rect 110 3239 116 3240
rect 112 3219 114 3239
rect 384 3219 386 3240
rect 496 3219 498 3240
rect 111 3218 115 3219
rect 111 3213 115 3214
rect 303 3218 307 3219
rect 303 3213 307 3214
rect 383 3218 387 3219
rect 383 3213 387 3214
rect 423 3218 427 3219
rect 423 3213 427 3214
rect 495 3218 499 3219
rect 495 3213 499 3214
rect 543 3218 547 3219
rect 543 3213 547 3214
rect 112 3197 114 3213
rect 110 3196 116 3197
rect 304 3196 306 3213
rect 424 3196 426 3213
rect 544 3196 546 3213
rect 110 3192 111 3196
rect 115 3192 116 3196
rect 110 3191 116 3192
rect 302 3195 308 3196
rect 302 3191 303 3195
rect 307 3191 308 3195
rect 302 3190 308 3191
rect 422 3195 428 3196
rect 422 3191 423 3195
rect 427 3191 428 3195
rect 422 3190 428 3191
rect 542 3195 548 3196
rect 542 3191 543 3195
rect 547 3191 548 3195
rect 542 3190 548 3191
rect 374 3183 380 3184
rect 110 3179 116 3180
rect 110 3175 111 3179
rect 115 3175 116 3179
rect 374 3179 375 3183
rect 379 3179 380 3183
rect 374 3178 380 3179
rect 494 3183 500 3184
rect 494 3179 495 3183
rect 499 3179 500 3183
rect 494 3178 500 3179
rect 110 3174 116 3175
rect 302 3176 308 3177
rect 112 3143 114 3174
rect 302 3172 303 3176
rect 307 3172 308 3176
rect 302 3171 308 3172
rect 304 3143 306 3171
rect 376 3160 378 3178
rect 422 3176 428 3177
rect 422 3172 423 3176
rect 427 3172 428 3176
rect 422 3171 428 3172
rect 374 3159 380 3160
rect 374 3155 375 3159
rect 379 3155 380 3159
rect 374 3154 380 3155
rect 424 3143 426 3171
rect 111 3142 115 3143
rect 111 3137 115 3138
rect 175 3142 179 3143
rect 175 3137 179 3138
rect 303 3142 307 3143
rect 303 3137 307 3138
rect 319 3142 323 3143
rect 319 3137 323 3138
rect 423 3142 427 3143
rect 423 3137 427 3138
rect 471 3142 475 3143
rect 471 3137 475 3138
rect 112 3118 114 3137
rect 176 3121 178 3137
rect 246 3135 252 3136
rect 246 3131 247 3135
rect 251 3131 252 3135
rect 246 3130 252 3131
rect 174 3120 180 3121
rect 110 3117 116 3118
rect 110 3113 111 3117
rect 115 3113 116 3117
rect 174 3116 175 3120
rect 179 3116 180 3120
rect 174 3115 180 3116
rect 110 3112 116 3113
rect 248 3112 250 3130
rect 320 3121 322 3137
rect 472 3121 474 3137
rect 496 3136 498 3178
rect 542 3176 548 3177
rect 542 3172 543 3176
rect 547 3172 548 3176
rect 542 3171 548 3172
rect 544 3143 546 3171
rect 568 3160 570 3250
rect 606 3245 612 3246
rect 606 3241 607 3245
rect 611 3241 612 3245
rect 606 3240 612 3241
rect 726 3245 732 3246
rect 726 3241 727 3245
rect 731 3241 732 3245
rect 726 3240 732 3241
rect 846 3245 852 3246
rect 846 3241 847 3245
rect 851 3241 852 3245
rect 846 3240 852 3241
rect 966 3245 972 3246
rect 966 3241 967 3245
rect 971 3241 972 3245
rect 966 3240 972 3241
rect 608 3219 610 3240
rect 728 3219 730 3240
rect 848 3219 850 3240
rect 968 3219 970 3240
rect 607 3218 611 3219
rect 607 3213 611 3214
rect 671 3218 675 3219
rect 671 3213 675 3214
rect 727 3218 731 3219
rect 727 3213 731 3214
rect 799 3218 803 3219
rect 799 3213 803 3214
rect 847 3218 851 3219
rect 847 3213 851 3214
rect 927 3218 931 3219
rect 927 3213 931 3214
rect 967 3218 971 3219
rect 967 3213 971 3214
rect 672 3196 674 3213
rect 800 3196 802 3213
rect 928 3196 930 3213
rect 670 3195 676 3196
rect 670 3191 671 3195
rect 675 3191 676 3195
rect 670 3190 676 3191
rect 798 3195 804 3196
rect 798 3191 799 3195
rect 803 3191 804 3195
rect 798 3190 804 3191
rect 926 3195 932 3196
rect 926 3191 927 3195
rect 931 3191 932 3195
rect 926 3190 932 3191
rect 1000 3188 1002 3274
rect 1040 3256 1042 3274
rect 1088 3265 1090 3281
rect 1158 3279 1164 3280
rect 1158 3275 1159 3279
rect 1163 3275 1164 3279
rect 1158 3274 1164 3275
rect 1086 3264 1092 3265
rect 1086 3260 1087 3264
rect 1091 3260 1092 3264
rect 1086 3259 1092 3260
rect 1160 3256 1162 3274
rect 1208 3265 1210 3281
rect 1278 3279 1284 3280
rect 1278 3275 1279 3279
rect 1283 3275 1284 3279
rect 1278 3274 1284 3275
rect 1206 3264 1212 3265
rect 1206 3260 1207 3264
rect 1211 3260 1212 3264
rect 1206 3259 1212 3260
rect 1280 3256 1282 3274
rect 1336 3265 1338 3281
rect 1334 3264 1340 3265
rect 1334 3260 1335 3264
rect 1339 3260 1340 3264
rect 1334 3259 1340 3260
rect 1400 3256 1402 3290
rect 1768 3287 1770 3310
rect 1807 3309 1811 3310
rect 1831 3314 1835 3315
rect 1831 3309 1835 3310
rect 1808 3290 1810 3309
rect 1832 3293 1834 3309
rect 1830 3292 1836 3293
rect 1806 3289 1812 3290
rect 1767 3286 1771 3287
rect 1806 3285 1807 3289
rect 1811 3285 1812 3289
rect 1830 3288 1831 3292
rect 1835 3288 1836 3292
rect 1830 3287 1836 3288
rect 1806 3284 1812 3285
rect 1896 3284 1898 3322
rect 1952 3315 1954 3339
rect 2024 3328 2026 3346
rect 2094 3344 2100 3345
rect 2094 3340 2095 3344
rect 2099 3340 2100 3344
rect 2094 3339 2100 3340
rect 2238 3344 2244 3345
rect 2238 3340 2239 3344
rect 2243 3340 2244 3344
rect 2238 3339 2244 3340
rect 2022 3327 2028 3328
rect 2022 3323 2023 3327
rect 2027 3323 2028 3327
rect 2022 3322 2028 3323
rect 2096 3315 2098 3339
rect 2240 3315 2242 3339
rect 2288 3328 2290 3422
rect 2350 3417 2356 3418
rect 2350 3413 2351 3417
rect 2355 3413 2356 3417
rect 2350 3412 2356 3413
rect 2478 3417 2484 3418
rect 2478 3413 2479 3417
rect 2483 3413 2484 3417
rect 2478 3412 2484 3413
rect 2352 3387 2354 3412
rect 2480 3387 2482 3412
rect 2351 3386 2355 3387
rect 2351 3381 2355 3382
rect 2383 3386 2387 3387
rect 2383 3381 2387 3382
rect 2479 3386 2483 3387
rect 2479 3381 2483 3382
rect 2519 3386 2523 3387
rect 2519 3381 2523 3382
rect 2384 3364 2386 3381
rect 2520 3364 2522 3381
rect 2382 3363 2388 3364
rect 2382 3359 2383 3363
rect 2387 3359 2388 3363
rect 2382 3358 2388 3359
rect 2518 3363 2524 3364
rect 2518 3359 2519 3363
rect 2523 3359 2524 3363
rect 2518 3358 2524 3359
rect 2592 3356 2594 3446
rect 2600 3437 2602 3453
rect 2670 3451 2676 3452
rect 2670 3447 2671 3451
rect 2675 3447 2676 3451
rect 2670 3446 2676 3447
rect 2598 3436 2604 3437
rect 2598 3432 2599 3436
rect 2603 3432 2604 3436
rect 2598 3431 2604 3432
rect 2672 3428 2674 3446
rect 2720 3437 2722 3453
rect 2790 3451 2796 3452
rect 2790 3447 2791 3451
rect 2795 3447 2796 3451
rect 2790 3446 2796 3447
rect 2718 3436 2724 3437
rect 2718 3432 2719 3436
rect 2723 3432 2724 3436
rect 2718 3431 2724 3432
rect 2792 3428 2794 3446
rect 2848 3437 2850 3453
rect 2918 3451 2924 3452
rect 2918 3447 2919 3451
rect 2923 3447 2924 3451
rect 2918 3446 2924 3447
rect 2846 3436 2852 3437
rect 2846 3432 2847 3436
rect 2851 3432 2852 3436
rect 2846 3431 2852 3432
rect 2920 3428 2922 3446
rect 2976 3437 2978 3453
rect 2974 3436 2980 3437
rect 2974 3432 2975 3436
rect 2979 3432 2980 3436
rect 3464 3434 3466 3453
rect 2974 3431 2980 3432
rect 3462 3433 3468 3434
rect 3462 3429 3463 3433
rect 3467 3429 3468 3433
rect 3462 3428 3468 3429
rect 2670 3427 2676 3428
rect 2670 3423 2671 3427
rect 2675 3423 2676 3427
rect 2670 3422 2676 3423
rect 2790 3427 2796 3428
rect 2790 3423 2791 3427
rect 2795 3423 2796 3427
rect 2790 3422 2796 3423
rect 2918 3427 2924 3428
rect 2918 3423 2919 3427
rect 2923 3423 2924 3427
rect 2918 3422 2924 3423
rect 2598 3417 2604 3418
rect 2598 3413 2599 3417
rect 2603 3413 2604 3417
rect 2598 3412 2604 3413
rect 2718 3417 2724 3418
rect 2718 3413 2719 3417
rect 2723 3413 2724 3417
rect 2718 3412 2724 3413
rect 2846 3417 2852 3418
rect 2846 3413 2847 3417
rect 2851 3413 2852 3417
rect 2846 3412 2852 3413
rect 2974 3417 2980 3418
rect 2974 3413 2975 3417
rect 2979 3413 2980 3417
rect 2974 3412 2980 3413
rect 3462 3416 3468 3417
rect 3462 3412 3463 3416
rect 3467 3412 3468 3416
rect 2600 3387 2602 3412
rect 2720 3387 2722 3412
rect 2848 3387 2850 3412
rect 2976 3387 2978 3412
rect 3462 3411 3468 3412
rect 3464 3387 3466 3411
rect 2599 3386 2603 3387
rect 2599 3381 2603 3382
rect 2647 3386 2651 3387
rect 2647 3381 2651 3382
rect 2719 3386 2723 3387
rect 2719 3381 2723 3382
rect 2775 3386 2779 3387
rect 2775 3381 2779 3382
rect 2847 3386 2851 3387
rect 2847 3381 2851 3382
rect 2903 3386 2907 3387
rect 2903 3381 2907 3382
rect 2975 3386 2979 3387
rect 2975 3381 2979 3382
rect 3039 3386 3043 3387
rect 3039 3381 3043 3382
rect 3463 3386 3467 3387
rect 3463 3381 3467 3382
rect 2648 3364 2650 3381
rect 2776 3364 2778 3381
rect 2904 3364 2906 3381
rect 3040 3364 3042 3381
rect 3464 3365 3466 3381
rect 3462 3364 3468 3365
rect 2646 3363 2652 3364
rect 2646 3359 2647 3363
rect 2651 3359 2652 3363
rect 2646 3358 2652 3359
rect 2774 3363 2780 3364
rect 2774 3359 2775 3363
rect 2779 3359 2780 3363
rect 2774 3358 2780 3359
rect 2902 3363 2908 3364
rect 2902 3359 2903 3363
rect 2907 3359 2908 3363
rect 2902 3358 2908 3359
rect 3038 3363 3044 3364
rect 3038 3359 3039 3363
rect 3043 3359 3044 3363
rect 3462 3360 3463 3364
rect 3467 3360 3468 3364
rect 3462 3359 3468 3360
rect 3038 3358 3044 3359
rect 2590 3355 2596 3356
rect 2310 3351 2316 3352
rect 2310 3347 2311 3351
rect 2315 3347 2316 3351
rect 2310 3346 2316 3347
rect 2454 3351 2460 3352
rect 2454 3347 2455 3351
rect 2459 3347 2460 3351
rect 2590 3351 2591 3355
rect 2595 3351 2596 3355
rect 2590 3350 2596 3351
rect 2598 3355 2604 3356
rect 2598 3351 2599 3355
rect 2603 3351 2604 3355
rect 2598 3350 2604 3351
rect 2726 3355 2732 3356
rect 2726 3351 2727 3355
rect 2731 3351 2732 3355
rect 2982 3355 2988 3356
rect 2726 3350 2732 3351
rect 2974 3351 2980 3352
rect 2454 3346 2460 3347
rect 2312 3328 2314 3346
rect 2382 3344 2388 3345
rect 2382 3340 2383 3344
rect 2387 3340 2388 3344
rect 2382 3339 2388 3340
rect 2286 3327 2292 3328
rect 2286 3323 2287 3327
rect 2291 3323 2292 3327
rect 2286 3322 2292 3323
rect 2310 3327 2316 3328
rect 2310 3323 2311 3327
rect 2315 3323 2316 3327
rect 2310 3322 2316 3323
rect 2384 3315 2386 3339
rect 1951 3314 1955 3315
rect 1951 3309 1955 3310
rect 1975 3314 1979 3315
rect 1975 3309 1979 3310
rect 2095 3314 2099 3315
rect 2095 3309 2099 3310
rect 2151 3314 2155 3315
rect 2151 3309 2155 3310
rect 2239 3314 2243 3315
rect 2239 3309 2243 3310
rect 2335 3314 2339 3315
rect 2335 3309 2339 3310
rect 2383 3314 2387 3315
rect 2383 3309 2387 3310
rect 1910 3307 1916 3308
rect 1910 3303 1911 3307
rect 1915 3303 1916 3307
rect 1910 3302 1916 3303
rect 1912 3284 1914 3302
rect 1976 3293 1978 3309
rect 2054 3307 2060 3308
rect 2054 3303 2055 3307
rect 2059 3303 2060 3307
rect 2054 3302 2060 3303
rect 2102 3307 2108 3308
rect 2102 3303 2103 3307
rect 2107 3303 2108 3307
rect 2102 3302 2108 3303
rect 1974 3292 1980 3293
rect 1974 3288 1975 3292
rect 1979 3288 1980 3292
rect 1974 3287 1980 3288
rect 2056 3284 2058 3302
rect 1767 3281 1771 3282
rect 1894 3283 1900 3284
rect 1768 3262 1770 3281
rect 1894 3279 1895 3283
rect 1899 3279 1900 3283
rect 1894 3278 1900 3279
rect 1910 3283 1916 3284
rect 1910 3279 1911 3283
rect 1915 3279 1916 3283
rect 1910 3278 1916 3279
rect 2054 3283 2060 3284
rect 2054 3279 2055 3283
rect 2059 3279 2060 3283
rect 2054 3278 2060 3279
rect 1830 3273 1836 3274
rect 1806 3272 1812 3273
rect 1806 3268 1807 3272
rect 1811 3268 1812 3272
rect 1830 3269 1831 3273
rect 1835 3269 1836 3273
rect 1830 3268 1836 3269
rect 1974 3273 1980 3274
rect 1974 3269 1975 3273
rect 1979 3269 1980 3273
rect 1974 3268 1980 3269
rect 1806 3267 1812 3268
rect 1766 3261 1772 3262
rect 1766 3257 1767 3261
rect 1771 3257 1772 3261
rect 1766 3256 1772 3257
rect 1038 3255 1044 3256
rect 1038 3251 1039 3255
rect 1043 3251 1044 3255
rect 1038 3250 1044 3251
rect 1158 3255 1164 3256
rect 1158 3251 1159 3255
rect 1163 3251 1164 3255
rect 1158 3250 1164 3251
rect 1278 3255 1284 3256
rect 1278 3251 1279 3255
rect 1283 3251 1284 3255
rect 1278 3250 1284 3251
rect 1398 3255 1404 3256
rect 1398 3251 1399 3255
rect 1403 3251 1404 3255
rect 1398 3250 1404 3251
rect 1086 3245 1092 3246
rect 1086 3241 1087 3245
rect 1091 3241 1092 3245
rect 1086 3240 1092 3241
rect 1206 3245 1212 3246
rect 1206 3241 1207 3245
rect 1211 3241 1212 3245
rect 1206 3240 1212 3241
rect 1334 3245 1340 3246
rect 1334 3241 1335 3245
rect 1339 3241 1340 3245
rect 1334 3240 1340 3241
rect 1766 3244 1772 3245
rect 1766 3240 1767 3244
rect 1771 3240 1772 3244
rect 1808 3243 1810 3267
rect 1832 3243 1834 3268
rect 1976 3243 1978 3268
rect 1088 3219 1090 3240
rect 1208 3219 1210 3240
rect 1336 3219 1338 3240
rect 1766 3239 1772 3240
rect 1807 3242 1811 3243
rect 1768 3219 1770 3239
rect 1807 3237 1811 3238
rect 1831 3242 1835 3243
rect 1831 3237 1835 3238
rect 1975 3242 1979 3243
rect 1975 3237 1979 3238
rect 2031 3242 2035 3243
rect 2031 3237 2035 3238
rect 1808 3221 1810 3237
rect 1806 3220 1812 3221
rect 1832 3220 1834 3237
rect 2032 3220 2034 3237
rect 1055 3218 1059 3219
rect 1055 3213 1059 3214
rect 1087 3218 1091 3219
rect 1087 3213 1091 3214
rect 1175 3218 1179 3219
rect 1175 3213 1179 3214
rect 1207 3218 1211 3219
rect 1207 3213 1211 3214
rect 1303 3218 1307 3219
rect 1303 3213 1307 3214
rect 1335 3218 1339 3219
rect 1335 3213 1339 3214
rect 1431 3218 1435 3219
rect 1431 3213 1435 3214
rect 1767 3218 1771 3219
rect 1806 3216 1807 3220
rect 1811 3216 1812 3220
rect 1806 3215 1812 3216
rect 1830 3219 1836 3220
rect 1830 3215 1831 3219
rect 1835 3215 1836 3219
rect 1830 3214 1836 3215
rect 2030 3219 2036 3220
rect 2030 3215 2031 3219
rect 2035 3215 2036 3219
rect 2030 3214 2036 3215
rect 1767 3213 1771 3214
rect 1056 3196 1058 3213
rect 1176 3196 1178 3213
rect 1304 3196 1306 3213
rect 1432 3196 1434 3213
rect 1768 3197 1770 3213
rect 2104 3212 2106 3302
rect 2152 3293 2154 3309
rect 2336 3293 2338 3309
rect 2456 3308 2458 3346
rect 2518 3344 2524 3345
rect 2518 3340 2519 3344
rect 2523 3340 2524 3344
rect 2518 3339 2524 3340
rect 2520 3315 2522 3339
rect 2600 3328 2602 3350
rect 2646 3344 2652 3345
rect 2646 3340 2647 3344
rect 2651 3340 2652 3344
rect 2646 3339 2652 3340
rect 2598 3327 2604 3328
rect 2598 3323 2599 3327
rect 2603 3323 2604 3327
rect 2598 3322 2604 3323
rect 2648 3315 2650 3339
rect 2728 3328 2730 3350
rect 2974 3347 2975 3351
rect 2979 3347 2980 3351
rect 2982 3351 2983 3355
rect 2987 3351 2988 3355
rect 2982 3350 2988 3351
rect 2974 3346 2980 3347
rect 2774 3344 2780 3345
rect 2774 3340 2775 3344
rect 2779 3340 2780 3344
rect 2774 3339 2780 3340
rect 2902 3344 2908 3345
rect 2902 3340 2903 3344
rect 2907 3340 2908 3344
rect 2902 3339 2908 3340
rect 2726 3327 2732 3328
rect 2726 3323 2727 3327
rect 2731 3323 2732 3327
rect 2726 3322 2732 3323
rect 2776 3315 2778 3339
rect 2904 3315 2906 3339
rect 2976 3328 2978 3346
rect 2984 3336 2986 3350
rect 3462 3347 3468 3348
rect 3038 3344 3044 3345
rect 3038 3340 3039 3344
rect 3043 3340 3044 3344
rect 3462 3343 3463 3347
rect 3467 3343 3468 3347
rect 3462 3342 3468 3343
rect 3038 3339 3044 3340
rect 2982 3335 2988 3336
rect 2982 3331 2983 3335
rect 2987 3331 2988 3335
rect 2982 3330 2988 3331
rect 2974 3327 2980 3328
rect 2974 3323 2975 3327
rect 2979 3323 2980 3327
rect 2974 3322 2980 3323
rect 3040 3315 3042 3339
rect 3464 3315 3466 3342
rect 2511 3314 2515 3315
rect 2511 3309 2515 3310
rect 2519 3314 2523 3315
rect 2519 3309 2523 3310
rect 2647 3314 2651 3315
rect 2647 3309 2651 3310
rect 2679 3314 2683 3315
rect 2679 3309 2683 3310
rect 2775 3314 2779 3315
rect 2775 3309 2779 3310
rect 2831 3314 2835 3315
rect 2831 3309 2835 3310
rect 2903 3314 2907 3315
rect 2903 3309 2907 3310
rect 2975 3314 2979 3315
rect 2975 3309 2979 3310
rect 3039 3314 3043 3315
rect 3039 3309 3043 3310
rect 3111 3314 3115 3315
rect 3111 3309 3115 3310
rect 3247 3314 3251 3315
rect 3247 3309 3251 3310
rect 3367 3314 3371 3315
rect 3367 3309 3371 3310
rect 3463 3314 3467 3315
rect 3463 3309 3467 3310
rect 2414 3307 2420 3308
rect 2414 3303 2415 3307
rect 2419 3303 2420 3307
rect 2414 3302 2420 3303
rect 2454 3307 2460 3308
rect 2454 3303 2455 3307
rect 2459 3303 2460 3307
rect 2454 3302 2460 3303
rect 2150 3292 2156 3293
rect 2150 3288 2151 3292
rect 2155 3288 2156 3292
rect 2150 3287 2156 3288
rect 2334 3292 2340 3293
rect 2334 3288 2335 3292
rect 2339 3288 2340 3292
rect 2334 3287 2340 3288
rect 2416 3284 2418 3302
rect 2512 3293 2514 3309
rect 2680 3293 2682 3309
rect 2750 3307 2756 3308
rect 2750 3303 2751 3307
rect 2755 3303 2756 3307
rect 2750 3302 2756 3303
rect 2510 3292 2516 3293
rect 2510 3288 2511 3292
rect 2515 3288 2516 3292
rect 2510 3287 2516 3288
rect 2678 3292 2684 3293
rect 2678 3288 2679 3292
rect 2683 3288 2684 3292
rect 2678 3287 2684 3288
rect 2752 3284 2754 3302
rect 2832 3293 2834 3309
rect 2976 3293 2978 3309
rect 3054 3307 3060 3308
rect 3054 3303 3055 3307
rect 3059 3303 3060 3307
rect 3054 3302 3060 3303
rect 2830 3292 2836 3293
rect 2830 3288 2831 3292
rect 2835 3288 2836 3292
rect 2830 3287 2836 3288
rect 2974 3292 2980 3293
rect 2974 3288 2975 3292
rect 2979 3288 2980 3292
rect 2974 3287 2980 3288
rect 3056 3284 3058 3302
rect 3112 3293 3114 3309
rect 3248 3293 3250 3309
rect 3326 3307 3332 3308
rect 3326 3303 3327 3307
rect 3331 3303 3332 3307
rect 3326 3302 3332 3303
rect 3110 3292 3116 3293
rect 3110 3288 3111 3292
rect 3115 3288 3116 3292
rect 3110 3287 3116 3288
rect 3246 3292 3252 3293
rect 3246 3288 3247 3292
rect 3251 3288 3252 3292
rect 3246 3287 3252 3288
rect 3328 3284 3330 3302
rect 3368 3293 3370 3309
rect 3438 3307 3444 3308
rect 3438 3303 3439 3307
rect 3443 3303 3444 3307
rect 3438 3302 3444 3303
rect 3366 3292 3372 3293
rect 3366 3288 3367 3292
rect 3371 3288 3372 3292
rect 3366 3287 3372 3288
rect 2302 3283 2308 3284
rect 2302 3279 2303 3283
rect 2307 3279 2308 3283
rect 2302 3278 2308 3279
rect 2414 3283 2420 3284
rect 2414 3279 2415 3283
rect 2419 3279 2420 3283
rect 2414 3278 2420 3279
rect 2750 3283 2756 3284
rect 2750 3279 2751 3283
rect 2755 3279 2756 3283
rect 2750 3278 2756 3279
rect 3054 3283 3060 3284
rect 3054 3279 3055 3283
rect 3059 3279 3060 3283
rect 3054 3278 3060 3279
rect 3326 3283 3332 3284
rect 3326 3279 3327 3283
rect 3331 3279 3332 3283
rect 3326 3278 3332 3279
rect 2150 3273 2156 3274
rect 2150 3269 2151 3273
rect 2155 3269 2156 3273
rect 2150 3268 2156 3269
rect 2152 3243 2154 3268
rect 2151 3242 2155 3243
rect 2151 3237 2155 3238
rect 2247 3242 2251 3243
rect 2247 3237 2251 3238
rect 2248 3220 2250 3237
rect 2246 3219 2252 3220
rect 2246 3215 2247 3219
rect 2251 3215 2252 3219
rect 2246 3214 2252 3215
rect 2102 3211 2108 3212
rect 2102 3207 2103 3211
rect 2107 3207 2108 3211
rect 2102 3206 2108 3207
rect 1806 3203 1812 3204
rect 1806 3199 1807 3203
rect 1811 3199 1812 3203
rect 1806 3198 1812 3199
rect 1830 3200 1836 3201
rect 1766 3196 1772 3197
rect 1054 3195 1060 3196
rect 1054 3191 1055 3195
rect 1059 3191 1060 3195
rect 1054 3190 1060 3191
rect 1174 3195 1180 3196
rect 1174 3191 1175 3195
rect 1179 3191 1180 3195
rect 1174 3190 1180 3191
rect 1302 3195 1308 3196
rect 1302 3191 1303 3195
rect 1307 3191 1308 3195
rect 1302 3190 1308 3191
rect 1430 3195 1436 3196
rect 1430 3191 1431 3195
rect 1435 3191 1436 3195
rect 1766 3192 1767 3196
rect 1771 3192 1772 3196
rect 1766 3191 1772 3192
rect 1430 3190 1436 3191
rect 758 3187 764 3188
rect 614 3183 620 3184
rect 614 3179 615 3183
rect 619 3179 620 3183
rect 614 3178 620 3179
rect 742 3183 748 3184
rect 742 3179 743 3183
rect 747 3179 748 3183
rect 758 3183 759 3187
rect 763 3183 764 3187
rect 758 3182 764 3183
rect 998 3187 1004 3188
rect 998 3183 999 3187
rect 1003 3183 1004 3187
rect 998 3182 1004 3183
rect 1006 3187 1012 3188
rect 1006 3183 1007 3187
rect 1011 3183 1012 3187
rect 1006 3182 1012 3183
rect 1134 3187 1140 3188
rect 1134 3183 1135 3187
rect 1139 3183 1140 3187
rect 1382 3187 1388 3188
rect 1134 3182 1140 3183
rect 1374 3183 1380 3184
rect 742 3178 748 3179
rect 616 3160 618 3178
rect 670 3176 676 3177
rect 670 3172 671 3176
rect 675 3172 676 3176
rect 670 3171 676 3172
rect 566 3159 572 3160
rect 566 3155 567 3159
rect 571 3155 572 3159
rect 566 3154 572 3155
rect 614 3159 620 3160
rect 614 3155 615 3159
rect 619 3155 620 3159
rect 614 3154 620 3155
rect 672 3143 674 3171
rect 744 3160 746 3178
rect 760 3168 762 3182
rect 798 3176 804 3177
rect 798 3172 799 3176
rect 803 3172 804 3176
rect 798 3171 804 3172
rect 926 3176 932 3177
rect 926 3172 927 3176
rect 931 3172 932 3176
rect 926 3171 932 3172
rect 758 3167 764 3168
rect 758 3163 759 3167
rect 763 3163 764 3167
rect 758 3162 764 3163
rect 742 3159 748 3160
rect 742 3155 743 3159
rect 747 3155 748 3159
rect 742 3154 748 3155
rect 800 3143 802 3171
rect 928 3143 930 3171
rect 1008 3160 1010 3182
rect 1054 3176 1060 3177
rect 1054 3172 1055 3176
rect 1059 3172 1060 3176
rect 1054 3171 1060 3172
rect 1006 3159 1012 3160
rect 1006 3155 1007 3159
rect 1011 3155 1012 3159
rect 1006 3154 1012 3155
rect 1056 3143 1058 3171
rect 1136 3160 1138 3182
rect 1374 3179 1375 3183
rect 1379 3179 1380 3183
rect 1382 3183 1383 3187
rect 1387 3183 1388 3187
rect 1382 3182 1388 3183
rect 1374 3178 1380 3179
rect 1174 3176 1180 3177
rect 1174 3172 1175 3176
rect 1179 3172 1180 3176
rect 1174 3171 1180 3172
rect 1302 3176 1308 3177
rect 1302 3172 1303 3176
rect 1307 3172 1308 3176
rect 1302 3171 1308 3172
rect 1134 3159 1140 3160
rect 1134 3155 1135 3159
rect 1139 3155 1140 3159
rect 1134 3154 1140 3155
rect 1176 3143 1178 3171
rect 1270 3159 1276 3160
rect 1270 3155 1271 3159
rect 1275 3155 1276 3159
rect 1270 3154 1276 3155
rect 543 3142 547 3143
rect 543 3137 547 3138
rect 623 3142 627 3143
rect 623 3137 627 3138
rect 671 3142 675 3143
rect 671 3137 675 3138
rect 775 3142 779 3143
rect 775 3137 779 3138
rect 799 3142 803 3143
rect 799 3137 803 3138
rect 919 3142 923 3143
rect 919 3137 923 3138
rect 927 3142 931 3143
rect 927 3137 931 3138
rect 1055 3142 1059 3143
rect 1055 3137 1059 3138
rect 1063 3142 1067 3143
rect 1063 3137 1067 3138
rect 1175 3142 1179 3143
rect 1175 3137 1179 3138
rect 1199 3142 1203 3143
rect 1199 3137 1203 3138
rect 494 3135 500 3136
rect 494 3131 495 3135
rect 499 3131 500 3135
rect 494 3130 500 3131
rect 624 3121 626 3137
rect 694 3135 700 3136
rect 694 3131 695 3135
rect 699 3131 700 3135
rect 694 3130 700 3131
rect 318 3120 324 3121
rect 318 3116 319 3120
rect 323 3116 324 3120
rect 318 3115 324 3116
rect 470 3120 476 3121
rect 470 3116 471 3120
rect 475 3116 476 3120
rect 470 3115 476 3116
rect 622 3120 628 3121
rect 622 3116 623 3120
rect 627 3116 628 3120
rect 622 3115 628 3116
rect 696 3112 698 3130
rect 776 3121 778 3137
rect 920 3121 922 3137
rect 990 3135 996 3136
rect 990 3131 991 3135
rect 995 3131 996 3135
rect 990 3130 996 3131
rect 774 3120 780 3121
rect 774 3116 775 3120
rect 779 3116 780 3120
rect 774 3115 780 3116
rect 918 3120 924 3121
rect 918 3116 919 3120
rect 923 3116 924 3120
rect 918 3115 924 3116
rect 992 3112 994 3130
rect 1064 3121 1066 3137
rect 1134 3135 1140 3136
rect 1134 3131 1135 3135
rect 1139 3131 1140 3135
rect 1134 3130 1140 3131
rect 1062 3120 1068 3121
rect 1062 3116 1063 3120
rect 1067 3116 1068 3120
rect 1062 3115 1068 3116
rect 1136 3112 1138 3130
rect 1200 3121 1202 3137
rect 1198 3120 1204 3121
rect 1198 3116 1199 3120
rect 1203 3116 1204 3120
rect 1198 3115 1204 3116
rect 1272 3112 1274 3154
rect 1304 3143 1306 3171
rect 1376 3160 1378 3178
rect 1384 3168 1386 3182
rect 1766 3179 1772 3180
rect 1808 3179 1810 3198
rect 1830 3196 1831 3200
rect 1835 3196 1836 3200
rect 1830 3195 1836 3196
rect 2030 3200 2036 3201
rect 2030 3196 2031 3200
rect 2035 3196 2036 3200
rect 2030 3195 2036 3196
rect 2246 3200 2252 3201
rect 2246 3196 2247 3200
rect 2251 3196 2252 3200
rect 2246 3195 2252 3196
rect 1832 3179 1834 3195
rect 1902 3183 1908 3184
rect 1902 3179 1903 3183
rect 1907 3179 1908 3183
rect 2032 3179 2034 3195
rect 2248 3179 2250 3195
rect 2304 3184 2306 3278
rect 2334 3273 2340 3274
rect 2334 3269 2335 3273
rect 2339 3269 2340 3273
rect 2334 3268 2340 3269
rect 2510 3273 2516 3274
rect 2510 3269 2511 3273
rect 2515 3269 2516 3273
rect 2510 3268 2516 3269
rect 2678 3273 2684 3274
rect 2678 3269 2679 3273
rect 2683 3269 2684 3273
rect 2678 3268 2684 3269
rect 2830 3273 2836 3274
rect 2830 3269 2831 3273
rect 2835 3269 2836 3273
rect 2830 3268 2836 3269
rect 2974 3273 2980 3274
rect 2974 3269 2975 3273
rect 2979 3269 2980 3273
rect 2974 3268 2980 3269
rect 3110 3273 3116 3274
rect 3110 3269 3111 3273
rect 3115 3269 3116 3273
rect 3110 3268 3116 3269
rect 3246 3273 3252 3274
rect 3246 3269 3247 3273
rect 3251 3269 3252 3273
rect 3246 3268 3252 3269
rect 3366 3273 3372 3274
rect 3366 3269 3367 3273
rect 3371 3269 3372 3273
rect 3366 3268 3372 3269
rect 2336 3243 2338 3268
rect 2512 3243 2514 3268
rect 2680 3243 2682 3268
rect 2832 3243 2834 3268
rect 2976 3243 2978 3268
rect 3112 3243 3114 3268
rect 3248 3243 3250 3268
rect 3368 3243 3370 3268
rect 2335 3242 2339 3243
rect 2335 3237 2339 3238
rect 2455 3242 2459 3243
rect 2455 3237 2459 3238
rect 2511 3242 2515 3243
rect 2511 3237 2515 3238
rect 2655 3242 2659 3243
rect 2655 3237 2659 3238
rect 2679 3242 2683 3243
rect 2679 3237 2683 3238
rect 2831 3242 2835 3243
rect 2831 3237 2835 3238
rect 2839 3242 2843 3243
rect 2839 3237 2843 3238
rect 2975 3242 2979 3243
rect 2975 3237 2979 3238
rect 3023 3242 3027 3243
rect 3023 3237 3027 3238
rect 3111 3242 3115 3243
rect 3111 3237 3115 3238
rect 3207 3242 3211 3243
rect 3207 3237 3211 3238
rect 3247 3242 3251 3243
rect 3247 3237 3251 3238
rect 3367 3242 3371 3243
rect 3367 3237 3371 3238
rect 2456 3220 2458 3237
rect 2656 3220 2658 3237
rect 2840 3220 2842 3237
rect 3024 3220 3026 3237
rect 3208 3220 3210 3237
rect 3368 3220 3370 3237
rect 2454 3219 2460 3220
rect 2454 3215 2455 3219
rect 2459 3215 2460 3219
rect 2454 3214 2460 3215
rect 2654 3219 2660 3220
rect 2654 3215 2655 3219
rect 2659 3215 2660 3219
rect 2654 3214 2660 3215
rect 2838 3219 2844 3220
rect 2838 3215 2839 3219
rect 2843 3215 2844 3219
rect 2838 3214 2844 3215
rect 3022 3219 3028 3220
rect 3022 3215 3023 3219
rect 3027 3215 3028 3219
rect 3022 3214 3028 3215
rect 3206 3219 3212 3220
rect 3206 3215 3207 3219
rect 3211 3215 3212 3219
rect 3206 3214 3212 3215
rect 3366 3219 3372 3220
rect 3366 3215 3367 3219
rect 3371 3215 3372 3219
rect 3366 3214 3372 3215
rect 3440 3212 3442 3302
rect 3464 3290 3466 3309
rect 3462 3289 3468 3290
rect 3462 3285 3463 3289
rect 3467 3285 3468 3289
rect 3462 3284 3468 3285
rect 3462 3272 3468 3273
rect 3462 3268 3463 3272
rect 3467 3268 3468 3272
rect 3462 3267 3468 3268
rect 3464 3243 3466 3267
rect 3463 3242 3467 3243
rect 3463 3237 3467 3238
rect 3464 3221 3466 3237
rect 3462 3220 3468 3221
rect 3462 3216 3463 3220
rect 3467 3216 3468 3220
rect 3462 3215 3468 3216
rect 3438 3211 3444 3212
rect 2318 3207 2324 3208
rect 2318 3203 2319 3207
rect 2323 3203 2324 3207
rect 2318 3202 2324 3203
rect 2726 3207 2732 3208
rect 2726 3203 2727 3207
rect 2731 3203 2732 3207
rect 2726 3202 2732 3203
rect 2910 3207 2916 3208
rect 2910 3203 2911 3207
rect 2915 3203 2916 3207
rect 2910 3202 2916 3203
rect 3094 3207 3100 3208
rect 3094 3203 3095 3207
rect 3099 3203 3100 3207
rect 3438 3207 3439 3211
rect 3443 3207 3444 3211
rect 3438 3206 3444 3207
rect 3094 3202 3100 3203
rect 3462 3203 3468 3204
rect 2320 3184 2322 3202
rect 2454 3200 2460 3201
rect 2454 3196 2455 3200
rect 2459 3196 2460 3200
rect 2454 3195 2460 3196
rect 2654 3200 2660 3201
rect 2654 3196 2655 3200
rect 2659 3196 2660 3200
rect 2654 3195 2660 3196
rect 2302 3183 2308 3184
rect 2302 3179 2303 3183
rect 2307 3179 2308 3183
rect 1430 3176 1436 3177
rect 1430 3172 1431 3176
rect 1435 3172 1436 3176
rect 1766 3175 1767 3179
rect 1771 3175 1772 3179
rect 1766 3174 1772 3175
rect 1807 3178 1811 3179
rect 1430 3171 1436 3172
rect 1382 3167 1388 3168
rect 1382 3163 1383 3167
rect 1387 3163 1388 3167
rect 1382 3162 1388 3163
rect 1374 3159 1380 3160
rect 1374 3155 1375 3159
rect 1379 3155 1380 3159
rect 1374 3154 1380 3155
rect 1432 3143 1434 3171
rect 1768 3143 1770 3174
rect 1807 3173 1811 3174
rect 1831 3178 1835 3179
rect 1831 3173 1835 3174
rect 1839 3178 1843 3179
rect 1902 3178 1908 3179
rect 2031 3178 2035 3179
rect 1839 3173 1843 3174
rect 1808 3154 1810 3173
rect 1840 3157 1842 3173
rect 1838 3156 1844 3157
rect 1806 3153 1812 3154
rect 1806 3149 1807 3153
rect 1811 3149 1812 3153
rect 1838 3152 1839 3156
rect 1843 3152 1844 3156
rect 1838 3151 1844 3152
rect 1806 3148 1812 3149
rect 1904 3148 1906 3178
rect 2031 3173 2035 3174
rect 2223 3178 2227 3179
rect 2223 3173 2227 3174
rect 2247 3178 2251 3179
rect 2302 3178 2308 3179
rect 2318 3183 2324 3184
rect 2318 3179 2319 3183
rect 2323 3179 2324 3183
rect 2456 3179 2458 3195
rect 2646 3183 2652 3184
rect 2646 3179 2647 3183
rect 2651 3179 2652 3183
rect 2656 3179 2658 3195
rect 2728 3184 2730 3202
rect 2838 3200 2844 3201
rect 2838 3196 2839 3200
rect 2843 3196 2844 3200
rect 2838 3195 2844 3196
rect 2726 3183 2732 3184
rect 2726 3179 2727 3183
rect 2731 3179 2732 3183
rect 2840 3179 2842 3195
rect 2912 3184 2914 3202
rect 3022 3200 3028 3201
rect 3022 3196 3023 3200
rect 3027 3196 3028 3200
rect 3022 3195 3028 3196
rect 3062 3195 3068 3196
rect 2910 3183 2916 3184
rect 2910 3179 2911 3183
rect 2915 3179 2916 3183
rect 3024 3179 3026 3195
rect 3062 3191 3063 3195
rect 3067 3191 3068 3195
rect 3062 3190 3068 3191
rect 2318 3178 2324 3179
rect 2407 3178 2411 3179
rect 2247 3173 2251 3174
rect 2407 3173 2411 3174
rect 2455 3178 2459 3179
rect 2455 3173 2459 3174
rect 2575 3178 2579 3179
rect 2646 3178 2652 3179
rect 2655 3178 2659 3179
rect 2726 3178 2732 3179
rect 2735 3178 2739 3179
rect 2575 3173 2579 3174
rect 1918 3171 1924 3172
rect 1918 3167 1919 3171
rect 1923 3167 1924 3171
rect 1918 3166 1924 3167
rect 1920 3148 1922 3166
rect 2032 3157 2034 3173
rect 2110 3171 2116 3172
rect 2110 3167 2111 3171
rect 2115 3167 2116 3171
rect 2110 3166 2116 3167
rect 2030 3156 2036 3157
rect 2030 3152 2031 3156
rect 2035 3152 2036 3156
rect 2030 3151 2036 3152
rect 2112 3148 2114 3166
rect 2224 3157 2226 3173
rect 2254 3171 2260 3172
rect 2254 3167 2255 3171
rect 2259 3167 2260 3171
rect 2254 3166 2260 3167
rect 2222 3156 2228 3157
rect 2222 3152 2223 3156
rect 2227 3152 2228 3156
rect 2222 3151 2228 3152
rect 1902 3147 1908 3148
rect 1902 3143 1903 3147
rect 1907 3143 1908 3147
rect 1303 3142 1307 3143
rect 1303 3137 1307 3138
rect 1343 3142 1347 3143
rect 1343 3137 1347 3138
rect 1431 3142 1435 3143
rect 1431 3137 1435 3138
rect 1487 3142 1491 3143
rect 1487 3137 1491 3138
rect 1767 3142 1771 3143
rect 1902 3142 1908 3143
rect 1918 3147 1924 3148
rect 1918 3143 1919 3147
rect 1923 3143 1924 3147
rect 1918 3142 1924 3143
rect 2110 3147 2116 3148
rect 2110 3143 2111 3147
rect 2115 3143 2116 3147
rect 2110 3142 2116 3143
rect 1767 3137 1771 3138
rect 1838 3137 1844 3138
rect 1344 3121 1346 3137
rect 1422 3135 1428 3136
rect 1422 3131 1423 3135
rect 1427 3131 1428 3135
rect 1422 3130 1428 3131
rect 1342 3120 1348 3121
rect 1342 3116 1343 3120
rect 1347 3116 1348 3120
rect 1342 3115 1348 3116
rect 1424 3112 1426 3130
rect 1488 3121 1490 3137
rect 1582 3135 1588 3136
rect 1582 3131 1583 3135
rect 1587 3131 1588 3135
rect 1582 3130 1588 3131
rect 1486 3120 1492 3121
rect 1486 3116 1487 3120
rect 1491 3116 1492 3120
rect 1486 3115 1492 3116
rect 246 3111 252 3112
rect 246 3107 247 3111
rect 251 3107 252 3111
rect 246 3106 252 3107
rect 390 3111 396 3112
rect 390 3107 391 3111
rect 395 3107 396 3111
rect 390 3106 396 3107
rect 694 3111 700 3112
rect 694 3107 695 3111
rect 699 3107 700 3111
rect 694 3106 700 3107
rect 990 3111 996 3112
rect 990 3107 991 3111
rect 995 3107 996 3111
rect 990 3106 996 3107
rect 1134 3111 1140 3112
rect 1134 3107 1135 3111
rect 1139 3107 1140 3111
rect 1134 3106 1140 3107
rect 1270 3111 1276 3112
rect 1270 3107 1271 3111
rect 1275 3107 1276 3111
rect 1270 3106 1276 3107
rect 1422 3111 1428 3112
rect 1422 3107 1423 3111
rect 1427 3107 1428 3111
rect 1422 3106 1428 3107
rect 174 3101 180 3102
rect 110 3100 116 3101
rect 110 3096 111 3100
rect 115 3096 116 3100
rect 174 3097 175 3101
rect 179 3097 180 3101
rect 174 3096 180 3097
rect 318 3101 324 3102
rect 318 3097 319 3101
rect 323 3097 324 3101
rect 318 3096 324 3097
rect 110 3095 116 3096
rect 112 3071 114 3095
rect 176 3071 178 3096
rect 320 3071 322 3096
rect 111 3070 115 3071
rect 111 3065 115 3066
rect 135 3070 139 3071
rect 135 3065 139 3066
rect 175 3070 179 3071
rect 175 3065 179 3066
rect 263 3070 267 3071
rect 263 3065 267 3066
rect 319 3070 323 3071
rect 319 3065 323 3066
rect 112 3049 114 3065
rect 110 3048 116 3049
rect 136 3048 138 3065
rect 264 3048 266 3065
rect 110 3044 111 3048
rect 115 3044 116 3048
rect 110 3043 116 3044
rect 134 3047 140 3048
rect 134 3043 135 3047
rect 139 3043 140 3047
rect 134 3042 140 3043
rect 262 3047 268 3048
rect 262 3043 263 3047
rect 267 3043 268 3047
rect 262 3042 268 3043
rect 206 3035 212 3036
rect 110 3031 116 3032
rect 110 3027 111 3031
rect 115 3027 116 3031
rect 206 3031 207 3035
rect 211 3031 212 3035
rect 206 3030 212 3031
rect 334 3035 340 3036
rect 334 3031 335 3035
rect 339 3031 340 3035
rect 334 3030 340 3031
rect 110 3026 116 3027
rect 134 3028 140 3029
rect 112 3003 114 3026
rect 134 3024 135 3028
rect 139 3024 140 3028
rect 134 3023 140 3024
rect 136 3003 138 3023
rect 208 3012 210 3030
rect 262 3028 268 3029
rect 262 3024 263 3028
rect 267 3024 268 3028
rect 262 3023 268 3024
rect 206 3011 212 3012
rect 206 3007 207 3011
rect 211 3007 212 3011
rect 206 3006 212 3007
rect 264 3003 266 3023
rect 111 3002 115 3003
rect 111 2997 115 2998
rect 135 3002 139 3003
rect 135 2997 139 2998
rect 263 3002 267 3003
rect 263 2997 267 2998
rect 327 3002 331 3003
rect 327 2997 331 2998
rect 112 2978 114 2997
rect 136 2981 138 2997
rect 328 2981 330 2997
rect 336 2996 338 3030
rect 392 3012 394 3106
rect 470 3101 476 3102
rect 470 3097 471 3101
rect 475 3097 476 3101
rect 470 3096 476 3097
rect 622 3101 628 3102
rect 622 3097 623 3101
rect 627 3097 628 3101
rect 622 3096 628 3097
rect 774 3101 780 3102
rect 774 3097 775 3101
rect 779 3097 780 3101
rect 774 3096 780 3097
rect 918 3101 924 3102
rect 918 3097 919 3101
rect 923 3097 924 3101
rect 918 3096 924 3097
rect 1062 3101 1068 3102
rect 1062 3097 1063 3101
rect 1067 3097 1068 3101
rect 1062 3096 1068 3097
rect 1198 3101 1204 3102
rect 1198 3097 1199 3101
rect 1203 3097 1204 3101
rect 1198 3096 1204 3097
rect 1342 3101 1348 3102
rect 1342 3097 1343 3101
rect 1347 3097 1348 3101
rect 1342 3096 1348 3097
rect 1486 3101 1492 3102
rect 1486 3097 1487 3101
rect 1491 3097 1492 3101
rect 1486 3096 1492 3097
rect 472 3071 474 3096
rect 624 3071 626 3096
rect 776 3071 778 3096
rect 920 3071 922 3096
rect 1064 3071 1066 3096
rect 1200 3071 1202 3096
rect 1344 3071 1346 3096
rect 1488 3071 1490 3096
rect 431 3070 435 3071
rect 431 3065 435 3066
rect 471 3070 475 3071
rect 471 3065 475 3066
rect 607 3070 611 3071
rect 607 3065 611 3066
rect 623 3070 627 3071
rect 623 3065 627 3066
rect 775 3070 779 3071
rect 775 3065 779 3066
rect 791 3070 795 3071
rect 791 3065 795 3066
rect 919 3070 923 3071
rect 919 3065 923 3066
rect 967 3070 971 3071
rect 967 3065 971 3066
rect 1063 3070 1067 3071
rect 1063 3065 1067 3066
rect 1143 3070 1147 3071
rect 1143 3065 1147 3066
rect 1199 3070 1203 3071
rect 1199 3065 1203 3066
rect 1327 3070 1331 3071
rect 1327 3065 1331 3066
rect 1343 3070 1347 3071
rect 1343 3065 1347 3066
rect 1487 3070 1491 3071
rect 1487 3065 1491 3066
rect 1511 3070 1515 3071
rect 1511 3065 1515 3066
rect 432 3048 434 3065
rect 608 3048 610 3065
rect 792 3048 794 3065
rect 968 3048 970 3065
rect 1144 3048 1146 3065
rect 1328 3048 1330 3065
rect 1512 3048 1514 3065
rect 430 3047 436 3048
rect 430 3043 431 3047
rect 435 3043 436 3047
rect 430 3042 436 3043
rect 606 3047 612 3048
rect 606 3043 607 3047
rect 611 3043 612 3047
rect 606 3042 612 3043
rect 790 3047 796 3048
rect 790 3043 791 3047
rect 795 3043 796 3047
rect 790 3042 796 3043
rect 966 3047 972 3048
rect 966 3043 967 3047
rect 971 3043 972 3047
rect 966 3042 972 3043
rect 1142 3047 1148 3048
rect 1142 3043 1143 3047
rect 1147 3043 1148 3047
rect 1142 3042 1148 3043
rect 1326 3047 1332 3048
rect 1326 3043 1327 3047
rect 1331 3043 1332 3047
rect 1326 3042 1332 3043
rect 1510 3047 1516 3048
rect 1510 3043 1511 3047
rect 1515 3043 1516 3047
rect 1510 3042 1516 3043
rect 1584 3040 1586 3130
rect 1768 3118 1770 3137
rect 1806 3136 1812 3137
rect 1806 3132 1807 3136
rect 1811 3132 1812 3136
rect 1838 3133 1839 3137
rect 1843 3133 1844 3137
rect 1838 3132 1844 3133
rect 2030 3137 2036 3138
rect 2030 3133 2031 3137
rect 2035 3133 2036 3137
rect 2030 3132 2036 3133
rect 2222 3137 2228 3138
rect 2222 3133 2223 3137
rect 2227 3133 2228 3137
rect 2222 3132 2228 3133
rect 1806 3131 1812 3132
rect 1766 3117 1772 3118
rect 1766 3113 1767 3117
rect 1771 3113 1772 3117
rect 1766 3112 1772 3113
rect 1808 3111 1810 3131
rect 1840 3111 1842 3132
rect 2032 3111 2034 3132
rect 2224 3111 2226 3132
rect 1807 3110 1811 3111
rect 1807 3105 1811 3106
rect 1839 3110 1843 3111
rect 1839 3105 1843 3106
rect 1935 3110 1939 3111
rect 1935 3105 1939 3106
rect 2031 3110 2035 3111
rect 2031 3105 2035 3106
rect 2055 3110 2059 3111
rect 2055 3105 2059 3106
rect 2175 3110 2179 3111
rect 2175 3105 2179 3106
rect 2223 3110 2227 3111
rect 2223 3105 2227 3106
rect 1766 3100 1772 3101
rect 1766 3096 1767 3100
rect 1771 3096 1772 3100
rect 1766 3095 1772 3096
rect 1768 3071 1770 3095
rect 1808 3089 1810 3105
rect 1806 3088 1812 3089
rect 1936 3088 1938 3105
rect 2056 3088 2058 3105
rect 2176 3088 2178 3105
rect 1806 3084 1807 3088
rect 1811 3084 1812 3088
rect 1806 3083 1812 3084
rect 1934 3087 1940 3088
rect 1934 3083 1935 3087
rect 1939 3083 1940 3087
rect 1934 3082 1940 3083
rect 2054 3087 2060 3088
rect 2054 3083 2055 3087
rect 2059 3083 2060 3087
rect 2054 3082 2060 3083
rect 2174 3087 2180 3088
rect 2174 3083 2175 3087
rect 2179 3083 2180 3087
rect 2174 3082 2180 3083
rect 2256 3080 2258 3166
rect 2408 3157 2410 3173
rect 2576 3157 2578 3173
rect 2406 3156 2412 3157
rect 2406 3152 2407 3156
rect 2411 3152 2412 3156
rect 2406 3151 2412 3152
rect 2574 3156 2580 3157
rect 2574 3152 2575 3156
rect 2579 3152 2580 3156
rect 2574 3151 2580 3152
rect 2648 3148 2650 3178
rect 2655 3173 2659 3174
rect 2735 3173 2739 3174
rect 2839 3178 2843 3179
rect 2839 3173 2843 3174
rect 2879 3178 2883 3179
rect 2910 3178 2916 3179
rect 3007 3178 3011 3179
rect 2879 3173 2883 3174
rect 3007 3173 3011 3174
rect 3023 3178 3027 3179
rect 3023 3173 3027 3174
rect 2736 3157 2738 3173
rect 2814 3171 2820 3172
rect 2814 3167 2815 3171
rect 2819 3167 2820 3171
rect 2814 3166 2820 3167
rect 2734 3156 2740 3157
rect 2734 3152 2735 3156
rect 2739 3152 2740 3156
rect 2734 3151 2740 3152
rect 2816 3148 2818 3166
rect 2880 3157 2882 3173
rect 2974 3171 2980 3172
rect 2974 3167 2975 3171
rect 2979 3167 2980 3171
rect 2974 3166 2980 3167
rect 2878 3156 2884 3157
rect 2878 3152 2879 3156
rect 2883 3152 2884 3156
rect 2878 3151 2884 3152
rect 2478 3147 2484 3148
rect 2478 3143 2479 3147
rect 2483 3143 2484 3147
rect 2478 3142 2484 3143
rect 2646 3147 2652 3148
rect 2646 3143 2647 3147
rect 2651 3143 2652 3147
rect 2646 3142 2652 3143
rect 2814 3147 2820 3148
rect 2814 3143 2815 3147
rect 2819 3143 2820 3147
rect 2814 3142 2820 3143
rect 2406 3137 2412 3138
rect 2406 3133 2407 3137
rect 2411 3133 2412 3137
rect 2406 3132 2412 3133
rect 2408 3111 2410 3132
rect 2303 3110 2307 3111
rect 2303 3105 2307 3106
rect 2407 3110 2411 3111
rect 2407 3105 2411 3106
rect 2431 3110 2435 3111
rect 2431 3105 2435 3106
rect 2304 3088 2306 3105
rect 2432 3088 2434 3105
rect 2302 3087 2308 3088
rect 2302 3083 2303 3087
rect 2307 3083 2308 3087
rect 2302 3082 2308 3083
rect 2430 3087 2436 3088
rect 2430 3083 2431 3087
rect 2435 3083 2436 3087
rect 2430 3082 2436 3083
rect 2254 3079 2260 3080
rect 2006 3075 2012 3076
rect 1806 3071 1812 3072
rect 1767 3070 1771 3071
rect 1806 3067 1807 3071
rect 1811 3067 1812 3071
rect 2006 3071 2007 3075
rect 2011 3071 2012 3075
rect 2006 3070 2012 3071
rect 2126 3075 2132 3076
rect 2126 3071 2127 3075
rect 2131 3071 2132 3075
rect 2254 3075 2255 3079
rect 2259 3075 2260 3079
rect 2414 3079 2420 3080
rect 2254 3074 2260 3075
rect 2374 3075 2380 3076
rect 2126 3070 2132 3071
rect 2374 3071 2375 3075
rect 2379 3071 2380 3075
rect 2414 3075 2415 3079
rect 2419 3075 2420 3079
rect 2414 3074 2420 3075
rect 2374 3070 2380 3071
rect 1806 3066 1812 3067
rect 1934 3068 1940 3069
rect 1767 3065 1771 3066
rect 1768 3049 1770 3065
rect 1766 3048 1772 3049
rect 1766 3044 1767 3048
rect 1771 3044 1772 3048
rect 1766 3043 1772 3044
rect 754 3039 760 3040
rect 502 3035 508 3036
rect 502 3031 503 3035
rect 507 3031 508 3035
rect 502 3030 508 3031
rect 678 3035 684 3036
rect 678 3031 679 3035
rect 683 3031 684 3035
rect 754 3035 755 3039
rect 759 3035 760 3039
rect 1582 3039 1588 3040
rect 1808 3039 1810 3066
rect 1934 3064 1935 3068
rect 1939 3064 1940 3068
rect 1934 3063 1940 3064
rect 1936 3039 1938 3063
rect 2008 3052 2010 3070
rect 2054 3068 2060 3069
rect 2054 3064 2055 3068
rect 2059 3064 2060 3068
rect 2054 3063 2060 3064
rect 1990 3051 1996 3052
rect 1990 3047 1991 3051
rect 1995 3047 1996 3051
rect 1990 3046 1996 3047
rect 2006 3051 2012 3052
rect 2006 3047 2007 3051
rect 2011 3047 2012 3051
rect 2006 3046 2012 3047
rect 754 3034 760 3035
rect 1038 3035 1044 3036
rect 678 3030 684 3031
rect 430 3028 436 3029
rect 430 3024 431 3028
rect 435 3024 436 3028
rect 430 3023 436 3024
rect 390 3011 396 3012
rect 390 3007 391 3011
rect 395 3007 396 3011
rect 390 3006 396 3007
rect 432 3003 434 3023
rect 504 3012 506 3030
rect 606 3028 612 3029
rect 606 3024 607 3028
rect 611 3024 612 3028
rect 606 3023 612 3024
rect 502 3011 508 3012
rect 502 3007 503 3011
rect 507 3007 508 3011
rect 502 3006 508 3007
rect 608 3003 610 3023
rect 680 3012 682 3030
rect 756 3020 758 3034
rect 1038 3031 1039 3035
rect 1043 3031 1044 3035
rect 1038 3030 1044 3031
rect 1214 3035 1220 3036
rect 1214 3031 1215 3035
rect 1219 3031 1220 3035
rect 1214 3030 1220 3031
rect 1398 3035 1404 3036
rect 1398 3031 1399 3035
rect 1403 3031 1404 3035
rect 1582 3035 1583 3039
rect 1587 3035 1588 3039
rect 1582 3034 1588 3035
rect 1807 3038 1811 3039
rect 1807 3033 1811 3034
rect 1935 3038 1939 3039
rect 1935 3033 1939 3034
rect 1398 3030 1404 3031
rect 1766 3031 1772 3032
rect 790 3028 796 3029
rect 790 3024 791 3028
rect 795 3024 796 3028
rect 790 3023 796 3024
rect 966 3028 972 3029
rect 966 3024 967 3028
rect 971 3024 972 3028
rect 966 3023 972 3024
rect 754 3019 760 3020
rect 754 3015 755 3019
rect 759 3015 760 3019
rect 754 3014 760 3015
rect 678 3011 684 3012
rect 678 3007 679 3011
rect 683 3007 684 3011
rect 678 3006 684 3007
rect 792 3003 794 3023
rect 968 3003 970 3023
rect 1040 3012 1042 3030
rect 1142 3028 1148 3029
rect 1142 3024 1143 3028
rect 1147 3024 1148 3028
rect 1142 3023 1148 3024
rect 998 3011 1004 3012
rect 998 3007 999 3011
rect 1003 3007 1004 3011
rect 998 3006 1004 3007
rect 1038 3011 1044 3012
rect 1038 3007 1039 3011
rect 1043 3007 1044 3011
rect 1038 3006 1044 3007
rect 431 3002 435 3003
rect 431 2997 435 2998
rect 535 3002 539 3003
rect 535 2997 539 2998
rect 607 3002 611 3003
rect 607 2997 611 2998
rect 735 3002 739 3003
rect 735 2997 739 2998
rect 791 3002 795 3003
rect 791 2997 795 2998
rect 927 3002 931 3003
rect 927 2997 931 2998
rect 967 3002 971 3003
rect 967 2997 971 2998
rect 334 2995 340 2996
rect 334 2991 335 2995
rect 339 2991 340 2995
rect 334 2990 340 2991
rect 398 2995 404 2996
rect 398 2991 399 2995
rect 403 2991 404 2995
rect 398 2990 404 2991
rect 134 2980 140 2981
rect 110 2977 116 2978
rect 110 2973 111 2977
rect 115 2973 116 2977
rect 134 2976 135 2980
rect 139 2976 140 2980
rect 134 2975 140 2976
rect 326 2980 332 2981
rect 326 2976 327 2980
rect 331 2976 332 2980
rect 326 2975 332 2976
rect 110 2972 116 2973
rect 400 2972 402 2990
rect 536 2981 538 2997
rect 710 2995 716 2996
rect 710 2991 711 2995
rect 715 2991 716 2995
rect 710 2990 716 2991
rect 534 2980 540 2981
rect 534 2976 535 2980
rect 539 2976 540 2980
rect 534 2975 540 2976
rect 712 2972 714 2990
rect 736 2981 738 2997
rect 928 2981 930 2997
rect 734 2980 740 2981
rect 734 2976 735 2980
rect 739 2976 740 2980
rect 734 2975 740 2976
rect 926 2980 932 2981
rect 926 2976 927 2980
rect 931 2976 932 2980
rect 926 2975 932 2976
rect 1000 2972 1002 3006
rect 1144 3003 1146 3023
rect 1216 3012 1218 3030
rect 1326 3028 1332 3029
rect 1326 3024 1327 3028
rect 1331 3024 1332 3028
rect 1326 3023 1332 3024
rect 1214 3011 1220 3012
rect 1214 3007 1215 3011
rect 1219 3007 1220 3011
rect 1214 3006 1220 3007
rect 1328 3003 1330 3023
rect 1400 3012 1402 3030
rect 1510 3028 1516 3029
rect 1510 3024 1511 3028
rect 1515 3024 1516 3028
rect 1766 3027 1767 3031
rect 1771 3027 1772 3031
rect 1766 3026 1772 3027
rect 1510 3023 1516 3024
rect 1398 3011 1404 3012
rect 1398 3007 1399 3011
rect 1403 3007 1404 3011
rect 1398 3006 1404 3007
rect 1512 3003 1514 3023
rect 1768 3003 1770 3026
rect 1808 3014 1810 3033
rect 1806 3013 1812 3014
rect 1806 3009 1807 3013
rect 1811 3009 1812 3013
rect 1806 3008 1812 3009
rect 1992 3008 1994 3046
rect 2056 3039 2058 3063
rect 2128 3052 2130 3070
rect 2174 3068 2180 3069
rect 2174 3064 2175 3068
rect 2179 3064 2180 3068
rect 2174 3063 2180 3064
rect 2302 3068 2308 3069
rect 2302 3064 2303 3068
rect 2307 3064 2308 3068
rect 2302 3063 2308 3064
rect 2126 3051 2132 3052
rect 2126 3047 2127 3051
rect 2131 3047 2132 3051
rect 2126 3046 2132 3047
rect 2176 3039 2178 3063
rect 2304 3039 2306 3063
rect 2023 3038 2027 3039
rect 2023 3033 2027 3034
rect 2055 3038 2059 3039
rect 2055 3033 2059 3034
rect 2127 3038 2131 3039
rect 2127 3033 2131 3034
rect 2175 3038 2179 3039
rect 2175 3033 2179 3034
rect 2231 3038 2235 3039
rect 2231 3033 2235 3034
rect 2303 3038 2307 3039
rect 2303 3033 2307 3034
rect 2335 3038 2339 3039
rect 2335 3033 2339 3034
rect 2024 3017 2026 3033
rect 2128 3017 2130 3033
rect 2134 3031 2140 3032
rect 2134 3027 2135 3031
rect 2139 3027 2140 3031
rect 2134 3026 2140 3027
rect 2198 3031 2204 3032
rect 2198 3027 2199 3031
rect 2203 3027 2204 3031
rect 2198 3026 2204 3027
rect 2022 3016 2028 3017
rect 2022 3012 2023 3016
rect 2027 3012 2028 3016
rect 2022 3011 2028 3012
rect 2126 3016 2132 3017
rect 2126 3012 2127 3016
rect 2131 3012 2132 3016
rect 2126 3011 2132 3012
rect 1990 3007 1996 3008
rect 1990 3003 1991 3007
rect 1995 3003 1996 3007
rect 1103 3002 1107 3003
rect 1103 2997 1107 2998
rect 1143 3002 1147 3003
rect 1143 2997 1147 2998
rect 1279 3002 1283 3003
rect 1279 2997 1283 2998
rect 1327 3002 1331 3003
rect 1327 2997 1331 2998
rect 1447 3002 1451 3003
rect 1447 2997 1451 2998
rect 1511 3002 1515 3003
rect 1511 2997 1515 2998
rect 1623 3002 1627 3003
rect 1623 2997 1627 2998
rect 1767 3002 1771 3003
rect 1990 3002 1996 3003
rect 1767 2997 1771 2998
rect 2022 2997 2028 2998
rect 1006 2995 1012 2996
rect 1006 2991 1007 2995
rect 1011 2991 1012 2995
rect 1006 2990 1012 2991
rect 1008 2972 1010 2990
rect 1104 2981 1106 2997
rect 1280 2981 1282 2997
rect 1410 2995 1416 2996
rect 1410 2991 1411 2995
rect 1415 2991 1416 2995
rect 1410 2990 1416 2991
rect 1102 2980 1108 2981
rect 1102 2976 1103 2980
rect 1107 2976 1108 2980
rect 1102 2975 1108 2976
rect 1278 2980 1284 2981
rect 1278 2976 1279 2980
rect 1283 2976 1284 2980
rect 1278 2975 1284 2976
rect 1412 2972 1414 2990
rect 1448 2981 1450 2997
rect 1554 2995 1560 2996
rect 1554 2991 1555 2995
rect 1559 2991 1560 2995
rect 1554 2990 1560 2991
rect 1446 2980 1452 2981
rect 1446 2976 1447 2980
rect 1451 2976 1452 2980
rect 1446 2975 1452 2976
rect 1556 2972 1558 2990
rect 1624 2981 1626 2997
rect 1662 2995 1668 2996
rect 1662 2991 1663 2995
rect 1667 2991 1668 2995
rect 1662 2990 1668 2991
rect 1622 2980 1628 2981
rect 1622 2976 1623 2980
rect 1627 2976 1628 2980
rect 1622 2975 1628 2976
rect 198 2971 204 2972
rect 198 2967 199 2971
rect 203 2967 204 2971
rect 198 2966 204 2967
rect 398 2971 404 2972
rect 398 2967 399 2971
rect 403 2967 404 2971
rect 398 2966 404 2967
rect 710 2971 716 2972
rect 710 2967 711 2971
rect 715 2967 716 2971
rect 710 2966 716 2967
rect 998 2971 1004 2972
rect 998 2967 999 2971
rect 1003 2967 1004 2971
rect 998 2966 1004 2967
rect 1006 2971 1012 2972
rect 1006 2967 1007 2971
rect 1011 2967 1012 2971
rect 1006 2966 1012 2967
rect 1410 2971 1416 2972
rect 1410 2967 1411 2971
rect 1415 2967 1416 2971
rect 1410 2966 1416 2967
rect 1554 2971 1560 2972
rect 1554 2967 1555 2971
rect 1559 2967 1560 2971
rect 1554 2966 1560 2967
rect 134 2961 140 2962
rect 110 2960 116 2961
rect 110 2956 111 2960
rect 115 2956 116 2960
rect 134 2957 135 2961
rect 139 2957 140 2961
rect 134 2956 140 2957
rect 110 2955 116 2956
rect 112 2931 114 2955
rect 136 2931 138 2956
rect 111 2930 115 2931
rect 111 2925 115 2926
rect 135 2930 139 2931
rect 135 2925 139 2926
rect 112 2909 114 2925
rect 110 2908 116 2909
rect 136 2908 138 2925
rect 110 2904 111 2908
rect 115 2904 116 2908
rect 110 2903 116 2904
rect 134 2907 140 2908
rect 134 2903 135 2907
rect 139 2903 140 2907
rect 134 2902 140 2903
rect 110 2891 116 2892
rect 110 2887 111 2891
rect 115 2887 116 2891
rect 110 2886 116 2887
rect 134 2888 140 2889
rect 112 2863 114 2886
rect 134 2884 135 2888
rect 139 2884 140 2888
rect 134 2883 140 2884
rect 136 2863 138 2883
rect 200 2872 202 2966
rect 326 2961 332 2962
rect 326 2957 327 2961
rect 331 2957 332 2961
rect 326 2956 332 2957
rect 534 2961 540 2962
rect 534 2957 535 2961
rect 539 2957 540 2961
rect 534 2956 540 2957
rect 734 2961 740 2962
rect 734 2957 735 2961
rect 739 2957 740 2961
rect 734 2956 740 2957
rect 926 2961 932 2962
rect 926 2957 927 2961
rect 931 2957 932 2961
rect 926 2956 932 2957
rect 1102 2961 1108 2962
rect 1102 2957 1103 2961
rect 1107 2957 1108 2961
rect 1102 2956 1108 2957
rect 1278 2961 1284 2962
rect 1278 2957 1279 2961
rect 1283 2957 1284 2961
rect 1278 2956 1284 2957
rect 1446 2961 1452 2962
rect 1446 2957 1447 2961
rect 1451 2957 1452 2961
rect 1446 2956 1452 2957
rect 1622 2961 1628 2962
rect 1622 2957 1623 2961
rect 1627 2957 1628 2961
rect 1622 2956 1628 2957
rect 328 2931 330 2956
rect 536 2931 538 2956
rect 736 2931 738 2956
rect 928 2931 930 2956
rect 1104 2931 1106 2956
rect 1280 2931 1282 2956
rect 1448 2931 1450 2956
rect 1624 2931 1626 2956
rect 263 2930 267 2931
rect 263 2925 267 2926
rect 327 2930 331 2931
rect 327 2925 331 2926
rect 431 2930 435 2931
rect 431 2925 435 2926
rect 535 2930 539 2931
rect 535 2925 539 2926
rect 607 2930 611 2931
rect 607 2925 611 2926
rect 735 2930 739 2931
rect 735 2925 739 2926
rect 783 2930 787 2931
rect 783 2925 787 2926
rect 927 2930 931 2931
rect 927 2925 931 2926
rect 951 2930 955 2931
rect 951 2925 955 2926
rect 1103 2930 1107 2931
rect 1103 2925 1107 2926
rect 1111 2930 1115 2931
rect 1111 2925 1115 2926
rect 1271 2930 1275 2931
rect 1271 2925 1275 2926
rect 1279 2930 1283 2931
rect 1279 2925 1283 2926
rect 1431 2930 1435 2931
rect 1431 2925 1435 2926
rect 1447 2930 1451 2931
rect 1447 2925 1451 2926
rect 1591 2930 1595 2931
rect 1591 2925 1595 2926
rect 1623 2930 1627 2931
rect 1623 2925 1627 2926
rect 264 2908 266 2925
rect 432 2908 434 2925
rect 608 2908 610 2925
rect 784 2908 786 2925
rect 952 2908 954 2925
rect 1112 2908 1114 2925
rect 1272 2908 1274 2925
rect 1432 2908 1434 2925
rect 1592 2908 1594 2925
rect 262 2907 268 2908
rect 262 2903 263 2907
rect 267 2903 268 2907
rect 262 2902 268 2903
rect 430 2907 436 2908
rect 430 2903 431 2907
rect 435 2903 436 2907
rect 430 2902 436 2903
rect 606 2907 612 2908
rect 606 2903 607 2907
rect 611 2903 612 2907
rect 606 2902 612 2903
rect 782 2907 788 2908
rect 782 2903 783 2907
rect 787 2903 788 2907
rect 782 2902 788 2903
rect 950 2907 956 2908
rect 950 2903 951 2907
rect 955 2903 956 2907
rect 950 2902 956 2903
rect 1110 2907 1116 2908
rect 1110 2903 1111 2907
rect 1115 2903 1116 2907
rect 1110 2902 1116 2903
rect 1270 2907 1276 2908
rect 1270 2903 1271 2907
rect 1275 2903 1276 2907
rect 1270 2902 1276 2903
rect 1430 2907 1436 2908
rect 1430 2903 1431 2907
rect 1435 2903 1436 2907
rect 1430 2902 1436 2903
rect 1590 2907 1596 2908
rect 1590 2903 1591 2907
rect 1595 2903 1596 2907
rect 1590 2902 1596 2903
rect 1664 2900 1666 2990
rect 1768 2978 1770 2997
rect 1806 2996 1812 2997
rect 1806 2992 1807 2996
rect 1811 2992 1812 2996
rect 2022 2993 2023 2997
rect 2027 2993 2028 2997
rect 2022 2992 2028 2993
rect 2126 2997 2132 2998
rect 2126 2993 2127 2997
rect 2131 2993 2132 2997
rect 2126 2992 2132 2993
rect 1806 2991 1812 2992
rect 1766 2977 1772 2978
rect 1766 2973 1767 2977
rect 1771 2973 1772 2977
rect 1808 2975 1810 2991
rect 2024 2975 2026 2992
rect 2128 2975 2130 2992
rect 1766 2972 1772 2973
rect 1807 2974 1811 2975
rect 1807 2969 1811 2970
rect 2023 2974 2027 2975
rect 2023 2969 2027 2970
rect 2055 2974 2059 2975
rect 2055 2969 2059 2970
rect 2127 2974 2131 2975
rect 2127 2969 2131 2970
rect 1766 2960 1772 2961
rect 1766 2956 1767 2960
rect 1771 2956 1772 2960
rect 1766 2955 1772 2956
rect 1768 2931 1770 2955
rect 1808 2953 1810 2969
rect 1806 2952 1812 2953
rect 2056 2952 2058 2969
rect 2136 2952 2138 3026
rect 2200 3008 2202 3026
rect 2232 3017 2234 3033
rect 2336 3017 2338 3033
rect 2376 3032 2378 3070
rect 2416 3052 2418 3074
rect 2430 3068 2436 3069
rect 2430 3064 2431 3068
rect 2435 3064 2436 3068
rect 2430 3063 2436 3064
rect 2414 3051 2420 3052
rect 2414 3047 2415 3051
rect 2419 3047 2420 3051
rect 2414 3046 2420 3047
rect 2432 3039 2434 3063
rect 2480 3052 2482 3142
rect 2574 3137 2580 3138
rect 2574 3133 2575 3137
rect 2579 3133 2580 3137
rect 2574 3132 2580 3133
rect 2734 3137 2740 3138
rect 2734 3133 2735 3137
rect 2739 3133 2740 3137
rect 2734 3132 2740 3133
rect 2878 3137 2884 3138
rect 2878 3133 2879 3137
rect 2883 3133 2884 3137
rect 2878 3132 2884 3133
rect 2576 3111 2578 3132
rect 2736 3111 2738 3132
rect 2880 3111 2882 3132
rect 2567 3110 2571 3111
rect 2567 3105 2571 3106
rect 2575 3110 2579 3111
rect 2575 3105 2579 3106
rect 2719 3110 2723 3111
rect 2719 3105 2723 3106
rect 2735 3110 2739 3111
rect 2735 3105 2739 3106
rect 2871 3110 2875 3111
rect 2871 3105 2875 3106
rect 2879 3110 2883 3111
rect 2879 3105 2883 3106
rect 2568 3088 2570 3105
rect 2720 3088 2722 3105
rect 2872 3088 2874 3105
rect 2566 3087 2572 3088
rect 2566 3083 2567 3087
rect 2571 3083 2572 3087
rect 2566 3082 2572 3083
rect 2718 3087 2724 3088
rect 2718 3083 2719 3087
rect 2723 3083 2724 3087
rect 2718 3082 2724 3083
rect 2870 3087 2876 3088
rect 2870 3083 2871 3087
rect 2875 3083 2876 3087
rect 2870 3082 2876 3083
rect 2976 3080 2978 3166
rect 3008 3157 3010 3173
rect 3064 3172 3066 3190
rect 3096 3184 3098 3202
rect 3206 3200 3212 3201
rect 3206 3196 3207 3200
rect 3211 3196 3212 3200
rect 3206 3195 3212 3196
rect 3366 3200 3372 3201
rect 3366 3196 3367 3200
rect 3371 3196 3372 3200
rect 3462 3199 3463 3203
rect 3467 3199 3468 3203
rect 3462 3198 3468 3199
rect 3366 3195 3372 3196
rect 3094 3183 3100 3184
rect 3094 3179 3095 3183
rect 3099 3179 3100 3183
rect 3208 3179 3210 3195
rect 3368 3179 3370 3195
rect 3430 3183 3436 3184
rect 3430 3179 3431 3183
rect 3435 3179 3436 3183
rect 3464 3179 3466 3198
rect 3094 3178 3100 3179
rect 3135 3178 3139 3179
rect 3135 3173 3139 3174
rect 3207 3178 3211 3179
rect 3207 3173 3211 3174
rect 3263 3178 3267 3179
rect 3263 3173 3267 3174
rect 3367 3178 3371 3179
rect 3430 3178 3436 3179
rect 3463 3178 3467 3179
rect 3367 3173 3371 3174
rect 3062 3171 3068 3172
rect 3062 3167 3063 3171
rect 3067 3167 3068 3171
rect 3062 3166 3068 3167
rect 3078 3171 3084 3172
rect 3078 3167 3079 3171
rect 3083 3167 3084 3171
rect 3078 3166 3084 3167
rect 3006 3156 3012 3157
rect 3006 3152 3007 3156
rect 3011 3152 3012 3156
rect 3006 3151 3012 3152
rect 3080 3148 3082 3166
rect 3136 3157 3138 3173
rect 3264 3157 3266 3173
rect 3350 3171 3356 3172
rect 3350 3167 3351 3171
rect 3355 3167 3356 3171
rect 3350 3166 3356 3167
rect 3134 3156 3140 3157
rect 3134 3152 3135 3156
rect 3139 3152 3140 3156
rect 3134 3151 3140 3152
rect 3262 3156 3268 3157
rect 3262 3152 3263 3156
rect 3267 3152 3268 3156
rect 3262 3151 3268 3152
rect 3078 3147 3084 3148
rect 3078 3143 3079 3147
rect 3083 3143 3084 3147
rect 3078 3142 3084 3143
rect 3206 3147 3212 3148
rect 3206 3143 3207 3147
rect 3211 3143 3212 3147
rect 3206 3142 3212 3143
rect 3006 3137 3012 3138
rect 3006 3133 3007 3137
rect 3011 3133 3012 3137
rect 3006 3132 3012 3133
rect 3134 3137 3140 3138
rect 3134 3133 3135 3137
rect 3139 3133 3140 3137
rect 3134 3132 3140 3133
rect 3008 3111 3010 3132
rect 3136 3111 3138 3132
rect 3007 3110 3011 3111
rect 3007 3105 3011 3106
rect 3031 3110 3035 3111
rect 3031 3105 3035 3106
rect 3135 3110 3139 3111
rect 3135 3105 3139 3106
rect 3199 3110 3203 3111
rect 3199 3105 3203 3106
rect 3032 3088 3034 3105
rect 3200 3088 3202 3105
rect 3030 3087 3036 3088
rect 3030 3083 3031 3087
rect 3035 3083 3036 3087
rect 3030 3082 3036 3083
rect 3198 3087 3204 3088
rect 3198 3083 3199 3087
rect 3203 3083 3204 3087
rect 3198 3082 3204 3083
rect 2974 3079 2980 3080
rect 2638 3075 2644 3076
rect 2638 3071 2639 3075
rect 2643 3071 2644 3075
rect 2638 3070 2644 3071
rect 2790 3075 2796 3076
rect 2790 3071 2791 3075
rect 2795 3071 2796 3075
rect 2790 3070 2796 3071
rect 2942 3075 2948 3076
rect 2942 3071 2943 3075
rect 2947 3071 2948 3075
rect 2974 3075 2975 3079
rect 2979 3075 2980 3079
rect 2974 3074 2980 3075
rect 2942 3070 2948 3071
rect 2566 3068 2572 3069
rect 2566 3064 2567 3068
rect 2571 3064 2572 3068
rect 2566 3063 2572 3064
rect 2478 3051 2484 3052
rect 2478 3047 2479 3051
rect 2483 3047 2484 3051
rect 2478 3046 2484 3047
rect 2568 3039 2570 3063
rect 2640 3052 2642 3070
rect 2718 3068 2724 3069
rect 2718 3064 2719 3068
rect 2723 3064 2724 3068
rect 2718 3063 2724 3064
rect 2638 3051 2644 3052
rect 2638 3047 2639 3051
rect 2643 3047 2644 3051
rect 2638 3046 2644 3047
rect 2720 3039 2722 3063
rect 2792 3052 2794 3070
rect 2870 3068 2876 3069
rect 2870 3064 2871 3068
rect 2875 3064 2876 3068
rect 2870 3063 2876 3064
rect 2790 3051 2796 3052
rect 2790 3047 2791 3051
rect 2795 3047 2796 3051
rect 2790 3046 2796 3047
rect 2822 3043 2828 3044
rect 2822 3039 2823 3043
rect 2827 3039 2828 3043
rect 2872 3039 2874 3063
rect 2944 3052 2946 3070
rect 3030 3068 3036 3069
rect 3030 3064 3031 3068
rect 3035 3064 3036 3068
rect 3030 3063 3036 3064
rect 3198 3068 3204 3069
rect 3198 3064 3199 3068
rect 3203 3064 3204 3068
rect 3198 3063 3204 3064
rect 2942 3051 2948 3052
rect 2942 3047 2943 3051
rect 2947 3047 2948 3051
rect 2942 3046 2948 3047
rect 3032 3039 3034 3063
rect 3200 3039 3202 3063
rect 3208 3052 3210 3142
rect 3262 3137 3268 3138
rect 3262 3133 3263 3137
rect 3267 3133 3268 3137
rect 3262 3132 3268 3133
rect 3264 3111 3266 3132
rect 3263 3110 3267 3111
rect 3263 3105 3267 3106
rect 3352 3080 3354 3166
rect 3368 3157 3370 3173
rect 3366 3156 3372 3157
rect 3366 3152 3367 3156
rect 3371 3152 3372 3156
rect 3366 3151 3372 3152
rect 3432 3148 3434 3178
rect 3463 3173 3467 3174
rect 3464 3154 3466 3173
rect 3462 3153 3468 3154
rect 3462 3149 3463 3153
rect 3467 3149 3468 3153
rect 3462 3148 3468 3149
rect 3430 3147 3436 3148
rect 3430 3143 3431 3147
rect 3435 3143 3436 3147
rect 3430 3142 3436 3143
rect 3366 3137 3372 3138
rect 3366 3133 3367 3137
rect 3371 3133 3372 3137
rect 3366 3132 3372 3133
rect 3462 3136 3468 3137
rect 3462 3132 3463 3136
rect 3467 3132 3468 3136
rect 3368 3111 3370 3132
rect 3462 3131 3468 3132
rect 3464 3111 3466 3131
rect 3367 3110 3371 3111
rect 3367 3105 3371 3106
rect 3463 3110 3467 3111
rect 3463 3105 3467 3106
rect 3368 3088 3370 3105
rect 3464 3089 3466 3105
rect 3462 3088 3468 3089
rect 3366 3087 3372 3088
rect 3366 3083 3367 3087
rect 3371 3083 3372 3087
rect 3462 3084 3463 3088
rect 3467 3084 3468 3088
rect 3462 3083 3468 3084
rect 3366 3082 3372 3083
rect 3350 3079 3356 3080
rect 3270 3075 3276 3076
rect 3270 3071 3271 3075
rect 3275 3071 3276 3075
rect 3350 3075 3351 3079
rect 3355 3075 3356 3079
rect 3350 3074 3356 3075
rect 3270 3070 3276 3071
rect 3462 3071 3468 3072
rect 3272 3052 3274 3070
rect 3366 3068 3372 3069
rect 3366 3064 3367 3068
rect 3371 3064 3372 3068
rect 3462 3067 3463 3071
rect 3467 3067 3468 3071
rect 3462 3066 3468 3067
rect 3366 3063 3372 3064
rect 3206 3051 3212 3052
rect 3206 3047 3207 3051
rect 3211 3047 3212 3051
rect 3206 3046 3212 3047
rect 3270 3051 3276 3052
rect 3270 3047 3271 3051
rect 3275 3047 3276 3051
rect 3270 3046 3276 3047
rect 3368 3039 3370 3063
rect 3464 3039 3466 3066
rect 2431 3038 2435 3039
rect 2431 3033 2435 3034
rect 2439 3038 2443 3039
rect 2439 3033 2443 3034
rect 2543 3038 2547 3039
rect 2543 3033 2547 3034
rect 2567 3038 2571 3039
rect 2567 3033 2571 3034
rect 2647 3038 2651 3039
rect 2647 3033 2651 3034
rect 2719 3038 2723 3039
rect 2719 3033 2723 3034
rect 2759 3038 2763 3039
rect 2822 3038 2828 3039
rect 2871 3038 2875 3039
rect 2759 3033 2763 3034
rect 2374 3031 2380 3032
rect 2374 3027 2375 3031
rect 2379 3027 2380 3031
rect 2374 3026 2380 3027
rect 2440 3017 2442 3033
rect 2510 3031 2516 3032
rect 2510 3027 2511 3031
rect 2515 3027 2516 3031
rect 2510 3026 2516 3027
rect 2230 3016 2236 3017
rect 2230 3012 2231 3016
rect 2235 3012 2236 3016
rect 2230 3011 2236 3012
rect 2334 3016 2340 3017
rect 2334 3012 2335 3016
rect 2339 3012 2340 3016
rect 2334 3011 2340 3012
rect 2438 3016 2444 3017
rect 2438 3012 2439 3016
rect 2443 3012 2444 3016
rect 2438 3011 2444 3012
rect 2512 3008 2514 3026
rect 2544 3017 2546 3033
rect 2614 3031 2620 3032
rect 2614 3027 2615 3031
rect 2619 3027 2620 3031
rect 2614 3026 2620 3027
rect 2542 3016 2548 3017
rect 2542 3012 2543 3016
rect 2547 3012 2548 3016
rect 2542 3011 2548 3012
rect 2616 3008 2618 3026
rect 2648 3017 2650 3033
rect 2750 3031 2756 3032
rect 2750 3027 2751 3031
rect 2755 3027 2756 3031
rect 2750 3026 2756 3027
rect 2662 3023 2668 3024
rect 2662 3019 2663 3023
rect 2667 3019 2668 3023
rect 2662 3018 2668 3019
rect 2646 3016 2652 3017
rect 2646 3012 2647 3016
rect 2651 3012 2652 3016
rect 2646 3011 2652 3012
rect 2198 3007 2204 3008
rect 2198 3003 2199 3007
rect 2203 3003 2204 3007
rect 2198 3002 2204 3003
rect 2398 3007 2404 3008
rect 2398 3003 2399 3007
rect 2403 3003 2404 3007
rect 2398 3002 2404 3003
rect 2510 3007 2516 3008
rect 2510 3003 2511 3007
rect 2515 3003 2516 3007
rect 2510 3002 2516 3003
rect 2614 3007 2620 3008
rect 2614 3003 2615 3007
rect 2619 3003 2620 3007
rect 2614 3002 2620 3003
rect 2230 2997 2236 2998
rect 2230 2993 2231 2997
rect 2235 2993 2236 2997
rect 2230 2992 2236 2993
rect 2334 2997 2340 2998
rect 2334 2993 2335 2997
rect 2339 2993 2340 2997
rect 2334 2992 2340 2993
rect 2232 2975 2234 2992
rect 2336 2975 2338 2992
rect 2143 2974 2147 2975
rect 2143 2969 2147 2970
rect 2231 2974 2235 2975
rect 2231 2969 2235 2970
rect 2319 2974 2323 2975
rect 2319 2969 2323 2970
rect 2335 2974 2339 2975
rect 2335 2969 2339 2970
rect 2144 2952 2146 2969
rect 2232 2952 2234 2969
rect 2320 2952 2322 2969
rect 1806 2948 1807 2952
rect 1811 2948 1812 2952
rect 1806 2947 1812 2948
rect 2054 2951 2060 2952
rect 2054 2947 2055 2951
rect 2059 2947 2060 2951
rect 2054 2946 2060 2947
rect 2134 2951 2140 2952
rect 2134 2947 2135 2951
rect 2139 2947 2140 2951
rect 2134 2946 2140 2947
rect 2142 2951 2148 2952
rect 2142 2947 2143 2951
rect 2147 2947 2148 2951
rect 2142 2946 2148 2947
rect 2230 2951 2236 2952
rect 2230 2947 2231 2951
rect 2235 2947 2236 2951
rect 2230 2946 2236 2947
rect 2318 2951 2324 2952
rect 2318 2947 2319 2951
rect 2323 2947 2324 2951
rect 2318 2946 2324 2947
rect 2134 2943 2140 2944
rect 2134 2939 2135 2943
rect 2139 2939 2140 2943
rect 2134 2938 2140 2939
rect 2302 2939 2308 2940
rect 1806 2935 1812 2936
rect 1806 2931 1807 2935
rect 1811 2931 1812 2935
rect 1767 2930 1771 2931
rect 1806 2930 1812 2931
rect 2054 2932 2060 2933
rect 1767 2925 1771 2926
rect 1768 2909 1770 2925
rect 1766 2908 1772 2909
rect 1766 2904 1767 2908
rect 1771 2904 1772 2908
rect 1766 2903 1772 2904
rect 1808 2903 1810 2930
rect 2054 2928 2055 2932
rect 2059 2928 2060 2932
rect 2054 2927 2060 2928
rect 2056 2903 2058 2927
rect 2136 2916 2138 2938
rect 2302 2935 2303 2939
rect 2307 2935 2308 2939
rect 2302 2934 2308 2935
rect 2390 2939 2396 2940
rect 2390 2935 2391 2939
rect 2395 2935 2396 2939
rect 2390 2934 2396 2935
rect 2142 2932 2148 2933
rect 2142 2928 2143 2932
rect 2147 2928 2148 2932
rect 2142 2927 2148 2928
rect 2230 2932 2236 2933
rect 2230 2928 2231 2932
rect 2235 2928 2236 2932
rect 2230 2927 2236 2928
rect 2134 2915 2140 2916
rect 2134 2911 2135 2915
rect 2139 2911 2140 2915
rect 2134 2910 2140 2911
rect 2144 2903 2146 2927
rect 2232 2903 2234 2927
rect 2254 2915 2260 2916
rect 2254 2911 2255 2915
rect 2259 2911 2260 2915
rect 2254 2910 2260 2911
rect 1807 2902 1811 2903
rect 750 2899 756 2900
rect 206 2895 212 2896
rect 206 2891 207 2895
rect 211 2891 212 2895
rect 206 2890 212 2891
rect 334 2895 340 2896
rect 334 2891 335 2895
rect 339 2891 340 2895
rect 334 2890 340 2891
rect 502 2895 508 2896
rect 502 2891 503 2895
rect 507 2891 508 2895
rect 502 2890 508 2891
rect 678 2895 684 2896
rect 678 2891 679 2895
rect 683 2891 684 2895
rect 750 2895 751 2899
rect 755 2895 756 2899
rect 1662 2899 1668 2900
rect 750 2894 756 2895
rect 1022 2895 1028 2896
rect 678 2890 684 2891
rect 208 2872 210 2890
rect 262 2888 268 2889
rect 262 2884 263 2888
rect 267 2884 268 2888
rect 262 2883 268 2884
rect 198 2871 204 2872
rect 198 2867 199 2871
rect 203 2867 204 2871
rect 198 2866 204 2867
rect 206 2871 212 2872
rect 206 2867 207 2871
rect 211 2867 212 2871
rect 206 2866 212 2867
rect 264 2863 266 2883
rect 336 2872 338 2890
rect 430 2888 436 2889
rect 430 2884 431 2888
rect 435 2884 436 2888
rect 430 2883 436 2884
rect 334 2871 340 2872
rect 334 2867 335 2871
rect 339 2867 340 2871
rect 334 2866 340 2867
rect 432 2863 434 2883
rect 504 2872 506 2890
rect 606 2888 612 2889
rect 606 2884 607 2888
rect 611 2884 612 2888
rect 606 2883 612 2884
rect 502 2871 508 2872
rect 502 2867 503 2871
rect 507 2867 508 2871
rect 502 2866 508 2867
rect 608 2863 610 2883
rect 680 2872 682 2890
rect 678 2871 684 2872
rect 678 2867 679 2871
rect 683 2867 684 2871
rect 678 2866 684 2867
rect 752 2864 754 2894
rect 1022 2891 1023 2895
rect 1027 2891 1028 2895
rect 1022 2890 1028 2891
rect 1182 2895 1188 2896
rect 1182 2891 1183 2895
rect 1187 2891 1188 2895
rect 1182 2890 1188 2891
rect 1342 2895 1348 2896
rect 1342 2891 1343 2895
rect 1347 2891 1348 2895
rect 1342 2890 1348 2891
rect 1502 2895 1508 2896
rect 1502 2891 1503 2895
rect 1507 2891 1508 2895
rect 1662 2895 1663 2899
rect 1667 2895 1668 2899
rect 1807 2897 1811 2898
rect 2055 2902 2059 2903
rect 2055 2897 2059 2898
rect 2071 2902 2075 2903
rect 2071 2897 2075 2898
rect 2143 2902 2147 2903
rect 2143 2897 2147 2898
rect 2175 2902 2179 2903
rect 2175 2897 2179 2898
rect 2231 2902 2235 2903
rect 2231 2897 2235 2898
rect 1662 2894 1668 2895
rect 1502 2890 1508 2891
rect 1766 2891 1772 2892
rect 782 2888 788 2889
rect 782 2884 783 2888
rect 787 2884 788 2888
rect 782 2883 788 2884
rect 950 2888 956 2889
rect 950 2884 951 2888
rect 955 2884 956 2888
rect 950 2883 956 2884
rect 750 2863 756 2864
rect 784 2863 786 2883
rect 952 2863 954 2883
rect 1024 2872 1026 2890
rect 1110 2888 1116 2889
rect 1110 2884 1111 2888
rect 1115 2884 1116 2888
rect 1110 2883 1116 2884
rect 1022 2871 1028 2872
rect 1022 2867 1023 2871
rect 1027 2867 1028 2871
rect 1022 2866 1028 2867
rect 1112 2863 1114 2883
rect 1184 2872 1186 2890
rect 1270 2888 1276 2889
rect 1270 2884 1271 2888
rect 1275 2884 1276 2888
rect 1270 2883 1276 2884
rect 1182 2871 1188 2872
rect 1182 2867 1183 2871
rect 1187 2867 1188 2871
rect 1182 2866 1188 2867
rect 1272 2863 1274 2883
rect 1344 2872 1346 2890
rect 1430 2888 1436 2889
rect 1430 2884 1431 2888
rect 1435 2884 1436 2888
rect 1430 2883 1436 2884
rect 1342 2871 1348 2872
rect 1342 2867 1343 2871
rect 1347 2867 1348 2871
rect 1342 2866 1348 2867
rect 1398 2863 1404 2864
rect 1432 2863 1434 2883
rect 1504 2872 1506 2890
rect 1590 2888 1596 2889
rect 1590 2884 1591 2888
rect 1595 2884 1596 2888
rect 1766 2887 1767 2891
rect 1771 2887 1772 2891
rect 1766 2886 1772 2887
rect 1590 2883 1596 2884
rect 1502 2871 1508 2872
rect 1502 2867 1503 2871
rect 1507 2867 1508 2871
rect 1502 2866 1508 2867
rect 1592 2863 1594 2883
rect 1768 2863 1770 2886
rect 1808 2878 1810 2897
rect 2054 2891 2060 2892
rect 2054 2887 2055 2891
rect 2059 2887 2060 2891
rect 2054 2886 2060 2887
rect 1806 2877 1812 2878
rect 1806 2873 1807 2877
rect 1811 2873 1812 2877
rect 1806 2872 1812 2873
rect 111 2862 115 2863
rect 111 2857 115 2858
rect 135 2862 139 2863
rect 135 2857 139 2858
rect 255 2862 259 2863
rect 255 2857 259 2858
rect 263 2862 267 2863
rect 263 2857 267 2858
rect 407 2862 411 2863
rect 407 2857 411 2858
rect 431 2862 435 2863
rect 431 2857 435 2858
rect 567 2862 571 2863
rect 567 2857 571 2858
rect 607 2862 611 2863
rect 607 2857 611 2858
rect 727 2862 731 2863
rect 750 2859 751 2863
rect 755 2859 756 2863
rect 750 2858 756 2859
rect 783 2862 787 2863
rect 727 2857 731 2858
rect 783 2857 787 2858
rect 879 2862 883 2863
rect 879 2857 883 2858
rect 951 2862 955 2863
rect 951 2857 955 2858
rect 1023 2862 1027 2863
rect 1023 2857 1027 2858
rect 1111 2862 1115 2863
rect 1111 2857 1115 2858
rect 1167 2862 1171 2863
rect 1167 2857 1171 2858
rect 1271 2862 1275 2863
rect 1271 2857 1275 2858
rect 1311 2862 1315 2863
rect 1398 2859 1399 2863
rect 1403 2859 1404 2863
rect 1398 2858 1404 2859
rect 1431 2862 1435 2863
rect 1311 2857 1315 2858
rect 112 2838 114 2857
rect 136 2841 138 2857
rect 206 2855 212 2856
rect 206 2851 207 2855
rect 211 2851 212 2855
rect 206 2850 212 2851
rect 134 2840 140 2841
rect 110 2837 116 2838
rect 110 2833 111 2837
rect 115 2833 116 2837
rect 134 2836 135 2840
rect 139 2836 140 2840
rect 134 2835 140 2836
rect 110 2832 116 2833
rect 208 2832 210 2850
rect 256 2841 258 2857
rect 326 2855 332 2856
rect 326 2851 327 2855
rect 331 2851 332 2855
rect 326 2850 332 2851
rect 254 2840 260 2841
rect 254 2836 255 2840
rect 259 2836 260 2840
rect 254 2835 260 2836
rect 328 2832 330 2850
rect 408 2841 410 2857
rect 478 2855 484 2856
rect 478 2851 479 2855
rect 483 2851 484 2855
rect 478 2850 484 2851
rect 406 2840 412 2841
rect 406 2836 407 2840
rect 411 2836 412 2840
rect 406 2835 412 2836
rect 480 2832 482 2850
rect 568 2841 570 2857
rect 638 2855 644 2856
rect 638 2851 639 2855
rect 643 2851 644 2855
rect 638 2850 644 2851
rect 566 2840 572 2841
rect 566 2836 567 2840
rect 571 2836 572 2840
rect 566 2835 572 2836
rect 640 2832 642 2850
rect 728 2841 730 2857
rect 880 2841 882 2857
rect 998 2855 1004 2856
rect 998 2851 999 2855
rect 1003 2851 1004 2855
rect 998 2850 1004 2851
rect 726 2840 732 2841
rect 726 2836 727 2840
rect 731 2836 732 2840
rect 726 2835 732 2836
rect 878 2840 884 2841
rect 878 2836 879 2840
rect 883 2836 884 2840
rect 878 2835 884 2836
rect 1000 2832 1002 2850
rect 1024 2841 1026 2857
rect 1094 2855 1100 2856
rect 1094 2851 1095 2855
rect 1099 2851 1100 2855
rect 1094 2850 1100 2851
rect 1022 2840 1028 2841
rect 1022 2836 1023 2840
rect 1027 2836 1028 2840
rect 1022 2835 1028 2836
rect 1096 2832 1098 2850
rect 1168 2841 1170 2857
rect 1238 2855 1244 2856
rect 1238 2851 1239 2855
rect 1243 2851 1244 2855
rect 1238 2850 1244 2851
rect 1166 2840 1172 2841
rect 1166 2836 1167 2840
rect 1171 2836 1172 2840
rect 1166 2835 1172 2836
rect 1240 2832 1242 2850
rect 1278 2847 1284 2848
rect 1278 2843 1279 2847
rect 1283 2843 1284 2847
rect 1278 2842 1284 2843
rect 206 2831 212 2832
rect 206 2827 207 2831
rect 211 2827 212 2831
rect 206 2826 212 2827
rect 326 2831 332 2832
rect 326 2827 327 2831
rect 331 2827 332 2831
rect 326 2826 332 2827
rect 478 2831 484 2832
rect 478 2827 479 2831
rect 483 2827 484 2831
rect 478 2826 484 2827
rect 638 2831 644 2832
rect 638 2827 639 2831
rect 643 2827 644 2831
rect 638 2826 644 2827
rect 646 2831 652 2832
rect 646 2827 647 2831
rect 651 2827 652 2831
rect 646 2826 652 2827
rect 998 2831 1004 2832
rect 998 2827 999 2831
rect 1003 2827 1004 2831
rect 998 2826 1004 2827
rect 1094 2831 1100 2832
rect 1094 2827 1095 2831
rect 1099 2827 1100 2831
rect 1094 2826 1100 2827
rect 1238 2831 1244 2832
rect 1238 2827 1239 2831
rect 1243 2827 1244 2831
rect 1238 2826 1244 2827
rect 134 2821 140 2822
rect 110 2820 116 2821
rect 110 2816 111 2820
rect 115 2816 116 2820
rect 134 2817 135 2821
rect 139 2817 140 2821
rect 134 2816 140 2817
rect 254 2821 260 2822
rect 254 2817 255 2821
rect 259 2817 260 2821
rect 254 2816 260 2817
rect 406 2821 412 2822
rect 406 2817 407 2821
rect 411 2817 412 2821
rect 406 2816 412 2817
rect 566 2821 572 2822
rect 566 2817 567 2821
rect 571 2817 572 2821
rect 566 2816 572 2817
rect 110 2815 116 2816
rect 112 2791 114 2815
rect 136 2791 138 2816
rect 256 2791 258 2816
rect 408 2791 410 2816
rect 568 2791 570 2816
rect 111 2790 115 2791
rect 111 2785 115 2786
rect 135 2790 139 2791
rect 135 2785 139 2786
rect 255 2790 259 2791
rect 255 2785 259 2786
rect 287 2790 291 2791
rect 287 2785 291 2786
rect 391 2790 395 2791
rect 391 2785 395 2786
rect 407 2790 411 2791
rect 407 2785 411 2786
rect 503 2790 507 2791
rect 503 2785 507 2786
rect 567 2790 571 2791
rect 567 2785 571 2786
rect 623 2790 627 2791
rect 623 2785 627 2786
rect 112 2769 114 2785
rect 110 2768 116 2769
rect 288 2768 290 2785
rect 392 2768 394 2785
rect 504 2768 506 2785
rect 624 2768 626 2785
rect 110 2764 111 2768
rect 115 2764 116 2768
rect 110 2763 116 2764
rect 286 2767 292 2768
rect 286 2763 287 2767
rect 291 2763 292 2767
rect 286 2762 292 2763
rect 390 2767 396 2768
rect 390 2763 391 2767
rect 395 2763 396 2767
rect 390 2762 396 2763
rect 502 2767 508 2768
rect 502 2763 503 2767
rect 507 2763 508 2767
rect 502 2762 508 2763
rect 622 2767 628 2768
rect 622 2763 623 2767
rect 627 2763 628 2767
rect 622 2762 628 2763
rect 358 2755 364 2756
rect 110 2751 116 2752
rect 110 2747 111 2751
rect 115 2747 116 2751
rect 358 2751 359 2755
rect 363 2751 364 2755
rect 358 2750 364 2751
rect 462 2755 468 2756
rect 462 2751 463 2755
rect 467 2751 468 2755
rect 462 2750 468 2751
rect 574 2755 580 2756
rect 574 2751 575 2755
rect 579 2751 580 2755
rect 574 2750 580 2751
rect 110 2746 116 2747
rect 286 2748 292 2749
rect 112 2723 114 2746
rect 286 2744 287 2748
rect 291 2744 292 2748
rect 286 2743 292 2744
rect 288 2723 290 2743
rect 360 2732 362 2750
rect 390 2748 396 2749
rect 390 2744 391 2748
rect 395 2744 396 2748
rect 390 2743 396 2744
rect 358 2731 364 2732
rect 358 2727 359 2731
rect 363 2727 364 2731
rect 358 2726 364 2727
rect 392 2723 394 2743
rect 464 2732 466 2750
rect 502 2748 508 2749
rect 502 2744 503 2748
rect 507 2744 508 2748
rect 502 2743 508 2744
rect 462 2731 468 2732
rect 462 2727 463 2731
rect 467 2727 468 2731
rect 462 2726 468 2727
rect 504 2723 506 2743
rect 576 2732 578 2750
rect 622 2748 628 2749
rect 622 2744 623 2748
rect 627 2744 628 2748
rect 622 2743 628 2744
rect 574 2731 580 2732
rect 574 2727 575 2731
rect 579 2727 580 2731
rect 574 2726 580 2727
rect 624 2723 626 2743
rect 648 2740 650 2826
rect 726 2821 732 2822
rect 726 2817 727 2821
rect 731 2817 732 2821
rect 726 2816 732 2817
rect 878 2821 884 2822
rect 878 2817 879 2821
rect 883 2817 884 2821
rect 878 2816 884 2817
rect 1022 2821 1028 2822
rect 1022 2817 1023 2821
rect 1027 2817 1028 2821
rect 1022 2816 1028 2817
rect 1166 2821 1172 2822
rect 1166 2817 1167 2821
rect 1171 2817 1172 2821
rect 1166 2816 1172 2817
rect 728 2791 730 2816
rect 880 2791 882 2816
rect 1024 2791 1026 2816
rect 1168 2791 1170 2816
rect 727 2790 731 2791
rect 727 2785 731 2786
rect 743 2790 747 2791
rect 743 2785 747 2786
rect 855 2790 859 2791
rect 855 2785 859 2786
rect 879 2790 883 2791
rect 879 2785 883 2786
rect 967 2790 971 2791
rect 967 2785 971 2786
rect 1023 2790 1027 2791
rect 1023 2785 1027 2786
rect 1079 2790 1083 2791
rect 1079 2785 1083 2786
rect 1167 2790 1171 2791
rect 1167 2785 1171 2786
rect 1199 2790 1203 2791
rect 1199 2785 1203 2786
rect 744 2768 746 2785
rect 856 2768 858 2785
rect 968 2768 970 2785
rect 1080 2768 1082 2785
rect 1200 2768 1202 2785
rect 742 2767 748 2768
rect 742 2763 743 2767
rect 747 2763 748 2767
rect 742 2762 748 2763
rect 854 2767 860 2768
rect 854 2763 855 2767
rect 859 2763 860 2767
rect 854 2762 860 2763
rect 966 2767 972 2768
rect 966 2763 967 2767
rect 971 2763 972 2767
rect 966 2762 972 2763
rect 1078 2767 1084 2768
rect 1078 2763 1079 2767
rect 1083 2763 1084 2767
rect 1078 2762 1084 2763
rect 1198 2767 1204 2768
rect 1198 2763 1199 2767
rect 1203 2763 1204 2767
rect 1198 2762 1204 2763
rect 1280 2760 1282 2842
rect 1312 2841 1314 2857
rect 1382 2855 1388 2856
rect 1382 2851 1383 2855
rect 1387 2851 1388 2855
rect 1382 2850 1388 2851
rect 1310 2840 1316 2841
rect 1310 2836 1311 2840
rect 1315 2836 1316 2840
rect 1310 2835 1316 2836
rect 1384 2832 1386 2850
rect 1400 2832 1402 2858
rect 1431 2857 1435 2858
rect 1463 2862 1467 2863
rect 1463 2857 1467 2858
rect 1591 2862 1595 2863
rect 1591 2857 1595 2858
rect 1767 2862 1771 2863
rect 1767 2857 1771 2858
rect 1806 2860 1812 2861
rect 1464 2841 1466 2857
rect 1462 2840 1468 2841
rect 1462 2836 1463 2840
rect 1467 2836 1468 2840
rect 1768 2838 1770 2857
rect 1806 2856 1807 2860
rect 1811 2856 1812 2860
rect 1806 2855 1812 2856
rect 1462 2835 1468 2836
rect 1766 2837 1772 2838
rect 1766 2833 1767 2837
rect 1771 2833 1772 2837
rect 1808 2835 1810 2855
rect 1766 2832 1772 2833
rect 1807 2834 1811 2835
rect 1382 2831 1388 2832
rect 1382 2827 1383 2831
rect 1387 2827 1388 2831
rect 1382 2826 1388 2827
rect 1398 2831 1404 2832
rect 1398 2827 1399 2831
rect 1403 2827 1404 2831
rect 1807 2829 1811 2830
rect 1983 2834 1987 2835
rect 1983 2829 1987 2830
rect 1398 2826 1404 2827
rect 1310 2821 1316 2822
rect 1310 2817 1311 2821
rect 1315 2817 1316 2821
rect 1310 2816 1316 2817
rect 1462 2821 1468 2822
rect 1462 2817 1463 2821
rect 1467 2817 1468 2821
rect 1462 2816 1468 2817
rect 1766 2820 1772 2821
rect 1766 2816 1767 2820
rect 1771 2816 1772 2820
rect 1312 2791 1314 2816
rect 1464 2791 1466 2816
rect 1766 2815 1772 2816
rect 1768 2791 1770 2815
rect 1808 2813 1810 2829
rect 1806 2812 1812 2813
rect 1984 2812 1986 2829
rect 1806 2808 1807 2812
rect 1811 2808 1812 2812
rect 1806 2807 1812 2808
rect 1982 2811 1988 2812
rect 1982 2807 1983 2811
rect 1987 2807 1988 2811
rect 1982 2806 1988 2807
rect 2056 2804 2058 2886
rect 2072 2881 2074 2897
rect 2176 2881 2178 2897
rect 2246 2895 2252 2896
rect 2246 2891 2247 2895
rect 2251 2891 2252 2895
rect 2246 2890 2252 2891
rect 2070 2880 2076 2881
rect 2070 2876 2071 2880
rect 2075 2876 2076 2880
rect 2070 2875 2076 2876
rect 2174 2880 2180 2881
rect 2174 2876 2175 2880
rect 2179 2876 2180 2880
rect 2174 2875 2180 2876
rect 2248 2872 2250 2890
rect 2256 2872 2258 2910
rect 2304 2908 2306 2934
rect 2318 2932 2324 2933
rect 2318 2928 2319 2932
rect 2323 2928 2324 2932
rect 2318 2927 2324 2928
rect 2302 2907 2308 2908
rect 2302 2903 2303 2907
rect 2307 2903 2308 2907
rect 2320 2903 2322 2927
rect 2271 2902 2275 2903
rect 2302 2902 2308 2903
rect 2319 2902 2323 2903
rect 2271 2897 2275 2898
rect 2319 2897 2323 2898
rect 2367 2902 2371 2903
rect 2367 2897 2371 2898
rect 2272 2881 2274 2897
rect 2368 2881 2370 2897
rect 2392 2896 2394 2934
rect 2400 2916 2402 3002
rect 2438 2997 2444 2998
rect 2438 2993 2439 2997
rect 2443 2993 2444 2997
rect 2438 2992 2444 2993
rect 2542 2997 2548 2998
rect 2542 2993 2543 2997
rect 2547 2993 2548 2997
rect 2542 2992 2548 2993
rect 2646 2997 2652 2998
rect 2646 2993 2647 2997
rect 2651 2993 2652 2997
rect 2646 2992 2652 2993
rect 2440 2975 2442 2992
rect 2544 2975 2546 2992
rect 2648 2975 2650 2992
rect 2407 2974 2411 2975
rect 2407 2969 2411 2970
rect 2439 2974 2443 2975
rect 2439 2969 2443 2970
rect 2495 2974 2499 2975
rect 2495 2969 2499 2970
rect 2543 2974 2547 2975
rect 2543 2969 2547 2970
rect 2583 2974 2587 2975
rect 2583 2969 2587 2970
rect 2647 2974 2651 2975
rect 2647 2969 2651 2970
rect 2408 2952 2410 2969
rect 2496 2952 2498 2969
rect 2584 2952 2586 2969
rect 2406 2951 2412 2952
rect 2406 2947 2407 2951
rect 2411 2947 2412 2951
rect 2406 2946 2412 2947
rect 2494 2951 2500 2952
rect 2494 2947 2495 2951
rect 2499 2947 2500 2951
rect 2494 2946 2500 2947
rect 2582 2951 2588 2952
rect 2582 2947 2583 2951
rect 2587 2947 2588 2951
rect 2582 2946 2588 2947
rect 2664 2944 2666 3018
rect 2752 3008 2754 3026
rect 2760 3017 2762 3033
rect 2758 3016 2764 3017
rect 2758 3012 2759 3016
rect 2763 3012 2764 3016
rect 2758 3011 2764 3012
rect 2824 3008 2826 3038
rect 2871 3033 2875 3034
rect 3031 3038 3035 3039
rect 3031 3033 3035 3034
rect 3199 3038 3203 3039
rect 3199 3033 3203 3034
rect 3367 3038 3371 3039
rect 3367 3033 3371 3034
rect 3463 3038 3467 3039
rect 3463 3033 3467 3034
rect 3464 3014 3466 3033
rect 3462 3013 3468 3014
rect 3462 3009 3463 3013
rect 3467 3009 3468 3013
rect 3462 3008 3468 3009
rect 2750 3007 2756 3008
rect 2750 3003 2751 3007
rect 2755 3003 2756 3007
rect 2750 3002 2756 3003
rect 2822 3007 2828 3008
rect 2822 3003 2823 3007
rect 2827 3003 2828 3007
rect 2822 3002 2828 3003
rect 2758 2997 2764 2998
rect 2758 2993 2759 2997
rect 2763 2993 2764 2997
rect 2758 2992 2764 2993
rect 3462 2996 3468 2997
rect 3462 2992 3463 2996
rect 3467 2992 3468 2996
rect 2760 2975 2762 2992
rect 3462 2991 3468 2992
rect 3464 2975 3466 2991
rect 2671 2974 2675 2975
rect 2671 2969 2675 2970
rect 2759 2974 2763 2975
rect 2759 2969 2763 2970
rect 2847 2974 2851 2975
rect 2847 2969 2851 2970
rect 3463 2974 3467 2975
rect 3463 2969 3467 2970
rect 2672 2952 2674 2969
rect 2760 2952 2762 2969
rect 2848 2952 2850 2969
rect 3464 2953 3466 2969
rect 3462 2952 3468 2953
rect 2670 2951 2676 2952
rect 2670 2947 2671 2951
rect 2675 2947 2676 2951
rect 2670 2946 2676 2947
rect 2758 2951 2764 2952
rect 2758 2947 2759 2951
rect 2763 2947 2764 2951
rect 2758 2946 2764 2947
rect 2846 2951 2852 2952
rect 2846 2947 2847 2951
rect 2851 2947 2852 2951
rect 3462 2948 3463 2952
rect 3467 2948 3468 2952
rect 3462 2947 3468 2948
rect 2846 2946 2852 2947
rect 2662 2943 2668 2944
rect 2478 2939 2484 2940
rect 2478 2935 2479 2939
rect 2483 2935 2484 2939
rect 2478 2934 2484 2935
rect 2566 2939 2572 2940
rect 2566 2935 2567 2939
rect 2571 2935 2572 2939
rect 2566 2934 2572 2935
rect 2654 2939 2660 2940
rect 2654 2935 2655 2939
rect 2659 2935 2660 2939
rect 2662 2939 2663 2943
rect 2667 2939 2668 2943
rect 2662 2938 2668 2939
rect 2750 2943 2756 2944
rect 2750 2939 2751 2943
rect 2755 2939 2756 2943
rect 2750 2938 2756 2939
rect 2838 2943 2844 2944
rect 2838 2939 2839 2943
rect 2843 2939 2844 2943
rect 2838 2938 2844 2939
rect 2654 2934 2660 2935
rect 2406 2932 2412 2933
rect 2406 2928 2407 2932
rect 2411 2928 2412 2932
rect 2406 2927 2412 2928
rect 2398 2915 2404 2916
rect 2398 2911 2399 2915
rect 2403 2911 2404 2915
rect 2398 2910 2404 2911
rect 2408 2903 2410 2927
rect 2480 2916 2482 2934
rect 2494 2932 2500 2933
rect 2494 2928 2495 2932
rect 2499 2928 2500 2932
rect 2494 2927 2500 2928
rect 2478 2915 2484 2916
rect 2478 2911 2479 2915
rect 2483 2911 2484 2915
rect 2478 2910 2484 2911
rect 2496 2903 2498 2927
rect 2568 2916 2570 2934
rect 2582 2932 2588 2933
rect 2582 2928 2583 2932
rect 2587 2928 2588 2932
rect 2582 2927 2588 2928
rect 2566 2915 2572 2916
rect 2566 2911 2567 2915
rect 2571 2911 2572 2915
rect 2566 2910 2572 2911
rect 2584 2903 2586 2927
rect 2656 2916 2658 2934
rect 2670 2932 2676 2933
rect 2670 2928 2671 2932
rect 2675 2928 2676 2932
rect 2670 2927 2676 2928
rect 2654 2915 2660 2916
rect 2654 2911 2655 2915
rect 2659 2911 2660 2915
rect 2654 2910 2660 2911
rect 2672 2903 2674 2927
rect 2752 2924 2754 2938
rect 2758 2932 2764 2933
rect 2758 2928 2759 2932
rect 2763 2928 2764 2932
rect 2758 2927 2764 2928
rect 2750 2923 2756 2924
rect 2750 2919 2751 2923
rect 2755 2919 2756 2923
rect 2750 2918 2756 2919
rect 2760 2903 2762 2927
rect 2840 2916 2842 2938
rect 3462 2935 3468 2936
rect 2846 2932 2852 2933
rect 2846 2928 2847 2932
rect 2851 2928 2852 2932
rect 3462 2931 3463 2935
rect 3467 2931 3468 2935
rect 3462 2930 3468 2931
rect 2846 2927 2852 2928
rect 2838 2915 2844 2916
rect 2838 2911 2839 2915
rect 2843 2911 2844 2915
rect 2838 2910 2844 2911
rect 2848 2903 2850 2927
rect 2854 2915 2860 2916
rect 2854 2911 2855 2915
rect 2859 2911 2860 2915
rect 2854 2910 2860 2911
rect 2407 2902 2411 2903
rect 2407 2897 2411 2898
rect 2471 2902 2475 2903
rect 2471 2897 2475 2898
rect 2495 2902 2499 2903
rect 2495 2897 2499 2898
rect 2575 2902 2579 2903
rect 2575 2897 2579 2898
rect 2583 2902 2587 2903
rect 2583 2897 2587 2898
rect 2671 2902 2675 2903
rect 2671 2897 2675 2898
rect 2679 2902 2683 2903
rect 2679 2897 2683 2898
rect 2759 2902 2763 2903
rect 2759 2897 2763 2898
rect 2783 2902 2787 2903
rect 2783 2897 2787 2898
rect 2847 2902 2851 2903
rect 2847 2897 2851 2898
rect 2390 2895 2396 2896
rect 2390 2891 2391 2895
rect 2395 2891 2396 2895
rect 2390 2890 2396 2891
rect 2472 2881 2474 2897
rect 2558 2895 2564 2896
rect 2558 2891 2559 2895
rect 2563 2891 2564 2895
rect 2558 2890 2564 2891
rect 2270 2880 2276 2881
rect 2270 2876 2271 2880
rect 2275 2876 2276 2880
rect 2270 2875 2276 2876
rect 2366 2880 2372 2881
rect 2366 2876 2367 2880
rect 2371 2876 2372 2880
rect 2366 2875 2372 2876
rect 2470 2880 2476 2881
rect 2470 2876 2471 2880
rect 2475 2876 2476 2880
rect 2470 2875 2476 2876
rect 2246 2871 2252 2872
rect 2246 2867 2247 2871
rect 2251 2867 2252 2871
rect 2246 2866 2252 2867
rect 2254 2871 2260 2872
rect 2254 2867 2255 2871
rect 2259 2867 2260 2871
rect 2254 2866 2260 2867
rect 2430 2871 2436 2872
rect 2430 2867 2431 2871
rect 2435 2867 2436 2871
rect 2430 2866 2436 2867
rect 2070 2861 2076 2862
rect 2070 2857 2071 2861
rect 2075 2857 2076 2861
rect 2070 2856 2076 2857
rect 2174 2861 2180 2862
rect 2174 2857 2175 2861
rect 2179 2857 2180 2861
rect 2174 2856 2180 2857
rect 2270 2861 2276 2862
rect 2270 2857 2271 2861
rect 2275 2857 2276 2861
rect 2270 2856 2276 2857
rect 2366 2861 2372 2862
rect 2366 2857 2367 2861
rect 2371 2857 2372 2861
rect 2366 2856 2372 2857
rect 2072 2835 2074 2856
rect 2176 2835 2178 2856
rect 2272 2835 2274 2856
rect 2368 2835 2370 2856
rect 2071 2834 2075 2835
rect 2071 2829 2075 2830
rect 2111 2834 2115 2835
rect 2111 2829 2115 2830
rect 2175 2834 2179 2835
rect 2175 2829 2179 2830
rect 2239 2834 2243 2835
rect 2239 2829 2243 2830
rect 2271 2834 2275 2835
rect 2271 2829 2275 2830
rect 2367 2834 2371 2835
rect 2367 2829 2371 2830
rect 2112 2812 2114 2829
rect 2240 2812 2242 2829
rect 2368 2812 2370 2829
rect 2110 2811 2116 2812
rect 2110 2807 2111 2811
rect 2115 2807 2116 2811
rect 2110 2806 2116 2807
rect 2238 2811 2244 2812
rect 2238 2807 2239 2811
rect 2243 2807 2244 2811
rect 2238 2806 2244 2807
rect 2366 2811 2372 2812
rect 2366 2807 2367 2811
rect 2371 2807 2372 2811
rect 2366 2806 2372 2807
rect 2054 2803 2060 2804
rect 2054 2799 2055 2803
rect 2059 2799 2060 2803
rect 2054 2798 2060 2799
rect 2062 2803 2068 2804
rect 2062 2799 2063 2803
rect 2067 2799 2068 2803
rect 2062 2798 2068 2799
rect 2190 2803 2196 2804
rect 2190 2799 2191 2803
rect 2195 2799 2196 2803
rect 2190 2798 2196 2799
rect 1806 2795 1812 2796
rect 1806 2791 1807 2795
rect 1811 2791 1812 2795
rect 1311 2790 1315 2791
rect 1311 2785 1315 2786
rect 1319 2790 1323 2791
rect 1319 2785 1323 2786
rect 1463 2790 1467 2791
rect 1463 2785 1467 2786
rect 1767 2790 1771 2791
rect 1806 2790 1812 2791
rect 1982 2792 1988 2793
rect 1767 2785 1771 2786
rect 1320 2768 1322 2785
rect 1768 2769 1770 2785
rect 1766 2768 1772 2769
rect 1318 2767 1324 2768
rect 1318 2763 1319 2767
rect 1323 2763 1324 2767
rect 1766 2764 1767 2768
rect 1771 2764 1772 2768
rect 1808 2767 1810 2790
rect 1982 2788 1983 2792
rect 1987 2788 1988 2792
rect 1982 2787 1988 2788
rect 1984 2767 1986 2787
rect 2064 2776 2066 2798
rect 2110 2792 2116 2793
rect 2110 2788 2111 2792
rect 2115 2788 2116 2792
rect 2110 2787 2116 2788
rect 2062 2775 2068 2776
rect 2062 2771 2063 2775
rect 2067 2771 2068 2775
rect 2062 2770 2068 2771
rect 2112 2767 2114 2787
rect 2192 2776 2194 2798
rect 2238 2792 2244 2793
rect 2238 2788 2239 2792
rect 2243 2788 2244 2792
rect 2238 2787 2244 2788
rect 2366 2792 2372 2793
rect 2366 2788 2367 2792
rect 2371 2788 2372 2792
rect 2366 2787 2372 2788
rect 2190 2775 2196 2776
rect 2190 2771 2191 2775
rect 2195 2771 2196 2775
rect 2190 2770 2196 2771
rect 2240 2767 2242 2787
rect 2254 2775 2260 2776
rect 2254 2771 2255 2775
rect 2259 2771 2260 2775
rect 2254 2770 2260 2771
rect 1766 2763 1772 2764
rect 1807 2766 1811 2767
rect 1318 2762 1324 2763
rect 1807 2761 1811 2762
rect 1887 2766 1891 2767
rect 1887 2761 1891 2762
rect 1983 2766 1987 2767
rect 1983 2761 1987 2762
rect 2031 2766 2035 2767
rect 2031 2761 2035 2762
rect 2111 2766 2115 2767
rect 2111 2761 2115 2762
rect 2183 2766 2187 2767
rect 2183 2761 2187 2762
rect 2239 2766 2243 2767
rect 2239 2761 2243 2762
rect 730 2759 736 2760
rect 694 2755 700 2756
rect 694 2751 695 2755
rect 699 2751 700 2755
rect 730 2755 731 2759
rect 735 2755 736 2759
rect 1278 2759 1284 2760
rect 730 2754 736 2755
rect 926 2755 932 2756
rect 694 2750 700 2751
rect 646 2739 652 2740
rect 646 2735 647 2739
rect 651 2735 652 2739
rect 646 2734 652 2735
rect 696 2732 698 2750
rect 694 2731 700 2732
rect 694 2727 695 2731
rect 699 2727 700 2731
rect 694 2726 700 2727
rect 732 2724 734 2754
rect 926 2751 927 2755
rect 931 2751 932 2755
rect 926 2750 932 2751
rect 1038 2755 1044 2756
rect 1038 2751 1039 2755
rect 1043 2751 1044 2755
rect 1038 2750 1044 2751
rect 1150 2755 1156 2756
rect 1150 2751 1151 2755
rect 1155 2751 1156 2755
rect 1150 2750 1156 2751
rect 1270 2755 1276 2756
rect 1270 2751 1271 2755
rect 1275 2751 1276 2755
rect 1278 2755 1279 2759
rect 1283 2755 1284 2759
rect 1278 2754 1284 2755
rect 1270 2750 1276 2751
rect 1766 2751 1772 2752
rect 742 2748 748 2749
rect 742 2744 743 2748
rect 747 2744 748 2748
rect 742 2743 748 2744
rect 854 2748 860 2749
rect 854 2744 855 2748
rect 859 2744 860 2748
rect 854 2743 860 2744
rect 730 2723 736 2724
rect 744 2723 746 2743
rect 856 2723 858 2743
rect 928 2732 930 2750
rect 966 2748 972 2749
rect 966 2744 967 2748
rect 971 2744 972 2748
rect 966 2743 972 2744
rect 926 2731 932 2732
rect 926 2727 927 2731
rect 931 2727 932 2731
rect 926 2726 932 2727
rect 968 2723 970 2743
rect 1040 2732 1042 2750
rect 1078 2748 1084 2749
rect 1078 2744 1079 2748
rect 1083 2744 1084 2748
rect 1078 2743 1084 2744
rect 1038 2731 1044 2732
rect 1038 2727 1039 2731
rect 1043 2727 1044 2731
rect 1038 2726 1044 2727
rect 1080 2723 1082 2743
rect 1152 2732 1154 2750
rect 1198 2748 1204 2749
rect 1198 2744 1199 2748
rect 1203 2744 1204 2748
rect 1198 2743 1204 2744
rect 1150 2731 1156 2732
rect 1150 2727 1151 2731
rect 1155 2727 1156 2731
rect 1150 2726 1156 2727
rect 1174 2723 1180 2724
rect 1200 2723 1202 2743
rect 1272 2732 1274 2750
rect 1318 2748 1324 2749
rect 1318 2744 1319 2748
rect 1323 2744 1324 2748
rect 1766 2747 1767 2751
rect 1771 2747 1772 2751
rect 1766 2746 1772 2747
rect 1318 2743 1324 2744
rect 1270 2731 1276 2732
rect 1270 2727 1271 2731
rect 1275 2727 1276 2731
rect 1270 2726 1276 2727
rect 1320 2723 1322 2743
rect 1768 2723 1770 2746
rect 1808 2742 1810 2761
rect 1888 2745 1890 2761
rect 1902 2759 1908 2760
rect 1902 2755 1903 2759
rect 1907 2755 1908 2759
rect 1902 2754 1908 2755
rect 1958 2759 1964 2760
rect 1958 2755 1959 2759
rect 1963 2755 1964 2759
rect 1958 2754 1964 2755
rect 1886 2744 1892 2745
rect 1806 2741 1812 2742
rect 1806 2737 1807 2741
rect 1811 2737 1812 2741
rect 1886 2740 1887 2744
rect 1891 2740 1892 2744
rect 1886 2739 1892 2740
rect 1806 2736 1812 2737
rect 1886 2725 1892 2726
rect 1806 2724 1812 2725
rect 111 2722 115 2723
rect 111 2717 115 2718
rect 287 2722 291 2723
rect 287 2717 291 2718
rect 391 2722 395 2723
rect 391 2717 395 2718
rect 479 2722 483 2723
rect 479 2717 483 2718
rect 503 2722 507 2723
rect 503 2717 507 2718
rect 567 2722 571 2723
rect 567 2717 571 2718
rect 623 2722 627 2723
rect 623 2717 627 2718
rect 655 2722 659 2723
rect 730 2719 731 2723
rect 735 2719 736 2723
rect 730 2718 736 2719
rect 743 2722 747 2723
rect 655 2717 659 2718
rect 743 2717 747 2718
rect 831 2722 835 2723
rect 831 2717 835 2718
rect 855 2722 859 2723
rect 855 2717 859 2718
rect 919 2722 923 2723
rect 919 2717 923 2718
rect 967 2722 971 2723
rect 967 2717 971 2718
rect 1007 2722 1011 2723
rect 1007 2717 1011 2718
rect 1079 2722 1083 2723
rect 1079 2717 1083 2718
rect 1095 2722 1099 2723
rect 1174 2719 1175 2723
rect 1179 2719 1180 2723
rect 1174 2718 1180 2719
rect 1183 2722 1187 2723
rect 1095 2717 1099 2718
rect 112 2698 114 2717
rect 480 2701 482 2717
rect 550 2715 556 2716
rect 550 2711 551 2715
rect 555 2711 556 2715
rect 550 2710 556 2711
rect 478 2700 484 2701
rect 110 2697 116 2698
rect 110 2693 111 2697
rect 115 2693 116 2697
rect 478 2696 479 2700
rect 483 2696 484 2700
rect 478 2695 484 2696
rect 110 2692 116 2693
rect 552 2692 554 2710
rect 568 2701 570 2717
rect 638 2715 644 2716
rect 638 2711 639 2715
rect 643 2711 644 2715
rect 638 2710 644 2711
rect 566 2700 572 2701
rect 566 2696 567 2700
rect 571 2696 572 2700
rect 566 2695 572 2696
rect 640 2692 642 2710
rect 656 2701 658 2717
rect 726 2715 732 2716
rect 726 2711 727 2715
rect 731 2711 732 2715
rect 726 2710 732 2711
rect 654 2700 660 2701
rect 654 2696 655 2700
rect 659 2696 660 2700
rect 654 2695 660 2696
rect 728 2692 730 2710
rect 744 2701 746 2717
rect 814 2715 820 2716
rect 814 2711 815 2715
rect 819 2711 820 2715
rect 814 2710 820 2711
rect 742 2700 748 2701
rect 742 2696 743 2700
rect 747 2696 748 2700
rect 742 2695 748 2696
rect 816 2692 818 2710
rect 832 2701 834 2717
rect 920 2701 922 2717
rect 990 2715 996 2716
rect 990 2711 991 2715
rect 995 2711 996 2715
rect 990 2710 996 2711
rect 830 2700 836 2701
rect 830 2696 831 2700
rect 835 2696 836 2700
rect 830 2695 836 2696
rect 918 2700 924 2701
rect 918 2696 919 2700
rect 923 2696 924 2700
rect 918 2695 924 2696
rect 992 2692 994 2710
rect 1008 2701 1010 2717
rect 1078 2707 1084 2708
rect 1078 2703 1079 2707
rect 1083 2703 1084 2707
rect 1078 2702 1084 2703
rect 1006 2700 1012 2701
rect 1006 2696 1007 2700
rect 1011 2696 1012 2700
rect 1006 2695 1012 2696
rect 550 2691 556 2692
rect 550 2687 551 2691
rect 555 2687 556 2691
rect 550 2686 556 2687
rect 638 2691 644 2692
rect 638 2687 639 2691
rect 643 2687 644 2691
rect 638 2686 644 2687
rect 726 2691 732 2692
rect 726 2687 727 2691
rect 731 2687 732 2691
rect 726 2686 732 2687
rect 814 2691 820 2692
rect 814 2687 815 2691
rect 819 2687 820 2691
rect 814 2686 820 2687
rect 902 2691 908 2692
rect 902 2687 903 2691
rect 907 2687 908 2691
rect 902 2686 908 2687
rect 990 2691 996 2692
rect 990 2687 991 2691
rect 995 2687 996 2691
rect 990 2686 996 2687
rect 478 2681 484 2682
rect 110 2680 116 2681
rect 110 2676 111 2680
rect 115 2676 116 2680
rect 478 2677 479 2681
rect 483 2677 484 2681
rect 478 2676 484 2677
rect 566 2681 572 2682
rect 566 2677 567 2681
rect 571 2677 572 2681
rect 566 2676 572 2677
rect 654 2681 660 2682
rect 654 2677 655 2681
rect 659 2677 660 2681
rect 654 2676 660 2677
rect 742 2681 748 2682
rect 742 2677 743 2681
rect 747 2677 748 2681
rect 742 2676 748 2677
rect 830 2681 836 2682
rect 830 2677 831 2681
rect 835 2677 836 2681
rect 830 2676 836 2677
rect 110 2675 116 2676
rect 112 2651 114 2675
rect 480 2651 482 2676
rect 568 2651 570 2676
rect 656 2651 658 2676
rect 744 2651 746 2676
rect 832 2651 834 2676
rect 111 2650 115 2651
rect 111 2645 115 2646
rect 471 2650 475 2651
rect 471 2645 475 2646
rect 479 2650 483 2651
rect 479 2645 483 2646
rect 559 2650 563 2651
rect 559 2645 563 2646
rect 567 2650 571 2651
rect 567 2645 571 2646
rect 647 2650 651 2651
rect 647 2645 651 2646
rect 655 2650 659 2651
rect 655 2645 659 2646
rect 735 2650 739 2651
rect 735 2645 739 2646
rect 743 2650 747 2651
rect 743 2645 747 2646
rect 823 2650 827 2651
rect 823 2645 827 2646
rect 831 2650 835 2651
rect 831 2645 835 2646
rect 112 2629 114 2645
rect 110 2628 116 2629
rect 472 2628 474 2645
rect 560 2628 562 2645
rect 648 2628 650 2645
rect 736 2628 738 2645
rect 824 2628 826 2645
rect 110 2624 111 2628
rect 115 2624 116 2628
rect 110 2623 116 2624
rect 470 2627 476 2628
rect 470 2623 471 2627
rect 475 2623 476 2627
rect 470 2622 476 2623
rect 558 2627 564 2628
rect 558 2623 559 2627
rect 563 2623 564 2627
rect 558 2622 564 2623
rect 646 2627 652 2628
rect 646 2623 647 2627
rect 651 2623 652 2627
rect 646 2622 652 2623
rect 734 2627 740 2628
rect 734 2623 735 2627
rect 739 2623 740 2627
rect 734 2622 740 2623
rect 822 2627 828 2628
rect 822 2623 823 2627
rect 827 2623 828 2627
rect 822 2622 828 2623
rect 550 2619 556 2620
rect 542 2615 548 2616
rect 110 2611 116 2612
rect 110 2607 111 2611
rect 115 2607 116 2611
rect 542 2611 543 2615
rect 547 2611 548 2615
rect 550 2615 551 2619
rect 555 2615 556 2619
rect 550 2614 556 2615
rect 638 2619 644 2620
rect 638 2615 639 2619
rect 643 2615 644 2619
rect 638 2614 644 2615
rect 726 2619 732 2620
rect 726 2615 727 2619
rect 731 2615 732 2619
rect 726 2614 732 2615
rect 814 2619 820 2620
rect 814 2615 815 2619
rect 819 2615 820 2619
rect 814 2614 820 2615
rect 542 2610 548 2611
rect 110 2606 116 2607
rect 470 2608 476 2609
rect 112 2575 114 2606
rect 470 2604 471 2608
rect 475 2604 476 2608
rect 470 2603 476 2604
rect 472 2575 474 2603
rect 111 2574 115 2575
rect 111 2569 115 2570
rect 223 2574 227 2575
rect 223 2569 227 2570
rect 311 2574 315 2575
rect 311 2569 315 2570
rect 407 2574 411 2575
rect 407 2569 411 2570
rect 471 2574 475 2575
rect 471 2569 475 2570
rect 503 2574 507 2575
rect 503 2569 507 2570
rect 112 2550 114 2569
rect 224 2553 226 2569
rect 294 2567 300 2568
rect 294 2563 295 2567
rect 299 2563 300 2567
rect 294 2562 300 2563
rect 222 2552 228 2553
rect 110 2549 116 2550
rect 110 2545 111 2549
rect 115 2545 116 2549
rect 222 2548 223 2552
rect 227 2548 228 2552
rect 222 2547 228 2548
rect 110 2544 116 2545
rect 296 2544 298 2562
rect 312 2553 314 2569
rect 408 2553 410 2569
rect 504 2553 506 2569
rect 544 2568 546 2610
rect 552 2592 554 2614
rect 558 2608 564 2609
rect 558 2604 559 2608
rect 563 2604 564 2608
rect 558 2603 564 2604
rect 550 2591 556 2592
rect 550 2587 551 2591
rect 555 2587 556 2591
rect 550 2586 556 2587
rect 560 2575 562 2603
rect 640 2592 642 2614
rect 646 2608 652 2609
rect 646 2604 647 2608
rect 651 2604 652 2608
rect 646 2603 652 2604
rect 638 2591 644 2592
rect 638 2587 639 2591
rect 643 2587 644 2591
rect 638 2586 644 2587
rect 648 2575 650 2603
rect 728 2592 730 2614
rect 734 2608 740 2609
rect 734 2604 735 2608
rect 739 2604 740 2608
rect 734 2603 740 2604
rect 726 2591 732 2592
rect 726 2587 727 2591
rect 731 2587 732 2591
rect 726 2586 732 2587
rect 736 2575 738 2603
rect 816 2592 818 2614
rect 822 2608 828 2609
rect 822 2604 823 2608
rect 827 2604 828 2608
rect 822 2603 828 2604
rect 814 2591 820 2592
rect 814 2587 815 2591
rect 819 2587 820 2591
rect 814 2586 820 2587
rect 824 2575 826 2603
rect 904 2592 906 2686
rect 918 2681 924 2682
rect 918 2677 919 2681
rect 923 2677 924 2681
rect 918 2676 924 2677
rect 1006 2681 1012 2682
rect 1006 2677 1007 2681
rect 1011 2677 1012 2681
rect 1006 2676 1012 2677
rect 920 2651 922 2676
rect 1008 2651 1010 2676
rect 911 2650 915 2651
rect 911 2645 915 2646
rect 919 2650 923 2651
rect 919 2645 923 2646
rect 999 2650 1003 2651
rect 999 2645 1003 2646
rect 1007 2650 1011 2651
rect 1007 2645 1011 2646
rect 912 2628 914 2645
rect 1000 2628 1002 2645
rect 910 2627 916 2628
rect 910 2623 911 2627
rect 915 2623 916 2627
rect 910 2622 916 2623
rect 998 2627 1004 2628
rect 998 2623 999 2627
rect 1003 2623 1004 2627
rect 998 2622 1004 2623
rect 1080 2620 1082 2702
rect 1096 2701 1098 2717
rect 1166 2715 1172 2716
rect 1166 2711 1167 2715
rect 1171 2711 1172 2715
rect 1166 2710 1172 2711
rect 1094 2700 1100 2701
rect 1094 2696 1095 2700
rect 1099 2696 1100 2700
rect 1094 2695 1100 2696
rect 1168 2692 1170 2710
rect 1176 2692 1178 2718
rect 1183 2717 1187 2718
rect 1199 2722 1203 2723
rect 1199 2717 1203 2718
rect 1319 2722 1323 2723
rect 1319 2717 1323 2718
rect 1767 2722 1771 2723
rect 1806 2720 1807 2724
rect 1811 2720 1812 2724
rect 1886 2721 1887 2725
rect 1891 2721 1892 2725
rect 1886 2720 1892 2721
rect 1806 2719 1812 2720
rect 1767 2717 1771 2718
rect 1184 2701 1186 2717
rect 1182 2700 1188 2701
rect 1182 2696 1183 2700
rect 1187 2696 1188 2700
rect 1768 2698 1770 2717
rect 1808 2703 1810 2719
rect 1888 2703 1890 2720
rect 1807 2702 1811 2703
rect 1182 2695 1188 2696
rect 1766 2697 1772 2698
rect 1807 2697 1811 2698
rect 1831 2702 1835 2703
rect 1831 2697 1835 2698
rect 1887 2702 1891 2703
rect 1887 2697 1891 2698
rect 1766 2693 1767 2697
rect 1771 2693 1772 2697
rect 1766 2692 1772 2693
rect 1166 2691 1172 2692
rect 1166 2687 1167 2691
rect 1171 2687 1172 2691
rect 1166 2686 1172 2687
rect 1174 2691 1180 2692
rect 1174 2687 1175 2691
rect 1179 2687 1180 2691
rect 1174 2686 1180 2687
rect 1094 2681 1100 2682
rect 1094 2677 1095 2681
rect 1099 2677 1100 2681
rect 1094 2676 1100 2677
rect 1182 2681 1188 2682
rect 1808 2681 1810 2697
rect 1182 2677 1183 2681
rect 1187 2677 1188 2681
rect 1182 2676 1188 2677
rect 1766 2680 1772 2681
rect 1766 2676 1767 2680
rect 1771 2676 1772 2680
rect 1096 2651 1098 2676
rect 1184 2651 1186 2676
rect 1766 2675 1772 2676
rect 1806 2680 1812 2681
rect 1832 2680 1834 2697
rect 1806 2676 1807 2680
rect 1811 2676 1812 2680
rect 1806 2675 1812 2676
rect 1830 2679 1836 2680
rect 1830 2675 1831 2679
rect 1835 2675 1836 2679
rect 1768 2651 1770 2675
rect 1830 2674 1836 2675
rect 1904 2672 1906 2754
rect 1960 2736 1962 2754
rect 2032 2745 2034 2761
rect 2102 2759 2108 2760
rect 2102 2755 2103 2759
rect 2107 2755 2108 2759
rect 2102 2754 2108 2755
rect 2030 2744 2036 2745
rect 2030 2740 2031 2744
rect 2035 2740 2036 2744
rect 2030 2739 2036 2740
rect 2104 2736 2106 2754
rect 2184 2745 2186 2761
rect 2182 2744 2188 2745
rect 2182 2740 2183 2744
rect 2187 2740 2188 2744
rect 2182 2739 2188 2740
rect 2256 2736 2258 2770
rect 2368 2767 2370 2787
rect 2432 2776 2434 2866
rect 2470 2861 2476 2862
rect 2470 2857 2471 2861
rect 2475 2857 2476 2861
rect 2470 2856 2476 2857
rect 2472 2835 2474 2856
rect 2471 2834 2475 2835
rect 2471 2829 2475 2830
rect 2487 2834 2491 2835
rect 2487 2829 2491 2830
rect 2488 2812 2490 2829
rect 2486 2811 2492 2812
rect 2486 2807 2487 2811
rect 2491 2807 2492 2811
rect 2486 2806 2492 2807
rect 2560 2804 2562 2890
rect 2576 2881 2578 2897
rect 2646 2895 2652 2896
rect 2646 2891 2647 2895
rect 2651 2891 2652 2895
rect 2646 2890 2652 2891
rect 2574 2880 2580 2881
rect 2574 2876 2575 2880
rect 2579 2876 2580 2880
rect 2574 2875 2580 2876
rect 2648 2872 2650 2890
rect 2680 2881 2682 2897
rect 2750 2895 2756 2896
rect 2750 2891 2751 2895
rect 2755 2891 2756 2895
rect 2750 2890 2756 2891
rect 2678 2880 2684 2881
rect 2678 2876 2679 2880
rect 2683 2876 2684 2880
rect 2678 2875 2684 2876
rect 2752 2872 2754 2890
rect 2784 2881 2786 2897
rect 2782 2880 2788 2881
rect 2782 2876 2783 2880
rect 2787 2876 2788 2880
rect 2782 2875 2788 2876
rect 2856 2872 2858 2910
rect 3464 2903 3466 2930
rect 3463 2902 3467 2903
rect 3463 2897 3467 2898
rect 3464 2878 3466 2897
rect 3462 2877 3468 2878
rect 3462 2873 3463 2877
rect 3467 2873 3468 2877
rect 3462 2872 3468 2873
rect 2646 2871 2652 2872
rect 2646 2867 2647 2871
rect 2651 2867 2652 2871
rect 2646 2866 2652 2867
rect 2750 2871 2756 2872
rect 2750 2867 2751 2871
rect 2755 2867 2756 2871
rect 2750 2866 2756 2867
rect 2854 2871 2860 2872
rect 2854 2867 2855 2871
rect 2859 2867 2860 2871
rect 2854 2866 2860 2867
rect 2574 2861 2580 2862
rect 2574 2857 2575 2861
rect 2579 2857 2580 2861
rect 2574 2856 2580 2857
rect 2678 2861 2684 2862
rect 2678 2857 2679 2861
rect 2683 2857 2684 2861
rect 2678 2856 2684 2857
rect 2782 2861 2788 2862
rect 2782 2857 2783 2861
rect 2787 2857 2788 2861
rect 2782 2856 2788 2857
rect 3462 2860 3468 2861
rect 3462 2856 3463 2860
rect 3467 2856 3468 2860
rect 2576 2835 2578 2856
rect 2680 2835 2682 2856
rect 2784 2835 2786 2856
rect 3462 2855 3468 2856
rect 3464 2835 3466 2855
rect 2575 2834 2579 2835
rect 2575 2829 2579 2830
rect 2607 2834 2611 2835
rect 2607 2829 2611 2830
rect 2679 2834 2683 2835
rect 2679 2829 2683 2830
rect 2719 2834 2723 2835
rect 2719 2829 2723 2830
rect 2783 2834 2787 2835
rect 2783 2829 2787 2830
rect 2839 2834 2843 2835
rect 2839 2829 2843 2830
rect 2959 2834 2963 2835
rect 2959 2829 2963 2830
rect 3463 2834 3467 2835
rect 3463 2829 3467 2830
rect 2608 2812 2610 2829
rect 2720 2812 2722 2829
rect 2840 2812 2842 2829
rect 2960 2812 2962 2829
rect 3464 2813 3466 2829
rect 3462 2812 3468 2813
rect 2606 2811 2612 2812
rect 2606 2807 2607 2811
rect 2611 2807 2612 2811
rect 2606 2806 2612 2807
rect 2718 2811 2724 2812
rect 2718 2807 2719 2811
rect 2723 2807 2724 2811
rect 2718 2806 2724 2807
rect 2838 2811 2844 2812
rect 2838 2807 2839 2811
rect 2843 2807 2844 2811
rect 2838 2806 2844 2807
rect 2958 2811 2964 2812
rect 2958 2807 2959 2811
rect 2963 2807 2964 2811
rect 3462 2808 3463 2812
rect 3467 2808 3468 2812
rect 3462 2807 3468 2808
rect 2958 2806 2964 2807
rect 2558 2803 2564 2804
rect 2438 2799 2444 2800
rect 2438 2795 2439 2799
rect 2443 2795 2444 2799
rect 2558 2799 2559 2803
rect 2563 2799 2564 2803
rect 2558 2798 2564 2799
rect 2686 2803 2692 2804
rect 2686 2799 2687 2803
rect 2691 2799 2692 2803
rect 2918 2803 2924 2804
rect 2686 2798 2692 2799
rect 2910 2799 2916 2800
rect 2438 2794 2444 2795
rect 2430 2775 2436 2776
rect 2430 2771 2431 2775
rect 2435 2771 2436 2775
rect 2430 2770 2436 2771
rect 2335 2766 2339 2767
rect 2335 2761 2339 2762
rect 2367 2766 2371 2767
rect 2367 2761 2371 2762
rect 2336 2745 2338 2761
rect 2440 2760 2442 2794
rect 2486 2792 2492 2793
rect 2486 2788 2487 2792
rect 2491 2788 2492 2792
rect 2486 2787 2492 2788
rect 2606 2792 2612 2793
rect 2606 2788 2607 2792
rect 2611 2788 2612 2792
rect 2606 2787 2612 2788
rect 2488 2767 2490 2787
rect 2608 2767 2610 2787
rect 2688 2776 2690 2798
rect 2910 2795 2911 2799
rect 2915 2795 2916 2799
rect 2918 2799 2919 2803
rect 2923 2799 2924 2803
rect 2918 2798 2924 2799
rect 2910 2794 2916 2795
rect 2718 2792 2724 2793
rect 2718 2788 2719 2792
rect 2723 2788 2724 2792
rect 2718 2787 2724 2788
rect 2838 2792 2844 2793
rect 2838 2788 2839 2792
rect 2843 2788 2844 2792
rect 2838 2787 2844 2788
rect 2686 2775 2692 2776
rect 2686 2771 2687 2775
rect 2691 2771 2692 2775
rect 2686 2770 2692 2771
rect 2720 2767 2722 2787
rect 2840 2767 2842 2787
rect 2912 2776 2914 2794
rect 2920 2784 2922 2798
rect 3462 2795 3468 2796
rect 2958 2792 2964 2793
rect 2958 2788 2959 2792
rect 2963 2788 2964 2792
rect 3462 2791 3463 2795
rect 3467 2791 3468 2795
rect 3462 2790 3468 2791
rect 2958 2787 2964 2788
rect 2918 2783 2924 2784
rect 2918 2779 2919 2783
rect 2923 2779 2924 2783
rect 2918 2778 2924 2779
rect 2910 2775 2916 2776
rect 2910 2771 2911 2775
rect 2915 2771 2916 2775
rect 2910 2770 2916 2771
rect 2960 2767 2962 2787
rect 3464 2767 3466 2790
rect 2479 2766 2483 2767
rect 2479 2761 2483 2762
rect 2487 2766 2491 2767
rect 2487 2761 2491 2762
rect 2607 2766 2611 2767
rect 2607 2761 2611 2762
rect 2623 2766 2627 2767
rect 2623 2761 2627 2762
rect 2719 2766 2723 2767
rect 2719 2761 2723 2762
rect 2767 2766 2771 2767
rect 2767 2761 2771 2762
rect 2839 2766 2843 2767
rect 2839 2761 2843 2762
rect 2911 2766 2915 2767
rect 2911 2761 2915 2762
rect 2959 2766 2963 2767
rect 2959 2761 2963 2762
rect 3055 2766 3059 2767
rect 3055 2761 3059 2762
rect 3463 2766 3467 2767
rect 3463 2761 3467 2762
rect 2438 2759 2444 2760
rect 2438 2755 2439 2759
rect 2443 2755 2444 2759
rect 2438 2754 2444 2755
rect 2454 2759 2460 2760
rect 2454 2755 2455 2759
rect 2459 2755 2460 2759
rect 2454 2754 2460 2755
rect 2334 2744 2340 2745
rect 2334 2740 2335 2744
rect 2339 2740 2340 2744
rect 2334 2739 2340 2740
rect 2456 2736 2458 2754
rect 2480 2745 2482 2761
rect 2624 2745 2626 2761
rect 2694 2759 2700 2760
rect 2694 2755 2695 2759
rect 2699 2755 2700 2759
rect 2694 2754 2700 2755
rect 2478 2744 2484 2745
rect 2478 2740 2479 2744
rect 2483 2740 2484 2744
rect 2478 2739 2484 2740
rect 2622 2744 2628 2745
rect 2622 2740 2623 2744
rect 2627 2740 2628 2744
rect 2622 2739 2628 2740
rect 2696 2736 2698 2754
rect 2768 2745 2770 2761
rect 2912 2745 2914 2761
rect 2990 2759 2996 2760
rect 2990 2755 2991 2759
rect 2995 2755 2996 2759
rect 2990 2754 2996 2755
rect 2766 2744 2772 2745
rect 2766 2740 2767 2744
rect 2771 2740 2772 2744
rect 2766 2739 2772 2740
rect 2910 2744 2916 2745
rect 2910 2740 2911 2744
rect 2915 2740 2916 2744
rect 2910 2739 2916 2740
rect 2992 2736 2994 2754
rect 3056 2745 3058 2761
rect 3166 2759 3172 2760
rect 3166 2755 3167 2759
rect 3171 2755 3172 2759
rect 3166 2754 3172 2755
rect 3054 2744 3060 2745
rect 3054 2740 3055 2744
rect 3059 2740 3060 2744
rect 3054 2739 3060 2740
rect 1958 2735 1964 2736
rect 1958 2731 1959 2735
rect 1963 2731 1964 2735
rect 1958 2730 1964 2731
rect 2102 2735 2108 2736
rect 2102 2731 2103 2735
rect 2107 2731 2108 2735
rect 2102 2730 2108 2731
rect 2254 2735 2260 2736
rect 2254 2731 2255 2735
rect 2259 2731 2260 2735
rect 2254 2730 2260 2731
rect 2454 2735 2460 2736
rect 2454 2731 2455 2735
rect 2459 2731 2460 2735
rect 2454 2730 2460 2731
rect 2542 2735 2548 2736
rect 2542 2731 2543 2735
rect 2547 2731 2548 2735
rect 2542 2730 2548 2731
rect 2694 2735 2700 2736
rect 2694 2731 2695 2735
rect 2699 2731 2700 2735
rect 2694 2730 2700 2731
rect 2990 2735 2996 2736
rect 2990 2731 2991 2735
rect 2995 2731 2996 2735
rect 2990 2730 2996 2731
rect 2030 2725 2036 2726
rect 2030 2721 2031 2725
rect 2035 2721 2036 2725
rect 2030 2720 2036 2721
rect 2182 2725 2188 2726
rect 2182 2721 2183 2725
rect 2187 2721 2188 2725
rect 2182 2720 2188 2721
rect 2334 2725 2340 2726
rect 2334 2721 2335 2725
rect 2339 2721 2340 2725
rect 2334 2720 2340 2721
rect 2478 2725 2484 2726
rect 2478 2721 2479 2725
rect 2483 2721 2484 2725
rect 2478 2720 2484 2721
rect 2032 2703 2034 2720
rect 2184 2703 2186 2720
rect 2336 2703 2338 2720
rect 2480 2703 2482 2720
rect 2023 2702 2027 2703
rect 2023 2697 2027 2698
rect 2031 2702 2035 2703
rect 2031 2697 2035 2698
rect 2183 2702 2187 2703
rect 2183 2697 2187 2698
rect 2231 2702 2235 2703
rect 2231 2697 2235 2698
rect 2335 2702 2339 2703
rect 2335 2697 2339 2698
rect 2431 2702 2435 2703
rect 2431 2697 2435 2698
rect 2479 2702 2483 2703
rect 2479 2697 2483 2698
rect 2024 2680 2026 2697
rect 2232 2680 2234 2697
rect 2432 2680 2434 2697
rect 2022 2679 2028 2680
rect 2022 2675 2023 2679
rect 2027 2675 2028 2679
rect 2022 2674 2028 2675
rect 2230 2679 2236 2680
rect 2230 2675 2231 2679
rect 2235 2675 2236 2679
rect 2230 2674 2236 2675
rect 2430 2679 2436 2680
rect 2430 2675 2431 2679
rect 2435 2675 2436 2679
rect 2430 2674 2436 2675
rect 1902 2671 1908 2672
rect 1902 2667 1903 2671
rect 1907 2667 1908 2671
rect 1902 2666 1908 2667
rect 1910 2671 1916 2672
rect 1910 2667 1911 2671
rect 1915 2667 1916 2671
rect 1910 2666 1916 2667
rect 2102 2671 2108 2672
rect 2102 2667 2103 2671
rect 2107 2667 2108 2671
rect 2102 2666 2108 2667
rect 2414 2671 2420 2672
rect 2414 2667 2415 2671
rect 2419 2667 2420 2671
rect 2414 2666 2420 2667
rect 1806 2663 1812 2664
rect 1806 2659 1807 2663
rect 1811 2659 1812 2663
rect 1806 2658 1812 2659
rect 1830 2660 1836 2661
rect 1087 2650 1091 2651
rect 1087 2645 1091 2646
rect 1095 2650 1099 2651
rect 1095 2645 1099 2646
rect 1183 2650 1187 2651
rect 1183 2645 1187 2646
rect 1767 2650 1771 2651
rect 1767 2645 1771 2646
rect 1088 2628 1090 2645
rect 1768 2629 1770 2645
rect 1808 2635 1810 2658
rect 1830 2656 1831 2660
rect 1835 2656 1836 2660
rect 1830 2655 1836 2656
rect 1832 2635 1834 2655
rect 1912 2644 1914 2666
rect 2022 2660 2028 2661
rect 2022 2656 2023 2660
rect 2027 2656 2028 2660
rect 2022 2655 2028 2656
rect 1910 2643 1916 2644
rect 1910 2639 1911 2643
rect 1915 2639 1916 2643
rect 1910 2638 1916 2639
rect 2024 2635 2026 2655
rect 2104 2644 2106 2666
rect 2230 2660 2236 2661
rect 2230 2656 2231 2660
rect 2235 2656 2236 2660
rect 2230 2655 2236 2656
rect 2102 2643 2108 2644
rect 2102 2639 2103 2643
rect 2107 2639 2108 2643
rect 2102 2638 2108 2639
rect 2232 2635 2234 2655
rect 2254 2643 2260 2644
rect 2254 2639 2255 2643
rect 2259 2639 2260 2643
rect 2254 2638 2260 2639
rect 1807 2634 1811 2635
rect 1807 2629 1811 2630
rect 1831 2634 1835 2635
rect 1831 2629 1835 2630
rect 1999 2634 2003 2635
rect 1999 2629 2003 2630
rect 2023 2634 2027 2635
rect 2023 2629 2027 2630
rect 2183 2634 2187 2635
rect 2183 2629 2187 2630
rect 2231 2634 2235 2635
rect 2231 2629 2235 2630
rect 1766 2628 1772 2629
rect 1086 2627 1092 2628
rect 1086 2623 1087 2627
rect 1091 2623 1092 2627
rect 1766 2624 1767 2628
rect 1771 2624 1772 2628
rect 1766 2623 1772 2624
rect 1798 2627 1804 2628
rect 1798 2623 1799 2627
rect 1803 2623 1804 2627
rect 1086 2622 1092 2623
rect 1798 2622 1804 2623
rect 1078 2619 1084 2620
rect 982 2615 988 2616
rect 982 2611 983 2615
rect 987 2611 988 2615
rect 982 2610 988 2611
rect 1070 2615 1076 2616
rect 1070 2611 1071 2615
rect 1075 2611 1076 2615
rect 1078 2615 1079 2619
rect 1083 2615 1084 2619
rect 1078 2614 1084 2615
rect 1070 2610 1076 2611
rect 1766 2611 1772 2612
rect 910 2608 916 2609
rect 910 2604 911 2608
rect 915 2604 916 2608
rect 910 2603 916 2604
rect 902 2591 908 2592
rect 902 2587 903 2591
rect 907 2587 908 2591
rect 902 2586 908 2587
rect 838 2583 844 2584
rect 838 2579 839 2583
rect 843 2579 844 2583
rect 838 2578 844 2579
rect 559 2574 563 2575
rect 559 2569 563 2570
rect 591 2574 595 2575
rect 591 2569 595 2570
rect 647 2574 651 2575
rect 647 2569 651 2570
rect 679 2574 683 2575
rect 679 2569 683 2570
rect 735 2574 739 2575
rect 735 2569 739 2570
rect 767 2574 771 2575
rect 767 2569 771 2570
rect 823 2574 827 2575
rect 823 2569 827 2570
rect 542 2567 548 2568
rect 542 2563 543 2567
rect 547 2563 548 2567
rect 542 2562 548 2563
rect 574 2567 580 2568
rect 574 2563 575 2567
rect 579 2563 580 2567
rect 574 2562 580 2563
rect 310 2552 316 2553
rect 310 2548 311 2552
rect 315 2548 316 2552
rect 310 2547 316 2548
rect 406 2552 412 2553
rect 406 2548 407 2552
rect 411 2548 412 2552
rect 406 2547 412 2548
rect 502 2552 508 2553
rect 502 2548 503 2552
rect 507 2548 508 2552
rect 502 2547 508 2548
rect 576 2544 578 2562
rect 592 2553 594 2569
rect 680 2553 682 2569
rect 750 2567 756 2568
rect 750 2563 751 2567
rect 755 2563 756 2567
rect 750 2562 756 2563
rect 590 2552 596 2553
rect 590 2548 591 2552
rect 595 2548 596 2552
rect 590 2547 596 2548
rect 678 2552 684 2553
rect 678 2548 679 2552
rect 683 2548 684 2552
rect 678 2547 684 2548
rect 752 2544 754 2562
rect 768 2553 770 2569
rect 806 2559 812 2560
rect 806 2555 807 2559
rect 811 2555 812 2559
rect 806 2554 812 2555
rect 766 2552 772 2553
rect 766 2548 767 2552
rect 771 2548 772 2552
rect 766 2547 772 2548
rect 294 2543 300 2544
rect 294 2539 295 2543
rect 299 2539 300 2543
rect 294 2538 300 2539
rect 382 2543 388 2544
rect 382 2539 383 2543
rect 387 2539 388 2543
rect 382 2538 388 2539
rect 574 2543 580 2544
rect 574 2539 575 2543
rect 579 2539 580 2543
rect 574 2538 580 2539
rect 750 2543 756 2544
rect 750 2539 751 2543
rect 755 2539 756 2543
rect 750 2538 756 2539
rect 222 2533 228 2534
rect 110 2532 116 2533
rect 110 2528 111 2532
rect 115 2528 116 2532
rect 222 2529 223 2533
rect 227 2529 228 2533
rect 222 2528 228 2529
rect 310 2533 316 2534
rect 310 2529 311 2533
rect 315 2529 316 2533
rect 310 2528 316 2529
rect 110 2527 116 2528
rect 112 2511 114 2527
rect 224 2511 226 2528
rect 312 2511 314 2528
rect 111 2510 115 2511
rect 111 2505 115 2506
rect 135 2510 139 2511
rect 135 2505 139 2506
rect 223 2510 227 2511
rect 223 2505 227 2506
rect 247 2510 251 2511
rect 247 2505 251 2506
rect 311 2510 315 2511
rect 311 2505 315 2506
rect 112 2489 114 2505
rect 110 2488 116 2489
rect 136 2488 138 2505
rect 248 2488 250 2505
rect 110 2484 111 2488
rect 115 2484 116 2488
rect 110 2483 116 2484
rect 134 2487 140 2488
rect 134 2483 135 2487
rect 139 2483 140 2487
rect 134 2482 140 2483
rect 246 2487 252 2488
rect 246 2483 247 2487
rect 251 2483 252 2487
rect 246 2482 252 2483
rect 214 2479 220 2480
rect 206 2475 212 2476
rect 110 2471 116 2472
rect 110 2467 111 2471
rect 115 2467 116 2471
rect 206 2471 207 2475
rect 211 2471 212 2475
rect 214 2475 215 2479
rect 219 2475 220 2479
rect 214 2474 220 2475
rect 206 2470 212 2471
rect 110 2466 116 2467
rect 134 2468 140 2469
rect 112 2431 114 2466
rect 134 2464 135 2468
rect 139 2464 140 2468
rect 134 2463 140 2464
rect 136 2431 138 2463
rect 111 2430 115 2431
rect 111 2425 115 2426
rect 135 2430 139 2431
rect 135 2425 139 2426
rect 112 2406 114 2425
rect 136 2409 138 2425
rect 208 2424 210 2470
rect 216 2452 218 2474
rect 246 2468 252 2469
rect 246 2464 247 2468
rect 251 2464 252 2468
rect 246 2463 252 2464
rect 214 2451 220 2452
rect 214 2447 215 2451
rect 219 2447 220 2451
rect 214 2446 220 2447
rect 248 2431 250 2463
rect 384 2452 386 2538
rect 406 2533 412 2534
rect 406 2529 407 2533
rect 411 2529 412 2533
rect 406 2528 412 2529
rect 502 2533 508 2534
rect 502 2529 503 2533
rect 507 2529 508 2533
rect 502 2528 508 2529
rect 590 2533 596 2534
rect 590 2529 591 2533
rect 595 2529 596 2533
rect 590 2528 596 2529
rect 678 2533 684 2534
rect 678 2529 679 2533
rect 683 2529 684 2533
rect 678 2528 684 2529
rect 766 2533 772 2534
rect 766 2529 767 2533
rect 771 2529 772 2533
rect 766 2528 772 2529
rect 408 2511 410 2528
rect 504 2511 506 2528
rect 592 2511 594 2528
rect 680 2511 682 2528
rect 768 2511 770 2528
rect 391 2510 395 2511
rect 391 2505 395 2506
rect 407 2510 411 2511
rect 407 2505 411 2506
rect 503 2510 507 2511
rect 503 2505 507 2506
rect 543 2510 547 2511
rect 543 2505 547 2506
rect 591 2510 595 2511
rect 591 2505 595 2506
rect 679 2510 683 2511
rect 679 2505 683 2506
rect 695 2510 699 2511
rect 695 2505 699 2506
rect 767 2510 771 2511
rect 767 2505 771 2506
rect 392 2488 394 2505
rect 544 2488 546 2505
rect 696 2488 698 2505
rect 390 2487 396 2488
rect 390 2483 391 2487
rect 395 2483 396 2487
rect 390 2482 396 2483
rect 542 2487 548 2488
rect 542 2483 543 2487
rect 547 2483 548 2487
rect 542 2482 548 2483
rect 694 2487 700 2488
rect 694 2483 695 2487
rect 699 2483 700 2487
rect 694 2482 700 2483
rect 808 2480 810 2554
rect 840 2544 842 2578
rect 912 2575 914 2603
rect 984 2592 986 2610
rect 998 2608 1004 2609
rect 998 2604 999 2608
rect 1003 2604 1004 2608
rect 998 2603 1004 2604
rect 982 2591 988 2592
rect 982 2587 983 2591
rect 987 2587 988 2591
rect 982 2586 988 2587
rect 1000 2575 1002 2603
rect 1072 2592 1074 2610
rect 1086 2608 1092 2609
rect 1086 2604 1087 2608
rect 1091 2604 1092 2608
rect 1766 2607 1767 2611
rect 1771 2607 1772 2611
rect 1766 2606 1772 2607
rect 1086 2603 1092 2604
rect 1070 2591 1076 2592
rect 1070 2587 1071 2591
rect 1075 2587 1076 2591
rect 1070 2586 1076 2587
rect 1088 2575 1090 2603
rect 1768 2575 1770 2606
rect 855 2574 859 2575
rect 855 2569 859 2570
rect 911 2574 915 2575
rect 911 2569 915 2570
rect 943 2574 947 2575
rect 943 2569 947 2570
rect 999 2574 1003 2575
rect 999 2569 1003 2570
rect 1031 2574 1035 2575
rect 1031 2569 1035 2570
rect 1087 2574 1091 2575
rect 1087 2569 1091 2570
rect 1119 2574 1123 2575
rect 1119 2569 1123 2570
rect 1215 2574 1219 2575
rect 1215 2569 1219 2570
rect 1311 2574 1315 2575
rect 1311 2569 1315 2570
rect 1407 2574 1411 2575
rect 1407 2569 1411 2570
rect 1495 2574 1499 2575
rect 1495 2569 1499 2570
rect 1583 2574 1587 2575
rect 1583 2569 1587 2570
rect 1671 2574 1675 2575
rect 1671 2569 1675 2570
rect 1767 2574 1771 2575
rect 1767 2569 1771 2570
rect 856 2553 858 2569
rect 926 2567 932 2568
rect 926 2563 927 2567
rect 931 2563 932 2567
rect 926 2562 932 2563
rect 854 2552 860 2553
rect 854 2548 855 2552
rect 859 2548 860 2552
rect 854 2547 860 2548
rect 928 2544 930 2562
rect 944 2553 946 2569
rect 1014 2567 1020 2568
rect 1014 2563 1015 2567
rect 1019 2563 1020 2567
rect 1014 2562 1020 2563
rect 942 2552 948 2553
rect 942 2548 943 2552
rect 947 2548 948 2552
rect 942 2547 948 2548
rect 1016 2544 1018 2562
rect 1032 2553 1034 2569
rect 1102 2567 1108 2568
rect 1102 2563 1103 2567
rect 1107 2563 1108 2567
rect 1102 2562 1108 2563
rect 1054 2559 1060 2560
rect 1054 2555 1055 2559
rect 1059 2555 1060 2559
rect 1054 2554 1060 2555
rect 1030 2552 1036 2553
rect 1030 2548 1031 2552
rect 1035 2548 1036 2552
rect 1030 2547 1036 2548
rect 838 2543 844 2544
rect 838 2539 839 2543
rect 843 2539 844 2543
rect 838 2538 844 2539
rect 926 2543 932 2544
rect 926 2539 927 2543
rect 931 2539 932 2543
rect 926 2538 932 2539
rect 1014 2543 1020 2544
rect 1014 2539 1015 2543
rect 1019 2539 1020 2543
rect 1014 2538 1020 2539
rect 854 2533 860 2534
rect 854 2529 855 2533
rect 859 2529 860 2533
rect 854 2528 860 2529
rect 942 2533 948 2534
rect 942 2529 943 2533
rect 947 2529 948 2533
rect 942 2528 948 2529
rect 1030 2533 1036 2534
rect 1030 2529 1031 2533
rect 1035 2529 1036 2533
rect 1030 2528 1036 2529
rect 856 2511 858 2528
rect 944 2511 946 2528
rect 1032 2511 1034 2528
rect 839 2510 843 2511
rect 839 2505 843 2506
rect 855 2510 859 2511
rect 855 2505 859 2506
rect 943 2510 947 2511
rect 943 2505 947 2506
rect 975 2510 979 2511
rect 975 2505 979 2506
rect 1031 2510 1035 2511
rect 1031 2505 1035 2506
rect 840 2488 842 2505
rect 976 2488 978 2505
rect 838 2487 844 2488
rect 838 2483 839 2487
rect 843 2483 844 2487
rect 838 2482 844 2483
rect 974 2487 980 2488
rect 974 2483 975 2487
rect 979 2483 980 2487
rect 974 2482 980 2483
rect 1056 2480 1058 2554
rect 1104 2544 1106 2562
rect 1120 2553 1122 2569
rect 1190 2567 1196 2568
rect 1190 2563 1191 2567
rect 1195 2563 1196 2567
rect 1190 2562 1196 2563
rect 1118 2552 1124 2553
rect 1118 2548 1119 2552
rect 1123 2548 1124 2552
rect 1118 2547 1124 2548
rect 1192 2544 1194 2562
rect 1216 2553 1218 2569
rect 1286 2567 1292 2568
rect 1286 2563 1287 2567
rect 1291 2563 1292 2567
rect 1286 2562 1292 2563
rect 1214 2552 1220 2553
rect 1214 2548 1215 2552
rect 1219 2548 1220 2552
rect 1214 2547 1220 2548
rect 1288 2544 1290 2562
rect 1312 2553 1314 2569
rect 1408 2553 1410 2569
rect 1496 2553 1498 2569
rect 1566 2567 1572 2568
rect 1566 2563 1567 2567
rect 1571 2563 1572 2567
rect 1566 2562 1572 2563
rect 1310 2552 1316 2553
rect 1310 2548 1311 2552
rect 1315 2548 1316 2552
rect 1310 2547 1316 2548
rect 1406 2552 1412 2553
rect 1406 2548 1407 2552
rect 1411 2548 1412 2552
rect 1406 2547 1412 2548
rect 1494 2552 1500 2553
rect 1494 2548 1495 2552
rect 1499 2548 1500 2552
rect 1494 2547 1500 2548
rect 1568 2544 1570 2562
rect 1584 2553 1586 2569
rect 1654 2567 1660 2568
rect 1654 2563 1655 2567
rect 1659 2563 1660 2567
rect 1654 2562 1660 2563
rect 1582 2552 1588 2553
rect 1582 2548 1583 2552
rect 1587 2548 1588 2552
rect 1582 2547 1588 2548
rect 1656 2544 1658 2562
rect 1662 2559 1668 2560
rect 1662 2555 1663 2559
rect 1667 2555 1668 2559
rect 1662 2554 1668 2555
rect 1102 2543 1108 2544
rect 1102 2539 1103 2543
rect 1107 2539 1108 2543
rect 1102 2538 1108 2539
rect 1190 2543 1196 2544
rect 1190 2539 1191 2543
rect 1195 2539 1196 2543
rect 1190 2538 1196 2539
rect 1286 2543 1292 2544
rect 1286 2539 1287 2543
rect 1291 2539 1292 2543
rect 1286 2538 1292 2539
rect 1382 2543 1388 2544
rect 1382 2539 1383 2543
rect 1387 2539 1388 2543
rect 1382 2538 1388 2539
rect 1566 2543 1572 2544
rect 1566 2539 1567 2543
rect 1571 2539 1572 2543
rect 1566 2538 1572 2539
rect 1654 2543 1660 2544
rect 1654 2539 1655 2543
rect 1659 2539 1660 2543
rect 1654 2538 1660 2539
rect 1118 2533 1124 2534
rect 1118 2529 1119 2533
rect 1123 2529 1124 2533
rect 1118 2528 1124 2529
rect 1214 2533 1220 2534
rect 1214 2529 1215 2533
rect 1219 2529 1220 2533
rect 1214 2528 1220 2529
rect 1310 2533 1316 2534
rect 1310 2529 1311 2533
rect 1315 2529 1316 2533
rect 1310 2528 1316 2529
rect 1120 2511 1122 2528
rect 1216 2511 1218 2528
rect 1312 2511 1314 2528
rect 1103 2510 1107 2511
rect 1103 2505 1107 2506
rect 1119 2510 1123 2511
rect 1119 2505 1123 2506
rect 1215 2510 1219 2511
rect 1215 2505 1219 2506
rect 1231 2510 1235 2511
rect 1231 2505 1235 2506
rect 1311 2510 1315 2511
rect 1311 2505 1315 2506
rect 1351 2510 1355 2511
rect 1351 2505 1355 2506
rect 1104 2488 1106 2505
rect 1232 2488 1234 2505
rect 1352 2488 1354 2505
rect 1102 2487 1108 2488
rect 1102 2483 1103 2487
rect 1107 2483 1108 2487
rect 1102 2482 1108 2483
rect 1230 2487 1236 2488
rect 1230 2483 1231 2487
rect 1235 2483 1236 2487
rect 1230 2482 1236 2483
rect 1350 2487 1356 2488
rect 1350 2483 1351 2487
rect 1355 2483 1356 2487
rect 1350 2482 1356 2483
rect 622 2479 628 2480
rect 462 2475 468 2476
rect 462 2471 463 2475
rect 467 2471 468 2475
rect 462 2470 468 2471
rect 614 2475 620 2476
rect 614 2471 615 2475
rect 619 2471 620 2475
rect 622 2475 623 2479
rect 627 2475 628 2479
rect 622 2474 628 2475
rect 806 2479 812 2480
rect 806 2475 807 2479
rect 811 2475 812 2479
rect 806 2474 812 2475
rect 918 2479 924 2480
rect 918 2475 919 2479
rect 923 2475 924 2479
rect 918 2474 924 2475
rect 1054 2479 1060 2480
rect 1054 2475 1055 2479
rect 1059 2475 1060 2479
rect 1054 2474 1060 2475
rect 1182 2479 1188 2480
rect 1182 2475 1183 2479
rect 1187 2475 1188 2479
rect 1182 2474 1188 2475
rect 1310 2479 1316 2480
rect 1310 2475 1311 2479
rect 1315 2475 1316 2479
rect 1310 2474 1316 2475
rect 614 2470 620 2471
rect 390 2468 396 2469
rect 390 2464 391 2468
rect 395 2464 396 2468
rect 390 2463 396 2464
rect 382 2451 388 2452
rect 382 2447 383 2451
rect 387 2447 388 2451
rect 382 2446 388 2447
rect 392 2431 394 2463
rect 464 2452 466 2470
rect 542 2468 548 2469
rect 542 2464 543 2468
rect 547 2464 548 2468
rect 542 2463 548 2464
rect 462 2451 468 2452
rect 462 2447 463 2451
rect 467 2447 468 2451
rect 462 2446 468 2447
rect 544 2431 546 2463
rect 616 2452 618 2470
rect 624 2460 626 2474
rect 694 2468 700 2469
rect 694 2464 695 2468
rect 699 2464 700 2468
rect 694 2463 700 2464
rect 838 2468 844 2469
rect 838 2464 839 2468
rect 843 2464 844 2468
rect 838 2463 844 2464
rect 622 2459 628 2460
rect 622 2455 623 2459
rect 627 2455 628 2459
rect 622 2454 628 2455
rect 614 2451 620 2452
rect 614 2447 615 2451
rect 619 2447 620 2451
rect 614 2446 620 2447
rect 696 2431 698 2463
rect 840 2431 842 2463
rect 920 2452 922 2474
rect 974 2468 980 2469
rect 974 2464 975 2468
rect 979 2464 980 2468
rect 974 2463 980 2464
rect 1102 2468 1108 2469
rect 1102 2464 1103 2468
rect 1107 2464 1108 2468
rect 1102 2463 1108 2464
rect 918 2451 924 2452
rect 918 2447 919 2451
rect 923 2447 924 2451
rect 918 2446 924 2447
rect 976 2431 978 2463
rect 1030 2451 1036 2452
rect 1030 2447 1031 2451
rect 1035 2447 1036 2451
rect 1030 2446 1036 2447
rect 239 2430 243 2431
rect 239 2425 243 2426
rect 247 2430 251 2431
rect 247 2425 251 2426
rect 391 2430 395 2431
rect 391 2425 395 2426
rect 543 2430 547 2431
rect 543 2425 547 2426
rect 551 2430 555 2431
rect 551 2425 555 2426
rect 695 2430 699 2431
rect 695 2425 699 2426
rect 719 2430 723 2431
rect 719 2425 723 2426
rect 839 2430 843 2431
rect 839 2425 843 2426
rect 895 2430 899 2431
rect 895 2425 899 2426
rect 975 2430 979 2431
rect 975 2425 979 2426
rect 206 2423 212 2424
rect 206 2419 207 2423
rect 211 2419 212 2423
rect 206 2418 212 2419
rect 240 2409 242 2425
rect 310 2423 316 2424
rect 310 2419 311 2423
rect 315 2419 316 2423
rect 310 2418 316 2419
rect 134 2408 140 2409
rect 110 2405 116 2406
rect 110 2401 111 2405
rect 115 2401 116 2405
rect 134 2404 135 2408
rect 139 2404 140 2408
rect 134 2403 140 2404
rect 238 2408 244 2409
rect 238 2404 239 2408
rect 243 2404 244 2408
rect 238 2403 244 2404
rect 110 2400 116 2401
rect 312 2400 314 2418
rect 392 2409 394 2425
rect 462 2423 468 2424
rect 462 2419 463 2423
rect 467 2419 468 2423
rect 462 2418 468 2419
rect 390 2408 396 2409
rect 390 2404 391 2408
rect 395 2404 396 2408
rect 390 2403 396 2404
rect 464 2400 466 2418
rect 552 2409 554 2425
rect 622 2423 628 2424
rect 622 2419 623 2423
rect 627 2419 628 2423
rect 622 2418 628 2419
rect 550 2408 556 2409
rect 550 2404 551 2408
rect 555 2404 556 2408
rect 550 2403 556 2404
rect 624 2400 626 2418
rect 720 2409 722 2425
rect 896 2409 898 2425
rect 918 2423 924 2424
rect 918 2419 919 2423
rect 923 2419 924 2423
rect 918 2418 924 2419
rect 966 2423 972 2424
rect 966 2419 967 2423
rect 971 2419 972 2423
rect 966 2418 972 2419
rect 718 2408 724 2409
rect 718 2404 719 2408
rect 723 2404 724 2408
rect 718 2403 724 2404
rect 894 2408 900 2409
rect 894 2404 895 2408
rect 899 2404 900 2408
rect 894 2403 900 2404
rect 310 2399 316 2400
rect 310 2395 311 2399
rect 315 2395 316 2399
rect 310 2394 316 2395
rect 462 2399 468 2400
rect 462 2395 463 2399
rect 467 2395 468 2399
rect 462 2394 468 2395
rect 622 2399 628 2400
rect 622 2395 623 2399
rect 627 2395 628 2399
rect 622 2394 628 2395
rect 630 2399 636 2400
rect 630 2395 631 2399
rect 635 2395 636 2399
rect 630 2394 636 2395
rect 134 2389 140 2390
rect 110 2388 116 2389
rect 110 2384 111 2388
rect 115 2384 116 2388
rect 134 2385 135 2389
rect 139 2385 140 2389
rect 134 2384 140 2385
rect 238 2389 244 2390
rect 238 2385 239 2389
rect 243 2385 244 2389
rect 238 2384 244 2385
rect 390 2389 396 2390
rect 390 2385 391 2389
rect 395 2385 396 2389
rect 390 2384 396 2385
rect 550 2389 556 2390
rect 550 2385 551 2389
rect 555 2385 556 2389
rect 550 2384 556 2385
rect 110 2383 116 2384
rect 112 2359 114 2383
rect 136 2359 138 2384
rect 240 2359 242 2384
rect 392 2359 394 2384
rect 552 2359 554 2384
rect 111 2358 115 2359
rect 111 2353 115 2354
rect 135 2358 139 2359
rect 135 2353 139 2354
rect 239 2358 243 2359
rect 239 2353 243 2354
rect 375 2358 379 2359
rect 375 2353 379 2354
rect 391 2358 395 2359
rect 391 2353 395 2354
rect 479 2358 483 2359
rect 479 2353 483 2354
rect 551 2358 555 2359
rect 551 2353 555 2354
rect 599 2358 603 2359
rect 599 2353 603 2354
rect 112 2337 114 2353
rect 110 2336 116 2337
rect 376 2336 378 2353
rect 480 2336 482 2353
rect 600 2336 602 2353
rect 110 2332 111 2336
rect 115 2332 116 2336
rect 110 2331 116 2332
rect 374 2335 380 2336
rect 374 2331 375 2335
rect 379 2331 380 2335
rect 374 2330 380 2331
rect 478 2335 484 2336
rect 478 2331 479 2335
rect 483 2331 484 2335
rect 478 2330 484 2331
rect 598 2335 604 2336
rect 598 2331 599 2335
rect 603 2331 604 2335
rect 598 2330 604 2331
rect 446 2323 452 2324
rect 110 2319 116 2320
rect 110 2315 111 2319
rect 115 2315 116 2319
rect 446 2319 447 2323
rect 451 2319 452 2323
rect 446 2318 452 2319
rect 550 2323 556 2324
rect 550 2319 551 2323
rect 555 2319 556 2323
rect 550 2318 556 2319
rect 110 2314 116 2315
rect 374 2316 380 2317
rect 112 2287 114 2314
rect 374 2312 375 2316
rect 379 2312 380 2316
rect 374 2311 380 2312
rect 376 2287 378 2311
rect 448 2300 450 2318
rect 478 2316 484 2317
rect 478 2312 479 2316
rect 483 2312 484 2316
rect 478 2311 484 2312
rect 446 2299 452 2300
rect 446 2295 447 2299
rect 451 2295 452 2299
rect 446 2294 452 2295
rect 480 2287 482 2311
rect 552 2300 554 2318
rect 598 2316 604 2317
rect 598 2312 599 2316
rect 603 2312 604 2316
rect 598 2311 604 2312
rect 550 2299 556 2300
rect 550 2295 551 2299
rect 555 2295 556 2299
rect 550 2294 556 2295
rect 600 2287 602 2311
rect 632 2308 634 2394
rect 718 2389 724 2390
rect 718 2385 719 2389
rect 723 2385 724 2389
rect 718 2384 724 2385
rect 894 2389 900 2390
rect 894 2385 895 2389
rect 899 2385 900 2389
rect 894 2384 900 2385
rect 720 2359 722 2384
rect 896 2359 898 2384
rect 719 2358 723 2359
rect 719 2353 723 2354
rect 847 2358 851 2359
rect 847 2353 851 2354
rect 895 2358 899 2359
rect 895 2353 899 2354
rect 720 2336 722 2353
rect 848 2336 850 2353
rect 718 2335 724 2336
rect 718 2331 719 2335
rect 723 2331 724 2335
rect 718 2330 724 2331
rect 846 2335 852 2336
rect 846 2331 847 2335
rect 851 2331 852 2335
rect 846 2330 852 2331
rect 920 2328 922 2418
rect 968 2400 970 2418
rect 1032 2400 1034 2446
rect 1104 2431 1106 2463
rect 1184 2452 1186 2474
rect 1230 2468 1236 2469
rect 1230 2464 1231 2468
rect 1235 2464 1236 2468
rect 1230 2463 1236 2464
rect 1182 2451 1188 2452
rect 1182 2447 1183 2451
rect 1187 2447 1188 2451
rect 1182 2446 1188 2447
rect 1232 2431 1234 2463
rect 1312 2452 1314 2474
rect 1350 2468 1356 2469
rect 1350 2464 1351 2468
rect 1355 2464 1356 2468
rect 1350 2463 1356 2464
rect 1310 2451 1316 2452
rect 1310 2447 1311 2451
rect 1315 2447 1316 2451
rect 1310 2446 1316 2447
rect 1334 2451 1340 2452
rect 1334 2447 1335 2451
rect 1339 2447 1340 2451
rect 1334 2446 1340 2447
rect 1063 2430 1067 2431
rect 1063 2425 1067 2426
rect 1103 2430 1107 2431
rect 1103 2425 1107 2426
rect 1231 2430 1235 2431
rect 1231 2425 1235 2426
rect 1239 2430 1243 2431
rect 1239 2425 1243 2426
rect 1064 2409 1066 2425
rect 1240 2409 1242 2425
rect 1318 2423 1324 2424
rect 1318 2419 1319 2423
rect 1323 2419 1324 2423
rect 1318 2418 1324 2419
rect 1062 2408 1068 2409
rect 1062 2404 1063 2408
rect 1067 2404 1068 2408
rect 1062 2403 1068 2404
rect 1238 2408 1244 2409
rect 1238 2404 1239 2408
rect 1243 2404 1244 2408
rect 1238 2403 1244 2404
rect 1320 2400 1322 2418
rect 1336 2408 1338 2446
rect 1352 2431 1354 2463
rect 1384 2460 1386 2538
rect 1406 2533 1412 2534
rect 1406 2529 1407 2533
rect 1411 2529 1412 2533
rect 1406 2528 1412 2529
rect 1494 2533 1500 2534
rect 1494 2529 1495 2533
rect 1499 2529 1500 2533
rect 1494 2528 1500 2529
rect 1582 2533 1588 2534
rect 1582 2529 1583 2533
rect 1587 2529 1588 2533
rect 1582 2528 1588 2529
rect 1408 2511 1410 2528
rect 1496 2511 1498 2528
rect 1584 2511 1586 2528
rect 1407 2510 1411 2511
rect 1407 2505 1411 2506
rect 1463 2510 1467 2511
rect 1463 2505 1467 2506
rect 1495 2510 1499 2511
rect 1495 2505 1499 2506
rect 1575 2510 1579 2511
rect 1575 2505 1579 2506
rect 1583 2510 1587 2511
rect 1583 2505 1587 2506
rect 1464 2488 1466 2505
rect 1576 2488 1578 2505
rect 1462 2487 1468 2488
rect 1462 2483 1463 2487
rect 1467 2483 1468 2487
rect 1462 2482 1468 2483
rect 1574 2487 1580 2488
rect 1574 2483 1575 2487
rect 1579 2483 1580 2487
rect 1574 2482 1580 2483
rect 1664 2480 1666 2554
rect 1672 2553 1674 2569
rect 1670 2552 1676 2553
rect 1670 2548 1671 2552
rect 1675 2548 1676 2552
rect 1768 2550 1770 2569
rect 1670 2547 1676 2548
rect 1766 2549 1772 2550
rect 1766 2545 1767 2549
rect 1771 2545 1772 2549
rect 1766 2544 1772 2545
rect 1800 2544 1802 2622
rect 1808 2610 1810 2629
rect 1832 2613 1834 2629
rect 1902 2627 1908 2628
rect 1902 2623 1903 2627
rect 1907 2623 1908 2627
rect 1902 2622 1908 2623
rect 1830 2612 1836 2613
rect 1806 2609 1812 2610
rect 1806 2605 1807 2609
rect 1811 2605 1812 2609
rect 1830 2608 1831 2612
rect 1835 2608 1836 2612
rect 1830 2607 1836 2608
rect 1806 2604 1812 2605
rect 1904 2604 1906 2622
rect 2000 2613 2002 2629
rect 2070 2627 2076 2628
rect 2070 2623 2071 2627
rect 2075 2623 2076 2627
rect 2070 2622 2076 2623
rect 1998 2612 2004 2613
rect 1998 2608 1999 2612
rect 2003 2608 2004 2612
rect 1998 2607 2004 2608
rect 2072 2604 2074 2622
rect 2184 2613 2186 2629
rect 2182 2612 2188 2613
rect 2182 2608 2183 2612
rect 2187 2608 2188 2612
rect 2182 2607 2188 2608
rect 2256 2604 2258 2638
rect 2359 2634 2363 2635
rect 2359 2629 2363 2630
rect 2360 2613 2362 2629
rect 2416 2628 2418 2666
rect 2430 2660 2436 2661
rect 2430 2656 2431 2660
rect 2435 2656 2436 2660
rect 2430 2655 2436 2656
rect 2432 2635 2434 2655
rect 2544 2644 2546 2730
rect 2622 2725 2628 2726
rect 2622 2721 2623 2725
rect 2627 2721 2628 2725
rect 2622 2720 2628 2721
rect 2766 2725 2772 2726
rect 2766 2721 2767 2725
rect 2771 2721 2772 2725
rect 2766 2720 2772 2721
rect 2910 2725 2916 2726
rect 2910 2721 2911 2725
rect 2915 2721 2916 2725
rect 2910 2720 2916 2721
rect 3054 2725 3060 2726
rect 3054 2721 3055 2725
rect 3059 2721 3060 2725
rect 3054 2720 3060 2721
rect 2624 2703 2626 2720
rect 2768 2703 2770 2720
rect 2912 2703 2914 2720
rect 3056 2703 3058 2720
rect 2615 2702 2619 2703
rect 2615 2697 2619 2698
rect 2623 2702 2627 2703
rect 2623 2697 2627 2698
rect 2767 2702 2771 2703
rect 2767 2697 2771 2698
rect 2783 2702 2787 2703
rect 2783 2697 2787 2698
rect 2911 2702 2915 2703
rect 2911 2697 2915 2698
rect 2943 2702 2947 2703
rect 2943 2697 2947 2698
rect 3055 2702 3059 2703
rect 3055 2697 3059 2698
rect 3095 2702 3099 2703
rect 3095 2697 3099 2698
rect 2616 2680 2618 2697
rect 2784 2680 2786 2697
rect 2944 2680 2946 2697
rect 3096 2680 3098 2697
rect 2614 2679 2620 2680
rect 2614 2675 2615 2679
rect 2619 2675 2620 2679
rect 2614 2674 2620 2675
rect 2782 2679 2788 2680
rect 2782 2675 2783 2679
rect 2787 2675 2788 2679
rect 2782 2674 2788 2675
rect 2942 2679 2948 2680
rect 2942 2675 2943 2679
rect 2947 2675 2948 2679
rect 2942 2674 2948 2675
rect 3094 2679 3100 2680
rect 3094 2675 3095 2679
rect 3099 2675 3100 2679
rect 3094 2674 3100 2675
rect 3168 2672 3170 2754
rect 3464 2742 3466 2761
rect 3462 2741 3468 2742
rect 3462 2737 3463 2741
rect 3467 2737 3468 2741
rect 3462 2736 3468 2737
rect 3462 2724 3468 2725
rect 3462 2720 3463 2724
rect 3467 2720 3468 2724
rect 3462 2719 3468 2720
rect 3464 2703 3466 2719
rect 3239 2702 3243 2703
rect 3239 2697 3243 2698
rect 3367 2702 3371 2703
rect 3367 2697 3371 2698
rect 3463 2702 3467 2703
rect 3463 2697 3467 2698
rect 3240 2680 3242 2697
rect 3368 2680 3370 2697
rect 3464 2681 3466 2697
rect 3462 2680 3468 2681
rect 3238 2679 3244 2680
rect 3238 2675 3239 2679
rect 3243 2675 3244 2679
rect 3238 2674 3244 2675
rect 3366 2679 3372 2680
rect 3366 2675 3367 2679
rect 3371 2675 3372 2679
rect 3462 2676 3463 2680
rect 3467 2676 3468 2680
rect 3462 2675 3468 2676
rect 3366 2674 3372 2675
rect 3166 2671 3172 2672
rect 2686 2667 2692 2668
rect 2686 2663 2687 2667
rect 2691 2663 2692 2667
rect 2686 2662 2692 2663
rect 2854 2667 2860 2668
rect 2854 2663 2855 2667
rect 2859 2663 2860 2667
rect 2854 2662 2860 2663
rect 3014 2667 3020 2668
rect 3014 2663 3015 2667
rect 3019 2663 3020 2667
rect 3166 2667 3167 2671
rect 3171 2667 3172 2671
rect 3318 2671 3324 2672
rect 3166 2666 3172 2667
rect 3310 2667 3316 2668
rect 3014 2662 3020 2663
rect 3310 2663 3311 2667
rect 3315 2663 3316 2667
rect 3318 2667 3319 2671
rect 3323 2667 3324 2671
rect 3318 2666 3324 2667
rect 3310 2662 3316 2663
rect 2614 2660 2620 2661
rect 2614 2656 2615 2660
rect 2619 2656 2620 2660
rect 2614 2655 2620 2656
rect 2542 2643 2548 2644
rect 2542 2639 2543 2643
rect 2547 2639 2548 2643
rect 2542 2638 2548 2639
rect 2590 2643 2596 2644
rect 2590 2639 2591 2643
rect 2595 2639 2596 2643
rect 2590 2638 2596 2639
rect 2431 2634 2435 2635
rect 2431 2629 2435 2630
rect 2519 2634 2523 2635
rect 2519 2629 2523 2630
rect 2414 2627 2420 2628
rect 2414 2623 2415 2627
rect 2419 2623 2420 2627
rect 2414 2622 2420 2623
rect 2520 2613 2522 2629
rect 2358 2612 2364 2613
rect 2358 2608 2359 2612
rect 2363 2608 2364 2612
rect 2358 2607 2364 2608
rect 2518 2612 2524 2613
rect 2518 2608 2519 2612
rect 2523 2608 2524 2612
rect 2518 2607 2524 2608
rect 2592 2604 2594 2638
rect 2616 2635 2618 2655
rect 2688 2644 2690 2662
rect 2782 2660 2788 2661
rect 2782 2656 2783 2660
rect 2787 2656 2788 2660
rect 2782 2655 2788 2656
rect 2686 2643 2692 2644
rect 2686 2639 2687 2643
rect 2691 2639 2692 2643
rect 2686 2638 2692 2639
rect 2784 2635 2786 2655
rect 2856 2644 2858 2662
rect 2942 2660 2948 2661
rect 2942 2656 2943 2660
rect 2947 2656 2948 2660
rect 2942 2655 2948 2656
rect 2854 2643 2860 2644
rect 2854 2639 2855 2643
rect 2859 2639 2860 2643
rect 2854 2638 2860 2639
rect 2944 2635 2946 2655
rect 3016 2644 3018 2662
rect 3094 2660 3100 2661
rect 3094 2656 3095 2660
rect 3099 2656 3100 2660
rect 3094 2655 3100 2656
rect 3238 2660 3244 2661
rect 3238 2656 3239 2660
rect 3243 2656 3244 2660
rect 3238 2655 3244 2656
rect 3014 2643 3020 2644
rect 3014 2639 3015 2643
rect 3019 2639 3020 2643
rect 3014 2638 3020 2639
rect 3096 2635 3098 2655
rect 3240 2635 3242 2655
rect 2615 2634 2619 2635
rect 2615 2629 2619 2630
rect 2671 2634 2675 2635
rect 2671 2629 2675 2630
rect 2783 2634 2787 2635
rect 2783 2629 2787 2630
rect 2807 2634 2811 2635
rect 2807 2629 2811 2630
rect 2927 2634 2931 2635
rect 2927 2629 2931 2630
rect 2943 2634 2947 2635
rect 2943 2629 2947 2630
rect 3047 2634 3051 2635
rect 3047 2629 3051 2630
rect 3095 2634 3099 2635
rect 3095 2629 3099 2630
rect 3159 2634 3163 2635
rect 3159 2629 3163 2630
rect 3239 2634 3243 2635
rect 3239 2629 3243 2630
rect 3271 2634 3275 2635
rect 3271 2629 3275 2630
rect 2672 2613 2674 2629
rect 2808 2613 2810 2629
rect 2914 2627 2920 2628
rect 2914 2623 2915 2627
rect 2919 2623 2920 2627
rect 2914 2622 2920 2623
rect 2870 2619 2876 2620
rect 2870 2615 2871 2619
rect 2875 2615 2876 2619
rect 2870 2614 2876 2615
rect 2670 2612 2676 2613
rect 2670 2608 2671 2612
rect 2675 2608 2676 2612
rect 2670 2607 2676 2608
rect 2806 2612 2812 2613
rect 2806 2608 2807 2612
rect 2811 2608 2812 2612
rect 2806 2607 2812 2608
rect 1902 2603 1908 2604
rect 1902 2599 1903 2603
rect 1907 2599 1908 2603
rect 1902 2598 1908 2599
rect 2070 2603 2076 2604
rect 2070 2599 2071 2603
rect 2075 2599 2076 2603
rect 2070 2598 2076 2599
rect 2254 2603 2260 2604
rect 2254 2599 2255 2603
rect 2259 2599 2260 2603
rect 2254 2598 2260 2599
rect 2262 2603 2268 2604
rect 2262 2599 2263 2603
rect 2267 2599 2268 2603
rect 2262 2598 2268 2599
rect 2590 2603 2596 2604
rect 2590 2599 2591 2603
rect 2595 2599 2596 2603
rect 2590 2598 2596 2599
rect 1830 2593 1836 2594
rect 1806 2592 1812 2593
rect 1806 2588 1807 2592
rect 1811 2588 1812 2592
rect 1830 2589 1831 2593
rect 1835 2589 1836 2593
rect 1830 2588 1836 2589
rect 1998 2593 2004 2594
rect 1998 2589 1999 2593
rect 2003 2589 2004 2593
rect 1998 2588 2004 2589
rect 2182 2593 2188 2594
rect 2182 2589 2183 2593
rect 2187 2589 2188 2593
rect 2182 2588 2188 2589
rect 1806 2587 1812 2588
rect 1808 2563 1810 2587
rect 1832 2563 1834 2588
rect 2000 2563 2002 2588
rect 2184 2563 2186 2588
rect 1807 2562 1811 2563
rect 1807 2557 1811 2558
rect 1831 2562 1835 2563
rect 1831 2557 1835 2558
rect 1999 2562 2003 2563
rect 1999 2557 2003 2558
rect 2183 2562 2187 2563
rect 2183 2557 2187 2558
rect 2207 2562 2211 2563
rect 2207 2557 2211 2558
rect 1798 2543 1804 2544
rect 1798 2539 1799 2543
rect 1803 2539 1804 2543
rect 1808 2541 1810 2557
rect 1798 2538 1804 2539
rect 1806 2540 1812 2541
rect 2208 2540 2210 2557
rect 1806 2536 1807 2540
rect 1811 2536 1812 2540
rect 1806 2535 1812 2536
rect 2206 2539 2212 2540
rect 2206 2535 2207 2539
rect 2211 2535 2212 2539
rect 2206 2534 2212 2535
rect 1670 2533 1676 2534
rect 1670 2529 1671 2533
rect 1675 2529 1676 2533
rect 1670 2528 1676 2529
rect 1766 2532 1772 2533
rect 1766 2528 1767 2532
rect 1771 2528 1772 2532
rect 1672 2511 1674 2528
rect 1766 2527 1772 2528
rect 2070 2531 2076 2532
rect 2070 2527 2071 2531
rect 2075 2527 2076 2531
rect 1768 2511 1770 2527
rect 2070 2526 2076 2527
rect 1806 2523 1812 2524
rect 1806 2519 1807 2523
rect 1811 2519 1812 2523
rect 1806 2518 1812 2519
rect 1671 2510 1675 2511
rect 1671 2505 1675 2506
rect 1767 2510 1771 2511
rect 1767 2505 1771 2506
rect 1672 2488 1674 2505
rect 1768 2489 1770 2505
rect 1766 2488 1772 2489
rect 1670 2487 1676 2488
rect 1670 2483 1671 2487
rect 1675 2483 1676 2487
rect 1766 2484 1767 2488
rect 1771 2484 1772 2488
rect 1766 2483 1772 2484
rect 1808 2483 1810 2518
rect 1670 2482 1676 2483
rect 1807 2482 1811 2483
rect 1662 2479 1668 2480
rect 1534 2475 1540 2476
rect 1534 2471 1535 2475
rect 1539 2471 1540 2475
rect 1534 2470 1540 2471
rect 1646 2475 1652 2476
rect 1646 2471 1647 2475
rect 1651 2471 1652 2475
rect 1662 2475 1663 2479
rect 1667 2475 1668 2479
rect 1807 2477 1811 2478
rect 2015 2482 2019 2483
rect 2015 2477 2019 2478
rect 1662 2474 1668 2475
rect 1646 2470 1652 2471
rect 1766 2471 1772 2472
rect 1462 2468 1468 2469
rect 1462 2464 1463 2468
rect 1467 2464 1468 2468
rect 1462 2463 1468 2464
rect 1382 2459 1388 2460
rect 1382 2455 1383 2459
rect 1387 2455 1388 2459
rect 1382 2454 1388 2455
rect 1464 2431 1466 2463
rect 1536 2452 1538 2470
rect 1574 2468 1580 2469
rect 1574 2464 1575 2468
rect 1579 2464 1580 2468
rect 1574 2463 1580 2464
rect 1534 2451 1540 2452
rect 1534 2447 1535 2451
rect 1539 2447 1540 2451
rect 1534 2446 1540 2447
rect 1576 2431 1578 2463
rect 1648 2452 1650 2470
rect 1670 2468 1676 2469
rect 1670 2464 1671 2468
rect 1675 2464 1676 2468
rect 1766 2467 1767 2471
rect 1771 2467 1772 2471
rect 1766 2466 1772 2467
rect 1670 2463 1676 2464
rect 1646 2451 1652 2452
rect 1646 2447 1647 2451
rect 1651 2447 1652 2451
rect 1646 2446 1652 2447
rect 1672 2431 1674 2463
rect 1768 2431 1770 2466
rect 1808 2458 1810 2477
rect 2016 2461 2018 2477
rect 2072 2476 2074 2526
rect 2206 2520 2212 2521
rect 2206 2516 2207 2520
rect 2211 2516 2212 2520
rect 2206 2515 2212 2516
rect 2208 2483 2210 2515
rect 2264 2504 2266 2598
rect 2358 2593 2364 2594
rect 2358 2589 2359 2593
rect 2363 2589 2364 2593
rect 2358 2588 2364 2589
rect 2518 2593 2524 2594
rect 2518 2589 2519 2593
rect 2523 2589 2524 2593
rect 2518 2588 2524 2589
rect 2670 2593 2676 2594
rect 2670 2589 2671 2593
rect 2675 2589 2676 2593
rect 2670 2588 2676 2589
rect 2806 2593 2812 2594
rect 2806 2589 2807 2593
rect 2811 2589 2812 2593
rect 2806 2588 2812 2589
rect 2360 2563 2362 2588
rect 2520 2563 2522 2588
rect 2672 2563 2674 2588
rect 2808 2563 2810 2588
rect 2359 2562 2363 2563
rect 2359 2557 2363 2558
rect 2519 2562 2523 2563
rect 2519 2557 2523 2558
rect 2671 2562 2675 2563
rect 2671 2557 2675 2558
rect 2799 2562 2803 2563
rect 2799 2557 2803 2558
rect 2807 2562 2811 2563
rect 2807 2557 2811 2558
rect 2800 2540 2802 2557
rect 2798 2539 2804 2540
rect 2798 2535 2799 2539
rect 2803 2535 2804 2539
rect 2798 2534 2804 2535
rect 2872 2532 2874 2614
rect 2916 2604 2918 2622
rect 2928 2613 2930 2629
rect 3034 2627 3040 2628
rect 3034 2623 3035 2627
rect 3039 2623 3040 2627
rect 3034 2622 3040 2623
rect 2926 2612 2932 2613
rect 2926 2608 2927 2612
rect 2931 2608 2932 2612
rect 2926 2607 2932 2608
rect 3036 2604 3038 2622
rect 3048 2613 3050 2629
rect 3150 2627 3156 2628
rect 3150 2623 3151 2627
rect 3155 2623 3156 2627
rect 3150 2622 3156 2623
rect 3046 2612 3052 2613
rect 3046 2608 3047 2612
rect 3051 2608 3052 2612
rect 3046 2607 3052 2608
rect 3152 2604 3154 2622
rect 3160 2613 3162 2629
rect 3272 2613 3274 2629
rect 3312 2628 3314 2662
rect 3320 2644 3322 2666
rect 3462 2663 3468 2664
rect 3366 2660 3372 2661
rect 3366 2656 3367 2660
rect 3371 2656 3372 2660
rect 3462 2659 3463 2663
rect 3467 2659 3468 2663
rect 3462 2658 3468 2659
rect 3366 2655 3372 2656
rect 3318 2643 3324 2644
rect 3318 2639 3319 2643
rect 3323 2639 3324 2643
rect 3318 2638 3324 2639
rect 3368 2635 3370 2655
rect 3430 2643 3436 2644
rect 3430 2639 3431 2643
rect 3435 2639 3436 2643
rect 3430 2638 3436 2639
rect 3367 2634 3371 2635
rect 3367 2629 3371 2630
rect 3310 2627 3316 2628
rect 3310 2623 3311 2627
rect 3315 2623 3316 2627
rect 3310 2622 3316 2623
rect 3368 2613 3370 2629
rect 3158 2612 3164 2613
rect 3158 2608 3159 2612
rect 3163 2608 3164 2612
rect 3158 2607 3164 2608
rect 3270 2612 3276 2613
rect 3270 2608 3271 2612
rect 3275 2608 3276 2612
rect 3270 2607 3276 2608
rect 3366 2612 3372 2613
rect 3366 2608 3367 2612
rect 3371 2608 3372 2612
rect 3366 2607 3372 2608
rect 3432 2604 3434 2638
rect 3464 2635 3466 2658
rect 3463 2634 3467 2635
rect 3463 2629 3467 2630
rect 3464 2610 3466 2629
rect 3462 2609 3468 2610
rect 3462 2605 3463 2609
rect 3467 2605 3468 2609
rect 3462 2604 3468 2605
rect 2914 2603 2920 2604
rect 2914 2599 2915 2603
rect 2919 2599 2920 2603
rect 2914 2598 2920 2599
rect 3034 2603 3040 2604
rect 3034 2599 3035 2603
rect 3039 2599 3040 2603
rect 3034 2598 3040 2599
rect 3150 2603 3156 2604
rect 3150 2599 3151 2603
rect 3155 2599 3156 2603
rect 3150 2598 3156 2599
rect 3430 2603 3436 2604
rect 3430 2599 3431 2603
rect 3435 2599 3436 2603
rect 3430 2598 3436 2599
rect 2926 2593 2932 2594
rect 2926 2589 2927 2593
rect 2931 2589 2932 2593
rect 2926 2588 2932 2589
rect 3046 2593 3052 2594
rect 3046 2589 3047 2593
rect 3051 2589 3052 2593
rect 3046 2588 3052 2589
rect 3158 2593 3164 2594
rect 3158 2589 3159 2593
rect 3163 2589 3164 2593
rect 3158 2588 3164 2589
rect 3270 2593 3276 2594
rect 3270 2589 3271 2593
rect 3275 2589 3276 2593
rect 3270 2588 3276 2589
rect 3366 2593 3372 2594
rect 3366 2589 3367 2593
rect 3371 2589 3372 2593
rect 3366 2588 3372 2589
rect 3462 2592 3468 2593
rect 3462 2588 3463 2592
rect 3467 2588 3468 2592
rect 2928 2563 2930 2588
rect 3048 2563 3050 2588
rect 3160 2563 3162 2588
rect 3272 2563 3274 2588
rect 3368 2563 3370 2588
rect 3462 2587 3468 2588
rect 3464 2563 3466 2587
rect 2927 2562 2931 2563
rect 2927 2557 2931 2558
rect 3047 2562 3051 2563
rect 3047 2557 3051 2558
rect 3159 2562 3163 2563
rect 3159 2557 3163 2558
rect 3271 2562 3275 2563
rect 3271 2557 3275 2558
rect 3367 2562 3371 2563
rect 3367 2557 3371 2558
rect 3463 2562 3467 2563
rect 3463 2557 3467 2558
rect 3368 2540 3370 2557
rect 3464 2541 3466 2557
rect 3462 2540 3468 2541
rect 3366 2539 3372 2540
rect 3366 2535 3367 2539
rect 3371 2535 3372 2539
rect 3462 2536 3463 2540
rect 3467 2536 3468 2540
rect 3462 2535 3468 2536
rect 3366 2534 3372 2535
rect 2870 2531 2876 2532
rect 2870 2527 2871 2531
rect 2875 2527 2876 2531
rect 2870 2526 2876 2527
rect 2878 2531 2884 2532
rect 2878 2527 2879 2531
rect 2883 2527 2884 2531
rect 2878 2526 2884 2527
rect 2798 2520 2804 2521
rect 2798 2516 2799 2520
rect 2803 2516 2804 2520
rect 2798 2515 2804 2516
rect 2262 2503 2268 2504
rect 2262 2499 2263 2503
rect 2267 2499 2268 2503
rect 2262 2498 2268 2499
rect 2800 2483 2802 2515
rect 2880 2504 2882 2526
rect 3462 2523 3468 2524
rect 3366 2520 3372 2521
rect 3366 2516 3367 2520
rect 3371 2516 3372 2520
rect 3462 2519 3463 2523
rect 3467 2519 3468 2523
rect 3462 2518 3468 2519
rect 3366 2515 3372 2516
rect 2878 2503 2884 2504
rect 2878 2499 2879 2503
rect 2883 2499 2884 2503
rect 2878 2498 2884 2499
rect 3368 2483 3370 2515
rect 3430 2503 3436 2504
rect 3430 2499 3431 2503
rect 3435 2499 3436 2503
rect 3430 2498 3436 2499
rect 2199 2482 2203 2483
rect 2199 2477 2203 2478
rect 2207 2482 2211 2483
rect 2207 2477 2211 2478
rect 2367 2482 2371 2483
rect 2367 2477 2371 2478
rect 2527 2482 2531 2483
rect 2527 2477 2531 2478
rect 2671 2482 2675 2483
rect 2671 2477 2675 2478
rect 2799 2482 2803 2483
rect 2799 2477 2803 2478
rect 2807 2482 2811 2483
rect 2807 2477 2811 2478
rect 2927 2482 2931 2483
rect 2927 2477 2931 2478
rect 3047 2482 3051 2483
rect 3047 2477 3051 2478
rect 3159 2482 3163 2483
rect 3159 2477 3163 2478
rect 3271 2482 3275 2483
rect 3271 2477 3275 2478
rect 3367 2482 3371 2483
rect 3367 2477 3371 2478
rect 2070 2475 2076 2476
rect 2070 2471 2071 2475
rect 2075 2471 2076 2475
rect 2070 2470 2076 2471
rect 2086 2475 2092 2476
rect 2086 2471 2087 2475
rect 2091 2471 2092 2475
rect 2086 2470 2092 2471
rect 2014 2460 2020 2461
rect 1806 2457 1812 2458
rect 1806 2453 1807 2457
rect 1811 2453 1812 2457
rect 2014 2456 2015 2460
rect 2019 2456 2020 2460
rect 2014 2455 2020 2456
rect 1806 2452 1812 2453
rect 2088 2452 2090 2470
rect 2200 2461 2202 2477
rect 2270 2475 2276 2476
rect 2270 2471 2271 2475
rect 2275 2471 2276 2475
rect 2270 2470 2276 2471
rect 2198 2460 2204 2461
rect 2198 2456 2199 2460
rect 2203 2456 2204 2460
rect 2198 2455 2204 2456
rect 2272 2452 2274 2470
rect 2368 2461 2370 2477
rect 2528 2461 2530 2477
rect 2630 2475 2636 2476
rect 2630 2471 2631 2475
rect 2635 2471 2636 2475
rect 2630 2470 2636 2471
rect 2646 2475 2652 2476
rect 2646 2471 2647 2475
rect 2651 2471 2652 2475
rect 2646 2470 2652 2471
rect 2366 2460 2372 2461
rect 2366 2456 2367 2460
rect 2371 2456 2372 2460
rect 2366 2455 2372 2456
rect 2526 2460 2532 2461
rect 2526 2456 2527 2460
rect 2531 2456 2532 2460
rect 2526 2455 2532 2456
rect 2086 2451 2092 2452
rect 2086 2447 2087 2451
rect 2091 2447 2092 2451
rect 2086 2446 2092 2447
rect 2270 2451 2276 2452
rect 2270 2447 2271 2451
rect 2275 2447 2276 2451
rect 2270 2446 2276 2447
rect 2430 2451 2436 2452
rect 2430 2447 2431 2451
rect 2435 2447 2436 2451
rect 2430 2446 2436 2447
rect 2014 2441 2020 2442
rect 1806 2440 1812 2441
rect 1806 2436 1807 2440
rect 1811 2436 1812 2440
rect 2014 2437 2015 2441
rect 2019 2437 2020 2441
rect 2014 2436 2020 2437
rect 2198 2441 2204 2442
rect 2198 2437 2199 2441
rect 2203 2437 2204 2441
rect 2198 2436 2204 2437
rect 2366 2441 2372 2442
rect 2366 2437 2367 2441
rect 2371 2437 2372 2441
rect 2366 2436 2372 2437
rect 1806 2435 1812 2436
rect 1351 2430 1355 2431
rect 1351 2425 1355 2426
rect 1415 2430 1419 2431
rect 1415 2425 1419 2426
rect 1463 2430 1467 2431
rect 1463 2425 1467 2426
rect 1575 2430 1579 2431
rect 1575 2425 1579 2426
rect 1591 2430 1595 2431
rect 1591 2425 1595 2426
rect 1671 2430 1675 2431
rect 1671 2425 1675 2426
rect 1767 2430 1771 2431
rect 1767 2425 1771 2426
rect 1416 2409 1418 2425
rect 1592 2409 1594 2425
rect 1598 2423 1604 2424
rect 1598 2419 1599 2423
rect 1603 2419 1604 2423
rect 1598 2418 1604 2419
rect 1414 2408 1420 2409
rect 1334 2407 1340 2408
rect 1334 2403 1335 2407
rect 1339 2403 1340 2407
rect 1414 2404 1415 2408
rect 1419 2404 1420 2408
rect 1414 2403 1420 2404
rect 1590 2408 1596 2409
rect 1590 2404 1591 2408
rect 1595 2404 1596 2408
rect 1590 2403 1596 2404
rect 1334 2402 1340 2403
rect 966 2399 972 2400
rect 966 2395 967 2399
rect 971 2395 972 2399
rect 966 2394 972 2395
rect 1030 2399 1036 2400
rect 1030 2395 1031 2399
rect 1035 2395 1036 2399
rect 1030 2394 1036 2395
rect 1318 2399 1324 2400
rect 1318 2395 1319 2399
rect 1323 2395 1324 2399
rect 1318 2394 1324 2395
rect 1062 2389 1068 2390
rect 1062 2385 1063 2389
rect 1067 2385 1068 2389
rect 1062 2384 1068 2385
rect 1238 2389 1244 2390
rect 1238 2385 1239 2389
rect 1243 2385 1244 2389
rect 1238 2384 1244 2385
rect 1414 2389 1420 2390
rect 1414 2385 1415 2389
rect 1419 2385 1420 2389
rect 1414 2384 1420 2385
rect 1590 2389 1596 2390
rect 1590 2385 1591 2389
rect 1595 2385 1596 2389
rect 1590 2384 1596 2385
rect 1064 2359 1066 2384
rect 1240 2359 1242 2384
rect 1416 2359 1418 2384
rect 1592 2359 1594 2384
rect 975 2358 979 2359
rect 975 2353 979 2354
rect 1063 2358 1067 2359
rect 1063 2353 1067 2354
rect 1103 2358 1107 2359
rect 1103 2353 1107 2354
rect 1239 2358 1243 2359
rect 1239 2353 1243 2354
rect 1375 2358 1379 2359
rect 1375 2353 1379 2354
rect 1415 2358 1419 2359
rect 1415 2353 1419 2354
rect 1511 2358 1515 2359
rect 1511 2353 1515 2354
rect 1591 2358 1595 2359
rect 1591 2353 1595 2354
rect 976 2336 978 2353
rect 1104 2336 1106 2353
rect 1240 2336 1242 2353
rect 1376 2336 1378 2353
rect 1512 2336 1514 2353
rect 974 2335 980 2336
rect 974 2331 975 2335
rect 979 2331 980 2335
rect 974 2330 980 2331
rect 1102 2335 1108 2336
rect 1102 2331 1103 2335
rect 1107 2331 1108 2335
rect 1102 2330 1108 2331
rect 1238 2335 1244 2336
rect 1238 2331 1239 2335
rect 1243 2331 1244 2335
rect 1238 2330 1244 2331
rect 1374 2335 1380 2336
rect 1374 2331 1375 2335
rect 1379 2331 1380 2335
rect 1374 2330 1380 2331
rect 1510 2335 1516 2336
rect 1510 2331 1511 2335
rect 1515 2331 1516 2335
rect 1510 2330 1516 2331
rect 1600 2328 1602 2418
rect 1768 2406 1770 2425
rect 1808 2415 1810 2435
rect 2016 2415 2018 2436
rect 2200 2415 2202 2436
rect 2368 2415 2370 2436
rect 1807 2414 1811 2415
rect 1807 2409 1811 2410
rect 1839 2414 1843 2415
rect 1839 2409 1843 2410
rect 2007 2414 2011 2415
rect 2007 2409 2011 2410
rect 2015 2414 2019 2415
rect 2015 2409 2019 2410
rect 2183 2414 2187 2415
rect 2183 2409 2187 2410
rect 2199 2414 2203 2415
rect 2199 2409 2203 2410
rect 2367 2414 2371 2415
rect 2367 2409 2371 2410
rect 1766 2405 1772 2406
rect 1766 2401 1767 2405
rect 1771 2401 1772 2405
rect 1766 2400 1772 2401
rect 1808 2393 1810 2409
rect 1806 2392 1812 2393
rect 1840 2392 1842 2409
rect 2008 2392 2010 2409
rect 2184 2392 2186 2409
rect 2368 2392 2370 2409
rect 1766 2388 1772 2389
rect 1766 2384 1767 2388
rect 1771 2384 1772 2388
rect 1806 2388 1807 2392
rect 1811 2388 1812 2392
rect 1806 2387 1812 2388
rect 1838 2391 1844 2392
rect 1838 2387 1839 2391
rect 1843 2387 1844 2391
rect 1838 2386 1844 2387
rect 2006 2391 2012 2392
rect 2006 2387 2007 2391
rect 2011 2387 2012 2391
rect 2006 2386 2012 2387
rect 2182 2391 2188 2392
rect 2182 2387 2183 2391
rect 2187 2387 2188 2391
rect 2182 2386 2188 2387
rect 2366 2391 2372 2392
rect 2366 2387 2367 2391
rect 2371 2387 2372 2391
rect 2366 2386 2372 2387
rect 1766 2383 1772 2384
rect 1918 2383 1924 2384
rect 1768 2359 1770 2383
rect 1910 2379 1916 2380
rect 1806 2375 1812 2376
rect 1806 2371 1807 2375
rect 1811 2371 1812 2375
rect 1910 2375 1911 2379
rect 1915 2375 1916 2379
rect 1918 2379 1919 2383
rect 1923 2379 1924 2383
rect 1918 2378 1924 2379
rect 2086 2383 2092 2384
rect 2086 2379 2087 2383
rect 2091 2379 2092 2383
rect 2086 2378 2092 2379
rect 2262 2383 2268 2384
rect 2262 2379 2263 2383
rect 2267 2379 2268 2383
rect 2262 2378 2268 2379
rect 1910 2374 1916 2375
rect 1806 2370 1812 2371
rect 1838 2372 1844 2373
rect 1767 2358 1771 2359
rect 1767 2353 1771 2354
rect 1768 2337 1770 2353
rect 1808 2351 1810 2370
rect 1838 2368 1839 2372
rect 1843 2368 1844 2372
rect 1838 2367 1844 2368
rect 1840 2351 1842 2367
rect 1807 2350 1811 2351
rect 1807 2345 1811 2346
rect 1839 2350 1843 2351
rect 1839 2345 1843 2346
rect 1887 2350 1891 2351
rect 1887 2345 1891 2346
rect 1766 2336 1772 2337
rect 1766 2332 1767 2336
rect 1771 2332 1772 2336
rect 1766 2331 1772 2332
rect 694 2327 700 2328
rect 670 2323 676 2324
rect 670 2319 671 2323
rect 675 2319 676 2323
rect 694 2323 695 2327
rect 699 2323 700 2327
rect 694 2322 700 2323
rect 918 2327 924 2328
rect 918 2323 919 2327
rect 923 2323 924 2327
rect 918 2322 924 2323
rect 926 2327 932 2328
rect 926 2323 927 2327
rect 931 2323 932 2327
rect 926 2322 932 2323
rect 1054 2327 1060 2328
rect 1054 2323 1055 2327
rect 1059 2323 1060 2327
rect 1598 2327 1604 2328
rect 1054 2322 1060 2323
rect 1310 2323 1316 2324
rect 670 2318 676 2319
rect 630 2307 636 2308
rect 630 2303 631 2307
rect 635 2303 636 2307
rect 630 2302 636 2303
rect 672 2300 674 2318
rect 670 2299 676 2300
rect 670 2295 671 2299
rect 675 2295 676 2299
rect 670 2294 676 2295
rect 696 2288 698 2322
rect 718 2316 724 2317
rect 718 2312 719 2316
rect 723 2312 724 2316
rect 718 2311 724 2312
rect 846 2316 852 2317
rect 846 2312 847 2316
rect 851 2312 852 2316
rect 846 2311 852 2312
rect 694 2287 700 2288
rect 720 2287 722 2311
rect 848 2287 850 2311
rect 928 2300 930 2322
rect 974 2316 980 2317
rect 974 2312 975 2316
rect 979 2312 980 2316
rect 974 2311 980 2312
rect 926 2299 932 2300
rect 926 2295 927 2299
rect 931 2295 932 2299
rect 926 2294 932 2295
rect 976 2287 978 2311
rect 1056 2300 1058 2322
rect 1310 2319 1311 2323
rect 1315 2319 1316 2323
rect 1310 2318 1316 2319
rect 1446 2323 1452 2324
rect 1446 2319 1447 2323
rect 1451 2319 1452 2323
rect 1598 2323 1599 2327
rect 1603 2323 1604 2327
rect 1808 2326 1810 2345
rect 1888 2329 1890 2345
rect 1912 2344 1914 2374
rect 1920 2356 1922 2378
rect 2006 2372 2012 2373
rect 2006 2368 2007 2372
rect 2011 2368 2012 2372
rect 2006 2367 2012 2368
rect 1918 2355 1924 2356
rect 1918 2351 1919 2355
rect 1923 2351 1924 2355
rect 2008 2351 2010 2367
rect 2088 2356 2090 2378
rect 2182 2372 2188 2373
rect 2182 2368 2183 2372
rect 2187 2368 2188 2372
rect 2182 2367 2188 2368
rect 2086 2355 2092 2356
rect 2086 2351 2087 2355
rect 2091 2351 2092 2355
rect 2184 2351 2186 2367
rect 2264 2356 2266 2378
rect 2366 2372 2372 2373
rect 2366 2368 2367 2372
rect 2371 2368 2372 2372
rect 2366 2367 2372 2368
rect 2262 2355 2268 2356
rect 2262 2351 2263 2355
rect 2267 2351 2268 2355
rect 2368 2351 2370 2367
rect 2432 2356 2434 2446
rect 2526 2441 2532 2442
rect 2526 2437 2527 2441
rect 2531 2437 2532 2441
rect 2526 2436 2532 2437
rect 2528 2415 2530 2436
rect 2527 2414 2531 2415
rect 2527 2409 2531 2410
rect 2559 2414 2563 2415
rect 2559 2409 2563 2410
rect 2560 2392 2562 2409
rect 2558 2391 2564 2392
rect 2558 2387 2559 2391
rect 2563 2387 2564 2391
rect 2558 2386 2564 2387
rect 2632 2384 2634 2470
rect 2648 2452 2650 2470
rect 2672 2461 2674 2477
rect 2742 2475 2748 2476
rect 2742 2471 2743 2475
rect 2747 2471 2748 2475
rect 2742 2470 2748 2471
rect 2670 2460 2676 2461
rect 2670 2456 2671 2460
rect 2675 2456 2676 2460
rect 2670 2455 2676 2456
rect 2744 2452 2746 2470
rect 2808 2461 2810 2477
rect 2878 2475 2884 2476
rect 2878 2471 2879 2475
rect 2883 2471 2884 2475
rect 2878 2470 2884 2471
rect 2806 2460 2812 2461
rect 2806 2456 2807 2460
rect 2811 2456 2812 2460
rect 2806 2455 2812 2456
rect 2880 2452 2882 2470
rect 2928 2461 2930 2477
rect 2998 2475 3004 2476
rect 2998 2471 2999 2475
rect 3003 2471 3004 2475
rect 2998 2470 3004 2471
rect 2926 2460 2932 2461
rect 2926 2456 2927 2460
rect 2931 2456 2932 2460
rect 2926 2455 2932 2456
rect 3000 2452 3002 2470
rect 3048 2461 3050 2477
rect 3118 2475 3124 2476
rect 3118 2471 3119 2475
rect 3123 2471 3124 2475
rect 3118 2470 3124 2471
rect 3046 2460 3052 2461
rect 3046 2456 3047 2460
rect 3051 2456 3052 2460
rect 3046 2455 3052 2456
rect 3120 2452 3122 2470
rect 3160 2461 3162 2477
rect 3230 2475 3236 2476
rect 3230 2471 3231 2475
rect 3235 2471 3236 2475
rect 3230 2470 3236 2471
rect 3158 2460 3164 2461
rect 3158 2456 3159 2460
rect 3163 2456 3164 2460
rect 3158 2455 3164 2456
rect 3232 2452 3234 2470
rect 3272 2461 3274 2477
rect 3368 2461 3370 2477
rect 3270 2460 3276 2461
rect 3270 2456 3271 2460
rect 3275 2456 3276 2460
rect 3270 2455 3276 2456
rect 3366 2460 3372 2461
rect 3366 2456 3367 2460
rect 3371 2456 3372 2460
rect 3366 2455 3372 2456
rect 3432 2452 3434 2498
rect 3464 2483 3466 2518
rect 3463 2482 3467 2483
rect 3463 2477 3467 2478
rect 3438 2475 3444 2476
rect 3438 2471 3439 2475
rect 3443 2471 3444 2475
rect 3438 2470 3444 2471
rect 2646 2451 2652 2452
rect 2646 2447 2647 2451
rect 2651 2447 2652 2451
rect 2646 2446 2652 2447
rect 2742 2451 2748 2452
rect 2742 2447 2743 2451
rect 2747 2447 2748 2451
rect 2742 2446 2748 2447
rect 2878 2451 2884 2452
rect 2878 2447 2879 2451
rect 2883 2447 2884 2451
rect 2878 2446 2884 2447
rect 2998 2451 3004 2452
rect 2998 2447 2999 2451
rect 3003 2447 3004 2451
rect 2998 2446 3004 2447
rect 3118 2451 3124 2452
rect 3118 2447 3119 2451
rect 3123 2447 3124 2451
rect 3118 2446 3124 2447
rect 3230 2451 3236 2452
rect 3230 2447 3231 2451
rect 3235 2447 3236 2451
rect 3230 2446 3236 2447
rect 3238 2451 3244 2452
rect 3238 2447 3239 2451
rect 3243 2447 3244 2451
rect 3238 2446 3244 2447
rect 3430 2451 3436 2452
rect 3430 2447 3431 2451
rect 3435 2447 3436 2451
rect 3430 2446 3436 2447
rect 2670 2441 2676 2442
rect 2670 2437 2671 2441
rect 2675 2437 2676 2441
rect 2670 2436 2676 2437
rect 2806 2441 2812 2442
rect 2806 2437 2807 2441
rect 2811 2437 2812 2441
rect 2806 2436 2812 2437
rect 2926 2441 2932 2442
rect 2926 2437 2927 2441
rect 2931 2437 2932 2441
rect 2926 2436 2932 2437
rect 3046 2441 3052 2442
rect 3046 2437 3047 2441
rect 3051 2437 3052 2441
rect 3046 2436 3052 2437
rect 3158 2441 3164 2442
rect 3158 2437 3159 2441
rect 3163 2437 3164 2441
rect 3158 2436 3164 2437
rect 2672 2415 2674 2436
rect 2808 2415 2810 2436
rect 2928 2415 2930 2436
rect 3048 2415 3050 2436
rect 3160 2415 3162 2436
rect 2671 2414 2675 2415
rect 2671 2409 2675 2410
rect 2759 2414 2763 2415
rect 2759 2409 2763 2410
rect 2807 2414 2811 2415
rect 2807 2409 2811 2410
rect 2927 2414 2931 2415
rect 2927 2409 2931 2410
rect 2967 2414 2971 2415
rect 2967 2409 2971 2410
rect 3047 2414 3051 2415
rect 3047 2409 3051 2410
rect 3159 2414 3163 2415
rect 3159 2409 3163 2410
rect 3175 2414 3179 2415
rect 3175 2409 3179 2410
rect 2760 2392 2762 2409
rect 2968 2392 2970 2409
rect 3176 2392 3178 2409
rect 2758 2391 2764 2392
rect 2758 2387 2759 2391
rect 2763 2387 2764 2391
rect 2758 2386 2764 2387
rect 2966 2391 2972 2392
rect 2966 2387 2967 2391
rect 2971 2387 2972 2391
rect 2966 2386 2972 2387
rect 3174 2391 3180 2392
rect 3174 2387 3175 2391
rect 3179 2387 3180 2391
rect 3174 2386 3180 2387
rect 2630 2383 2636 2384
rect 2630 2379 2631 2383
rect 2635 2379 2636 2383
rect 2630 2378 2636 2379
rect 2638 2383 2644 2384
rect 2638 2379 2639 2383
rect 2643 2379 2644 2383
rect 2638 2378 2644 2379
rect 2558 2372 2564 2373
rect 2558 2368 2559 2372
rect 2563 2368 2564 2372
rect 2558 2367 2564 2368
rect 2430 2355 2436 2356
rect 2430 2351 2431 2355
rect 2435 2351 2436 2355
rect 2560 2351 2562 2367
rect 2640 2356 2642 2378
rect 2758 2372 2764 2373
rect 2758 2368 2759 2372
rect 2763 2368 2764 2372
rect 2758 2367 2764 2368
rect 2966 2372 2972 2373
rect 2966 2368 2967 2372
rect 2971 2368 2972 2372
rect 2966 2367 2972 2368
rect 3174 2372 3180 2373
rect 3174 2368 3175 2372
rect 3179 2368 3180 2372
rect 3174 2367 3180 2368
rect 2638 2355 2644 2356
rect 2638 2351 2639 2355
rect 2643 2351 2644 2355
rect 2760 2351 2762 2367
rect 2968 2351 2970 2367
rect 3038 2355 3044 2356
rect 3038 2351 3039 2355
rect 3043 2351 3044 2355
rect 3176 2351 3178 2367
rect 3240 2356 3242 2446
rect 3270 2441 3276 2442
rect 3270 2437 3271 2441
rect 3275 2437 3276 2441
rect 3270 2436 3276 2437
rect 3366 2441 3372 2442
rect 3366 2437 3367 2441
rect 3371 2437 3372 2441
rect 3366 2436 3372 2437
rect 3272 2415 3274 2436
rect 3368 2415 3370 2436
rect 3271 2414 3275 2415
rect 3271 2409 3275 2410
rect 3367 2414 3371 2415
rect 3367 2409 3371 2410
rect 3368 2392 3370 2409
rect 3366 2391 3372 2392
rect 3366 2387 3367 2391
rect 3371 2387 3372 2391
rect 3366 2386 3372 2387
rect 3440 2384 3442 2470
rect 3464 2458 3466 2477
rect 3462 2457 3468 2458
rect 3462 2453 3463 2457
rect 3467 2453 3468 2457
rect 3462 2452 3468 2453
rect 3462 2440 3468 2441
rect 3462 2436 3463 2440
rect 3467 2436 3468 2440
rect 3462 2435 3468 2436
rect 3464 2415 3466 2435
rect 3463 2414 3467 2415
rect 3463 2409 3467 2410
rect 3464 2393 3466 2409
rect 3462 2392 3468 2393
rect 3462 2388 3463 2392
rect 3467 2388 3468 2392
rect 3462 2387 3468 2388
rect 3438 2383 3444 2384
rect 3246 2379 3252 2380
rect 3246 2375 3247 2379
rect 3251 2375 3252 2379
rect 3438 2379 3439 2383
rect 3443 2379 3444 2383
rect 3438 2378 3444 2379
rect 3246 2374 3252 2375
rect 3462 2375 3468 2376
rect 3238 2355 3244 2356
rect 3238 2351 3239 2355
rect 3243 2351 3244 2355
rect 1918 2350 1924 2351
rect 2007 2350 2011 2351
rect 2007 2345 2011 2346
rect 2015 2350 2019 2351
rect 2086 2350 2092 2351
rect 2151 2350 2155 2351
rect 2015 2345 2019 2346
rect 2151 2345 2155 2346
rect 2183 2350 2187 2351
rect 2262 2350 2268 2351
rect 2303 2350 2307 2351
rect 2183 2345 2187 2346
rect 2303 2345 2307 2346
rect 2367 2350 2371 2351
rect 2430 2350 2436 2351
rect 2463 2350 2467 2351
rect 2367 2345 2371 2346
rect 2463 2345 2467 2346
rect 2559 2350 2563 2351
rect 2638 2350 2644 2351
rect 2647 2350 2651 2351
rect 2559 2345 2563 2346
rect 2647 2345 2651 2346
rect 2759 2350 2763 2351
rect 2759 2345 2763 2346
rect 2839 2350 2843 2351
rect 2839 2345 2843 2346
rect 2967 2350 2971 2351
rect 3038 2350 3044 2351
rect 3047 2350 3051 2351
rect 2967 2345 2971 2346
rect 1910 2343 1916 2344
rect 1910 2339 1911 2343
rect 1915 2339 1916 2343
rect 1910 2338 1916 2339
rect 1958 2343 1964 2344
rect 1958 2339 1959 2343
rect 1963 2339 1964 2343
rect 1958 2338 1964 2339
rect 1886 2328 1892 2329
rect 1598 2322 1604 2323
rect 1806 2325 1812 2326
rect 1806 2321 1807 2325
rect 1811 2321 1812 2325
rect 1886 2324 1887 2328
rect 1891 2324 1892 2328
rect 1886 2323 1892 2324
rect 1806 2320 1812 2321
rect 1960 2320 1962 2338
rect 2016 2329 2018 2345
rect 2086 2343 2092 2344
rect 2086 2339 2087 2343
rect 2091 2339 2092 2343
rect 2086 2338 2092 2339
rect 2014 2328 2020 2329
rect 2014 2324 2015 2328
rect 2019 2324 2020 2328
rect 2014 2323 2020 2324
rect 2088 2320 2090 2338
rect 2152 2329 2154 2345
rect 2222 2343 2228 2344
rect 2222 2339 2223 2343
rect 2227 2339 2228 2343
rect 2222 2338 2228 2339
rect 2150 2328 2156 2329
rect 2150 2324 2151 2328
rect 2155 2324 2156 2328
rect 2150 2323 2156 2324
rect 2224 2320 2226 2338
rect 2304 2329 2306 2345
rect 2464 2329 2466 2345
rect 2648 2329 2650 2345
rect 2718 2343 2724 2344
rect 2718 2339 2719 2343
rect 2723 2339 2724 2343
rect 2718 2338 2724 2339
rect 2302 2328 2308 2329
rect 2302 2324 2303 2328
rect 2307 2324 2308 2328
rect 2302 2323 2308 2324
rect 2462 2328 2468 2329
rect 2462 2324 2463 2328
rect 2467 2324 2468 2328
rect 2462 2323 2468 2324
rect 2646 2328 2652 2329
rect 2646 2324 2647 2328
rect 2651 2324 2652 2328
rect 2646 2323 2652 2324
rect 2720 2320 2722 2338
rect 2840 2329 2842 2345
rect 2910 2343 2916 2344
rect 2910 2339 2911 2343
rect 2915 2339 2916 2343
rect 2910 2338 2916 2339
rect 2838 2328 2844 2329
rect 2838 2324 2839 2328
rect 2843 2324 2844 2328
rect 2838 2323 2844 2324
rect 2912 2320 2914 2338
rect 3040 2320 3042 2350
rect 3047 2345 3051 2346
rect 3175 2350 3179 2351
rect 3238 2350 3244 2351
rect 3175 2345 3179 2346
rect 3048 2329 3050 2345
rect 3248 2344 3250 2374
rect 3366 2372 3372 2373
rect 3366 2368 3367 2372
rect 3371 2368 3372 2372
rect 3462 2371 3463 2375
rect 3467 2371 3468 2375
rect 3462 2370 3468 2371
rect 3366 2367 3372 2368
rect 3368 2351 3370 2367
rect 3438 2355 3444 2356
rect 3438 2351 3439 2355
rect 3443 2351 3444 2355
rect 3464 2351 3466 2370
rect 3255 2350 3259 2351
rect 3255 2345 3259 2346
rect 3367 2350 3371 2351
rect 3438 2350 3444 2351
rect 3463 2350 3467 2351
rect 3367 2345 3371 2346
rect 3246 2343 3252 2344
rect 3246 2339 3247 2343
rect 3251 2339 3252 2343
rect 3246 2338 3252 2339
rect 3256 2329 3258 2345
rect 3046 2328 3052 2329
rect 3046 2324 3047 2328
rect 3051 2324 3052 2328
rect 3046 2323 3052 2324
rect 3254 2328 3260 2329
rect 3254 2324 3255 2328
rect 3259 2324 3260 2328
rect 3254 2323 3260 2324
rect 1446 2318 1452 2319
rect 1766 2319 1772 2320
rect 1102 2316 1108 2317
rect 1102 2312 1103 2316
rect 1107 2312 1108 2316
rect 1102 2311 1108 2312
rect 1238 2316 1244 2317
rect 1238 2312 1239 2316
rect 1243 2312 1244 2316
rect 1238 2311 1244 2312
rect 1054 2299 1060 2300
rect 1054 2295 1055 2299
rect 1059 2295 1060 2299
rect 1054 2294 1060 2295
rect 1104 2287 1106 2311
rect 1150 2299 1156 2300
rect 1150 2295 1151 2299
rect 1155 2295 1156 2299
rect 1150 2294 1156 2295
rect 111 2286 115 2287
rect 111 2281 115 2282
rect 375 2286 379 2287
rect 375 2281 379 2282
rect 479 2286 483 2287
rect 479 2281 483 2282
rect 575 2286 579 2287
rect 575 2281 579 2282
rect 599 2286 603 2287
rect 599 2281 603 2282
rect 663 2286 667 2287
rect 694 2283 695 2287
rect 699 2283 700 2287
rect 694 2282 700 2283
rect 719 2286 723 2287
rect 663 2281 667 2282
rect 719 2281 723 2282
rect 759 2286 763 2287
rect 759 2281 763 2282
rect 847 2286 851 2287
rect 847 2281 851 2282
rect 863 2286 867 2287
rect 863 2281 867 2282
rect 967 2286 971 2287
rect 967 2281 971 2282
rect 975 2286 979 2287
rect 975 2281 979 2282
rect 1079 2286 1083 2287
rect 1079 2281 1083 2282
rect 1103 2286 1107 2287
rect 1103 2281 1107 2282
rect 112 2262 114 2281
rect 576 2265 578 2281
rect 646 2279 652 2280
rect 646 2275 647 2279
rect 651 2275 652 2279
rect 646 2274 652 2275
rect 574 2264 580 2265
rect 110 2261 116 2262
rect 110 2257 111 2261
rect 115 2257 116 2261
rect 574 2260 575 2264
rect 579 2260 580 2264
rect 574 2259 580 2260
rect 110 2256 116 2257
rect 648 2256 650 2274
rect 664 2265 666 2281
rect 760 2265 762 2281
rect 854 2279 860 2280
rect 854 2275 855 2279
rect 859 2275 860 2279
rect 854 2274 860 2275
rect 662 2264 668 2265
rect 662 2260 663 2264
rect 667 2260 668 2264
rect 662 2259 668 2260
rect 758 2264 764 2265
rect 758 2260 759 2264
rect 763 2260 764 2264
rect 758 2259 764 2260
rect 646 2255 652 2256
rect 646 2251 647 2255
rect 651 2251 652 2255
rect 646 2250 652 2251
rect 734 2255 740 2256
rect 734 2251 735 2255
rect 739 2251 740 2255
rect 734 2250 740 2251
rect 574 2245 580 2246
rect 110 2244 116 2245
rect 110 2240 111 2244
rect 115 2240 116 2244
rect 574 2241 575 2245
rect 579 2241 580 2245
rect 574 2240 580 2241
rect 662 2245 668 2246
rect 662 2241 663 2245
rect 667 2241 668 2245
rect 662 2240 668 2241
rect 110 2239 116 2240
rect 112 2223 114 2239
rect 576 2223 578 2240
rect 664 2223 666 2240
rect 111 2222 115 2223
rect 111 2217 115 2218
rect 439 2222 443 2223
rect 439 2217 443 2218
rect 527 2222 531 2223
rect 527 2217 531 2218
rect 575 2222 579 2223
rect 575 2217 579 2218
rect 615 2222 619 2223
rect 615 2217 619 2218
rect 663 2222 667 2223
rect 663 2217 667 2218
rect 703 2222 707 2223
rect 703 2217 707 2218
rect 112 2201 114 2217
rect 110 2200 116 2201
rect 440 2200 442 2217
rect 528 2200 530 2217
rect 616 2200 618 2217
rect 704 2200 706 2217
rect 110 2196 111 2200
rect 115 2196 116 2200
rect 110 2195 116 2196
rect 438 2199 444 2200
rect 438 2195 439 2199
rect 443 2195 444 2199
rect 438 2194 444 2195
rect 526 2199 532 2200
rect 526 2195 527 2199
rect 531 2195 532 2199
rect 526 2194 532 2195
rect 614 2199 620 2200
rect 614 2195 615 2199
rect 619 2195 620 2199
rect 614 2194 620 2195
rect 702 2199 708 2200
rect 702 2195 703 2199
rect 707 2195 708 2199
rect 702 2194 708 2195
rect 510 2187 516 2188
rect 110 2183 116 2184
rect 110 2179 111 2183
rect 115 2179 116 2183
rect 510 2183 511 2187
rect 515 2183 516 2187
rect 510 2182 516 2183
rect 598 2187 604 2188
rect 598 2183 599 2187
rect 603 2183 604 2187
rect 598 2182 604 2183
rect 686 2187 692 2188
rect 686 2183 687 2187
rect 691 2183 692 2187
rect 686 2182 692 2183
rect 110 2178 116 2179
rect 438 2180 444 2181
rect 112 2143 114 2178
rect 438 2176 439 2180
rect 443 2176 444 2180
rect 438 2175 444 2176
rect 440 2143 442 2175
rect 512 2164 514 2182
rect 526 2180 532 2181
rect 526 2176 527 2180
rect 531 2176 532 2180
rect 526 2175 532 2176
rect 510 2163 516 2164
rect 510 2159 511 2163
rect 515 2159 516 2163
rect 510 2158 516 2159
rect 528 2143 530 2175
rect 600 2164 602 2182
rect 614 2180 620 2181
rect 614 2176 615 2180
rect 619 2176 620 2180
rect 614 2175 620 2176
rect 598 2163 604 2164
rect 598 2159 599 2163
rect 603 2159 604 2163
rect 598 2158 604 2159
rect 598 2155 604 2156
rect 598 2151 599 2155
rect 603 2151 604 2155
rect 598 2150 604 2151
rect 111 2142 115 2143
rect 111 2137 115 2138
rect 303 2142 307 2143
rect 303 2137 307 2138
rect 407 2142 411 2143
rect 407 2137 411 2138
rect 439 2142 443 2143
rect 439 2137 443 2138
rect 519 2142 523 2143
rect 519 2137 523 2138
rect 527 2142 531 2143
rect 527 2137 531 2138
rect 112 2118 114 2137
rect 304 2121 306 2137
rect 326 2135 332 2136
rect 326 2131 327 2135
rect 331 2131 332 2135
rect 326 2130 332 2131
rect 374 2135 380 2136
rect 374 2131 375 2135
rect 379 2131 380 2135
rect 374 2130 380 2131
rect 302 2120 308 2121
rect 110 2117 116 2118
rect 110 2113 111 2117
rect 115 2113 116 2117
rect 302 2116 303 2120
rect 307 2116 308 2120
rect 302 2115 308 2116
rect 110 2112 116 2113
rect 302 2101 308 2102
rect 110 2100 116 2101
rect 110 2096 111 2100
rect 115 2096 116 2100
rect 302 2097 303 2101
rect 307 2097 308 2101
rect 302 2096 308 2097
rect 110 2095 116 2096
rect 112 2079 114 2095
rect 304 2079 306 2096
rect 111 2078 115 2079
rect 111 2073 115 2074
rect 255 2078 259 2079
rect 255 2073 259 2074
rect 303 2078 307 2079
rect 303 2073 307 2074
rect 112 2057 114 2073
rect 110 2056 116 2057
rect 256 2056 258 2073
rect 110 2052 111 2056
rect 115 2052 116 2056
rect 110 2051 116 2052
rect 254 2055 260 2056
rect 254 2051 255 2055
rect 259 2051 260 2055
rect 254 2050 260 2051
rect 328 2048 330 2130
rect 376 2112 378 2130
rect 408 2121 410 2137
rect 478 2135 484 2136
rect 478 2131 479 2135
rect 483 2131 484 2135
rect 478 2130 484 2131
rect 406 2120 412 2121
rect 406 2116 407 2120
rect 411 2116 412 2120
rect 406 2115 412 2116
rect 480 2112 482 2130
rect 520 2121 522 2137
rect 590 2135 596 2136
rect 590 2131 591 2135
rect 595 2131 596 2135
rect 590 2130 596 2131
rect 518 2120 524 2121
rect 518 2116 519 2120
rect 523 2116 524 2120
rect 518 2115 524 2116
rect 592 2112 594 2130
rect 600 2112 602 2150
rect 616 2143 618 2175
rect 688 2164 690 2182
rect 702 2180 708 2181
rect 702 2176 703 2180
rect 707 2176 708 2180
rect 702 2175 708 2176
rect 686 2163 692 2164
rect 686 2159 687 2163
rect 691 2159 692 2163
rect 686 2158 692 2159
rect 704 2143 706 2175
rect 736 2172 738 2250
rect 758 2245 764 2246
rect 758 2241 759 2245
rect 763 2241 764 2245
rect 758 2240 764 2241
rect 760 2223 762 2240
rect 759 2222 763 2223
rect 759 2217 763 2218
rect 791 2222 795 2223
rect 791 2217 795 2218
rect 792 2200 794 2217
rect 790 2199 796 2200
rect 790 2195 791 2199
rect 795 2195 796 2199
rect 856 2196 858 2274
rect 864 2265 866 2281
rect 934 2279 940 2280
rect 934 2275 935 2279
rect 939 2275 940 2279
rect 934 2274 940 2275
rect 862 2264 868 2265
rect 862 2260 863 2264
rect 867 2260 868 2264
rect 862 2259 868 2260
rect 936 2256 938 2274
rect 968 2265 970 2281
rect 1038 2279 1044 2280
rect 1038 2275 1039 2279
rect 1043 2275 1044 2279
rect 1038 2274 1044 2275
rect 966 2264 972 2265
rect 966 2260 967 2264
rect 971 2260 972 2264
rect 966 2259 972 2260
rect 1040 2256 1042 2274
rect 1080 2265 1082 2281
rect 1078 2264 1084 2265
rect 1078 2260 1079 2264
rect 1083 2260 1084 2264
rect 1078 2259 1084 2260
rect 1152 2256 1154 2294
rect 1240 2287 1242 2311
rect 1312 2300 1314 2318
rect 1374 2316 1380 2317
rect 1374 2312 1375 2316
rect 1379 2312 1380 2316
rect 1374 2311 1380 2312
rect 1262 2299 1268 2300
rect 1262 2295 1263 2299
rect 1267 2295 1268 2299
rect 1262 2294 1268 2295
rect 1310 2299 1316 2300
rect 1310 2295 1311 2299
rect 1315 2295 1316 2299
rect 1310 2294 1316 2295
rect 1191 2286 1195 2287
rect 1191 2281 1195 2282
rect 1239 2286 1243 2287
rect 1239 2281 1243 2282
rect 1192 2265 1194 2281
rect 1190 2264 1196 2265
rect 1190 2260 1191 2264
rect 1195 2260 1196 2264
rect 1190 2259 1196 2260
rect 1264 2256 1266 2294
rect 1376 2287 1378 2311
rect 1448 2300 1450 2318
rect 1510 2316 1516 2317
rect 1510 2312 1511 2316
rect 1515 2312 1516 2316
rect 1766 2315 1767 2319
rect 1771 2315 1772 2319
rect 1766 2314 1772 2315
rect 1958 2319 1964 2320
rect 1958 2315 1959 2319
rect 1963 2315 1964 2319
rect 1958 2314 1964 2315
rect 2086 2319 2092 2320
rect 2086 2315 2087 2319
rect 2091 2315 2092 2319
rect 2086 2314 2092 2315
rect 2222 2319 2228 2320
rect 2222 2315 2223 2319
rect 2227 2315 2228 2319
rect 2222 2314 2228 2315
rect 2230 2319 2236 2320
rect 2230 2315 2231 2319
rect 2235 2315 2236 2319
rect 2230 2314 2236 2315
rect 2718 2319 2724 2320
rect 2718 2315 2719 2319
rect 2723 2315 2724 2319
rect 2718 2314 2724 2315
rect 2910 2319 2916 2320
rect 2910 2315 2911 2319
rect 2915 2315 2916 2319
rect 2910 2314 2916 2315
rect 3038 2319 3044 2320
rect 3038 2315 3039 2319
rect 3043 2315 3044 2319
rect 3038 2314 3044 2315
rect 3318 2319 3324 2320
rect 3318 2315 3319 2319
rect 3323 2315 3324 2319
rect 3318 2314 3324 2315
rect 1510 2311 1516 2312
rect 1446 2299 1452 2300
rect 1446 2295 1447 2299
rect 1451 2295 1452 2299
rect 1446 2294 1452 2295
rect 1512 2287 1514 2311
rect 1768 2287 1770 2314
rect 1886 2309 1892 2310
rect 1806 2308 1812 2309
rect 1806 2304 1807 2308
rect 1811 2304 1812 2308
rect 1886 2305 1887 2309
rect 1891 2305 1892 2309
rect 1886 2304 1892 2305
rect 2014 2309 2020 2310
rect 2014 2305 2015 2309
rect 2019 2305 2020 2309
rect 2014 2304 2020 2305
rect 2150 2309 2156 2310
rect 2150 2305 2151 2309
rect 2155 2305 2156 2309
rect 2150 2304 2156 2305
rect 1806 2303 1812 2304
rect 1303 2286 1307 2287
rect 1303 2281 1307 2282
rect 1375 2286 1379 2287
rect 1375 2281 1379 2282
rect 1415 2286 1419 2287
rect 1415 2281 1419 2282
rect 1511 2286 1515 2287
rect 1511 2281 1515 2282
rect 1767 2286 1771 2287
rect 1808 2283 1810 2303
rect 1888 2283 1890 2304
rect 2016 2283 2018 2304
rect 2152 2283 2154 2304
rect 1767 2281 1771 2282
rect 1807 2282 1811 2283
rect 1304 2265 1306 2281
rect 1416 2265 1418 2281
rect 1302 2264 1308 2265
rect 1302 2260 1303 2264
rect 1307 2260 1308 2264
rect 1302 2259 1308 2260
rect 1414 2264 1420 2265
rect 1414 2260 1415 2264
rect 1419 2260 1420 2264
rect 1768 2262 1770 2281
rect 1807 2277 1811 2278
rect 1887 2282 1891 2283
rect 1887 2277 1891 2278
rect 2015 2282 2019 2283
rect 2015 2277 2019 2278
rect 2039 2282 2043 2283
rect 2039 2277 2043 2278
rect 2135 2282 2139 2283
rect 2135 2277 2139 2278
rect 2151 2282 2155 2283
rect 2151 2277 2155 2278
rect 1414 2259 1420 2260
rect 1766 2261 1772 2262
rect 1808 2261 1810 2277
rect 1766 2257 1767 2261
rect 1771 2257 1772 2261
rect 1766 2256 1772 2257
rect 1806 2260 1812 2261
rect 2040 2260 2042 2277
rect 2136 2260 2138 2277
rect 1806 2256 1807 2260
rect 1811 2256 1812 2260
rect 934 2255 940 2256
rect 934 2251 935 2255
rect 939 2251 940 2255
rect 934 2250 940 2251
rect 1038 2255 1044 2256
rect 1038 2251 1039 2255
rect 1043 2251 1044 2255
rect 1038 2250 1044 2251
rect 1150 2255 1156 2256
rect 1150 2251 1151 2255
rect 1155 2251 1156 2255
rect 1150 2250 1156 2251
rect 1262 2255 1268 2256
rect 1806 2255 1812 2256
rect 2038 2259 2044 2260
rect 2038 2255 2039 2259
rect 2043 2255 2044 2259
rect 1262 2251 1263 2255
rect 1267 2251 1268 2255
rect 2038 2254 2044 2255
rect 2134 2259 2140 2260
rect 2134 2255 2135 2259
rect 2139 2255 2140 2259
rect 2134 2254 2140 2255
rect 1262 2250 1268 2251
rect 2110 2247 2116 2248
rect 862 2245 868 2246
rect 862 2241 863 2245
rect 867 2241 868 2245
rect 862 2240 868 2241
rect 966 2245 972 2246
rect 966 2241 967 2245
rect 971 2241 972 2245
rect 966 2240 972 2241
rect 1078 2245 1084 2246
rect 1078 2241 1079 2245
rect 1083 2241 1084 2245
rect 1078 2240 1084 2241
rect 1190 2245 1196 2246
rect 1190 2241 1191 2245
rect 1195 2241 1196 2245
rect 1190 2240 1196 2241
rect 1302 2245 1308 2246
rect 1302 2241 1303 2245
rect 1307 2241 1308 2245
rect 1302 2240 1308 2241
rect 1414 2245 1420 2246
rect 1414 2241 1415 2245
rect 1419 2241 1420 2245
rect 1414 2240 1420 2241
rect 1766 2244 1772 2245
rect 1766 2240 1767 2244
rect 1771 2240 1772 2244
rect 864 2223 866 2240
rect 968 2223 970 2240
rect 1080 2223 1082 2240
rect 1192 2223 1194 2240
rect 1304 2223 1306 2240
rect 1416 2223 1418 2240
rect 1766 2239 1772 2240
rect 1806 2243 1812 2244
rect 1806 2239 1807 2243
rect 1811 2239 1812 2243
rect 2110 2243 2111 2247
rect 2115 2243 2116 2247
rect 2110 2242 2116 2243
rect 2206 2247 2212 2248
rect 2206 2243 2207 2247
rect 2211 2243 2212 2247
rect 2206 2242 2212 2243
rect 1768 2223 1770 2239
rect 1806 2238 1812 2239
rect 2038 2240 2044 2241
rect 863 2222 867 2223
rect 863 2217 867 2218
rect 879 2222 883 2223
rect 879 2217 883 2218
rect 967 2222 971 2223
rect 967 2217 971 2218
rect 1055 2222 1059 2223
rect 1055 2217 1059 2218
rect 1079 2222 1083 2223
rect 1079 2217 1083 2218
rect 1143 2222 1147 2223
rect 1143 2217 1147 2218
rect 1191 2222 1195 2223
rect 1191 2217 1195 2218
rect 1231 2222 1235 2223
rect 1231 2217 1235 2218
rect 1303 2222 1307 2223
rect 1303 2217 1307 2218
rect 1319 2222 1323 2223
rect 1319 2217 1323 2218
rect 1415 2222 1419 2223
rect 1415 2217 1419 2218
rect 1767 2222 1771 2223
rect 1767 2217 1771 2218
rect 880 2200 882 2217
rect 968 2200 970 2217
rect 1056 2200 1058 2217
rect 1144 2200 1146 2217
rect 1232 2200 1234 2217
rect 1320 2200 1322 2217
rect 1768 2201 1770 2217
rect 1808 2207 1810 2238
rect 2038 2236 2039 2240
rect 2043 2236 2044 2240
rect 2038 2235 2044 2236
rect 2040 2207 2042 2235
rect 2112 2224 2114 2242
rect 2134 2240 2140 2241
rect 2134 2236 2135 2240
rect 2139 2236 2140 2240
rect 2134 2235 2140 2236
rect 2110 2223 2116 2224
rect 2110 2219 2111 2223
rect 2115 2219 2116 2223
rect 2110 2218 2116 2219
rect 2136 2207 2138 2235
rect 2208 2224 2210 2242
rect 2232 2232 2234 2314
rect 2302 2309 2308 2310
rect 2302 2305 2303 2309
rect 2307 2305 2308 2309
rect 2302 2304 2308 2305
rect 2462 2309 2468 2310
rect 2462 2305 2463 2309
rect 2467 2305 2468 2309
rect 2462 2304 2468 2305
rect 2646 2309 2652 2310
rect 2646 2305 2647 2309
rect 2651 2305 2652 2309
rect 2646 2304 2652 2305
rect 2838 2309 2844 2310
rect 2838 2305 2839 2309
rect 2843 2305 2844 2309
rect 2838 2304 2844 2305
rect 3046 2309 3052 2310
rect 3046 2305 3047 2309
rect 3051 2305 3052 2309
rect 3046 2304 3052 2305
rect 3254 2309 3260 2310
rect 3254 2305 3255 2309
rect 3259 2305 3260 2309
rect 3254 2304 3260 2305
rect 2304 2283 2306 2304
rect 2464 2283 2466 2304
rect 2648 2283 2650 2304
rect 2840 2283 2842 2304
rect 3048 2283 3050 2304
rect 3256 2283 3258 2304
rect 2239 2282 2243 2283
rect 2239 2277 2243 2278
rect 2303 2282 2307 2283
rect 2303 2277 2307 2278
rect 2343 2282 2347 2283
rect 2343 2277 2347 2278
rect 2463 2282 2467 2283
rect 2463 2277 2467 2278
rect 2591 2282 2595 2283
rect 2591 2277 2595 2278
rect 2647 2282 2651 2283
rect 2647 2277 2651 2278
rect 2735 2282 2739 2283
rect 2735 2277 2739 2278
rect 2839 2282 2843 2283
rect 2839 2277 2843 2278
rect 2887 2282 2891 2283
rect 2887 2277 2891 2278
rect 3047 2282 3051 2283
rect 3047 2277 3051 2278
rect 3215 2282 3219 2283
rect 3215 2277 3219 2278
rect 3255 2282 3259 2283
rect 3255 2277 3259 2278
rect 2240 2260 2242 2277
rect 2344 2260 2346 2277
rect 2464 2260 2466 2277
rect 2592 2260 2594 2277
rect 2736 2260 2738 2277
rect 2888 2260 2890 2277
rect 3048 2260 3050 2277
rect 3216 2260 3218 2277
rect 2238 2259 2244 2260
rect 2238 2255 2239 2259
rect 2243 2255 2244 2259
rect 2238 2254 2244 2255
rect 2342 2259 2348 2260
rect 2342 2255 2343 2259
rect 2347 2255 2348 2259
rect 2342 2254 2348 2255
rect 2462 2259 2468 2260
rect 2462 2255 2463 2259
rect 2467 2255 2468 2259
rect 2462 2254 2468 2255
rect 2590 2259 2596 2260
rect 2590 2255 2591 2259
rect 2595 2255 2596 2259
rect 2590 2254 2596 2255
rect 2734 2259 2740 2260
rect 2734 2255 2735 2259
rect 2739 2255 2740 2259
rect 2734 2254 2740 2255
rect 2886 2259 2892 2260
rect 2886 2255 2887 2259
rect 2891 2255 2892 2259
rect 2886 2254 2892 2255
rect 3046 2259 3052 2260
rect 3046 2255 3047 2259
rect 3051 2255 3052 2259
rect 3046 2254 3052 2255
rect 3214 2259 3220 2260
rect 3214 2255 3215 2259
rect 3219 2255 3220 2259
rect 3214 2254 3220 2255
rect 2430 2251 2436 2252
rect 2310 2247 2316 2248
rect 2310 2243 2311 2247
rect 2315 2243 2316 2247
rect 2310 2242 2316 2243
rect 2414 2247 2420 2248
rect 2414 2243 2415 2247
rect 2419 2243 2420 2247
rect 2430 2247 2431 2251
rect 2435 2247 2436 2251
rect 2430 2246 2436 2247
rect 2670 2251 2676 2252
rect 2670 2247 2671 2251
rect 2675 2247 2676 2251
rect 2670 2246 2676 2247
rect 2814 2251 2820 2252
rect 2814 2247 2815 2251
rect 2819 2247 2820 2251
rect 2814 2246 2820 2247
rect 2966 2251 2972 2252
rect 2966 2247 2967 2251
rect 2971 2247 2972 2251
rect 2966 2246 2972 2247
rect 2414 2242 2420 2243
rect 2238 2240 2244 2241
rect 2238 2236 2239 2240
rect 2243 2236 2244 2240
rect 2238 2235 2244 2236
rect 2230 2231 2236 2232
rect 2230 2227 2231 2231
rect 2235 2227 2236 2231
rect 2230 2226 2236 2227
rect 2206 2223 2212 2224
rect 2206 2219 2207 2223
rect 2211 2219 2212 2223
rect 2206 2218 2212 2219
rect 2240 2207 2242 2235
rect 2312 2224 2314 2242
rect 2342 2240 2348 2241
rect 2342 2236 2343 2240
rect 2347 2236 2348 2240
rect 2342 2235 2348 2236
rect 2310 2223 2316 2224
rect 2310 2219 2311 2223
rect 2315 2219 2316 2223
rect 2310 2218 2316 2219
rect 2344 2207 2346 2235
rect 2416 2224 2418 2242
rect 2414 2223 2420 2224
rect 2414 2219 2415 2223
rect 2419 2219 2420 2223
rect 2414 2218 2420 2219
rect 2432 2208 2434 2246
rect 2462 2240 2468 2241
rect 2462 2236 2463 2240
rect 2467 2236 2468 2240
rect 2462 2235 2468 2236
rect 2590 2240 2596 2241
rect 2590 2236 2591 2240
rect 2595 2236 2596 2240
rect 2590 2235 2596 2236
rect 2430 2207 2436 2208
rect 2464 2207 2466 2235
rect 2592 2207 2594 2235
rect 2672 2224 2674 2246
rect 2734 2240 2740 2241
rect 2734 2236 2735 2240
rect 2739 2236 2740 2240
rect 2734 2235 2740 2236
rect 2670 2223 2676 2224
rect 2670 2219 2671 2223
rect 2675 2219 2676 2223
rect 2670 2218 2676 2219
rect 2736 2207 2738 2235
rect 2816 2224 2818 2246
rect 2886 2240 2892 2241
rect 2886 2236 2887 2240
rect 2891 2236 2892 2240
rect 2886 2235 2892 2236
rect 2814 2223 2820 2224
rect 2814 2219 2815 2223
rect 2819 2219 2820 2223
rect 2814 2218 2820 2219
rect 2888 2207 2890 2235
rect 2968 2224 2970 2246
rect 3046 2240 3052 2241
rect 3046 2236 3047 2240
rect 3051 2236 3052 2240
rect 3046 2235 3052 2236
rect 3214 2240 3220 2241
rect 3214 2236 3215 2240
rect 3219 2236 3220 2240
rect 3214 2235 3220 2236
rect 2966 2223 2972 2224
rect 2966 2219 2967 2223
rect 2971 2219 2972 2223
rect 2966 2218 2972 2219
rect 3038 2223 3044 2224
rect 3038 2219 3039 2223
rect 3043 2219 3044 2223
rect 3038 2218 3044 2219
rect 1807 2206 1811 2207
rect 1807 2201 1811 2202
rect 2039 2206 2043 2207
rect 2039 2201 2043 2202
rect 2135 2206 2139 2207
rect 2135 2201 2139 2202
rect 2183 2206 2187 2207
rect 2183 2201 2187 2202
rect 2239 2206 2243 2207
rect 2239 2201 2243 2202
rect 2279 2206 2283 2207
rect 2279 2201 2283 2202
rect 2343 2206 2347 2207
rect 2343 2201 2347 2202
rect 2383 2206 2387 2207
rect 2430 2203 2431 2207
rect 2435 2203 2436 2207
rect 2430 2202 2436 2203
rect 2463 2206 2467 2207
rect 2383 2201 2387 2202
rect 2463 2201 2467 2202
rect 2495 2206 2499 2207
rect 2495 2201 2499 2202
rect 2591 2206 2595 2207
rect 2591 2201 2595 2202
rect 2607 2206 2611 2207
rect 2607 2201 2611 2202
rect 2719 2206 2723 2207
rect 2719 2201 2723 2202
rect 2735 2206 2739 2207
rect 2735 2201 2739 2202
rect 2839 2206 2843 2207
rect 2839 2201 2843 2202
rect 2887 2206 2891 2207
rect 2887 2201 2891 2202
rect 2967 2206 2971 2207
rect 2967 2201 2971 2202
rect 1766 2200 1772 2201
rect 878 2199 884 2200
rect 790 2194 796 2195
rect 854 2195 860 2196
rect 854 2191 855 2195
rect 859 2191 860 2195
rect 878 2195 879 2199
rect 883 2195 884 2199
rect 878 2194 884 2195
rect 966 2199 972 2200
rect 966 2195 967 2199
rect 971 2195 972 2199
rect 966 2194 972 2195
rect 1054 2199 1060 2200
rect 1054 2195 1055 2199
rect 1059 2195 1060 2199
rect 1054 2194 1060 2195
rect 1142 2199 1148 2200
rect 1142 2195 1143 2199
rect 1147 2195 1148 2199
rect 1142 2194 1148 2195
rect 1230 2199 1236 2200
rect 1230 2195 1231 2199
rect 1235 2195 1236 2199
rect 1230 2194 1236 2195
rect 1318 2199 1324 2200
rect 1318 2195 1319 2199
rect 1323 2195 1324 2199
rect 1766 2196 1767 2200
rect 1771 2196 1772 2200
rect 1766 2195 1772 2196
rect 1318 2194 1324 2195
rect 854 2190 860 2191
rect 774 2187 780 2188
rect 774 2183 775 2187
rect 779 2183 780 2187
rect 774 2182 780 2183
rect 950 2187 956 2188
rect 950 2183 951 2187
rect 955 2183 956 2187
rect 950 2182 956 2183
rect 1038 2187 1044 2188
rect 1038 2183 1039 2187
rect 1043 2183 1044 2187
rect 1038 2182 1044 2183
rect 1126 2187 1132 2188
rect 1126 2183 1127 2187
rect 1131 2183 1132 2187
rect 1126 2182 1132 2183
rect 1214 2187 1220 2188
rect 1214 2183 1215 2187
rect 1219 2183 1220 2187
rect 1214 2182 1220 2183
rect 1302 2187 1308 2188
rect 1302 2183 1303 2187
rect 1307 2183 1308 2187
rect 1302 2182 1308 2183
rect 1766 2183 1772 2184
rect 734 2171 740 2172
rect 734 2167 735 2171
rect 739 2167 740 2171
rect 734 2166 740 2167
rect 776 2164 778 2182
rect 790 2180 796 2181
rect 790 2176 791 2180
rect 795 2176 796 2180
rect 790 2175 796 2176
rect 878 2180 884 2181
rect 878 2176 879 2180
rect 883 2176 884 2180
rect 878 2175 884 2176
rect 774 2163 780 2164
rect 774 2159 775 2163
rect 779 2159 780 2163
rect 774 2158 780 2159
rect 792 2143 794 2175
rect 880 2143 882 2175
rect 952 2164 954 2182
rect 966 2180 972 2181
rect 966 2176 967 2180
rect 971 2176 972 2180
rect 966 2175 972 2176
rect 950 2163 956 2164
rect 950 2159 951 2163
rect 955 2159 956 2163
rect 950 2158 956 2159
rect 968 2143 970 2175
rect 1040 2164 1042 2182
rect 1054 2180 1060 2181
rect 1054 2176 1055 2180
rect 1059 2176 1060 2180
rect 1054 2175 1060 2176
rect 1038 2163 1044 2164
rect 1038 2159 1039 2163
rect 1043 2159 1044 2163
rect 1038 2158 1044 2159
rect 1056 2143 1058 2175
rect 1128 2164 1130 2182
rect 1142 2180 1148 2181
rect 1142 2176 1143 2180
rect 1147 2176 1148 2180
rect 1142 2175 1148 2176
rect 1126 2163 1132 2164
rect 1126 2159 1127 2163
rect 1131 2159 1132 2163
rect 1126 2158 1132 2159
rect 1144 2143 1146 2175
rect 1216 2164 1218 2182
rect 1230 2180 1236 2181
rect 1230 2176 1231 2180
rect 1235 2176 1236 2180
rect 1230 2175 1236 2176
rect 1214 2163 1220 2164
rect 1214 2159 1215 2163
rect 1219 2159 1220 2163
rect 1214 2158 1220 2159
rect 1232 2143 1234 2175
rect 1304 2164 1306 2182
rect 1318 2180 1324 2181
rect 1318 2176 1319 2180
rect 1323 2176 1324 2180
rect 1766 2179 1767 2183
rect 1771 2179 1772 2183
rect 1808 2182 1810 2201
rect 2184 2185 2186 2201
rect 2254 2199 2260 2200
rect 2254 2195 2255 2199
rect 2259 2195 2260 2199
rect 2254 2194 2260 2195
rect 2182 2184 2188 2185
rect 1766 2178 1772 2179
rect 1806 2181 1812 2182
rect 1318 2175 1324 2176
rect 1302 2163 1308 2164
rect 1302 2159 1303 2163
rect 1307 2159 1308 2163
rect 1302 2158 1308 2159
rect 1320 2143 1322 2175
rect 1768 2143 1770 2178
rect 1806 2177 1807 2181
rect 1811 2177 1812 2181
rect 2182 2180 2183 2184
rect 2187 2180 2188 2184
rect 2182 2179 2188 2180
rect 1806 2176 1812 2177
rect 2256 2176 2258 2194
rect 2280 2185 2282 2201
rect 2350 2199 2356 2200
rect 2350 2195 2351 2199
rect 2355 2195 2356 2199
rect 2350 2194 2356 2195
rect 2278 2184 2284 2185
rect 2278 2180 2279 2184
rect 2283 2180 2284 2184
rect 2278 2179 2284 2180
rect 2352 2176 2354 2194
rect 2384 2185 2386 2201
rect 2454 2199 2460 2200
rect 2454 2195 2455 2199
rect 2459 2195 2460 2199
rect 2454 2194 2460 2195
rect 2382 2184 2388 2185
rect 2382 2180 2383 2184
rect 2387 2180 2388 2184
rect 2382 2179 2388 2180
rect 2456 2176 2458 2194
rect 2496 2185 2498 2201
rect 2566 2199 2572 2200
rect 2566 2195 2567 2199
rect 2571 2195 2572 2199
rect 2566 2194 2572 2195
rect 2494 2184 2500 2185
rect 2494 2180 2495 2184
rect 2499 2180 2500 2184
rect 2494 2179 2500 2180
rect 2568 2176 2570 2194
rect 2608 2185 2610 2201
rect 2720 2185 2722 2201
rect 2790 2199 2796 2200
rect 2790 2195 2791 2199
rect 2795 2195 2796 2199
rect 2790 2194 2796 2195
rect 2606 2184 2612 2185
rect 2606 2180 2607 2184
rect 2611 2180 2612 2184
rect 2606 2179 2612 2180
rect 2718 2184 2724 2185
rect 2718 2180 2719 2184
rect 2723 2180 2724 2184
rect 2718 2179 2724 2180
rect 2792 2176 2794 2194
rect 2840 2185 2842 2201
rect 2910 2199 2916 2200
rect 2910 2195 2911 2199
rect 2915 2195 2916 2199
rect 2910 2194 2916 2195
rect 2838 2184 2844 2185
rect 2838 2180 2839 2184
rect 2843 2180 2844 2184
rect 2838 2179 2844 2180
rect 2912 2176 2914 2194
rect 2968 2185 2970 2201
rect 2966 2184 2972 2185
rect 2966 2180 2967 2184
rect 2971 2180 2972 2184
rect 2966 2179 2972 2180
rect 3040 2176 3042 2218
rect 3048 2207 3050 2235
rect 3216 2207 3218 2235
rect 3320 2224 3322 2314
rect 3367 2282 3371 2283
rect 3367 2277 3371 2278
rect 3368 2260 3370 2277
rect 3366 2259 3372 2260
rect 3366 2255 3367 2259
rect 3371 2255 3372 2259
rect 3366 2254 3372 2255
rect 3440 2252 3442 2350
rect 3463 2345 3467 2346
rect 3464 2326 3466 2345
rect 3462 2325 3468 2326
rect 3462 2321 3463 2325
rect 3467 2321 3468 2325
rect 3462 2320 3468 2321
rect 3462 2308 3468 2309
rect 3462 2304 3463 2308
rect 3467 2304 3468 2308
rect 3462 2303 3468 2304
rect 3464 2283 3466 2303
rect 3463 2282 3467 2283
rect 3463 2277 3467 2278
rect 3464 2261 3466 2277
rect 3462 2260 3468 2261
rect 3462 2256 3463 2260
rect 3467 2256 3468 2260
rect 3462 2255 3468 2256
rect 3438 2251 3444 2252
rect 3338 2247 3344 2248
rect 3338 2243 3339 2247
rect 3343 2243 3344 2247
rect 3438 2247 3439 2251
rect 3443 2247 3444 2251
rect 3438 2246 3444 2247
rect 3338 2242 3344 2243
rect 3462 2243 3468 2244
rect 3318 2223 3324 2224
rect 3318 2219 3319 2223
rect 3323 2219 3324 2223
rect 3318 2218 3324 2219
rect 3047 2206 3051 2207
rect 3047 2201 3051 2202
rect 3103 2206 3107 2207
rect 3103 2201 3107 2202
rect 3215 2206 3219 2207
rect 3215 2201 3219 2202
rect 3247 2206 3251 2207
rect 3247 2201 3251 2202
rect 3104 2185 3106 2201
rect 3114 2199 3120 2200
rect 3114 2195 3115 2199
rect 3119 2195 3120 2199
rect 3114 2194 3120 2195
rect 3174 2199 3180 2200
rect 3174 2195 3175 2199
rect 3179 2195 3180 2199
rect 3174 2194 3180 2195
rect 3102 2184 3108 2185
rect 3102 2180 3103 2184
rect 3107 2180 3108 2184
rect 3102 2179 3108 2180
rect 2254 2175 2260 2176
rect 2254 2171 2255 2175
rect 2259 2171 2260 2175
rect 2254 2170 2260 2171
rect 2350 2175 2356 2176
rect 2350 2171 2351 2175
rect 2355 2171 2356 2175
rect 2350 2170 2356 2171
rect 2454 2175 2460 2176
rect 2454 2171 2455 2175
rect 2459 2171 2460 2175
rect 2454 2170 2460 2171
rect 2566 2175 2572 2176
rect 2566 2171 2567 2175
rect 2571 2171 2572 2175
rect 2566 2170 2572 2171
rect 2678 2175 2684 2176
rect 2678 2171 2679 2175
rect 2683 2171 2684 2175
rect 2678 2170 2684 2171
rect 2790 2175 2796 2176
rect 2790 2171 2791 2175
rect 2795 2171 2796 2175
rect 2790 2170 2796 2171
rect 2910 2175 2916 2176
rect 2910 2171 2911 2175
rect 2915 2171 2916 2175
rect 2910 2170 2916 2171
rect 3038 2175 3044 2176
rect 3038 2171 3039 2175
rect 3043 2171 3044 2175
rect 3038 2170 3044 2171
rect 2182 2165 2188 2166
rect 1806 2164 1812 2165
rect 1806 2160 1807 2164
rect 1811 2160 1812 2164
rect 2182 2161 2183 2165
rect 2187 2161 2188 2165
rect 2182 2160 2188 2161
rect 2278 2165 2284 2166
rect 2278 2161 2279 2165
rect 2283 2161 2284 2165
rect 2278 2160 2284 2161
rect 2382 2165 2388 2166
rect 2382 2161 2383 2165
rect 2387 2161 2388 2165
rect 2382 2160 2388 2161
rect 2494 2165 2500 2166
rect 2494 2161 2495 2165
rect 2499 2161 2500 2165
rect 2494 2160 2500 2161
rect 2606 2165 2612 2166
rect 2606 2161 2607 2165
rect 2611 2161 2612 2165
rect 2606 2160 2612 2161
rect 1806 2159 1812 2160
rect 615 2142 619 2143
rect 615 2137 619 2138
rect 631 2142 635 2143
rect 631 2137 635 2138
rect 703 2142 707 2143
rect 703 2137 707 2138
rect 743 2142 747 2143
rect 743 2137 747 2138
rect 791 2142 795 2143
rect 791 2137 795 2138
rect 863 2142 867 2143
rect 863 2137 867 2138
rect 879 2142 883 2143
rect 879 2137 883 2138
rect 967 2142 971 2143
rect 967 2137 971 2138
rect 983 2142 987 2143
rect 983 2137 987 2138
rect 1055 2142 1059 2143
rect 1055 2137 1059 2138
rect 1143 2142 1147 2143
rect 1143 2137 1147 2138
rect 1231 2142 1235 2143
rect 1231 2137 1235 2138
rect 1319 2142 1323 2143
rect 1319 2137 1323 2138
rect 1767 2142 1771 2143
rect 1767 2137 1771 2138
rect 632 2121 634 2137
rect 744 2121 746 2137
rect 822 2135 828 2136
rect 822 2131 823 2135
rect 827 2131 828 2135
rect 822 2130 828 2131
rect 630 2120 636 2121
rect 630 2116 631 2120
rect 635 2116 636 2120
rect 630 2115 636 2116
rect 742 2120 748 2121
rect 742 2116 743 2120
rect 747 2116 748 2120
rect 742 2115 748 2116
rect 824 2112 826 2130
rect 864 2121 866 2137
rect 984 2121 986 2137
rect 1006 2135 1012 2136
rect 1006 2131 1007 2135
rect 1011 2131 1012 2135
rect 1006 2130 1012 2131
rect 862 2120 868 2121
rect 862 2116 863 2120
rect 867 2116 868 2120
rect 862 2115 868 2116
rect 982 2120 988 2121
rect 982 2116 983 2120
rect 987 2116 988 2120
rect 982 2115 988 2116
rect 374 2111 380 2112
rect 374 2107 375 2111
rect 379 2107 380 2111
rect 374 2106 380 2107
rect 478 2111 484 2112
rect 478 2107 479 2111
rect 483 2107 484 2111
rect 478 2106 484 2107
rect 590 2111 596 2112
rect 590 2107 591 2111
rect 595 2107 596 2111
rect 590 2106 596 2107
rect 598 2111 604 2112
rect 598 2107 599 2111
rect 603 2107 604 2111
rect 598 2106 604 2107
rect 718 2111 724 2112
rect 718 2107 719 2111
rect 723 2107 724 2111
rect 718 2106 724 2107
rect 822 2111 828 2112
rect 822 2107 823 2111
rect 827 2107 828 2111
rect 822 2106 828 2107
rect 406 2101 412 2102
rect 406 2097 407 2101
rect 411 2097 412 2101
rect 406 2096 412 2097
rect 518 2101 524 2102
rect 518 2097 519 2101
rect 523 2097 524 2101
rect 518 2096 524 2097
rect 630 2101 636 2102
rect 630 2097 631 2101
rect 635 2097 636 2101
rect 630 2096 636 2097
rect 408 2079 410 2096
rect 520 2079 522 2096
rect 632 2079 634 2096
rect 375 2078 379 2079
rect 375 2073 379 2074
rect 407 2078 411 2079
rect 407 2073 411 2074
rect 495 2078 499 2079
rect 495 2073 499 2074
rect 519 2078 523 2079
rect 519 2073 523 2074
rect 615 2078 619 2079
rect 615 2073 619 2074
rect 631 2078 635 2079
rect 631 2073 635 2074
rect 376 2056 378 2073
rect 496 2056 498 2073
rect 616 2056 618 2073
rect 374 2055 380 2056
rect 374 2051 375 2055
rect 379 2051 380 2055
rect 374 2050 380 2051
rect 494 2055 500 2056
rect 494 2051 495 2055
rect 499 2051 500 2055
rect 494 2050 500 2051
rect 614 2055 620 2056
rect 614 2051 615 2055
rect 619 2051 620 2055
rect 614 2050 620 2051
rect 326 2047 332 2048
rect 326 2043 327 2047
rect 331 2043 332 2047
rect 326 2042 332 2043
rect 334 2047 340 2048
rect 334 2043 335 2047
rect 339 2043 340 2047
rect 334 2042 340 2043
rect 454 2047 460 2048
rect 454 2043 455 2047
rect 459 2043 460 2047
rect 454 2042 460 2043
rect 686 2043 692 2044
rect 110 2039 116 2040
rect 110 2035 111 2039
rect 115 2035 116 2039
rect 110 2034 116 2035
rect 254 2036 260 2037
rect 112 2015 114 2034
rect 254 2032 255 2036
rect 259 2032 260 2036
rect 254 2031 260 2032
rect 256 2015 258 2031
rect 336 2020 338 2042
rect 374 2036 380 2037
rect 374 2032 375 2036
rect 379 2032 380 2036
rect 374 2031 380 2032
rect 334 2019 340 2020
rect 334 2015 335 2019
rect 339 2015 340 2019
rect 376 2015 378 2031
rect 456 2020 458 2042
rect 686 2039 687 2043
rect 691 2039 692 2043
rect 686 2038 692 2039
rect 494 2036 500 2037
rect 494 2032 495 2036
rect 499 2032 500 2036
rect 494 2031 500 2032
rect 614 2036 620 2037
rect 614 2032 615 2036
rect 619 2032 620 2036
rect 614 2031 620 2032
rect 454 2019 460 2020
rect 454 2015 455 2019
rect 459 2015 460 2019
rect 496 2015 498 2031
rect 550 2019 556 2020
rect 550 2015 551 2019
rect 555 2015 556 2019
rect 616 2015 618 2031
rect 688 2020 690 2038
rect 720 2028 722 2106
rect 742 2101 748 2102
rect 742 2097 743 2101
rect 747 2097 748 2101
rect 742 2096 748 2097
rect 862 2101 868 2102
rect 862 2097 863 2101
rect 867 2097 868 2101
rect 862 2096 868 2097
rect 982 2101 988 2102
rect 982 2097 983 2101
rect 987 2097 988 2101
rect 982 2096 988 2097
rect 744 2079 746 2096
rect 864 2079 866 2096
rect 984 2079 986 2096
rect 727 2078 731 2079
rect 727 2073 731 2074
rect 743 2078 747 2079
rect 743 2073 747 2074
rect 831 2078 835 2079
rect 831 2073 835 2074
rect 863 2078 867 2079
rect 863 2073 867 2074
rect 935 2078 939 2079
rect 935 2073 939 2074
rect 983 2078 987 2079
rect 983 2073 987 2074
rect 728 2056 730 2073
rect 832 2056 834 2073
rect 936 2056 938 2073
rect 726 2055 732 2056
rect 726 2051 727 2055
rect 731 2051 732 2055
rect 726 2050 732 2051
rect 830 2055 836 2056
rect 830 2051 831 2055
rect 835 2051 836 2055
rect 830 2050 836 2051
rect 934 2055 940 2056
rect 934 2051 935 2055
rect 939 2051 940 2055
rect 934 2050 940 2051
rect 1008 2048 1010 2130
rect 1768 2118 1770 2137
rect 1808 2135 1810 2159
rect 2184 2135 2186 2160
rect 2280 2135 2282 2160
rect 2384 2135 2386 2160
rect 2496 2135 2498 2160
rect 2608 2135 2610 2160
rect 1807 2134 1811 2135
rect 1807 2129 1811 2130
rect 2135 2134 2139 2135
rect 2135 2129 2139 2130
rect 2183 2134 2187 2135
rect 2183 2129 2187 2130
rect 2255 2134 2259 2135
rect 2255 2129 2259 2130
rect 2279 2134 2283 2135
rect 2279 2129 2283 2130
rect 2383 2134 2387 2135
rect 2383 2129 2387 2130
rect 2495 2134 2499 2135
rect 2495 2129 2499 2130
rect 2519 2134 2523 2135
rect 2519 2129 2523 2130
rect 2607 2134 2611 2135
rect 2607 2129 2611 2130
rect 2655 2134 2659 2135
rect 2655 2129 2659 2130
rect 1766 2117 1772 2118
rect 1766 2113 1767 2117
rect 1771 2113 1772 2117
rect 1808 2113 1810 2129
rect 1766 2112 1772 2113
rect 1806 2112 1812 2113
rect 2136 2112 2138 2129
rect 2256 2112 2258 2129
rect 2384 2112 2386 2129
rect 2520 2112 2522 2129
rect 2656 2112 2658 2129
rect 1806 2108 1807 2112
rect 1811 2108 1812 2112
rect 1806 2107 1812 2108
rect 2134 2111 2140 2112
rect 2134 2107 2135 2111
rect 2139 2107 2140 2111
rect 2134 2106 2140 2107
rect 2254 2111 2260 2112
rect 2254 2107 2255 2111
rect 2259 2107 2260 2111
rect 2254 2106 2260 2107
rect 2382 2111 2388 2112
rect 2382 2107 2383 2111
rect 2387 2107 2388 2111
rect 2382 2106 2388 2107
rect 2518 2111 2524 2112
rect 2518 2107 2519 2111
rect 2523 2107 2524 2111
rect 2518 2106 2524 2107
rect 2654 2111 2660 2112
rect 2654 2107 2655 2111
rect 2659 2107 2660 2111
rect 2654 2106 2660 2107
rect 2214 2103 2220 2104
rect 1766 2100 1772 2101
rect 1766 2096 1767 2100
rect 1771 2096 1772 2100
rect 2206 2099 2212 2100
rect 1766 2095 1772 2096
rect 1806 2095 1812 2096
rect 1768 2079 1770 2095
rect 1806 2091 1807 2095
rect 1811 2091 1812 2095
rect 2206 2095 2207 2099
rect 2211 2095 2212 2099
rect 2214 2099 2215 2103
rect 2219 2099 2220 2103
rect 2214 2098 2220 2099
rect 2334 2103 2340 2104
rect 2334 2099 2335 2103
rect 2339 2099 2340 2103
rect 2334 2098 2340 2099
rect 2462 2103 2468 2104
rect 2462 2099 2463 2103
rect 2467 2099 2468 2103
rect 2462 2098 2468 2099
rect 2598 2103 2604 2104
rect 2598 2099 2599 2103
rect 2603 2099 2604 2103
rect 2598 2098 2604 2099
rect 2206 2094 2212 2095
rect 1806 2090 1812 2091
rect 2134 2092 2140 2093
rect 1039 2078 1043 2079
rect 1039 2073 1043 2074
rect 1143 2078 1147 2079
rect 1143 2073 1147 2074
rect 1255 2078 1259 2079
rect 1255 2073 1259 2074
rect 1767 2078 1771 2079
rect 1767 2073 1771 2074
rect 1040 2056 1042 2073
rect 1144 2056 1146 2073
rect 1256 2056 1258 2073
rect 1768 2057 1770 2073
rect 1808 2063 1810 2090
rect 2134 2088 2135 2092
rect 2139 2088 2140 2092
rect 2134 2087 2140 2088
rect 2136 2063 2138 2087
rect 1807 2062 1811 2063
rect 1807 2057 1811 2058
rect 2135 2062 2139 2063
rect 2135 2057 2139 2058
rect 1766 2056 1772 2057
rect 1038 2055 1044 2056
rect 1038 2051 1039 2055
rect 1043 2051 1044 2055
rect 1038 2050 1044 2051
rect 1142 2055 1148 2056
rect 1142 2051 1143 2055
rect 1147 2051 1148 2055
rect 1142 2050 1148 2051
rect 1254 2055 1260 2056
rect 1254 2051 1255 2055
rect 1259 2051 1260 2055
rect 1766 2052 1767 2056
rect 1771 2052 1772 2056
rect 1766 2051 1772 2052
rect 1254 2050 1260 2051
rect 1006 2047 1012 2048
rect 798 2043 804 2044
rect 798 2039 799 2043
rect 803 2039 804 2043
rect 798 2038 804 2039
rect 902 2043 908 2044
rect 902 2039 903 2043
rect 907 2039 908 2043
rect 1006 2043 1007 2047
rect 1011 2043 1012 2047
rect 1006 2042 1012 2043
rect 1014 2047 1020 2048
rect 1014 2043 1015 2047
rect 1019 2043 1020 2047
rect 1014 2042 1020 2043
rect 1118 2047 1124 2048
rect 1118 2043 1119 2047
rect 1123 2043 1124 2047
rect 1118 2042 1124 2043
rect 1222 2047 1228 2048
rect 1222 2043 1223 2047
rect 1227 2043 1228 2047
rect 1222 2042 1228 2043
rect 902 2038 908 2039
rect 726 2036 732 2037
rect 726 2032 727 2036
rect 731 2032 732 2036
rect 726 2031 732 2032
rect 718 2027 724 2028
rect 718 2023 719 2027
rect 723 2023 724 2027
rect 718 2022 724 2023
rect 686 2019 692 2020
rect 686 2015 687 2019
rect 691 2015 692 2019
rect 728 2015 730 2031
rect 111 2014 115 2015
rect 111 2009 115 2010
rect 255 2014 259 2015
rect 334 2014 340 2015
rect 359 2014 363 2015
rect 255 2009 259 2010
rect 359 2009 363 2010
rect 375 2014 379 2015
rect 454 2014 460 2015
rect 487 2014 491 2015
rect 375 2009 379 2010
rect 487 2009 491 2010
rect 495 2014 499 2015
rect 550 2014 556 2015
rect 615 2014 619 2015
rect 495 2009 499 2010
rect 112 1990 114 2009
rect 360 1993 362 2009
rect 430 2007 436 2008
rect 430 2003 431 2007
rect 435 2003 436 2007
rect 430 2002 436 2003
rect 358 1992 364 1993
rect 110 1989 116 1990
rect 110 1985 111 1989
rect 115 1985 116 1989
rect 358 1988 359 1992
rect 363 1988 364 1992
rect 358 1987 364 1988
rect 110 1984 116 1985
rect 432 1984 434 2002
rect 488 1993 490 2009
rect 486 1992 492 1993
rect 486 1988 487 1992
rect 491 1988 492 1992
rect 486 1987 492 1988
rect 552 1984 554 2014
rect 615 2009 619 2010
rect 623 2014 627 2015
rect 686 2014 692 2015
rect 727 2014 731 2015
rect 623 2009 627 2010
rect 727 2009 731 2010
rect 759 2014 763 2015
rect 759 2009 763 2010
rect 624 1993 626 2009
rect 702 2007 708 2008
rect 702 2003 703 2007
rect 707 2003 708 2007
rect 702 2002 708 2003
rect 622 1992 628 1993
rect 622 1988 623 1992
rect 627 1988 628 1992
rect 622 1987 628 1988
rect 430 1983 436 1984
rect 430 1979 431 1983
rect 435 1979 436 1983
rect 430 1978 436 1979
rect 550 1983 556 1984
rect 550 1979 551 1983
rect 555 1979 556 1983
rect 550 1978 556 1979
rect 358 1973 364 1974
rect 110 1972 116 1973
rect 110 1968 111 1972
rect 115 1968 116 1972
rect 358 1969 359 1973
rect 363 1969 364 1973
rect 358 1968 364 1969
rect 486 1973 492 1974
rect 486 1969 487 1973
rect 491 1969 492 1973
rect 486 1968 492 1969
rect 622 1973 628 1974
rect 622 1969 623 1973
rect 627 1969 628 1973
rect 622 1968 628 1969
rect 110 1967 116 1968
rect 112 1951 114 1967
rect 360 1951 362 1968
rect 488 1951 490 1968
rect 624 1951 626 1968
rect 111 1950 115 1951
rect 111 1945 115 1946
rect 359 1950 363 1951
rect 359 1945 363 1946
rect 447 1950 451 1951
rect 447 1945 451 1946
rect 487 1950 491 1951
rect 487 1945 491 1946
rect 575 1950 579 1951
rect 575 1945 579 1946
rect 623 1950 627 1951
rect 623 1945 627 1946
rect 112 1929 114 1945
rect 110 1928 116 1929
rect 448 1928 450 1945
rect 576 1928 578 1945
rect 110 1924 111 1928
rect 115 1924 116 1928
rect 110 1923 116 1924
rect 446 1927 452 1928
rect 446 1923 447 1927
rect 451 1923 452 1927
rect 446 1922 452 1923
rect 574 1927 580 1928
rect 574 1923 575 1927
rect 579 1923 580 1927
rect 574 1922 580 1923
rect 704 1920 706 2002
rect 760 1993 762 2009
rect 800 2008 802 2038
rect 830 2036 836 2037
rect 830 2032 831 2036
rect 835 2032 836 2036
rect 830 2031 836 2032
rect 832 2015 834 2031
rect 904 2020 906 2038
rect 934 2036 940 2037
rect 934 2032 935 2036
rect 939 2032 940 2036
rect 934 2031 940 2032
rect 902 2019 908 2020
rect 902 2015 903 2019
rect 907 2015 908 2019
rect 936 2015 938 2031
rect 1016 2028 1018 2042
rect 1038 2036 1044 2037
rect 1038 2032 1039 2036
rect 1043 2032 1044 2036
rect 1038 2031 1044 2032
rect 1014 2027 1020 2028
rect 1014 2023 1015 2027
rect 1019 2023 1020 2027
rect 1014 2022 1020 2023
rect 1040 2015 1042 2031
rect 1120 2020 1122 2042
rect 1142 2036 1148 2037
rect 1142 2032 1143 2036
rect 1147 2032 1148 2036
rect 1142 2031 1148 2032
rect 1118 2019 1124 2020
rect 1118 2015 1119 2019
rect 1123 2015 1124 2019
rect 1144 2015 1146 2031
rect 1224 2020 1226 2042
rect 1766 2039 1772 2040
rect 1254 2036 1260 2037
rect 1254 2032 1255 2036
rect 1259 2032 1260 2036
rect 1766 2035 1767 2039
rect 1771 2035 1772 2039
rect 1808 2038 1810 2057
rect 2208 2056 2210 2094
rect 2216 2076 2218 2098
rect 2254 2092 2260 2093
rect 2254 2088 2255 2092
rect 2259 2088 2260 2092
rect 2254 2087 2260 2088
rect 2214 2075 2220 2076
rect 2214 2071 2215 2075
rect 2219 2071 2220 2075
rect 2214 2070 2220 2071
rect 2256 2063 2258 2087
rect 2336 2076 2338 2098
rect 2382 2092 2388 2093
rect 2382 2088 2383 2092
rect 2387 2088 2388 2092
rect 2382 2087 2388 2088
rect 2334 2075 2340 2076
rect 2334 2071 2335 2075
rect 2339 2071 2340 2075
rect 2334 2070 2340 2071
rect 2384 2063 2386 2087
rect 2464 2076 2466 2098
rect 2518 2092 2524 2093
rect 2518 2088 2519 2092
rect 2523 2088 2524 2092
rect 2518 2087 2524 2088
rect 2462 2075 2468 2076
rect 2462 2071 2463 2075
rect 2467 2071 2468 2075
rect 2462 2070 2468 2071
rect 2520 2063 2522 2087
rect 2600 2076 2602 2098
rect 2654 2092 2660 2093
rect 2654 2088 2655 2092
rect 2659 2088 2660 2092
rect 2654 2087 2660 2088
rect 2598 2075 2604 2076
rect 2598 2071 2599 2075
rect 2603 2071 2604 2075
rect 2598 2070 2604 2071
rect 2656 2063 2658 2087
rect 2680 2076 2682 2170
rect 2718 2165 2724 2166
rect 2718 2161 2719 2165
rect 2723 2161 2724 2165
rect 2718 2160 2724 2161
rect 2838 2165 2844 2166
rect 2838 2161 2839 2165
rect 2843 2161 2844 2165
rect 2838 2160 2844 2161
rect 2966 2165 2972 2166
rect 2966 2161 2967 2165
rect 2971 2161 2972 2165
rect 2966 2160 2972 2161
rect 3102 2165 3108 2166
rect 3102 2161 3103 2165
rect 3107 2161 3108 2165
rect 3102 2160 3108 2161
rect 2720 2135 2722 2160
rect 2840 2135 2842 2160
rect 2968 2135 2970 2160
rect 3104 2135 3106 2160
rect 2719 2134 2723 2135
rect 2719 2129 2723 2130
rect 2783 2134 2787 2135
rect 2783 2129 2787 2130
rect 2839 2134 2843 2135
rect 2839 2129 2843 2130
rect 2911 2134 2915 2135
rect 2911 2129 2915 2130
rect 2967 2134 2971 2135
rect 2967 2129 2971 2130
rect 3031 2134 3035 2135
rect 3031 2129 3035 2130
rect 3103 2134 3107 2135
rect 3103 2129 3107 2130
rect 2784 2112 2786 2129
rect 2912 2112 2914 2129
rect 3032 2112 3034 2129
rect 2782 2111 2788 2112
rect 2782 2107 2783 2111
rect 2787 2107 2788 2111
rect 2782 2106 2788 2107
rect 2910 2111 2916 2112
rect 2910 2107 2911 2111
rect 2915 2107 2916 2111
rect 2910 2106 2916 2107
rect 3030 2111 3036 2112
rect 3030 2107 3031 2111
rect 3035 2107 3036 2111
rect 3030 2106 3036 2107
rect 3116 2104 3118 2194
rect 3176 2176 3178 2194
rect 3248 2185 3250 2201
rect 3246 2184 3252 2185
rect 3246 2180 3247 2184
rect 3251 2180 3252 2184
rect 3246 2179 3252 2180
rect 3174 2175 3180 2176
rect 3174 2171 3175 2175
rect 3179 2171 3180 2175
rect 3174 2170 3180 2171
rect 3246 2165 3252 2166
rect 3246 2161 3247 2165
rect 3251 2161 3252 2165
rect 3246 2160 3252 2161
rect 3248 2135 3250 2160
rect 3151 2134 3155 2135
rect 3151 2129 3155 2130
rect 3247 2134 3251 2135
rect 3247 2129 3251 2130
rect 3271 2134 3275 2135
rect 3271 2129 3275 2130
rect 3152 2112 3154 2129
rect 3272 2112 3274 2129
rect 3150 2111 3156 2112
rect 3150 2107 3151 2111
rect 3155 2107 3156 2111
rect 3150 2106 3156 2107
rect 3270 2111 3276 2112
rect 3270 2107 3271 2111
rect 3275 2107 3276 2111
rect 3270 2106 3276 2107
rect 3114 2103 3120 2104
rect 2854 2099 2860 2100
rect 2854 2095 2855 2099
rect 2859 2095 2860 2099
rect 2854 2094 2860 2095
rect 2982 2099 2988 2100
rect 2982 2095 2983 2099
rect 2987 2095 2988 2099
rect 3114 2099 3115 2103
rect 3119 2099 3120 2103
rect 3114 2098 3120 2099
rect 3122 2103 3128 2104
rect 3122 2099 3123 2103
rect 3127 2099 3128 2103
rect 3122 2098 3128 2099
rect 3230 2103 3236 2104
rect 3230 2099 3231 2103
rect 3235 2099 3236 2103
rect 3230 2098 3236 2099
rect 2982 2094 2988 2095
rect 2782 2092 2788 2093
rect 2782 2088 2783 2092
rect 2787 2088 2788 2092
rect 2782 2087 2788 2088
rect 2678 2075 2684 2076
rect 2678 2071 2679 2075
rect 2683 2071 2684 2075
rect 2678 2070 2684 2071
rect 2784 2063 2786 2087
rect 2856 2076 2858 2094
rect 2910 2092 2916 2093
rect 2910 2088 2911 2092
rect 2915 2088 2916 2092
rect 2910 2087 2916 2088
rect 2854 2075 2860 2076
rect 2854 2071 2855 2075
rect 2859 2071 2860 2075
rect 2854 2070 2860 2071
rect 2912 2063 2914 2087
rect 2984 2076 2986 2094
rect 3030 2092 3036 2093
rect 3030 2088 3031 2092
rect 3035 2088 3036 2092
rect 3030 2087 3036 2088
rect 2982 2075 2988 2076
rect 2982 2071 2983 2075
rect 2987 2071 2988 2075
rect 2982 2070 2988 2071
rect 3032 2063 3034 2087
rect 3124 2084 3126 2098
rect 3150 2092 3156 2093
rect 3150 2088 3151 2092
rect 3155 2088 3156 2092
rect 3150 2087 3156 2088
rect 3122 2083 3128 2084
rect 3122 2079 3123 2083
rect 3127 2079 3128 2083
rect 3122 2078 3128 2079
rect 3152 2063 3154 2087
rect 3232 2076 3234 2098
rect 3270 2092 3276 2093
rect 3270 2088 3271 2092
rect 3275 2088 3276 2092
rect 3270 2087 3276 2088
rect 3230 2075 3236 2076
rect 3230 2071 3231 2075
rect 3235 2071 3236 2075
rect 3230 2070 3236 2071
rect 3272 2063 3274 2087
rect 3340 2076 3342 2242
rect 3366 2240 3372 2241
rect 3366 2236 3367 2240
rect 3371 2236 3372 2240
rect 3462 2239 3463 2243
rect 3467 2239 3468 2243
rect 3462 2238 3468 2239
rect 3366 2235 3372 2236
rect 3368 2207 3370 2235
rect 3430 2223 3436 2224
rect 3430 2219 3431 2223
rect 3435 2219 3436 2223
rect 3430 2218 3436 2219
rect 3367 2206 3371 2207
rect 3367 2201 3371 2202
rect 3368 2185 3370 2201
rect 3366 2184 3372 2185
rect 3366 2180 3367 2184
rect 3371 2180 3372 2184
rect 3366 2179 3372 2180
rect 3432 2176 3434 2218
rect 3464 2207 3466 2238
rect 3463 2206 3467 2207
rect 3463 2201 3467 2202
rect 3438 2199 3444 2200
rect 3438 2195 3439 2199
rect 3443 2195 3444 2199
rect 3438 2194 3444 2195
rect 3430 2175 3436 2176
rect 3430 2171 3431 2175
rect 3435 2171 3436 2175
rect 3430 2170 3436 2171
rect 3366 2165 3372 2166
rect 3366 2161 3367 2165
rect 3371 2161 3372 2165
rect 3366 2160 3372 2161
rect 3368 2135 3370 2160
rect 3367 2134 3371 2135
rect 3367 2129 3371 2130
rect 3368 2112 3370 2129
rect 3366 2111 3372 2112
rect 3366 2107 3367 2111
rect 3371 2107 3372 2111
rect 3366 2106 3372 2107
rect 3358 2103 3364 2104
rect 3358 2099 3359 2103
rect 3363 2099 3364 2103
rect 3358 2098 3364 2099
rect 3326 2075 3332 2076
rect 3326 2071 3327 2075
rect 3331 2071 3332 2075
rect 3326 2070 3332 2071
rect 3338 2075 3344 2076
rect 3338 2071 3339 2075
rect 3343 2071 3344 2075
rect 3338 2070 3344 2071
rect 2247 2062 2251 2063
rect 2247 2057 2251 2058
rect 2255 2062 2259 2063
rect 2255 2057 2259 2058
rect 2383 2062 2387 2063
rect 2383 2057 2387 2058
rect 2415 2062 2419 2063
rect 2415 2057 2419 2058
rect 2519 2062 2523 2063
rect 2519 2057 2523 2058
rect 2575 2062 2579 2063
rect 2575 2057 2579 2058
rect 2655 2062 2659 2063
rect 2655 2057 2659 2058
rect 2727 2062 2731 2063
rect 2727 2057 2731 2058
rect 2783 2062 2787 2063
rect 2783 2057 2787 2058
rect 2871 2062 2875 2063
rect 2871 2057 2875 2058
rect 2911 2062 2915 2063
rect 2911 2057 2915 2058
rect 3007 2062 3011 2063
rect 3007 2057 3011 2058
rect 3031 2062 3035 2063
rect 3031 2057 3035 2058
rect 3135 2062 3139 2063
rect 3135 2057 3139 2058
rect 3151 2062 3155 2063
rect 3151 2057 3155 2058
rect 3263 2062 3267 2063
rect 3263 2057 3267 2058
rect 3271 2062 3275 2063
rect 3271 2057 3275 2058
rect 2206 2055 2212 2056
rect 2206 2051 2207 2055
rect 2211 2051 2212 2055
rect 2206 2050 2212 2051
rect 2248 2041 2250 2057
rect 2318 2055 2324 2056
rect 2318 2051 2319 2055
rect 2323 2051 2324 2055
rect 2318 2050 2324 2051
rect 2246 2040 2252 2041
rect 1766 2034 1772 2035
rect 1806 2037 1812 2038
rect 1254 2031 1260 2032
rect 1222 2019 1228 2020
rect 1222 2015 1223 2019
rect 1227 2015 1228 2019
rect 1256 2015 1258 2031
rect 1768 2015 1770 2034
rect 1806 2033 1807 2037
rect 1811 2033 1812 2037
rect 2246 2036 2247 2040
rect 2251 2036 2252 2040
rect 2246 2035 2252 2036
rect 1806 2032 1812 2033
rect 2320 2032 2322 2050
rect 2416 2041 2418 2057
rect 2486 2055 2492 2056
rect 2486 2051 2487 2055
rect 2491 2051 2492 2055
rect 2486 2050 2492 2051
rect 2414 2040 2420 2041
rect 2414 2036 2415 2040
rect 2419 2036 2420 2040
rect 2414 2035 2420 2036
rect 2488 2032 2490 2050
rect 2576 2041 2578 2057
rect 2728 2041 2730 2057
rect 2798 2055 2804 2056
rect 2798 2051 2799 2055
rect 2803 2051 2804 2055
rect 2798 2050 2804 2051
rect 2574 2040 2580 2041
rect 2574 2036 2575 2040
rect 2579 2036 2580 2040
rect 2574 2035 2580 2036
rect 2726 2040 2732 2041
rect 2726 2036 2727 2040
rect 2731 2036 2732 2040
rect 2726 2035 2732 2036
rect 2800 2032 2802 2050
rect 2872 2041 2874 2057
rect 2942 2055 2948 2056
rect 2942 2051 2943 2055
rect 2947 2051 2948 2055
rect 2942 2050 2948 2051
rect 2870 2040 2876 2041
rect 2870 2036 2871 2040
rect 2875 2036 2876 2040
rect 2870 2035 2876 2036
rect 2944 2032 2946 2050
rect 3008 2041 3010 2057
rect 3078 2055 3084 2056
rect 3078 2051 3079 2055
rect 3083 2051 3084 2055
rect 3078 2050 3084 2051
rect 3006 2040 3012 2041
rect 3006 2036 3007 2040
rect 3011 2036 3012 2040
rect 3006 2035 3012 2036
rect 3080 2032 3082 2050
rect 3110 2047 3116 2048
rect 3110 2043 3111 2047
rect 3115 2043 3116 2047
rect 3110 2042 3116 2043
rect 2318 2031 2324 2032
rect 2318 2027 2319 2031
rect 2323 2027 2324 2031
rect 2318 2026 2324 2027
rect 2486 2031 2492 2032
rect 2486 2027 2487 2031
rect 2491 2027 2492 2031
rect 2486 2026 2492 2027
rect 2526 2031 2532 2032
rect 2526 2027 2527 2031
rect 2531 2027 2532 2031
rect 2526 2026 2532 2027
rect 2798 2031 2804 2032
rect 2798 2027 2799 2031
rect 2803 2027 2804 2031
rect 2798 2026 2804 2027
rect 2942 2031 2948 2032
rect 2942 2027 2943 2031
rect 2947 2027 2948 2031
rect 2942 2026 2948 2027
rect 3078 2031 3084 2032
rect 3078 2027 3079 2031
rect 3083 2027 3084 2031
rect 3078 2026 3084 2027
rect 2246 2021 2252 2022
rect 1806 2020 1812 2021
rect 1806 2016 1807 2020
rect 1811 2016 1812 2020
rect 2246 2017 2247 2021
rect 2251 2017 2252 2021
rect 2246 2016 2252 2017
rect 2414 2021 2420 2022
rect 2414 2017 2415 2021
rect 2419 2017 2420 2021
rect 2414 2016 2420 2017
rect 1806 2015 1812 2016
rect 831 2014 835 2015
rect 831 2009 835 2010
rect 895 2014 899 2015
rect 902 2014 908 2015
rect 935 2014 939 2015
rect 895 2009 899 2010
rect 935 2009 939 2010
rect 1023 2014 1027 2015
rect 1023 2009 1027 2010
rect 1039 2014 1043 2015
rect 1118 2014 1124 2015
rect 1143 2014 1147 2015
rect 1039 2009 1043 2010
rect 1143 2009 1147 2010
rect 1151 2014 1155 2015
rect 1222 2014 1228 2015
rect 1255 2014 1259 2015
rect 1151 2009 1155 2010
rect 1255 2009 1259 2010
rect 1271 2014 1275 2015
rect 1271 2009 1275 2010
rect 1399 2014 1403 2015
rect 1399 2009 1403 2010
rect 1527 2014 1531 2015
rect 1527 2009 1531 2010
rect 1767 2014 1771 2015
rect 1767 2009 1771 2010
rect 798 2007 804 2008
rect 798 2003 799 2007
rect 803 2003 804 2007
rect 798 2002 804 2003
rect 896 1993 898 2009
rect 1024 1993 1026 2009
rect 1094 2007 1100 2008
rect 1094 2003 1095 2007
rect 1099 2003 1100 2007
rect 1094 2002 1100 2003
rect 758 1992 764 1993
rect 758 1988 759 1992
rect 763 1988 764 1992
rect 758 1987 764 1988
rect 894 1992 900 1993
rect 894 1988 895 1992
rect 899 1988 900 1992
rect 894 1987 900 1988
rect 1022 1992 1028 1993
rect 1022 1988 1023 1992
rect 1027 1988 1028 1992
rect 1022 1987 1028 1988
rect 1096 1984 1098 2002
rect 1152 1993 1154 2009
rect 1272 1993 1274 2009
rect 1350 2007 1356 2008
rect 1350 2003 1351 2007
rect 1355 2003 1356 2007
rect 1350 2002 1356 2003
rect 1150 1992 1156 1993
rect 1150 1988 1151 1992
rect 1155 1988 1156 1992
rect 1150 1987 1156 1988
rect 1270 1992 1276 1993
rect 1270 1988 1271 1992
rect 1275 1988 1276 1992
rect 1270 1987 1276 1988
rect 1352 1984 1354 2002
rect 1400 1993 1402 2009
rect 1486 2007 1492 2008
rect 1486 2003 1487 2007
rect 1491 2003 1492 2007
rect 1486 2002 1492 2003
rect 1398 1992 1404 1993
rect 1398 1988 1399 1992
rect 1403 1988 1404 1992
rect 1398 1987 1404 1988
rect 1488 1984 1490 2002
rect 1528 1993 1530 2009
rect 1598 2007 1604 2008
rect 1598 2003 1599 2007
rect 1603 2003 1604 2007
rect 1598 2002 1604 2003
rect 1526 1992 1532 1993
rect 1526 1988 1527 1992
rect 1531 1988 1532 1992
rect 1526 1987 1532 1988
rect 966 1983 972 1984
rect 966 1979 967 1983
rect 971 1979 972 1983
rect 966 1978 972 1979
rect 1094 1983 1100 1984
rect 1094 1979 1095 1983
rect 1099 1979 1100 1983
rect 1094 1978 1100 1979
rect 1350 1983 1356 1984
rect 1350 1979 1351 1983
rect 1355 1979 1356 1983
rect 1350 1978 1356 1979
rect 1486 1983 1492 1984
rect 1486 1979 1487 1983
rect 1491 1979 1492 1983
rect 1486 1978 1492 1979
rect 758 1973 764 1974
rect 758 1969 759 1973
rect 763 1969 764 1973
rect 758 1968 764 1969
rect 894 1973 900 1974
rect 894 1969 895 1973
rect 899 1969 900 1973
rect 894 1968 900 1969
rect 760 1951 762 1968
rect 896 1951 898 1968
rect 711 1950 715 1951
rect 711 1945 715 1946
rect 759 1950 763 1951
rect 759 1945 763 1946
rect 847 1950 851 1951
rect 847 1945 851 1946
rect 895 1950 899 1951
rect 895 1945 899 1946
rect 712 1928 714 1945
rect 848 1928 850 1945
rect 710 1927 716 1928
rect 710 1923 711 1927
rect 715 1923 716 1927
rect 710 1922 716 1923
rect 846 1927 852 1928
rect 846 1923 847 1927
rect 851 1923 852 1927
rect 846 1922 852 1923
rect 702 1919 708 1920
rect 646 1915 652 1916
rect 110 1911 116 1912
rect 110 1907 111 1911
rect 115 1907 116 1911
rect 646 1911 647 1915
rect 651 1911 652 1915
rect 702 1915 703 1919
rect 707 1915 708 1919
rect 926 1919 932 1920
rect 702 1914 708 1915
rect 918 1915 924 1916
rect 646 1910 652 1911
rect 918 1911 919 1915
rect 923 1911 924 1915
rect 926 1915 927 1919
rect 931 1915 932 1919
rect 926 1914 932 1915
rect 918 1910 924 1911
rect 110 1906 116 1907
rect 446 1908 452 1909
rect 112 1887 114 1906
rect 446 1904 447 1908
rect 451 1904 452 1908
rect 446 1903 452 1904
rect 574 1908 580 1909
rect 574 1904 575 1908
rect 579 1904 580 1908
rect 574 1903 580 1904
rect 448 1887 450 1903
rect 538 1891 544 1892
rect 538 1887 539 1891
rect 543 1887 544 1891
rect 576 1887 578 1903
rect 648 1892 650 1910
rect 710 1908 716 1909
rect 710 1904 711 1908
rect 715 1904 716 1908
rect 710 1903 716 1904
rect 846 1908 852 1909
rect 846 1904 847 1908
rect 851 1904 852 1908
rect 846 1903 852 1904
rect 646 1891 652 1892
rect 646 1887 647 1891
rect 651 1887 652 1891
rect 712 1887 714 1903
rect 848 1887 850 1903
rect 111 1886 115 1887
rect 111 1881 115 1882
rect 447 1886 451 1887
rect 538 1886 544 1887
rect 559 1886 563 1887
rect 447 1881 451 1882
rect 112 1862 114 1881
rect 110 1861 116 1862
rect 110 1857 111 1861
rect 115 1857 116 1861
rect 110 1856 116 1857
rect 540 1856 542 1886
rect 559 1881 563 1882
rect 575 1886 579 1887
rect 646 1886 652 1887
rect 695 1886 699 1887
rect 575 1881 579 1882
rect 695 1881 699 1882
rect 711 1886 715 1887
rect 711 1881 715 1882
rect 831 1886 835 1887
rect 831 1881 835 1882
rect 847 1886 851 1887
rect 847 1881 851 1882
rect 560 1865 562 1881
rect 646 1879 652 1880
rect 646 1875 647 1879
rect 651 1875 652 1879
rect 646 1874 652 1875
rect 558 1864 564 1865
rect 558 1860 559 1864
rect 563 1860 564 1864
rect 558 1859 564 1860
rect 648 1856 650 1874
rect 696 1865 698 1881
rect 774 1879 780 1880
rect 774 1875 775 1879
rect 779 1875 780 1879
rect 774 1874 780 1875
rect 694 1864 700 1865
rect 694 1860 695 1864
rect 699 1860 700 1864
rect 694 1859 700 1860
rect 776 1856 778 1874
rect 832 1865 834 1881
rect 920 1880 922 1910
rect 928 1892 930 1914
rect 968 1892 970 1978
rect 1022 1973 1028 1974
rect 1022 1969 1023 1973
rect 1027 1969 1028 1973
rect 1022 1968 1028 1969
rect 1150 1973 1156 1974
rect 1150 1969 1151 1973
rect 1155 1969 1156 1973
rect 1150 1968 1156 1969
rect 1270 1973 1276 1974
rect 1270 1969 1271 1973
rect 1275 1969 1276 1973
rect 1270 1968 1276 1969
rect 1398 1973 1404 1974
rect 1398 1969 1399 1973
rect 1403 1969 1404 1973
rect 1398 1968 1404 1969
rect 1526 1973 1532 1974
rect 1526 1969 1527 1973
rect 1531 1969 1532 1973
rect 1526 1968 1532 1969
rect 1024 1951 1026 1968
rect 1152 1951 1154 1968
rect 1272 1951 1274 1968
rect 1400 1951 1402 1968
rect 1528 1951 1530 1968
rect 983 1950 987 1951
rect 983 1945 987 1946
rect 1023 1950 1027 1951
rect 1023 1945 1027 1946
rect 1119 1950 1123 1951
rect 1119 1945 1123 1946
rect 1151 1950 1155 1951
rect 1151 1945 1155 1946
rect 1255 1950 1259 1951
rect 1255 1945 1259 1946
rect 1271 1950 1275 1951
rect 1271 1945 1275 1946
rect 1383 1950 1387 1951
rect 1383 1945 1387 1946
rect 1399 1950 1403 1951
rect 1399 1945 1403 1946
rect 1519 1950 1523 1951
rect 1519 1945 1523 1946
rect 1527 1950 1531 1951
rect 1527 1945 1531 1946
rect 984 1928 986 1945
rect 1120 1928 1122 1945
rect 1256 1928 1258 1945
rect 1384 1928 1386 1945
rect 1520 1928 1522 1945
rect 982 1927 988 1928
rect 982 1923 983 1927
rect 987 1923 988 1927
rect 982 1922 988 1923
rect 1118 1927 1124 1928
rect 1118 1923 1119 1927
rect 1123 1923 1124 1927
rect 1118 1922 1124 1923
rect 1254 1927 1260 1928
rect 1254 1923 1255 1927
rect 1259 1923 1260 1927
rect 1254 1922 1260 1923
rect 1382 1927 1388 1928
rect 1382 1923 1383 1927
rect 1387 1923 1388 1927
rect 1382 1922 1388 1923
rect 1518 1927 1524 1928
rect 1518 1923 1519 1927
rect 1523 1923 1524 1927
rect 1518 1922 1524 1923
rect 1600 1920 1602 2002
rect 1768 1990 1770 2009
rect 1766 1989 1772 1990
rect 1766 1985 1767 1989
rect 1771 1985 1772 1989
rect 1766 1984 1772 1985
rect 1808 1983 1810 2015
rect 2248 1983 2250 2016
rect 2416 1983 2418 2016
rect 1807 1982 1811 1983
rect 1807 1977 1811 1978
rect 1831 1982 1835 1983
rect 1831 1977 1835 1978
rect 1919 1982 1923 1983
rect 1919 1977 1923 1978
rect 2047 1982 2051 1983
rect 2047 1977 2051 1978
rect 2183 1982 2187 1983
rect 2183 1977 2187 1978
rect 2247 1982 2251 1983
rect 2247 1977 2251 1978
rect 2327 1982 2331 1983
rect 2327 1977 2331 1978
rect 2415 1982 2419 1983
rect 2415 1977 2419 1978
rect 2471 1982 2475 1983
rect 2471 1977 2475 1978
rect 1766 1972 1772 1973
rect 1766 1968 1767 1972
rect 1771 1968 1772 1972
rect 1766 1967 1772 1968
rect 1768 1951 1770 1967
rect 1808 1961 1810 1977
rect 1806 1960 1812 1961
rect 1832 1960 1834 1977
rect 1920 1960 1922 1977
rect 2048 1960 2050 1977
rect 2184 1960 2186 1977
rect 2328 1960 2330 1977
rect 2472 1960 2474 1977
rect 1806 1956 1807 1960
rect 1811 1956 1812 1960
rect 1806 1955 1812 1956
rect 1830 1959 1836 1960
rect 1830 1955 1831 1959
rect 1835 1955 1836 1959
rect 1830 1954 1836 1955
rect 1918 1959 1924 1960
rect 1918 1955 1919 1959
rect 1923 1955 1924 1959
rect 1918 1954 1924 1955
rect 2046 1959 2052 1960
rect 2046 1955 2047 1959
rect 2051 1955 2052 1959
rect 2046 1954 2052 1955
rect 2182 1959 2188 1960
rect 2182 1955 2183 1959
rect 2187 1955 2188 1959
rect 2182 1954 2188 1955
rect 2326 1959 2332 1960
rect 2326 1955 2327 1959
rect 2331 1955 2332 1959
rect 2326 1954 2332 1955
rect 2470 1959 2476 1960
rect 2470 1955 2471 1959
rect 2475 1955 2476 1959
rect 2470 1954 2476 1955
rect 1910 1951 1916 1952
rect 1655 1950 1659 1951
rect 1655 1945 1659 1946
rect 1767 1950 1771 1951
rect 1767 1945 1771 1946
rect 1902 1947 1908 1948
rect 1656 1928 1658 1945
rect 1768 1929 1770 1945
rect 1806 1943 1812 1944
rect 1806 1939 1807 1943
rect 1811 1939 1812 1943
rect 1902 1943 1903 1947
rect 1907 1943 1908 1947
rect 1910 1947 1911 1951
rect 1915 1947 1916 1951
rect 1910 1946 1916 1947
rect 1998 1951 2004 1952
rect 1998 1947 1999 1951
rect 2003 1947 2004 1951
rect 1998 1946 2004 1947
rect 2126 1951 2132 1952
rect 2126 1947 2127 1951
rect 2131 1947 2132 1951
rect 2126 1946 2132 1947
rect 2262 1951 2268 1952
rect 2262 1947 2263 1951
rect 2267 1947 2268 1951
rect 2262 1946 2268 1947
rect 1902 1942 1908 1943
rect 1806 1938 1812 1939
rect 1830 1940 1836 1941
rect 1766 1928 1772 1929
rect 1654 1927 1660 1928
rect 1654 1923 1655 1927
rect 1659 1923 1660 1927
rect 1766 1924 1767 1928
rect 1771 1924 1772 1928
rect 1766 1923 1772 1924
rect 1654 1922 1660 1923
rect 1598 1919 1604 1920
rect 1190 1915 1196 1916
rect 1190 1911 1191 1915
rect 1195 1911 1196 1915
rect 1190 1910 1196 1911
rect 1366 1915 1372 1916
rect 1366 1911 1367 1915
rect 1371 1911 1372 1915
rect 1366 1910 1372 1911
rect 1470 1915 1476 1916
rect 1470 1911 1471 1915
rect 1475 1911 1476 1915
rect 1470 1910 1476 1911
rect 1590 1915 1596 1916
rect 1590 1911 1591 1915
rect 1595 1911 1596 1915
rect 1598 1915 1599 1919
rect 1603 1915 1604 1919
rect 1808 1915 1810 1938
rect 1830 1936 1831 1940
rect 1835 1936 1836 1940
rect 1830 1935 1836 1936
rect 1832 1915 1834 1935
rect 1904 1916 1906 1942
rect 1912 1924 1914 1946
rect 1918 1940 1924 1941
rect 1918 1936 1919 1940
rect 1923 1936 1924 1940
rect 1918 1935 1924 1936
rect 1910 1923 1916 1924
rect 1910 1919 1911 1923
rect 1915 1919 1916 1923
rect 1910 1918 1916 1919
rect 1902 1915 1908 1916
rect 1920 1915 1922 1935
rect 2000 1924 2002 1946
rect 2046 1940 2052 1941
rect 2046 1936 2047 1940
rect 2051 1936 2052 1940
rect 2046 1935 2052 1936
rect 1998 1923 2004 1924
rect 1998 1919 1999 1923
rect 2003 1919 2004 1923
rect 1998 1918 2004 1919
rect 2048 1915 2050 1935
rect 2128 1924 2130 1946
rect 2182 1940 2188 1941
rect 2182 1936 2183 1940
rect 2187 1936 2188 1940
rect 2182 1935 2188 1936
rect 2126 1923 2132 1924
rect 2126 1919 2127 1923
rect 2131 1919 2132 1923
rect 2126 1918 2132 1919
rect 2184 1915 2186 1935
rect 2264 1924 2266 1946
rect 2326 1940 2332 1941
rect 2326 1936 2327 1940
rect 2331 1936 2332 1940
rect 2326 1935 2332 1936
rect 2470 1940 2476 1941
rect 2470 1936 2471 1940
rect 2475 1936 2476 1940
rect 2470 1935 2476 1936
rect 2262 1923 2268 1924
rect 2262 1919 2263 1923
rect 2267 1919 2268 1923
rect 2262 1918 2268 1919
rect 2328 1915 2330 1935
rect 2374 1923 2380 1924
rect 2374 1919 2375 1923
rect 2379 1919 2380 1923
rect 2374 1918 2380 1919
rect 1598 1914 1604 1915
rect 1807 1914 1811 1915
rect 1590 1910 1596 1911
rect 1766 1911 1772 1912
rect 982 1908 988 1909
rect 982 1904 983 1908
rect 987 1904 988 1908
rect 982 1903 988 1904
rect 1118 1908 1124 1909
rect 1118 1904 1119 1908
rect 1123 1904 1124 1908
rect 1118 1903 1124 1904
rect 926 1891 932 1892
rect 926 1887 927 1891
rect 931 1887 932 1891
rect 966 1891 972 1892
rect 966 1887 967 1891
rect 971 1887 972 1891
rect 984 1887 986 1903
rect 1120 1887 1122 1903
rect 1192 1892 1194 1910
rect 1254 1908 1260 1909
rect 1254 1904 1255 1908
rect 1259 1904 1260 1908
rect 1254 1903 1260 1904
rect 1190 1891 1196 1892
rect 1190 1887 1191 1891
rect 1195 1887 1196 1891
rect 1256 1887 1258 1903
rect 1368 1892 1370 1910
rect 1382 1908 1388 1909
rect 1382 1904 1383 1908
rect 1387 1904 1388 1908
rect 1382 1903 1388 1904
rect 1366 1891 1372 1892
rect 1366 1887 1367 1891
rect 1371 1887 1372 1891
rect 1384 1887 1386 1903
rect 1406 1899 1412 1900
rect 1406 1895 1407 1899
rect 1411 1895 1412 1899
rect 1406 1894 1412 1895
rect 926 1886 932 1887
rect 959 1886 963 1887
rect 966 1886 972 1887
rect 983 1886 987 1887
rect 959 1881 963 1882
rect 983 1881 987 1882
rect 1079 1886 1083 1887
rect 1079 1881 1083 1882
rect 1119 1886 1123 1887
rect 1190 1886 1196 1887
rect 1199 1886 1203 1887
rect 1119 1881 1123 1882
rect 1199 1881 1203 1882
rect 1255 1886 1259 1887
rect 1255 1881 1259 1882
rect 1327 1886 1331 1887
rect 1366 1886 1372 1887
rect 1383 1886 1387 1887
rect 1327 1881 1331 1882
rect 1383 1881 1387 1882
rect 918 1879 924 1880
rect 918 1875 919 1879
rect 923 1875 924 1879
rect 918 1874 924 1875
rect 960 1865 962 1881
rect 1030 1879 1036 1880
rect 1030 1875 1031 1879
rect 1035 1875 1036 1879
rect 1030 1874 1036 1875
rect 830 1864 836 1865
rect 830 1860 831 1864
rect 835 1860 836 1864
rect 830 1859 836 1860
rect 958 1864 964 1865
rect 958 1860 959 1864
rect 963 1860 964 1864
rect 958 1859 964 1860
rect 1032 1856 1034 1874
rect 1080 1865 1082 1881
rect 1150 1879 1156 1880
rect 1150 1875 1151 1879
rect 1155 1875 1156 1879
rect 1150 1874 1156 1875
rect 1078 1864 1084 1865
rect 1078 1860 1079 1864
rect 1083 1860 1084 1864
rect 1078 1859 1084 1860
rect 1152 1856 1154 1874
rect 1166 1871 1172 1872
rect 1166 1867 1167 1871
rect 1171 1867 1172 1871
rect 1166 1866 1172 1867
rect 538 1855 544 1856
rect 538 1851 539 1855
rect 543 1851 544 1855
rect 538 1850 544 1851
rect 646 1855 652 1856
rect 646 1851 647 1855
rect 651 1851 652 1855
rect 646 1850 652 1851
rect 774 1855 780 1856
rect 774 1851 775 1855
rect 779 1851 780 1855
rect 774 1850 780 1851
rect 1030 1855 1036 1856
rect 1030 1851 1031 1855
rect 1035 1851 1036 1855
rect 1030 1850 1036 1851
rect 1150 1855 1156 1856
rect 1150 1851 1151 1855
rect 1155 1851 1156 1855
rect 1150 1850 1156 1851
rect 558 1845 564 1846
rect 110 1844 116 1845
rect 110 1840 111 1844
rect 115 1840 116 1844
rect 558 1841 559 1845
rect 563 1841 564 1845
rect 558 1840 564 1841
rect 694 1845 700 1846
rect 694 1841 695 1845
rect 699 1841 700 1845
rect 694 1840 700 1841
rect 830 1845 836 1846
rect 830 1841 831 1845
rect 835 1841 836 1845
rect 830 1840 836 1841
rect 958 1845 964 1846
rect 958 1841 959 1845
rect 963 1841 964 1845
rect 958 1840 964 1841
rect 1078 1845 1084 1846
rect 1078 1841 1079 1845
rect 1083 1841 1084 1845
rect 1078 1840 1084 1841
rect 110 1839 116 1840
rect 112 1815 114 1839
rect 560 1815 562 1840
rect 696 1815 698 1840
rect 832 1815 834 1840
rect 960 1815 962 1840
rect 1080 1815 1082 1840
rect 111 1814 115 1815
rect 111 1809 115 1810
rect 135 1814 139 1815
rect 135 1809 139 1810
rect 223 1814 227 1815
rect 223 1809 227 1810
rect 311 1814 315 1815
rect 311 1809 315 1810
rect 407 1814 411 1815
rect 407 1809 411 1810
rect 527 1814 531 1815
rect 527 1809 531 1810
rect 559 1814 563 1815
rect 559 1809 563 1810
rect 655 1814 659 1815
rect 655 1809 659 1810
rect 695 1814 699 1815
rect 695 1809 699 1810
rect 799 1814 803 1815
rect 799 1809 803 1810
rect 831 1814 835 1815
rect 831 1809 835 1810
rect 943 1814 947 1815
rect 943 1809 947 1810
rect 959 1814 963 1815
rect 959 1809 963 1810
rect 1079 1814 1083 1815
rect 1079 1809 1083 1810
rect 1087 1814 1091 1815
rect 1087 1809 1091 1810
rect 112 1793 114 1809
rect 110 1792 116 1793
rect 136 1792 138 1809
rect 224 1792 226 1809
rect 312 1792 314 1809
rect 408 1792 410 1809
rect 528 1792 530 1809
rect 656 1792 658 1809
rect 800 1792 802 1809
rect 944 1792 946 1809
rect 1088 1792 1090 1809
rect 110 1788 111 1792
rect 115 1788 116 1792
rect 110 1787 116 1788
rect 134 1791 140 1792
rect 134 1787 135 1791
rect 139 1787 140 1791
rect 134 1786 140 1787
rect 222 1791 228 1792
rect 222 1787 223 1791
rect 227 1787 228 1791
rect 222 1786 228 1787
rect 310 1791 316 1792
rect 310 1787 311 1791
rect 315 1787 316 1791
rect 310 1786 316 1787
rect 406 1791 412 1792
rect 406 1787 407 1791
rect 411 1787 412 1791
rect 406 1786 412 1787
rect 526 1791 532 1792
rect 526 1787 527 1791
rect 531 1787 532 1791
rect 526 1786 532 1787
rect 654 1791 660 1792
rect 654 1787 655 1791
rect 659 1787 660 1791
rect 654 1786 660 1787
rect 798 1791 804 1792
rect 798 1787 799 1791
rect 803 1787 804 1791
rect 798 1786 804 1787
rect 942 1791 948 1792
rect 942 1787 943 1791
rect 947 1787 948 1791
rect 942 1786 948 1787
rect 1086 1791 1092 1792
rect 1086 1787 1087 1791
rect 1091 1787 1092 1791
rect 1086 1786 1092 1787
rect 1168 1784 1170 1866
rect 1200 1865 1202 1881
rect 1270 1879 1276 1880
rect 1270 1875 1271 1879
rect 1275 1875 1276 1879
rect 1270 1874 1276 1875
rect 1198 1864 1204 1865
rect 1198 1860 1199 1864
rect 1203 1860 1204 1864
rect 1198 1859 1204 1860
rect 1272 1856 1274 1874
rect 1328 1865 1330 1881
rect 1398 1879 1404 1880
rect 1398 1875 1399 1879
rect 1403 1875 1404 1879
rect 1398 1874 1404 1875
rect 1326 1864 1332 1865
rect 1326 1860 1327 1864
rect 1331 1860 1332 1864
rect 1326 1859 1332 1860
rect 1400 1856 1402 1874
rect 1408 1856 1410 1894
rect 1472 1892 1474 1910
rect 1518 1908 1524 1909
rect 1518 1904 1519 1908
rect 1523 1904 1524 1908
rect 1518 1903 1524 1904
rect 1470 1891 1476 1892
rect 1470 1887 1471 1891
rect 1475 1887 1476 1891
rect 1520 1887 1522 1903
rect 1592 1892 1594 1910
rect 1654 1908 1660 1909
rect 1654 1904 1655 1908
rect 1659 1904 1660 1908
rect 1766 1907 1767 1911
rect 1771 1907 1772 1911
rect 1807 1909 1811 1910
rect 1831 1914 1835 1915
rect 1902 1911 1903 1915
rect 1907 1911 1908 1915
rect 1902 1910 1908 1911
rect 1919 1914 1923 1915
rect 1831 1909 1835 1910
rect 1919 1909 1923 1910
rect 2039 1914 2043 1915
rect 2039 1909 2043 1910
rect 2047 1914 2051 1915
rect 2047 1909 2051 1910
rect 2167 1914 2171 1915
rect 2167 1909 2171 1910
rect 2183 1914 2187 1915
rect 2183 1909 2187 1910
rect 2303 1914 2307 1915
rect 2303 1909 2307 1910
rect 2327 1914 2331 1915
rect 2327 1909 2331 1910
rect 1766 1906 1772 1907
rect 1654 1903 1660 1904
rect 1590 1891 1596 1892
rect 1590 1887 1591 1891
rect 1595 1887 1596 1891
rect 1656 1887 1658 1903
rect 1768 1887 1770 1906
rect 1808 1890 1810 1909
rect 1832 1893 1834 1909
rect 1910 1907 1916 1908
rect 1910 1903 1911 1907
rect 1915 1903 1916 1907
rect 1910 1902 1916 1903
rect 1830 1892 1836 1893
rect 1806 1889 1812 1890
rect 1455 1886 1459 1887
rect 1470 1886 1476 1887
rect 1519 1886 1523 1887
rect 1590 1886 1596 1887
rect 1655 1886 1659 1887
rect 1455 1881 1459 1882
rect 1519 1881 1523 1882
rect 1655 1881 1659 1882
rect 1767 1886 1771 1887
rect 1806 1885 1807 1889
rect 1811 1885 1812 1889
rect 1830 1888 1831 1892
rect 1835 1888 1836 1892
rect 1830 1887 1836 1888
rect 1806 1884 1812 1885
rect 1912 1884 1914 1902
rect 1920 1893 1922 1909
rect 2040 1893 2042 1909
rect 2094 1907 2100 1908
rect 2094 1903 2095 1907
rect 2099 1903 2100 1907
rect 2094 1902 2100 1903
rect 2110 1907 2116 1908
rect 2110 1903 2111 1907
rect 2115 1903 2116 1907
rect 2110 1902 2116 1903
rect 1918 1892 1924 1893
rect 1918 1888 1919 1892
rect 1923 1888 1924 1892
rect 1918 1887 1924 1888
rect 2038 1892 2044 1893
rect 2038 1888 2039 1892
rect 2043 1888 2044 1892
rect 2038 1887 2044 1888
rect 1767 1881 1771 1882
rect 1894 1883 1900 1884
rect 1456 1865 1458 1881
rect 1454 1864 1460 1865
rect 1454 1860 1455 1864
rect 1459 1860 1460 1864
rect 1768 1862 1770 1881
rect 1894 1879 1895 1883
rect 1899 1879 1900 1883
rect 1894 1878 1900 1879
rect 1910 1883 1916 1884
rect 1910 1879 1911 1883
rect 1915 1879 1916 1883
rect 1910 1878 1916 1879
rect 1830 1873 1836 1874
rect 1806 1872 1812 1873
rect 1806 1868 1807 1872
rect 1811 1868 1812 1872
rect 1830 1869 1831 1873
rect 1835 1869 1836 1873
rect 1830 1868 1836 1869
rect 1806 1867 1812 1868
rect 1454 1859 1460 1860
rect 1766 1861 1772 1862
rect 1766 1857 1767 1861
rect 1771 1857 1772 1861
rect 1766 1856 1772 1857
rect 1270 1855 1276 1856
rect 1270 1851 1271 1855
rect 1275 1851 1276 1855
rect 1270 1850 1276 1851
rect 1398 1855 1404 1856
rect 1398 1851 1399 1855
rect 1403 1851 1404 1855
rect 1398 1850 1404 1851
rect 1406 1855 1412 1856
rect 1406 1851 1407 1855
rect 1411 1851 1412 1855
rect 1406 1850 1412 1851
rect 1808 1847 1810 1867
rect 1832 1847 1834 1868
rect 1807 1846 1811 1847
rect 1198 1845 1204 1846
rect 1198 1841 1199 1845
rect 1203 1841 1204 1845
rect 1198 1840 1204 1841
rect 1326 1845 1332 1846
rect 1326 1841 1327 1845
rect 1331 1841 1332 1845
rect 1326 1840 1332 1841
rect 1454 1845 1460 1846
rect 1454 1841 1455 1845
rect 1459 1841 1460 1845
rect 1454 1840 1460 1841
rect 1766 1844 1772 1845
rect 1766 1840 1767 1844
rect 1771 1840 1772 1844
rect 1807 1841 1811 1842
rect 1831 1846 1835 1847
rect 1831 1841 1835 1842
rect 1200 1815 1202 1840
rect 1328 1815 1330 1840
rect 1456 1815 1458 1840
rect 1766 1839 1772 1840
rect 1726 1815 1732 1816
rect 1768 1815 1770 1839
rect 1808 1825 1810 1841
rect 1806 1824 1812 1825
rect 1832 1824 1834 1841
rect 1806 1820 1807 1824
rect 1811 1820 1812 1824
rect 1806 1819 1812 1820
rect 1830 1823 1836 1824
rect 1830 1819 1831 1823
rect 1835 1819 1836 1823
rect 1830 1818 1836 1819
rect 1199 1814 1203 1815
rect 1199 1809 1203 1810
rect 1239 1814 1243 1815
rect 1239 1809 1243 1810
rect 1327 1814 1331 1815
rect 1327 1809 1331 1810
rect 1391 1814 1395 1815
rect 1391 1809 1395 1810
rect 1455 1814 1459 1815
rect 1455 1809 1459 1810
rect 1543 1814 1547 1815
rect 1543 1809 1547 1810
rect 1671 1814 1675 1815
rect 1726 1811 1727 1815
rect 1731 1811 1732 1815
rect 1726 1810 1732 1811
rect 1767 1814 1771 1815
rect 1671 1809 1675 1810
rect 1240 1792 1242 1809
rect 1392 1792 1394 1809
rect 1544 1792 1546 1809
rect 1672 1792 1674 1809
rect 1238 1791 1244 1792
rect 1238 1787 1239 1791
rect 1243 1787 1244 1791
rect 1238 1786 1244 1787
rect 1390 1791 1396 1792
rect 1390 1787 1391 1791
rect 1395 1787 1396 1791
rect 1390 1786 1396 1787
rect 1542 1791 1548 1792
rect 1542 1787 1543 1791
rect 1547 1787 1548 1791
rect 1542 1786 1548 1787
rect 1670 1791 1676 1792
rect 1670 1787 1671 1791
rect 1675 1787 1676 1791
rect 1670 1786 1676 1787
rect 1166 1783 1172 1784
rect 206 1779 212 1780
rect 110 1775 116 1776
rect 110 1771 111 1775
rect 115 1771 116 1775
rect 206 1775 207 1779
rect 211 1775 212 1779
rect 206 1774 212 1775
rect 294 1779 300 1780
rect 294 1775 295 1779
rect 299 1775 300 1779
rect 294 1774 300 1775
rect 382 1779 388 1780
rect 382 1775 383 1779
rect 387 1775 388 1779
rect 382 1774 388 1775
rect 478 1779 484 1780
rect 478 1775 479 1779
rect 483 1775 484 1779
rect 478 1774 484 1775
rect 598 1779 604 1780
rect 598 1775 599 1779
rect 603 1775 604 1779
rect 598 1774 604 1775
rect 726 1779 732 1780
rect 726 1775 727 1779
rect 731 1775 732 1779
rect 726 1774 732 1775
rect 1014 1779 1020 1780
rect 1014 1775 1015 1779
rect 1019 1775 1020 1779
rect 1014 1774 1020 1775
rect 1158 1779 1164 1780
rect 1158 1775 1159 1779
rect 1163 1775 1164 1779
rect 1166 1779 1167 1783
rect 1171 1779 1172 1783
rect 1166 1778 1172 1779
rect 1366 1783 1372 1784
rect 1366 1779 1367 1783
rect 1371 1779 1372 1783
rect 1366 1778 1372 1779
rect 1622 1783 1628 1784
rect 1622 1779 1623 1783
rect 1627 1779 1628 1783
rect 1622 1778 1628 1779
rect 1158 1774 1164 1775
rect 110 1770 116 1771
rect 134 1772 140 1773
rect 112 1739 114 1770
rect 134 1768 135 1772
rect 139 1768 140 1772
rect 134 1767 140 1768
rect 136 1739 138 1767
rect 208 1756 210 1774
rect 222 1772 228 1773
rect 222 1768 223 1772
rect 227 1768 228 1772
rect 222 1767 228 1768
rect 198 1755 204 1756
rect 198 1751 199 1755
rect 203 1751 204 1755
rect 198 1750 204 1751
rect 206 1755 212 1756
rect 206 1751 207 1755
rect 211 1751 212 1755
rect 206 1750 212 1751
rect 111 1738 115 1739
rect 111 1733 115 1734
rect 135 1738 139 1739
rect 135 1733 139 1734
rect 112 1714 114 1733
rect 136 1717 138 1733
rect 134 1716 140 1717
rect 110 1713 116 1714
rect 110 1709 111 1713
rect 115 1709 116 1713
rect 134 1712 135 1716
rect 139 1712 140 1716
rect 134 1711 140 1712
rect 110 1708 116 1709
rect 200 1708 202 1750
rect 224 1739 226 1767
rect 296 1756 298 1774
rect 310 1772 316 1773
rect 310 1768 311 1772
rect 315 1768 316 1772
rect 310 1767 316 1768
rect 294 1755 300 1756
rect 294 1751 295 1755
rect 299 1751 300 1755
rect 294 1750 300 1751
rect 312 1739 314 1767
rect 384 1756 386 1774
rect 406 1772 412 1773
rect 406 1768 407 1772
rect 411 1768 412 1772
rect 406 1767 412 1768
rect 382 1755 388 1756
rect 382 1751 383 1755
rect 387 1751 388 1755
rect 382 1750 388 1751
rect 408 1739 410 1767
rect 480 1756 482 1774
rect 526 1772 532 1773
rect 526 1768 527 1772
rect 531 1768 532 1772
rect 526 1767 532 1768
rect 478 1755 484 1756
rect 478 1751 479 1755
rect 483 1751 484 1755
rect 478 1750 484 1751
rect 528 1739 530 1767
rect 600 1756 602 1774
rect 654 1772 660 1773
rect 654 1768 655 1772
rect 659 1768 660 1772
rect 654 1767 660 1768
rect 598 1755 604 1756
rect 598 1751 599 1755
rect 603 1751 604 1755
rect 598 1750 604 1751
rect 656 1739 658 1767
rect 728 1756 730 1774
rect 798 1772 804 1773
rect 798 1768 799 1772
rect 803 1768 804 1772
rect 798 1767 804 1768
rect 942 1772 948 1773
rect 942 1768 943 1772
rect 947 1768 948 1772
rect 942 1767 948 1768
rect 726 1755 732 1756
rect 726 1751 727 1755
rect 731 1751 732 1755
rect 726 1750 732 1751
rect 800 1739 802 1767
rect 944 1739 946 1767
rect 1016 1756 1018 1774
rect 1086 1772 1092 1773
rect 1086 1768 1087 1772
rect 1091 1768 1092 1772
rect 1086 1767 1092 1768
rect 998 1755 1004 1756
rect 998 1751 999 1755
rect 1003 1751 1004 1755
rect 998 1750 1004 1751
rect 1014 1755 1020 1756
rect 1014 1751 1015 1755
rect 1019 1751 1020 1755
rect 1014 1750 1020 1751
rect 223 1738 227 1739
rect 223 1733 227 1734
rect 247 1738 251 1739
rect 247 1733 251 1734
rect 311 1738 315 1739
rect 311 1733 315 1734
rect 399 1738 403 1739
rect 399 1733 403 1734
rect 407 1738 411 1739
rect 407 1733 411 1734
rect 527 1738 531 1739
rect 527 1733 531 1734
rect 567 1738 571 1739
rect 567 1733 571 1734
rect 655 1738 659 1739
rect 655 1733 659 1734
rect 751 1738 755 1739
rect 751 1733 755 1734
rect 799 1738 803 1739
rect 799 1733 803 1734
rect 935 1738 939 1739
rect 935 1733 939 1734
rect 943 1738 947 1739
rect 943 1733 947 1734
rect 214 1731 220 1732
rect 214 1727 215 1731
rect 219 1727 220 1731
rect 214 1726 220 1727
rect 216 1708 218 1726
rect 248 1717 250 1733
rect 326 1731 332 1732
rect 326 1727 327 1731
rect 331 1727 332 1731
rect 326 1726 332 1727
rect 246 1716 252 1717
rect 246 1712 247 1716
rect 251 1712 252 1716
rect 246 1711 252 1712
rect 328 1708 330 1726
rect 400 1717 402 1733
rect 478 1731 484 1732
rect 478 1727 479 1731
rect 483 1727 484 1731
rect 478 1726 484 1727
rect 398 1716 404 1717
rect 398 1712 399 1716
rect 403 1712 404 1716
rect 398 1711 404 1712
rect 198 1707 204 1708
rect 198 1703 199 1707
rect 203 1703 204 1707
rect 198 1702 204 1703
rect 214 1707 220 1708
rect 214 1703 215 1707
rect 219 1703 220 1707
rect 214 1702 220 1703
rect 326 1707 332 1708
rect 326 1703 327 1707
rect 331 1703 332 1707
rect 326 1702 332 1703
rect 134 1697 140 1698
rect 110 1696 116 1697
rect 110 1692 111 1696
rect 115 1692 116 1696
rect 134 1693 135 1697
rect 139 1693 140 1697
rect 134 1692 140 1693
rect 246 1697 252 1698
rect 246 1693 247 1697
rect 251 1693 252 1697
rect 246 1692 252 1693
rect 398 1697 404 1698
rect 398 1693 399 1697
rect 403 1693 404 1697
rect 398 1692 404 1693
rect 110 1691 116 1692
rect 112 1671 114 1691
rect 136 1671 138 1692
rect 248 1671 250 1692
rect 400 1671 402 1692
rect 111 1670 115 1671
rect 111 1665 115 1666
rect 135 1670 139 1671
rect 135 1665 139 1666
rect 191 1670 195 1671
rect 191 1665 195 1666
rect 247 1670 251 1671
rect 247 1665 251 1666
rect 295 1670 299 1671
rect 295 1665 299 1666
rect 399 1670 403 1671
rect 399 1665 403 1666
rect 407 1670 411 1671
rect 407 1665 411 1666
rect 112 1649 114 1665
rect 110 1648 116 1649
rect 192 1648 194 1665
rect 296 1648 298 1665
rect 408 1648 410 1665
rect 110 1644 111 1648
rect 115 1644 116 1648
rect 110 1643 116 1644
rect 190 1647 196 1648
rect 190 1643 191 1647
rect 195 1643 196 1647
rect 190 1642 196 1643
rect 294 1647 300 1648
rect 294 1643 295 1647
rect 299 1643 300 1647
rect 294 1642 300 1643
rect 406 1647 412 1648
rect 406 1643 407 1647
rect 411 1643 412 1647
rect 406 1642 412 1643
rect 480 1640 482 1726
rect 568 1717 570 1733
rect 734 1731 740 1732
rect 734 1727 735 1731
rect 739 1727 740 1731
rect 734 1726 740 1727
rect 566 1716 572 1717
rect 566 1712 567 1716
rect 571 1712 572 1716
rect 566 1711 572 1712
rect 736 1708 738 1726
rect 752 1717 754 1733
rect 936 1717 938 1733
rect 750 1716 756 1717
rect 750 1712 751 1716
rect 755 1712 756 1716
rect 750 1711 756 1712
rect 934 1716 940 1717
rect 934 1712 935 1716
rect 939 1712 940 1716
rect 934 1711 940 1712
rect 1000 1708 1002 1750
rect 1088 1739 1090 1767
rect 1160 1756 1162 1774
rect 1238 1772 1244 1773
rect 1238 1768 1239 1772
rect 1243 1768 1244 1772
rect 1238 1767 1244 1768
rect 1158 1755 1164 1756
rect 1158 1751 1159 1755
rect 1163 1751 1164 1755
rect 1158 1750 1164 1751
rect 1240 1739 1242 1767
rect 1087 1738 1091 1739
rect 1087 1733 1091 1734
rect 1119 1738 1123 1739
rect 1119 1733 1123 1734
rect 1239 1738 1243 1739
rect 1239 1733 1243 1734
rect 1311 1738 1315 1739
rect 1311 1733 1315 1734
rect 1014 1731 1020 1732
rect 1014 1727 1015 1731
rect 1019 1727 1020 1731
rect 1014 1726 1020 1727
rect 1016 1708 1018 1726
rect 1120 1717 1122 1733
rect 1174 1731 1180 1732
rect 1174 1727 1175 1731
rect 1179 1727 1180 1731
rect 1174 1726 1180 1727
rect 1118 1716 1124 1717
rect 1118 1712 1119 1716
rect 1123 1712 1124 1716
rect 1118 1711 1124 1712
rect 722 1707 728 1708
rect 722 1703 723 1707
rect 727 1703 728 1707
rect 722 1702 728 1703
rect 734 1707 740 1708
rect 734 1703 735 1707
rect 739 1703 740 1707
rect 734 1702 740 1703
rect 998 1707 1004 1708
rect 998 1703 999 1707
rect 1003 1703 1004 1707
rect 998 1702 1004 1703
rect 1014 1707 1020 1708
rect 1014 1703 1015 1707
rect 1019 1703 1020 1707
rect 1014 1702 1020 1703
rect 566 1697 572 1698
rect 566 1693 567 1697
rect 571 1693 572 1697
rect 566 1692 572 1693
rect 568 1671 570 1692
rect 535 1670 539 1671
rect 535 1665 539 1666
rect 567 1670 571 1671
rect 567 1665 571 1666
rect 687 1670 691 1671
rect 687 1665 691 1666
rect 536 1648 538 1665
rect 688 1648 690 1665
rect 534 1647 540 1648
rect 534 1643 535 1647
rect 539 1643 540 1647
rect 534 1642 540 1643
rect 686 1647 692 1648
rect 686 1643 687 1647
rect 691 1643 692 1647
rect 686 1642 692 1643
rect 478 1639 484 1640
rect 262 1635 268 1636
rect 110 1631 116 1632
rect 110 1627 111 1631
rect 115 1627 116 1631
rect 262 1631 263 1635
rect 267 1631 268 1635
rect 262 1630 268 1631
rect 366 1635 372 1636
rect 366 1631 367 1635
rect 371 1631 372 1635
rect 478 1635 479 1639
rect 483 1635 484 1639
rect 614 1639 620 1640
rect 478 1634 484 1635
rect 606 1635 612 1636
rect 366 1630 372 1631
rect 606 1631 607 1635
rect 611 1631 612 1635
rect 614 1635 615 1639
rect 619 1635 620 1639
rect 614 1634 620 1635
rect 606 1630 612 1631
rect 110 1626 116 1627
rect 190 1628 196 1629
rect 112 1603 114 1626
rect 190 1624 191 1628
rect 195 1624 196 1628
rect 190 1623 196 1624
rect 192 1603 194 1623
rect 264 1612 266 1630
rect 294 1628 300 1629
rect 294 1624 295 1628
rect 299 1624 300 1628
rect 294 1623 300 1624
rect 246 1611 252 1612
rect 246 1607 247 1611
rect 251 1607 252 1611
rect 246 1606 252 1607
rect 262 1611 268 1612
rect 262 1607 263 1611
rect 267 1607 268 1611
rect 262 1606 268 1607
rect 111 1602 115 1603
rect 111 1597 115 1598
rect 191 1602 195 1603
rect 191 1597 195 1598
rect 112 1578 114 1597
rect 110 1577 116 1578
rect 110 1573 111 1577
rect 115 1573 116 1577
rect 110 1572 116 1573
rect 248 1572 250 1606
rect 296 1603 298 1623
rect 368 1612 370 1630
rect 406 1628 412 1629
rect 406 1624 407 1628
rect 411 1624 412 1628
rect 406 1623 412 1624
rect 534 1628 540 1629
rect 534 1624 535 1628
rect 539 1624 540 1628
rect 534 1623 540 1624
rect 366 1611 372 1612
rect 366 1607 367 1611
rect 371 1607 372 1611
rect 366 1606 372 1607
rect 408 1603 410 1623
rect 536 1603 538 1623
rect 295 1602 299 1603
rect 295 1597 299 1598
rect 327 1602 331 1603
rect 327 1597 331 1598
rect 407 1602 411 1603
rect 407 1597 411 1598
rect 431 1602 435 1603
rect 431 1597 435 1598
rect 535 1602 539 1603
rect 535 1597 539 1598
rect 543 1602 547 1603
rect 543 1597 547 1598
rect 328 1581 330 1597
rect 432 1581 434 1597
rect 462 1595 468 1596
rect 462 1591 463 1595
rect 467 1591 468 1595
rect 462 1590 468 1591
rect 326 1580 332 1581
rect 326 1576 327 1580
rect 331 1576 332 1580
rect 326 1575 332 1576
rect 430 1580 436 1581
rect 430 1576 431 1580
rect 435 1576 436 1580
rect 430 1575 436 1576
rect 246 1571 252 1572
rect 246 1567 247 1571
rect 251 1567 252 1571
rect 246 1566 252 1567
rect 326 1561 332 1562
rect 110 1560 116 1561
rect 110 1556 111 1560
rect 115 1556 116 1560
rect 326 1557 327 1561
rect 331 1557 332 1561
rect 326 1556 332 1557
rect 430 1561 436 1562
rect 430 1557 431 1561
rect 435 1557 436 1561
rect 430 1556 436 1557
rect 110 1555 116 1556
rect 112 1535 114 1555
rect 328 1535 330 1556
rect 432 1535 434 1556
rect 111 1534 115 1535
rect 111 1529 115 1530
rect 223 1534 227 1535
rect 223 1529 227 1530
rect 327 1534 331 1535
rect 327 1529 331 1530
rect 343 1534 347 1535
rect 343 1529 347 1530
rect 431 1534 435 1535
rect 431 1529 435 1530
rect 112 1513 114 1529
rect 110 1512 116 1513
rect 224 1512 226 1529
rect 344 1512 346 1529
rect 110 1508 111 1512
rect 115 1508 116 1512
rect 110 1507 116 1508
rect 222 1511 228 1512
rect 222 1507 223 1511
rect 227 1507 228 1511
rect 222 1506 228 1507
rect 342 1511 348 1512
rect 342 1507 343 1511
rect 347 1507 348 1511
rect 342 1506 348 1507
rect 464 1504 466 1590
rect 544 1581 546 1597
rect 608 1596 610 1630
rect 616 1612 618 1634
rect 686 1628 692 1629
rect 686 1624 687 1628
rect 691 1624 692 1628
rect 686 1623 692 1624
rect 614 1611 620 1612
rect 614 1607 615 1611
rect 619 1607 620 1611
rect 614 1606 620 1607
rect 688 1603 690 1623
rect 724 1612 726 1702
rect 750 1697 756 1698
rect 750 1693 751 1697
rect 755 1693 756 1697
rect 750 1692 756 1693
rect 934 1697 940 1698
rect 934 1693 935 1697
rect 939 1693 940 1697
rect 934 1692 940 1693
rect 1118 1697 1124 1698
rect 1118 1693 1119 1697
rect 1123 1693 1124 1697
rect 1118 1692 1124 1693
rect 752 1671 754 1692
rect 936 1671 938 1692
rect 1120 1671 1122 1692
rect 751 1670 755 1671
rect 751 1665 755 1666
rect 855 1670 859 1671
rect 855 1665 859 1666
rect 935 1670 939 1671
rect 935 1665 939 1666
rect 1039 1670 1043 1671
rect 1039 1665 1043 1666
rect 1119 1670 1123 1671
rect 1119 1665 1123 1666
rect 856 1648 858 1665
rect 1040 1648 1042 1665
rect 854 1647 860 1648
rect 854 1643 855 1647
rect 859 1643 860 1647
rect 854 1642 860 1643
rect 1038 1647 1044 1648
rect 1038 1643 1039 1647
rect 1043 1643 1044 1647
rect 1038 1642 1044 1643
rect 1176 1640 1178 1726
rect 1312 1717 1314 1733
rect 1368 1732 1370 1778
rect 1390 1772 1396 1773
rect 1390 1768 1391 1772
rect 1395 1768 1396 1772
rect 1390 1767 1396 1768
rect 1542 1772 1548 1773
rect 1542 1768 1543 1772
rect 1547 1768 1548 1772
rect 1542 1767 1548 1768
rect 1392 1739 1394 1767
rect 1544 1739 1546 1767
rect 1624 1756 1626 1778
rect 1670 1772 1676 1773
rect 1670 1768 1671 1772
rect 1675 1768 1676 1772
rect 1670 1767 1676 1768
rect 1622 1755 1628 1756
rect 1622 1751 1623 1755
rect 1627 1751 1628 1755
rect 1622 1750 1628 1751
rect 1672 1739 1674 1767
rect 1728 1756 1730 1810
rect 1767 1809 1771 1810
rect 1768 1793 1770 1809
rect 1806 1807 1812 1808
rect 1806 1803 1807 1807
rect 1811 1803 1812 1807
rect 1806 1802 1812 1803
rect 1830 1804 1836 1805
rect 1766 1792 1772 1793
rect 1766 1788 1767 1792
rect 1771 1788 1772 1792
rect 1766 1787 1772 1788
rect 1766 1775 1772 1776
rect 1766 1771 1767 1775
rect 1771 1771 1772 1775
rect 1808 1771 1810 1802
rect 1830 1800 1831 1804
rect 1835 1800 1836 1804
rect 1830 1799 1836 1800
rect 1832 1771 1834 1799
rect 1896 1788 1898 1878
rect 1918 1873 1924 1874
rect 1918 1869 1919 1873
rect 1923 1869 1924 1873
rect 1918 1868 1924 1869
rect 2038 1873 2044 1874
rect 2038 1869 2039 1873
rect 2043 1869 2044 1873
rect 2038 1868 2044 1869
rect 1920 1847 1922 1868
rect 2040 1847 2042 1868
rect 1919 1846 1923 1847
rect 1919 1841 1923 1842
rect 1959 1846 1963 1847
rect 1959 1841 1963 1842
rect 2039 1846 2043 1847
rect 2039 1841 2043 1842
rect 1960 1824 1962 1841
rect 1958 1823 1964 1824
rect 1958 1819 1959 1823
rect 1963 1819 1964 1823
rect 1958 1818 1964 1819
rect 2096 1816 2098 1902
rect 2112 1884 2114 1902
rect 2168 1893 2170 1909
rect 2238 1907 2244 1908
rect 2238 1903 2239 1907
rect 2243 1903 2244 1907
rect 2238 1902 2244 1903
rect 2166 1892 2172 1893
rect 2166 1888 2167 1892
rect 2171 1888 2172 1892
rect 2166 1887 2172 1888
rect 2240 1884 2242 1902
rect 2304 1893 2306 1909
rect 2302 1892 2308 1893
rect 2302 1888 2303 1892
rect 2307 1888 2308 1892
rect 2302 1887 2308 1888
rect 2376 1884 2378 1918
rect 2472 1915 2474 1935
rect 2528 1924 2530 2026
rect 2574 2021 2580 2022
rect 2574 2017 2575 2021
rect 2579 2017 2580 2021
rect 2574 2016 2580 2017
rect 2726 2021 2732 2022
rect 2726 2017 2727 2021
rect 2731 2017 2732 2021
rect 2726 2016 2732 2017
rect 2870 2021 2876 2022
rect 2870 2017 2871 2021
rect 2875 2017 2876 2021
rect 2870 2016 2876 2017
rect 3006 2021 3012 2022
rect 3006 2017 3007 2021
rect 3011 2017 3012 2021
rect 3006 2016 3012 2017
rect 2576 1983 2578 2016
rect 2728 1983 2730 2016
rect 2872 1983 2874 2016
rect 3008 1983 3010 2016
rect 2575 1982 2579 1983
rect 2575 1977 2579 1978
rect 2615 1982 2619 1983
rect 2615 1977 2619 1978
rect 2727 1982 2731 1983
rect 2727 1977 2731 1978
rect 2751 1982 2755 1983
rect 2751 1977 2755 1978
rect 2871 1982 2875 1983
rect 2871 1977 2875 1978
rect 2887 1982 2891 1983
rect 2887 1977 2891 1978
rect 3007 1982 3011 1983
rect 3007 1977 3011 1978
rect 3031 1982 3035 1983
rect 3031 1977 3035 1978
rect 2616 1960 2618 1977
rect 2752 1960 2754 1977
rect 2888 1960 2890 1977
rect 3032 1960 3034 1977
rect 2614 1959 2620 1960
rect 2614 1955 2615 1959
rect 2619 1955 2620 1959
rect 2614 1954 2620 1955
rect 2750 1959 2756 1960
rect 2750 1955 2751 1959
rect 2755 1955 2756 1959
rect 2750 1954 2756 1955
rect 2886 1959 2892 1960
rect 2886 1955 2887 1959
rect 2891 1955 2892 1959
rect 2886 1954 2892 1955
rect 3030 1959 3036 1960
rect 3030 1955 3031 1959
rect 3035 1955 3036 1959
rect 3030 1954 3036 1955
rect 3112 1952 3114 2042
rect 3136 2041 3138 2057
rect 3206 2055 3212 2056
rect 3206 2051 3207 2055
rect 3211 2051 3212 2055
rect 3206 2050 3212 2051
rect 3134 2040 3140 2041
rect 3134 2036 3135 2040
rect 3139 2036 3140 2040
rect 3134 2035 3140 2036
rect 3208 2032 3210 2050
rect 3264 2041 3266 2057
rect 3262 2040 3268 2041
rect 3262 2036 3263 2040
rect 3267 2036 3268 2040
rect 3262 2035 3268 2036
rect 3328 2032 3330 2070
rect 3206 2031 3212 2032
rect 3206 2027 3207 2031
rect 3211 2027 3212 2031
rect 3206 2026 3212 2027
rect 3326 2031 3332 2032
rect 3326 2027 3327 2031
rect 3331 2027 3332 2031
rect 3326 2026 3332 2027
rect 3134 2021 3140 2022
rect 3134 2017 3135 2021
rect 3139 2017 3140 2021
rect 3134 2016 3140 2017
rect 3262 2021 3268 2022
rect 3262 2017 3263 2021
rect 3267 2017 3268 2021
rect 3262 2016 3268 2017
rect 3136 1983 3138 2016
rect 3264 1983 3266 2016
rect 3135 1982 3139 1983
rect 3135 1977 3139 1978
rect 3175 1982 3179 1983
rect 3175 1977 3179 1978
rect 3263 1982 3267 1983
rect 3263 1977 3267 1978
rect 3319 1982 3323 1983
rect 3319 1977 3323 1978
rect 3176 1960 3178 1977
rect 3320 1960 3322 1977
rect 3174 1959 3180 1960
rect 3174 1955 3175 1959
rect 3179 1955 3180 1959
rect 3174 1954 3180 1955
rect 3318 1959 3324 1960
rect 3318 1955 3319 1959
rect 3323 1955 3324 1959
rect 3318 1954 3324 1955
rect 3110 1951 3116 1952
rect 2542 1947 2548 1948
rect 2542 1943 2543 1947
rect 2547 1943 2548 1947
rect 2542 1942 2548 1943
rect 2686 1947 2692 1948
rect 2686 1943 2687 1947
rect 2691 1943 2692 1947
rect 2686 1942 2692 1943
rect 2822 1947 2828 1948
rect 2822 1943 2823 1947
rect 2827 1943 2828 1947
rect 2822 1942 2828 1943
rect 2958 1947 2964 1948
rect 2958 1943 2959 1947
rect 2963 1943 2964 1947
rect 2958 1942 2964 1943
rect 3102 1947 3108 1948
rect 3102 1943 3103 1947
rect 3107 1943 3108 1947
rect 3110 1947 3111 1951
rect 3115 1947 3116 1951
rect 3110 1946 3116 1947
rect 3102 1942 3108 1943
rect 2526 1923 2532 1924
rect 2526 1919 2527 1923
rect 2531 1919 2532 1923
rect 2526 1918 2532 1919
rect 2455 1914 2459 1915
rect 2455 1909 2459 1910
rect 2471 1914 2475 1915
rect 2471 1909 2475 1910
rect 2456 1893 2458 1909
rect 2544 1908 2546 1942
rect 2614 1940 2620 1941
rect 2614 1936 2615 1940
rect 2619 1936 2620 1940
rect 2614 1935 2620 1936
rect 2616 1915 2618 1935
rect 2688 1924 2690 1942
rect 2750 1940 2756 1941
rect 2750 1936 2751 1940
rect 2755 1936 2756 1940
rect 2750 1935 2756 1936
rect 2686 1923 2692 1924
rect 2686 1919 2687 1923
rect 2691 1919 2692 1923
rect 2686 1918 2692 1919
rect 2752 1915 2754 1935
rect 2824 1924 2826 1942
rect 2886 1940 2892 1941
rect 2886 1936 2887 1940
rect 2891 1936 2892 1940
rect 2886 1935 2892 1936
rect 2822 1923 2828 1924
rect 2822 1919 2823 1923
rect 2827 1919 2828 1923
rect 2822 1918 2828 1919
rect 2888 1915 2890 1935
rect 2960 1924 2962 1942
rect 3030 1940 3036 1941
rect 3030 1936 3031 1940
rect 3035 1936 3036 1940
rect 3030 1935 3036 1936
rect 2958 1923 2964 1924
rect 2958 1919 2959 1923
rect 2963 1919 2964 1923
rect 2958 1918 2964 1919
rect 3032 1915 3034 1935
rect 3104 1924 3106 1942
rect 3174 1940 3180 1941
rect 3174 1936 3175 1940
rect 3179 1936 3180 1940
rect 3174 1935 3180 1936
rect 3318 1940 3324 1941
rect 3318 1936 3319 1940
rect 3323 1936 3324 1940
rect 3318 1935 3324 1936
rect 3102 1923 3108 1924
rect 3102 1919 3103 1923
rect 3107 1919 3108 1923
rect 3102 1918 3108 1919
rect 3166 1915 3172 1916
rect 3176 1915 3178 1935
rect 3320 1915 3322 1935
rect 3360 1924 3362 2098
rect 3366 2092 3372 2093
rect 3366 2088 3367 2092
rect 3371 2088 3372 2092
rect 3366 2087 3372 2088
rect 3368 2063 3370 2087
rect 3367 2062 3371 2063
rect 3367 2057 3371 2058
rect 3368 2041 3370 2057
rect 3430 2055 3436 2056
rect 3430 2051 3431 2055
rect 3435 2051 3436 2055
rect 3430 2050 3436 2051
rect 3366 2040 3372 2041
rect 3366 2036 3367 2040
rect 3371 2036 3372 2040
rect 3366 2035 3372 2036
rect 3366 2021 3372 2022
rect 3366 2017 3367 2021
rect 3371 2017 3372 2021
rect 3366 2016 3372 2017
rect 3368 1983 3370 2016
rect 3367 1982 3371 1983
rect 3367 1977 3371 1978
rect 3390 1947 3396 1948
rect 3390 1943 3391 1947
rect 3395 1943 3396 1947
rect 3390 1942 3396 1943
rect 3358 1923 3364 1924
rect 3358 1919 3359 1923
rect 3363 1919 3364 1923
rect 3358 1918 3364 1919
rect 2615 1914 2619 1915
rect 2615 1909 2619 1910
rect 2751 1914 2755 1915
rect 2751 1909 2755 1910
rect 2791 1914 2795 1915
rect 2791 1909 2795 1910
rect 2887 1914 2891 1915
rect 2887 1909 2891 1910
rect 2983 1914 2987 1915
rect 2983 1909 2987 1910
rect 3031 1914 3035 1915
rect 3166 1911 3167 1915
rect 3171 1911 3172 1915
rect 3166 1910 3172 1911
rect 3175 1914 3179 1915
rect 3031 1909 3035 1910
rect 2542 1907 2548 1908
rect 2542 1903 2543 1907
rect 2547 1903 2548 1907
rect 2542 1902 2548 1903
rect 2616 1893 2618 1909
rect 2686 1907 2692 1908
rect 2686 1903 2687 1907
rect 2691 1903 2692 1907
rect 2686 1902 2692 1903
rect 2454 1892 2460 1893
rect 2454 1888 2455 1892
rect 2459 1888 2460 1892
rect 2454 1887 2460 1888
rect 2614 1892 2620 1893
rect 2614 1888 2615 1892
rect 2619 1888 2620 1892
rect 2614 1887 2620 1888
rect 2688 1884 2690 1902
rect 2792 1893 2794 1909
rect 2862 1907 2868 1908
rect 2862 1903 2863 1907
rect 2867 1903 2868 1907
rect 2862 1902 2868 1903
rect 2790 1892 2796 1893
rect 2790 1888 2791 1892
rect 2795 1888 2796 1892
rect 2790 1887 2796 1888
rect 2864 1884 2866 1902
rect 2984 1893 2986 1909
rect 3054 1907 3060 1908
rect 3054 1903 3055 1907
rect 3059 1903 3060 1907
rect 3054 1902 3060 1903
rect 2982 1892 2988 1893
rect 2982 1888 2983 1892
rect 2987 1888 2988 1892
rect 2982 1887 2988 1888
rect 3056 1884 3058 1902
rect 3078 1899 3084 1900
rect 3078 1895 3079 1899
rect 3083 1895 3084 1899
rect 3078 1894 3084 1895
rect 2110 1883 2116 1884
rect 2110 1879 2111 1883
rect 2115 1879 2116 1883
rect 2110 1878 2116 1879
rect 2238 1883 2244 1884
rect 2238 1879 2239 1883
rect 2243 1879 2244 1883
rect 2238 1878 2244 1879
rect 2374 1883 2380 1884
rect 2374 1879 2375 1883
rect 2379 1879 2380 1883
rect 2374 1878 2380 1879
rect 2426 1883 2432 1884
rect 2426 1879 2427 1883
rect 2431 1879 2432 1883
rect 2426 1878 2432 1879
rect 2686 1883 2692 1884
rect 2686 1879 2687 1883
rect 2691 1879 2692 1883
rect 2686 1878 2692 1879
rect 2862 1883 2868 1884
rect 2862 1879 2863 1883
rect 2867 1879 2868 1883
rect 2862 1878 2868 1879
rect 3054 1883 3060 1884
rect 3054 1879 3055 1883
rect 3059 1879 3060 1883
rect 3054 1878 3060 1879
rect 2166 1873 2172 1874
rect 2166 1869 2167 1873
rect 2171 1869 2172 1873
rect 2166 1868 2172 1869
rect 2302 1873 2308 1874
rect 2302 1869 2303 1873
rect 2307 1869 2308 1873
rect 2302 1868 2308 1869
rect 2168 1847 2170 1868
rect 2304 1847 2306 1868
rect 2111 1846 2115 1847
rect 2111 1841 2115 1842
rect 2167 1846 2171 1847
rect 2167 1841 2171 1842
rect 2255 1846 2259 1847
rect 2255 1841 2259 1842
rect 2303 1846 2307 1847
rect 2303 1841 2307 1842
rect 2407 1846 2411 1847
rect 2407 1841 2411 1842
rect 2112 1824 2114 1841
rect 2256 1824 2258 1841
rect 2408 1824 2410 1841
rect 2110 1823 2116 1824
rect 2110 1819 2111 1823
rect 2115 1819 2116 1823
rect 2110 1818 2116 1819
rect 2254 1823 2260 1824
rect 2254 1819 2255 1823
rect 2259 1819 2260 1823
rect 2254 1818 2260 1819
rect 2406 1823 2412 1824
rect 2406 1819 2407 1823
rect 2411 1819 2412 1823
rect 2406 1818 2412 1819
rect 2094 1815 2100 1816
rect 2030 1811 2036 1812
rect 2030 1807 2031 1811
rect 2035 1807 2036 1811
rect 2094 1811 2095 1815
rect 2099 1811 2100 1815
rect 2094 1810 2100 1811
rect 2326 1811 2332 1812
rect 2030 1806 2036 1807
rect 2326 1807 2327 1811
rect 2331 1807 2332 1811
rect 2326 1806 2332 1807
rect 1958 1804 1964 1805
rect 1958 1800 1959 1804
rect 1963 1800 1964 1804
rect 1958 1799 1964 1800
rect 1894 1787 1900 1788
rect 1894 1783 1895 1787
rect 1899 1783 1900 1787
rect 1894 1782 1900 1783
rect 1950 1787 1956 1788
rect 1950 1783 1951 1787
rect 1955 1783 1956 1787
rect 1950 1782 1956 1783
rect 1766 1770 1772 1771
rect 1807 1770 1811 1771
rect 1726 1755 1732 1756
rect 1726 1751 1727 1755
rect 1731 1751 1732 1755
rect 1726 1750 1732 1751
rect 1768 1739 1770 1770
rect 1807 1765 1811 1766
rect 1831 1770 1835 1771
rect 1831 1765 1835 1766
rect 1879 1770 1883 1771
rect 1879 1765 1883 1766
rect 1808 1746 1810 1765
rect 1880 1749 1882 1765
rect 1878 1748 1884 1749
rect 1806 1745 1812 1746
rect 1806 1741 1807 1745
rect 1811 1741 1812 1745
rect 1878 1744 1879 1748
rect 1883 1744 1884 1748
rect 1878 1743 1884 1744
rect 1806 1740 1812 1741
rect 1952 1740 1954 1782
rect 1960 1771 1962 1799
rect 2032 1788 2034 1806
rect 2110 1804 2116 1805
rect 2110 1800 2111 1804
rect 2115 1800 2116 1804
rect 2110 1799 2116 1800
rect 2254 1804 2260 1805
rect 2254 1800 2255 1804
rect 2259 1800 2260 1804
rect 2254 1799 2260 1800
rect 2030 1787 2036 1788
rect 2030 1783 2031 1787
rect 2035 1783 2036 1787
rect 2030 1782 2036 1783
rect 2112 1771 2114 1799
rect 2256 1771 2258 1799
rect 1959 1770 1963 1771
rect 1959 1765 1963 1766
rect 2015 1770 2019 1771
rect 2015 1765 2019 1766
rect 2111 1770 2115 1771
rect 2111 1765 2115 1766
rect 2151 1770 2155 1771
rect 2151 1765 2155 1766
rect 2255 1770 2259 1771
rect 2255 1765 2259 1766
rect 2303 1770 2307 1771
rect 2303 1765 2307 1766
rect 2016 1749 2018 1765
rect 2094 1763 2100 1764
rect 2094 1759 2095 1763
rect 2099 1759 2100 1763
rect 2094 1758 2100 1759
rect 2014 1748 2020 1749
rect 2014 1744 2015 1748
rect 2019 1744 2020 1748
rect 2014 1743 2020 1744
rect 2096 1740 2098 1758
rect 2152 1749 2154 1765
rect 2254 1759 2260 1760
rect 2254 1755 2255 1759
rect 2259 1755 2260 1759
rect 2254 1754 2260 1755
rect 2150 1748 2156 1749
rect 2150 1744 2151 1748
rect 2155 1744 2156 1748
rect 2150 1743 2156 1744
rect 1950 1739 1956 1740
rect 1391 1738 1395 1739
rect 1391 1733 1395 1734
rect 1503 1738 1507 1739
rect 1503 1733 1507 1734
rect 1543 1738 1547 1739
rect 1543 1733 1547 1734
rect 1671 1738 1675 1739
rect 1671 1733 1675 1734
rect 1767 1738 1771 1739
rect 1950 1735 1951 1739
rect 1955 1735 1956 1739
rect 1950 1734 1956 1735
rect 2094 1739 2100 1740
rect 2094 1735 2095 1739
rect 2099 1735 2100 1739
rect 2094 1734 2100 1735
rect 1767 1733 1771 1734
rect 1366 1731 1372 1732
rect 1366 1727 1367 1731
rect 1371 1727 1372 1731
rect 1366 1726 1372 1727
rect 1382 1731 1388 1732
rect 1382 1727 1383 1731
rect 1387 1727 1388 1731
rect 1382 1726 1388 1727
rect 1310 1716 1316 1717
rect 1310 1712 1311 1716
rect 1315 1712 1316 1716
rect 1310 1711 1316 1712
rect 1384 1708 1386 1726
rect 1504 1717 1506 1733
rect 1574 1731 1580 1732
rect 1574 1727 1575 1731
rect 1579 1727 1580 1731
rect 1574 1726 1580 1727
rect 1502 1716 1508 1717
rect 1502 1712 1503 1716
rect 1507 1712 1508 1716
rect 1502 1711 1508 1712
rect 1576 1708 1578 1726
rect 1672 1717 1674 1733
rect 1670 1716 1676 1717
rect 1670 1712 1671 1716
rect 1675 1712 1676 1716
rect 1768 1714 1770 1733
rect 1878 1729 1884 1730
rect 1806 1728 1812 1729
rect 1806 1724 1807 1728
rect 1811 1724 1812 1728
rect 1878 1725 1879 1729
rect 1883 1725 1884 1729
rect 1878 1724 1884 1725
rect 2014 1729 2020 1730
rect 2014 1725 2015 1729
rect 2019 1725 2020 1729
rect 2014 1724 2020 1725
rect 2150 1729 2156 1730
rect 2150 1725 2151 1729
rect 2155 1725 2156 1729
rect 2150 1724 2156 1725
rect 1806 1723 1812 1724
rect 1670 1711 1676 1712
rect 1766 1713 1772 1714
rect 1766 1709 1767 1713
rect 1771 1709 1772 1713
rect 1766 1708 1772 1709
rect 1382 1707 1388 1708
rect 1382 1703 1383 1707
rect 1387 1703 1388 1707
rect 1382 1702 1388 1703
rect 1574 1707 1580 1708
rect 1574 1703 1575 1707
rect 1579 1703 1580 1707
rect 1574 1702 1580 1703
rect 1734 1707 1740 1708
rect 1734 1703 1735 1707
rect 1739 1703 1740 1707
rect 1734 1702 1740 1703
rect 1310 1697 1316 1698
rect 1310 1693 1311 1697
rect 1315 1693 1316 1697
rect 1310 1692 1316 1693
rect 1502 1697 1508 1698
rect 1502 1693 1503 1697
rect 1507 1693 1508 1697
rect 1502 1692 1508 1693
rect 1670 1697 1676 1698
rect 1670 1693 1671 1697
rect 1675 1693 1676 1697
rect 1670 1692 1676 1693
rect 1312 1671 1314 1692
rect 1504 1671 1506 1692
rect 1672 1671 1674 1692
rect 1231 1670 1235 1671
rect 1231 1665 1235 1666
rect 1311 1670 1315 1671
rect 1311 1665 1315 1666
rect 1431 1670 1435 1671
rect 1431 1665 1435 1666
rect 1503 1670 1507 1671
rect 1503 1665 1507 1666
rect 1639 1670 1643 1671
rect 1639 1665 1643 1666
rect 1671 1670 1675 1671
rect 1671 1665 1675 1666
rect 1232 1648 1234 1665
rect 1432 1648 1434 1665
rect 1640 1648 1642 1665
rect 1230 1647 1236 1648
rect 1230 1643 1231 1647
rect 1235 1643 1236 1647
rect 1230 1642 1236 1643
rect 1430 1647 1436 1648
rect 1430 1643 1431 1647
rect 1435 1643 1436 1647
rect 1430 1642 1436 1643
rect 1638 1647 1644 1648
rect 1638 1643 1639 1647
rect 1643 1643 1644 1647
rect 1638 1642 1644 1643
rect 1174 1639 1180 1640
rect 926 1635 932 1636
rect 926 1631 927 1635
rect 931 1631 932 1635
rect 926 1630 932 1631
rect 1110 1635 1116 1636
rect 1110 1631 1111 1635
rect 1115 1631 1116 1635
rect 1174 1635 1175 1639
rect 1179 1635 1180 1639
rect 1510 1639 1516 1640
rect 1174 1634 1180 1635
rect 1502 1635 1508 1636
rect 1110 1630 1116 1631
rect 1502 1631 1503 1635
rect 1507 1631 1508 1635
rect 1510 1635 1511 1639
rect 1515 1635 1516 1639
rect 1510 1634 1516 1635
rect 1502 1630 1508 1631
rect 854 1628 860 1629
rect 854 1624 855 1628
rect 859 1624 860 1628
rect 854 1623 860 1624
rect 722 1611 728 1612
rect 722 1607 723 1611
rect 727 1607 728 1611
rect 722 1606 728 1607
rect 856 1603 858 1623
rect 928 1612 930 1630
rect 1038 1628 1044 1629
rect 1038 1624 1039 1628
rect 1043 1624 1044 1628
rect 1038 1623 1044 1624
rect 910 1611 916 1612
rect 910 1607 911 1611
rect 915 1607 916 1611
rect 910 1606 916 1607
rect 926 1611 932 1612
rect 926 1607 927 1611
rect 931 1607 932 1611
rect 926 1606 932 1607
rect 671 1602 675 1603
rect 671 1597 675 1598
rect 687 1602 691 1603
rect 687 1597 691 1598
rect 815 1602 819 1603
rect 815 1597 819 1598
rect 855 1602 859 1603
rect 855 1597 859 1598
rect 606 1595 612 1596
rect 606 1591 607 1595
rect 611 1591 612 1595
rect 606 1590 612 1591
rect 614 1595 620 1596
rect 614 1591 615 1595
rect 619 1591 620 1595
rect 614 1590 620 1591
rect 542 1580 548 1581
rect 542 1576 543 1580
rect 547 1576 548 1580
rect 542 1575 548 1576
rect 616 1572 618 1590
rect 672 1581 674 1597
rect 742 1595 748 1596
rect 742 1591 743 1595
rect 747 1591 748 1595
rect 742 1590 748 1591
rect 670 1580 676 1581
rect 670 1576 671 1580
rect 675 1576 676 1580
rect 670 1575 676 1576
rect 744 1572 746 1590
rect 816 1581 818 1597
rect 814 1580 820 1581
rect 814 1576 815 1580
rect 819 1576 820 1580
rect 814 1575 820 1576
rect 912 1572 914 1606
rect 1040 1603 1042 1623
rect 1112 1612 1114 1630
rect 1230 1628 1236 1629
rect 1230 1624 1231 1628
rect 1235 1624 1236 1628
rect 1230 1623 1236 1624
rect 1430 1628 1436 1629
rect 1430 1624 1431 1628
rect 1435 1624 1436 1628
rect 1430 1623 1436 1624
rect 1110 1611 1116 1612
rect 1110 1607 1111 1611
rect 1115 1607 1116 1611
rect 1110 1606 1116 1607
rect 1232 1603 1234 1623
rect 1432 1603 1434 1623
rect 967 1602 971 1603
rect 967 1597 971 1598
rect 1039 1602 1043 1603
rect 1039 1597 1043 1598
rect 1119 1602 1123 1603
rect 1119 1597 1123 1598
rect 1231 1602 1235 1603
rect 1231 1597 1235 1598
rect 1279 1602 1283 1603
rect 1279 1597 1283 1598
rect 1431 1602 1435 1603
rect 1431 1597 1435 1598
rect 1439 1602 1443 1603
rect 1439 1597 1443 1598
rect 968 1581 970 1597
rect 1120 1581 1122 1597
rect 1190 1595 1196 1596
rect 1190 1591 1191 1595
rect 1195 1591 1196 1595
rect 1190 1590 1196 1591
rect 966 1580 972 1581
rect 966 1576 967 1580
rect 971 1576 972 1580
rect 966 1575 972 1576
rect 1118 1580 1124 1581
rect 1118 1576 1119 1580
rect 1123 1576 1124 1580
rect 1118 1575 1124 1576
rect 614 1571 620 1572
rect 614 1567 615 1571
rect 619 1567 620 1571
rect 614 1566 620 1567
rect 742 1571 748 1572
rect 742 1567 743 1571
rect 747 1567 748 1571
rect 742 1566 748 1567
rect 806 1571 812 1572
rect 806 1567 807 1571
rect 811 1567 812 1571
rect 806 1566 812 1567
rect 910 1571 916 1572
rect 910 1567 911 1571
rect 915 1567 916 1571
rect 910 1566 916 1567
rect 542 1561 548 1562
rect 542 1557 543 1561
rect 547 1557 548 1561
rect 542 1556 548 1557
rect 670 1561 676 1562
rect 670 1557 671 1561
rect 675 1557 676 1561
rect 670 1556 676 1557
rect 544 1535 546 1556
rect 672 1535 674 1556
rect 471 1534 475 1535
rect 471 1529 475 1530
rect 543 1534 547 1535
rect 543 1529 547 1530
rect 607 1534 611 1535
rect 607 1529 611 1530
rect 671 1534 675 1535
rect 671 1529 675 1530
rect 751 1534 755 1535
rect 751 1529 755 1530
rect 472 1512 474 1529
rect 608 1512 610 1529
rect 752 1512 754 1529
rect 470 1511 476 1512
rect 470 1507 471 1511
rect 475 1507 476 1511
rect 470 1506 476 1507
rect 606 1511 612 1512
rect 606 1507 607 1511
rect 611 1507 612 1511
rect 606 1506 612 1507
rect 750 1511 756 1512
rect 750 1507 751 1511
rect 755 1507 756 1511
rect 750 1506 756 1507
rect 462 1503 468 1504
rect 294 1499 300 1500
rect 110 1495 116 1496
rect 110 1491 111 1495
rect 115 1491 116 1495
rect 294 1495 295 1499
rect 299 1495 300 1499
rect 294 1494 300 1495
rect 414 1499 420 1500
rect 414 1495 415 1499
rect 419 1495 420 1499
rect 462 1499 463 1503
rect 467 1499 468 1503
rect 462 1498 468 1499
rect 550 1503 556 1504
rect 550 1499 551 1503
rect 555 1499 556 1503
rect 550 1498 556 1499
rect 414 1494 420 1495
rect 110 1490 116 1491
rect 222 1492 228 1493
rect 112 1463 114 1490
rect 222 1488 223 1492
rect 227 1488 228 1492
rect 222 1487 228 1488
rect 206 1475 212 1476
rect 206 1471 207 1475
rect 211 1471 212 1475
rect 206 1470 212 1471
rect 111 1462 115 1463
rect 111 1457 115 1458
rect 135 1462 139 1463
rect 135 1457 139 1458
rect 112 1438 114 1457
rect 136 1441 138 1457
rect 134 1440 140 1441
rect 110 1437 116 1438
rect 110 1433 111 1437
rect 115 1433 116 1437
rect 134 1436 135 1440
rect 139 1436 140 1440
rect 134 1435 140 1436
rect 110 1432 116 1433
rect 208 1432 210 1470
rect 224 1463 226 1487
rect 296 1476 298 1494
rect 342 1492 348 1493
rect 342 1488 343 1492
rect 347 1488 348 1492
rect 342 1487 348 1488
rect 294 1475 300 1476
rect 294 1471 295 1475
rect 299 1471 300 1475
rect 294 1470 300 1471
rect 344 1463 346 1487
rect 416 1476 418 1494
rect 470 1492 476 1493
rect 470 1488 471 1492
rect 475 1488 476 1492
rect 470 1487 476 1488
rect 414 1475 420 1476
rect 414 1471 415 1475
rect 419 1471 420 1475
rect 414 1470 420 1471
rect 472 1463 474 1487
rect 223 1462 227 1463
rect 223 1457 227 1458
rect 303 1462 307 1463
rect 303 1457 307 1458
rect 343 1462 347 1463
rect 343 1457 347 1458
rect 471 1462 475 1463
rect 471 1457 475 1458
rect 304 1441 306 1457
rect 358 1455 364 1456
rect 358 1451 359 1455
rect 363 1451 364 1455
rect 358 1450 364 1451
rect 302 1440 308 1441
rect 302 1436 303 1440
rect 307 1436 308 1440
rect 302 1435 308 1436
rect 206 1431 212 1432
rect 206 1427 207 1431
rect 211 1427 212 1431
rect 206 1426 212 1427
rect 134 1421 140 1422
rect 110 1420 116 1421
rect 110 1416 111 1420
rect 115 1416 116 1420
rect 134 1417 135 1421
rect 139 1417 140 1421
rect 134 1416 140 1417
rect 302 1421 308 1422
rect 302 1417 303 1421
rect 307 1417 308 1421
rect 302 1416 308 1417
rect 110 1415 116 1416
rect 112 1395 114 1415
rect 136 1395 138 1416
rect 304 1395 306 1416
rect 111 1394 115 1395
rect 111 1389 115 1390
rect 135 1394 139 1395
rect 135 1389 139 1390
rect 279 1394 283 1395
rect 279 1389 283 1390
rect 303 1394 307 1395
rect 303 1389 307 1390
rect 112 1373 114 1389
rect 110 1372 116 1373
rect 136 1372 138 1389
rect 280 1372 282 1389
rect 110 1368 111 1372
rect 115 1368 116 1372
rect 110 1367 116 1368
rect 134 1371 140 1372
rect 134 1367 135 1371
rect 139 1367 140 1371
rect 134 1366 140 1367
rect 278 1371 284 1372
rect 278 1367 279 1371
rect 283 1367 284 1371
rect 278 1366 284 1367
rect 360 1364 362 1450
rect 472 1441 474 1457
rect 552 1456 554 1498
rect 606 1492 612 1493
rect 606 1488 607 1492
rect 611 1488 612 1492
rect 606 1487 612 1488
rect 750 1492 756 1493
rect 750 1488 751 1492
rect 755 1488 756 1492
rect 750 1487 756 1488
rect 608 1463 610 1487
rect 752 1463 754 1487
rect 808 1476 810 1566
rect 814 1561 820 1562
rect 814 1557 815 1561
rect 819 1557 820 1561
rect 814 1556 820 1557
rect 966 1561 972 1562
rect 966 1557 967 1561
rect 971 1557 972 1561
rect 966 1556 972 1557
rect 1118 1561 1124 1562
rect 1118 1557 1119 1561
rect 1123 1557 1124 1561
rect 1118 1556 1124 1557
rect 816 1535 818 1556
rect 968 1535 970 1556
rect 1120 1535 1122 1556
rect 815 1534 819 1535
rect 815 1529 819 1530
rect 895 1534 899 1535
rect 895 1529 899 1530
rect 967 1534 971 1535
rect 967 1529 971 1530
rect 1047 1534 1051 1535
rect 1047 1529 1051 1530
rect 1119 1534 1123 1535
rect 1119 1529 1123 1530
rect 896 1512 898 1529
rect 1048 1512 1050 1529
rect 894 1511 900 1512
rect 894 1507 895 1511
rect 899 1507 900 1511
rect 894 1506 900 1507
rect 1046 1511 1052 1512
rect 1046 1507 1047 1511
rect 1051 1507 1052 1511
rect 1046 1506 1052 1507
rect 1192 1504 1194 1590
rect 1280 1581 1282 1597
rect 1440 1581 1442 1597
rect 1504 1596 1506 1630
rect 1512 1612 1514 1634
rect 1638 1628 1644 1629
rect 1638 1624 1639 1628
rect 1643 1624 1644 1628
rect 1638 1623 1644 1624
rect 1510 1611 1516 1612
rect 1510 1607 1511 1611
rect 1515 1607 1516 1611
rect 1510 1606 1516 1607
rect 1640 1603 1642 1623
rect 1736 1612 1738 1702
rect 1808 1699 1810 1723
rect 1880 1699 1882 1724
rect 2016 1699 2018 1724
rect 2152 1699 2154 1724
rect 1807 1698 1811 1699
rect 1766 1696 1772 1697
rect 1766 1692 1767 1696
rect 1771 1692 1772 1696
rect 1807 1693 1811 1694
rect 1831 1698 1835 1699
rect 1831 1693 1835 1694
rect 1879 1698 1883 1699
rect 1879 1693 1883 1694
rect 1935 1698 1939 1699
rect 1935 1693 1939 1694
rect 2015 1698 2019 1699
rect 2015 1693 2019 1694
rect 2063 1698 2067 1699
rect 2063 1693 2067 1694
rect 2151 1698 2155 1699
rect 2151 1693 2155 1694
rect 2183 1698 2187 1699
rect 2183 1693 2187 1694
rect 1766 1691 1772 1692
rect 1768 1671 1770 1691
rect 1808 1677 1810 1693
rect 1806 1676 1812 1677
rect 1832 1676 1834 1693
rect 1936 1676 1938 1693
rect 2064 1676 2066 1693
rect 2184 1676 2186 1693
rect 1806 1672 1807 1676
rect 1811 1672 1812 1676
rect 1806 1671 1812 1672
rect 1830 1675 1836 1676
rect 1830 1671 1831 1675
rect 1835 1671 1836 1675
rect 1767 1670 1771 1671
rect 1830 1670 1836 1671
rect 1934 1675 1940 1676
rect 1934 1671 1935 1675
rect 1939 1671 1940 1675
rect 1934 1670 1940 1671
rect 2062 1675 2068 1676
rect 2062 1671 2063 1675
rect 2067 1671 2068 1675
rect 2062 1670 2068 1671
rect 2182 1675 2188 1676
rect 2182 1671 2183 1675
rect 2187 1671 2188 1675
rect 2182 1670 2188 1671
rect 2256 1668 2258 1754
rect 2304 1749 2306 1765
rect 2328 1764 2330 1806
rect 2406 1804 2412 1805
rect 2406 1800 2407 1804
rect 2411 1800 2412 1804
rect 2406 1799 2412 1800
rect 2408 1771 2410 1799
rect 2428 1788 2430 1878
rect 2454 1873 2460 1874
rect 2454 1869 2455 1873
rect 2459 1869 2460 1873
rect 2454 1868 2460 1869
rect 2614 1873 2620 1874
rect 2614 1869 2615 1873
rect 2619 1869 2620 1873
rect 2614 1868 2620 1869
rect 2790 1873 2796 1874
rect 2790 1869 2791 1873
rect 2795 1869 2796 1873
rect 2790 1868 2796 1869
rect 2982 1873 2988 1874
rect 2982 1869 2983 1873
rect 2987 1869 2988 1873
rect 2982 1868 2988 1869
rect 2456 1847 2458 1868
rect 2616 1847 2618 1868
rect 2792 1847 2794 1868
rect 2984 1847 2986 1868
rect 2455 1846 2459 1847
rect 2455 1841 2459 1842
rect 2567 1846 2571 1847
rect 2567 1841 2571 1842
rect 2615 1846 2619 1847
rect 2615 1841 2619 1842
rect 2743 1846 2747 1847
rect 2743 1841 2747 1842
rect 2791 1846 2795 1847
rect 2791 1841 2795 1842
rect 2935 1846 2939 1847
rect 2935 1841 2939 1842
rect 2983 1846 2987 1847
rect 2983 1841 2987 1842
rect 2568 1824 2570 1841
rect 2744 1824 2746 1841
rect 2936 1824 2938 1841
rect 2566 1823 2572 1824
rect 2566 1819 2567 1823
rect 2571 1819 2572 1823
rect 2566 1818 2572 1819
rect 2742 1823 2748 1824
rect 2742 1819 2743 1823
rect 2747 1819 2748 1823
rect 2742 1818 2748 1819
rect 2934 1823 2940 1824
rect 2934 1819 2935 1823
rect 2939 1819 2940 1823
rect 2934 1818 2940 1819
rect 3080 1816 3082 1894
rect 3168 1884 3170 1910
rect 3175 1909 3179 1910
rect 3183 1914 3187 1915
rect 3183 1909 3187 1910
rect 3319 1914 3323 1915
rect 3319 1909 3323 1910
rect 3367 1914 3371 1915
rect 3367 1909 3371 1910
rect 3184 1893 3186 1909
rect 3368 1893 3370 1909
rect 3182 1892 3188 1893
rect 3182 1888 3183 1892
rect 3187 1888 3188 1892
rect 3182 1887 3188 1888
rect 3366 1892 3372 1893
rect 3366 1888 3367 1892
rect 3371 1888 3372 1892
rect 3366 1887 3372 1888
rect 3166 1883 3172 1884
rect 3166 1879 3167 1883
rect 3171 1879 3172 1883
rect 3166 1878 3172 1879
rect 3182 1873 3188 1874
rect 3182 1869 3183 1873
rect 3187 1869 3188 1873
rect 3182 1868 3188 1869
rect 3366 1873 3372 1874
rect 3366 1869 3367 1873
rect 3371 1869 3372 1873
rect 3366 1868 3372 1869
rect 3184 1847 3186 1868
rect 3368 1847 3370 1868
rect 3135 1846 3139 1847
rect 3135 1841 3139 1842
rect 3183 1846 3187 1847
rect 3183 1841 3187 1842
rect 3343 1846 3347 1847
rect 3343 1841 3347 1842
rect 3367 1846 3371 1847
rect 3367 1841 3371 1842
rect 3136 1824 3138 1841
rect 3344 1824 3346 1841
rect 3134 1823 3140 1824
rect 3134 1819 3135 1823
rect 3139 1819 3140 1823
rect 3134 1818 3140 1819
rect 3342 1823 3348 1824
rect 3342 1819 3343 1823
rect 3347 1819 3348 1823
rect 3342 1818 3348 1819
rect 3078 1815 3084 1816
rect 2478 1811 2484 1812
rect 2478 1807 2479 1811
rect 2483 1807 2484 1811
rect 2478 1806 2484 1807
rect 2638 1811 2644 1812
rect 2638 1807 2639 1811
rect 2643 1807 2644 1811
rect 2638 1806 2644 1807
rect 2814 1811 2820 1812
rect 2814 1807 2815 1811
rect 2819 1807 2820 1811
rect 2814 1806 2820 1807
rect 3006 1811 3012 1812
rect 3006 1807 3007 1811
rect 3011 1807 3012 1811
rect 3078 1811 3079 1815
rect 3083 1811 3084 1815
rect 3078 1810 3084 1811
rect 3270 1815 3276 1816
rect 3270 1811 3271 1815
rect 3275 1811 3276 1815
rect 3270 1810 3276 1811
rect 3006 1806 3012 1807
rect 2480 1788 2482 1806
rect 2566 1804 2572 1805
rect 2566 1800 2567 1804
rect 2571 1800 2572 1804
rect 2566 1799 2572 1800
rect 2426 1787 2432 1788
rect 2426 1783 2427 1787
rect 2431 1783 2432 1787
rect 2426 1782 2432 1783
rect 2462 1787 2468 1788
rect 2462 1783 2463 1787
rect 2467 1783 2468 1787
rect 2462 1782 2468 1783
rect 2478 1787 2484 1788
rect 2478 1783 2479 1787
rect 2483 1783 2484 1787
rect 2478 1782 2484 1783
rect 2407 1770 2411 1771
rect 2407 1765 2411 1766
rect 2326 1763 2332 1764
rect 2326 1759 2327 1763
rect 2331 1759 2332 1763
rect 2326 1758 2332 1759
rect 2302 1748 2308 1749
rect 2302 1744 2303 1748
rect 2307 1744 2308 1748
rect 2302 1743 2308 1744
rect 2464 1740 2466 1782
rect 2568 1771 2570 1799
rect 2640 1788 2642 1806
rect 2742 1804 2748 1805
rect 2742 1800 2743 1804
rect 2747 1800 2748 1804
rect 2742 1799 2748 1800
rect 2638 1787 2644 1788
rect 2638 1783 2639 1787
rect 2643 1783 2644 1787
rect 2638 1782 2644 1783
rect 2744 1771 2746 1799
rect 2816 1788 2818 1806
rect 2934 1804 2940 1805
rect 2934 1800 2935 1804
rect 2939 1800 2940 1804
rect 2934 1799 2940 1800
rect 2814 1787 2820 1788
rect 2814 1783 2815 1787
rect 2819 1783 2820 1787
rect 2814 1782 2820 1783
rect 2798 1771 2804 1772
rect 2936 1771 2938 1799
rect 3008 1788 3010 1806
rect 3134 1804 3140 1805
rect 3134 1800 3135 1804
rect 3139 1800 3140 1804
rect 3134 1799 3140 1800
rect 3006 1787 3012 1788
rect 3006 1783 3007 1787
rect 3011 1783 3012 1787
rect 3006 1782 3012 1783
rect 3136 1771 3138 1799
rect 2479 1770 2483 1771
rect 2479 1765 2483 1766
rect 2567 1770 2571 1771
rect 2567 1765 2571 1766
rect 2687 1770 2691 1771
rect 2687 1765 2691 1766
rect 2743 1770 2747 1771
rect 2798 1767 2799 1771
rect 2803 1767 2804 1771
rect 2798 1766 2804 1767
rect 2911 1770 2915 1771
rect 2743 1765 2747 1766
rect 2480 1749 2482 1765
rect 2558 1763 2564 1764
rect 2558 1759 2559 1763
rect 2563 1759 2564 1763
rect 2558 1758 2564 1759
rect 2478 1748 2484 1749
rect 2478 1744 2479 1748
rect 2483 1744 2484 1748
rect 2478 1743 2484 1744
rect 2560 1740 2562 1758
rect 2688 1749 2690 1765
rect 2686 1748 2692 1749
rect 2686 1744 2687 1748
rect 2691 1744 2692 1748
rect 2686 1743 2692 1744
rect 2366 1739 2372 1740
rect 2366 1735 2367 1739
rect 2371 1735 2372 1739
rect 2366 1734 2372 1735
rect 2462 1739 2468 1740
rect 2462 1735 2463 1739
rect 2467 1735 2468 1739
rect 2462 1734 2468 1735
rect 2558 1739 2564 1740
rect 2558 1735 2559 1739
rect 2563 1735 2564 1739
rect 2558 1734 2564 1735
rect 2302 1729 2308 1730
rect 2302 1725 2303 1729
rect 2307 1725 2308 1729
rect 2302 1724 2308 1725
rect 2304 1699 2306 1724
rect 2303 1698 2307 1699
rect 2303 1693 2307 1694
rect 2311 1698 2315 1699
rect 2311 1693 2315 1694
rect 2312 1676 2314 1693
rect 2310 1675 2316 1676
rect 2310 1671 2311 1675
rect 2315 1671 2316 1675
rect 2310 1670 2316 1671
rect 1767 1665 1771 1666
rect 2254 1667 2260 1668
rect 1768 1649 1770 1665
rect 1902 1663 1908 1664
rect 1806 1659 1812 1660
rect 1806 1655 1807 1659
rect 1811 1655 1812 1659
rect 1902 1659 1903 1663
rect 1907 1659 1908 1663
rect 1902 1658 1908 1659
rect 2006 1663 2012 1664
rect 2006 1659 2007 1663
rect 2011 1659 2012 1663
rect 2006 1658 2012 1659
rect 2134 1663 2140 1664
rect 2134 1659 2135 1663
rect 2139 1659 2140 1663
rect 2254 1663 2255 1667
rect 2259 1663 2260 1667
rect 2254 1662 2260 1663
rect 2134 1658 2140 1659
rect 1806 1654 1812 1655
rect 1830 1656 1836 1657
rect 1766 1648 1772 1649
rect 1766 1644 1767 1648
rect 1771 1644 1772 1648
rect 1766 1643 1772 1644
rect 1766 1631 1772 1632
rect 1766 1627 1767 1631
rect 1771 1627 1772 1631
rect 1808 1627 1810 1654
rect 1830 1652 1831 1656
rect 1835 1652 1836 1656
rect 1830 1651 1836 1652
rect 1832 1627 1834 1651
rect 1904 1640 1906 1658
rect 1934 1656 1940 1657
rect 1934 1652 1935 1656
rect 1939 1652 1940 1656
rect 1934 1651 1940 1652
rect 1894 1639 1900 1640
rect 1894 1635 1895 1639
rect 1899 1635 1900 1639
rect 1894 1634 1900 1635
rect 1902 1639 1908 1640
rect 1902 1635 1903 1639
rect 1907 1635 1908 1639
rect 1902 1634 1908 1635
rect 1766 1626 1772 1627
rect 1807 1626 1811 1627
rect 1734 1611 1740 1612
rect 1734 1607 1735 1611
rect 1739 1607 1740 1611
rect 1734 1606 1740 1607
rect 1768 1603 1770 1626
rect 1807 1621 1811 1622
rect 1831 1626 1835 1627
rect 1831 1621 1835 1622
rect 1607 1602 1611 1603
rect 1607 1597 1611 1598
rect 1639 1602 1643 1603
rect 1639 1597 1643 1598
rect 1767 1602 1771 1603
rect 1808 1602 1810 1621
rect 1832 1605 1834 1621
rect 1830 1604 1836 1605
rect 1767 1597 1771 1598
rect 1806 1601 1812 1602
rect 1806 1597 1807 1601
rect 1811 1597 1812 1601
rect 1830 1600 1831 1604
rect 1835 1600 1836 1604
rect 1830 1599 1836 1600
rect 1502 1595 1508 1596
rect 1502 1591 1503 1595
rect 1507 1591 1508 1595
rect 1502 1590 1508 1591
rect 1510 1595 1516 1596
rect 1510 1591 1511 1595
rect 1515 1591 1516 1595
rect 1510 1590 1516 1591
rect 1278 1580 1284 1581
rect 1278 1576 1279 1580
rect 1283 1576 1284 1580
rect 1278 1575 1284 1576
rect 1438 1580 1444 1581
rect 1438 1576 1439 1580
rect 1443 1576 1444 1580
rect 1438 1575 1444 1576
rect 1512 1572 1514 1590
rect 1608 1581 1610 1597
rect 1606 1580 1612 1581
rect 1606 1576 1607 1580
rect 1611 1576 1612 1580
rect 1768 1578 1770 1597
rect 1806 1596 1812 1597
rect 1896 1596 1898 1634
rect 1936 1627 1938 1651
rect 2008 1640 2010 1658
rect 2062 1656 2068 1657
rect 2062 1652 2063 1656
rect 2067 1652 2068 1656
rect 2062 1651 2068 1652
rect 2006 1639 2012 1640
rect 2006 1635 2007 1639
rect 2011 1635 2012 1639
rect 2006 1634 2012 1635
rect 2064 1627 2066 1651
rect 2136 1640 2138 1658
rect 2182 1656 2188 1657
rect 2182 1652 2183 1656
rect 2187 1652 2188 1656
rect 2182 1651 2188 1652
rect 2310 1656 2316 1657
rect 2310 1652 2311 1656
rect 2315 1652 2316 1656
rect 2310 1651 2316 1652
rect 2134 1639 2140 1640
rect 2134 1635 2135 1639
rect 2139 1635 2140 1639
rect 2134 1634 2140 1635
rect 2184 1627 2186 1651
rect 2312 1627 2314 1651
rect 2368 1640 2370 1734
rect 2478 1729 2484 1730
rect 2478 1725 2479 1729
rect 2483 1725 2484 1729
rect 2478 1724 2484 1725
rect 2686 1729 2692 1730
rect 2686 1725 2687 1729
rect 2691 1725 2692 1729
rect 2686 1724 2692 1725
rect 2480 1699 2482 1724
rect 2688 1699 2690 1724
rect 2439 1698 2443 1699
rect 2439 1693 2443 1694
rect 2479 1698 2483 1699
rect 2479 1693 2483 1694
rect 2575 1698 2579 1699
rect 2575 1693 2579 1694
rect 2687 1698 2691 1699
rect 2687 1693 2691 1694
rect 2727 1698 2731 1699
rect 2727 1693 2731 1694
rect 2440 1676 2442 1693
rect 2576 1676 2578 1693
rect 2728 1676 2730 1693
rect 2438 1675 2444 1676
rect 2438 1671 2439 1675
rect 2443 1671 2444 1675
rect 2438 1670 2444 1671
rect 2574 1675 2580 1676
rect 2574 1671 2575 1675
rect 2579 1671 2580 1675
rect 2574 1670 2580 1671
rect 2726 1675 2732 1676
rect 2726 1671 2727 1675
rect 2731 1671 2732 1675
rect 2726 1670 2732 1671
rect 2800 1668 2802 1766
rect 2911 1765 2915 1766
rect 2935 1770 2939 1771
rect 2935 1765 2939 1766
rect 3135 1770 3139 1771
rect 3135 1765 3139 1766
rect 3151 1770 3155 1771
rect 3151 1765 3155 1766
rect 2912 1749 2914 1765
rect 2982 1763 2988 1764
rect 2982 1759 2983 1763
rect 2987 1759 2988 1763
rect 2982 1758 2988 1759
rect 2910 1748 2916 1749
rect 2910 1744 2911 1748
rect 2915 1744 2916 1748
rect 2910 1743 2916 1744
rect 2984 1740 2986 1758
rect 3152 1749 3154 1765
rect 3150 1748 3156 1749
rect 3150 1744 3151 1748
rect 3155 1744 3156 1748
rect 3150 1743 3156 1744
rect 2982 1739 2988 1740
rect 2982 1735 2983 1739
rect 2987 1735 2988 1739
rect 2982 1734 2988 1735
rect 2910 1729 2916 1730
rect 2910 1725 2911 1729
rect 2915 1725 2916 1729
rect 2910 1724 2916 1725
rect 3150 1729 3156 1730
rect 3150 1725 3151 1729
rect 3155 1725 3156 1729
rect 3150 1724 3156 1725
rect 2912 1699 2914 1724
rect 3152 1699 3154 1724
rect 2887 1698 2891 1699
rect 2887 1693 2891 1694
rect 2911 1698 2915 1699
rect 2911 1693 2915 1694
rect 3047 1698 3051 1699
rect 3047 1693 3051 1694
rect 3151 1698 3155 1699
rect 3151 1693 3155 1694
rect 3215 1698 3219 1699
rect 3215 1693 3219 1694
rect 2888 1676 2890 1693
rect 3048 1676 3050 1693
rect 3216 1676 3218 1693
rect 2886 1675 2892 1676
rect 2886 1671 2887 1675
rect 2891 1671 2892 1675
rect 2886 1670 2892 1671
rect 3046 1675 3052 1676
rect 3046 1671 3047 1675
rect 3051 1671 3052 1675
rect 3046 1670 3052 1671
rect 3214 1675 3220 1676
rect 3214 1671 3215 1675
rect 3219 1671 3220 1675
rect 3214 1670 3220 1671
rect 2798 1667 2804 1668
rect 2382 1663 2388 1664
rect 2382 1659 2383 1663
rect 2387 1659 2388 1663
rect 2382 1658 2388 1659
rect 2510 1663 2516 1664
rect 2510 1659 2511 1663
rect 2515 1659 2516 1663
rect 2510 1658 2516 1659
rect 2646 1663 2652 1664
rect 2646 1659 2647 1663
rect 2651 1659 2652 1663
rect 2798 1663 2799 1667
rect 2803 1663 2804 1667
rect 2798 1662 2804 1663
rect 2806 1667 2812 1668
rect 2806 1663 2807 1667
rect 2811 1663 2812 1667
rect 2806 1662 2812 1663
rect 2966 1667 2972 1668
rect 2966 1663 2967 1667
rect 2971 1663 2972 1667
rect 2966 1662 2972 1663
rect 3186 1667 3192 1668
rect 3186 1663 3187 1667
rect 3191 1663 3192 1667
rect 3186 1662 3192 1663
rect 2646 1658 2652 1659
rect 2366 1639 2372 1640
rect 2366 1635 2367 1639
rect 2371 1635 2372 1639
rect 2366 1634 2372 1635
rect 1935 1626 1939 1627
rect 1935 1621 1939 1622
rect 1943 1626 1947 1627
rect 1943 1621 1947 1622
rect 2063 1626 2067 1627
rect 2063 1621 2067 1622
rect 2087 1626 2091 1627
rect 2087 1621 2091 1622
rect 2183 1626 2187 1627
rect 2183 1621 2187 1622
rect 2231 1626 2235 1627
rect 2231 1621 2235 1622
rect 2311 1626 2315 1627
rect 2311 1621 2315 1622
rect 2367 1626 2371 1627
rect 2367 1621 2371 1622
rect 1910 1619 1916 1620
rect 1910 1615 1911 1619
rect 1915 1615 1916 1619
rect 1910 1614 1916 1615
rect 1912 1596 1914 1614
rect 1944 1605 1946 1621
rect 2022 1619 2028 1620
rect 2022 1615 2023 1619
rect 2027 1615 2028 1619
rect 2022 1614 2028 1615
rect 1942 1604 1948 1605
rect 1942 1600 1943 1604
rect 1947 1600 1948 1604
rect 1942 1599 1948 1600
rect 2024 1596 2026 1614
rect 2088 1605 2090 1621
rect 2166 1619 2172 1620
rect 2166 1615 2167 1619
rect 2171 1615 2172 1619
rect 2166 1614 2172 1615
rect 2086 1604 2092 1605
rect 2086 1600 2087 1604
rect 2091 1600 2092 1604
rect 2086 1599 2092 1600
rect 2168 1596 2170 1614
rect 2232 1605 2234 1621
rect 2286 1619 2292 1620
rect 2286 1615 2287 1619
rect 2291 1615 2292 1619
rect 2286 1614 2292 1615
rect 2230 1604 2236 1605
rect 2230 1600 2231 1604
rect 2235 1600 2236 1604
rect 2230 1599 2236 1600
rect 1894 1595 1900 1596
rect 1894 1591 1895 1595
rect 1899 1591 1900 1595
rect 1894 1590 1900 1591
rect 1910 1595 1916 1596
rect 1910 1591 1911 1595
rect 1915 1591 1916 1595
rect 1910 1590 1916 1591
rect 2022 1595 2028 1596
rect 2022 1591 2023 1595
rect 2027 1591 2028 1595
rect 2022 1590 2028 1591
rect 2166 1595 2172 1596
rect 2166 1591 2167 1595
rect 2171 1591 2172 1595
rect 2166 1590 2172 1591
rect 1830 1585 1836 1586
rect 1806 1584 1812 1585
rect 1806 1580 1807 1584
rect 1811 1580 1812 1584
rect 1830 1581 1831 1585
rect 1835 1581 1836 1585
rect 1830 1580 1836 1581
rect 1942 1585 1948 1586
rect 1942 1581 1943 1585
rect 1947 1581 1948 1585
rect 1942 1580 1948 1581
rect 2086 1585 2092 1586
rect 2086 1581 2087 1585
rect 2091 1581 2092 1585
rect 2086 1580 2092 1581
rect 2230 1585 2236 1586
rect 2230 1581 2231 1585
rect 2235 1581 2236 1585
rect 2230 1580 2236 1581
rect 1806 1579 1812 1580
rect 1606 1575 1612 1576
rect 1766 1577 1772 1578
rect 1766 1573 1767 1577
rect 1771 1573 1772 1577
rect 1766 1572 1772 1573
rect 1362 1571 1368 1572
rect 1362 1567 1363 1571
rect 1367 1567 1368 1571
rect 1362 1566 1368 1567
rect 1510 1571 1516 1572
rect 1510 1567 1511 1571
rect 1515 1567 1516 1571
rect 1510 1566 1516 1567
rect 1278 1561 1284 1562
rect 1278 1557 1279 1561
rect 1283 1557 1284 1561
rect 1278 1556 1284 1557
rect 1280 1535 1282 1556
rect 1199 1534 1203 1535
rect 1199 1529 1203 1530
rect 1279 1534 1283 1535
rect 1279 1529 1283 1530
rect 1351 1534 1355 1535
rect 1351 1529 1355 1530
rect 1200 1512 1202 1529
rect 1352 1512 1354 1529
rect 1198 1511 1204 1512
rect 1198 1507 1199 1511
rect 1203 1507 1204 1511
rect 1198 1506 1204 1507
rect 1350 1511 1356 1512
rect 1350 1507 1351 1511
rect 1355 1507 1356 1511
rect 1350 1506 1356 1507
rect 1190 1503 1196 1504
rect 966 1499 972 1500
rect 966 1495 967 1499
rect 971 1495 972 1499
rect 966 1494 972 1495
rect 1118 1499 1124 1500
rect 1118 1495 1119 1499
rect 1123 1495 1124 1499
rect 1190 1499 1191 1503
rect 1195 1499 1196 1503
rect 1190 1498 1196 1499
rect 1118 1494 1124 1495
rect 894 1492 900 1493
rect 894 1488 895 1492
rect 899 1488 900 1492
rect 894 1487 900 1488
rect 806 1475 812 1476
rect 806 1471 807 1475
rect 811 1471 812 1475
rect 806 1470 812 1471
rect 896 1463 898 1487
rect 968 1476 970 1494
rect 1046 1492 1052 1493
rect 1046 1488 1047 1492
rect 1051 1488 1052 1492
rect 1046 1487 1052 1488
rect 966 1475 972 1476
rect 966 1471 967 1475
rect 971 1471 972 1475
rect 966 1470 972 1471
rect 1010 1467 1016 1468
rect 1010 1463 1011 1467
rect 1015 1463 1016 1467
rect 1048 1463 1050 1487
rect 1120 1476 1122 1494
rect 1198 1492 1204 1493
rect 1198 1488 1199 1492
rect 1203 1488 1204 1492
rect 1198 1487 1204 1488
rect 1350 1492 1356 1493
rect 1350 1488 1351 1492
rect 1355 1488 1356 1492
rect 1350 1487 1356 1488
rect 1118 1475 1124 1476
rect 1118 1471 1119 1475
rect 1123 1471 1124 1475
rect 1118 1470 1124 1471
rect 1200 1463 1202 1487
rect 1352 1463 1354 1487
rect 1364 1476 1366 1566
rect 1438 1561 1444 1562
rect 1438 1557 1439 1561
rect 1443 1557 1444 1561
rect 1438 1556 1444 1557
rect 1606 1561 1612 1562
rect 1606 1557 1607 1561
rect 1611 1557 1612 1561
rect 1606 1556 1612 1557
rect 1766 1560 1772 1561
rect 1766 1556 1767 1560
rect 1771 1556 1772 1560
rect 1440 1535 1442 1556
rect 1608 1535 1610 1556
rect 1766 1555 1772 1556
rect 1808 1555 1810 1579
rect 1832 1555 1834 1580
rect 1944 1555 1946 1580
rect 2088 1555 2090 1580
rect 2232 1555 2234 1580
rect 1768 1535 1770 1555
rect 1807 1554 1811 1555
rect 1807 1549 1811 1550
rect 1831 1554 1835 1555
rect 1831 1549 1835 1550
rect 1839 1554 1843 1555
rect 1839 1549 1843 1550
rect 1943 1554 1947 1555
rect 1943 1549 1947 1550
rect 1991 1554 1995 1555
rect 1991 1549 1995 1550
rect 2087 1554 2091 1555
rect 2087 1549 2091 1550
rect 2151 1554 2155 1555
rect 2151 1549 2155 1550
rect 2231 1554 2235 1555
rect 2231 1549 2235 1550
rect 1439 1534 1443 1535
rect 1439 1529 1443 1530
rect 1503 1534 1507 1535
rect 1503 1529 1507 1530
rect 1607 1534 1611 1535
rect 1607 1529 1611 1530
rect 1767 1534 1771 1535
rect 1808 1533 1810 1549
rect 1767 1529 1771 1530
rect 1806 1532 1812 1533
rect 1840 1532 1842 1549
rect 1992 1532 1994 1549
rect 2152 1532 2154 1549
rect 1504 1512 1506 1529
rect 1768 1513 1770 1529
rect 1806 1528 1807 1532
rect 1811 1528 1812 1532
rect 1806 1527 1812 1528
rect 1838 1531 1844 1532
rect 1838 1527 1839 1531
rect 1843 1527 1844 1531
rect 1838 1526 1844 1527
rect 1990 1531 1996 1532
rect 1990 1527 1991 1531
rect 1995 1527 1996 1531
rect 1990 1526 1996 1527
rect 2150 1531 2156 1532
rect 2150 1527 2151 1531
rect 2155 1527 2156 1531
rect 2150 1526 2156 1527
rect 2288 1524 2290 1614
rect 2368 1605 2370 1621
rect 2384 1620 2386 1658
rect 2438 1656 2444 1657
rect 2438 1652 2439 1656
rect 2443 1652 2444 1656
rect 2438 1651 2444 1652
rect 2440 1627 2442 1651
rect 2512 1640 2514 1658
rect 2574 1656 2580 1657
rect 2574 1652 2575 1656
rect 2579 1652 2580 1656
rect 2574 1651 2580 1652
rect 2510 1639 2516 1640
rect 2510 1635 2511 1639
rect 2515 1635 2516 1639
rect 2510 1634 2516 1635
rect 2576 1627 2578 1651
rect 2648 1640 2650 1658
rect 2726 1656 2732 1657
rect 2726 1652 2727 1656
rect 2731 1652 2732 1656
rect 2726 1651 2732 1652
rect 2646 1639 2652 1640
rect 2646 1635 2647 1639
rect 2651 1635 2652 1639
rect 2646 1634 2652 1635
rect 2728 1627 2730 1651
rect 2808 1648 2810 1662
rect 2886 1656 2892 1657
rect 2886 1652 2887 1656
rect 2891 1652 2892 1656
rect 2886 1651 2892 1652
rect 2806 1647 2812 1648
rect 2806 1643 2807 1647
rect 2811 1643 2812 1647
rect 2806 1642 2812 1643
rect 2888 1627 2890 1651
rect 2968 1640 2970 1662
rect 3046 1656 3052 1657
rect 3046 1652 3047 1656
rect 3051 1652 3052 1656
rect 3046 1651 3052 1652
rect 2966 1639 2972 1640
rect 2966 1635 2967 1639
rect 2971 1635 2972 1639
rect 2966 1634 2972 1635
rect 3048 1627 3050 1651
rect 3086 1639 3092 1640
rect 3086 1635 3087 1639
rect 3091 1635 3092 1639
rect 3086 1634 3092 1635
rect 2439 1626 2443 1627
rect 2439 1621 2443 1622
rect 2503 1626 2507 1627
rect 2503 1621 2507 1622
rect 2575 1626 2579 1627
rect 2575 1621 2579 1622
rect 2639 1626 2643 1627
rect 2639 1621 2643 1622
rect 2727 1626 2731 1627
rect 2727 1621 2731 1622
rect 2767 1626 2771 1627
rect 2767 1621 2771 1622
rect 2887 1626 2891 1627
rect 2887 1621 2891 1622
rect 2895 1626 2899 1627
rect 2895 1621 2899 1622
rect 3015 1626 3019 1627
rect 3015 1621 3019 1622
rect 3047 1626 3051 1627
rect 3047 1621 3051 1622
rect 2382 1619 2388 1620
rect 2382 1615 2383 1619
rect 2387 1615 2388 1619
rect 2382 1614 2388 1615
rect 2504 1605 2506 1621
rect 2558 1619 2564 1620
rect 2558 1615 2559 1619
rect 2563 1615 2564 1619
rect 2558 1614 2564 1615
rect 2366 1604 2372 1605
rect 2366 1600 2367 1604
rect 2371 1600 2372 1604
rect 2366 1599 2372 1600
rect 2502 1604 2508 1605
rect 2502 1600 2503 1604
rect 2507 1600 2508 1604
rect 2502 1599 2508 1600
rect 2438 1595 2444 1596
rect 2438 1591 2439 1595
rect 2443 1591 2444 1595
rect 2438 1590 2444 1591
rect 2366 1585 2372 1586
rect 2366 1581 2367 1585
rect 2371 1581 2372 1585
rect 2366 1580 2372 1581
rect 2368 1555 2370 1580
rect 2303 1554 2307 1555
rect 2303 1549 2307 1550
rect 2367 1554 2371 1555
rect 2367 1549 2371 1550
rect 2304 1532 2306 1549
rect 2302 1531 2308 1532
rect 2302 1527 2303 1531
rect 2307 1527 2308 1531
rect 2302 1526 2308 1527
rect 2286 1523 2292 1524
rect 1910 1519 1916 1520
rect 1806 1515 1812 1516
rect 1766 1512 1772 1513
rect 1502 1511 1508 1512
rect 1502 1507 1503 1511
rect 1507 1507 1508 1511
rect 1766 1508 1767 1512
rect 1771 1508 1772 1512
rect 1806 1511 1807 1515
rect 1811 1511 1812 1515
rect 1910 1515 1911 1519
rect 1915 1515 1916 1519
rect 1910 1514 1916 1515
rect 2062 1519 2068 1520
rect 2062 1515 2063 1519
rect 2067 1515 2068 1519
rect 2062 1514 2068 1515
rect 2222 1519 2228 1520
rect 2222 1515 2223 1519
rect 2227 1515 2228 1519
rect 2286 1519 2287 1523
rect 2291 1519 2292 1523
rect 2286 1518 2292 1519
rect 2222 1514 2228 1515
rect 1806 1510 1812 1511
rect 1838 1512 1844 1513
rect 1766 1507 1772 1508
rect 1502 1506 1508 1507
rect 1422 1499 1428 1500
rect 1422 1495 1423 1499
rect 1427 1495 1428 1499
rect 1422 1494 1428 1495
rect 1574 1499 1580 1500
rect 1574 1495 1575 1499
rect 1579 1495 1580 1499
rect 1574 1494 1580 1495
rect 1766 1495 1772 1496
rect 1424 1476 1426 1494
rect 1502 1492 1508 1493
rect 1502 1488 1503 1492
rect 1507 1488 1508 1492
rect 1502 1487 1508 1488
rect 1362 1475 1368 1476
rect 1362 1471 1363 1475
rect 1367 1471 1368 1475
rect 1362 1470 1368 1471
rect 1422 1475 1428 1476
rect 1422 1471 1423 1475
rect 1427 1471 1428 1475
rect 1422 1470 1428 1471
rect 1504 1463 1506 1487
rect 607 1462 611 1463
rect 607 1457 611 1458
rect 631 1462 635 1463
rect 631 1457 635 1458
rect 751 1462 755 1463
rect 751 1457 755 1458
rect 783 1462 787 1463
rect 783 1457 787 1458
rect 895 1462 899 1463
rect 895 1457 899 1458
rect 927 1462 931 1463
rect 1010 1462 1016 1463
rect 1047 1462 1051 1463
rect 927 1457 931 1458
rect 550 1455 556 1456
rect 550 1451 551 1455
rect 555 1451 556 1455
rect 550 1450 556 1451
rect 598 1455 604 1456
rect 598 1451 599 1455
rect 603 1451 604 1455
rect 598 1450 604 1451
rect 470 1440 476 1441
rect 470 1436 471 1440
rect 475 1436 476 1440
rect 470 1435 476 1436
rect 600 1432 602 1450
rect 632 1441 634 1457
rect 702 1455 708 1456
rect 702 1451 703 1455
rect 707 1451 708 1455
rect 702 1450 708 1451
rect 630 1440 636 1441
rect 630 1436 631 1440
rect 635 1436 636 1440
rect 630 1435 636 1436
rect 704 1432 706 1450
rect 784 1441 786 1457
rect 928 1441 930 1457
rect 974 1455 980 1456
rect 974 1451 975 1455
rect 979 1451 980 1455
rect 974 1450 980 1451
rect 998 1455 1004 1456
rect 998 1451 999 1455
rect 1003 1451 1004 1455
rect 998 1450 1004 1451
rect 782 1440 788 1441
rect 782 1436 783 1440
rect 787 1436 788 1440
rect 782 1435 788 1436
rect 926 1440 932 1441
rect 926 1436 927 1440
rect 931 1436 932 1440
rect 926 1435 932 1436
rect 598 1431 604 1432
rect 598 1427 599 1431
rect 603 1427 604 1431
rect 598 1426 604 1427
rect 702 1431 708 1432
rect 702 1427 703 1431
rect 707 1427 708 1431
rect 702 1426 708 1427
rect 846 1431 852 1432
rect 846 1427 847 1431
rect 851 1427 852 1431
rect 846 1426 852 1427
rect 470 1421 476 1422
rect 470 1417 471 1421
rect 475 1417 476 1421
rect 470 1416 476 1417
rect 630 1421 636 1422
rect 630 1417 631 1421
rect 635 1417 636 1421
rect 630 1416 636 1417
rect 782 1421 788 1422
rect 782 1417 783 1421
rect 787 1417 788 1421
rect 782 1416 788 1417
rect 472 1395 474 1416
rect 632 1395 634 1416
rect 784 1395 786 1416
rect 447 1394 451 1395
rect 447 1389 451 1390
rect 471 1394 475 1395
rect 471 1389 475 1390
rect 607 1394 611 1395
rect 607 1389 611 1390
rect 631 1394 635 1395
rect 631 1389 635 1390
rect 759 1394 763 1395
rect 759 1389 763 1390
rect 783 1394 787 1395
rect 783 1389 787 1390
rect 448 1372 450 1389
rect 608 1372 610 1389
rect 760 1372 762 1389
rect 446 1371 452 1372
rect 446 1367 447 1371
rect 451 1367 452 1371
rect 446 1366 452 1367
rect 606 1371 612 1372
rect 606 1367 607 1371
rect 611 1367 612 1371
rect 606 1366 612 1367
rect 758 1371 764 1372
rect 758 1367 759 1371
rect 763 1367 764 1371
rect 758 1366 764 1367
rect 358 1363 364 1364
rect 206 1359 212 1360
rect 110 1355 116 1356
rect 110 1351 111 1355
rect 115 1351 116 1355
rect 206 1355 207 1359
rect 211 1355 212 1359
rect 206 1354 212 1355
rect 350 1359 356 1360
rect 350 1355 351 1359
rect 355 1355 356 1359
rect 358 1359 359 1363
rect 363 1359 364 1363
rect 358 1358 364 1359
rect 558 1363 564 1364
rect 558 1359 559 1363
rect 563 1359 564 1363
rect 558 1358 564 1359
rect 738 1363 744 1364
rect 738 1359 739 1363
rect 743 1359 744 1363
rect 738 1358 744 1359
rect 350 1354 356 1355
rect 110 1350 116 1351
rect 134 1352 140 1353
rect 112 1327 114 1350
rect 134 1348 135 1352
rect 139 1348 140 1352
rect 134 1347 140 1348
rect 136 1327 138 1347
rect 208 1336 210 1354
rect 278 1352 284 1353
rect 278 1348 279 1352
rect 283 1348 284 1352
rect 278 1347 284 1348
rect 198 1335 204 1336
rect 198 1331 199 1335
rect 203 1331 204 1335
rect 198 1330 204 1331
rect 206 1335 212 1336
rect 206 1331 207 1335
rect 211 1331 212 1335
rect 206 1330 212 1331
rect 111 1326 115 1327
rect 111 1321 115 1322
rect 135 1326 139 1327
rect 135 1321 139 1322
rect 112 1302 114 1321
rect 136 1305 138 1321
rect 134 1304 140 1305
rect 110 1301 116 1302
rect 110 1297 111 1301
rect 115 1297 116 1301
rect 134 1300 135 1304
rect 139 1300 140 1304
rect 134 1299 140 1300
rect 110 1296 116 1297
rect 200 1296 202 1330
rect 280 1327 282 1347
rect 352 1336 354 1354
rect 446 1352 452 1353
rect 446 1348 447 1352
rect 451 1348 452 1352
rect 446 1347 452 1348
rect 350 1335 356 1336
rect 350 1331 351 1335
rect 355 1331 356 1335
rect 350 1330 356 1331
rect 448 1327 450 1347
rect 560 1328 562 1358
rect 606 1352 612 1353
rect 606 1348 607 1352
rect 611 1348 612 1352
rect 606 1347 612 1348
rect 558 1327 564 1328
rect 608 1327 610 1347
rect 740 1336 742 1358
rect 758 1352 764 1353
rect 758 1348 759 1352
rect 763 1348 764 1352
rect 758 1347 764 1348
rect 738 1335 744 1336
rect 738 1331 739 1335
rect 743 1331 744 1335
rect 738 1330 744 1331
rect 760 1327 762 1347
rect 848 1336 850 1426
rect 926 1421 932 1422
rect 926 1417 927 1421
rect 931 1417 932 1421
rect 926 1416 932 1417
rect 928 1395 930 1416
rect 903 1394 907 1395
rect 903 1389 907 1390
rect 927 1394 931 1395
rect 927 1389 931 1390
rect 904 1372 906 1389
rect 902 1371 908 1372
rect 902 1367 903 1371
rect 907 1367 908 1371
rect 902 1366 908 1367
rect 976 1364 978 1450
rect 1000 1432 1002 1450
rect 1012 1432 1014 1462
rect 1047 1457 1051 1458
rect 1063 1462 1067 1463
rect 1063 1457 1067 1458
rect 1199 1462 1203 1463
rect 1199 1457 1203 1458
rect 1335 1462 1339 1463
rect 1335 1457 1339 1458
rect 1351 1462 1355 1463
rect 1351 1457 1355 1458
rect 1471 1462 1475 1463
rect 1471 1457 1475 1458
rect 1503 1462 1507 1463
rect 1503 1457 1507 1458
rect 1064 1441 1066 1457
rect 1200 1441 1202 1457
rect 1278 1455 1284 1456
rect 1278 1451 1279 1455
rect 1283 1451 1284 1455
rect 1278 1450 1284 1451
rect 1062 1440 1068 1441
rect 1062 1436 1063 1440
rect 1067 1436 1068 1440
rect 1062 1435 1068 1436
rect 1198 1440 1204 1441
rect 1198 1436 1199 1440
rect 1203 1436 1204 1440
rect 1198 1435 1204 1436
rect 1280 1432 1282 1450
rect 1336 1441 1338 1457
rect 1414 1455 1420 1456
rect 1414 1451 1415 1455
rect 1419 1451 1420 1455
rect 1414 1450 1420 1451
rect 1334 1440 1340 1441
rect 1334 1436 1335 1440
rect 1339 1436 1340 1440
rect 1334 1435 1340 1436
rect 1416 1432 1418 1450
rect 1472 1441 1474 1457
rect 1576 1456 1578 1494
rect 1766 1491 1767 1495
rect 1771 1491 1772 1495
rect 1766 1490 1772 1491
rect 1768 1463 1770 1490
rect 1808 1483 1810 1510
rect 1838 1508 1839 1512
rect 1843 1508 1844 1512
rect 1838 1507 1844 1508
rect 1840 1483 1842 1507
rect 1912 1496 1914 1514
rect 1990 1512 1996 1513
rect 1990 1508 1991 1512
rect 1995 1508 1996 1512
rect 1990 1507 1996 1508
rect 1894 1495 1900 1496
rect 1894 1491 1895 1495
rect 1899 1491 1900 1495
rect 1894 1490 1900 1491
rect 1910 1495 1916 1496
rect 1910 1491 1911 1495
rect 1915 1491 1916 1495
rect 1910 1490 1916 1491
rect 1807 1482 1811 1483
rect 1807 1477 1811 1478
rect 1839 1482 1843 1483
rect 1839 1477 1843 1478
rect 1767 1462 1771 1463
rect 1808 1458 1810 1477
rect 1767 1457 1771 1458
rect 1806 1457 1812 1458
rect 1574 1455 1580 1456
rect 1574 1451 1575 1455
rect 1579 1451 1580 1455
rect 1574 1450 1580 1451
rect 1470 1440 1476 1441
rect 1470 1436 1471 1440
rect 1475 1436 1476 1440
rect 1768 1438 1770 1457
rect 1806 1453 1807 1457
rect 1811 1453 1812 1457
rect 1806 1452 1812 1453
rect 1896 1452 1898 1490
rect 1992 1483 1994 1507
rect 2064 1496 2066 1514
rect 2150 1512 2156 1513
rect 2150 1508 2151 1512
rect 2155 1508 2156 1512
rect 2150 1507 2156 1508
rect 2062 1495 2068 1496
rect 2062 1491 2063 1495
rect 2067 1491 2068 1495
rect 2062 1490 2068 1491
rect 2152 1483 2154 1507
rect 2224 1496 2226 1514
rect 2302 1512 2308 1513
rect 2302 1508 2303 1512
rect 2307 1508 2308 1512
rect 2302 1507 2308 1508
rect 2222 1495 2228 1496
rect 2222 1491 2223 1495
rect 2227 1491 2228 1495
rect 2222 1490 2228 1491
rect 2304 1483 2306 1507
rect 2440 1496 2442 1590
rect 2502 1585 2508 1586
rect 2502 1581 2503 1585
rect 2507 1581 2508 1585
rect 2502 1580 2508 1581
rect 2504 1555 2506 1580
rect 2455 1554 2459 1555
rect 2455 1549 2459 1550
rect 2503 1554 2507 1555
rect 2503 1549 2507 1550
rect 2456 1532 2458 1549
rect 2454 1531 2460 1532
rect 2454 1527 2455 1531
rect 2459 1527 2460 1531
rect 2454 1526 2460 1527
rect 2560 1524 2562 1614
rect 2640 1605 2642 1621
rect 2710 1619 2716 1620
rect 2710 1615 2711 1619
rect 2715 1615 2716 1619
rect 2710 1614 2716 1615
rect 2638 1604 2644 1605
rect 2638 1600 2639 1604
rect 2643 1600 2644 1604
rect 2638 1599 2644 1600
rect 2712 1596 2714 1614
rect 2768 1605 2770 1621
rect 2838 1619 2844 1620
rect 2838 1615 2839 1619
rect 2843 1615 2844 1619
rect 2838 1614 2844 1615
rect 2766 1604 2772 1605
rect 2766 1600 2767 1604
rect 2771 1600 2772 1604
rect 2766 1599 2772 1600
rect 2840 1596 2842 1614
rect 2896 1605 2898 1621
rect 2966 1619 2972 1620
rect 2966 1615 2967 1619
rect 2971 1615 2972 1619
rect 2966 1614 2972 1615
rect 2894 1604 2900 1605
rect 2894 1600 2895 1604
rect 2899 1600 2900 1604
rect 2894 1599 2900 1600
rect 2968 1596 2970 1614
rect 3016 1605 3018 1621
rect 3014 1604 3020 1605
rect 3014 1600 3015 1604
rect 3019 1600 3020 1604
rect 3014 1599 3020 1600
rect 3088 1596 3090 1634
rect 3135 1626 3139 1627
rect 3135 1621 3139 1622
rect 3136 1605 3138 1621
rect 3188 1620 3190 1662
rect 3214 1656 3220 1657
rect 3214 1652 3215 1656
rect 3219 1652 3220 1656
rect 3214 1651 3220 1652
rect 3216 1627 3218 1651
rect 3272 1640 3274 1810
rect 3342 1804 3348 1805
rect 3342 1800 3343 1804
rect 3347 1800 3348 1804
rect 3342 1799 3348 1800
rect 3344 1771 3346 1799
rect 3392 1788 3394 1942
rect 3432 1884 3434 2050
rect 3440 2032 3442 2194
rect 3464 2182 3466 2201
rect 3462 2181 3468 2182
rect 3462 2177 3463 2181
rect 3467 2177 3468 2181
rect 3462 2176 3468 2177
rect 3462 2164 3468 2165
rect 3462 2160 3463 2164
rect 3467 2160 3468 2164
rect 3462 2159 3468 2160
rect 3464 2135 3466 2159
rect 3463 2134 3467 2135
rect 3463 2129 3467 2130
rect 3464 2113 3466 2129
rect 3462 2112 3468 2113
rect 3462 2108 3463 2112
rect 3467 2108 3468 2112
rect 3462 2107 3468 2108
rect 3462 2095 3468 2096
rect 3462 2091 3463 2095
rect 3467 2091 3468 2095
rect 3462 2090 3468 2091
rect 3464 2063 3466 2090
rect 3463 2062 3467 2063
rect 3463 2057 3467 2058
rect 3464 2038 3466 2057
rect 3462 2037 3468 2038
rect 3462 2033 3463 2037
rect 3467 2033 3468 2037
rect 3462 2032 3468 2033
rect 3438 2031 3444 2032
rect 3438 2027 3439 2031
rect 3443 2027 3444 2031
rect 3438 2026 3444 2027
rect 3462 2020 3468 2021
rect 3462 2016 3463 2020
rect 3467 2016 3468 2020
rect 3462 2015 3468 2016
rect 3464 1983 3466 2015
rect 3463 1982 3467 1983
rect 3463 1977 3467 1978
rect 3464 1961 3466 1977
rect 3462 1960 3468 1961
rect 3462 1956 3463 1960
rect 3467 1956 3468 1960
rect 3462 1955 3468 1956
rect 3462 1943 3468 1944
rect 3462 1939 3463 1943
rect 3467 1939 3468 1943
rect 3462 1938 3468 1939
rect 3464 1915 3466 1938
rect 3463 1914 3467 1915
rect 3463 1909 3467 1910
rect 3446 1907 3452 1908
rect 3446 1903 3447 1907
rect 3451 1903 3452 1907
rect 3446 1902 3452 1903
rect 3430 1883 3436 1884
rect 3430 1879 3431 1883
rect 3435 1879 3436 1883
rect 3430 1878 3436 1879
rect 3390 1787 3396 1788
rect 3390 1783 3391 1787
rect 3395 1783 3396 1787
rect 3390 1782 3396 1783
rect 3343 1770 3347 1771
rect 3343 1765 3347 1766
rect 3367 1770 3371 1771
rect 3367 1765 3371 1766
rect 3368 1749 3370 1765
rect 3430 1763 3436 1764
rect 3430 1759 3431 1763
rect 3435 1759 3436 1763
rect 3430 1758 3436 1759
rect 3366 1748 3372 1749
rect 3366 1744 3367 1748
rect 3371 1744 3372 1748
rect 3366 1743 3372 1744
rect 3366 1729 3372 1730
rect 3366 1725 3367 1729
rect 3371 1725 3372 1729
rect 3366 1724 3372 1725
rect 3368 1699 3370 1724
rect 3367 1698 3371 1699
rect 3367 1693 3371 1694
rect 3368 1676 3370 1693
rect 3366 1675 3372 1676
rect 3366 1671 3367 1675
rect 3371 1671 3372 1675
rect 3432 1672 3434 1758
rect 3448 1740 3450 1902
rect 3464 1890 3466 1909
rect 3462 1889 3468 1890
rect 3462 1885 3463 1889
rect 3467 1885 3468 1889
rect 3462 1884 3468 1885
rect 3462 1872 3468 1873
rect 3462 1868 3463 1872
rect 3467 1868 3468 1872
rect 3462 1867 3468 1868
rect 3464 1847 3466 1867
rect 3463 1846 3467 1847
rect 3463 1841 3467 1842
rect 3464 1825 3466 1841
rect 3462 1824 3468 1825
rect 3462 1820 3463 1824
rect 3467 1820 3468 1824
rect 3462 1819 3468 1820
rect 3462 1807 3468 1808
rect 3462 1803 3463 1807
rect 3467 1803 3468 1807
rect 3462 1802 3468 1803
rect 3464 1771 3466 1802
rect 3463 1770 3467 1771
rect 3463 1765 3467 1766
rect 3464 1746 3466 1765
rect 3462 1745 3468 1746
rect 3462 1741 3463 1745
rect 3467 1741 3468 1745
rect 3462 1740 3468 1741
rect 3446 1739 3452 1740
rect 3446 1735 3447 1739
rect 3451 1735 3452 1739
rect 3446 1734 3452 1735
rect 3462 1728 3468 1729
rect 3462 1724 3463 1728
rect 3467 1724 3468 1728
rect 3462 1723 3468 1724
rect 3464 1699 3466 1723
rect 3463 1698 3467 1699
rect 3463 1693 3467 1694
rect 3464 1677 3466 1693
rect 3462 1676 3468 1677
rect 3462 1672 3463 1676
rect 3467 1672 3468 1676
rect 3366 1670 3372 1671
rect 3430 1671 3436 1672
rect 3462 1671 3468 1672
rect 3430 1667 3431 1671
rect 3435 1667 3436 1671
rect 3430 1666 3436 1667
rect 3462 1659 3468 1660
rect 3366 1656 3372 1657
rect 3366 1652 3367 1656
rect 3371 1652 3372 1656
rect 3462 1655 3463 1659
rect 3467 1655 3468 1659
rect 3462 1654 3468 1655
rect 3366 1651 3372 1652
rect 3270 1639 3276 1640
rect 3270 1635 3271 1639
rect 3275 1635 3276 1639
rect 3270 1634 3276 1635
rect 3368 1627 3370 1651
rect 3430 1639 3436 1640
rect 3430 1635 3431 1639
rect 3435 1635 3436 1639
rect 3430 1634 3436 1635
rect 3215 1626 3219 1627
rect 3215 1621 3219 1622
rect 3263 1626 3267 1627
rect 3263 1621 3267 1622
rect 3367 1626 3371 1627
rect 3367 1621 3371 1622
rect 3186 1619 3192 1620
rect 3186 1615 3187 1619
rect 3191 1615 3192 1619
rect 3186 1614 3192 1615
rect 3206 1619 3212 1620
rect 3206 1615 3207 1619
rect 3211 1615 3212 1619
rect 3206 1614 3212 1615
rect 3134 1604 3140 1605
rect 3134 1600 3135 1604
rect 3139 1600 3140 1604
rect 3134 1599 3140 1600
rect 3208 1596 3210 1614
rect 3264 1605 3266 1621
rect 3334 1619 3340 1620
rect 3334 1615 3335 1619
rect 3339 1615 3340 1619
rect 3334 1614 3340 1615
rect 3262 1604 3268 1605
rect 3262 1600 3263 1604
rect 3267 1600 3268 1604
rect 3262 1599 3268 1600
rect 3336 1596 3338 1614
rect 3368 1605 3370 1621
rect 3366 1604 3372 1605
rect 3366 1600 3367 1604
rect 3371 1600 3372 1604
rect 3366 1599 3372 1600
rect 3432 1596 3434 1634
rect 3464 1627 3466 1654
rect 3463 1626 3467 1627
rect 3463 1621 3467 1622
rect 3464 1602 3466 1621
rect 3462 1601 3468 1602
rect 3462 1597 3463 1601
rect 3467 1597 3468 1601
rect 3462 1596 3468 1597
rect 2710 1595 2716 1596
rect 2710 1591 2711 1595
rect 2715 1591 2716 1595
rect 2710 1590 2716 1591
rect 2838 1595 2844 1596
rect 2838 1591 2839 1595
rect 2843 1591 2844 1595
rect 2838 1590 2844 1591
rect 2966 1595 2972 1596
rect 2966 1591 2967 1595
rect 2971 1591 2972 1595
rect 2966 1590 2972 1591
rect 3086 1595 3092 1596
rect 3086 1591 3087 1595
rect 3091 1591 3092 1595
rect 3086 1590 3092 1591
rect 3206 1595 3212 1596
rect 3206 1591 3207 1595
rect 3211 1591 3212 1595
rect 3206 1590 3212 1591
rect 3334 1595 3340 1596
rect 3334 1591 3335 1595
rect 3339 1591 3340 1595
rect 3334 1590 3340 1591
rect 3430 1595 3436 1596
rect 3430 1591 3431 1595
rect 3435 1591 3436 1595
rect 3430 1590 3436 1591
rect 2638 1585 2644 1586
rect 2638 1581 2639 1585
rect 2643 1581 2644 1585
rect 2638 1580 2644 1581
rect 2766 1585 2772 1586
rect 2766 1581 2767 1585
rect 2771 1581 2772 1585
rect 2766 1580 2772 1581
rect 2894 1585 2900 1586
rect 2894 1581 2895 1585
rect 2899 1581 2900 1585
rect 2894 1580 2900 1581
rect 3014 1585 3020 1586
rect 3014 1581 3015 1585
rect 3019 1581 3020 1585
rect 3014 1580 3020 1581
rect 3134 1585 3140 1586
rect 3134 1581 3135 1585
rect 3139 1581 3140 1585
rect 3134 1580 3140 1581
rect 3262 1585 3268 1586
rect 3262 1581 3263 1585
rect 3267 1581 3268 1585
rect 3262 1580 3268 1581
rect 3366 1585 3372 1586
rect 3366 1581 3367 1585
rect 3371 1581 3372 1585
rect 3366 1580 3372 1581
rect 3462 1584 3468 1585
rect 3462 1580 3463 1584
rect 3467 1580 3468 1584
rect 2640 1555 2642 1580
rect 2768 1555 2770 1580
rect 2896 1555 2898 1580
rect 3016 1555 3018 1580
rect 3136 1555 3138 1580
rect 3264 1555 3266 1580
rect 3368 1555 3370 1580
rect 3462 1579 3468 1580
rect 3464 1555 3466 1579
rect 2599 1554 2603 1555
rect 2599 1549 2603 1550
rect 2639 1554 2643 1555
rect 2639 1549 2643 1550
rect 2735 1554 2739 1555
rect 2735 1549 2739 1550
rect 2767 1554 2771 1555
rect 2767 1549 2771 1550
rect 2871 1554 2875 1555
rect 2871 1549 2875 1550
rect 2895 1554 2899 1555
rect 2895 1549 2899 1550
rect 3007 1554 3011 1555
rect 3007 1549 3011 1550
rect 3015 1554 3019 1555
rect 3015 1549 3019 1550
rect 3135 1554 3139 1555
rect 3135 1549 3139 1550
rect 3143 1554 3147 1555
rect 3143 1549 3147 1550
rect 3263 1554 3267 1555
rect 3263 1549 3267 1550
rect 3367 1554 3371 1555
rect 3367 1549 3371 1550
rect 3463 1554 3467 1555
rect 3463 1549 3467 1550
rect 2600 1532 2602 1549
rect 2736 1532 2738 1549
rect 2872 1532 2874 1549
rect 3008 1532 3010 1549
rect 3144 1532 3146 1549
rect 3464 1533 3466 1549
rect 3462 1532 3468 1533
rect 2598 1531 2604 1532
rect 2598 1527 2599 1531
rect 2603 1527 2604 1531
rect 2598 1526 2604 1527
rect 2734 1531 2740 1532
rect 2734 1527 2735 1531
rect 2739 1527 2740 1531
rect 2734 1526 2740 1527
rect 2870 1531 2876 1532
rect 2870 1527 2871 1531
rect 2875 1527 2876 1531
rect 2870 1526 2876 1527
rect 3006 1531 3012 1532
rect 3006 1527 3007 1531
rect 3011 1527 3012 1531
rect 3006 1526 3012 1527
rect 3142 1531 3148 1532
rect 3142 1527 3143 1531
rect 3147 1527 3148 1531
rect 3462 1528 3463 1532
rect 3467 1528 3468 1532
rect 3462 1527 3468 1528
rect 3142 1526 3148 1527
rect 2558 1523 2564 1524
rect 2550 1519 2556 1520
rect 2550 1515 2551 1519
rect 2555 1515 2556 1519
rect 2558 1519 2559 1523
rect 2563 1519 2564 1523
rect 2558 1518 2564 1519
rect 2678 1523 2684 1524
rect 2678 1519 2679 1523
rect 2683 1519 2684 1523
rect 2678 1518 2684 1519
rect 2814 1523 2820 1524
rect 2814 1519 2815 1523
rect 2819 1519 2820 1523
rect 2814 1518 2820 1519
rect 2950 1523 2956 1524
rect 2950 1519 2951 1523
rect 2955 1519 2956 1523
rect 2950 1518 2956 1519
rect 3086 1523 3092 1524
rect 3086 1519 3087 1523
rect 3091 1519 3092 1523
rect 3086 1518 3092 1519
rect 2550 1514 2556 1515
rect 2454 1512 2460 1513
rect 2454 1508 2455 1512
rect 2459 1508 2460 1512
rect 2454 1507 2460 1508
rect 2438 1495 2444 1496
rect 2438 1491 2439 1495
rect 2443 1491 2444 1495
rect 2438 1490 2444 1491
rect 2456 1483 2458 1507
rect 1943 1482 1947 1483
rect 1943 1477 1947 1478
rect 1991 1482 1995 1483
rect 1991 1477 1995 1478
rect 2055 1482 2059 1483
rect 2055 1477 2059 1478
rect 2151 1482 2155 1483
rect 2151 1477 2155 1478
rect 2191 1482 2195 1483
rect 2191 1477 2195 1478
rect 2303 1482 2307 1483
rect 2303 1477 2307 1478
rect 2335 1482 2339 1483
rect 2335 1477 2339 1478
rect 2455 1482 2459 1483
rect 2455 1477 2459 1478
rect 2479 1482 2483 1483
rect 2479 1477 2483 1478
rect 1944 1461 1946 1477
rect 2056 1461 2058 1477
rect 2134 1475 2140 1476
rect 2134 1471 2135 1475
rect 2139 1471 2140 1475
rect 2134 1470 2140 1471
rect 1942 1460 1948 1461
rect 1942 1456 1943 1460
rect 1947 1456 1948 1460
rect 1942 1455 1948 1456
rect 2054 1460 2060 1461
rect 2054 1456 2055 1460
rect 2059 1456 2060 1460
rect 2054 1455 2060 1456
rect 2136 1452 2138 1470
rect 2192 1461 2194 1477
rect 2336 1461 2338 1477
rect 2390 1475 2396 1476
rect 2390 1471 2391 1475
rect 2395 1471 2396 1475
rect 2390 1470 2396 1471
rect 2406 1475 2412 1476
rect 2406 1471 2407 1475
rect 2411 1471 2412 1475
rect 2406 1470 2412 1471
rect 2190 1460 2196 1461
rect 2190 1456 2191 1460
rect 2195 1456 2196 1460
rect 2190 1455 2196 1456
rect 2334 1460 2340 1461
rect 2334 1456 2335 1460
rect 2339 1456 2340 1460
rect 2334 1455 2340 1456
rect 1894 1451 1900 1452
rect 1894 1447 1895 1451
rect 1899 1447 1900 1451
rect 1894 1446 1900 1447
rect 2134 1451 2140 1452
rect 2134 1447 2135 1451
rect 2139 1447 2140 1451
rect 2134 1446 2140 1447
rect 1942 1441 1948 1442
rect 1806 1440 1812 1441
rect 1470 1435 1476 1436
rect 1766 1437 1772 1438
rect 1766 1433 1767 1437
rect 1771 1433 1772 1437
rect 1806 1436 1807 1440
rect 1811 1436 1812 1440
rect 1942 1437 1943 1441
rect 1947 1437 1948 1441
rect 1942 1436 1948 1437
rect 2054 1441 2060 1442
rect 2054 1437 2055 1441
rect 2059 1437 2060 1441
rect 2054 1436 2060 1437
rect 2190 1441 2196 1442
rect 2190 1437 2191 1441
rect 2195 1437 2196 1441
rect 2190 1436 2196 1437
rect 2334 1441 2340 1442
rect 2334 1437 2335 1441
rect 2339 1437 2340 1441
rect 2334 1436 2340 1437
rect 1806 1435 1812 1436
rect 1766 1432 1772 1433
rect 998 1431 1004 1432
rect 998 1427 999 1431
rect 1003 1427 1004 1431
rect 998 1426 1004 1427
rect 1010 1431 1016 1432
rect 1010 1427 1011 1431
rect 1015 1427 1016 1431
rect 1010 1426 1016 1427
rect 1270 1431 1276 1432
rect 1270 1427 1271 1431
rect 1275 1427 1276 1431
rect 1270 1426 1276 1427
rect 1278 1431 1284 1432
rect 1278 1427 1279 1431
rect 1283 1427 1284 1431
rect 1278 1426 1284 1427
rect 1414 1431 1420 1432
rect 1414 1427 1415 1431
rect 1419 1427 1420 1431
rect 1414 1426 1420 1427
rect 1062 1421 1068 1422
rect 1062 1417 1063 1421
rect 1067 1417 1068 1421
rect 1062 1416 1068 1417
rect 1198 1421 1204 1422
rect 1198 1417 1199 1421
rect 1203 1417 1204 1421
rect 1198 1416 1204 1417
rect 1064 1395 1066 1416
rect 1200 1395 1202 1416
rect 1031 1394 1035 1395
rect 1031 1389 1035 1390
rect 1063 1394 1067 1395
rect 1063 1389 1067 1390
rect 1159 1394 1163 1395
rect 1159 1389 1163 1390
rect 1199 1394 1203 1395
rect 1199 1389 1203 1390
rect 1032 1372 1034 1389
rect 1160 1372 1162 1389
rect 1030 1371 1036 1372
rect 1030 1367 1031 1371
rect 1035 1367 1036 1371
rect 1030 1366 1036 1367
rect 1158 1371 1164 1372
rect 1158 1367 1159 1371
rect 1163 1367 1164 1371
rect 1158 1366 1164 1367
rect 974 1363 980 1364
rect 974 1359 975 1363
rect 979 1359 980 1363
rect 974 1358 980 1359
rect 982 1363 988 1364
rect 982 1359 983 1363
rect 987 1359 988 1363
rect 982 1358 988 1359
rect 1110 1363 1116 1364
rect 1110 1359 1111 1363
rect 1115 1359 1116 1363
rect 1110 1358 1116 1359
rect 902 1352 908 1353
rect 902 1348 903 1352
rect 907 1348 908 1352
rect 902 1347 908 1348
rect 846 1335 852 1336
rect 846 1331 847 1335
rect 851 1331 852 1335
rect 846 1330 852 1331
rect 904 1327 906 1347
rect 984 1336 986 1358
rect 1030 1352 1036 1353
rect 1030 1348 1031 1352
rect 1035 1348 1036 1352
rect 1030 1347 1036 1348
rect 982 1335 988 1336
rect 982 1331 983 1335
rect 987 1331 988 1335
rect 982 1330 988 1331
rect 1032 1327 1034 1347
rect 1112 1336 1114 1358
rect 1158 1352 1164 1353
rect 1158 1348 1159 1352
rect 1163 1348 1164 1352
rect 1158 1347 1164 1348
rect 1110 1335 1116 1336
rect 1110 1331 1111 1335
rect 1115 1331 1116 1335
rect 1110 1330 1116 1331
rect 1160 1327 1162 1347
rect 1272 1336 1274 1426
rect 1334 1421 1340 1422
rect 1334 1417 1335 1421
rect 1339 1417 1340 1421
rect 1334 1416 1340 1417
rect 1470 1421 1476 1422
rect 1470 1417 1471 1421
rect 1475 1417 1476 1421
rect 1470 1416 1476 1417
rect 1766 1420 1772 1421
rect 1766 1416 1767 1420
rect 1771 1416 1772 1420
rect 1336 1395 1338 1416
rect 1472 1395 1474 1416
rect 1766 1415 1772 1416
rect 1768 1395 1770 1415
rect 1808 1411 1810 1435
rect 1944 1411 1946 1436
rect 2056 1411 2058 1436
rect 2192 1411 2194 1436
rect 2336 1411 2338 1436
rect 1807 1410 1811 1411
rect 1807 1405 1811 1406
rect 1943 1410 1947 1411
rect 1943 1405 1947 1406
rect 2055 1410 2059 1411
rect 2055 1405 2059 1406
rect 2095 1410 2099 1411
rect 2095 1405 2099 1406
rect 2191 1410 2195 1411
rect 2191 1405 2195 1406
rect 2199 1410 2203 1411
rect 2199 1405 2203 1406
rect 2319 1410 2323 1411
rect 2319 1405 2323 1406
rect 2335 1410 2339 1411
rect 2335 1405 2339 1406
rect 1287 1394 1291 1395
rect 1287 1389 1291 1390
rect 1335 1394 1339 1395
rect 1335 1389 1339 1390
rect 1415 1394 1419 1395
rect 1415 1389 1419 1390
rect 1471 1394 1475 1395
rect 1471 1389 1475 1390
rect 1767 1394 1771 1395
rect 1767 1389 1771 1390
rect 1808 1389 1810 1405
rect 1288 1372 1290 1389
rect 1416 1372 1418 1389
rect 1768 1373 1770 1389
rect 1806 1388 1812 1389
rect 2096 1388 2098 1405
rect 2200 1388 2202 1405
rect 2320 1388 2322 1405
rect 1806 1384 1807 1388
rect 1811 1384 1812 1388
rect 1806 1383 1812 1384
rect 2094 1387 2100 1388
rect 2094 1383 2095 1387
rect 2099 1383 2100 1387
rect 2094 1382 2100 1383
rect 2198 1387 2204 1388
rect 2198 1383 2199 1387
rect 2203 1383 2204 1387
rect 2198 1382 2204 1383
rect 2318 1387 2324 1388
rect 2318 1383 2319 1387
rect 2323 1383 2324 1387
rect 2318 1382 2324 1383
rect 2392 1380 2394 1470
rect 2408 1452 2410 1470
rect 2480 1461 2482 1477
rect 2552 1476 2554 1514
rect 2598 1512 2604 1513
rect 2598 1508 2599 1512
rect 2603 1508 2604 1512
rect 2598 1507 2604 1508
rect 2600 1483 2602 1507
rect 2680 1496 2682 1518
rect 2734 1512 2740 1513
rect 2734 1508 2735 1512
rect 2739 1508 2740 1512
rect 2734 1507 2740 1508
rect 2678 1495 2684 1496
rect 2678 1491 2679 1495
rect 2683 1491 2684 1495
rect 2678 1490 2684 1491
rect 2736 1483 2738 1507
rect 2816 1496 2818 1518
rect 2870 1512 2876 1513
rect 2870 1508 2871 1512
rect 2875 1508 2876 1512
rect 2870 1507 2876 1508
rect 2814 1495 2820 1496
rect 2814 1491 2815 1495
rect 2819 1491 2820 1495
rect 2814 1490 2820 1491
rect 2872 1483 2874 1507
rect 2952 1496 2954 1518
rect 3006 1512 3012 1513
rect 3006 1508 3007 1512
rect 3011 1508 3012 1512
rect 3006 1507 3012 1508
rect 2950 1495 2956 1496
rect 2950 1491 2951 1495
rect 2955 1491 2956 1495
rect 2950 1490 2956 1491
rect 3008 1483 3010 1507
rect 3088 1496 3090 1518
rect 3462 1515 3468 1516
rect 3142 1512 3148 1513
rect 3142 1508 3143 1512
rect 3147 1508 3148 1512
rect 3462 1511 3463 1515
rect 3467 1511 3468 1515
rect 3462 1510 3468 1511
rect 3142 1507 3148 1508
rect 3086 1495 3092 1496
rect 3086 1491 3087 1495
rect 3091 1491 3092 1495
rect 3086 1490 3092 1491
rect 3144 1483 3146 1507
rect 3198 1495 3204 1496
rect 3198 1491 3199 1495
rect 3203 1491 3204 1495
rect 3198 1490 3204 1491
rect 2599 1482 2603 1483
rect 2599 1477 2603 1478
rect 2631 1482 2635 1483
rect 2631 1477 2635 1478
rect 2735 1482 2739 1483
rect 2735 1477 2739 1478
rect 2783 1482 2787 1483
rect 2783 1477 2787 1478
rect 2871 1482 2875 1483
rect 2871 1477 2875 1478
rect 2935 1482 2939 1483
rect 2935 1477 2939 1478
rect 3007 1482 3011 1483
rect 3007 1477 3011 1478
rect 3087 1482 3091 1483
rect 3087 1477 3091 1478
rect 3143 1482 3147 1483
rect 3143 1477 3147 1478
rect 2550 1475 2556 1476
rect 2550 1471 2551 1475
rect 2555 1471 2556 1475
rect 2550 1470 2556 1471
rect 2632 1461 2634 1477
rect 2784 1461 2786 1477
rect 2838 1475 2844 1476
rect 2838 1471 2839 1475
rect 2843 1471 2844 1475
rect 2838 1470 2844 1471
rect 2854 1475 2860 1476
rect 2854 1471 2855 1475
rect 2859 1471 2860 1475
rect 2854 1470 2860 1471
rect 2478 1460 2484 1461
rect 2478 1456 2479 1460
rect 2483 1456 2484 1460
rect 2478 1455 2484 1456
rect 2630 1460 2636 1461
rect 2630 1456 2631 1460
rect 2635 1456 2636 1460
rect 2630 1455 2636 1456
rect 2782 1460 2788 1461
rect 2782 1456 2783 1460
rect 2787 1456 2788 1460
rect 2782 1455 2788 1456
rect 2406 1451 2412 1452
rect 2406 1447 2407 1451
rect 2411 1447 2412 1451
rect 2406 1446 2412 1447
rect 2702 1451 2708 1452
rect 2702 1447 2703 1451
rect 2707 1447 2708 1451
rect 2702 1446 2708 1447
rect 2478 1441 2484 1442
rect 2478 1437 2479 1441
rect 2483 1437 2484 1441
rect 2478 1436 2484 1437
rect 2630 1441 2636 1442
rect 2630 1437 2631 1441
rect 2635 1437 2636 1441
rect 2630 1436 2636 1437
rect 2480 1411 2482 1436
rect 2632 1411 2634 1436
rect 2455 1410 2459 1411
rect 2455 1405 2459 1406
rect 2479 1410 2483 1411
rect 2479 1405 2483 1406
rect 2599 1410 2603 1411
rect 2599 1405 2603 1406
rect 2631 1410 2635 1411
rect 2631 1405 2635 1406
rect 2456 1388 2458 1405
rect 2600 1388 2602 1405
rect 2454 1387 2460 1388
rect 2454 1383 2455 1387
rect 2459 1383 2460 1387
rect 2454 1382 2460 1383
rect 2598 1387 2604 1388
rect 2598 1383 2599 1387
rect 2603 1383 2604 1387
rect 2598 1382 2604 1383
rect 2390 1379 2396 1380
rect 2166 1375 2172 1376
rect 1766 1372 1772 1373
rect 1286 1371 1292 1372
rect 1286 1367 1287 1371
rect 1291 1367 1292 1371
rect 1286 1366 1292 1367
rect 1414 1371 1420 1372
rect 1414 1367 1415 1371
rect 1419 1367 1420 1371
rect 1766 1368 1767 1372
rect 1771 1368 1772 1372
rect 1766 1367 1772 1368
rect 1806 1371 1812 1372
rect 1806 1367 1807 1371
rect 1811 1367 1812 1371
rect 2166 1371 2167 1375
rect 2171 1371 2172 1375
rect 2166 1370 2172 1371
rect 2270 1375 2276 1376
rect 2270 1371 2271 1375
rect 2275 1371 2276 1375
rect 2390 1375 2391 1379
rect 2395 1375 2396 1379
rect 2390 1374 2396 1375
rect 2426 1379 2432 1380
rect 2426 1375 2427 1379
rect 2431 1375 2432 1379
rect 2426 1374 2432 1375
rect 2534 1379 2540 1380
rect 2534 1375 2535 1379
rect 2539 1375 2540 1379
rect 2534 1374 2540 1375
rect 2270 1370 2276 1371
rect 1414 1366 1420 1367
rect 1806 1366 1812 1367
rect 2094 1368 2100 1369
rect 1366 1363 1372 1364
rect 1358 1359 1364 1360
rect 1358 1355 1359 1359
rect 1363 1355 1364 1359
rect 1366 1359 1367 1363
rect 1371 1359 1372 1363
rect 1366 1358 1372 1359
rect 1358 1354 1364 1355
rect 1286 1352 1292 1353
rect 1286 1348 1287 1352
rect 1291 1348 1292 1352
rect 1286 1347 1292 1348
rect 1254 1335 1260 1336
rect 1254 1331 1255 1335
rect 1259 1331 1260 1335
rect 1254 1330 1260 1331
rect 1270 1335 1276 1336
rect 1270 1331 1271 1335
rect 1275 1331 1276 1335
rect 1270 1330 1276 1331
rect 279 1326 283 1327
rect 279 1321 283 1322
rect 439 1326 443 1327
rect 439 1321 443 1322
rect 447 1326 451 1327
rect 558 1323 559 1327
rect 563 1323 564 1327
rect 558 1322 564 1323
rect 583 1326 587 1327
rect 447 1321 451 1322
rect 583 1321 587 1322
rect 607 1326 611 1327
rect 607 1321 611 1322
rect 719 1326 723 1327
rect 719 1321 723 1322
rect 759 1326 763 1327
rect 759 1321 763 1322
rect 847 1326 851 1327
rect 847 1321 851 1322
rect 903 1326 907 1327
rect 903 1321 907 1322
rect 967 1326 971 1327
rect 967 1321 971 1322
rect 1031 1326 1035 1327
rect 1031 1321 1035 1322
rect 1079 1326 1083 1327
rect 1079 1321 1083 1322
rect 1159 1326 1163 1327
rect 1159 1321 1163 1322
rect 1191 1326 1195 1327
rect 1191 1321 1195 1322
rect 206 1319 212 1320
rect 206 1315 207 1319
rect 211 1315 212 1319
rect 206 1314 212 1315
rect 198 1295 204 1296
rect 198 1291 199 1295
rect 203 1291 204 1295
rect 198 1290 204 1291
rect 134 1285 140 1286
rect 110 1284 116 1285
rect 110 1280 111 1284
rect 115 1280 116 1284
rect 134 1281 135 1285
rect 139 1281 140 1285
rect 134 1280 140 1281
rect 110 1279 116 1280
rect 112 1259 114 1279
rect 136 1259 138 1280
rect 111 1258 115 1259
rect 111 1253 115 1254
rect 135 1258 139 1259
rect 135 1253 139 1254
rect 112 1237 114 1253
rect 110 1236 116 1237
rect 136 1236 138 1253
rect 110 1232 111 1236
rect 115 1232 116 1236
rect 110 1231 116 1232
rect 134 1235 140 1236
rect 134 1231 135 1235
rect 139 1231 140 1235
rect 134 1230 140 1231
rect 208 1228 210 1314
rect 280 1305 282 1321
rect 350 1319 356 1320
rect 350 1315 351 1319
rect 355 1315 356 1319
rect 350 1314 356 1315
rect 278 1304 284 1305
rect 278 1300 279 1304
rect 283 1300 284 1304
rect 278 1299 284 1300
rect 352 1296 354 1314
rect 440 1305 442 1321
rect 510 1319 516 1320
rect 510 1315 511 1319
rect 515 1315 516 1319
rect 510 1314 516 1315
rect 438 1304 444 1305
rect 438 1300 439 1304
rect 443 1300 444 1304
rect 438 1299 444 1300
rect 512 1296 514 1314
rect 584 1305 586 1321
rect 686 1319 692 1320
rect 686 1315 687 1319
rect 691 1315 692 1319
rect 686 1314 692 1315
rect 582 1304 588 1305
rect 582 1300 583 1304
rect 587 1300 588 1304
rect 582 1299 588 1300
rect 350 1295 356 1296
rect 350 1291 351 1295
rect 355 1291 356 1295
rect 350 1290 356 1291
rect 510 1295 516 1296
rect 510 1291 511 1295
rect 515 1291 516 1295
rect 510 1290 516 1291
rect 654 1295 660 1296
rect 654 1291 655 1295
rect 659 1291 660 1295
rect 654 1290 660 1291
rect 278 1285 284 1286
rect 278 1281 279 1285
rect 283 1281 284 1285
rect 278 1280 284 1281
rect 438 1285 444 1286
rect 438 1281 439 1285
rect 443 1281 444 1285
rect 438 1280 444 1281
rect 582 1285 588 1286
rect 582 1281 583 1285
rect 587 1281 588 1285
rect 582 1280 588 1281
rect 280 1259 282 1280
rect 440 1259 442 1280
rect 584 1259 586 1280
rect 239 1258 243 1259
rect 239 1253 243 1254
rect 279 1258 283 1259
rect 279 1253 283 1254
rect 367 1258 371 1259
rect 367 1253 371 1254
rect 439 1258 443 1259
rect 439 1253 443 1254
rect 495 1258 499 1259
rect 495 1253 499 1254
rect 583 1258 587 1259
rect 583 1253 587 1254
rect 615 1258 619 1259
rect 615 1253 619 1254
rect 240 1236 242 1253
rect 368 1236 370 1253
rect 496 1236 498 1253
rect 616 1236 618 1253
rect 238 1235 244 1236
rect 238 1231 239 1235
rect 243 1231 244 1235
rect 238 1230 244 1231
rect 366 1235 372 1236
rect 366 1231 367 1235
rect 371 1231 372 1235
rect 366 1230 372 1231
rect 494 1235 500 1236
rect 494 1231 495 1235
rect 499 1231 500 1235
rect 494 1230 500 1231
rect 614 1235 620 1236
rect 614 1231 615 1235
rect 619 1231 620 1235
rect 614 1230 620 1231
rect 206 1227 212 1228
rect 206 1223 207 1227
rect 211 1223 212 1227
rect 206 1222 212 1223
rect 214 1227 220 1228
rect 214 1223 215 1227
rect 219 1223 220 1227
rect 214 1222 220 1223
rect 318 1227 324 1228
rect 318 1223 319 1227
rect 323 1223 324 1227
rect 318 1222 324 1223
rect 446 1227 452 1228
rect 446 1223 447 1227
rect 451 1223 452 1227
rect 446 1222 452 1223
rect 110 1219 116 1220
rect 110 1215 111 1219
rect 115 1215 116 1219
rect 110 1214 116 1215
rect 134 1216 140 1217
rect 112 1191 114 1214
rect 134 1212 135 1216
rect 139 1212 140 1216
rect 134 1211 140 1212
rect 136 1191 138 1211
rect 216 1200 218 1222
rect 238 1216 244 1217
rect 238 1212 239 1216
rect 243 1212 244 1216
rect 238 1211 244 1212
rect 214 1199 220 1200
rect 214 1195 215 1199
rect 219 1195 220 1199
rect 214 1194 220 1195
rect 240 1191 242 1211
rect 320 1200 322 1222
rect 366 1216 372 1217
rect 366 1212 367 1216
rect 371 1212 372 1216
rect 366 1211 372 1212
rect 318 1199 324 1200
rect 318 1195 319 1199
rect 323 1195 324 1199
rect 318 1194 324 1195
rect 368 1191 370 1211
rect 448 1200 450 1222
rect 494 1216 500 1217
rect 494 1212 495 1216
rect 499 1212 500 1216
rect 494 1211 500 1212
rect 614 1216 620 1217
rect 614 1212 615 1216
rect 619 1212 620 1216
rect 614 1211 620 1212
rect 446 1199 452 1200
rect 446 1195 447 1199
rect 451 1195 452 1199
rect 446 1194 452 1195
rect 496 1191 498 1211
rect 616 1191 618 1211
rect 656 1200 658 1290
rect 688 1228 690 1314
rect 720 1305 722 1321
rect 790 1319 796 1320
rect 790 1315 791 1319
rect 795 1315 796 1319
rect 790 1314 796 1315
rect 718 1304 724 1305
rect 718 1300 719 1304
rect 723 1300 724 1304
rect 718 1299 724 1300
rect 792 1296 794 1314
rect 848 1305 850 1321
rect 918 1319 924 1320
rect 918 1315 919 1319
rect 923 1315 924 1319
rect 918 1314 924 1315
rect 846 1304 852 1305
rect 846 1300 847 1304
rect 851 1300 852 1304
rect 846 1299 852 1300
rect 920 1296 922 1314
rect 968 1305 970 1321
rect 1038 1319 1044 1320
rect 1038 1315 1039 1319
rect 1043 1315 1044 1319
rect 1038 1314 1044 1315
rect 966 1304 972 1305
rect 966 1300 967 1304
rect 971 1300 972 1304
rect 966 1299 972 1300
rect 1040 1296 1042 1314
rect 1080 1305 1082 1321
rect 1192 1305 1194 1321
rect 1078 1304 1084 1305
rect 1078 1300 1079 1304
rect 1083 1300 1084 1304
rect 1078 1299 1084 1300
rect 1190 1304 1196 1305
rect 1190 1300 1191 1304
rect 1195 1300 1196 1304
rect 1190 1299 1196 1300
rect 1256 1296 1258 1330
rect 1288 1327 1290 1347
rect 1360 1336 1362 1354
rect 1358 1335 1364 1336
rect 1358 1331 1359 1335
rect 1363 1331 1364 1335
rect 1358 1330 1364 1331
rect 1287 1326 1291 1327
rect 1287 1321 1291 1322
rect 1311 1326 1315 1327
rect 1311 1321 1315 1322
rect 1298 1319 1304 1320
rect 1298 1315 1299 1319
rect 1303 1315 1304 1319
rect 1298 1314 1304 1315
rect 1300 1296 1302 1314
rect 1312 1305 1314 1321
rect 1368 1320 1370 1358
rect 1766 1355 1772 1356
rect 1414 1352 1420 1353
rect 1414 1348 1415 1352
rect 1419 1348 1420 1352
rect 1766 1351 1767 1355
rect 1771 1351 1772 1355
rect 1766 1350 1772 1351
rect 1414 1347 1420 1348
rect 1416 1327 1418 1347
rect 1768 1327 1770 1350
rect 1808 1343 1810 1366
rect 2094 1364 2095 1368
rect 2099 1364 2100 1368
rect 2094 1363 2100 1364
rect 2096 1343 2098 1363
rect 2168 1352 2170 1370
rect 2198 1368 2204 1369
rect 2198 1364 2199 1368
rect 2203 1364 2204 1368
rect 2198 1363 2204 1364
rect 2166 1351 2172 1352
rect 2166 1347 2167 1351
rect 2171 1347 2172 1351
rect 2166 1346 2172 1347
rect 2200 1343 2202 1363
rect 2272 1352 2274 1370
rect 2318 1368 2324 1369
rect 2318 1364 2319 1368
rect 2323 1364 2324 1368
rect 2318 1363 2324 1364
rect 2270 1351 2276 1352
rect 2270 1347 2271 1351
rect 2275 1347 2276 1351
rect 2270 1346 2276 1347
rect 2320 1343 2322 1363
rect 2428 1360 2430 1374
rect 2454 1368 2460 1369
rect 2454 1364 2455 1368
rect 2459 1364 2460 1368
rect 2454 1363 2460 1364
rect 2426 1359 2432 1360
rect 2426 1355 2427 1359
rect 2431 1355 2432 1359
rect 2426 1354 2432 1355
rect 2456 1343 2458 1363
rect 2536 1352 2538 1374
rect 2598 1368 2604 1369
rect 2598 1364 2599 1368
rect 2603 1364 2604 1368
rect 2598 1363 2604 1364
rect 2534 1351 2540 1352
rect 2534 1347 2535 1351
rect 2539 1347 2540 1351
rect 2534 1346 2540 1347
rect 2600 1343 2602 1363
rect 2704 1352 2706 1446
rect 2782 1441 2788 1442
rect 2782 1437 2783 1441
rect 2787 1437 2788 1441
rect 2782 1436 2788 1437
rect 2784 1411 2786 1436
rect 2743 1410 2747 1411
rect 2743 1405 2747 1406
rect 2783 1410 2787 1411
rect 2783 1405 2787 1406
rect 2744 1388 2746 1405
rect 2742 1387 2748 1388
rect 2742 1383 2743 1387
rect 2747 1383 2748 1387
rect 2742 1382 2748 1383
rect 2840 1380 2842 1470
rect 2856 1452 2858 1470
rect 2936 1461 2938 1477
rect 3088 1461 3090 1477
rect 3158 1475 3164 1476
rect 3158 1471 3159 1475
rect 3163 1471 3164 1475
rect 3158 1470 3164 1471
rect 2934 1460 2940 1461
rect 2934 1456 2935 1460
rect 2939 1456 2940 1460
rect 2934 1455 2940 1456
rect 3086 1460 3092 1461
rect 3086 1456 3087 1460
rect 3091 1456 3092 1460
rect 3086 1455 3092 1456
rect 3160 1452 3162 1470
rect 3200 1452 3202 1490
rect 3464 1483 3466 1510
rect 3239 1482 3243 1483
rect 3239 1477 3243 1478
rect 3463 1482 3467 1483
rect 3463 1477 3467 1478
rect 3240 1461 3242 1477
rect 3238 1460 3244 1461
rect 3238 1456 3239 1460
rect 3243 1456 3244 1460
rect 3464 1458 3466 1477
rect 3238 1455 3244 1456
rect 3462 1457 3468 1458
rect 3462 1453 3463 1457
rect 3467 1453 3468 1457
rect 3462 1452 3468 1453
rect 2854 1451 2860 1452
rect 2854 1447 2855 1451
rect 2859 1447 2860 1451
rect 2854 1446 2860 1447
rect 3158 1451 3164 1452
rect 3158 1447 3159 1451
rect 3163 1447 3164 1451
rect 3158 1446 3164 1447
rect 3198 1451 3204 1452
rect 3198 1447 3199 1451
rect 3203 1447 3204 1451
rect 3198 1446 3204 1447
rect 2934 1441 2940 1442
rect 2934 1437 2935 1441
rect 2939 1437 2940 1441
rect 2934 1436 2940 1437
rect 3086 1441 3092 1442
rect 3086 1437 3087 1441
rect 3091 1437 3092 1441
rect 3086 1436 3092 1437
rect 3238 1441 3244 1442
rect 3238 1437 3239 1441
rect 3243 1437 3244 1441
rect 3238 1436 3244 1437
rect 3462 1440 3468 1441
rect 3462 1436 3463 1440
rect 3467 1436 3468 1440
rect 2936 1411 2938 1436
rect 3088 1411 3090 1436
rect 3240 1411 3242 1436
rect 3462 1435 3468 1436
rect 3464 1411 3466 1435
rect 2887 1410 2891 1411
rect 2887 1405 2891 1406
rect 2935 1410 2939 1411
rect 2935 1405 2939 1406
rect 3031 1410 3035 1411
rect 3031 1405 3035 1406
rect 3087 1410 3091 1411
rect 3087 1405 3091 1406
rect 3175 1410 3179 1411
rect 3175 1405 3179 1406
rect 3239 1410 3243 1411
rect 3239 1405 3243 1406
rect 3327 1410 3331 1411
rect 3327 1405 3331 1406
rect 3463 1410 3467 1411
rect 3463 1405 3467 1406
rect 2888 1388 2890 1405
rect 3032 1388 3034 1405
rect 3176 1388 3178 1405
rect 3328 1388 3330 1405
rect 3464 1389 3466 1405
rect 3462 1388 3468 1389
rect 2886 1387 2892 1388
rect 2886 1383 2887 1387
rect 2891 1383 2892 1387
rect 2886 1382 2892 1383
rect 3030 1387 3036 1388
rect 3030 1383 3031 1387
rect 3035 1383 3036 1387
rect 3030 1382 3036 1383
rect 3174 1387 3180 1388
rect 3174 1383 3175 1387
rect 3179 1383 3180 1387
rect 3174 1382 3180 1383
rect 3326 1387 3332 1388
rect 3326 1383 3327 1387
rect 3331 1383 3332 1387
rect 3462 1384 3463 1388
rect 3467 1384 3468 1388
rect 3462 1383 3468 1384
rect 3326 1382 3332 1383
rect 2734 1379 2740 1380
rect 2734 1375 2735 1379
rect 2739 1375 2740 1379
rect 2734 1374 2740 1375
rect 2838 1379 2844 1380
rect 2838 1375 2839 1379
rect 2843 1375 2844 1379
rect 2838 1374 2844 1375
rect 2966 1379 2972 1380
rect 2966 1375 2967 1379
rect 2971 1375 2972 1379
rect 2966 1374 2972 1375
rect 3254 1379 3260 1380
rect 3254 1375 3255 1379
rect 3259 1375 3260 1379
rect 3254 1374 3260 1375
rect 2606 1351 2612 1352
rect 2606 1347 2607 1351
rect 2611 1347 2612 1351
rect 2606 1346 2612 1347
rect 2702 1351 2708 1352
rect 2702 1347 2703 1351
rect 2707 1347 2708 1351
rect 2702 1346 2708 1347
rect 1807 1342 1811 1343
rect 1807 1337 1811 1338
rect 2095 1342 2099 1343
rect 2095 1337 2099 1338
rect 2103 1342 2107 1343
rect 2103 1337 2107 1338
rect 2199 1342 2203 1343
rect 2199 1337 2203 1338
rect 2239 1342 2243 1343
rect 2239 1337 2243 1338
rect 2319 1342 2323 1343
rect 2319 1337 2323 1338
rect 2383 1342 2387 1343
rect 2383 1337 2387 1338
rect 2455 1342 2459 1343
rect 2455 1337 2459 1338
rect 2535 1342 2539 1343
rect 2535 1337 2539 1338
rect 2599 1342 2603 1343
rect 2599 1337 2603 1338
rect 1415 1326 1419 1327
rect 1415 1321 1419 1322
rect 1767 1326 1771 1327
rect 1767 1321 1771 1322
rect 1366 1319 1372 1320
rect 1366 1315 1367 1319
rect 1371 1315 1372 1319
rect 1366 1314 1372 1315
rect 1310 1304 1316 1305
rect 1310 1300 1311 1304
rect 1315 1300 1316 1304
rect 1768 1302 1770 1321
rect 1808 1318 1810 1337
rect 2104 1321 2106 1337
rect 2174 1335 2180 1336
rect 2174 1331 2175 1335
rect 2179 1331 2180 1335
rect 2174 1330 2180 1331
rect 2102 1320 2108 1321
rect 1806 1317 1812 1318
rect 1806 1313 1807 1317
rect 1811 1313 1812 1317
rect 2102 1316 2103 1320
rect 2107 1316 2108 1320
rect 2102 1315 2108 1316
rect 1806 1312 1812 1313
rect 2176 1312 2178 1330
rect 2240 1321 2242 1337
rect 2310 1335 2316 1336
rect 2310 1331 2311 1335
rect 2315 1331 2316 1335
rect 2310 1330 2316 1331
rect 2238 1320 2244 1321
rect 2238 1316 2239 1320
rect 2243 1316 2244 1320
rect 2238 1315 2244 1316
rect 2312 1312 2314 1330
rect 2322 1327 2328 1328
rect 2322 1323 2323 1327
rect 2327 1323 2328 1327
rect 2322 1322 2328 1323
rect 2174 1311 2180 1312
rect 2174 1307 2175 1311
rect 2179 1307 2180 1311
rect 2174 1306 2180 1307
rect 2310 1311 2316 1312
rect 2310 1307 2311 1311
rect 2315 1307 2316 1311
rect 2310 1306 2316 1307
rect 1310 1299 1316 1300
rect 1766 1301 1772 1302
rect 2102 1301 2108 1302
rect 1766 1297 1767 1301
rect 1771 1297 1772 1301
rect 1766 1296 1772 1297
rect 1806 1300 1812 1301
rect 1806 1296 1807 1300
rect 1811 1296 1812 1300
rect 2102 1297 2103 1301
rect 2107 1297 2108 1301
rect 2102 1296 2108 1297
rect 2238 1301 2244 1302
rect 2238 1297 2239 1301
rect 2243 1297 2244 1301
rect 2238 1296 2244 1297
rect 790 1295 796 1296
rect 790 1291 791 1295
rect 795 1291 796 1295
rect 790 1290 796 1291
rect 918 1295 924 1296
rect 918 1291 919 1295
rect 923 1291 924 1295
rect 918 1290 924 1291
rect 1038 1295 1044 1296
rect 1038 1291 1039 1295
rect 1043 1291 1044 1295
rect 1038 1290 1044 1291
rect 1046 1295 1052 1296
rect 1046 1291 1047 1295
rect 1051 1291 1052 1295
rect 1046 1290 1052 1291
rect 1254 1295 1260 1296
rect 1254 1291 1255 1295
rect 1259 1291 1260 1295
rect 1254 1290 1260 1291
rect 1298 1295 1304 1296
rect 1806 1295 1812 1296
rect 1298 1291 1299 1295
rect 1303 1291 1304 1295
rect 1298 1290 1304 1291
rect 718 1285 724 1286
rect 718 1281 719 1285
rect 723 1281 724 1285
rect 718 1280 724 1281
rect 846 1285 852 1286
rect 846 1281 847 1285
rect 851 1281 852 1285
rect 846 1280 852 1281
rect 966 1285 972 1286
rect 966 1281 967 1285
rect 971 1281 972 1285
rect 966 1280 972 1281
rect 720 1259 722 1280
rect 848 1259 850 1280
rect 968 1259 970 1280
rect 719 1258 723 1259
rect 719 1253 723 1254
rect 735 1258 739 1259
rect 735 1253 739 1254
rect 847 1258 851 1259
rect 847 1253 851 1254
rect 959 1258 963 1259
rect 959 1253 963 1254
rect 967 1258 971 1259
rect 967 1253 971 1254
rect 736 1236 738 1253
rect 848 1236 850 1253
rect 960 1236 962 1253
rect 734 1235 740 1236
rect 734 1231 735 1235
rect 739 1231 740 1235
rect 734 1230 740 1231
rect 846 1235 852 1236
rect 846 1231 847 1235
rect 851 1231 852 1235
rect 846 1230 852 1231
rect 958 1235 964 1236
rect 958 1231 959 1235
rect 963 1231 964 1235
rect 958 1230 964 1231
rect 686 1227 692 1228
rect 686 1223 687 1227
rect 691 1223 692 1227
rect 686 1222 692 1223
rect 806 1223 812 1224
rect 806 1219 807 1223
rect 811 1219 812 1223
rect 806 1218 812 1219
rect 918 1223 924 1224
rect 918 1219 919 1223
rect 923 1219 924 1223
rect 918 1218 924 1219
rect 1030 1223 1036 1224
rect 1030 1219 1031 1223
rect 1035 1219 1036 1223
rect 1030 1218 1036 1219
rect 734 1216 740 1217
rect 734 1212 735 1216
rect 739 1212 740 1216
rect 734 1211 740 1212
rect 622 1199 628 1200
rect 622 1195 623 1199
rect 627 1195 628 1199
rect 622 1194 628 1195
rect 654 1199 660 1200
rect 654 1195 655 1199
rect 659 1195 660 1199
rect 654 1194 660 1195
rect 111 1190 115 1191
rect 111 1185 115 1186
rect 135 1190 139 1191
rect 135 1185 139 1186
rect 239 1190 243 1191
rect 239 1185 243 1186
rect 367 1190 371 1191
rect 367 1185 371 1186
rect 375 1190 379 1191
rect 375 1185 379 1186
rect 495 1190 499 1191
rect 495 1185 499 1186
rect 511 1190 515 1191
rect 511 1185 515 1186
rect 615 1190 619 1191
rect 615 1185 619 1186
rect 112 1166 114 1185
rect 136 1169 138 1185
rect 182 1183 188 1184
rect 182 1179 183 1183
rect 187 1179 188 1183
rect 182 1178 188 1179
rect 206 1183 212 1184
rect 206 1179 207 1183
rect 211 1179 212 1183
rect 206 1178 212 1179
rect 134 1168 140 1169
rect 110 1165 116 1166
rect 110 1161 111 1165
rect 115 1161 116 1165
rect 134 1164 135 1168
rect 139 1164 140 1168
rect 134 1163 140 1164
rect 110 1160 116 1161
rect 134 1149 140 1150
rect 110 1148 116 1149
rect 110 1144 111 1148
rect 115 1144 116 1148
rect 134 1145 135 1149
rect 139 1145 140 1149
rect 134 1144 140 1145
rect 110 1143 116 1144
rect 112 1123 114 1143
rect 136 1123 138 1144
rect 111 1122 115 1123
rect 111 1117 115 1118
rect 135 1122 139 1123
rect 135 1117 139 1118
rect 112 1101 114 1117
rect 110 1100 116 1101
rect 110 1096 111 1100
rect 115 1096 116 1100
rect 110 1095 116 1096
rect 184 1092 186 1178
rect 208 1160 210 1178
rect 240 1169 242 1185
rect 310 1183 316 1184
rect 310 1179 311 1183
rect 315 1179 316 1183
rect 310 1178 316 1179
rect 238 1168 244 1169
rect 238 1164 239 1168
rect 243 1164 244 1168
rect 238 1163 244 1164
rect 312 1160 314 1178
rect 376 1169 378 1185
rect 446 1183 452 1184
rect 446 1179 447 1183
rect 451 1179 452 1183
rect 446 1178 452 1179
rect 374 1168 380 1169
rect 374 1164 375 1168
rect 379 1164 380 1168
rect 374 1163 380 1164
rect 448 1160 450 1178
rect 512 1169 514 1185
rect 582 1183 588 1184
rect 582 1179 583 1183
rect 587 1179 588 1183
rect 582 1178 588 1179
rect 510 1168 516 1169
rect 510 1164 511 1168
rect 515 1164 516 1168
rect 510 1163 516 1164
rect 584 1160 586 1178
rect 624 1160 626 1194
rect 736 1191 738 1211
rect 808 1200 810 1218
rect 846 1216 852 1217
rect 846 1212 847 1216
rect 851 1212 852 1216
rect 846 1211 852 1212
rect 806 1199 812 1200
rect 806 1195 807 1199
rect 811 1195 812 1199
rect 806 1194 812 1195
rect 848 1191 850 1211
rect 920 1200 922 1218
rect 958 1216 964 1217
rect 958 1212 959 1216
rect 963 1212 964 1216
rect 958 1211 964 1212
rect 918 1199 924 1200
rect 918 1195 919 1199
rect 923 1195 924 1199
rect 918 1194 924 1195
rect 960 1191 962 1211
rect 1032 1200 1034 1218
rect 1048 1208 1050 1290
rect 1078 1285 1084 1286
rect 1078 1281 1079 1285
rect 1083 1281 1084 1285
rect 1078 1280 1084 1281
rect 1190 1285 1196 1286
rect 1190 1281 1191 1285
rect 1195 1281 1196 1285
rect 1190 1280 1196 1281
rect 1310 1285 1316 1286
rect 1310 1281 1311 1285
rect 1315 1281 1316 1285
rect 1310 1280 1316 1281
rect 1766 1284 1772 1285
rect 1766 1280 1767 1284
rect 1771 1280 1772 1284
rect 1080 1259 1082 1280
rect 1192 1259 1194 1280
rect 1312 1259 1314 1280
rect 1766 1279 1772 1280
rect 1808 1279 1810 1295
rect 2104 1279 2106 1296
rect 2240 1279 2242 1296
rect 1768 1259 1770 1279
rect 1807 1278 1811 1279
rect 1807 1273 1811 1274
rect 1935 1278 1939 1279
rect 1935 1273 1939 1274
rect 2063 1278 2067 1279
rect 2063 1273 2067 1274
rect 2103 1278 2107 1279
rect 2103 1273 2107 1274
rect 2199 1278 2203 1279
rect 2199 1273 2203 1274
rect 2239 1278 2243 1279
rect 2239 1273 2243 1274
rect 1071 1258 1075 1259
rect 1071 1253 1075 1254
rect 1079 1258 1083 1259
rect 1079 1253 1083 1254
rect 1191 1258 1195 1259
rect 1191 1253 1195 1254
rect 1311 1258 1315 1259
rect 1311 1253 1315 1254
rect 1767 1258 1771 1259
rect 1808 1257 1810 1273
rect 1767 1253 1771 1254
rect 1806 1256 1812 1257
rect 1936 1256 1938 1273
rect 2064 1256 2066 1273
rect 2200 1256 2202 1273
rect 1072 1236 1074 1253
rect 1192 1236 1194 1253
rect 1768 1237 1770 1253
rect 1806 1252 1807 1256
rect 1811 1252 1812 1256
rect 1806 1251 1812 1252
rect 1934 1255 1940 1256
rect 1934 1251 1935 1255
rect 1939 1251 1940 1255
rect 1934 1250 1940 1251
rect 2062 1255 2068 1256
rect 2062 1251 2063 1255
rect 2067 1251 2068 1255
rect 2062 1250 2068 1251
rect 2198 1255 2204 1256
rect 2198 1251 2199 1255
rect 2203 1251 2204 1255
rect 2198 1250 2204 1251
rect 2324 1248 2326 1322
rect 2384 1321 2386 1337
rect 2536 1321 2538 1337
rect 2382 1320 2388 1321
rect 2382 1316 2383 1320
rect 2387 1316 2388 1320
rect 2382 1315 2388 1316
rect 2534 1320 2540 1321
rect 2534 1316 2535 1320
rect 2539 1316 2540 1320
rect 2534 1315 2540 1316
rect 2608 1312 2610 1346
rect 2687 1342 2691 1343
rect 2687 1337 2691 1338
rect 2688 1321 2690 1337
rect 2736 1336 2738 1374
rect 2742 1368 2748 1369
rect 2742 1364 2743 1368
rect 2747 1364 2748 1368
rect 2742 1363 2748 1364
rect 2886 1368 2892 1369
rect 2886 1364 2887 1368
rect 2891 1364 2892 1368
rect 2886 1363 2892 1364
rect 2744 1343 2746 1363
rect 2888 1343 2890 1363
rect 2968 1352 2970 1374
rect 3030 1368 3036 1369
rect 3030 1364 3031 1368
rect 3035 1364 3036 1368
rect 3030 1363 3036 1364
rect 3174 1368 3180 1369
rect 3174 1364 3175 1368
rect 3179 1364 3180 1368
rect 3174 1363 3180 1364
rect 2966 1351 2972 1352
rect 2966 1347 2967 1351
rect 2971 1347 2972 1351
rect 2966 1346 2972 1347
rect 3032 1343 3034 1363
rect 3176 1343 3178 1363
rect 3256 1352 3258 1374
rect 3462 1371 3468 1372
rect 3326 1368 3332 1369
rect 3326 1364 3327 1368
rect 3331 1364 3332 1368
rect 3462 1367 3463 1371
rect 3467 1367 3468 1371
rect 3462 1366 3468 1367
rect 3326 1363 3332 1364
rect 3254 1351 3260 1352
rect 3254 1347 3255 1351
rect 3259 1347 3260 1351
rect 3254 1346 3260 1347
rect 3328 1343 3330 1363
rect 3374 1351 3380 1352
rect 3374 1347 3375 1351
rect 3379 1347 3380 1351
rect 3374 1346 3380 1347
rect 2743 1342 2747 1343
rect 2743 1337 2747 1338
rect 2839 1342 2843 1343
rect 2839 1337 2843 1338
rect 2887 1342 2891 1343
rect 2887 1337 2891 1338
rect 2991 1342 2995 1343
rect 2991 1337 2995 1338
rect 3031 1342 3035 1343
rect 3031 1337 3035 1338
rect 3143 1342 3147 1343
rect 3143 1337 3147 1338
rect 3175 1342 3179 1343
rect 3175 1337 3179 1338
rect 3303 1342 3307 1343
rect 3303 1337 3307 1338
rect 3327 1342 3331 1343
rect 3327 1337 3331 1338
rect 2734 1335 2740 1336
rect 2734 1331 2735 1335
rect 2739 1331 2740 1335
rect 2734 1330 2740 1331
rect 2840 1321 2842 1337
rect 2910 1335 2916 1336
rect 2910 1331 2911 1335
rect 2915 1331 2916 1335
rect 2910 1330 2916 1331
rect 2686 1320 2692 1321
rect 2686 1316 2687 1320
rect 2691 1316 2692 1320
rect 2686 1315 2692 1316
rect 2838 1320 2844 1321
rect 2838 1316 2839 1320
rect 2843 1316 2844 1320
rect 2838 1315 2844 1316
rect 2912 1312 2914 1330
rect 2992 1321 2994 1337
rect 3062 1335 3068 1336
rect 3062 1331 3063 1335
rect 3067 1331 3068 1335
rect 3062 1330 3068 1331
rect 3054 1327 3060 1328
rect 3054 1323 3055 1327
rect 3059 1323 3060 1327
rect 3054 1322 3060 1323
rect 2990 1320 2996 1321
rect 2990 1316 2991 1320
rect 2995 1316 2996 1320
rect 2990 1315 2996 1316
rect 2606 1311 2612 1312
rect 2606 1307 2607 1311
rect 2611 1307 2612 1311
rect 2606 1306 2612 1307
rect 2750 1311 2756 1312
rect 2750 1307 2751 1311
rect 2755 1307 2756 1311
rect 2750 1306 2756 1307
rect 2910 1311 2916 1312
rect 2910 1307 2911 1311
rect 2915 1307 2916 1311
rect 2910 1306 2916 1307
rect 2382 1301 2388 1302
rect 2382 1297 2383 1301
rect 2387 1297 2388 1301
rect 2382 1296 2388 1297
rect 2534 1301 2540 1302
rect 2534 1297 2535 1301
rect 2539 1297 2540 1301
rect 2534 1296 2540 1297
rect 2686 1301 2692 1302
rect 2686 1297 2687 1301
rect 2691 1297 2692 1301
rect 2686 1296 2692 1297
rect 2384 1279 2386 1296
rect 2536 1279 2538 1296
rect 2688 1279 2690 1296
rect 2343 1278 2347 1279
rect 2343 1273 2347 1274
rect 2383 1278 2387 1279
rect 2383 1273 2387 1274
rect 2495 1278 2499 1279
rect 2495 1273 2499 1274
rect 2535 1278 2539 1279
rect 2535 1273 2539 1274
rect 2655 1278 2659 1279
rect 2655 1273 2659 1274
rect 2687 1278 2691 1279
rect 2687 1273 2691 1274
rect 2344 1256 2346 1273
rect 2496 1256 2498 1273
rect 2656 1256 2658 1273
rect 2342 1255 2348 1256
rect 2342 1251 2343 1255
rect 2347 1251 2348 1255
rect 2342 1250 2348 1251
rect 2494 1255 2500 1256
rect 2494 1251 2495 1255
rect 2499 1251 2500 1255
rect 2494 1250 2500 1251
rect 2654 1255 2660 1256
rect 2654 1251 2655 1255
rect 2659 1251 2660 1255
rect 2654 1250 2660 1251
rect 2322 1247 2328 1248
rect 2006 1243 2012 1244
rect 1806 1239 1812 1240
rect 1766 1236 1772 1237
rect 1070 1235 1076 1236
rect 1070 1231 1071 1235
rect 1075 1231 1076 1235
rect 1070 1230 1076 1231
rect 1190 1235 1196 1236
rect 1190 1231 1191 1235
rect 1195 1231 1196 1235
rect 1766 1232 1767 1236
rect 1771 1232 1772 1236
rect 1806 1235 1807 1239
rect 1811 1235 1812 1239
rect 2006 1239 2007 1243
rect 2011 1239 2012 1243
rect 2006 1238 2012 1239
rect 2134 1243 2140 1244
rect 2134 1239 2135 1243
rect 2139 1239 2140 1243
rect 2134 1238 2140 1239
rect 2270 1243 2276 1244
rect 2270 1239 2271 1243
rect 2275 1239 2276 1243
rect 2322 1243 2323 1247
rect 2327 1243 2328 1247
rect 2574 1247 2580 1248
rect 2322 1242 2328 1243
rect 2566 1243 2572 1244
rect 2270 1238 2276 1239
rect 2566 1239 2567 1243
rect 2571 1239 2572 1243
rect 2574 1243 2575 1247
rect 2579 1243 2580 1247
rect 2574 1242 2580 1243
rect 2566 1238 2572 1239
rect 1806 1234 1812 1235
rect 1934 1236 1940 1237
rect 1766 1231 1772 1232
rect 1190 1230 1196 1231
rect 1150 1227 1156 1228
rect 1142 1223 1148 1224
rect 1142 1219 1143 1223
rect 1147 1219 1148 1223
rect 1150 1223 1151 1227
rect 1155 1223 1156 1227
rect 1150 1222 1156 1223
rect 1142 1218 1148 1219
rect 1070 1216 1076 1217
rect 1070 1212 1071 1216
rect 1075 1212 1076 1216
rect 1070 1211 1076 1212
rect 1046 1207 1052 1208
rect 1046 1203 1047 1207
rect 1051 1203 1052 1207
rect 1046 1202 1052 1203
rect 1030 1199 1036 1200
rect 1030 1195 1031 1199
rect 1035 1195 1036 1199
rect 1030 1194 1036 1195
rect 1072 1191 1074 1211
rect 1144 1200 1146 1218
rect 1142 1199 1148 1200
rect 1142 1195 1143 1199
rect 1147 1195 1148 1199
rect 1142 1194 1148 1195
rect 1152 1192 1154 1222
rect 1766 1219 1772 1220
rect 1190 1216 1196 1217
rect 1190 1212 1191 1216
rect 1195 1212 1196 1216
rect 1766 1215 1767 1219
rect 1771 1215 1772 1219
rect 1808 1215 1810 1234
rect 1934 1232 1935 1236
rect 1939 1232 1940 1236
rect 1934 1231 1940 1232
rect 1936 1215 1938 1231
rect 2008 1220 2010 1238
rect 2062 1236 2068 1237
rect 2062 1232 2063 1236
rect 2067 1232 2068 1236
rect 2062 1231 2068 1232
rect 2006 1219 2012 1220
rect 2006 1215 2007 1219
rect 2011 1215 2012 1219
rect 2064 1215 2066 1231
rect 2136 1220 2138 1238
rect 2198 1236 2204 1237
rect 2198 1232 2199 1236
rect 2203 1232 2204 1236
rect 2198 1231 2204 1232
rect 2134 1219 2140 1220
rect 2134 1215 2135 1219
rect 2139 1215 2140 1219
rect 2200 1215 2202 1231
rect 2272 1220 2274 1238
rect 2342 1236 2348 1237
rect 2342 1232 2343 1236
rect 2347 1232 2348 1236
rect 2342 1231 2348 1232
rect 2494 1236 2500 1237
rect 2494 1232 2495 1236
rect 2499 1232 2500 1236
rect 2494 1231 2500 1232
rect 2310 1227 2316 1228
rect 2310 1223 2311 1227
rect 2315 1223 2316 1227
rect 2310 1222 2316 1223
rect 2270 1219 2276 1220
rect 2270 1215 2271 1219
rect 2275 1215 2276 1219
rect 1766 1214 1772 1215
rect 1807 1214 1811 1215
rect 1190 1211 1196 1212
rect 1150 1191 1156 1192
rect 1192 1191 1194 1211
rect 1768 1191 1770 1214
rect 1807 1209 1811 1210
rect 1831 1214 1835 1215
rect 1831 1209 1835 1210
rect 1935 1214 1939 1215
rect 2006 1214 2012 1215
rect 2063 1214 2067 1215
rect 1935 1209 1939 1210
rect 2063 1209 2067 1210
rect 2079 1214 2083 1215
rect 2134 1214 2140 1215
rect 2199 1214 2203 1215
rect 2079 1209 2083 1210
rect 2199 1209 2203 1210
rect 2231 1214 2235 1215
rect 2270 1214 2276 1215
rect 2231 1209 2235 1210
rect 655 1190 659 1191
rect 655 1185 659 1186
rect 735 1190 739 1191
rect 735 1185 739 1186
rect 791 1190 795 1191
rect 791 1185 795 1186
rect 847 1190 851 1191
rect 847 1185 851 1186
rect 927 1190 931 1191
rect 927 1185 931 1186
rect 959 1190 963 1191
rect 959 1185 963 1186
rect 1063 1190 1067 1191
rect 1063 1185 1067 1186
rect 1071 1190 1075 1191
rect 1150 1187 1151 1191
rect 1155 1187 1156 1191
rect 1150 1186 1156 1187
rect 1191 1190 1195 1191
rect 1071 1185 1075 1186
rect 1191 1185 1195 1186
rect 1199 1190 1203 1191
rect 1199 1185 1203 1186
rect 1335 1190 1339 1191
rect 1335 1185 1339 1186
rect 1767 1190 1771 1191
rect 1808 1190 1810 1209
rect 1832 1193 1834 1209
rect 1926 1207 1932 1208
rect 1926 1203 1927 1207
rect 1931 1203 1932 1207
rect 1926 1202 1932 1203
rect 1830 1192 1836 1193
rect 1767 1185 1771 1186
rect 1806 1189 1812 1190
rect 1806 1185 1807 1189
rect 1811 1185 1812 1189
rect 1830 1188 1831 1192
rect 1835 1188 1836 1192
rect 1830 1187 1836 1188
rect 656 1169 658 1185
rect 792 1169 794 1185
rect 862 1183 868 1184
rect 862 1179 863 1183
rect 867 1179 868 1183
rect 862 1178 868 1179
rect 654 1168 660 1169
rect 654 1164 655 1168
rect 659 1164 660 1168
rect 654 1163 660 1164
rect 790 1168 796 1169
rect 790 1164 791 1168
rect 795 1164 796 1168
rect 790 1163 796 1164
rect 864 1160 866 1178
rect 928 1169 930 1185
rect 998 1183 1004 1184
rect 998 1179 999 1183
rect 1003 1179 1004 1183
rect 998 1178 1004 1179
rect 926 1168 932 1169
rect 926 1164 927 1168
rect 931 1164 932 1168
rect 926 1163 932 1164
rect 1000 1160 1002 1178
rect 1064 1169 1066 1185
rect 1134 1183 1140 1184
rect 1134 1179 1135 1183
rect 1139 1179 1140 1183
rect 1134 1178 1140 1179
rect 1062 1168 1068 1169
rect 1062 1164 1063 1168
rect 1067 1164 1068 1168
rect 1062 1163 1068 1164
rect 1136 1160 1138 1178
rect 1200 1169 1202 1185
rect 1270 1183 1276 1184
rect 1270 1179 1271 1183
rect 1275 1179 1276 1183
rect 1270 1178 1276 1179
rect 1198 1168 1204 1169
rect 1198 1164 1199 1168
rect 1203 1164 1204 1168
rect 1198 1163 1204 1164
rect 1272 1160 1274 1178
rect 1336 1169 1338 1185
rect 1334 1168 1340 1169
rect 1334 1164 1335 1168
rect 1339 1164 1340 1168
rect 1768 1166 1770 1185
rect 1806 1184 1812 1185
rect 1830 1173 1836 1174
rect 1806 1172 1812 1173
rect 1806 1168 1807 1172
rect 1811 1168 1812 1172
rect 1830 1169 1831 1173
rect 1835 1169 1836 1173
rect 1830 1168 1836 1169
rect 1806 1167 1812 1168
rect 1334 1163 1340 1164
rect 1766 1165 1772 1166
rect 1766 1161 1767 1165
rect 1771 1161 1772 1165
rect 1766 1160 1772 1161
rect 206 1159 212 1160
rect 206 1155 207 1159
rect 211 1155 212 1159
rect 206 1154 212 1155
rect 310 1159 316 1160
rect 310 1155 311 1159
rect 315 1155 316 1159
rect 310 1154 316 1155
rect 446 1159 452 1160
rect 446 1155 447 1159
rect 451 1155 452 1159
rect 446 1154 452 1155
rect 582 1159 588 1160
rect 582 1155 583 1159
rect 587 1155 588 1159
rect 582 1154 588 1155
rect 622 1159 628 1160
rect 622 1155 623 1159
rect 627 1155 628 1159
rect 622 1154 628 1155
rect 862 1159 868 1160
rect 862 1155 863 1159
rect 867 1155 868 1159
rect 862 1154 868 1155
rect 998 1159 1004 1160
rect 998 1155 999 1159
rect 1003 1155 1004 1159
rect 998 1154 1004 1155
rect 1134 1159 1140 1160
rect 1134 1155 1135 1159
rect 1139 1155 1140 1159
rect 1134 1154 1140 1155
rect 1270 1159 1276 1160
rect 1270 1155 1271 1159
rect 1275 1155 1276 1159
rect 1270 1154 1276 1155
rect 1278 1159 1284 1160
rect 1278 1155 1279 1159
rect 1283 1155 1284 1159
rect 1278 1154 1284 1155
rect 238 1149 244 1150
rect 238 1145 239 1149
rect 243 1145 244 1149
rect 238 1144 244 1145
rect 374 1149 380 1150
rect 374 1145 375 1149
rect 379 1145 380 1149
rect 374 1144 380 1145
rect 510 1149 516 1150
rect 510 1145 511 1149
rect 515 1145 516 1149
rect 510 1144 516 1145
rect 654 1149 660 1150
rect 654 1145 655 1149
rect 659 1145 660 1149
rect 654 1144 660 1145
rect 790 1149 796 1150
rect 790 1145 791 1149
rect 795 1145 796 1149
rect 790 1144 796 1145
rect 926 1149 932 1150
rect 926 1145 927 1149
rect 931 1145 932 1149
rect 926 1144 932 1145
rect 1062 1149 1068 1150
rect 1062 1145 1063 1149
rect 1067 1145 1068 1149
rect 1062 1144 1068 1145
rect 1198 1149 1204 1150
rect 1198 1145 1199 1149
rect 1203 1145 1204 1149
rect 1198 1144 1204 1145
rect 240 1123 242 1144
rect 376 1123 378 1144
rect 512 1123 514 1144
rect 656 1123 658 1144
rect 792 1123 794 1144
rect 928 1123 930 1144
rect 1064 1123 1066 1144
rect 1200 1123 1202 1144
rect 191 1122 195 1123
rect 191 1117 195 1118
rect 239 1122 243 1123
rect 239 1117 243 1118
rect 335 1122 339 1123
rect 335 1117 339 1118
rect 375 1122 379 1123
rect 375 1117 379 1118
rect 495 1122 499 1123
rect 495 1117 499 1118
rect 511 1122 515 1123
rect 511 1117 515 1118
rect 655 1122 659 1123
rect 655 1117 659 1118
rect 791 1122 795 1123
rect 791 1117 795 1118
rect 815 1122 819 1123
rect 815 1117 819 1118
rect 927 1122 931 1123
rect 927 1117 931 1118
rect 967 1122 971 1123
rect 967 1117 971 1118
rect 1063 1122 1067 1123
rect 1063 1117 1067 1118
rect 1119 1122 1123 1123
rect 1119 1117 1123 1118
rect 1199 1122 1203 1123
rect 1199 1117 1203 1118
rect 1263 1122 1267 1123
rect 1263 1117 1267 1118
rect 192 1100 194 1117
rect 336 1100 338 1117
rect 496 1100 498 1117
rect 656 1100 658 1117
rect 816 1100 818 1117
rect 968 1100 970 1117
rect 1120 1100 1122 1117
rect 1264 1100 1266 1117
rect 190 1099 196 1100
rect 190 1095 191 1099
rect 195 1095 196 1099
rect 190 1094 196 1095
rect 334 1099 340 1100
rect 334 1095 335 1099
rect 339 1095 340 1099
rect 334 1094 340 1095
rect 494 1099 500 1100
rect 494 1095 495 1099
rect 499 1095 500 1099
rect 494 1094 500 1095
rect 654 1099 660 1100
rect 654 1095 655 1099
rect 659 1095 660 1099
rect 654 1094 660 1095
rect 814 1099 820 1100
rect 814 1095 815 1099
rect 819 1095 820 1099
rect 814 1094 820 1095
rect 966 1099 972 1100
rect 966 1095 967 1099
rect 971 1095 972 1099
rect 966 1094 972 1095
rect 1118 1099 1124 1100
rect 1118 1095 1119 1099
rect 1123 1095 1124 1099
rect 1118 1094 1124 1095
rect 1262 1099 1268 1100
rect 1262 1095 1263 1099
rect 1267 1095 1268 1099
rect 1262 1094 1268 1095
rect 182 1091 188 1092
rect 182 1087 183 1091
rect 187 1087 188 1091
rect 182 1086 188 1087
rect 270 1091 276 1092
rect 270 1087 271 1091
rect 275 1087 276 1091
rect 270 1086 276 1087
rect 414 1091 420 1092
rect 414 1087 415 1091
rect 419 1087 420 1091
rect 766 1091 772 1092
rect 414 1086 420 1087
rect 726 1087 732 1088
rect 110 1083 116 1084
rect 110 1079 111 1083
rect 115 1079 116 1083
rect 110 1078 116 1079
rect 190 1080 196 1081
rect 112 1051 114 1078
rect 190 1076 191 1080
rect 195 1076 196 1080
rect 190 1075 196 1076
rect 192 1051 194 1075
rect 272 1064 274 1086
rect 334 1080 340 1081
rect 334 1076 335 1080
rect 339 1076 340 1080
rect 334 1075 340 1076
rect 270 1063 276 1064
rect 270 1059 271 1063
rect 275 1059 276 1063
rect 270 1058 276 1059
rect 336 1051 338 1075
rect 416 1064 418 1086
rect 726 1083 727 1087
rect 731 1083 732 1087
rect 766 1087 767 1091
rect 771 1087 772 1091
rect 766 1086 772 1087
rect 1038 1087 1044 1088
rect 726 1082 732 1083
rect 494 1080 500 1081
rect 494 1076 495 1080
rect 499 1076 500 1080
rect 494 1075 500 1076
rect 654 1080 660 1081
rect 654 1076 655 1080
rect 659 1076 660 1080
rect 654 1075 660 1076
rect 414 1063 420 1064
rect 414 1059 415 1063
rect 419 1059 420 1063
rect 414 1058 420 1059
rect 398 1051 404 1052
rect 496 1051 498 1075
rect 656 1051 658 1075
rect 728 1064 730 1082
rect 768 1072 770 1086
rect 1038 1083 1039 1087
rect 1043 1083 1044 1087
rect 1038 1082 1044 1083
rect 1190 1087 1196 1088
rect 1190 1083 1191 1087
rect 1195 1083 1196 1087
rect 1190 1082 1196 1083
rect 814 1080 820 1081
rect 814 1076 815 1080
rect 819 1076 820 1080
rect 814 1075 820 1076
rect 966 1080 972 1081
rect 966 1076 967 1080
rect 971 1076 972 1080
rect 966 1075 972 1076
rect 766 1071 772 1072
rect 766 1067 767 1071
rect 771 1067 772 1071
rect 766 1066 772 1067
rect 678 1063 684 1064
rect 678 1059 679 1063
rect 683 1059 684 1063
rect 678 1058 684 1059
rect 726 1063 732 1064
rect 726 1059 727 1063
rect 731 1059 732 1063
rect 726 1058 732 1059
rect 111 1050 115 1051
rect 111 1045 115 1046
rect 191 1050 195 1051
rect 191 1045 195 1046
rect 327 1050 331 1051
rect 327 1045 331 1046
rect 335 1050 339 1051
rect 398 1047 399 1051
rect 403 1047 404 1051
rect 398 1046 404 1047
rect 463 1050 467 1051
rect 335 1045 339 1046
rect 112 1026 114 1045
rect 328 1029 330 1045
rect 326 1028 332 1029
rect 110 1025 116 1026
rect 110 1021 111 1025
rect 115 1021 116 1025
rect 326 1024 327 1028
rect 331 1024 332 1028
rect 326 1023 332 1024
rect 110 1020 116 1021
rect 400 1020 402 1046
rect 463 1045 467 1046
rect 495 1050 499 1051
rect 495 1045 499 1046
rect 607 1050 611 1051
rect 607 1045 611 1046
rect 655 1050 659 1051
rect 655 1045 659 1046
rect 464 1029 466 1045
rect 534 1043 540 1044
rect 534 1039 535 1043
rect 539 1039 540 1043
rect 534 1038 540 1039
rect 462 1028 468 1029
rect 462 1024 463 1028
rect 467 1024 468 1028
rect 462 1023 468 1024
rect 536 1020 538 1038
rect 608 1029 610 1045
rect 606 1028 612 1029
rect 606 1024 607 1028
rect 611 1024 612 1028
rect 606 1023 612 1024
rect 680 1020 682 1058
rect 816 1051 818 1075
rect 968 1051 970 1075
rect 1040 1064 1042 1082
rect 1118 1080 1124 1081
rect 1118 1076 1119 1080
rect 1123 1076 1124 1080
rect 1118 1075 1124 1076
rect 1038 1063 1044 1064
rect 1038 1059 1039 1063
rect 1043 1059 1044 1063
rect 1038 1058 1044 1059
rect 1120 1051 1122 1075
rect 1192 1064 1194 1082
rect 1262 1080 1268 1081
rect 1262 1076 1263 1080
rect 1267 1076 1268 1080
rect 1262 1075 1268 1076
rect 1190 1063 1196 1064
rect 1190 1059 1191 1063
rect 1195 1059 1196 1063
rect 1190 1058 1196 1059
rect 1264 1051 1266 1075
rect 1280 1072 1282 1154
rect 1334 1149 1340 1150
rect 1334 1145 1335 1149
rect 1339 1145 1340 1149
rect 1334 1144 1340 1145
rect 1766 1148 1772 1149
rect 1766 1144 1767 1148
rect 1771 1144 1772 1148
rect 1336 1123 1338 1144
rect 1766 1143 1772 1144
rect 1768 1123 1770 1143
rect 1808 1139 1810 1167
rect 1832 1139 1834 1168
rect 1807 1138 1811 1139
rect 1807 1133 1811 1134
rect 1831 1138 1835 1139
rect 1831 1133 1835 1134
rect 1863 1138 1867 1139
rect 1863 1133 1867 1134
rect 1335 1122 1339 1123
rect 1335 1117 1339 1118
rect 1407 1122 1411 1123
rect 1407 1117 1411 1118
rect 1559 1122 1563 1123
rect 1559 1117 1563 1118
rect 1767 1122 1771 1123
rect 1767 1117 1771 1118
rect 1808 1117 1810 1133
rect 1408 1100 1410 1117
rect 1560 1100 1562 1117
rect 1768 1101 1770 1117
rect 1806 1116 1812 1117
rect 1864 1116 1866 1133
rect 1806 1112 1807 1116
rect 1811 1112 1812 1116
rect 1806 1111 1812 1112
rect 1862 1115 1868 1116
rect 1862 1111 1863 1115
rect 1867 1111 1868 1115
rect 1928 1112 1930 1202
rect 1936 1193 1938 1209
rect 2006 1207 2012 1208
rect 2006 1203 2007 1207
rect 2011 1203 2012 1207
rect 2006 1202 2012 1203
rect 1934 1192 1940 1193
rect 1934 1188 1935 1192
rect 1939 1188 1940 1192
rect 1934 1187 1940 1188
rect 2008 1184 2010 1202
rect 2080 1193 2082 1209
rect 2150 1207 2156 1208
rect 2150 1203 2151 1207
rect 2155 1203 2156 1207
rect 2150 1202 2156 1203
rect 2078 1192 2084 1193
rect 2078 1188 2079 1192
rect 2083 1188 2084 1192
rect 2078 1187 2084 1188
rect 2152 1184 2154 1202
rect 2232 1193 2234 1209
rect 2302 1207 2308 1208
rect 2302 1203 2303 1207
rect 2307 1203 2308 1207
rect 2302 1202 2308 1203
rect 2230 1192 2236 1193
rect 2230 1188 2231 1192
rect 2235 1188 2236 1192
rect 2230 1187 2236 1188
rect 2304 1184 2306 1202
rect 2312 1184 2314 1222
rect 2344 1215 2346 1231
rect 2496 1215 2498 1231
rect 2343 1214 2347 1215
rect 2343 1209 2347 1210
rect 2391 1214 2395 1215
rect 2391 1209 2395 1210
rect 2495 1214 2499 1215
rect 2495 1209 2499 1210
rect 2543 1214 2547 1215
rect 2543 1209 2547 1210
rect 2392 1193 2394 1209
rect 2544 1193 2546 1209
rect 2568 1208 2570 1238
rect 2576 1220 2578 1242
rect 2654 1236 2660 1237
rect 2654 1232 2655 1236
rect 2659 1232 2660 1236
rect 2654 1231 2660 1232
rect 2574 1219 2580 1220
rect 2574 1215 2575 1219
rect 2579 1215 2580 1219
rect 2656 1215 2658 1231
rect 2752 1220 2754 1306
rect 2838 1301 2844 1302
rect 2838 1297 2839 1301
rect 2843 1297 2844 1301
rect 2838 1296 2844 1297
rect 2990 1301 2996 1302
rect 2990 1297 2991 1301
rect 2995 1297 2996 1301
rect 2990 1296 2996 1297
rect 2840 1279 2842 1296
rect 2992 1279 2994 1296
rect 2815 1278 2819 1279
rect 2815 1273 2819 1274
rect 2839 1278 2843 1279
rect 2839 1273 2843 1274
rect 2975 1278 2979 1279
rect 2975 1273 2979 1274
rect 2991 1278 2995 1279
rect 2991 1273 2995 1274
rect 2816 1256 2818 1273
rect 2976 1256 2978 1273
rect 2814 1255 2820 1256
rect 2814 1251 2815 1255
rect 2819 1251 2820 1255
rect 2814 1250 2820 1251
rect 2974 1255 2980 1256
rect 2974 1251 2975 1255
rect 2979 1251 2980 1255
rect 2974 1250 2980 1251
rect 3056 1248 3058 1322
rect 3064 1312 3066 1330
rect 3144 1321 3146 1337
rect 3214 1335 3220 1336
rect 3214 1331 3215 1335
rect 3219 1331 3220 1335
rect 3214 1330 3220 1331
rect 3142 1320 3148 1321
rect 3142 1316 3143 1320
rect 3147 1316 3148 1320
rect 3142 1315 3148 1316
rect 3216 1312 3218 1330
rect 3304 1321 3306 1337
rect 3302 1320 3308 1321
rect 3302 1316 3303 1320
rect 3307 1316 3308 1320
rect 3302 1315 3308 1316
rect 3376 1312 3378 1346
rect 3464 1343 3466 1366
rect 3463 1342 3467 1343
rect 3463 1337 3467 1338
rect 3464 1318 3466 1337
rect 3462 1317 3468 1318
rect 3462 1313 3463 1317
rect 3467 1313 3468 1317
rect 3462 1312 3468 1313
rect 3062 1311 3068 1312
rect 3062 1307 3063 1311
rect 3067 1307 3068 1311
rect 3062 1306 3068 1307
rect 3214 1311 3220 1312
rect 3214 1307 3215 1311
rect 3219 1307 3220 1311
rect 3214 1306 3220 1307
rect 3374 1311 3380 1312
rect 3374 1307 3375 1311
rect 3379 1307 3380 1311
rect 3374 1306 3380 1307
rect 3142 1301 3148 1302
rect 3142 1297 3143 1301
rect 3147 1297 3148 1301
rect 3142 1296 3148 1297
rect 3302 1301 3308 1302
rect 3302 1297 3303 1301
rect 3307 1297 3308 1301
rect 3302 1296 3308 1297
rect 3462 1300 3468 1301
rect 3462 1296 3463 1300
rect 3467 1296 3468 1300
rect 3144 1279 3146 1296
rect 3304 1279 3306 1296
rect 3462 1295 3468 1296
rect 3464 1279 3466 1295
rect 3143 1278 3147 1279
rect 3143 1273 3147 1274
rect 3303 1278 3307 1279
rect 3303 1273 3307 1274
rect 3463 1278 3467 1279
rect 3463 1273 3467 1274
rect 3144 1256 3146 1273
rect 3464 1257 3466 1273
rect 3462 1256 3468 1257
rect 3142 1255 3148 1256
rect 3142 1251 3143 1255
rect 3147 1251 3148 1255
rect 3462 1252 3463 1256
rect 3467 1252 3468 1256
rect 3462 1251 3468 1252
rect 3142 1250 3148 1251
rect 3054 1247 3060 1248
rect 2886 1243 2892 1244
rect 2886 1239 2887 1243
rect 2891 1239 2892 1243
rect 2886 1238 2892 1239
rect 3046 1243 3052 1244
rect 3046 1239 3047 1243
rect 3051 1239 3052 1243
rect 3054 1243 3055 1247
rect 3059 1243 3060 1247
rect 3054 1242 3060 1243
rect 3046 1238 3052 1239
rect 3462 1239 3468 1240
rect 2814 1236 2820 1237
rect 2814 1232 2815 1236
rect 2819 1232 2820 1236
rect 2814 1231 2820 1232
rect 2750 1219 2756 1220
rect 2750 1215 2751 1219
rect 2755 1215 2756 1219
rect 2574 1214 2580 1215
rect 2655 1214 2659 1215
rect 2655 1209 2659 1210
rect 2695 1214 2699 1215
rect 2750 1214 2756 1215
rect 2766 1219 2772 1220
rect 2766 1215 2767 1219
rect 2771 1215 2772 1219
rect 2816 1215 2818 1231
rect 2888 1220 2890 1238
rect 2974 1236 2980 1237
rect 2974 1232 2975 1236
rect 2979 1232 2980 1236
rect 2974 1231 2980 1232
rect 2886 1219 2892 1220
rect 2886 1215 2887 1219
rect 2891 1215 2892 1219
rect 2976 1215 2978 1231
rect 3048 1220 3050 1238
rect 3142 1236 3148 1237
rect 3142 1232 3143 1236
rect 3147 1232 3148 1236
rect 3462 1235 3463 1239
rect 3467 1235 3468 1239
rect 3462 1234 3468 1235
rect 3142 1231 3148 1232
rect 3046 1219 3052 1220
rect 3046 1215 3047 1219
rect 3051 1215 3052 1219
rect 3144 1215 3146 1231
rect 3464 1215 3466 1234
rect 2766 1214 2772 1215
rect 2815 1214 2819 1215
rect 2695 1209 2699 1210
rect 2566 1207 2572 1208
rect 2566 1203 2567 1207
rect 2571 1203 2572 1207
rect 2566 1202 2572 1203
rect 2696 1193 2698 1209
rect 2390 1192 2396 1193
rect 2390 1188 2391 1192
rect 2395 1188 2396 1192
rect 2390 1187 2396 1188
rect 2542 1192 2548 1193
rect 2542 1188 2543 1192
rect 2547 1188 2548 1192
rect 2542 1187 2548 1188
rect 2694 1192 2700 1193
rect 2694 1188 2695 1192
rect 2699 1188 2700 1192
rect 2694 1187 2700 1188
rect 2768 1184 2770 1214
rect 2815 1209 2819 1210
rect 2847 1214 2851 1215
rect 2886 1214 2892 1215
rect 2975 1214 2979 1215
rect 2847 1209 2851 1210
rect 2975 1209 2979 1210
rect 2999 1214 3003 1215
rect 3046 1214 3052 1215
rect 3143 1214 3147 1215
rect 2999 1209 3003 1210
rect 3143 1209 3147 1210
rect 3159 1214 3163 1215
rect 3159 1209 3163 1210
rect 3463 1214 3467 1215
rect 3463 1209 3467 1210
rect 2774 1207 2780 1208
rect 2774 1203 2775 1207
rect 2779 1203 2780 1207
rect 2774 1202 2780 1203
rect 2776 1184 2778 1202
rect 2848 1193 2850 1209
rect 2942 1207 2948 1208
rect 2942 1203 2943 1207
rect 2947 1203 2948 1207
rect 2942 1202 2948 1203
rect 2846 1192 2852 1193
rect 2846 1188 2847 1192
rect 2851 1188 2852 1192
rect 2846 1187 2852 1188
rect 2006 1183 2012 1184
rect 2006 1179 2007 1183
rect 2011 1179 2012 1183
rect 2006 1178 2012 1179
rect 2150 1183 2156 1184
rect 2150 1179 2151 1183
rect 2155 1179 2156 1183
rect 2150 1178 2156 1179
rect 2302 1183 2308 1184
rect 2302 1179 2303 1183
rect 2307 1179 2308 1183
rect 2302 1178 2308 1179
rect 2310 1183 2316 1184
rect 2310 1179 2311 1183
rect 2315 1179 2316 1183
rect 2310 1178 2316 1179
rect 2606 1183 2612 1184
rect 2606 1179 2607 1183
rect 2611 1179 2612 1183
rect 2606 1178 2612 1179
rect 2766 1183 2772 1184
rect 2766 1179 2767 1183
rect 2771 1179 2772 1183
rect 2766 1178 2772 1179
rect 2774 1183 2780 1184
rect 2774 1179 2775 1183
rect 2779 1179 2780 1183
rect 2774 1178 2780 1179
rect 1934 1173 1940 1174
rect 1934 1169 1935 1173
rect 1939 1169 1940 1173
rect 1934 1168 1940 1169
rect 2078 1173 2084 1174
rect 2078 1169 2079 1173
rect 2083 1169 2084 1173
rect 2078 1168 2084 1169
rect 2230 1173 2236 1174
rect 2230 1169 2231 1173
rect 2235 1169 2236 1173
rect 2230 1168 2236 1169
rect 2390 1173 2396 1174
rect 2390 1169 2391 1173
rect 2395 1169 2396 1173
rect 2390 1168 2396 1169
rect 2542 1173 2548 1174
rect 2542 1169 2543 1173
rect 2547 1169 2548 1173
rect 2542 1168 2548 1169
rect 1936 1139 1938 1168
rect 2080 1139 2082 1168
rect 2232 1139 2234 1168
rect 2392 1139 2394 1168
rect 2544 1139 2546 1168
rect 1935 1138 1939 1139
rect 1935 1133 1939 1134
rect 1983 1138 1987 1139
rect 1983 1133 1987 1134
rect 2079 1138 2083 1139
rect 2079 1133 2083 1134
rect 2111 1138 2115 1139
rect 2111 1133 2115 1134
rect 2231 1138 2235 1139
rect 2231 1133 2235 1134
rect 2247 1138 2251 1139
rect 2247 1133 2251 1134
rect 2383 1138 2387 1139
rect 2383 1133 2387 1134
rect 2391 1138 2395 1139
rect 2391 1133 2395 1134
rect 2511 1138 2515 1139
rect 2511 1133 2515 1134
rect 2543 1138 2547 1139
rect 2543 1133 2547 1134
rect 1984 1116 1986 1133
rect 2112 1116 2114 1133
rect 2248 1116 2250 1133
rect 2384 1116 2386 1133
rect 2512 1116 2514 1133
rect 1982 1115 1988 1116
rect 1862 1110 1868 1111
rect 1926 1111 1932 1112
rect 1926 1107 1927 1111
rect 1931 1107 1932 1111
rect 1982 1111 1983 1115
rect 1987 1111 1988 1115
rect 1982 1110 1988 1111
rect 2110 1115 2116 1116
rect 2110 1111 2111 1115
rect 2115 1111 2116 1115
rect 2110 1110 2116 1111
rect 2246 1115 2252 1116
rect 2246 1111 2247 1115
rect 2251 1111 2252 1115
rect 2246 1110 2252 1111
rect 2382 1115 2388 1116
rect 2382 1111 2383 1115
rect 2387 1111 2388 1115
rect 2382 1110 2388 1111
rect 2510 1115 2516 1116
rect 2510 1111 2511 1115
rect 2515 1111 2516 1115
rect 2510 1110 2516 1111
rect 1926 1106 1932 1107
rect 1942 1107 1948 1108
rect 1942 1103 1943 1107
rect 1947 1103 1948 1107
rect 1942 1102 1948 1103
rect 2062 1107 2068 1108
rect 2062 1103 2063 1107
rect 2067 1103 2068 1107
rect 2062 1102 2068 1103
rect 2190 1107 2196 1108
rect 2190 1103 2191 1107
rect 2195 1103 2196 1107
rect 2190 1102 2196 1103
rect 2582 1103 2588 1104
rect 1766 1100 1772 1101
rect 1406 1099 1412 1100
rect 1406 1095 1407 1099
rect 1411 1095 1412 1099
rect 1406 1094 1412 1095
rect 1558 1099 1564 1100
rect 1558 1095 1559 1099
rect 1563 1095 1564 1099
rect 1766 1096 1767 1100
rect 1771 1096 1772 1100
rect 1766 1095 1772 1096
rect 1806 1099 1812 1100
rect 1806 1095 1807 1099
rect 1811 1095 1812 1099
rect 1558 1094 1564 1095
rect 1806 1094 1812 1095
rect 1862 1096 1868 1097
rect 1334 1087 1340 1088
rect 1334 1083 1335 1087
rect 1339 1083 1340 1087
rect 1334 1082 1340 1083
rect 1478 1087 1484 1088
rect 1478 1083 1479 1087
rect 1483 1083 1484 1087
rect 1478 1082 1484 1083
rect 1766 1083 1772 1084
rect 1278 1071 1284 1072
rect 1278 1067 1279 1071
rect 1283 1067 1284 1071
rect 1278 1066 1284 1067
rect 1336 1064 1338 1082
rect 1406 1080 1412 1081
rect 1406 1076 1407 1080
rect 1411 1076 1412 1080
rect 1406 1075 1412 1076
rect 1334 1063 1340 1064
rect 1334 1059 1335 1063
rect 1339 1059 1340 1063
rect 1334 1058 1340 1059
rect 1408 1051 1410 1075
rect 1480 1064 1482 1082
rect 1558 1080 1564 1081
rect 1558 1076 1559 1080
rect 1563 1076 1564 1080
rect 1766 1079 1767 1083
rect 1771 1079 1772 1083
rect 1766 1078 1772 1079
rect 1558 1075 1564 1076
rect 1478 1063 1484 1064
rect 1478 1059 1479 1063
rect 1483 1059 1484 1063
rect 1478 1058 1484 1059
rect 1560 1051 1562 1075
rect 1768 1051 1770 1078
rect 1808 1067 1810 1094
rect 1862 1092 1863 1096
rect 1867 1092 1868 1096
rect 1862 1091 1868 1092
rect 1864 1067 1866 1091
rect 1944 1080 1946 1102
rect 1982 1096 1988 1097
rect 1982 1092 1983 1096
rect 1987 1092 1988 1096
rect 1982 1091 1988 1092
rect 1942 1079 1948 1080
rect 1942 1075 1943 1079
rect 1947 1075 1948 1079
rect 1942 1074 1948 1075
rect 1984 1067 1986 1091
rect 2064 1080 2066 1102
rect 2110 1096 2116 1097
rect 2110 1092 2111 1096
rect 2115 1092 2116 1096
rect 2110 1091 2116 1092
rect 2062 1079 2068 1080
rect 2062 1075 2063 1079
rect 2067 1075 2068 1079
rect 2062 1074 2068 1075
rect 2112 1067 2114 1091
rect 2192 1080 2194 1102
rect 2582 1099 2583 1103
rect 2587 1099 2588 1103
rect 2582 1098 2588 1099
rect 2246 1096 2252 1097
rect 2246 1092 2247 1096
rect 2251 1092 2252 1096
rect 2246 1091 2252 1092
rect 2382 1096 2388 1097
rect 2382 1092 2383 1096
rect 2387 1092 2388 1096
rect 2382 1091 2388 1092
rect 2510 1096 2516 1097
rect 2510 1092 2511 1096
rect 2515 1092 2516 1096
rect 2510 1091 2516 1092
rect 2190 1079 2196 1080
rect 2190 1075 2191 1079
rect 2195 1075 2196 1079
rect 2190 1074 2196 1075
rect 2174 1067 2180 1068
rect 2248 1067 2250 1091
rect 2350 1079 2356 1080
rect 2350 1075 2351 1079
rect 2355 1075 2356 1079
rect 2350 1074 2356 1075
rect 1807 1066 1811 1067
rect 1807 1061 1811 1062
rect 1863 1066 1867 1067
rect 1863 1061 1867 1062
rect 1983 1066 1987 1067
rect 1983 1061 1987 1062
rect 2103 1066 2107 1067
rect 2103 1061 2107 1062
rect 2111 1066 2115 1067
rect 2174 1063 2175 1067
rect 2179 1063 2180 1067
rect 2174 1062 2180 1063
rect 2191 1066 2195 1067
rect 2111 1061 2115 1062
rect 767 1050 771 1051
rect 767 1045 771 1046
rect 815 1050 819 1051
rect 815 1045 819 1046
rect 927 1050 931 1051
rect 927 1045 931 1046
rect 967 1050 971 1051
rect 967 1045 971 1046
rect 1079 1050 1083 1051
rect 1079 1045 1083 1046
rect 1119 1050 1123 1051
rect 1119 1045 1123 1046
rect 1231 1050 1235 1051
rect 1231 1045 1235 1046
rect 1263 1050 1267 1051
rect 1263 1045 1267 1046
rect 1383 1050 1387 1051
rect 1383 1045 1387 1046
rect 1407 1050 1411 1051
rect 1407 1045 1411 1046
rect 1535 1050 1539 1051
rect 1535 1045 1539 1046
rect 1559 1050 1563 1051
rect 1559 1045 1563 1046
rect 1671 1050 1675 1051
rect 1671 1045 1675 1046
rect 1767 1050 1771 1051
rect 1767 1045 1771 1046
rect 768 1029 770 1045
rect 846 1043 852 1044
rect 846 1039 847 1043
rect 851 1039 852 1043
rect 846 1038 852 1039
rect 766 1028 772 1029
rect 766 1024 767 1028
rect 771 1024 772 1028
rect 766 1023 772 1024
rect 848 1020 850 1038
rect 928 1029 930 1045
rect 958 1043 964 1044
rect 958 1039 959 1043
rect 963 1039 964 1043
rect 958 1038 964 1039
rect 926 1028 932 1029
rect 926 1024 927 1028
rect 931 1024 932 1028
rect 926 1023 932 1024
rect 398 1019 404 1020
rect 398 1015 399 1019
rect 403 1015 404 1019
rect 398 1014 404 1015
rect 534 1019 540 1020
rect 534 1015 535 1019
rect 539 1015 540 1019
rect 534 1014 540 1015
rect 678 1019 684 1020
rect 678 1015 679 1019
rect 683 1015 684 1019
rect 678 1014 684 1015
rect 846 1019 852 1020
rect 846 1015 847 1019
rect 851 1015 852 1019
rect 846 1014 852 1015
rect 326 1009 332 1010
rect 110 1008 116 1009
rect 110 1004 111 1008
rect 115 1004 116 1008
rect 326 1005 327 1009
rect 331 1005 332 1009
rect 326 1004 332 1005
rect 462 1009 468 1010
rect 462 1005 463 1009
rect 467 1005 468 1009
rect 462 1004 468 1005
rect 606 1009 612 1010
rect 606 1005 607 1009
rect 611 1005 612 1009
rect 606 1004 612 1005
rect 766 1009 772 1010
rect 766 1005 767 1009
rect 771 1005 772 1009
rect 766 1004 772 1005
rect 926 1009 932 1010
rect 926 1005 927 1009
rect 931 1005 932 1009
rect 926 1004 932 1005
rect 110 1003 116 1004
rect 112 983 114 1003
rect 328 983 330 1004
rect 464 983 466 1004
rect 608 983 610 1004
rect 768 983 770 1004
rect 928 983 930 1004
rect 111 982 115 983
rect 111 977 115 978
rect 327 982 331 983
rect 327 977 331 978
rect 463 982 467 983
rect 463 977 467 978
rect 471 982 475 983
rect 471 977 475 978
rect 567 982 571 983
rect 567 977 571 978
rect 607 982 611 983
rect 607 977 611 978
rect 671 982 675 983
rect 671 977 675 978
rect 767 982 771 983
rect 767 977 771 978
rect 783 982 787 983
rect 783 977 787 978
rect 887 982 891 983
rect 887 977 891 978
rect 927 982 931 983
rect 927 977 931 978
rect 112 961 114 977
rect 110 960 116 961
rect 472 960 474 977
rect 568 960 570 977
rect 672 960 674 977
rect 784 960 786 977
rect 888 960 890 977
rect 110 956 111 960
rect 115 956 116 960
rect 110 955 116 956
rect 470 959 476 960
rect 470 955 471 959
rect 475 955 476 959
rect 470 954 476 955
rect 566 959 572 960
rect 566 955 567 959
rect 571 955 572 959
rect 566 954 572 955
rect 670 959 676 960
rect 670 955 671 959
rect 675 955 676 959
rect 670 954 676 955
rect 782 959 788 960
rect 782 955 783 959
rect 787 955 788 959
rect 782 954 788 955
rect 886 959 892 960
rect 886 955 887 959
rect 891 955 892 959
rect 886 954 892 955
rect 960 952 962 1038
rect 1080 1029 1082 1045
rect 1158 1043 1164 1044
rect 1158 1039 1159 1043
rect 1163 1039 1164 1043
rect 1158 1038 1164 1039
rect 1078 1028 1084 1029
rect 1078 1024 1079 1028
rect 1083 1024 1084 1028
rect 1078 1023 1084 1024
rect 1160 1020 1162 1038
rect 1232 1029 1234 1045
rect 1384 1029 1386 1045
rect 1462 1043 1468 1044
rect 1462 1039 1463 1043
rect 1467 1039 1468 1043
rect 1462 1038 1468 1039
rect 1470 1043 1476 1044
rect 1470 1039 1471 1043
rect 1475 1039 1476 1043
rect 1470 1038 1476 1039
rect 1230 1028 1236 1029
rect 1230 1024 1231 1028
rect 1235 1024 1236 1028
rect 1230 1023 1236 1024
rect 1382 1028 1388 1029
rect 1382 1024 1383 1028
rect 1387 1024 1388 1028
rect 1382 1023 1388 1024
rect 1046 1019 1052 1020
rect 1046 1015 1047 1019
rect 1051 1015 1052 1019
rect 1046 1014 1052 1015
rect 1158 1019 1164 1020
rect 1158 1015 1159 1019
rect 1163 1015 1164 1019
rect 1158 1014 1164 1015
rect 991 982 995 983
rect 991 977 995 978
rect 992 960 994 977
rect 990 959 996 960
rect 990 955 991 959
rect 995 955 996 959
rect 990 954 996 955
rect 958 951 964 952
rect 542 947 548 948
rect 110 943 116 944
rect 110 939 111 943
rect 115 939 116 943
rect 542 943 543 947
rect 547 943 548 947
rect 542 942 548 943
rect 638 947 644 948
rect 638 943 639 947
rect 643 943 644 947
rect 638 942 644 943
rect 742 947 748 948
rect 742 943 743 947
rect 747 943 748 947
rect 742 942 748 943
rect 854 947 860 948
rect 854 943 855 947
rect 859 943 860 947
rect 958 947 959 951
rect 963 947 964 951
rect 958 946 964 947
rect 854 942 860 943
rect 110 938 116 939
rect 470 940 476 941
rect 112 915 114 938
rect 470 936 471 940
rect 475 936 476 940
rect 470 935 476 936
rect 472 915 474 935
rect 544 924 546 942
rect 566 940 572 941
rect 566 936 567 940
rect 571 936 572 940
rect 566 935 572 936
rect 526 923 532 924
rect 526 919 527 923
rect 531 919 532 923
rect 526 918 532 919
rect 542 923 548 924
rect 542 919 543 923
rect 547 919 548 923
rect 542 918 548 919
rect 111 914 115 915
rect 111 909 115 910
rect 471 914 475 915
rect 471 909 475 910
rect 112 890 114 909
rect 110 889 116 890
rect 110 885 111 889
rect 115 885 116 889
rect 110 884 116 885
rect 528 884 530 918
rect 568 915 570 935
rect 640 924 642 942
rect 670 940 676 941
rect 670 936 671 940
rect 675 936 676 940
rect 670 935 676 936
rect 638 923 644 924
rect 638 919 639 923
rect 643 919 644 923
rect 638 918 644 919
rect 672 915 674 935
rect 744 924 746 942
rect 782 940 788 941
rect 782 936 783 940
rect 787 936 788 940
rect 782 935 788 936
rect 742 923 748 924
rect 742 919 743 923
rect 747 919 748 923
rect 742 918 748 919
rect 784 915 786 935
rect 856 924 858 942
rect 886 940 892 941
rect 886 936 887 940
rect 891 936 892 940
rect 886 935 892 936
rect 990 940 996 941
rect 990 936 991 940
rect 995 936 996 940
rect 990 935 996 936
rect 854 923 860 924
rect 854 919 855 923
rect 859 919 860 923
rect 854 918 860 919
rect 888 915 890 935
rect 992 915 994 935
rect 1048 924 1050 1014
rect 1078 1009 1084 1010
rect 1078 1005 1079 1009
rect 1083 1005 1084 1009
rect 1078 1004 1084 1005
rect 1230 1009 1236 1010
rect 1230 1005 1231 1009
rect 1235 1005 1236 1009
rect 1230 1004 1236 1005
rect 1382 1009 1388 1010
rect 1382 1005 1383 1009
rect 1387 1005 1388 1009
rect 1382 1004 1388 1005
rect 1080 983 1082 1004
rect 1232 983 1234 1004
rect 1384 983 1386 1004
rect 1079 982 1083 983
rect 1079 977 1083 978
rect 1095 982 1099 983
rect 1095 977 1099 978
rect 1199 982 1203 983
rect 1199 977 1203 978
rect 1231 982 1235 983
rect 1231 977 1235 978
rect 1295 982 1299 983
rect 1295 977 1299 978
rect 1383 982 1387 983
rect 1383 977 1387 978
rect 1391 982 1395 983
rect 1391 977 1395 978
rect 1096 960 1098 977
rect 1200 960 1202 977
rect 1296 960 1298 977
rect 1392 960 1394 977
rect 1094 959 1100 960
rect 1094 955 1095 959
rect 1099 955 1100 959
rect 1094 954 1100 955
rect 1198 959 1204 960
rect 1198 955 1199 959
rect 1203 955 1204 959
rect 1198 954 1204 955
rect 1294 959 1300 960
rect 1294 955 1295 959
rect 1299 955 1300 959
rect 1294 954 1300 955
rect 1390 959 1396 960
rect 1390 955 1391 959
rect 1395 955 1396 959
rect 1390 954 1396 955
rect 1464 952 1466 1038
rect 1472 1020 1474 1038
rect 1536 1029 1538 1045
rect 1606 1043 1612 1044
rect 1606 1039 1607 1043
rect 1611 1039 1612 1043
rect 1606 1038 1612 1039
rect 1534 1028 1540 1029
rect 1534 1024 1535 1028
rect 1539 1024 1540 1028
rect 1534 1023 1540 1024
rect 1608 1020 1610 1038
rect 1672 1029 1674 1045
rect 1670 1028 1676 1029
rect 1670 1024 1671 1028
rect 1675 1024 1676 1028
rect 1768 1026 1770 1045
rect 1808 1042 1810 1061
rect 2104 1045 2106 1061
rect 2102 1044 2108 1045
rect 1806 1041 1812 1042
rect 1806 1037 1807 1041
rect 1811 1037 1812 1041
rect 2102 1040 2103 1044
rect 2107 1040 2108 1044
rect 2102 1039 2108 1040
rect 1806 1036 1812 1037
rect 2176 1036 2178 1062
rect 2191 1061 2195 1062
rect 2247 1066 2251 1067
rect 2247 1061 2251 1062
rect 2279 1066 2283 1067
rect 2279 1061 2283 1062
rect 2192 1045 2194 1061
rect 2262 1059 2268 1060
rect 2262 1055 2263 1059
rect 2267 1055 2268 1059
rect 2262 1054 2268 1055
rect 2190 1044 2196 1045
rect 2190 1040 2191 1044
rect 2195 1040 2196 1044
rect 2190 1039 2196 1040
rect 2264 1036 2266 1054
rect 2280 1045 2282 1061
rect 2278 1044 2284 1045
rect 2278 1040 2279 1044
rect 2283 1040 2284 1044
rect 2278 1039 2284 1040
rect 2352 1036 2354 1074
rect 2384 1067 2386 1091
rect 2512 1067 2514 1091
rect 2367 1066 2371 1067
rect 2367 1061 2371 1062
rect 2383 1066 2387 1067
rect 2383 1061 2387 1062
rect 2455 1066 2459 1067
rect 2455 1061 2459 1062
rect 2511 1066 2515 1067
rect 2511 1061 2515 1062
rect 2543 1066 2547 1067
rect 2543 1061 2547 1062
rect 2368 1045 2370 1061
rect 2446 1059 2452 1060
rect 2446 1055 2447 1059
rect 2451 1055 2452 1059
rect 2446 1054 2452 1055
rect 2366 1044 2372 1045
rect 2366 1040 2367 1044
rect 2371 1040 2372 1044
rect 2366 1039 2372 1040
rect 2448 1036 2450 1054
rect 2456 1045 2458 1061
rect 2502 1059 2508 1060
rect 2502 1055 2503 1059
rect 2507 1055 2508 1059
rect 2502 1054 2508 1055
rect 2454 1044 2460 1045
rect 2454 1040 2455 1044
rect 2459 1040 2460 1044
rect 2454 1039 2460 1040
rect 2174 1035 2180 1036
rect 2174 1031 2175 1035
rect 2179 1031 2180 1035
rect 2174 1030 2180 1031
rect 2262 1035 2268 1036
rect 2262 1031 2263 1035
rect 2267 1031 2268 1035
rect 2262 1030 2268 1031
rect 2350 1035 2356 1036
rect 2350 1031 2351 1035
rect 2355 1031 2356 1035
rect 2350 1030 2356 1031
rect 2446 1035 2452 1036
rect 2446 1031 2447 1035
rect 2451 1031 2452 1035
rect 2446 1030 2452 1031
rect 1670 1023 1676 1024
rect 1766 1025 1772 1026
rect 2102 1025 2108 1026
rect 1766 1021 1767 1025
rect 1771 1021 1772 1025
rect 1766 1020 1772 1021
rect 1806 1024 1812 1025
rect 1806 1020 1807 1024
rect 1811 1020 1812 1024
rect 2102 1021 2103 1025
rect 2107 1021 2108 1025
rect 2102 1020 2108 1021
rect 2190 1025 2196 1026
rect 2190 1021 2191 1025
rect 2195 1021 2196 1025
rect 2190 1020 2196 1021
rect 2278 1025 2284 1026
rect 2278 1021 2279 1025
rect 2283 1021 2284 1025
rect 2278 1020 2284 1021
rect 2366 1025 2372 1026
rect 2366 1021 2367 1025
rect 2371 1021 2372 1025
rect 2366 1020 2372 1021
rect 2454 1025 2460 1026
rect 2454 1021 2455 1025
rect 2459 1021 2460 1025
rect 2454 1020 2460 1021
rect 1470 1019 1476 1020
rect 1470 1015 1471 1019
rect 1475 1015 1476 1019
rect 1470 1014 1476 1015
rect 1606 1019 1612 1020
rect 1606 1015 1607 1019
rect 1611 1015 1612 1019
rect 1606 1014 1612 1015
rect 1614 1019 1620 1020
rect 1806 1019 1812 1020
rect 1614 1015 1615 1019
rect 1619 1015 1620 1019
rect 1614 1014 1620 1015
rect 1534 1009 1540 1010
rect 1534 1005 1535 1009
rect 1539 1005 1540 1009
rect 1534 1004 1540 1005
rect 1536 983 1538 1004
rect 1487 982 1491 983
rect 1487 977 1491 978
rect 1535 982 1539 983
rect 1535 977 1539 978
rect 1583 982 1587 983
rect 1583 977 1587 978
rect 1488 960 1490 977
rect 1584 960 1586 977
rect 1486 959 1492 960
rect 1486 955 1487 959
rect 1491 955 1492 959
rect 1486 954 1492 955
rect 1582 959 1588 960
rect 1582 955 1583 959
rect 1587 955 1588 959
rect 1582 954 1588 955
rect 1462 951 1468 952
rect 1062 947 1068 948
rect 1062 943 1063 947
rect 1067 943 1068 947
rect 1062 942 1068 943
rect 1166 947 1172 948
rect 1166 943 1167 947
rect 1171 943 1172 947
rect 1166 942 1172 943
rect 1270 947 1276 948
rect 1270 943 1271 947
rect 1275 943 1276 947
rect 1270 942 1276 943
rect 1366 947 1372 948
rect 1366 943 1367 947
rect 1371 943 1372 947
rect 1462 947 1463 951
rect 1467 947 1468 951
rect 1462 946 1468 947
rect 1558 947 1564 948
rect 1366 942 1372 943
rect 1558 943 1559 947
rect 1563 943 1564 947
rect 1558 942 1564 943
rect 1046 923 1052 924
rect 1046 919 1047 923
rect 1051 919 1052 923
rect 1046 918 1052 919
rect 567 914 571 915
rect 567 909 571 910
rect 607 914 611 915
rect 607 909 611 910
rect 671 914 675 915
rect 671 909 675 910
rect 695 914 699 915
rect 695 909 699 910
rect 783 914 787 915
rect 783 909 787 910
rect 791 914 795 915
rect 791 909 795 910
rect 887 914 891 915
rect 887 909 891 910
rect 895 914 899 915
rect 895 909 899 910
rect 991 914 995 915
rect 991 909 995 910
rect 999 914 1003 915
rect 999 909 1003 910
rect 608 893 610 909
rect 696 893 698 909
rect 774 907 780 908
rect 774 903 775 907
rect 779 903 780 907
rect 774 902 780 903
rect 606 892 612 893
rect 606 888 607 892
rect 611 888 612 892
rect 606 887 612 888
rect 694 892 700 893
rect 694 888 695 892
rect 699 888 700 892
rect 694 887 700 888
rect 776 884 778 902
rect 792 893 794 909
rect 870 907 876 908
rect 870 903 871 907
rect 875 903 876 907
rect 870 902 876 903
rect 790 892 796 893
rect 790 888 791 892
rect 795 888 796 892
rect 790 887 796 888
rect 872 884 874 902
rect 896 893 898 909
rect 1000 893 1002 909
rect 1064 908 1066 942
rect 1094 940 1100 941
rect 1094 936 1095 940
rect 1099 936 1100 940
rect 1094 935 1100 936
rect 1096 915 1098 935
rect 1168 924 1170 942
rect 1198 940 1204 941
rect 1198 936 1199 940
rect 1203 936 1204 940
rect 1198 935 1204 936
rect 1166 923 1172 924
rect 1166 919 1167 923
rect 1171 919 1172 923
rect 1166 918 1172 919
rect 1200 915 1202 935
rect 1272 924 1274 942
rect 1294 940 1300 941
rect 1294 936 1295 940
rect 1299 936 1300 940
rect 1294 935 1300 936
rect 1270 923 1276 924
rect 1270 919 1271 923
rect 1275 919 1276 923
rect 1270 918 1276 919
rect 1296 915 1298 935
rect 1368 924 1370 942
rect 1390 940 1396 941
rect 1390 936 1391 940
rect 1395 936 1396 940
rect 1390 935 1396 936
rect 1486 940 1492 941
rect 1486 936 1487 940
rect 1491 936 1492 940
rect 1486 935 1492 936
rect 1366 923 1372 924
rect 1366 919 1367 923
rect 1371 919 1372 923
rect 1366 918 1372 919
rect 1302 915 1308 916
rect 1392 915 1394 935
rect 1488 915 1490 935
rect 1560 924 1562 942
rect 1582 940 1588 941
rect 1582 936 1583 940
rect 1587 936 1588 940
rect 1582 935 1588 936
rect 1558 923 1564 924
rect 1558 919 1559 923
rect 1563 919 1564 923
rect 1558 918 1564 919
rect 1584 915 1586 935
rect 1616 932 1618 1014
rect 1670 1009 1676 1010
rect 1670 1005 1671 1009
rect 1675 1005 1676 1009
rect 1670 1004 1676 1005
rect 1766 1008 1772 1009
rect 1766 1004 1767 1008
rect 1771 1004 1772 1008
rect 1672 983 1674 1004
rect 1766 1003 1772 1004
rect 1808 1003 1810 1019
rect 2104 1003 2106 1020
rect 2192 1003 2194 1020
rect 2280 1003 2282 1020
rect 2368 1003 2370 1020
rect 2456 1003 2458 1020
rect 1768 983 1770 1003
rect 1807 1002 1811 1003
rect 1807 997 1811 998
rect 2103 1002 2107 1003
rect 2103 997 2107 998
rect 2191 1002 2195 1003
rect 2191 997 2195 998
rect 2279 1002 2283 1003
rect 2279 997 2283 998
rect 2311 1002 2315 1003
rect 2311 997 2315 998
rect 2367 1002 2371 1003
rect 2367 997 2371 998
rect 2407 1002 2411 1003
rect 2407 997 2411 998
rect 2455 1002 2459 1003
rect 2455 997 2459 998
rect 1671 982 1675 983
rect 1671 977 1675 978
rect 1767 982 1771 983
rect 1808 981 1810 997
rect 1767 977 1771 978
rect 1806 980 1812 981
rect 2312 980 2314 997
rect 2408 980 2410 997
rect 1672 960 1674 977
rect 1768 961 1770 977
rect 1806 976 1807 980
rect 1811 976 1812 980
rect 1806 975 1812 976
rect 2310 979 2316 980
rect 2310 975 2311 979
rect 2315 975 2316 979
rect 2310 974 2316 975
rect 2406 979 2412 980
rect 2406 975 2407 979
rect 2411 975 2412 979
rect 2406 974 2412 975
rect 2504 972 2506 1054
rect 2544 1045 2546 1061
rect 2584 1060 2586 1098
rect 2608 1080 2610 1178
rect 2694 1173 2700 1174
rect 2694 1169 2695 1173
rect 2699 1169 2700 1173
rect 2694 1168 2700 1169
rect 2846 1173 2852 1174
rect 2846 1169 2847 1173
rect 2851 1169 2852 1173
rect 2846 1168 2852 1169
rect 2696 1139 2698 1168
rect 2848 1139 2850 1168
rect 2639 1138 2643 1139
rect 2639 1133 2643 1134
rect 2695 1138 2699 1139
rect 2695 1133 2699 1134
rect 2759 1138 2763 1139
rect 2759 1133 2763 1134
rect 2847 1138 2851 1139
rect 2847 1133 2851 1134
rect 2871 1138 2875 1139
rect 2871 1133 2875 1134
rect 2640 1116 2642 1133
rect 2760 1116 2762 1133
rect 2872 1116 2874 1133
rect 2638 1115 2644 1116
rect 2638 1111 2639 1115
rect 2643 1111 2644 1115
rect 2638 1110 2644 1111
rect 2758 1115 2764 1116
rect 2758 1111 2759 1115
rect 2763 1111 2764 1115
rect 2758 1110 2764 1111
rect 2870 1115 2876 1116
rect 2870 1111 2871 1115
rect 2875 1111 2876 1115
rect 2870 1110 2876 1111
rect 2944 1108 2946 1202
rect 3000 1193 3002 1209
rect 3070 1207 3076 1208
rect 3070 1203 3071 1207
rect 3075 1203 3076 1207
rect 3070 1202 3076 1203
rect 2998 1192 3004 1193
rect 2998 1188 2999 1192
rect 3003 1188 3004 1192
rect 2998 1187 3004 1188
rect 3072 1184 3074 1202
rect 3160 1193 3162 1209
rect 3158 1192 3164 1193
rect 3158 1188 3159 1192
rect 3163 1188 3164 1192
rect 3464 1190 3466 1209
rect 3158 1187 3164 1188
rect 3462 1189 3468 1190
rect 3462 1185 3463 1189
rect 3467 1185 3468 1189
rect 3462 1184 3468 1185
rect 3070 1183 3076 1184
rect 3070 1179 3071 1183
rect 3075 1179 3076 1183
rect 3070 1178 3076 1179
rect 2998 1173 3004 1174
rect 2998 1169 2999 1173
rect 3003 1169 3004 1173
rect 2998 1168 3004 1169
rect 3158 1173 3164 1174
rect 3158 1169 3159 1173
rect 3163 1169 3164 1173
rect 3158 1168 3164 1169
rect 3462 1172 3468 1173
rect 3462 1168 3463 1172
rect 3467 1168 3468 1172
rect 3000 1139 3002 1168
rect 3160 1139 3162 1168
rect 3462 1167 3468 1168
rect 3464 1139 3466 1167
rect 2975 1138 2979 1139
rect 2975 1133 2979 1134
rect 2999 1138 3003 1139
rect 2999 1133 3003 1134
rect 3079 1138 3083 1139
rect 3079 1133 3083 1134
rect 3159 1138 3163 1139
rect 3159 1133 3163 1134
rect 3183 1138 3187 1139
rect 3183 1133 3187 1134
rect 3279 1138 3283 1139
rect 3279 1133 3283 1134
rect 3367 1138 3371 1139
rect 3367 1133 3371 1134
rect 3463 1138 3467 1139
rect 3463 1133 3467 1134
rect 2976 1116 2978 1133
rect 3080 1116 3082 1133
rect 3184 1116 3186 1133
rect 3280 1116 3282 1133
rect 3368 1116 3370 1133
rect 3464 1117 3466 1133
rect 3462 1116 3468 1117
rect 2974 1115 2980 1116
rect 2974 1111 2975 1115
rect 2979 1111 2980 1115
rect 2974 1110 2980 1111
rect 3078 1115 3084 1116
rect 3078 1111 3079 1115
rect 3083 1111 3084 1115
rect 3078 1110 3084 1111
rect 3182 1115 3188 1116
rect 3182 1111 3183 1115
rect 3187 1111 3188 1115
rect 3182 1110 3188 1111
rect 3278 1115 3284 1116
rect 3278 1111 3279 1115
rect 3283 1111 3284 1115
rect 3278 1110 3284 1111
rect 3366 1115 3372 1116
rect 3366 1111 3367 1115
rect 3371 1111 3372 1115
rect 3462 1112 3463 1116
rect 3467 1112 3468 1116
rect 3462 1111 3468 1112
rect 3366 1110 3372 1111
rect 2942 1107 2948 1108
rect 2710 1103 2716 1104
rect 2710 1099 2711 1103
rect 2715 1099 2716 1103
rect 2710 1098 2716 1099
rect 2830 1103 2836 1104
rect 2830 1099 2831 1103
rect 2835 1099 2836 1103
rect 2942 1103 2943 1107
rect 2947 1103 2948 1107
rect 2942 1102 2948 1103
rect 2950 1107 2956 1108
rect 2950 1103 2951 1107
rect 2955 1103 2956 1107
rect 2950 1102 2956 1103
rect 3054 1107 3060 1108
rect 3054 1103 3055 1107
rect 3059 1103 3060 1107
rect 3054 1102 3060 1103
rect 3158 1107 3164 1108
rect 3158 1103 3159 1107
rect 3163 1103 3164 1107
rect 3158 1102 3164 1103
rect 3262 1107 3268 1108
rect 3262 1103 3263 1107
rect 3267 1103 3268 1107
rect 3262 1102 3268 1103
rect 2830 1098 2836 1099
rect 2638 1096 2644 1097
rect 2638 1092 2639 1096
rect 2643 1092 2644 1096
rect 2638 1091 2644 1092
rect 2606 1079 2612 1080
rect 2606 1075 2607 1079
rect 2611 1075 2612 1079
rect 2606 1074 2612 1075
rect 2640 1067 2642 1091
rect 2712 1080 2714 1098
rect 2758 1096 2764 1097
rect 2758 1092 2759 1096
rect 2763 1092 2764 1096
rect 2758 1091 2764 1092
rect 2710 1079 2716 1080
rect 2710 1075 2711 1079
rect 2715 1075 2716 1079
rect 2710 1074 2716 1075
rect 2760 1067 2762 1091
rect 2832 1080 2834 1098
rect 2870 1096 2876 1097
rect 2870 1092 2871 1096
rect 2875 1092 2876 1096
rect 2870 1091 2876 1092
rect 2830 1079 2836 1080
rect 2830 1075 2831 1079
rect 2835 1075 2836 1079
rect 2830 1074 2836 1075
rect 2872 1067 2874 1091
rect 2952 1088 2954 1102
rect 2974 1096 2980 1097
rect 2974 1092 2975 1096
rect 2979 1092 2980 1096
rect 2974 1091 2980 1092
rect 2950 1087 2956 1088
rect 2950 1083 2951 1087
rect 2955 1083 2956 1087
rect 2950 1082 2956 1083
rect 2976 1067 2978 1091
rect 3056 1080 3058 1102
rect 3078 1096 3084 1097
rect 3078 1092 3079 1096
rect 3083 1092 3084 1096
rect 3078 1091 3084 1092
rect 3054 1079 3060 1080
rect 3054 1075 3055 1079
rect 3059 1075 3060 1079
rect 3054 1074 3060 1075
rect 3080 1067 3082 1091
rect 3160 1080 3162 1102
rect 3182 1096 3188 1097
rect 3182 1092 3183 1096
rect 3187 1092 3188 1096
rect 3182 1091 3188 1092
rect 3158 1079 3164 1080
rect 3158 1075 3159 1079
rect 3163 1075 3164 1079
rect 3158 1074 3164 1075
rect 3184 1067 3186 1091
rect 3264 1080 3266 1102
rect 3462 1099 3468 1100
rect 3278 1096 3284 1097
rect 3278 1092 3279 1096
rect 3283 1092 3284 1096
rect 3278 1091 3284 1092
rect 3366 1096 3372 1097
rect 3366 1092 3367 1096
rect 3371 1092 3372 1096
rect 3462 1095 3463 1099
rect 3467 1095 3468 1099
rect 3462 1094 3468 1095
rect 3366 1091 3372 1092
rect 3262 1079 3268 1080
rect 3262 1075 3263 1079
rect 3267 1075 3268 1079
rect 3262 1074 3268 1075
rect 3280 1067 3282 1091
rect 3368 1067 3370 1091
rect 3438 1079 3444 1080
rect 3438 1075 3439 1079
rect 3443 1075 3444 1079
rect 3438 1074 3444 1075
rect 2631 1066 2635 1067
rect 2631 1061 2635 1062
rect 2639 1066 2643 1067
rect 2639 1061 2643 1062
rect 2719 1066 2723 1067
rect 2719 1061 2723 1062
rect 2759 1066 2763 1067
rect 2759 1061 2763 1062
rect 2807 1066 2811 1067
rect 2807 1061 2811 1062
rect 2871 1066 2875 1067
rect 2871 1061 2875 1062
rect 2975 1066 2979 1067
rect 2975 1061 2979 1062
rect 3079 1066 3083 1067
rect 3079 1061 3083 1062
rect 3183 1066 3187 1067
rect 3183 1061 3187 1062
rect 3279 1066 3283 1067
rect 3279 1061 3283 1062
rect 3367 1066 3371 1067
rect 3367 1061 3371 1062
rect 2582 1059 2588 1060
rect 2582 1055 2583 1059
rect 2587 1055 2588 1059
rect 2582 1054 2588 1055
rect 2614 1059 2620 1060
rect 2614 1055 2615 1059
rect 2619 1055 2620 1059
rect 2614 1054 2620 1055
rect 2542 1044 2548 1045
rect 2542 1040 2543 1044
rect 2547 1040 2548 1044
rect 2542 1039 2548 1040
rect 2616 1036 2618 1054
rect 2632 1045 2634 1061
rect 2702 1059 2708 1060
rect 2702 1055 2703 1059
rect 2707 1055 2708 1059
rect 2702 1054 2708 1055
rect 2630 1044 2636 1045
rect 2630 1040 2631 1044
rect 2635 1040 2636 1044
rect 2630 1039 2636 1040
rect 2704 1036 2706 1054
rect 2720 1045 2722 1061
rect 2790 1059 2796 1060
rect 2790 1055 2791 1059
rect 2795 1055 2796 1059
rect 2790 1054 2796 1055
rect 2718 1044 2724 1045
rect 2718 1040 2719 1044
rect 2723 1040 2724 1044
rect 2718 1039 2724 1040
rect 2792 1036 2794 1054
rect 2808 1045 2810 1061
rect 2806 1044 2812 1045
rect 2806 1040 2807 1044
rect 2811 1040 2812 1044
rect 2806 1039 2812 1040
rect 2614 1035 2620 1036
rect 2614 1031 2615 1035
rect 2619 1031 2620 1035
rect 2614 1030 2620 1031
rect 2702 1035 2708 1036
rect 2702 1031 2703 1035
rect 2707 1031 2708 1035
rect 2702 1030 2708 1031
rect 2790 1035 2796 1036
rect 2790 1031 2791 1035
rect 2795 1031 2796 1035
rect 2790 1030 2796 1031
rect 2878 1035 2884 1036
rect 2878 1031 2879 1035
rect 2883 1031 2884 1035
rect 2878 1030 2884 1031
rect 2542 1025 2548 1026
rect 2542 1021 2543 1025
rect 2547 1021 2548 1025
rect 2542 1020 2548 1021
rect 2630 1025 2636 1026
rect 2630 1021 2631 1025
rect 2635 1021 2636 1025
rect 2630 1020 2636 1021
rect 2718 1025 2724 1026
rect 2718 1021 2719 1025
rect 2723 1021 2724 1025
rect 2718 1020 2724 1021
rect 2806 1025 2812 1026
rect 2806 1021 2807 1025
rect 2811 1021 2812 1025
rect 2806 1020 2812 1021
rect 2544 1003 2546 1020
rect 2632 1003 2634 1020
rect 2720 1003 2722 1020
rect 2808 1003 2810 1020
rect 2511 1002 2515 1003
rect 2511 997 2515 998
rect 2543 1002 2547 1003
rect 2543 997 2547 998
rect 2623 1002 2627 1003
rect 2623 997 2627 998
rect 2631 1002 2635 1003
rect 2631 997 2635 998
rect 2719 1002 2723 1003
rect 2719 997 2723 998
rect 2751 1002 2755 1003
rect 2751 997 2755 998
rect 2807 1002 2811 1003
rect 2807 997 2811 998
rect 2512 980 2514 997
rect 2624 980 2626 997
rect 2752 980 2754 997
rect 2510 979 2516 980
rect 2510 975 2511 979
rect 2515 975 2516 979
rect 2510 974 2516 975
rect 2622 979 2628 980
rect 2622 975 2623 979
rect 2627 975 2628 979
rect 2622 974 2628 975
rect 2750 979 2756 980
rect 2750 975 2751 979
rect 2755 975 2756 979
rect 2750 974 2756 975
rect 2502 971 2508 972
rect 2382 967 2388 968
rect 1806 963 1812 964
rect 1766 960 1772 961
rect 1670 959 1676 960
rect 1670 955 1671 959
rect 1675 955 1676 959
rect 1766 956 1767 960
rect 1771 956 1772 960
rect 1806 959 1807 963
rect 1811 959 1812 963
rect 2382 963 2383 967
rect 2387 963 2388 967
rect 2382 962 2388 963
rect 2478 967 2484 968
rect 2478 963 2479 967
rect 2483 963 2484 967
rect 2502 967 2503 971
rect 2507 967 2508 971
rect 2502 966 2508 967
rect 2694 967 2700 968
rect 2478 962 2484 963
rect 2694 963 2695 967
rect 2699 963 2700 967
rect 2694 962 2700 963
rect 2822 967 2828 968
rect 2822 963 2823 967
rect 2827 963 2828 967
rect 2822 962 2828 963
rect 1806 958 1812 959
rect 2310 960 2316 961
rect 1766 955 1772 956
rect 1670 954 1676 955
rect 1654 947 1660 948
rect 1654 943 1655 947
rect 1659 943 1660 947
rect 1654 942 1660 943
rect 1742 947 1748 948
rect 1742 943 1743 947
rect 1747 943 1748 947
rect 1742 942 1748 943
rect 1766 943 1772 944
rect 1614 931 1620 932
rect 1614 927 1615 931
rect 1619 927 1620 931
rect 1614 926 1620 927
rect 1656 924 1658 942
rect 1670 940 1676 941
rect 1670 936 1671 940
rect 1675 936 1676 940
rect 1670 935 1676 936
rect 1654 923 1660 924
rect 1654 919 1655 923
rect 1659 919 1660 923
rect 1654 918 1660 919
rect 1672 915 1674 935
rect 1744 920 1746 942
rect 1766 939 1767 943
rect 1771 939 1772 943
rect 1766 938 1772 939
rect 1742 919 1748 920
rect 1742 915 1743 919
rect 1747 915 1748 919
rect 1768 915 1770 938
rect 1808 927 1810 958
rect 2310 956 2311 960
rect 2315 956 2316 960
rect 2310 955 2316 956
rect 2222 943 2228 944
rect 2222 939 2223 943
rect 2227 939 2228 943
rect 2222 938 2228 939
rect 1807 926 1811 927
rect 1807 921 1811 922
rect 1831 926 1835 927
rect 1831 921 1835 922
rect 1983 926 1987 927
rect 1983 921 1987 922
rect 2151 926 2155 927
rect 2151 921 2155 922
rect 1095 914 1099 915
rect 1095 909 1099 910
rect 1111 914 1115 915
rect 1111 909 1115 910
rect 1199 914 1203 915
rect 1199 909 1203 910
rect 1223 914 1227 915
rect 1223 909 1227 910
rect 1295 914 1299 915
rect 1302 911 1303 915
rect 1307 911 1308 915
rect 1302 910 1308 911
rect 1343 914 1347 915
rect 1295 909 1299 910
rect 1022 907 1028 908
rect 1022 903 1023 907
rect 1027 903 1028 907
rect 1022 902 1028 903
rect 1062 907 1068 908
rect 1062 903 1063 907
rect 1067 903 1068 907
rect 1062 902 1068 903
rect 894 892 900 893
rect 894 888 895 892
rect 899 888 900 892
rect 894 887 900 888
rect 998 892 1004 893
rect 998 888 999 892
rect 1003 888 1004 892
rect 998 887 1004 888
rect 526 883 532 884
rect 526 879 527 883
rect 531 879 532 883
rect 526 878 532 879
rect 774 883 780 884
rect 774 879 775 883
rect 779 879 780 883
rect 774 878 780 879
rect 870 883 876 884
rect 870 879 871 883
rect 875 879 876 883
rect 870 878 876 879
rect 606 873 612 874
rect 110 872 116 873
rect 110 868 111 872
rect 115 868 116 872
rect 606 869 607 873
rect 611 869 612 873
rect 606 868 612 869
rect 694 873 700 874
rect 694 869 695 873
rect 699 869 700 873
rect 694 868 700 869
rect 790 873 796 874
rect 790 869 791 873
rect 795 869 796 873
rect 790 868 796 869
rect 894 873 900 874
rect 894 869 895 873
rect 899 869 900 873
rect 894 868 900 869
rect 998 873 1004 874
rect 998 869 999 873
rect 1003 869 1004 873
rect 998 868 1004 869
rect 110 867 116 868
rect 112 847 114 867
rect 608 847 610 868
rect 696 847 698 868
rect 792 847 794 868
rect 896 847 898 868
rect 1000 847 1002 868
rect 111 846 115 847
rect 111 841 115 842
rect 519 846 523 847
rect 519 841 523 842
rect 607 846 611 847
rect 607 841 611 842
rect 615 846 619 847
rect 615 841 619 842
rect 695 846 699 847
rect 695 841 699 842
rect 719 846 723 847
rect 719 841 723 842
rect 791 846 795 847
rect 791 841 795 842
rect 831 846 835 847
rect 831 841 835 842
rect 895 846 899 847
rect 895 841 899 842
rect 951 846 955 847
rect 951 841 955 842
rect 999 846 1003 847
rect 999 841 1003 842
rect 112 825 114 841
rect 110 824 116 825
rect 520 824 522 841
rect 616 824 618 841
rect 720 824 722 841
rect 832 824 834 841
rect 952 824 954 841
rect 110 820 111 824
rect 115 820 116 824
rect 110 819 116 820
rect 518 823 524 824
rect 518 819 519 823
rect 523 819 524 823
rect 518 818 524 819
rect 614 823 620 824
rect 614 819 615 823
rect 619 819 620 823
rect 614 818 620 819
rect 718 823 724 824
rect 718 819 719 823
rect 723 819 724 823
rect 718 818 724 819
rect 830 823 836 824
rect 830 819 831 823
rect 835 819 836 823
rect 830 818 836 819
rect 950 823 956 824
rect 950 819 951 823
rect 955 819 956 823
rect 950 818 956 819
rect 1024 816 1026 902
rect 1112 893 1114 909
rect 1182 907 1188 908
rect 1182 903 1183 907
rect 1187 903 1188 907
rect 1182 902 1188 903
rect 1110 892 1116 893
rect 1110 888 1111 892
rect 1115 888 1116 892
rect 1110 887 1116 888
rect 1184 884 1186 902
rect 1224 893 1226 909
rect 1222 892 1228 893
rect 1222 888 1223 892
rect 1227 888 1228 892
rect 1222 887 1228 888
rect 1304 884 1306 910
rect 1343 909 1347 910
rect 1391 914 1395 915
rect 1391 909 1395 910
rect 1463 914 1467 915
rect 1463 909 1467 910
rect 1487 914 1491 915
rect 1487 909 1491 910
rect 1583 914 1587 915
rect 1583 909 1587 910
rect 1671 914 1675 915
rect 1742 914 1748 915
rect 1767 914 1771 915
rect 1671 909 1675 910
rect 1767 909 1771 910
rect 1344 893 1346 909
rect 1464 893 1466 909
rect 1566 907 1572 908
rect 1566 903 1567 907
rect 1571 903 1572 907
rect 1566 902 1572 903
rect 1342 892 1348 893
rect 1342 888 1343 892
rect 1347 888 1348 892
rect 1342 887 1348 888
rect 1462 892 1468 893
rect 1462 888 1463 892
rect 1467 888 1468 892
rect 1462 887 1468 888
rect 1568 884 1570 902
rect 1584 893 1586 909
rect 1630 907 1636 908
rect 1630 903 1631 907
rect 1635 903 1636 907
rect 1630 902 1636 903
rect 1582 892 1588 893
rect 1582 888 1583 892
rect 1587 888 1588 892
rect 1582 887 1588 888
rect 1182 883 1188 884
rect 1182 879 1183 883
rect 1187 879 1188 883
rect 1182 878 1188 879
rect 1198 883 1204 884
rect 1198 879 1199 883
rect 1203 879 1204 883
rect 1198 878 1204 879
rect 1302 883 1308 884
rect 1302 879 1303 883
rect 1307 879 1308 883
rect 1302 878 1308 879
rect 1566 883 1572 884
rect 1566 879 1567 883
rect 1571 879 1572 883
rect 1566 878 1572 879
rect 1110 873 1116 874
rect 1110 869 1111 873
rect 1115 869 1116 873
rect 1110 868 1116 869
rect 1112 847 1114 868
rect 1071 846 1075 847
rect 1071 841 1075 842
rect 1111 846 1115 847
rect 1111 841 1115 842
rect 1191 846 1195 847
rect 1191 841 1195 842
rect 1072 824 1074 841
rect 1192 824 1194 841
rect 1070 823 1076 824
rect 1070 819 1071 823
rect 1075 819 1076 823
rect 1070 818 1076 819
rect 1190 823 1196 824
rect 1190 819 1191 823
rect 1195 819 1196 823
rect 1190 818 1196 819
rect 1022 815 1028 816
rect 686 811 692 812
rect 110 807 116 808
rect 110 803 111 807
rect 115 803 116 807
rect 686 807 687 811
rect 691 807 692 811
rect 686 806 692 807
rect 790 811 796 812
rect 790 807 791 811
rect 795 807 796 811
rect 790 806 796 807
rect 902 811 908 812
rect 902 807 903 811
rect 907 807 908 811
rect 1022 811 1023 815
rect 1027 811 1028 815
rect 1022 810 1028 811
rect 1142 811 1148 812
rect 902 806 908 807
rect 1142 807 1143 811
rect 1147 807 1148 811
rect 1142 806 1148 807
rect 110 802 116 803
rect 518 804 524 805
rect 112 779 114 802
rect 518 800 519 804
rect 523 800 524 804
rect 518 799 524 800
rect 614 804 620 805
rect 614 800 615 804
rect 619 800 620 804
rect 614 799 620 800
rect 520 779 522 799
rect 616 779 618 799
rect 688 788 690 806
rect 718 804 724 805
rect 718 800 719 804
rect 723 800 724 804
rect 718 799 724 800
rect 686 787 692 788
rect 686 783 687 787
rect 691 783 692 787
rect 686 782 692 783
rect 720 779 722 799
rect 792 788 794 806
rect 830 804 836 805
rect 830 800 831 804
rect 835 800 836 804
rect 830 799 836 800
rect 790 787 796 788
rect 790 783 791 787
rect 795 783 796 787
rect 790 782 796 783
rect 758 779 764 780
rect 832 779 834 799
rect 904 788 906 806
rect 950 804 956 805
rect 950 800 951 804
rect 955 800 956 804
rect 950 799 956 800
rect 1070 804 1076 805
rect 1070 800 1071 804
rect 1075 800 1076 804
rect 1070 799 1076 800
rect 902 787 908 788
rect 902 783 903 787
rect 907 783 908 787
rect 902 782 908 783
rect 952 779 954 799
rect 1072 779 1074 799
rect 111 778 115 779
rect 111 773 115 774
rect 383 778 387 779
rect 383 773 387 774
rect 471 778 475 779
rect 471 773 475 774
rect 519 778 523 779
rect 519 773 523 774
rect 575 778 579 779
rect 575 773 579 774
rect 615 778 619 779
rect 615 773 619 774
rect 679 778 683 779
rect 679 773 683 774
rect 719 778 723 779
rect 758 775 759 779
rect 763 775 764 779
rect 758 774 764 775
rect 791 778 795 779
rect 719 773 723 774
rect 112 754 114 773
rect 384 757 386 773
rect 454 771 460 772
rect 454 767 455 771
rect 459 767 460 771
rect 454 766 460 767
rect 382 756 388 757
rect 110 753 116 754
rect 110 749 111 753
rect 115 749 116 753
rect 382 752 383 756
rect 387 752 388 756
rect 382 751 388 752
rect 110 748 116 749
rect 456 748 458 766
rect 472 757 474 773
rect 542 771 548 772
rect 542 767 543 771
rect 547 767 548 771
rect 542 766 548 767
rect 470 756 476 757
rect 470 752 471 756
rect 475 752 476 756
rect 470 751 476 752
rect 544 748 546 766
rect 576 757 578 773
rect 646 771 652 772
rect 646 767 647 771
rect 651 767 652 771
rect 646 766 652 767
rect 574 756 580 757
rect 574 752 575 756
rect 579 752 580 756
rect 574 751 580 752
rect 648 748 650 766
rect 654 763 660 764
rect 654 759 655 763
rect 659 759 660 763
rect 654 758 660 759
rect 454 747 460 748
rect 454 743 455 747
rect 459 743 460 747
rect 454 742 460 743
rect 542 747 548 748
rect 542 743 543 747
rect 547 743 548 747
rect 542 742 548 743
rect 646 747 652 748
rect 646 743 647 747
rect 651 743 652 747
rect 646 742 652 743
rect 382 737 388 738
rect 110 736 116 737
rect 110 732 111 736
rect 115 732 116 736
rect 382 733 383 737
rect 387 733 388 737
rect 382 732 388 733
rect 470 737 476 738
rect 470 733 471 737
rect 475 733 476 737
rect 470 732 476 733
rect 574 737 580 738
rect 574 733 575 737
rect 579 733 580 737
rect 574 732 580 733
rect 110 731 116 732
rect 112 707 114 731
rect 384 707 386 732
rect 472 707 474 732
rect 576 707 578 732
rect 111 706 115 707
rect 111 701 115 702
rect 247 706 251 707
rect 247 701 251 702
rect 343 706 347 707
rect 343 701 347 702
rect 383 706 387 707
rect 383 701 387 702
rect 455 706 459 707
rect 455 701 459 702
rect 471 706 475 707
rect 471 701 475 702
rect 567 706 571 707
rect 567 701 571 702
rect 575 706 579 707
rect 575 701 579 702
rect 112 685 114 701
rect 110 684 116 685
rect 248 684 250 701
rect 344 684 346 701
rect 456 684 458 701
rect 568 684 570 701
rect 110 680 111 684
rect 115 680 116 684
rect 110 679 116 680
rect 246 683 252 684
rect 246 679 247 683
rect 251 679 252 683
rect 246 678 252 679
rect 342 683 348 684
rect 342 679 343 683
rect 347 679 348 683
rect 342 678 348 679
rect 454 683 460 684
rect 454 679 455 683
rect 459 679 460 683
rect 454 678 460 679
rect 566 683 572 684
rect 566 679 567 683
rect 571 679 572 683
rect 566 678 572 679
rect 656 676 658 758
rect 680 757 682 773
rect 750 771 756 772
rect 750 767 751 771
rect 755 767 756 771
rect 750 766 756 767
rect 678 756 684 757
rect 678 752 679 756
rect 683 752 684 756
rect 678 751 684 752
rect 752 748 754 766
rect 760 748 762 774
rect 791 773 795 774
rect 831 778 835 779
rect 831 773 835 774
rect 911 778 915 779
rect 911 773 915 774
rect 951 778 955 779
rect 951 773 955 774
rect 1031 778 1035 779
rect 1031 773 1035 774
rect 1071 778 1075 779
rect 1071 773 1075 774
rect 792 757 794 773
rect 912 757 914 773
rect 990 771 996 772
rect 990 767 991 771
rect 995 767 996 771
rect 990 766 996 767
rect 790 756 796 757
rect 790 752 791 756
rect 795 752 796 756
rect 790 751 796 752
rect 910 756 916 757
rect 910 752 911 756
rect 915 752 916 756
rect 910 751 916 752
rect 992 748 994 766
rect 1032 757 1034 773
rect 1144 772 1146 806
rect 1190 804 1196 805
rect 1190 800 1191 804
rect 1195 800 1196 804
rect 1190 799 1196 800
rect 1192 779 1194 799
rect 1200 788 1202 878
rect 1222 873 1228 874
rect 1222 869 1223 873
rect 1227 869 1228 873
rect 1222 868 1228 869
rect 1342 873 1348 874
rect 1342 869 1343 873
rect 1347 869 1348 873
rect 1342 868 1348 869
rect 1462 873 1468 874
rect 1462 869 1463 873
rect 1467 869 1468 873
rect 1462 868 1468 869
rect 1582 873 1588 874
rect 1582 869 1583 873
rect 1587 869 1588 873
rect 1582 868 1588 869
rect 1224 847 1226 868
rect 1344 847 1346 868
rect 1464 847 1466 868
rect 1584 847 1586 868
rect 1223 846 1227 847
rect 1223 841 1227 842
rect 1311 846 1315 847
rect 1311 841 1315 842
rect 1343 846 1347 847
rect 1343 841 1347 842
rect 1431 846 1435 847
rect 1431 841 1435 842
rect 1463 846 1467 847
rect 1463 841 1467 842
rect 1559 846 1563 847
rect 1559 841 1563 842
rect 1583 846 1587 847
rect 1583 841 1587 842
rect 1312 824 1314 841
rect 1432 824 1434 841
rect 1560 824 1562 841
rect 1310 823 1316 824
rect 1310 819 1311 823
rect 1315 819 1316 823
rect 1310 818 1316 819
rect 1430 823 1436 824
rect 1430 819 1431 823
rect 1435 819 1436 823
rect 1430 818 1436 819
rect 1558 823 1564 824
rect 1558 819 1559 823
rect 1563 819 1564 823
rect 1558 818 1564 819
rect 1632 816 1634 902
rect 1768 890 1770 909
rect 1808 902 1810 921
rect 1832 905 1834 921
rect 1984 905 1986 921
rect 2038 919 2044 920
rect 2038 915 2039 919
rect 2043 915 2044 919
rect 2038 914 2044 915
rect 2054 919 2060 920
rect 2054 915 2055 919
rect 2059 915 2060 919
rect 2054 914 2060 915
rect 1830 904 1836 905
rect 1806 901 1812 902
rect 1806 897 1807 901
rect 1811 897 1812 901
rect 1830 900 1831 904
rect 1835 900 1836 904
rect 1830 899 1836 900
rect 1982 904 1988 905
rect 1982 900 1983 904
rect 1987 900 1988 904
rect 1982 899 1988 900
rect 1806 896 1812 897
rect 1894 895 1900 896
rect 1894 891 1895 895
rect 1899 891 1900 895
rect 1894 890 1900 891
rect 1766 889 1772 890
rect 1766 885 1767 889
rect 1771 885 1772 889
rect 1830 885 1836 886
rect 1766 884 1772 885
rect 1806 884 1812 885
rect 1806 880 1807 884
rect 1811 880 1812 884
rect 1830 881 1831 885
rect 1835 881 1836 885
rect 1830 880 1836 881
rect 1806 879 1812 880
rect 1766 872 1772 873
rect 1766 868 1767 872
rect 1771 868 1772 872
rect 1766 867 1772 868
rect 1768 847 1770 867
rect 1808 859 1810 879
rect 1832 859 1834 880
rect 1807 858 1811 859
rect 1807 853 1811 854
rect 1831 858 1835 859
rect 1831 853 1835 854
rect 1767 846 1771 847
rect 1767 841 1771 842
rect 1768 825 1770 841
rect 1808 837 1810 853
rect 1806 836 1812 837
rect 1832 836 1834 853
rect 1806 832 1807 836
rect 1811 832 1812 836
rect 1806 831 1812 832
rect 1830 835 1836 836
rect 1830 831 1831 835
rect 1835 831 1836 835
rect 1830 830 1836 831
rect 1766 824 1772 825
rect 1766 820 1767 824
rect 1771 820 1772 824
rect 1766 819 1772 820
rect 1806 819 1812 820
rect 1630 815 1636 816
rect 1262 811 1268 812
rect 1262 807 1263 811
rect 1267 807 1268 811
rect 1262 806 1268 807
rect 1382 811 1388 812
rect 1382 807 1383 811
rect 1387 807 1388 811
rect 1382 806 1388 807
rect 1502 811 1508 812
rect 1502 807 1503 811
rect 1507 807 1508 811
rect 1630 811 1631 815
rect 1635 811 1636 815
rect 1806 815 1807 819
rect 1811 815 1812 819
rect 1806 814 1812 815
rect 1830 816 1836 817
rect 1630 810 1636 811
rect 1502 806 1508 807
rect 1766 807 1772 808
rect 1264 788 1266 806
rect 1310 804 1316 805
rect 1310 800 1311 804
rect 1315 800 1316 804
rect 1310 799 1316 800
rect 1198 787 1204 788
rect 1198 783 1199 787
rect 1203 783 1204 787
rect 1198 782 1204 783
rect 1230 787 1236 788
rect 1230 783 1231 787
rect 1235 783 1236 787
rect 1230 782 1236 783
rect 1262 787 1268 788
rect 1262 783 1263 787
rect 1267 783 1268 787
rect 1262 782 1268 783
rect 1159 778 1163 779
rect 1159 773 1163 774
rect 1191 778 1195 779
rect 1191 773 1195 774
rect 1142 771 1148 772
rect 1142 767 1143 771
rect 1147 767 1148 771
rect 1142 766 1148 767
rect 1160 757 1162 773
rect 1030 756 1036 757
rect 1030 752 1031 756
rect 1035 752 1036 756
rect 1030 751 1036 752
rect 1158 756 1164 757
rect 1158 752 1159 756
rect 1163 752 1164 756
rect 1158 751 1164 752
rect 1232 748 1234 782
rect 1312 779 1314 799
rect 1384 788 1386 806
rect 1430 804 1436 805
rect 1430 800 1431 804
rect 1435 800 1436 804
rect 1430 799 1436 800
rect 1382 787 1388 788
rect 1382 783 1383 787
rect 1387 783 1388 787
rect 1382 782 1388 783
rect 1432 779 1434 799
rect 1504 788 1506 806
rect 1558 804 1564 805
rect 1558 800 1559 804
rect 1563 800 1564 804
rect 1766 803 1767 807
rect 1771 803 1772 807
rect 1766 802 1772 803
rect 1558 799 1564 800
rect 1502 787 1508 788
rect 1502 783 1503 787
rect 1507 783 1508 787
rect 1502 782 1508 783
rect 1560 779 1562 799
rect 1768 779 1770 802
rect 1808 791 1810 814
rect 1830 812 1831 816
rect 1835 812 1836 816
rect 1830 811 1836 812
rect 1832 791 1834 811
rect 1896 800 1898 890
rect 1982 885 1988 886
rect 1982 881 1983 885
rect 1987 881 1988 885
rect 1982 880 1988 881
rect 1984 859 1986 880
rect 1959 858 1963 859
rect 1959 853 1963 854
rect 1983 858 1987 859
rect 1983 853 1987 854
rect 1960 836 1962 853
rect 1958 835 1964 836
rect 1958 831 1959 835
rect 1963 831 1964 835
rect 1958 830 1964 831
rect 2040 828 2042 914
rect 2056 896 2058 914
rect 2152 905 2154 921
rect 2150 904 2156 905
rect 2150 900 2151 904
rect 2155 900 2156 904
rect 2150 899 2156 900
rect 2224 896 2226 938
rect 2312 927 2314 955
rect 2384 944 2386 962
rect 2406 960 2412 961
rect 2406 956 2407 960
rect 2411 956 2412 960
rect 2406 955 2412 956
rect 2382 943 2388 944
rect 2382 939 2383 943
rect 2387 939 2388 943
rect 2382 938 2388 939
rect 2408 927 2410 955
rect 2480 944 2482 962
rect 2510 960 2516 961
rect 2510 956 2511 960
rect 2515 956 2516 960
rect 2510 955 2516 956
rect 2622 960 2628 961
rect 2622 956 2623 960
rect 2627 956 2628 960
rect 2622 955 2628 956
rect 2478 943 2484 944
rect 2478 939 2479 943
rect 2483 939 2484 943
rect 2478 938 2484 939
rect 2512 927 2514 955
rect 2624 927 2626 955
rect 2696 944 2698 962
rect 2750 960 2756 961
rect 2750 956 2751 960
rect 2755 956 2756 960
rect 2750 955 2756 956
rect 2694 943 2700 944
rect 2694 939 2695 943
rect 2699 939 2700 943
rect 2694 938 2700 939
rect 2752 927 2754 955
rect 2824 928 2826 962
rect 2880 944 2882 1030
rect 2895 1002 2899 1003
rect 2895 997 2899 998
rect 3055 1002 3059 1003
rect 3055 997 3059 998
rect 3223 1002 3227 1003
rect 3223 997 3227 998
rect 3367 1002 3371 1003
rect 3367 997 3371 998
rect 2896 980 2898 997
rect 3056 980 3058 997
rect 3224 980 3226 997
rect 3368 980 3370 997
rect 2894 979 2900 980
rect 2894 975 2895 979
rect 2899 975 2900 979
rect 2894 974 2900 975
rect 3054 979 3060 980
rect 3054 975 3055 979
rect 3059 975 3060 979
rect 3054 974 3060 975
rect 3222 979 3228 980
rect 3222 975 3223 979
rect 3227 975 3228 979
rect 3222 974 3228 975
rect 3366 979 3372 980
rect 3366 975 3367 979
rect 3371 975 3372 979
rect 3366 974 3372 975
rect 3440 972 3442 1074
rect 3464 1067 3466 1094
rect 3463 1066 3467 1067
rect 3463 1061 3467 1062
rect 3464 1042 3466 1061
rect 3462 1041 3468 1042
rect 3462 1037 3463 1041
rect 3467 1037 3468 1041
rect 3462 1036 3468 1037
rect 3462 1024 3468 1025
rect 3462 1020 3463 1024
rect 3467 1020 3468 1024
rect 3462 1019 3468 1020
rect 3464 1003 3466 1019
rect 3463 1002 3467 1003
rect 3463 997 3467 998
rect 3464 981 3466 997
rect 3462 980 3468 981
rect 3462 976 3463 980
rect 3467 976 3468 980
rect 3462 975 3468 976
rect 3138 971 3144 972
rect 2966 967 2972 968
rect 2966 963 2967 967
rect 2971 963 2972 967
rect 2966 962 2972 963
rect 3126 967 3132 968
rect 3126 963 3127 967
rect 3131 963 3132 967
rect 3138 967 3139 971
rect 3143 967 3144 971
rect 3138 966 3144 967
rect 3438 971 3444 972
rect 3438 967 3439 971
rect 3443 967 3444 971
rect 3438 966 3444 967
rect 3126 962 3132 963
rect 2894 960 2900 961
rect 2894 956 2895 960
rect 2899 956 2900 960
rect 2894 955 2900 956
rect 2878 943 2884 944
rect 2878 939 2879 943
rect 2883 939 2884 943
rect 2878 938 2884 939
rect 2822 927 2828 928
rect 2896 927 2898 955
rect 2968 944 2970 962
rect 3054 960 3060 961
rect 3054 956 3055 960
rect 3059 956 3060 960
rect 3054 955 3060 956
rect 2966 943 2972 944
rect 2966 939 2967 943
rect 2971 939 2972 943
rect 2966 938 2972 939
rect 3056 927 3058 955
rect 3128 944 3130 962
rect 3140 952 3142 966
rect 3462 963 3468 964
rect 3222 960 3228 961
rect 3222 956 3223 960
rect 3227 956 3228 960
rect 3222 955 3228 956
rect 3366 960 3372 961
rect 3366 956 3367 960
rect 3371 956 3372 960
rect 3462 959 3463 963
rect 3467 959 3468 963
rect 3462 958 3468 959
rect 3366 955 3372 956
rect 3138 951 3144 952
rect 3138 947 3139 951
rect 3143 947 3144 951
rect 3138 946 3144 947
rect 3126 943 3132 944
rect 3126 939 3127 943
rect 3131 939 3132 943
rect 3126 938 3132 939
rect 3224 927 3226 955
rect 3368 927 3370 955
rect 3430 943 3436 944
rect 3430 939 3431 943
rect 3435 939 3436 943
rect 3430 938 3436 939
rect 2311 926 2315 927
rect 2311 921 2315 922
rect 2327 926 2331 927
rect 2327 921 2331 922
rect 2407 926 2411 927
rect 2407 921 2411 922
rect 2511 926 2515 927
rect 2511 921 2515 922
rect 2519 926 2523 927
rect 2519 921 2523 922
rect 2623 926 2627 927
rect 2623 921 2627 922
rect 2719 926 2723 927
rect 2719 921 2723 922
rect 2751 926 2755 927
rect 2822 923 2823 927
rect 2827 923 2828 927
rect 2822 922 2828 923
rect 2895 926 2899 927
rect 2751 921 2755 922
rect 2895 921 2899 922
rect 2935 926 2939 927
rect 2935 921 2939 922
rect 3055 926 3059 927
rect 3055 921 3059 922
rect 3159 926 3163 927
rect 3159 921 3163 922
rect 3223 926 3227 927
rect 3223 921 3227 922
rect 3367 926 3371 927
rect 3367 921 3371 922
rect 2328 905 2330 921
rect 2520 905 2522 921
rect 2598 919 2604 920
rect 2598 915 2599 919
rect 2603 915 2604 919
rect 2598 914 2604 915
rect 2326 904 2332 905
rect 2326 900 2327 904
rect 2331 900 2332 904
rect 2326 899 2332 900
rect 2518 904 2524 905
rect 2518 900 2519 904
rect 2523 900 2524 904
rect 2518 899 2524 900
rect 2600 896 2602 914
rect 2720 905 2722 921
rect 2936 905 2938 921
rect 3006 919 3012 920
rect 3006 915 3007 919
rect 3011 915 3012 919
rect 3006 914 3012 915
rect 2718 904 2724 905
rect 2718 900 2719 904
rect 2723 900 2724 904
rect 2718 899 2724 900
rect 2934 904 2940 905
rect 2934 900 2935 904
rect 2939 900 2940 904
rect 2934 899 2940 900
rect 3008 896 3010 914
rect 3160 905 3162 921
rect 3368 905 3370 921
rect 3158 904 3164 905
rect 3158 900 3159 904
rect 3163 900 3164 904
rect 3158 899 3164 900
rect 3366 904 3372 905
rect 3366 900 3367 904
rect 3371 900 3372 904
rect 3366 899 3372 900
rect 3432 896 3434 938
rect 3464 927 3466 958
rect 3463 926 3467 927
rect 3463 921 3467 922
rect 3438 919 3444 920
rect 3438 915 3439 919
rect 3443 915 3444 919
rect 3438 914 3444 915
rect 2054 895 2060 896
rect 2054 891 2055 895
rect 2059 891 2060 895
rect 2054 890 2060 891
rect 2222 895 2228 896
rect 2222 891 2223 895
rect 2227 891 2228 895
rect 2222 890 2228 891
rect 2398 895 2404 896
rect 2398 891 2399 895
rect 2403 891 2404 895
rect 2398 890 2404 891
rect 2598 895 2604 896
rect 2598 891 2599 895
rect 2603 891 2604 895
rect 2598 890 2604 891
rect 3006 895 3012 896
rect 3006 891 3007 895
rect 3011 891 3012 895
rect 3006 890 3012 891
rect 3430 895 3436 896
rect 3430 891 3431 895
rect 3435 891 3436 895
rect 3430 890 3436 891
rect 2150 885 2156 886
rect 2150 881 2151 885
rect 2155 881 2156 885
rect 2150 880 2156 881
rect 2326 885 2332 886
rect 2326 881 2327 885
rect 2331 881 2332 885
rect 2326 880 2332 881
rect 2152 859 2154 880
rect 2328 859 2330 880
rect 2087 858 2091 859
rect 2087 853 2091 854
rect 2151 858 2155 859
rect 2151 853 2155 854
rect 2207 858 2211 859
rect 2207 853 2211 854
rect 2327 858 2331 859
rect 2327 853 2331 854
rect 2088 836 2090 853
rect 2208 836 2210 853
rect 2328 836 2330 853
rect 2086 835 2092 836
rect 2086 831 2087 835
rect 2091 831 2092 835
rect 2086 830 2092 831
rect 2206 835 2212 836
rect 2206 831 2207 835
rect 2211 831 2212 835
rect 2206 830 2212 831
rect 2326 835 2332 836
rect 2326 831 2327 835
rect 2331 831 2332 835
rect 2326 830 2332 831
rect 2038 827 2044 828
rect 1902 823 1908 824
rect 1902 819 1903 823
rect 1907 819 1908 823
rect 1902 818 1908 819
rect 2030 823 2036 824
rect 2030 819 2031 823
rect 2035 819 2036 823
rect 2038 823 2039 827
rect 2043 823 2044 827
rect 2286 827 2292 828
rect 2038 822 2044 823
rect 2278 823 2284 824
rect 2030 818 2036 819
rect 2278 819 2279 823
rect 2283 819 2284 823
rect 2286 823 2287 827
rect 2291 823 2292 827
rect 2286 822 2292 823
rect 2278 818 2284 819
rect 1904 800 1906 818
rect 1958 816 1964 817
rect 1958 812 1959 816
rect 1963 812 1964 816
rect 1958 811 1964 812
rect 1894 799 1900 800
rect 1894 795 1895 799
rect 1899 795 1900 799
rect 1894 794 1900 795
rect 1902 799 1908 800
rect 1902 795 1903 799
rect 1907 795 1908 799
rect 1902 794 1908 795
rect 1960 791 1962 811
rect 1807 790 1811 791
rect 1807 785 1811 786
rect 1831 790 1835 791
rect 1831 785 1835 786
rect 1879 790 1883 791
rect 1879 785 1883 786
rect 1959 790 1963 791
rect 1959 785 1963 786
rect 2015 790 2019 791
rect 2015 785 2019 786
rect 1287 778 1291 779
rect 1287 773 1291 774
rect 1311 778 1315 779
rect 1311 773 1315 774
rect 1415 778 1419 779
rect 1415 773 1419 774
rect 1431 778 1435 779
rect 1431 773 1435 774
rect 1559 778 1563 779
rect 1559 773 1563 774
rect 1767 778 1771 779
rect 1767 773 1771 774
rect 1238 771 1244 772
rect 1238 767 1239 771
rect 1243 767 1244 771
rect 1238 766 1244 767
rect 1240 748 1242 766
rect 1288 757 1290 773
rect 1366 771 1372 772
rect 1366 767 1367 771
rect 1371 767 1372 771
rect 1366 766 1372 767
rect 1286 756 1292 757
rect 1286 752 1287 756
rect 1291 752 1292 756
rect 1286 751 1292 752
rect 1368 748 1370 766
rect 1416 757 1418 773
rect 1414 756 1420 757
rect 1414 752 1415 756
rect 1419 752 1420 756
rect 1768 754 1770 773
rect 1808 766 1810 785
rect 1880 769 1882 785
rect 2016 769 2018 785
rect 2032 784 2034 818
rect 2086 816 2092 817
rect 2086 812 2087 816
rect 2091 812 2092 816
rect 2086 811 2092 812
rect 2206 816 2212 817
rect 2206 812 2207 816
rect 2211 812 2212 816
rect 2206 811 2212 812
rect 2088 791 2090 811
rect 2208 791 2210 811
rect 2280 800 2282 818
rect 2288 808 2290 822
rect 2326 816 2332 817
rect 2326 812 2327 816
rect 2331 812 2332 816
rect 2326 811 2332 812
rect 2286 807 2292 808
rect 2286 803 2287 807
rect 2291 803 2292 807
rect 2286 802 2292 803
rect 2222 799 2228 800
rect 2222 795 2223 799
rect 2227 795 2228 799
rect 2222 794 2228 795
rect 2278 799 2284 800
rect 2278 795 2279 799
rect 2283 795 2284 799
rect 2278 794 2284 795
rect 2087 790 2091 791
rect 2087 785 2091 786
rect 2151 790 2155 791
rect 2151 785 2155 786
rect 2207 790 2211 791
rect 2207 785 2211 786
rect 2030 783 2036 784
rect 2030 779 2031 783
rect 2035 779 2036 783
rect 2030 778 2036 779
rect 2152 769 2154 785
rect 1878 768 1884 769
rect 1806 765 1812 766
rect 1806 761 1807 765
rect 1811 761 1812 765
rect 1878 764 1879 768
rect 1883 764 1884 768
rect 1878 763 1884 764
rect 2014 768 2020 769
rect 2014 764 2015 768
rect 2019 764 2020 768
rect 2014 763 2020 764
rect 2150 768 2156 769
rect 2150 764 2151 768
rect 2155 764 2156 768
rect 2150 763 2156 764
rect 1806 760 1812 761
rect 2224 760 2226 794
rect 2328 791 2330 811
rect 2400 800 2402 890
rect 2518 885 2524 886
rect 2518 881 2519 885
rect 2523 881 2524 885
rect 2518 880 2524 881
rect 2718 885 2724 886
rect 2718 881 2719 885
rect 2723 881 2724 885
rect 2718 880 2724 881
rect 2934 885 2940 886
rect 2934 881 2935 885
rect 2939 881 2940 885
rect 2934 880 2940 881
rect 3158 885 3164 886
rect 3158 881 3159 885
rect 3163 881 3164 885
rect 3158 880 3164 881
rect 3366 885 3372 886
rect 3366 881 3367 885
rect 3371 881 3372 885
rect 3366 880 3372 881
rect 2520 859 2522 880
rect 2720 859 2722 880
rect 2936 859 2938 880
rect 3160 859 3162 880
rect 3368 859 3370 880
rect 2463 858 2467 859
rect 2463 853 2467 854
rect 2519 858 2523 859
rect 2519 853 2523 854
rect 2615 858 2619 859
rect 2615 853 2619 854
rect 2719 858 2723 859
rect 2719 853 2723 854
rect 2791 858 2795 859
rect 2791 853 2795 854
rect 2935 858 2939 859
rect 2935 853 2939 854
rect 2983 858 2987 859
rect 2983 853 2987 854
rect 3159 858 3163 859
rect 3159 853 3163 854
rect 3183 858 3187 859
rect 3183 853 3187 854
rect 3367 858 3371 859
rect 3367 853 3371 854
rect 2464 836 2466 853
rect 2616 836 2618 853
rect 2792 836 2794 853
rect 2984 836 2986 853
rect 3184 836 3186 853
rect 3368 836 3370 853
rect 2462 835 2468 836
rect 2462 831 2463 835
rect 2467 831 2468 835
rect 2462 830 2468 831
rect 2614 835 2620 836
rect 2614 831 2615 835
rect 2619 831 2620 835
rect 2614 830 2620 831
rect 2790 835 2796 836
rect 2790 831 2791 835
rect 2795 831 2796 835
rect 2790 830 2796 831
rect 2982 835 2988 836
rect 2982 831 2983 835
rect 2987 831 2988 835
rect 2982 830 2988 831
rect 3182 835 3188 836
rect 3182 831 3183 835
rect 3187 831 3188 835
rect 3182 830 3188 831
rect 3366 835 3372 836
rect 3366 831 3367 835
rect 3371 831 3372 835
rect 3366 830 3372 831
rect 3440 828 3442 914
rect 3464 902 3466 921
rect 3462 901 3468 902
rect 3462 897 3463 901
rect 3467 897 3468 901
rect 3462 896 3468 897
rect 3462 884 3468 885
rect 3462 880 3463 884
rect 3467 880 3468 884
rect 3462 879 3468 880
rect 3464 859 3466 879
rect 3463 858 3467 859
rect 3463 853 3467 854
rect 3464 837 3466 853
rect 3462 836 3468 837
rect 3462 832 3463 836
rect 3467 832 3468 836
rect 3462 831 3468 832
rect 3138 827 3144 828
rect 2534 823 2540 824
rect 2534 819 2535 823
rect 2539 819 2540 823
rect 2534 818 2540 819
rect 2686 823 2692 824
rect 2686 819 2687 823
rect 2691 819 2692 823
rect 2686 818 2692 819
rect 2862 823 2868 824
rect 2862 819 2863 823
rect 2867 819 2868 823
rect 2862 818 2868 819
rect 3054 823 3060 824
rect 3054 819 3055 823
rect 3059 819 3060 823
rect 3138 823 3139 827
rect 3143 823 3144 827
rect 3138 822 3144 823
rect 3438 827 3444 828
rect 3438 823 3439 827
rect 3443 823 3444 827
rect 3438 822 3444 823
rect 3054 818 3060 819
rect 2462 816 2468 817
rect 2462 812 2463 816
rect 2467 812 2468 816
rect 2462 811 2468 812
rect 2398 799 2404 800
rect 2398 795 2399 799
rect 2403 795 2404 799
rect 2398 794 2404 795
rect 2464 791 2466 811
rect 2536 800 2538 818
rect 2614 816 2620 817
rect 2614 812 2615 816
rect 2619 812 2620 816
rect 2614 811 2620 812
rect 2534 799 2540 800
rect 2534 795 2535 799
rect 2539 795 2540 799
rect 2534 794 2540 795
rect 2616 791 2618 811
rect 2688 800 2690 818
rect 2790 816 2796 817
rect 2790 812 2791 816
rect 2795 812 2796 816
rect 2790 811 2796 812
rect 2686 799 2692 800
rect 2686 795 2687 799
rect 2691 795 2692 799
rect 2686 794 2692 795
rect 2792 791 2794 811
rect 2864 800 2866 818
rect 2982 816 2988 817
rect 2982 812 2983 816
rect 2987 812 2988 816
rect 2982 811 2988 812
rect 2862 799 2868 800
rect 2862 795 2863 799
rect 2867 795 2868 799
rect 2862 794 2868 795
rect 2984 791 2986 811
rect 3056 800 3058 818
rect 3054 799 3060 800
rect 3054 795 3055 799
rect 3059 795 3060 799
rect 3054 794 3060 795
rect 3140 792 3142 822
rect 3462 819 3468 820
rect 3182 816 3188 817
rect 3182 812 3183 816
rect 3187 812 3188 816
rect 3182 811 3188 812
rect 3366 816 3372 817
rect 3366 812 3367 816
rect 3371 812 3372 816
rect 3462 815 3463 819
rect 3467 815 3468 819
rect 3462 814 3468 815
rect 3366 811 3372 812
rect 3138 791 3144 792
rect 3184 791 3186 811
rect 3368 791 3370 811
rect 3430 799 3436 800
rect 3430 795 3431 799
rect 3435 795 3436 799
rect 3430 794 3436 795
rect 2287 790 2291 791
rect 2287 785 2291 786
rect 2327 790 2331 791
rect 2327 785 2331 786
rect 2423 790 2427 791
rect 2423 785 2427 786
rect 2463 790 2467 791
rect 2463 785 2467 786
rect 2559 790 2563 791
rect 2559 785 2563 786
rect 2615 790 2619 791
rect 2615 785 2619 786
rect 2711 790 2715 791
rect 2711 785 2715 786
rect 2791 790 2795 791
rect 2791 785 2795 786
rect 2871 790 2875 791
rect 2871 785 2875 786
rect 2983 790 2987 791
rect 2983 785 2987 786
rect 3039 790 3043 791
rect 3138 787 3139 791
rect 3143 787 3144 791
rect 3138 786 3144 787
rect 3183 790 3187 791
rect 3039 785 3043 786
rect 3183 785 3187 786
rect 3215 790 3219 791
rect 3215 785 3219 786
rect 3367 790 3371 791
rect 3367 785 3371 786
rect 2230 783 2236 784
rect 2230 779 2231 783
rect 2235 779 2236 783
rect 2230 778 2236 779
rect 2232 760 2234 778
rect 2288 769 2290 785
rect 2366 783 2372 784
rect 2366 779 2367 783
rect 2371 779 2372 783
rect 2366 778 2372 779
rect 2286 768 2292 769
rect 2286 764 2287 768
rect 2291 764 2292 768
rect 2286 763 2292 764
rect 2368 760 2370 778
rect 2424 769 2426 785
rect 2486 783 2492 784
rect 2486 779 2487 783
rect 2491 779 2492 783
rect 2486 778 2492 779
rect 2422 768 2428 769
rect 2422 764 2423 768
rect 2427 764 2428 768
rect 2422 763 2428 764
rect 2222 759 2228 760
rect 2222 755 2223 759
rect 2227 755 2228 759
rect 2222 754 2228 755
rect 2230 759 2236 760
rect 2230 755 2231 759
rect 2235 755 2236 759
rect 2230 754 2236 755
rect 2366 759 2372 760
rect 2366 755 2367 759
rect 2371 755 2372 759
rect 2366 754 2372 755
rect 1414 751 1420 752
rect 1766 753 1772 754
rect 1766 749 1767 753
rect 1771 749 1772 753
rect 1962 751 1968 752
rect 1878 749 1884 750
rect 1766 748 1772 749
rect 1806 748 1812 749
rect 750 747 756 748
rect 750 743 751 747
rect 755 743 756 747
rect 750 742 756 743
rect 758 747 764 748
rect 758 743 759 747
rect 763 743 764 747
rect 758 742 764 743
rect 990 747 996 748
rect 990 743 991 747
rect 995 743 996 747
rect 990 742 996 743
rect 1230 747 1236 748
rect 1230 743 1231 747
rect 1235 743 1236 747
rect 1230 742 1236 743
rect 1238 747 1244 748
rect 1238 743 1239 747
rect 1243 743 1244 747
rect 1238 742 1244 743
rect 1366 747 1372 748
rect 1366 743 1367 747
rect 1371 743 1372 747
rect 1806 744 1807 748
rect 1811 744 1812 748
rect 1878 745 1879 749
rect 1883 745 1884 749
rect 1962 747 1963 751
rect 1967 747 1968 751
rect 1962 746 1968 747
rect 2014 749 2020 750
rect 1878 744 1884 745
rect 1806 743 1812 744
rect 1366 742 1372 743
rect 994 739 1000 740
rect 678 737 684 738
rect 678 733 679 737
rect 683 733 684 737
rect 678 732 684 733
rect 790 737 796 738
rect 790 733 791 737
rect 795 733 796 737
rect 790 732 796 733
rect 910 737 916 738
rect 910 733 911 737
rect 915 733 916 737
rect 994 735 995 739
rect 999 735 1000 739
rect 994 734 1000 735
rect 1030 737 1036 738
rect 910 732 916 733
rect 680 707 682 732
rect 792 707 794 732
rect 912 707 914 732
rect 679 706 683 707
rect 679 701 683 702
rect 695 706 699 707
rect 695 701 699 702
rect 791 706 795 707
rect 791 701 795 702
rect 831 706 835 707
rect 831 701 835 702
rect 911 706 915 707
rect 911 701 915 702
rect 983 706 987 707
rect 983 701 987 702
rect 696 684 698 701
rect 832 684 834 701
rect 984 684 986 701
rect 694 683 700 684
rect 694 679 695 683
rect 699 679 700 683
rect 694 678 700 679
rect 830 683 836 684
rect 830 679 831 683
rect 835 679 836 683
rect 830 678 836 679
rect 982 683 988 684
rect 982 679 983 683
rect 987 679 988 683
rect 982 678 988 679
rect 654 675 660 676
rect 318 671 324 672
rect 110 667 116 668
rect 110 663 111 667
rect 115 663 116 667
rect 318 667 319 671
rect 323 667 324 671
rect 318 666 324 667
rect 414 671 420 672
rect 414 667 415 671
rect 419 667 420 671
rect 414 666 420 667
rect 526 671 532 672
rect 526 667 527 671
rect 531 667 532 671
rect 526 666 532 667
rect 638 671 644 672
rect 638 667 639 671
rect 643 667 644 671
rect 654 671 655 675
rect 659 671 660 675
rect 654 670 660 671
rect 822 675 828 676
rect 822 671 823 675
rect 827 671 828 675
rect 822 670 828 671
rect 910 675 916 676
rect 910 671 911 675
rect 915 671 916 675
rect 910 670 916 671
rect 638 666 644 667
rect 110 662 116 663
rect 246 664 252 665
rect 112 639 114 662
rect 246 660 247 664
rect 251 660 252 664
rect 246 659 252 660
rect 248 639 250 659
rect 320 648 322 666
rect 342 664 348 665
rect 342 660 343 664
rect 347 660 348 664
rect 342 659 348 660
rect 318 647 324 648
rect 318 643 319 647
rect 323 643 324 647
rect 318 642 324 643
rect 344 639 346 659
rect 416 648 418 666
rect 454 664 460 665
rect 454 660 455 664
rect 459 660 460 664
rect 454 659 460 660
rect 414 647 420 648
rect 414 643 415 647
rect 419 643 420 647
rect 414 642 420 643
rect 456 639 458 659
rect 528 648 530 666
rect 566 664 572 665
rect 566 660 567 664
rect 571 660 572 664
rect 566 659 572 660
rect 526 647 532 648
rect 526 643 527 647
rect 531 643 532 647
rect 526 642 532 643
rect 568 639 570 659
rect 640 648 642 666
rect 694 664 700 665
rect 694 660 695 664
rect 699 660 700 664
rect 694 659 700 660
rect 638 647 644 648
rect 638 643 639 647
rect 643 643 644 647
rect 638 642 644 643
rect 696 639 698 659
rect 111 638 115 639
rect 111 633 115 634
rect 135 638 139 639
rect 135 633 139 634
rect 231 638 235 639
rect 231 633 235 634
rect 247 638 251 639
rect 247 633 251 634
rect 343 638 347 639
rect 343 633 347 634
rect 359 638 363 639
rect 359 633 363 634
rect 455 638 459 639
rect 455 633 459 634
rect 487 638 491 639
rect 487 633 491 634
rect 567 638 571 639
rect 567 633 571 634
rect 623 638 627 639
rect 623 633 627 634
rect 695 638 699 639
rect 695 633 699 634
rect 767 638 771 639
rect 767 633 771 634
rect 112 614 114 633
rect 136 617 138 633
rect 198 631 204 632
rect 198 627 199 631
rect 203 627 204 631
rect 198 626 204 627
rect 206 631 212 632
rect 206 627 207 631
rect 211 627 212 631
rect 206 626 212 627
rect 134 616 140 617
rect 110 613 116 614
rect 110 609 111 613
rect 115 609 116 613
rect 134 612 135 616
rect 139 612 140 616
rect 134 611 140 612
rect 110 608 116 609
rect 134 597 140 598
rect 110 596 116 597
rect 110 592 111 596
rect 115 592 116 596
rect 134 593 135 597
rect 139 593 140 597
rect 134 592 140 593
rect 110 591 116 592
rect 112 571 114 591
rect 136 571 138 592
rect 111 570 115 571
rect 111 565 115 566
rect 135 570 139 571
rect 135 565 139 566
rect 112 549 114 565
rect 110 548 116 549
rect 136 548 138 565
rect 110 544 111 548
rect 115 544 116 548
rect 110 543 116 544
rect 134 547 140 548
rect 134 543 135 547
rect 139 543 140 547
rect 200 544 202 626
rect 208 608 210 626
rect 232 617 234 633
rect 302 631 308 632
rect 302 627 303 631
rect 307 627 308 631
rect 302 626 308 627
rect 230 616 236 617
rect 230 612 231 616
rect 235 612 236 616
rect 230 611 236 612
rect 304 608 306 626
rect 360 617 362 633
rect 430 631 436 632
rect 430 627 431 631
rect 435 627 436 631
rect 430 626 436 627
rect 358 616 364 617
rect 358 612 359 616
rect 363 612 364 616
rect 358 611 364 612
rect 432 608 434 626
rect 488 617 490 633
rect 558 631 564 632
rect 558 627 559 631
rect 563 627 564 631
rect 558 626 564 627
rect 486 616 492 617
rect 486 612 487 616
rect 491 612 492 616
rect 486 611 492 612
rect 560 608 562 626
rect 624 617 626 633
rect 768 617 770 633
rect 824 632 826 670
rect 830 664 836 665
rect 830 660 831 664
rect 835 660 836 664
rect 830 659 836 660
rect 832 639 834 659
rect 912 648 914 670
rect 982 664 988 665
rect 982 660 983 664
rect 987 660 988 664
rect 982 659 988 660
rect 910 647 916 648
rect 910 643 911 647
rect 915 643 916 647
rect 910 642 916 643
rect 984 639 986 659
rect 996 648 998 734
rect 1030 733 1031 737
rect 1035 733 1036 737
rect 1030 732 1036 733
rect 1158 737 1164 738
rect 1158 733 1159 737
rect 1163 733 1164 737
rect 1158 732 1164 733
rect 1286 737 1292 738
rect 1286 733 1287 737
rect 1291 733 1292 737
rect 1286 732 1292 733
rect 1414 737 1420 738
rect 1414 733 1415 737
rect 1419 733 1420 737
rect 1414 732 1420 733
rect 1766 736 1772 737
rect 1766 732 1767 736
rect 1771 732 1772 736
rect 1032 707 1034 732
rect 1160 707 1162 732
rect 1288 707 1290 732
rect 1416 707 1418 732
rect 1766 731 1772 732
rect 1768 707 1770 731
rect 1808 723 1810 743
rect 1880 723 1882 744
rect 1807 722 1811 723
rect 1807 717 1811 718
rect 1831 722 1835 723
rect 1831 717 1835 718
rect 1879 722 1883 723
rect 1879 717 1883 718
rect 1951 722 1955 723
rect 1951 717 1955 718
rect 1031 706 1035 707
rect 1031 701 1035 702
rect 1151 706 1155 707
rect 1151 701 1155 702
rect 1159 706 1163 707
rect 1159 701 1163 702
rect 1287 706 1291 707
rect 1287 701 1291 702
rect 1327 706 1331 707
rect 1327 701 1331 702
rect 1415 706 1419 707
rect 1415 701 1419 702
rect 1511 706 1515 707
rect 1511 701 1515 702
rect 1671 706 1675 707
rect 1671 701 1675 702
rect 1767 706 1771 707
rect 1767 701 1771 702
rect 1808 701 1810 717
rect 1152 684 1154 701
rect 1328 684 1330 701
rect 1512 684 1514 701
rect 1672 684 1674 701
rect 1750 691 1756 692
rect 1750 687 1751 691
rect 1755 687 1756 691
rect 1750 686 1756 687
rect 1150 683 1156 684
rect 1150 679 1151 683
rect 1155 679 1156 683
rect 1150 678 1156 679
rect 1326 683 1332 684
rect 1326 679 1327 683
rect 1331 679 1332 683
rect 1326 678 1332 679
rect 1510 683 1516 684
rect 1510 679 1511 683
rect 1515 679 1516 683
rect 1510 678 1516 679
rect 1670 683 1676 684
rect 1670 679 1671 683
rect 1675 679 1676 683
rect 1670 678 1676 679
rect 1294 671 1300 672
rect 1294 667 1295 671
rect 1299 667 1300 671
rect 1294 666 1300 667
rect 1398 671 1404 672
rect 1398 667 1399 671
rect 1403 667 1404 671
rect 1398 666 1404 667
rect 1742 671 1748 672
rect 1742 667 1743 671
rect 1747 667 1748 671
rect 1742 666 1748 667
rect 1150 664 1156 665
rect 1150 660 1151 664
rect 1155 660 1156 664
rect 1150 659 1156 660
rect 994 647 1000 648
rect 994 643 995 647
rect 999 643 1000 647
rect 994 642 1000 643
rect 1152 639 1154 659
rect 1296 648 1298 666
rect 1326 664 1332 665
rect 1326 660 1327 664
rect 1331 660 1332 664
rect 1326 659 1332 660
rect 1286 647 1292 648
rect 1286 643 1287 647
rect 1291 643 1292 647
rect 1286 642 1292 643
rect 1294 647 1300 648
rect 1294 643 1295 647
rect 1299 643 1300 647
rect 1294 642 1300 643
rect 831 638 835 639
rect 831 633 835 634
rect 911 638 915 639
rect 911 633 915 634
rect 983 638 987 639
rect 983 633 987 634
rect 1055 638 1059 639
rect 1055 633 1059 634
rect 1151 638 1155 639
rect 1151 633 1155 634
rect 1207 638 1211 639
rect 1207 633 1211 634
rect 822 631 828 632
rect 822 627 823 631
rect 827 627 828 631
rect 822 626 828 627
rect 912 617 914 633
rect 1056 617 1058 633
rect 1110 631 1116 632
rect 1110 627 1111 631
rect 1115 627 1116 631
rect 1110 626 1116 627
rect 1126 631 1132 632
rect 1126 627 1127 631
rect 1131 627 1132 631
rect 1126 626 1132 627
rect 622 616 628 617
rect 622 612 623 616
rect 627 612 628 616
rect 622 611 628 612
rect 766 616 772 617
rect 766 612 767 616
rect 771 612 772 616
rect 766 611 772 612
rect 910 616 916 617
rect 910 612 911 616
rect 915 612 916 616
rect 910 611 916 612
rect 1054 616 1060 617
rect 1054 612 1055 616
rect 1059 612 1060 616
rect 1054 611 1060 612
rect 206 607 212 608
rect 206 603 207 607
rect 211 603 212 607
rect 206 602 212 603
rect 302 607 308 608
rect 302 603 303 607
rect 307 603 308 607
rect 302 602 308 603
rect 430 607 436 608
rect 430 603 431 607
rect 435 603 436 607
rect 430 602 436 603
rect 558 607 564 608
rect 558 603 559 607
rect 563 603 564 607
rect 558 602 564 603
rect 982 607 988 608
rect 982 603 983 607
rect 987 603 988 607
rect 982 602 988 603
rect 230 597 236 598
rect 230 593 231 597
rect 235 593 236 597
rect 230 592 236 593
rect 358 597 364 598
rect 358 593 359 597
rect 363 593 364 597
rect 358 592 364 593
rect 486 597 492 598
rect 486 593 487 597
rect 491 593 492 597
rect 486 592 492 593
rect 622 597 628 598
rect 622 593 623 597
rect 627 593 628 597
rect 622 592 628 593
rect 766 597 772 598
rect 766 593 767 597
rect 771 593 772 597
rect 766 592 772 593
rect 910 597 916 598
rect 910 593 911 597
rect 915 593 916 597
rect 910 592 916 593
rect 232 571 234 592
rect 360 571 362 592
rect 488 571 490 592
rect 624 571 626 592
rect 768 571 770 592
rect 912 571 914 592
rect 231 570 235 571
rect 231 565 235 566
rect 247 570 251 571
rect 247 565 251 566
rect 359 570 363 571
rect 359 565 363 566
rect 407 570 411 571
rect 407 565 411 566
rect 487 570 491 571
rect 487 565 491 566
rect 583 570 587 571
rect 583 565 587 566
rect 623 570 627 571
rect 623 565 627 566
rect 767 570 771 571
rect 767 565 771 566
rect 911 570 915 571
rect 911 565 915 566
rect 951 570 955 571
rect 951 565 955 566
rect 248 548 250 565
rect 408 548 410 565
rect 584 548 586 565
rect 768 548 770 565
rect 952 548 954 565
rect 246 547 252 548
rect 134 542 140 543
rect 198 543 204 544
rect 198 539 199 543
rect 203 539 204 543
rect 246 543 247 547
rect 251 543 252 547
rect 246 542 252 543
rect 406 547 412 548
rect 406 543 407 547
rect 411 543 412 547
rect 406 542 412 543
rect 582 547 588 548
rect 582 543 583 547
rect 587 543 588 547
rect 582 542 588 543
rect 766 547 772 548
rect 766 543 767 547
rect 771 543 772 547
rect 766 542 772 543
rect 950 547 956 548
rect 950 543 951 547
rect 955 543 956 547
rect 950 542 956 543
rect 198 538 204 539
rect 214 539 220 540
rect 214 535 215 539
rect 219 535 220 539
rect 214 534 220 535
rect 326 539 332 540
rect 326 535 327 539
rect 331 535 332 539
rect 742 539 748 540
rect 326 534 332 535
rect 654 535 660 536
rect 110 531 116 532
rect 110 527 111 531
rect 115 527 116 531
rect 110 526 116 527
rect 134 528 140 529
rect 112 503 114 526
rect 134 524 135 528
rect 139 524 140 528
rect 134 523 140 524
rect 136 503 138 523
rect 216 512 218 534
rect 246 528 252 529
rect 246 524 247 528
rect 251 524 252 528
rect 246 523 252 524
rect 214 511 220 512
rect 214 507 215 511
rect 219 507 220 511
rect 214 506 220 507
rect 248 503 250 523
rect 328 512 330 534
rect 654 531 655 535
rect 659 531 660 535
rect 742 535 743 539
rect 747 535 748 539
rect 742 534 748 535
rect 654 530 660 531
rect 406 528 412 529
rect 406 524 407 528
rect 411 524 412 528
rect 406 523 412 524
rect 582 528 588 529
rect 582 524 583 528
rect 587 524 588 528
rect 582 523 588 524
rect 326 511 332 512
rect 326 507 327 511
rect 331 507 332 511
rect 326 506 332 507
rect 408 503 410 523
rect 584 503 586 523
rect 656 512 658 530
rect 744 520 746 534
rect 766 528 772 529
rect 766 524 767 528
rect 771 524 772 528
rect 766 523 772 524
rect 950 528 956 529
rect 950 524 951 528
rect 955 524 956 528
rect 950 523 956 524
rect 742 519 748 520
rect 742 515 743 519
rect 747 515 748 519
rect 742 514 748 515
rect 634 511 640 512
rect 634 507 635 511
rect 639 507 640 511
rect 634 506 640 507
rect 654 511 660 512
rect 654 507 655 511
rect 659 507 660 511
rect 654 506 660 507
rect 111 502 115 503
rect 111 497 115 498
rect 135 502 139 503
rect 135 497 139 498
rect 247 502 251 503
rect 247 497 251 498
rect 399 502 403 503
rect 399 497 403 498
rect 407 502 411 503
rect 407 497 411 498
rect 567 502 571 503
rect 567 497 571 498
rect 583 502 587 503
rect 583 497 587 498
rect 112 478 114 497
rect 248 481 250 497
rect 318 495 324 496
rect 318 491 319 495
rect 323 491 324 495
rect 318 490 324 491
rect 246 480 252 481
rect 110 477 116 478
rect 110 473 111 477
rect 115 473 116 477
rect 246 476 247 480
rect 251 476 252 480
rect 246 475 252 476
rect 110 472 116 473
rect 320 472 322 490
rect 400 481 402 497
rect 470 495 476 496
rect 470 491 471 495
rect 475 491 476 495
rect 470 490 476 491
rect 398 480 404 481
rect 398 476 399 480
rect 403 476 404 480
rect 398 475 404 476
rect 472 472 474 490
rect 568 481 570 497
rect 566 480 572 481
rect 566 476 567 480
rect 571 476 572 480
rect 566 475 572 476
rect 636 472 638 506
rect 768 503 770 523
rect 952 503 954 523
rect 984 512 986 602
rect 1054 597 1060 598
rect 1054 593 1055 597
rect 1059 593 1060 597
rect 1054 592 1060 593
rect 1056 571 1058 592
rect 1055 570 1059 571
rect 1055 565 1059 566
rect 1112 540 1114 626
rect 1128 608 1130 626
rect 1208 617 1210 633
rect 1278 631 1284 632
rect 1278 627 1279 631
rect 1283 627 1284 631
rect 1278 626 1284 627
rect 1206 616 1212 617
rect 1206 612 1207 616
rect 1211 612 1212 616
rect 1206 611 1212 612
rect 1280 608 1282 626
rect 1288 608 1290 642
rect 1328 639 1330 659
rect 1400 648 1402 666
rect 1510 664 1516 665
rect 1510 660 1511 664
rect 1515 660 1516 664
rect 1510 659 1516 660
rect 1670 664 1676 665
rect 1670 660 1671 664
rect 1675 660 1676 664
rect 1670 659 1676 660
rect 1398 647 1404 648
rect 1398 643 1399 647
rect 1403 643 1404 647
rect 1398 642 1404 643
rect 1512 639 1514 659
rect 1672 639 1674 659
rect 1327 638 1331 639
rect 1327 633 1331 634
rect 1367 638 1371 639
rect 1367 633 1371 634
rect 1511 638 1515 639
rect 1511 633 1515 634
rect 1527 638 1531 639
rect 1527 633 1531 634
rect 1671 638 1675 639
rect 1671 633 1675 634
rect 1368 617 1370 633
rect 1528 617 1530 633
rect 1606 631 1612 632
rect 1606 627 1607 631
rect 1611 627 1612 631
rect 1606 626 1612 627
rect 1366 616 1372 617
rect 1366 612 1367 616
rect 1371 612 1372 616
rect 1366 611 1372 612
rect 1526 616 1532 617
rect 1526 612 1527 616
rect 1531 612 1532 616
rect 1526 611 1532 612
rect 1608 608 1610 626
rect 1672 617 1674 633
rect 1744 632 1746 666
rect 1752 648 1754 686
rect 1768 685 1770 701
rect 1806 700 1812 701
rect 1832 700 1834 717
rect 1952 700 1954 717
rect 1806 696 1807 700
rect 1811 696 1812 700
rect 1806 695 1812 696
rect 1830 699 1836 700
rect 1830 695 1831 699
rect 1835 695 1836 699
rect 1830 694 1836 695
rect 1950 699 1956 700
rect 1950 695 1951 699
rect 1955 695 1956 699
rect 1950 694 1956 695
rect 1910 691 1916 692
rect 1910 687 1911 691
rect 1915 687 1916 691
rect 1910 686 1916 687
rect 1766 684 1772 685
rect 1766 680 1767 684
rect 1771 680 1772 684
rect 1766 679 1772 680
rect 1806 683 1812 684
rect 1806 679 1807 683
rect 1811 679 1812 683
rect 1806 678 1812 679
rect 1830 680 1836 681
rect 1766 667 1772 668
rect 1766 663 1767 667
rect 1771 663 1772 667
rect 1766 662 1772 663
rect 1750 647 1756 648
rect 1750 643 1751 647
rect 1755 643 1756 647
rect 1750 642 1756 643
rect 1768 639 1770 662
rect 1808 659 1810 678
rect 1830 676 1831 680
rect 1835 676 1836 680
rect 1830 675 1836 676
rect 1832 659 1834 675
rect 1912 664 1914 686
rect 1950 680 1956 681
rect 1950 676 1951 680
rect 1955 676 1956 680
rect 1950 675 1956 676
rect 1910 663 1916 664
rect 1910 659 1911 663
rect 1915 659 1916 663
rect 1952 659 1954 675
rect 1964 664 1966 746
rect 2014 745 2015 749
rect 2019 745 2020 749
rect 2014 744 2020 745
rect 2150 749 2156 750
rect 2150 745 2151 749
rect 2155 745 2156 749
rect 2150 744 2156 745
rect 2286 749 2292 750
rect 2286 745 2287 749
rect 2291 745 2292 749
rect 2286 744 2292 745
rect 2422 749 2428 750
rect 2422 745 2423 749
rect 2427 745 2428 749
rect 2422 744 2428 745
rect 2016 723 2018 744
rect 2152 723 2154 744
rect 2288 723 2290 744
rect 2424 723 2426 744
rect 2015 722 2019 723
rect 2015 717 2019 718
rect 2103 722 2107 723
rect 2103 717 2107 718
rect 2151 722 2155 723
rect 2151 717 2155 718
rect 2263 722 2267 723
rect 2263 717 2267 718
rect 2287 722 2291 723
rect 2287 717 2291 718
rect 2415 722 2419 723
rect 2415 717 2419 718
rect 2423 722 2427 723
rect 2423 717 2427 718
rect 2104 700 2106 717
rect 2264 700 2266 717
rect 2416 700 2418 717
rect 2102 699 2108 700
rect 2102 695 2103 699
rect 2107 695 2108 699
rect 2102 694 2108 695
rect 2262 699 2268 700
rect 2262 695 2263 699
rect 2267 695 2268 699
rect 2262 694 2268 695
rect 2414 699 2420 700
rect 2414 695 2415 699
rect 2419 695 2420 699
rect 2414 694 2420 695
rect 2488 692 2490 778
rect 2560 769 2562 785
rect 2630 783 2636 784
rect 2630 779 2631 783
rect 2635 779 2636 783
rect 2630 778 2636 779
rect 2558 768 2564 769
rect 2558 764 2559 768
rect 2563 764 2564 768
rect 2558 763 2564 764
rect 2632 760 2634 778
rect 2712 769 2714 785
rect 2782 783 2788 784
rect 2782 779 2783 783
rect 2787 779 2788 783
rect 2782 778 2788 779
rect 2710 768 2716 769
rect 2710 764 2711 768
rect 2715 764 2716 768
rect 2710 763 2716 764
rect 2784 760 2786 778
rect 2872 769 2874 785
rect 2942 783 2948 784
rect 2942 779 2943 783
rect 2947 779 2948 783
rect 2942 778 2948 779
rect 2870 768 2876 769
rect 2870 764 2871 768
rect 2875 764 2876 768
rect 2870 763 2876 764
rect 2944 760 2946 778
rect 3040 769 3042 785
rect 3110 783 3116 784
rect 3110 779 3111 783
rect 3115 779 3116 783
rect 3110 778 3116 779
rect 3038 768 3044 769
rect 3038 764 3039 768
rect 3043 764 3044 768
rect 3038 763 3044 764
rect 3112 760 3114 778
rect 3216 769 3218 785
rect 3368 769 3370 785
rect 3214 768 3220 769
rect 3214 764 3215 768
rect 3219 764 3220 768
rect 3214 763 3220 764
rect 3366 768 3372 769
rect 3366 764 3367 768
rect 3371 764 3372 768
rect 3366 763 3372 764
rect 3432 760 3434 794
rect 3464 791 3466 814
rect 3463 790 3467 791
rect 3463 785 3467 786
rect 3438 783 3444 784
rect 3438 779 3439 783
rect 3443 779 3444 783
rect 3438 778 3444 779
rect 2630 759 2636 760
rect 2630 755 2631 759
rect 2635 755 2636 759
rect 2630 754 2636 755
rect 2782 759 2788 760
rect 2782 755 2783 759
rect 2787 755 2788 759
rect 2782 754 2788 755
rect 2942 759 2948 760
rect 2942 755 2943 759
rect 2947 755 2948 759
rect 2942 754 2948 755
rect 3110 759 3116 760
rect 3110 755 3111 759
rect 3115 755 3116 759
rect 3110 754 3116 755
rect 3278 759 3284 760
rect 3278 755 3279 759
rect 3283 755 3284 759
rect 3278 754 3284 755
rect 3430 759 3436 760
rect 3430 755 3431 759
rect 3435 755 3436 759
rect 3430 754 3436 755
rect 2558 749 2564 750
rect 2558 745 2559 749
rect 2563 745 2564 749
rect 2558 744 2564 745
rect 2710 749 2716 750
rect 2710 745 2711 749
rect 2715 745 2716 749
rect 2710 744 2716 745
rect 2870 749 2876 750
rect 2870 745 2871 749
rect 2875 745 2876 749
rect 2870 744 2876 745
rect 3038 749 3044 750
rect 3038 745 3039 749
rect 3043 745 3044 749
rect 3038 744 3044 745
rect 3214 749 3220 750
rect 3214 745 3215 749
rect 3219 745 3220 749
rect 3214 744 3220 745
rect 2560 723 2562 744
rect 2712 723 2714 744
rect 2872 723 2874 744
rect 3040 723 3042 744
rect 3216 723 3218 744
rect 2559 722 2563 723
rect 2559 717 2563 718
rect 2567 722 2571 723
rect 2567 717 2571 718
rect 2711 722 2715 723
rect 2711 717 2715 718
rect 2719 722 2723 723
rect 2719 717 2723 718
rect 2871 722 2875 723
rect 2871 717 2875 718
rect 2879 722 2883 723
rect 2879 717 2883 718
rect 3039 722 3043 723
rect 3039 717 3043 718
rect 3199 722 3203 723
rect 3199 717 3203 718
rect 3215 722 3219 723
rect 3215 717 3219 718
rect 2568 700 2570 717
rect 2720 700 2722 717
rect 2880 700 2882 717
rect 3040 700 3042 717
rect 3200 700 3202 717
rect 2566 699 2572 700
rect 2566 695 2567 699
rect 2571 695 2572 699
rect 2566 694 2572 695
rect 2718 699 2724 700
rect 2718 695 2719 699
rect 2723 695 2724 699
rect 2718 694 2724 695
rect 2878 699 2884 700
rect 2878 695 2879 699
rect 2883 695 2884 699
rect 2878 694 2884 695
rect 3038 699 3044 700
rect 3038 695 3039 699
rect 3043 695 3044 699
rect 3038 694 3044 695
rect 3198 699 3204 700
rect 3198 695 3199 699
rect 3203 695 3204 699
rect 3198 694 3204 695
rect 2486 691 2492 692
rect 2174 687 2180 688
rect 2174 683 2175 687
rect 2179 683 2180 687
rect 2174 682 2180 683
rect 2334 687 2340 688
rect 2334 683 2335 687
rect 2339 683 2340 687
rect 2486 687 2487 691
rect 2491 687 2492 691
rect 2486 686 2492 687
rect 2646 691 2652 692
rect 2646 687 2647 691
rect 2651 687 2652 691
rect 2646 686 2652 687
rect 2798 691 2804 692
rect 2798 687 2799 691
rect 2803 687 2804 691
rect 3138 691 3144 692
rect 2798 686 2804 687
rect 3110 687 3116 688
rect 2334 682 2340 683
rect 2630 683 2636 684
rect 2102 680 2108 681
rect 2102 676 2103 680
rect 2107 676 2108 680
rect 2102 675 2108 676
rect 1962 663 1968 664
rect 1962 659 1963 663
rect 1967 659 1968 663
rect 2104 659 2106 675
rect 2176 664 2178 682
rect 2262 680 2268 681
rect 2262 676 2263 680
rect 2267 676 2268 680
rect 2262 675 2268 676
rect 2158 663 2164 664
rect 2158 659 2159 663
rect 2163 659 2164 663
rect 1807 658 1811 659
rect 1807 653 1811 654
rect 1831 658 1835 659
rect 1910 658 1916 659
rect 1951 658 1955 659
rect 1962 658 1968 659
rect 1975 658 1979 659
rect 1831 653 1835 654
rect 1951 653 1955 654
rect 1975 653 1979 654
rect 2103 658 2107 659
rect 2158 658 2164 659
rect 2174 663 2180 664
rect 2174 659 2175 663
rect 2179 659 2180 663
rect 2264 659 2266 675
rect 2336 664 2338 682
rect 2414 680 2420 681
rect 2414 676 2415 680
rect 2419 676 2420 680
rect 2414 675 2420 676
rect 2566 680 2572 681
rect 2566 676 2567 680
rect 2571 676 2572 680
rect 2630 679 2631 683
rect 2635 679 2636 683
rect 2630 678 2636 679
rect 2566 675 2572 676
rect 2334 663 2340 664
rect 2334 659 2335 663
rect 2339 659 2340 663
rect 2416 659 2418 675
rect 2568 659 2570 675
rect 2174 658 2180 659
rect 2239 658 2243 659
rect 2103 653 2107 654
rect 1767 638 1771 639
rect 1808 634 1810 653
rect 1966 651 1972 652
rect 1966 647 1967 651
rect 1971 647 1972 651
rect 1966 646 1972 647
rect 1767 633 1771 634
rect 1806 633 1812 634
rect 1742 631 1748 632
rect 1742 627 1743 631
rect 1747 627 1748 631
rect 1742 626 1748 627
rect 1670 616 1676 617
rect 1670 612 1671 616
rect 1675 612 1676 616
rect 1768 614 1770 633
rect 1806 629 1807 633
rect 1811 629 1812 633
rect 1806 628 1812 629
rect 1806 616 1812 617
rect 1670 611 1676 612
rect 1766 613 1772 614
rect 1766 609 1767 613
rect 1771 609 1772 613
rect 1806 612 1807 616
rect 1811 612 1812 616
rect 1806 611 1812 612
rect 1766 608 1772 609
rect 1126 607 1132 608
rect 1126 603 1127 607
rect 1131 603 1132 607
rect 1126 602 1132 603
rect 1278 607 1284 608
rect 1278 603 1279 607
rect 1283 603 1284 607
rect 1278 602 1284 603
rect 1286 607 1292 608
rect 1286 603 1287 607
rect 1291 603 1292 607
rect 1286 602 1292 603
rect 1446 607 1452 608
rect 1446 603 1447 607
rect 1451 603 1452 607
rect 1446 602 1452 603
rect 1606 607 1612 608
rect 1606 603 1607 607
rect 1611 603 1612 607
rect 1606 602 1612 603
rect 1206 597 1212 598
rect 1206 593 1207 597
rect 1211 593 1212 597
rect 1206 592 1212 593
rect 1366 597 1372 598
rect 1366 593 1367 597
rect 1371 593 1372 597
rect 1366 592 1372 593
rect 1208 571 1210 592
rect 1368 571 1370 592
rect 1135 570 1139 571
rect 1135 565 1139 566
rect 1207 570 1211 571
rect 1207 565 1211 566
rect 1319 570 1323 571
rect 1319 565 1323 566
rect 1367 570 1371 571
rect 1367 565 1371 566
rect 1136 548 1138 565
rect 1320 548 1322 565
rect 1134 547 1140 548
rect 1134 543 1135 547
rect 1139 543 1140 547
rect 1134 542 1140 543
rect 1318 547 1324 548
rect 1318 543 1319 547
rect 1323 543 1324 547
rect 1318 542 1324 543
rect 1110 539 1116 540
rect 1022 535 1028 536
rect 1022 531 1023 535
rect 1027 531 1028 535
rect 1110 535 1111 539
rect 1115 535 1116 539
rect 1110 534 1116 535
rect 1390 535 1396 536
rect 1022 530 1028 531
rect 1390 531 1391 535
rect 1395 531 1396 535
rect 1390 530 1396 531
rect 1024 512 1026 530
rect 1134 528 1140 529
rect 1134 524 1135 528
rect 1139 524 1140 528
rect 1134 523 1140 524
rect 1318 528 1324 529
rect 1318 524 1319 528
rect 1323 524 1324 528
rect 1318 523 1324 524
rect 982 511 988 512
rect 982 507 983 511
rect 987 507 988 511
rect 982 506 988 507
rect 1022 511 1028 512
rect 1022 507 1023 511
rect 1027 507 1028 511
rect 1022 506 1028 507
rect 1136 503 1138 523
rect 1320 503 1322 523
rect 1392 512 1394 530
rect 1448 520 1450 602
rect 1526 597 1532 598
rect 1526 593 1527 597
rect 1531 593 1532 597
rect 1526 592 1532 593
rect 1670 597 1676 598
rect 1670 593 1671 597
rect 1675 593 1676 597
rect 1670 592 1676 593
rect 1766 596 1772 597
rect 1766 592 1767 596
rect 1771 592 1772 596
rect 1528 571 1530 592
rect 1672 571 1674 592
rect 1766 591 1772 592
rect 1768 571 1770 591
rect 1808 587 1810 611
rect 1807 586 1811 587
rect 1807 581 1811 582
rect 1895 586 1899 587
rect 1895 581 1899 582
rect 1503 570 1507 571
rect 1503 565 1507 566
rect 1527 570 1531 571
rect 1527 565 1531 566
rect 1671 570 1675 571
rect 1671 565 1675 566
rect 1767 570 1771 571
rect 1767 565 1771 566
rect 1808 565 1810 581
rect 1504 548 1506 565
rect 1672 548 1674 565
rect 1768 549 1770 565
rect 1806 564 1812 565
rect 1896 564 1898 581
rect 1806 560 1807 564
rect 1811 560 1812 564
rect 1806 559 1812 560
rect 1894 563 1900 564
rect 1894 559 1895 563
rect 1899 559 1900 563
rect 1894 558 1900 559
rect 1968 556 1970 646
rect 1976 637 1978 653
rect 2046 651 2052 652
rect 2046 647 2047 651
rect 2051 647 2052 651
rect 2046 646 2052 647
rect 1974 636 1980 637
rect 1974 632 1975 636
rect 1979 632 1980 636
rect 1974 631 1980 632
rect 2048 628 2050 646
rect 2160 628 2162 658
rect 2239 653 2243 654
rect 2263 658 2267 659
rect 2334 658 2340 659
rect 2415 658 2419 659
rect 2263 653 2267 654
rect 2415 653 2419 654
rect 2479 658 2483 659
rect 2479 653 2483 654
rect 2567 658 2571 659
rect 2567 653 2571 654
rect 2240 637 2242 653
rect 2480 637 2482 653
rect 2550 651 2556 652
rect 2550 647 2551 651
rect 2555 647 2556 651
rect 2550 646 2556 647
rect 2238 636 2244 637
rect 2238 632 2239 636
rect 2243 632 2244 636
rect 2238 631 2244 632
rect 2478 636 2484 637
rect 2478 632 2479 636
rect 2483 632 2484 636
rect 2478 631 2484 632
rect 2552 628 2554 646
rect 2046 627 2052 628
rect 2046 623 2047 627
rect 2051 623 2052 627
rect 2046 622 2052 623
rect 2158 627 2164 628
rect 2158 623 2159 627
rect 2163 623 2164 627
rect 2158 622 2164 623
rect 2550 627 2556 628
rect 2550 623 2551 627
rect 2555 623 2556 627
rect 2550 622 2556 623
rect 1974 617 1980 618
rect 1974 613 1975 617
rect 1979 613 1980 617
rect 1974 612 1980 613
rect 2238 617 2244 618
rect 2238 613 2239 617
rect 2243 613 2244 617
rect 2238 612 2244 613
rect 2478 617 2484 618
rect 2478 613 2479 617
rect 2483 613 2484 617
rect 2478 612 2484 613
rect 1976 587 1978 612
rect 2240 587 2242 612
rect 2480 587 2482 612
rect 1975 586 1979 587
rect 1975 581 1979 582
rect 2015 586 2019 587
rect 2015 581 2019 582
rect 2143 586 2147 587
rect 2143 581 2147 582
rect 2239 586 2243 587
rect 2239 581 2243 582
rect 2279 586 2283 587
rect 2279 581 2283 582
rect 2423 586 2427 587
rect 2423 581 2427 582
rect 2479 586 2483 587
rect 2479 581 2483 582
rect 2567 586 2571 587
rect 2567 581 2571 582
rect 2016 564 2018 581
rect 2144 564 2146 581
rect 2280 564 2282 581
rect 2424 564 2426 581
rect 2568 564 2570 581
rect 2014 563 2020 564
rect 2014 559 2015 563
rect 2019 559 2020 563
rect 2014 558 2020 559
rect 2142 563 2148 564
rect 2142 559 2143 563
rect 2147 559 2148 563
rect 2142 558 2148 559
rect 2278 563 2284 564
rect 2278 559 2279 563
rect 2283 559 2284 563
rect 2278 558 2284 559
rect 2422 563 2428 564
rect 2422 559 2423 563
rect 2427 559 2428 563
rect 2422 558 2428 559
rect 2566 563 2572 564
rect 2566 559 2567 563
rect 2571 559 2572 563
rect 2566 558 2572 559
rect 1966 555 1972 556
rect 1966 551 1967 555
rect 1971 551 1972 555
rect 1966 550 1972 551
rect 1974 555 1980 556
rect 1974 551 1975 555
rect 1979 551 1980 555
rect 1974 550 1980 551
rect 2094 555 2100 556
rect 2094 551 2095 555
rect 2099 551 2100 555
rect 2094 550 2100 551
rect 2222 555 2228 556
rect 2222 551 2223 555
rect 2227 551 2228 555
rect 2222 550 2228 551
rect 2410 555 2416 556
rect 2410 551 2411 555
rect 2415 551 2416 555
rect 2410 550 2416 551
rect 1766 548 1772 549
rect 1502 547 1508 548
rect 1502 543 1503 547
rect 1507 543 1508 547
rect 1502 542 1508 543
rect 1670 547 1676 548
rect 1670 543 1671 547
rect 1675 543 1676 547
rect 1766 544 1767 548
rect 1771 544 1772 548
rect 1766 543 1772 544
rect 1806 547 1812 548
rect 1806 543 1807 547
rect 1811 543 1812 547
rect 1670 542 1676 543
rect 1806 542 1812 543
rect 1894 544 1900 545
rect 1574 535 1580 536
rect 1574 531 1575 535
rect 1579 531 1580 535
rect 1574 530 1580 531
rect 1742 535 1748 536
rect 1742 531 1743 535
rect 1747 531 1748 535
rect 1742 530 1748 531
rect 1766 531 1772 532
rect 1502 528 1508 529
rect 1502 524 1503 528
rect 1507 524 1508 528
rect 1502 523 1508 524
rect 1446 519 1452 520
rect 1446 515 1447 519
rect 1451 515 1452 519
rect 1446 514 1452 515
rect 1390 511 1396 512
rect 1390 507 1391 511
rect 1395 507 1396 511
rect 1390 506 1396 507
rect 1504 503 1506 523
rect 1576 512 1578 530
rect 1670 528 1676 529
rect 1670 524 1671 528
rect 1675 524 1676 528
rect 1670 523 1676 524
rect 1574 511 1580 512
rect 1574 507 1575 511
rect 1579 507 1580 511
rect 1574 506 1580 507
rect 1672 503 1674 523
rect 735 502 739 503
rect 735 497 739 498
rect 767 502 771 503
rect 767 497 771 498
rect 903 502 907 503
rect 903 497 907 498
rect 951 502 955 503
rect 951 497 955 498
rect 1063 502 1067 503
rect 1063 497 1067 498
rect 1135 502 1139 503
rect 1135 497 1139 498
rect 1223 502 1227 503
rect 1223 497 1227 498
rect 1319 502 1323 503
rect 1319 497 1323 498
rect 1375 502 1379 503
rect 1375 497 1379 498
rect 1503 502 1507 503
rect 1503 497 1507 498
rect 1527 502 1531 503
rect 1527 497 1531 498
rect 1671 502 1675 503
rect 1671 497 1675 498
rect 736 481 738 497
rect 814 495 820 496
rect 814 491 815 495
rect 819 491 820 495
rect 814 490 820 491
rect 734 480 740 481
rect 734 476 735 480
rect 739 476 740 480
rect 734 475 740 476
rect 816 472 818 490
rect 904 481 906 497
rect 998 495 1004 496
rect 998 491 999 495
rect 1003 491 1004 495
rect 998 490 1004 491
rect 902 480 908 481
rect 902 476 903 480
rect 907 476 908 480
rect 902 475 908 476
rect 318 471 324 472
rect 318 467 319 471
rect 323 467 324 471
rect 318 466 324 467
rect 470 471 476 472
rect 470 467 471 471
rect 475 467 476 471
rect 470 466 476 467
rect 634 471 640 472
rect 634 467 635 471
rect 639 467 640 471
rect 634 466 640 467
rect 814 471 820 472
rect 814 467 815 471
rect 819 467 820 471
rect 814 466 820 467
rect 246 461 252 462
rect 110 460 116 461
rect 110 456 111 460
rect 115 456 116 460
rect 246 457 247 461
rect 251 457 252 461
rect 246 456 252 457
rect 398 461 404 462
rect 398 457 399 461
rect 403 457 404 461
rect 398 456 404 457
rect 566 461 572 462
rect 566 457 567 461
rect 571 457 572 461
rect 566 456 572 457
rect 734 461 740 462
rect 734 457 735 461
rect 739 457 740 461
rect 734 456 740 457
rect 902 461 908 462
rect 902 457 903 461
rect 907 457 908 461
rect 902 456 908 457
rect 110 455 116 456
rect 112 435 114 455
rect 248 435 250 456
rect 400 435 402 456
rect 568 435 570 456
rect 736 435 738 456
rect 904 435 906 456
rect 111 434 115 435
rect 111 429 115 430
rect 247 434 251 435
rect 247 429 251 430
rect 399 434 403 435
rect 399 429 403 430
rect 519 434 523 435
rect 519 429 523 430
rect 567 434 571 435
rect 567 429 571 430
rect 615 434 619 435
rect 615 429 619 430
rect 719 434 723 435
rect 719 429 723 430
rect 735 434 739 435
rect 735 429 739 430
rect 823 434 827 435
rect 823 429 827 430
rect 903 434 907 435
rect 903 429 907 430
rect 927 434 931 435
rect 927 429 931 430
rect 112 413 114 429
rect 110 412 116 413
rect 520 412 522 429
rect 616 412 618 429
rect 720 412 722 429
rect 824 412 826 429
rect 928 412 930 429
rect 110 408 111 412
rect 115 408 116 412
rect 110 407 116 408
rect 518 411 524 412
rect 518 407 519 411
rect 523 407 524 411
rect 518 406 524 407
rect 614 411 620 412
rect 614 407 615 411
rect 619 407 620 411
rect 614 406 620 407
rect 718 411 724 412
rect 718 407 719 411
rect 723 407 724 411
rect 718 406 724 407
rect 822 411 828 412
rect 822 407 823 411
rect 827 407 828 411
rect 822 406 828 407
rect 926 411 932 412
rect 926 407 927 411
rect 931 407 932 411
rect 926 406 932 407
rect 1000 404 1002 490
rect 1064 481 1066 497
rect 1186 495 1192 496
rect 1186 491 1187 495
rect 1191 491 1192 495
rect 1186 490 1192 491
rect 1062 480 1068 481
rect 1062 476 1063 480
rect 1067 476 1068 480
rect 1062 475 1068 476
rect 1188 472 1190 490
rect 1224 481 1226 497
rect 1376 481 1378 497
rect 1528 481 1530 497
rect 1606 495 1612 496
rect 1606 491 1607 495
rect 1611 491 1612 495
rect 1606 490 1612 491
rect 1222 480 1228 481
rect 1222 476 1223 480
rect 1227 476 1228 480
rect 1222 475 1228 476
rect 1374 480 1380 481
rect 1374 476 1375 480
rect 1379 476 1380 480
rect 1374 475 1380 476
rect 1526 480 1532 481
rect 1526 476 1527 480
rect 1531 476 1532 480
rect 1526 475 1532 476
rect 1608 472 1610 490
rect 1672 481 1674 497
rect 1744 496 1746 530
rect 1766 527 1767 531
rect 1771 527 1772 531
rect 1766 526 1772 527
rect 1768 503 1770 526
rect 1808 519 1810 542
rect 1894 540 1895 544
rect 1899 540 1900 544
rect 1894 539 1900 540
rect 1896 519 1898 539
rect 1976 528 1978 550
rect 2014 544 2020 545
rect 2014 540 2015 544
rect 2019 540 2020 544
rect 2014 539 2020 540
rect 1974 527 1980 528
rect 1974 523 1975 527
rect 1979 523 1980 527
rect 1974 522 1980 523
rect 2016 519 2018 539
rect 2096 528 2098 550
rect 2142 544 2148 545
rect 2142 540 2143 544
rect 2147 540 2148 544
rect 2142 539 2148 540
rect 2094 527 2100 528
rect 2094 523 2095 527
rect 2099 523 2100 527
rect 2094 522 2100 523
rect 2144 519 2146 539
rect 2224 528 2226 550
rect 2278 544 2284 545
rect 2278 540 2279 544
rect 2283 540 2284 544
rect 2278 539 2284 540
rect 2222 527 2228 528
rect 2222 523 2223 527
rect 2227 523 2228 527
rect 2222 522 2228 523
rect 2206 519 2212 520
rect 2280 519 2282 539
rect 2412 528 2414 550
rect 2422 544 2428 545
rect 2422 540 2423 544
rect 2427 540 2428 544
rect 2422 539 2428 540
rect 2566 544 2572 545
rect 2566 540 2567 544
rect 2571 540 2572 544
rect 2566 539 2572 540
rect 2410 527 2416 528
rect 2410 523 2411 527
rect 2415 523 2416 527
rect 2410 522 2416 523
rect 2424 519 2426 539
rect 2430 527 2436 528
rect 2430 523 2431 527
rect 2435 523 2436 527
rect 2430 522 2436 523
rect 1807 518 1811 519
rect 1807 513 1811 514
rect 1895 518 1899 519
rect 1895 513 1899 514
rect 2015 518 2019 519
rect 2015 513 2019 514
rect 2135 518 2139 519
rect 2135 513 2139 514
rect 2143 518 2147 519
rect 2206 515 2207 519
rect 2211 515 2212 519
rect 2206 514 2212 515
rect 2239 518 2243 519
rect 2143 513 2147 514
rect 1767 502 1771 503
rect 1767 497 1771 498
rect 1742 495 1748 496
rect 1742 491 1743 495
rect 1747 491 1748 495
rect 1742 490 1748 491
rect 1670 480 1676 481
rect 1670 476 1671 480
rect 1675 476 1676 480
rect 1768 478 1770 497
rect 1808 494 1810 513
rect 2136 497 2138 513
rect 2134 496 2140 497
rect 1806 493 1812 494
rect 1806 489 1807 493
rect 1811 489 1812 493
rect 2134 492 2135 496
rect 2139 492 2140 496
rect 2134 491 2140 492
rect 1806 488 1812 489
rect 2208 488 2210 514
rect 2239 513 2243 514
rect 2279 518 2283 519
rect 2279 513 2283 514
rect 2359 518 2363 519
rect 2359 513 2363 514
rect 2423 518 2427 519
rect 2423 513 2427 514
rect 2240 497 2242 513
rect 2310 511 2316 512
rect 2310 507 2311 511
rect 2315 507 2316 511
rect 2310 506 2316 507
rect 2238 496 2244 497
rect 2238 492 2239 496
rect 2243 492 2244 496
rect 2238 491 2244 492
rect 2312 488 2314 506
rect 2360 497 2362 513
rect 2358 496 2364 497
rect 2358 492 2359 496
rect 2363 492 2364 496
rect 2358 491 2364 492
rect 2432 488 2434 522
rect 2568 519 2570 539
rect 2632 528 2634 678
rect 2648 664 2650 686
rect 2718 680 2724 681
rect 2718 676 2719 680
rect 2723 676 2724 680
rect 2718 675 2724 676
rect 2646 663 2652 664
rect 2646 659 2647 663
rect 2651 659 2652 663
rect 2720 659 2722 675
rect 2800 664 2802 686
rect 3110 683 3111 687
rect 3115 683 3116 687
rect 3138 687 3139 691
rect 3143 687 3144 691
rect 3138 686 3144 687
rect 3110 682 3116 683
rect 2878 680 2884 681
rect 2878 676 2879 680
rect 2883 676 2884 680
rect 2878 675 2884 676
rect 3038 680 3044 681
rect 3038 676 3039 680
rect 3043 676 3044 680
rect 3038 675 3044 676
rect 2798 663 2804 664
rect 2798 659 2799 663
rect 2803 659 2804 663
rect 2880 659 2882 675
rect 2950 663 2956 664
rect 2950 659 2951 663
rect 2955 659 2956 663
rect 3040 659 3042 675
rect 2646 658 2652 659
rect 2687 658 2691 659
rect 2687 653 2691 654
rect 2719 658 2723 659
rect 2798 658 2804 659
rect 2879 658 2883 659
rect 2950 658 2956 659
rect 3039 658 3043 659
rect 2719 653 2723 654
rect 2879 653 2883 654
rect 2688 637 2690 653
rect 2758 651 2764 652
rect 2758 647 2759 651
rect 2763 647 2764 651
rect 2758 646 2764 647
rect 2686 636 2692 637
rect 2686 632 2687 636
rect 2691 632 2692 636
rect 2686 631 2692 632
rect 2760 628 2762 646
rect 2838 643 2844 644
rect 2838 639 2839 643
rect 2843 639 2844 643
rect 2838 638 2844 639
rect 2758 627 2764 628
rect 2758 623 2759 627
rect 2763 623 2764 627
rect 2758 622 2764 623
rect 2686 617 2692 618
rect 2686 613 2687 617
rect 2691 613 2692 617
rect 2686 612 2692 613
rect 2688 587 2690 612
rect 2687 586 2691 587
rect 2687 581 2691 582
rect 2719 586 2723 587
rect 2719 581 2723 582
rect 2720 564 2722 581
rect 2718 563 2724 564
rect 2718 559 2719 563
rect 2723 559 2724 563
rect 2718 558 2724 559
rect 2840 556 2842 638
rect 2880 637 2882 653
rect 2878 636 2884 637
rect 2878 632 2879 636
rect 2883 632 2884 636
rect 2878 631 2884 632
rect 2952 628 2954 658
rect 3039 653 3043 654
rect 3055 658 3059 659
rect 3055 653 3059 654
rect 3056 637 3058 653
rect 3112 652 3114 682
rect 3140 672 3142 686
rect 3198 680 3204 681
rect 3198 676 3199 680
rect 3203 676 3204 680
rect 3198 675 3204 676
rect 3138 671 3144 672
rect 3138 667 3139 671
rect 3143 667 3144 671
rect 3138 666 3144 667
rect 3200 659 3202 675
rect 3280 664 3282 754
rect 3366 749 3372 750
rect 3366 745 3367 749
rect 3371 745 3372 749
rect 3366 744 3372 745
rect 3368 723 3370 744
rect 3367 722 3371 723
rect 3367 717 3371 718
rect 3278 663 3284 664
rect 3278 659 3279 663
rect 3283 659 3284 663
rect 3199 658 3203 659
rect 3199 653 3203 654
rect 3223 658 3227 659
rect 3278 658 3284 659
rect 3367 658 3371 659
rect 3223 653 3227 654
rect 3367 653 3371 654
rect 3110 651 3116 652
rect 3110 647 3111 651
rect 3115 647 3116 651
rect 3110 646 3116 647
rect 3126 651 3132 652
rect 3126 647 3127 651
rect 3131 647 3132 651
rect 3126 646 3132 647
rect 3054 636 3060 637
rect 3054 632 3055 636
rect 3059 632 3060 636
rect 3054 631 3060 632
rect 3128 628 3130 646
rect 3224 637 3226 653
rect 3368 637 3370 653
rect 3430 651 3436 652
rect 3430 647 3431 651
rect 3435 647 3436 651
rect 3430 646 3436 647
rect 3222 636 3228 637
rect 3222 632 3223 636
rect 3227 632 3228 636
rect 3222 631 3228 632
rect 3366 636 3372 637
rect 3366 632 3367 636
rect 3371 632 3372 636
rect 3366 631 3372 632
rect 2950 627 2956 628
rect 2950 623 2951 627
rect 2955 623 2956 627
rect 2950 622 2956 623
rect 3126 627 3132 628
rect 3126 623 3127 627
rect 3131 623 3132 627
rect 3126 622 3132 623
rect 3190 627 3196 628
rect 3190 623 3191 627
rect 3195 623 3196 627
rect 3190 622 3196 623
rect 2878 617 2884 618
rect 2878 613 2879 617
rect 2883 613 2884 617
rect 2878 612 2884 613
rect 3054 617 3060 618
rect 3054 613 3055 617
rect 3059 613 3060 617
rect 3054 612 3060 613
rect 2880 587 2882 612
rect 3056 587 3058 612
rect 2871 586 2875 587
rect 2871 581 2875 582
rect 2879 586 2883 587
rect 2879 581 2883 582
rect 3031 586 3035 587
rect 3031 581 3035 582
rect 3055 586 3059 587
rect 3055 581 3059 582
rect 2872 564 2874 581
rect 3032 564 3034 581
rect 2870 563 2876 564
rect 2870 559 2871 563
rect 2875 559 2876 563
rect 2870 558 2876 559
rect 3030 563 3036 564
rect 3030 559 3031 563
rect 3035 559 3036 563
rect 3030 558 3036 559
rect 2838 555 2844 556
rect 2638 551 2644 552
rect 2638 547 2639 551
rect 2643 547 2644 551
rect 2638 546 2644 547
rect 2790 551 2796 552
rect 2790 547 2791 551
rect 2795 547 2796 551
rect 2838 551 2839 555
rect 2843 551 2844 555
rect 3138 555 3144 556
rect 2838 550 2844 551
rect 3102 551 3108 552
rect 2790 546 2796 547
rect 3102 547 3103 551
rect 3107 547 3108 551
rect 3138 551 3139 555
rect 3143 551 3144 555
rect 3138 550 3144 551
rect 3102 546 3108 547
rect 2640 528 2642 546
rect 2718 544 2724 545
rect 2718 540 2719 544
rect 2723 540 2724 544
rect 2718 539 2724 540
rect 2630 527 2636 528
rect 2630 523 2631 527
rect 2635 523 2636 527
rect 2630 522 2636 523
rect 2638 527 2644 528
rect 2638 523 2639 527
rect 2643 523 2644 527
rect 2638 522 2644 523
rect 2720 519 2722 539
rect 2487 518 2491 519
rect 2487 513 2491 514
rect 2567 518 2571 519
rect 2567 513 2571 514
rect 2615 518 2619 519
rect 2615 513 2619 514
rect 2719 518 2723 519
rect 2719 513 2723 514
rect 2751 518 2755 519
rect 2751 513 2755 514
rect 2488 497 2490 513
rect 2616 497 2618 513
rect 2670 511 2676 512
rect 2670 507 2671 511
rect 2675 507 2676 511
rect 2670 506 2676 507
rect 2486 496 2492 497
rect 2486 492 2487 496
rect 2491 492 2492 496
rect 2486 491 2492 492
rect 2614 496 2620 497
rect 2614 492 2615 496
rect 2619 492 2620 496
rect 2614 491 2620 492
rect 2206 487 2212 488
rect 2206 483 2207 487
rect 2211 483 2212 487
rect 2206 482 2212 483
rect 2310 487 2316 488
rect 2310 483 2311 487
rect 2315 483 2316 487
rect 2310 482 2316 483
rect 2430 487 2436 488
rect 2430 483 2431 487
rect 2435 483 2436 487
rect 2430 482 2436 483
rect 1670 475 1676 476
rect 1766 477 1772 478
rect 2134 477 2140 478
rect 1766 473 1767 477
rect 1771 473 1772 477
rect 1766 472 1772 473
rect 1806 476 1812 477
rect 1806 472 1807 476
rect 1811 472 1812 476
rect 2134 473 2135 477
rect 2139 473 2140 477
rect 2134 472 2140 473
rect 2238 477 2244 478
rect 2238 473 2239 477
rect 2243 473 2244 477
rect 2238 472 2244 473
rect 2358 477 2364 478
rect 2358 473 2359 477
rect 2363 473 2364 477
rect 2358 472 2364 473
rect 2486 477 2492 478
rect 2486 473 2487 477
rect 2491 473 2492 477
rect 2486 472 2492 473
rect 2614 477 2620 478
rect 2614 473 2615 477
rect 2619 473 2620 477
rect 2614 472 2620 473
rect 1186 471 1192 472
rect 1186 467 1187 471
rect 1191 467 1192 471
rect 1186 466 1192 467
rect 1294 471 1300 472
rect 1294 467 1295 471
rect 1299 467 1300 471
rect 1294 466 1300 467
rect 1606 471 1612 472
rect 1806 471 1812 472
rect 1606 467 1607 471
rect 1611 467 1612 471
rect 1606 466 1612 467
rect 1062 461 1068 462
rect 1062 457 1063 461
rect 1067 457 1068 461
rect 1062 456 1068 457
rect 1222 461 1228 462
rect 1222 457 1223 461
rect 1227 457 1228 461
rect 1222 456 1228 457
rect 1064 435 1066 456
rect 1224 435 1226 456
rect 1023 434 1027 435
rect 1023 429 1027 430
rect 1063 434 1067 435
rect 1063 429 1067 430
rect 1127 434 1131 435
rect 1127 429 1131 430
rect 1223 434 1227 435
rect 1223 429 1227 430
rect 1231 434 1235 435
rect 1231 429 1235 430
rect 1024 412 1026 429
rect 1128 412 1130 429
rect 1232 412 1234 429
rect 1022 411 1028 412
rect 1022 407 1023 411
rect 1027 407 1028 411
rect 1022 406 1028 407
rect 1126 411 1132 412
rect 1126 407 1127 411
rect 1131 407 1132 411
rect 1126 406 1132 407
rect 1230 411 1236 412
rect 1230 407 1231 411
rect 1235 407 1236 411
rect 1230 406 1236 407
rect 798 403 804 404
rect 590 399 596 400
rect 110 395 116 396
rect 110 391 111 395
rect 115 391 116 395
rect 590 395 591 399
rect 595 395 596 399
rect 590 394 596 395
rect 686 399 692 400
rect 686 395 687 399
rect 691 395 692 399
rect 798 399 799 403
rect 803 399 804 403
rect 798 398 804 399
rect 998 403 1004 404
rect 998 399 999 403
rect 1003 399 1004 403
rect 1206 403 1212 404
rect 998 398 1004 399
rect 1094 399 1100 400
rect 686 394 692 395
rect 110 390 116 391
rect 518 392 524 393
rect 112 367 114 390
rect 518 388 519 392
rect 523 388 524 392
rect 518 387 524 388
rect 520 367 522 387
rect 592 376 594 394
rect 614 392 620 393
rect 614 388 615 392
rect 619 388 620 392
rect 614 387 620 388
rect 590 375 596 376
rect 590 371 591 375
rect 595 371 596 375
rect 590 370 596 371
rect 616 367 618 387
rect 688 376 690 394
rect 718 392 724 393
rect 718 388 719 392
rect 723 388 724 392
rect 718 387 724 388
rect 686 375 692 376
rect 686 371 687 375
rect 691 371 692 375
rect 686 370 692 371
rect 720 367 722 387
rect 800 384 802 398
rect 1094 395 1095 399
rect 1099 395 1100 399
rect 1094 394 1100 395
rect 1198 399 1204 400
rect 1198 395 1199 399
rect 1203 395 1204 399
rect 1206 399 1207 403
rect 1211 399 1212 403
rect 1206 398 1212 399
rect 1198 394 1204 395
rect 822 392 828 393
rect 822 388 823 392
rect 827 388 828 392
rect 822 387 828 388
rect 926 392 932 393
rect 926 388 927 392
rect 931 388 932 392
rect 926 387 932 388
rect 1022 392 1028 393
rect 1022 388 1023 392
rect 1027 388 1028 392
rect 1022 387 1028 388
rect 798 383 804 384
rect 798 379 799 383
rect 803 379 804 383
rect 798 378 804 379
rect 824 367 826 387
rect 886 375 892 376
rect 886 371 887 375
rect 891 371 892 375
rect 886 370 892 371
rect 111 366 115 367
rect 111 361 115 362
rect 471 366 475 367
rect 471 361 475 362
rect 519 366 523 367
rect 519 361 523 362
rect 559 366 563 367
rect 559 361 563 362
rect 615 366 619 367
rect 615 361 619 362
rect 647 366 651 367
rect 647 361 651 362
rect 719 366 723 367
rect 719 361 723 362
rect 735 366 739 367
rect 735 361 739 362
rect 823 366 827 367
rect 823 361 827 362
rect 112 342 114 361
rect 472 345 474 361
rect 542 359 548 360
rect 542 355 543 359
rect 547 355 548 359
rect 542 354 548 355
rect 470 344 476 345
rect 110 341 116 342
rect 110 337 111 341
rect 115 337 116 341
rect 470 340 471 344
rect 475 340 476 344
rect 470 339 476 340
rect 110 336 116 337
rect 544 336 546 354
rect 560 345 562 361
rect 630 359 636 360
rect 630 355 631 359
rect 635 355 636 359
rect 630 354 636 355
rect 558 344 564 345
rect 558 340 559 344
rect 563 340 564 344
rect 558 339 564 340
rect 632 336 634 354
rect 638 351 644 352
rect 638 347 639 351
rect 643 347 644 351
rect 638 346 644 347
rect 542 335 548 336
rect 542 331 543 335
rect 547 331 548 335
rect 542 330 548 331
rect 630 335 636 336
rect 630 331 631 335
rect 635 331 636 335
rect 630 330 636 331
rect 470 325 476 326
rect 110 324 116 325
rect 110 320 111 324
rect 115 320 116 324
rect 470 321 471 325
rect 475 321 476 325
rect 470 320 476 321
rect 558 325 564 326
rect 558 321 559 325
rect 563 321 564 325
rect 558 320 564 321
rect 110 319 116 320
rect 112 299 114 319
rect 472 299 474 320
rect 560 299 562 320
rect 111 298 115 299
rect 111 293 115 294
rect 279 298 283 299
rect 279 293 283 294
rect 367 298 371 299
rect 367 293 371 294
rect 463 298 467 299
rect 463 293 467 294
rect 471 298 475 299
rect 471 293 475 294
rect 559 298 563 299
rect 559 293 563 294
rect 112 277 114 293
rect 110 276 116 277
rect 280 276 282 293
rect 368 276 370 293
rect 464 276 466 293
rect 560 276 562 293
rect 110 272 111 276
rect 115 272 116 276
rect 110 271 116 272
rect 278 275 284 276
rect 278 271 279 275
rect 283 271 284 275
rect 278 270 284 271
rect 366 275 372 276
rect 366 271 367 275
rect 371 271 372 275
rect 366 270 372 271
rect 462 275 468 276
rect 462 271 463 275
rect 467 271 468 275
rect 462 270 468 271
rect 558 275 564 276
rect 558 271 559 275
rect 563 271 564 275
rect 558 270 564 271
rect 640 268 642 346
rect 648 345 650 361
rect 736 345 738 361
rect 806 359 812 360
rect 806 355 807 359
rect 811 355 812 359
rect 806 354 812 355
rect 646 344 652 345
rect 646 340 647 344
rect 651 340 652 344
rect 646 339 652 340
rect 734 344 740 345
rect 734 340 735 344
rect 739 340 740 344
rect 734 339 740 340
rect 808 336 810 354
rect 824 345 826 361
rect 822 344 828 345
rect 822 340 823 344
rect 827 340 828 344
rect 822 339 828 340
rect 888 336 890 370
rect 928 367 930 387
rect 1024 367 1026 387
rect 1096 376 1098 394
rect 1126 392 1132 393
rect 1126 388 1127 392
rect 1131 388 1132 392
rect 1126 387 1132 388
rect 1094 375 1100 376
rect 1094 371 1095 375
rect 1099 371 1100 375
rect 1094 370 1100 371
rect 1128 367 1130 387
rect 911 366 915 367
rect 911 361 915 362
rect 927 366 931 367
rect 927 361 931 362
rect 999 366 1003 367
rect 999 361 1003 362
rect 1023 366 1027 367
rect 1023 361 1027 362
rect 1087 366 1091 367
rect 1087 361 1091 362
rect 1127 366 1131 367
rect 1127 361 1131 362
rect 1175 366 1179 367
rect 1175 361 1179 362
rect 912 345 914 361
rect 990 359 996 360
rect 990 355 991 359
rect 995 355 996 359
rect 990 354 996 355
rect 910 344 916 345
rect 910 340 911 344
rect 915 340 916 344
rect 910 339 916 340
rect 992 336 994 354
rect 1000 345 1002 361
rect 1078 359 1084 360
rect 1078 355 1079 359
rect 1083 355 1084 359
rect 1078 354 1084 355
rect 998 344 1004 345
rect 998 340 999 344
rect 1003 340 1004 344
rect 998 339 1004 340
rect 1080 336 1082 354
rect 1088 345 1090 361
rect 1176 345 1178 361
rect 1200 360 1202 394
rect 1208 384 1210 398
rect 1230 392 1236 393
rect 1230 388 1231 392
rect 1235 388 1236 392
rect 1230 387 1236 388
rect 1206 383 1212 384
rect 1206 379 1207 383
rect 1211 379 1212 383
rect 1206 378 1212 379
rect 1232 367 1234 387
rect 1296 376 1298 466
rect 1374 461 1380 462
rect 1374 457 1375 461
rect 1379 457 1380 461
rect 1374 456 1380 457
rect 1526 461 1532 462
rect 1526 457 1527 461
rect 1531 457 1532 461
rect 1526 456 1532 457
rect 1670 461 1676 462
rect 1670 457 1671 461
rect 1675 457 1676 461
rect 1670 456 1676 457
rect 1766 460 1772 461
rect 1766 456 1767 460
rect 1771 456 1772 460
rect 1376 435 1378 456
rect 1528 435 1530 456
rect 1672 435 1674 456
rect 1766 455 1772 456
rect 1768 435 1770 455
rect 1808 447 1810 471
rect 2136 447 2138 472
rect 2240 447 2242 472
rect 2360 447 2362 472
rect 2488 447 2490 472
rect 2616 447 2618 472
rect 1807 446 1811 447
rect 1807 441 1811 442
rect 2135 446 2139 447
rect 2135 441 2139 442
rect 2239 446 2243 447
rect 2239 441 2243 442
rect 2335 446 2339 447
rect 2335 441 2339 442
rect 2359 446 2363 447
rect 2359 441 2363 442
rect 2447 446 2451 447
rect 2447 441 2451 442
rect 2487 446 2491 447
rect 2487 441 2491 442
rect 2559 446 2563 447
rect 2559 441 2563 442
rect 2615 446 2619 447
rect 2615 441 2619 442
rect 1335 434 1339 435
rect 1335 429 1339 430
rect 1375 434 1379 435
rect 1375 429 1379 430
rect 1439 434 1443 435
rect 1439 429 1443 430
rect 1527 434 1531 435
rect 1527 429 1531 430
rect 1671 434 1675 435
rect 1671 429 1675 430
rect 1767 434 1771 435
rect 1767 429 1771 430
rect 1336 412 1338 429
rect 1440 412 1442 429
rect 1768 413 1770 429
rect 1808 425 1810 441
rect 1806 424 1812 425
rect 2240 424 2242 441
rect 2336 424 2338 441
rect 2448 424 2450 441
rect 2560 424 2562 441
rect 1806 420 1807 424
rect 1811 420 1812 424
rect 1806 419 1812 420
rect 2238 423 2244 424
rect 2238 419 2239 423
rect 2243 419 2244 423
rect 2238 418 2244 419
rect 2334 423 2340 424
rect 2334 419 2335 423
rect 2339 419 2340 423
rect 2334 418 2340 419
rect 2446 423 2452 424
rect 2446 419 2447 423
rect 2451 419 2452 423
rect 2446 418 2452 419
rect 2558 423 2564 424
rect 2558 419 2559 423
rect 2563 419 2564 423
rect 2558 418 2564 419
rect 2672 416 2674 506
rect 2752 497 2754 513
rect 2792 512 2794 546
rect 2870 544 2876 545
rect 2870 540 2871 544
rect 2875 540 2876 544
rect 2870 539 2876 540
rect 3030 544 3036 545
rect 3030 540 3031 544
rect 3035 540 3036 544
rect 3030 539 3036 540
rect 2872 519 2874 539
rect 3032 519 3034 539
rect 3104 528 3106 546
rect 3140 536 3142 550
rect 3138 535 3144 536
rect 3138 531 3139 535
rect 3143 531 3144 535
rect 3138 530 3144 531
rect 3078 527 3084 528
rect 3078 523 3079 527
rect 3083 523 3084 527
rect 3078 522 3084 523
rect 3102 527 3108 528
rect 3102 523 3103 527
rect 3107 523 3108 527
rect 3102 522 3108 523
rect 2871 518 2875 519
rect 2871 513 2875 514
rect 2879 518 2883 519
rect 2879 513 2883 514
rect 3007 518 3011 519
rect 3007 513 3011 514
rect 3031 518 3035 519
rect 3031 513 3035 514
rect 2790 511 2796 512
rect 2790 507 2791 511
rect 2795 507 2796 511
rect 2790 506 2796 507
rect 2880 497 2882 513
rect 2950 511 2956 512
rect 2950 507 2951 511
rect 2955 507 2956 511
rect 2950 506 2956 507
rect 2750 496 2756 497
rect 2750 492 2751 496
rect 2755 492 2756 496
rect 2750 491 2756 492
rect 2878 496 2884 497
rect 2878 492 2879 496
rect 2883 492 2884 496
rect 2878 491 2884 492
rect 2952 488 2954 506
rect 3008 497 3010 513
rect 3006 496 3012 497
rect 3006 492 3007 496
rect 3011 492 3012 496
rect 3006 491 3012 492
rect 3080 488 3082 522
rect 3135 518 3139 519
rect 3135 513 3139 514
rect 3102 503 3108 504
rect 3102 499 3103 503
rect 3107 499 3108 503
rect 3102 498 3108 499
rect 2822 487 2828 488
rect 2822 483 2823 487
rect 2827 483 2828 487
rect 2822 482 2828 483
rect 2950 487 2956 488
rect 2950 483 2951 487
rect 2955 483 2956 487
rect 2950 482 2956 483
rect 3078 487 3084 488
rect 3078 483 3079 487
rect 3083 483 3084 487
rect 3078 482 3084 483
rect 2750 477 2756 478
rect 2750 473 2751 477
rect 2755 473 2756 477
rect 2750 472 2756 473
rect 2752 447 2754 472
rect 2679 446 2683 447
rect 2679 441 2683 442
rect 2751 446 2755 447
rect 2751 441 2755 442
rect 2799 446 2803 447
rect 2799 441 2803 442
rect 2680 424 2682 441
rect 2800 424 2802 441
rect 2678 423 2684 424
rect 2678 419 2679 423
rect 2683 419 2684 423
rect 2678 418 2684 419
rect 2798 423 2804 424
rect 2798 419 2799 423
rect 2803 419 2804 423
rect 2798 418 2804 419
rect 2670 415 2676 416
rect 1766 412 1772 413
rect 1334 411 1340 412
rect 1334 407 1335 411
rect 1339 407 1340 411
rect 1334 406 1340 407
rect 1438 411 1444 412
rect 1438 407 1439 411
rect 1443 407 1444 411
rect 1766 408 1767 412
rect 1771 408 1772 412
rect 2406 411 2412 412
rect 1766 407 1772 408
rect 1806 407 1812 408
rect 1438 406 1444 407
rect 1414 403 1420 404
rect 1406 399 1412 400
rect 1406 395 1407 399
rect 1411 395 1412 399
rect 1414 399 1415 403
rect 1419 399 1420 403
rect 1806 403 1807 407
rect 1811 403 1812 407
rect 2406 407 2407 411
rect 2411 407 2412 411
rect 2406 406 2412 407
rect 2518 411 2524 412
rect 2518 407 2519 411
rect 2523 407 2524 411
rect 2518 406 2524 407
rect 2630 411 2636 412
rect 2630 407 2631 411
rect 2635 407 2636 411
rect 2670 411 2671 415
rect 2675 411 2676 415
rect 2670 410 2676 411
rect 2630 406 2636 407
rect 1806 402 1812 403
rect 2238 404 2244 405
rect 1414 398 1420 399
rect 1406 394 1412 395
rect 1334 392 1340 393
rect 1334 388 1335 392
rect 1339 388 1340 392
rect 1334 387 1340 388
rect 1294 375 1300 376
rect 1294 371 1295 375
rect 1299 371 1300 375
rect 1294 370 1300 371
rect 1336 367 1338 387
rect 1408 376 1410 394
rect 1416 384 1418 398
rect 1766 395 1772 396
rect 1438 392 1444 393
rect 1438 388 1439 392
rect 1443 388 1444 392
rect 1766 391 1767 395
rect 1771 391 1772 395
rect 1766 390 1772 391
rect 1438 387 1444 388
rect 1414 383 1420 384
rect 1414 379 1415 383
rect 1419 379 1420 383
rect 1414 378 1420 379
rect 1406 375 1412 376
rect 1406 371 1407 375
rect 1411 371 1412 375
rect 1406 370 1412 371
rect 1440 367 1442 387
rect 1768 367 1770 390
rect 1808 379 1810 402
rect 2238 400 2239 404
rect 2243 400 2244 404
rect 2238 399 2244 400
rect 2334 404 2340 405
rect 2334 400 2335 404
rect 2339 400 2340 404
rect 2334 399 2340 400
rect 2240 379 2242 399
rect 2336 379 2338 399
rect 2408 388 2410 406
rect 2446 404 2452 405
rect 2446 400 2447 404
rect 2451 400 2452 404
rect 2446 399 2452 400
rect 2406 387 2412 388
rect 2406 383 2407 387
rect 2411 383 2412 387
rect 2406 382 2412 383
rect 2438 379 2444 380
rect 2448 379 2450 399
rect 2520 388 2522 406
rect 2558 404 2564 405
rect 2558 400 2559 404
rect 2563 400 2564 404
rect 2558 399 2564 400
rect 2518 387 2524 388
rect 2518 383 2519 387
rect 2523 383 2524 387
rect 2518 382 2524 383
rect 2560 379 2562 399
rect 2632 388 2634 406
rect 2678 404 2684 405
rect 2678 400 2679 404
rect 2683 400 2684 404
rect 2678 399 2684 400
rect 2798 404 2804 405
rect 2798 400 2799 404
rect 2803 400 2804 404
rect 2798 399 2804 400
rect 2630 387 2636 388
rect 2630 383 2631 387
rect 2635 383 2636 387
rect 2630 382 2636 383
rect 2680 379 2682 399
rect 2800 379 2802 399
rect 2824 388 2826 482
rect 2878 477 2884 478
rect 2878 473 2879 477
rect 2883 473 2884 477
rect 2878 472 2884 473
rect 3006 477 3012 478
rect 3006 473 3007 477
rect 3011 473 3012 477
rect 3006 472 3012 473
rect 2880 447 2882 472
rect 3008 447 3010 472
rect 2879 446 2883 447
rect 2879 441 2883 442
rect 2911 446 2915 447
rect 2911 441 2915 442
rect 3007 446 3011 447
rect 3007 441 3011 442
rect 3023 446 3027 447
rect 3023 441 3027 442
rect 2912 424 2914 441
rect 3024 424 3026 441
rect 2910 423 2916 424
rect 2910 419 2911 423
rect 2915 419 2916 423
rect 2910 418 2916 419
rect 3022 423 3028 424
rect 3022 419 3023 423
rect 3027 419 3028 423
rect 3022 418 3028 419
rect 3104 416 3106 498
rect 3136 497 3138 513
rect 3192 512 3194 622
rect 3222 617 3228 618
rect 3222 613 3223 617
rect 3227 613 3228 617
rect 3222 612 3228 613
rect 3366 617 3372 618
rect 3366 613 3367 617
rect 3371 613 3372 617
rect 3366 612 3372 613
rect 3224 587 3226 612
rect 3368 587 3370 612
rect 3199 586 3203 587
rect 3199 581 3203 582
rect 3223 586 3227 587
rect 3223 581 3227 582
rect 3367 586 3371 587
rect 3367 581 3371 582
rect 3200 564 3202 581
rect 3368 564 3370 581
rect 3198 563 3204 564
rect 3198 559 3199 563
rect 3203 559 3204 563
rect 3198 558 3204 559
rect 3366 563 3372 564
rect 3366 559 3367 563
rect 3371 559 3372 563
rect 3432 560 3434 646
rect 3440 628 3442 778
rect 3464 766 3466 785
rect 3462 765 3468 766
rect 3462 761 3463 765
rect 3467 761 3468 765
rect 3462 760 3468 761
rect 3462 748 3468 749
rect 3462 744 3463 748
rect 3467 744 3468 748
rect 3462 743 3468 744
rect 3464 723 3466 743
rect 3463 722 3467 723
rect 3463 717 3467 718
rect 3464 701 3466 717
rect 3462 700 3468 701
rect 3462 696 3463 700
rect 3467 696 3468 700
rect 3462 695 3468 696
rect 3462 683 3468 684
rect 3462 679 3463 683
rect 3467 679 3468 683
rect 3462 678 3468 679
rect 3464 659 3466 678
rect 3463 658 3467 659
rect 3463 653 3467 654
rect 3464 634 3466 653
rect 3462 633 3468 634
rect 3462 629 3463 633
rect 3467 629 3468 633
rect 3462 628 3468 629
rect 3438 627 3444 628
rect 3438 623 3439 627
rect 3443 623 3444 627
rect 3438 622 3444 623
rect 3462 616 3468 617
rect 3462 612 3463 616
rect 3467 612 3468 616
rect 3462 611 3468 612
rect 3464 587 3466 611
rect 3463 586 3467 587
rect 3463 581 3467 582
rect 3464 565 3466 581
rect 3462 564 3468 565
rect 3462 560 3463 564
rect 3467 560 3468 564
rect 3366 558 3372 559
rect 3430 559 3436 560
rect 3462 559 3468 560
rect 3430 555 3431 559
rect 3435 555 3436 559
rect 3430 554 3436 555
rect 3462 547 3468 548
rect 3198 544 3204 545
rect 3198 540 3199 544
rect 3203 540 3204 544
rect 3198 539 3204 540
rect 3366 544 3372 545
rect 3366 540 3367 544
rect 3371 540 3372 544
rect 3462 543 3463 547
rect 3467 543 3468 547
rect 3462 542 3468 543
rect 3366 539 3372 540
rect 3200 519 3202 539
rect 3368 519 3370 539
rect 3430 527 3436 528
rect 3430 523 3431 527
rect 3435 523 3436 527
rect 3430 522 3436 523
rect 3199 518 3203 519
rect 3199 513 3203 514
rect 3263 518 3267 519
rect 3263 513 3267 514
rect 3367 518 3371 519
rect 3367 513 3371 514
rect 3190 511 3196 512
rect 3190 507 3191 511
rect 3195 507 3196 511
rect 3190 506 3196 507
rect 3206 511 3212 512
rect 3206 507 3207 511
rect 3211 507 3212 511
rect 3206 506 3212 507
rect 3134 496 3140 497
rect 3134 492 3135 496
rect 3139 492 3140 496
rect 3134 491 3140 492
rect 3208 488 3210 506
rect 3264 497 3266 513
rect 3368 497 3370 513
rect 3262 496 3268 497
rect 3262 492 3263 496
rect 3267 492 3268 496
rect 3262 491 3268 492
rect 3366 496 3372 497
rect 3366 492 3367 496
rect 3371 492 3372 496
rect 3366 491 3372 492
rect 3432 488 3434 522
rect 3464 519 3466 542
rect 3463 518 3467 519
rect 3463 513 3467 514
rect 3438 511 3444 512
rect 3438 507 3439 511
rect 3443 507 3444 511
rect 3438 506 3444 507
rect 3206 487 3212 488
rect 3206 483 3207 487
rect 3211 483 3212 487
rect 3206 482 3212 483
rect 3326 487 3332 488
rect 3326 483 3327 487
rect 3331 483 3332 487
rect 3326 482 3332 483
rect 3430 487 3436 488
rect 3430 483 3431 487
rect 3435 483 3436 487
rect 3430 482 3436 483
rect 3134 477 3140 478
rect 3134 473 3135 477
rect 3139 473 3140 477
rect 3134 472 3140 473
rect 3262 477 3268 478
rect 3262 473 3263 477
rect 3267 473 3268 477
rect 3262 472 3268 473
rect 3136 447 3138 472
rect 3264 447 3266 472
rect 3135 446 3139 447
rect 3135 441 3139 442
rect 3143 446 3147 447
rect 3143 441 3147 442
rect 3263 446 3267 447
rect 3263 441 3267 442
rect 3144 424 3146 441
rect 3264 424 3266 441
rect 3142 423 3148 424
rect 3142 419 3143 423
rect 3147 419 3148 423
rect 3142 418 3148 419
rect 3262 423 3268 424
rect 3262 419 3263 423
rect 3267 419 3268 423
rect 3262 418 3268 419
rect 3102 415 3108 416
rect 2870 411 2876 412
rect 2870 407 2871 411
rect 2875 407 2876 411
rect 2870 406 2876 407
rect 2982 411 2988 412
rect 2982 407 2983 411
rect 2987 407 2988 411
rect 2982 406 2988 407
rect 3094 411 3100 412
rect 3094 407 3095 411
rect 3099 407 3100 411
rect 3102 411 3103 415
rect 3107 411 3108 415
rect 3102 410 3108 411
rect 3094 406 3100 407
rect 2822 387 2828 388
rect 2822 383 2823 387
rect 2827 383 2828 387
rect 2822 382 2828 383
rect 1807 378 1811 379
rect 1807 373 1811 374
rect 2063 378 2067 379
rect 2063 373 2067 374
rect 2151 378 2155 379
rect 2151 373 2155 374
rect 2239 378 2243 379
rect 2239 373 2243 374
rect 2247 378 2251 379
rect 2247 373 2251 374
rect 2335 378 2339 379
rect 2335 373 2339 374
rect 2359 378 2363 379
rect 2438 375 2439 379
rect 2443 375 2444 379
rect 2438 374 2444 375
rect 2447 378 2451 379
rect 2359 373 2363 374
rect 1231 366 1235 367
rect 1231 361 1235 362
rect 1263 366 1267 367
rect 1263 361 1267 362
rect 1335 366 1339 367
rect 1335 361 1339 362
rect 1439 366 1443 367
rect 1439 361 1443 362
rect 1767 366 1771 367
rect 1767 361 1771 362
rect 1198 359 1204 360
rect 1198 355 1199 359
rect 1203 355 1204 359
rect 1198 354 1204 355
rect 1246 359 1252 360
rect 1246 355 1247 359
rect 1251 355 1252 359
rect 1246 354 1252 355
rect 1086 344 1092 345
rect 1086 340 1087 344
rect 1091 340 1092 344
rect 1086 339 1092 340
rect 1174 344 1180 345
rect 1174 340 1175 344
rect 1179 340 1180 344
rect 1174 339 1180 340
rect 1248 336 1250 354
rect 1264 345 1266 361
rect 1262 344 1268 345
rect 1262 340 1263 344
rect 1267 340 1268 344
rect 1768 342 1770 361
rect 1808 354 1810 373
rect 2064 357 2066 373
rect 2134 371 2140 372
rect 2134 367 2135 371
rect 2139 367 2140 371
rect 2134 366 2140 367
rect 2062 356 2068 357
rect 1806 353 1812 354
rect 1806 349 1807 353
rect 1811 349 1812 353
rect 2062 352 2063 356
rect 2067 352 2068 356
rect 2062 351 2068 352
rect 1806 348 1812 349
rect 2136 348 2138 366
rect 2152 357 2154 373
rect 2222 371 2228 372
rect 2222 367 2223 371
rect 2227 367 2228 371
rect 2222 366 2228 367
rect 2150 356 2156 357
rect 2150 352 2151 356
rect 2155 352 2156 356
rect 2150 351 2156 352
rect 2224 348 2226 366
rect 2248 357 2250 373
rect 2318 371 2324 372
rect 2318 367 2319 371
rect 2323 367 2324 371
rect 2318 366 2324 367
rect 2246 356 2252 357
rect 2246 352 2247 356
rect 2251 352 2252 356
rect 2246 351 2252 352
rect 2320 348 2322 366
rect 2360 357 2362 373
rect 2430 371 2436 372
rect 2430 367 2431 371
rect 2435 367 2436 371
rect 2430 366 2436 367
rect 2422 363 2428 364
rect 2422 359 2423 363
rect 2427 359 2428 363
rect 2422 358 2428 359
rect 2358 356 2364 357
rect 2358 352 2359 356
rect 2363 352 2364 356
rect 2358 351 2364 352
rect 2134 347 2140 348
rect 2134 343 2135 347
rect 2139 343 2140 347
rect 2134 342 2140 343
rect 2222 347 2228 348
rect 2222 343 2223 347
rect 2227 343 2228 347
rect 2222 342 2228 343
rect 2318 347 2324 348
rect 2318 343 2319 347
rect 2323 343 2324 347
rect 2318 342 2324 343
rect 1262 339 1268 340
rect 1766 341 1772 342
rect 1766 337 1767 341
rect 1771 337 1772 341
rect 2062 337 2068 338
rect 1766 336 1772 337
rect 1806 336 1812 337
rect 806 335 812 336
rect 806 331 807 335
rect 811 331 812 335
rect 806 330 812 331
rect 886 335 892 336
rect 886 331 887 335
rect 891 331 892 335
rect 886 330 892 331
rect 902 335 908 336
rect 902 331 903 335
rect 907 331 908 335
rect 902 330 908 331
rect 990 335 996 336
rect 990 331 991 335
rect 995 331 996 335
rect 990 330 996 331
rect 1078 335 1084 336
rect 1078 331 1079 335
rect 1083 331 1084 335
rect 1078 330 1084 331
rect 1246 335 1252 336
rect 1246 331 1247 335
rect 1251 331 1252 335
rect 1806 332 1807 336
rect 1811 332 1812 336
rect 2062 333 2063 337
rect 2067 333 2068 337
rect 2062 332 2068 333
rect 2150 337 2156 338
rect 2150 333 2151 337
rect 2155 333 2156 337
rect 2150 332 2156 333
rect 2246 337 2252 338
rect 2246 333 2247 337
rect 2251 333 2252 337
rect 2246 332 2252 333
rect 2358 337 2364 338
rect 2358 333 2359 337
rect 2363 333 2364 337
rect 2358 332 2364 333
rect 1806 331 1812 332
rect 1246 330 1252 331
rect 646 325 652 326
rect 646 321 647 325
rect 651 321 652 325
rect 646 320 652 321
rect 734 325 740 326
rect 734 321 735 325
rect 739 321 740 325
rect 734 320 740 321
rect 822 325 828 326
rect 822 321 823 325
rect 827 321 828 325
rect 822 320 828 321
rect 648 299 650 320
rect 736 299 738 320
rect 824 299 826 320
rect 647 298 651 299
rect 647 293 651 294
rect 655 298 659 299
rect 655 293 659 294
rect 735 298 739 299
rect 735 293 739 294
rect 751 298 755 299
rect 751 293 755 294
rect 823 298 827 299
rect 823 293 827 294
rect 847 298 851 299
rect 847 293 851 294
rect 656 276 658 293
rect 752 276 754 293
rect 848 276 850 293
rect 654 275 660 276
rect 654 271 655 275
rect 659 271 660 275
rect 654 270 660 271
rect 750 275 756 276
rect 750 271 751 275
rect 755 271 756 275
rect 750 270 756 271
rect 846 275 852 276
rect 846 271 847 275
rect 851 271 852 275
rect 846 270 852 271
rect 638 267 644 268
rect 350 263 356 264
rect 110 259 116 260
rect 110 255 111 259
rect 115 255 116 259
rect 350 259 351 263
rect 355 259 356 263
rect 350 258 356 259
rect 438 263 444 264
rect 438 259 439 263
rect 443 259 444 263
rect 438 258 444 259
rect 534 263 540 264
rect 534 259 535 263
rect 539 259 540 263
rect 534 258 540 259
rect 630 263 636 264
rect 630 259 631 263
rect 635 259 636 263
rect 638 263 639 267
rect 643 263 644 267
rect 638 262 644 263
rect 822 263 828 264
rect 630 258 636 259
rect 822 259 823 263
rect 827 259 828 263
rect 822 258 828 259
rect 110 254 116 255
rect 278 256 284 257
rect 112 231 114 254
rect 278 252 279 256
rect 283 252 284 256
rect 278 251 284 252
rect 280 231 282 251
rect 352 240 354 258
rect 366 256 372 257
rect 366 252 367 256
rect 371 252 372 256
rect 366 251 372 252
rect 350 239 356 240
rect 350 235 351 239
rect 355 235 356 239
rect 350 234 356 235
rect 368 231 370 251
rect 440 240 442 258
rect 462 256 468 257
rect 462 252 463 256
rect 467 252 468 256
rect 462 251 468 252
rect 438 239 444 240
rect 438 235 439 239
rect 443 235 444 239
rect 438 234 444 235
rect 464 231 466 251
rect 536 240 538 258
rect 558 256 564 257
rect 558 252 559 256
rect 563 252 564 256
rect 558 251 564 252
rect 534 239 540 240
rect 534 235 535 239
rect 539 235 540 239
rect 534 234 540 235
rect 560 231 562 251
rect 632 240 634 258
rect 654 256 660 257
rect 654 252 655 256
rect 659 252 660 256
rect 654 251 660 252
rect 750 256 756 257
rect 750 252 751 256
rect 755 252 756 256
rect 750 251 756 252
rect 630 239 636 240
rect 630 235 631 239
rect 635 235 636 239
rect 630 234 636 235
rect 590 231 596 232
rect 656 231 658 251
rect 752 231 754 251
rect 824 240 826 258
rect 846 256 852 257
rect 846 252 847 256
rect 851 252 852 256
rect 846 251 852 252
rect 822 239 828 240
rect 822 235 823 239
rect 827 235 828 239
rect 822 234 828 235
rect 848 231 850 251
rect 904 248 906 330
rect 910 325 916 326
rect 910 321 911 325
rect 915 321 916 325
rect 910 320 916 321
rect 998 325 1004 326
rect 998 321 999 325
rect 1003 321 1004 325
rect 998 320 1004 321
rect 1086 325 1092 326
rect 1086 321 1087 325
rect 1091 321 1092 325
rect 1086 320 1092 321
rect 1174 325 1180 326
rect 1174 321 1175 325
rect 1179 321 1180 325
rect 1174 320 1180 321
rect 1262 325 1268 326
rect 1262 321 1263 325
rect 1267 321 1268 325
rect 1262 320 1268 321
rect 1766 324 1772 325
rect 1766 320 1767 324
rect 1771 320 1772 324
rect 912 299 914 320
rect 1000 299 1002 320
rect 1088 299 1090 320
rect 1176 299 1178 320
rect 1264 299 1266 320
rect 1766 319 1772 320
rect 1768 299 1770 319
rect 1808 311 1810 331
rect 2064 311 2066 332
rect 2152 311 2154 332
rect 2248 311 2250 332
rect 2360 311 2362 332
rect 1807 310 1811 311
rect 1807 305 1811 306
rect 1927 310 1931 311
rect 1927 305 1931 306
rect 2039 310 2043 311
rect 2039 305 2043 306
rect 2063 310 2067 311
rect 2063 305 2067 306
rect 2151 310 2155 311
rect 2151 305 2155 306
rect 2167 310 2171 311
rect 2167 305 2171 306
rect 2247 310 2251 311
rect 2247 305 2251 306
rect 2303 310 2307 311
rect 2303 305 2307 306
rect 2359 310 2363 311
rect 2359 305 2363 306
rect 911 298 915 299
rect 911 293 915 294
rect 943 298 947 299
rect 943 293 947 294
rect 999 298 1003 299
rect 999 293 1003 294
rect 1047 298 1051 299
rect 1047 293 1051 294
rect 1087 298 1091 299
rect 1087 293 1091 294
rect 1151 298 1155 299
rect 1151 293 1155 294
rect 1175 298 1179 299
rect 1175 293 1179 294
rect 1263 298 1267 299
rect 1263 293 1267 294
rect 1767 298 1771 299
rect 1767 293 1771 294
rect 944 276 946 293
rect 1048 276 1050 293
rect 1152 276 1154 293
rect 1768 277 1770 293
rect 1808 289 1810 305
rect 1806 288 1812 289
rect 1928 288 1930 305
rect 2040 288 2042 305
rect 2168 288 2170 305
rect 2304 288 2306 305
rect 1806 284 1807 288
rect 1811 284 1812 288
rect 1806 283 1812 284
rect 1926 287 1932 288
rect 1926 283 1927 287
rect 1931 283 1932 287
rect 1926 282 1932 283
rect 2038 287 2044 288
rect 2038 283 2039 287
rect 2043 283 2044 287
rect 2038 282 2044 283
rect 2166 287 2172 288
rect 2166 283 2167 287
rect 2171 283 2172 287
rect 2166 282 2172 283
rect 2302 287 2308 288
rect 2302 283 2303 287
rect 2307 283 2308 287
rect 2302 282 2308 283
rect 2424 280 2426 358
rect 2432 348 2434 366
rect 2440 348 2442 374
rect 2447 373 2451 374
rect 2479 378 2483 379
rect 2479 373 2483 374
rect 2559 378 2563 379
rect 2559 373 2563 374
rect 2615 378 2619 379
rect 2615 373 2619 374
rect 2679 378 2683 379
rect 2679 373 2683 374
rect 2759 378 2763 379
rect 2759 373 2763 374
rect 2799 378 2803 379
rect 2799 373 2803 374
rect 2480 357 2482 373
rect 2616 357 2618 373
rect 2694 371 2700 372
rect 2694 367 2695 371
rect 2699 367 2700 371
rect 2694 366 2700 367
rect 2478 356 2484 357
rect 2478 352 2479 356
rect 2483 352 2484 356
rect 2478 351 2484 352
rect 2614 356 2620 357
rect 2614 352 2615 356
rect 2619 352 2620 356
rect 2614 351 2620 352
rect 2696 348 2698 366
rect 2760 357 2762 373
rect 2872 372 2874 406
rect 2910 404 2916 405
rect 2910 400 2911 404
rect 2915 400 2916 404
rect 2910 399 2916 400
rect 2912 379 2914 399
rect 2984 388 2986 406
rect 3022 404 3028 405
rect 3022 400 3023 404
rect 3027 400 3028 404
rect 3022 399 3028 400
rect 2974 387 2980 388
rect 2974 383 2975 387
rect 2979 383 2980 387
rect 2974 382 2980 383
rect 2982 387 2988 388
rect 2982 383 2983 387
rect 2987 383 2988 387
rect 2982 382 2988 383
rect 2911 378 2915 379
rect 2911 373 2915 374
rect 2870 371 2876 372
rect 2870 367 2871 371
rect 2875 367 2876 371
rect 2870 366 2876 367
rect 2912 357 2914 373
rect 2758 356 2764 357
rect 2758 352 2759 356
rect 2763 352 2764 356
rect 2758 351 2764 352
rect 2910 356 2916 357
rect 2910 352 2911 356
rect 2915 352 2916 356
rect 2910 351 2916 352
rect 2976 348 2978 382
rect 3024 379 3026 399
rect 3096 388 3098 406
rect 3142 404 3148 405
rect 3142 400 3143 404
rect 3147 400 3148 404
rect 3142 399 3148 400
rect 3262 404 3268 405
rect 3262 400 3263 404
rect 3267 400 3268 404
rect 3262 399 3268 400
rect 3094 387 3100 388
rect 3094 383 3095 387
rect 3099 383 3100 387
rect 3094 382 3100 383
rect 3144 379 3146 399
rect 3264 379 3266 399
rect 3328 388 3330 482
rect 3366 477 3372 478
rect 3366 473 3367 477
rect 3371 473 3372 477
rect 3366 472 3372 473
rect 3368 447 3370 472
rect 3367 446 3371 447
rect 3367 441 3371 442
rect 3368 424 3370 441
rect 3366 423 3372 424
rect 3366 419 3367 423
rect 3371 419 3372 423
rect 3366 418 3372 419
rect 3440 416 3442 506
rect 3464 494 3466 513
rect 3462 493 3468 494
rect 3462 489 3463 493
rect 3467 489 3468 493
rect 3462 488 3468 489
rect 3462 476 3468 477
rect 3462 472 3463 476
rect 3467 472 3468 476
rect 3462 471 3468 472
rect 3464 447 3466 471
rect 3463 446 3467 447
rect 3463 441 3467 442
rect 3464 425 3466 441
rect 3462 424 3468 425
rect 3462 420 3463 424
rect 3467 420 3468 424
rect 3462 419 3468 420
rect 3438 415 3444 416
rect 3334 411 3340 412
rect 3334 407 3335 411
rect 3339 407 3340 411
rect 3438 411 3439 415
rect 3443 411 3444 415
rect 3438 410 3444 411
rect 3334 406 3340 407
rect 3462 407 3468 408
rect 3326 387 3332 388
rect 3326 383 3327 387
rect 3331 383 3332 387
rect 3326 382 3332 383
rect 3023 378 3027 379
rect 3023 373 3027 374
rect 3063 378 3067 379
rect 3063 373 3067 374
rect 3143 378 3147 379
rect 3143 373 3147 374
rect 3223 378 3227 379
rect 3223 373 3227 374
rect 3263 378 3267 379
rect 3263 373 3267 374
rect 2990 371 2996 372
rect 2990 367 2991 371
rect 2995 367 2996 371
rect 2990 366 2996 367
rect 2992 348 2994 366
rect 3064 357 3066 373
rect 3158 371 3164 372
rect 3158 367 3159 371
rect 3163 367 3164 371
rect 3158 366 3164 367
rect 3166 371 3172 372
rect 3166 367 3167 371
rect 3171 367 3172 371
rect 3166 366 3172 367
rect 3062 356 3068 357
rect 3062 352 3063 356
rect 3067 352 3068 356
rect 3062 351 3068 352
rect 3160 348 3162 366
rect 2430 347 2436 348
rect 2430 343 2431 347
rect 2435 343 2436 347
rect 2430 342 2436 343
rect 2438 347 2444 348
rect 2438 343 2439 347
rect 2443 343 2444 347
rect 2438 342 2444 343
rect 2678 347 2684 348
rect 2678 343 2679 347
rect 2683 343 2684 347
rect 2678 342 2684 343
rect 2694 347 2700 348
rect 2694 343 2695 347
rect 2699 343 2700 347
rect 2694 342 2700 343
rect 2974 347 2980 348
rect 2974 343 2975 347
rect 2979 343 2980 347
rect 2974 342 2980 343
rect 2990 347 2996 348
rect 2990 343 2991 347
rect 2995 343 2996 347
rect 2990 342 2996 343
rect 3158 347 3164 348
rect 3158 343 3159 347
rect 3163 343 3164 347
rect 3158 342 3164 343
rect 2478 337 2484 338
rect 2478 333 2479 337
rect 2483 333 2484 337
rect 2478 332 2484 333
rect 2614 337 2620 338
rect 2614 333 2615 337
rect 2619 333 2620 337
rect 2614 332 2620 333
rect 2480 311 2482 332
rect 2616 311 2618 332
rect 2447 310 2451 311
rect 2447 305 2451 306
rect 2479 310 2483 311
rect 2479 305 2483 306
rect 2599 310 2603 311
rect 2599 305 2603 306
rect 2615 310 2619 311
rect 2615 305 2619 306
rect 2448 288 2450 305
rect 2600 288 2602 305
rect 2446 287 2452 288
rect 2446 283 2447 287
rect 2451 283 2452 287
rect 2446 282 2452 283
rect 2598 287 2604 288
rect 2598 283 2599 287
rect 2603 283 2604 287
rect 2598 282 2604 283
rect 2422 279 2428 280
rect 1766 276 1772 277
rect 942 275 948 276
rect 942 271 943 275
rect 947 271 948 275
rect 942 270 948 271
rect 1046 275 1052 276
rect 1046 271 1047 275
rect 1051 271 1052 275
rect 1046 270 1052 271
rect 1150 275 1156 276
rect 1150 271 1151 275
rect 1155 271 1156 275
rect 1766 272 1767 276
rect 1771 272 1772 276
rect 1998 275 2004 276
rect 1766 271 1772 272
rect 1806 271 1812 272
rect 1150 270 1156 271
rect 1126 267 1132 268
rect 918 263 924 264
rect 918 259 919 263
rect 923 259 924 263
rect 918 258 924 259
rect 1014 263 1020 264
rect 1014 259 1015 263
rect 1019 259 1020 263
rect 1014 258 1020 259
rect 1118 263 1124 264
rect 1118 259 1119 263
rect 1123 259 1124 263
rect 1126 263 1127 267
rect 1131 263 1132 267
rect 1806 267 1807 271
rect 1811 267 1812 271
rect 1998 271 1999 275
rect 2003 271 2004 275
rect 1998 270 2004 271
rect 2110 275 2116 276
rect 2110 271 2111 275
rect 2115 271 2116 275
rect 2110 270 2116 271
rect 2238 275 2244 276
rect 2238 271 2239 275
rect 2243 271 2244 275
rect 2238 270 2244 271
rect 2374 275 2380 276
rect 2374 271 2375 275
rect 2379 271 2380 275
rect 2422 275 2423 279
rect 2427 275 2428 279
rect 2422 274 2428 275
rect 2670 275 2676 276
rect 2374 270 2380 271
rect 2670 271 2671 275
rect 2675 271 2676 275
rect 2670 270 2676 271
rect 1806 266 1812 267
rect 1926 268 1932 269
rect 1126 262 1132 263
rect 1118 258 1124 259
rect 902 247 908 248
rect 902 243 903 247
rect 907 243 908 247
rect 902 242 908 243
rect 920 240 922 258
rect 942 256 948 257
rect 942 252 943 256
rect 947 252 948 256
rect 942 251 948 252
rect 918 239 924 240
rect 918 235 919 239
rect 923 235 924 239
rect 918 234 924 235
rect 944 231 946 251
rect 1016 240 1018 258
rect 1046 256 1052 257
rect 1046 252 1047 256
rect 1051 252 1052 256
rect 1046 251 1052 252
rect 1014 239 1020 240
rect 1014 235 1015 239
rect 1019 235 1020 239
rect 1014 234 1020 235
rect 1048 231 1050 251
rect 1120 240 1122 258
rect 1118 239 1124 240
rect 1118 235 1119 239
rect 1123 235 1124 239
rect 1118 234 1124 235
rect 1128 232 1130 262
rect 1766 259 1772 260
rect 1150 256 1156 257
rect 1150 252 1151 256
rect 1155 252 1156 256
rect 1766 255 1767 259
rect 1771 255 1772 259
rect 1766 254 1772 255
rect 1150 251 1156 252
rect 1126 231 1132 232
rect 1152 231 1154 251
rect 1768 231 1770 254
rect 1808 243 1810 266
rect 1926 264 1927 268
rect 1931 264 1932 268
rect 1926 263 1932 264
rect 1928 243 1930 263
rect 2000 252 2002 270
rect 2038 268 2044 269
rect 2038 264 2039 268
rect 2043 264 2044 268
rect 2038 263 2044 264
rect 1998 251 2004 252
rect 1998 247 1999 251
rect 2003 247 2004 251
rect 1998 246 2004 247
rect 2040 243 2042 263
rect 2112 252 2114 270
rect 2166 268 2172 269
rect 2166 264 2167 268
rect 2171 264 2172 268
rect 2166 263 2172 264
rect 2110 251 2116 252
rect 2110 247 2111 251
rect 2115 247 2116 251
rect 2110 246 2116 247
rect 2168 243 2170 263
rect 2240 252 2242 270
rect 2302 268 2308 269
rect 2302 264 2303 268
rect 2307 264 2308 268
rect 2302 263 2308 264
rect 2238 251 2244 252
rect 2238 247 2239 251
rect 2243 247 2244 251
rect 2238 246 2244 247
rect 2304 243 2306 263
rect 2376 252 2378 270
rect 2446 268 2452 269
rect 2446 264 2447 268
rect 2451 264 2452 268
rect 2446 263 2452 264
rect 2598 268 2604 269
rect 2598 264 2599 268
rect 2603 264 2604 268
rect 2598 263 2604 264
rect 2374 251 2380 252
rect 2374 247 2375 251
rect 2379 247 2380 251
rect 2374 246 2380 247
rect 2322 243 2328 244
rect 2448 243 2450 263
rect 2600 243 2602 263
rect 1807 242 1811 243
rect 1807 237 1811 238
rect 1831 242 1835 243
rect 1831 237 1835 238
rect 1927 242 1931 243
rect 1927 237 1931 238
rect 2039 242 2043 243
rect 2039 237 2043 238
rect 2055 242 2059 243
rect 2055 237 2059 238
rect 2167 242 2171 243
rect 2167 237 2171 238
rect 2199 242 2203 243
rect 2199 237 2203 238
rect 2303 242 2307 243
rect 2322 239 2323 243
rect 2327 239 2328 243
rect 2322 238 2328 239
rect 2351 242 2355 243
rect 2303 237 2307 238
rect 111 230 115 231
rect 111 225 115 226
rect 167 230 171 231
rect 167 225 171 226
rect 279 230 283 231
rect 279 225 283 226
rect 343 230 347 231
rect 343 225 347 226
rect 367 230 371 231
rect 367 225 371 226
rect 463 230 467 231
rect 463 225 467 226
rect 511 230 515 231
rect 511 225 515 226
rect 559 230 563 231
rect 590 227 591 231
rect 595 227 596 231
rect 590 226 596 227
rect 655 230 659 231
rect 559 225 563 226
rect 112 206 114 225
rect 168 209 170 225
rect 230 223 236 224
rect 230 219 231 223
rect 235 219 236 223
rect 230 218 236 219
rect 238 223 244 224
rect 238 219 239 223
rect 243 219 244 223
rect 238 218 244 219
rect 166 208 172 209
rect 110 205 116 206
rect 110 201 111 205
rect 115 201 116 205
rect 166 204 167 208
rect 171 204 172 208
rect 166 203 172 204
rect 110 200 116 201
rect 166 189 172 190
rect 110 188 116 189
rect 110 184 111 188
rect 115 184 116 188
rect 166 185 167 189
rect 171 185 172 189
rect 166 184 172 185
rect 110 183 116 184
rect 112 143 114 183
rect 168 143 170 184
rect 232 165 234 218
rect 240 200 242 218
rect 344 209 346 225
rect 414 223 420 224
rect 414 219 415 223
rect 419 219 420 223
rect 414 218 420 219
rect 342 208 348 209
rect 342 204 343 208
rect 347 204 348 208
rect 342 203 348 204
rect 416 200 418 218
rect 512 209 514 225
rect 582 223 588 224
rect 582 219 583 223
rect 587 219 588 223
rect 582 218 588 219
rect 510 208 516 209
rect 510 204 511 208
rect 515 204 516 208
rect 510 203 516 204
rect 584 200 586 218
rect 592 200 594 226
rect 655 225 659 226
rect 679 230 683 231
rect 679 225 683 226
rect 751 230 755 231
rect 751 225 755 226
rect 839 230 843 231
rect 839 225 843 226
rect 847 230 851 231
rect 847 225 851 226
rect 943 230 947 231
rect 943 225 947 226
rect 991 230 995 231
rect 991 225 995 226
rect 1047 230 1051 231
rect 1126 227 1127 231
rect 1131 227 1132 231
rect 1126 226 1132 227
rect 1135 230 1139 231
rect 1047 225 1051 226
rect 1135 225 1139 226
rect 1151 230 1155 231
rect 1151 225 1155 226
rect 1279 230 1283 231
rect 1279 225 1283 226
rect 1431 230 1435 231
rect 1431 225 1435 226
rect 1767 230 1771 231
rect 1767 225 1771 226
rect 680 209 682 225
rect 840 209 842 225
rect 910 223 916 224
rect 910 219 911 223
rect 915 219 916 223
rect 910 218 916 219
rect 678 208 684 209
rect 678 204 679 208
rect 683 204 684 208
rect 678 203 684 204
rect 838 208 844 209
rect 838 204 839 208
rect 843 204 844 208
rect 838 203 844 204
rect 912 200 914 218
rect 992 209 994 225
rect 1062 223 1068 224
rect 1062 219 1063 223
rect 1067 219 1068 223
rect 1062 218 1068 219
rect 990 208 996 209
rect 990 204 991 208
rect 995 204 996 208
rect 990 203 996 204
rect 1064 200 1066 218
rect 1136 209 1138 225
rect 1206 223 1212 224
rect 1206 219 1207 223
rect 1211 219 1212 223
rect 1206 218 1212 219
rect 1134 208 1140 209
rect 1134 204 1135 208
rect 1139 204 1140 208
rect 1134 203 1140 204
rect 1208 200 1210 218
rect 1280 209 1282 225
rect 1350 223 1356 224
rect 1350 219 1351 223
rect 1355 219 1356 223
rect 1350 218 1356 219
rect 1278 208 1284 209
rect 1278 204 1279 208
rect 1283 204 1284 208
rect 1278 203 1284 204
rect 1352 200 1354 218
rect 1432 209 1434 225
rect 1430 208 1436 209
rect 1430 204 1431 208
rect 1435 204 1436 208
rect 1768 206 1770 225
rect 1808 218 1810 237
rect 1832 221 1834 237
rect 1902 235 1908 236
rect 1902 231 1903 235
rect 1907 231 1908 235
rect 1902 230 1908 231
rect 1830 220 1836 221
rect 1806 217 1812 218
rect 1806 213 1807 217
rect 1811 213 1812 217
rect 1830 216 1831 220
rect 1835 216 1836 220
rect 1830 215 1836 216
rect 1806 212 1812 213
rect 1904 212 1906 230
rect 1928 221 1930 237
rect 1998 235 2004 236
rect 1998 231 1999 235
rect 2003 231 2004 235
rect 1998 230 2004 231
rect 1926 220 1932 221
rect 1926 216 1927 220
rect 1931 216 1932 220
rect 1926 215 1932 216
rect 2000 212 2002 230
rect 2056 221 2058 237
rect 2126 235 2132 236
rect 2126 231 2127 235
rect 2131 231 2132 235
rect 2126 230 2132 231
rect 2054 220 2060 221
rect 2054 216 2055 220
rect 2059 216 2060 220
rect 2054 215 2060 216
rect 2128 212 2130 230
rect 2200 221 2202 237
rect 2270 235 2276 236
rect 2270 231 2271 235
rect 2275 231 2276 235
rect 2270 230 2276 231
rect 2238 227 2244 228
rect 2238 223 2239 227
rect 2243 223 2244 227
rect 2238 222 2244 223
rect 2198 220 2204 221
rect 2198 216 2199 220
rect 2203 216 2204 220
rect 2198 215 2204 216
rect 1902 211 1908 212
rect 1902 207 1903 211
rect 1907 207 1908 211
rect 1902 206 1908 207
rect 1998 211 2004 212
rect 1998 207 1999 211
rect 2003 207 2004 211
rect 1998 206 2004 207
rect 2126 211 2132 212
rect 2126 207 2127 211
rect 2131 207 2132 211
rect 2126 206 2132 207
rect 1430 203 1436 204
rect 1766 205 1772 206
rect 1766 201 1767 205
rect 1771 201 1772 205
rect 1830 201 1836 202
rect 1766 200 1772 201
rect 1806 200 1812 201
rect 238 199 244 200
rect 238 195 239 199
rect 243 195 244 199
rect 238 194 244 195
rect 414 199 420 200
rect 414 195 415 199
rect 419 195 420 199
rect 414 194 420 195
rect 582 199 588 200
rect 582 195 583 199
rect 587 195 588 199
rect 582 194 588 195
rect 590 199 596 200
rect 590 195 591 199
rect 595 195 596 199
rect 590 194 596 195
rect 910 199 916 200
rect 910 195 911 199
rect 915 195 916 199
rect 910 194 916 195
rect 1062 199 1068 200
rect 1062 195 1063 199
rect 1067 195 1068 199
rect 1062 194 1068 195
rect 1206 199 1212 200
rect 1206 195 1207 199
rect 1211 195 1212 199
rect 1206 194 1212 195
rect 1350 199 1356 200
rect 1350 195 1351 199
rect 1355 195 1356 199
rect 1350 194 1356 195
rect 1398 199 1404 200
rect 1398 195 1399 199
rect 1403 195 1404 199
rect 1806 196 1807 200
rect 1811 196 1812 200
rect 1830 197 1831 201
rect 1835 197 1836 201
rect 1830 196 1836 197
rect 1926 201 1932 202
rect 1926 197 1927 201
rect 1931 197 1932 201
rect 1926 196 1932 197
rect 2054 201 2060 202
rect 2054 197 2055 201
rect 2059 197 2060 201
rect 2054 196 2060 197
rect 2198 201 2204 202
rect 2198 197 2199 201
rect 2203 197 2204 201
rect 2198 196 2204 197
rect 1806 195 1812 196
rect 1398 194 1404 195
rect 342 189 348 190
rect 342 185 343 189
rect 347 185 348 189
rect 342 184 348 185
rect 510 189 516 190
rect 510 185 511 189
rect 515 185 516 189
rect 510 184 516 185
rect 678 189 684 190
rect 678 185 679 189
rect 683 185 684 189
rect 678 184 684 185
rect 838 189 844 190
rect 838 185 839 189
rect 843 185 844 189
rect 838 184 844 185
rect 990 189 996 190
rect 990 185 991 189
rect 995 185 996 189
rect 990 184 996 185
rect 1134 189 1140 190
rect 1134 185 1135 189
rect 1139 185 1140 189
rect 1134 184 1140 185
rect 1278 189 1284 190
rect 1278 185 1279 189
rect 1283 185 1284 189
rect 1278 184 1284 185
rect 231 164 235 165
rect 231 159 235 160
rect 344 143 346 184
rect 512 143 514 184
rect 680 143 682 184
rect 743 164 747 165
rect 743 159 747 160
rect 111 142 115 143
rect 111 137 115 138
rect 135 142 139 143
rect 135 137 139 138
rect 167 142 171 143
rect 167 137 171 138
rect 223 142 227 143
rect 223 137 227 138
rect 311 142 315 143
rect 311 137 315 138
rect 343 142 347 143
rect 343 137 347 138
rect 399 142 403 143
rect 399 137 403 138
rect 487 142 491 143
rect 487 137 491 138
rect 511 142 515 143
rect 511 137 515 138
rect 575 142 579 143
rect 575 137 579 138
rect 663 142 667 143
rect 663 137 667 138
rect 679 142 683 143
rect 679 137 683 138
rect 112 121 114 137
rect 110 120 116 121
rect 136 120 138 137
rect 224 120 226 137
rect 312 120 314 137
rect 400 120 402 137
rect 488 120 490 137
rect 576 120 578 137
rect 664 120 666 137
rect 110 116 111 120
rect 115 116 116 120
rect 110 115 116 116
rect 134 119 140 120
rect 134 115 135 119
rect 139 115 140 119
rect 134 114 140 115
rect 222 119 228 120
rect 222 115 223 119
rect 227 115 228 119
rect 222 114 228 115
rect 310 119 316 120
rect 310 115 311 119
rect 315 115 316 119
rect 310 114 316 115
rect 398 119 404 120
rect 398 115 399 119
rect 403 115 404 119
rect 398 114 404 115
rect 486 119 492 120
rect 486 115 487 119
rect 491 115 492 119
rect 486 114 492 115
rect 574 119 580 120
rect 574 115 575 119
rect 579 115 580 119
rect 574 114 580 115
rect 662 119 668 120
rect 662 115 663 119
rect 667 115 668 119
rect 662 114 668 115
rect 744 112 746 159
rect 840 143 842 184
rect 992 143 994 184
rect 1136 143 1138 184
rect 1280 143 1282 184
rect 751 142 755 143
rect 751 137 755 138
rect 839 142 843 143
rect 839 137 843 138
rect 847 142 851 143
rect 847 137 851 138
rect 943 142 947 143
rect 943 137 947 138
rect 991 142 995 143
rect 991 137 995 138
rect 1031 142 1035 143
rect 1031 137 1035 138
rect 1119 142 1123 143
rect 1119 137 1123 138
rect 1135 142 1139 143
rect 1135 137 1139 138
rect 1215 142 1219 143
rect 1215 137 1219 138
rect 1279 142 1283 143
rect 1279 137 1283 138
rect 1311 142 1315 143
rect 1311 137 1315 138
rect 752 120 754 137
rect 848 120 850 137
rect 944 120 946 137
rect 1032 120 1034 137
rect 1120 120 1122 137
rect 1216 120 1218 137
rect 1312 120 1314 137
rect 750 119 756 120
rect 750 115 751 119
rect 755 115 756 119
rect 750 114 756 115
rect 846 119 852 120
rect 846 115 847 119
rect 851 115 852 119
rect 846 114 852 115
rect 942 119 948 120
rect 942 115 943 119
rect 947 115 948 119
rect 942 114 948 115
rect 1030 119 1036 120
rect 1030 115 1031 119
rect 1035 115 1036 119
rect 1030 114 1036 115
rect 1118 119 1124 120
rect 1118 115 1119 119
rect 1123 115 1124 119
rect 1118 114 1124 115
rect 1214 119 1220 120
rect 1214 115 1215 119
rect 1219 115 1220 119
rect 1214 114 1220 115
rect 1310 119 1316 120
rect 1310 115 1311 119
rect 1315 115 1316 119
rect 1310 114 1316 115
rect 742 111 748 112
rect 206 107 212 108
rect 110 103 116 104
rect 110 99 111 103
rect 115 99 116 103
rect 206 103 207 107
rect 211 103 212 107
rect 206 102 212 103
rect 294 107 300 108
rect 294 103 295 107
rect 299 103 300 107
rect 294 102 300 103
rect 382 107 388 108
rect 382 103 383 107
rect 387 103 388 107
rect 382 102 388 103
rect 470 107 476 108
rect 470 103 471 107
rect 475 103 476 107
rect 470 102 476 103
rect 558 107 564 108
rect 558 103 559 107
rect 563 103 564 107
rect 558 102 564 103
rect 646 107 652 108
rect 646 103 647 107
rect 651 103 652 107
rect 646 102 652 103
rect 734 107 740 108
rect 734 103 735 107
rect 739 103 740 107
rect 742 107 743 111
rect 747 107 748 111
rect 742 106 748 107
rect 918 107 924 108
rect 734 102 740 103
rect 918 103 919 107
rect 923 103 924 107
rect 918 102 924 103
rect 1014 107 1020 108
rect 1014 103 1015 107
rect 1019 103 1020 107
rect 1014 102 1020 103
rect 1102 107 1108 108
rect 1102 103 1103 107
rect 1107 103 1108 107
rect 1102 102 1108 103
rect 1190 107 1196 108
rect 1190 103 1191 107
rect 1195 103 1196 107
rect 1190 102 1196 103
rect 1286 107 1292 108
rect 1286 103 1287 107
rect 1291 103 1292 107
rect 1286 102 1292 103
rect 1382 107 1388 108
rect 1382 103 1383 107
rect 1387 103 1388 107
rect 1382 102 1388 103
rect 110 98 116 99
rect 134 100 140 101
rect 112 79 114 98
rect 134 96 135 100
rect 139 96 140 100
rect 134 95 140 96
rect 136 79 138 95
rect 208 84 210 102
rect 222 100 228 101
rect 222 96 223 100
rect 227 96 228 100
rect 222 95 228 96
rect 206 83 212 84
rect 206 79 207 83
rect 211 79 212 83
rect 224 79 226 95
rect 296 84 298 102
rect 310 100 316 101
rect 310 96 311 100
rect 315 96 316 100
rect 310 95 316 96
rect 294 83 300 84
rect 294 79 295 83
rect 299 79 300 83
rect 312 79 314 95
rect 384 84 386 102
rect 398 100 404 101
rect 398 96 399 100
rect 403 96 404 100
rect 398 95 404 96
rect 382 83 388 84
rect 382 79 383 83
rect 387 79 388 83
rect 400 79 402 95
rect 472 84 474 102
rect 486 100 492 101
rect 486 96 487 100
rect 491 96 492 100
rect 486 95 492 96
rect 470 83 476 84
rect 470 79 471 83
rect 475 79 476 83
rect 488 79 490 95
rect 560 84 562 102
rect 574 100 580 101
rect 574 96 575 100
rect 579 96 580 100
rect 574 95 580 96
rect 558 83 564 84
rect 558 79 559 83
rect 563 79 564 83
rect 576 79 578 95
rect 648 84 650 102
rect 662 100 668 101
rect 662 96 663 100
rect 667 96 668 100
rect 662 95 668 96
rect 646 83 652 84
rect 646 79 647 83
rect 651 79 652 83
rect 664 79 666 95
rect 736 84 738 102
rect 750 100 756 101
rect 750 96 751 100
rect 755 96 756 100
rect 750 95 756 96
rect 846 100 852 101
rect 846 96 847 100
rect 851 96 852 100
rect 846 95 852 96
rect 734 83 740 84
rect 734 79 735 83
rect 739 79 740 83
rect 752 79 754 95
rect 848 79 850 95
rect 903 92 907 93
rect 903 87 907 88
rect 904 84 906 87
rect 920 84 922 102
rect 942 100 948 101
rect 942 96 943 100
rect 947 96 948 100
rect 942 95 948 96
rect 902 83 908 84
rect 902 79 903 83
rect 907 79 908 83
rect 111 78 115 79
rect 111 73 115 74
rect 135 78 139 79
rect 206 78 212 79
rect 223 78 227 79
rect 294 78 300 79
rect 311 78 315 79
rect 382 78 388 79
rect 399 78 403 79
rect 470 78 476 79
rect 487 78 491 79
rect 558 78 564 79
rect 575 78 579 79
rect 646 78 652 79
rect 663 78 667 79
rect 734 78 740 79
rect 751 78 755 79
rect 135 73 139 74
rect 223 73 227 74
rect 311 73 315 74
rect 399 73 403 74
rect 487 73 491 74
rect 575 73 579 74
rect 663 73 667 74
rect 751 73 755 74
rect 847 78 851 79
rect 902 78 908 79
rect 918 83 924 84
rect 918 79 919 83
rect 923 79 924 83
rect 944 79 946 95
rect 1016 84 1018 102
rect 1030 100 1036 101
rect 1030 96 1031 100
rect 1035 96 1036 100
rect 1030 95 1036 96
rect 1014 83 1020 84
rect 1014 79 1015 83
rect 1019 79 1020 83
rect 1032 79 1034 95
rect 1104 84 1106 102
rect 1118 100 1124 101
rect 1118 96 1119 100
rect 1123 96 1124 100
rect 1118 95 1124 96
rect 1102 83 1108 84
rect 1102 79 1103 83
rect 1107 79 1108 83
rect 1120 79 1122 95
rect 1192 84 1194 102
rect 1214 100 1220 101
rect 1214 96 1215 100
rect 1219 96 1220 100
rect 1214 95 1220 96
rect 1190 83 1196 84
rect 1190 79 1191 83
rect 1195 79 1196 83
rect 1216 79 1218 95
rect 1288 84 1290 102
rect 1310 100 1316 101
rect 1310 96 1311 100
rect 1315 96 1316 100
rect 1310 95 1316 96
rect 1286 83 1292 84
rect 1286 79 1287 83
rect 1291 79 1292 83
rect 1312 79 1314 95
rect 1384 84 1386 102
rect 1400 93 1402 194
rect 1430 189 1436 190
rect 1430 185 1431 189
rect 1435 185 1436 189
rect 1430 184 1436 185
rect 1766 188 1772 189
rect 1766 184 1767 188
rect 1771 184 1772 188
rect 1432 143 1434 184
rect 1766 183 1772 184
rect 1768 143 1770 183
rect 1808 159 1810 195
rect 1832 159 1834 196
rect 1928 159 1930 196
rect 2056 159 2058 196
rect 2200 159 2202 196
rect 1807 158 1811 159
rect 1807 153 1811 154
rect 1831 158 1835 159
rect 1831 153 1835 154
rect 1919 158 1923 159
rect 1919 153 1923 154
rect 1927 158 1931 159
rect 1927 153 1931 154
rect 2039 158 2043 159
rect 2039 153 2043 154
rect 2055 158 2059 159
rect 2055 153 2059 154
rect 2159 158 2163 159
rect 2159 153 2163 154
rect 2199 158 2203 159
rect 2199 153 2203 154
rect 1407 142 1411 143
rect 1407 137 1411 138
rect 1431 142 1435 143
rect 1431 137 1435 138
rect 1495 142 1499 143
rect 1495 137 1499 138
rect 1583 142 1587 143
rect 1583 137 1587 138
rect 1671 142 1675 143
rect 1671 137 1675 138
rect 1767 142 1771 143
rect 1767 137 1771 138
rect 1808 137 1810 153
rect 1408 120 1410 137
rect 1496 120 1498 137
rect 1584 120 1586 137
rect 1672 120 1674 137
rect 1768 121 1770 137
rect 1806 136 1812 137
rect 1832 136 1834 153
rect 1920 136 1922 153
rect 2040 136 2042 153
rect 2160 136 2162 153
rect 1806 132 1807 136
rect 1811 132 1812 136
rect 1806 131 1812 132
rect 1830 135 1836 136
rect 1830 131 1831 135
rect 1835 131 1836 135
rect 1830 130 1836 131
rect 1918 135 1924 136
rect 1918 131 1919 135
rect 1923 131 1924 135
rect 1918 130 1924 131
rect 2038 135 2044 136
rect 2038 131 2039 135
rect 2043 131 2044 135
rect 2038 130 2044 131
rect 2158 135 2164 136
rect 2158 131 2159 135
rect 2163 131 2164 135
rect 2158 130 2164 131
rect 2240 128 2242 222
rect 2272 212 2274 230
rect 2324 212 2326 238
rect 2351 237 2355 238
rect 2447 242 2451 243
rect 2447 237 2451 238
rect 2511 242 2515 243
rect 2511 237 2515 238
rect 2599 242 2603 243
rect 2599 237 2603 238
rect 2352 221 2354 237
rect 2512 221 2514 237
rect 2672 236 2674 270
rect 2680 252 2682 342
rect 2758 337 2764 338
rect 2758 333 2759 337
rect 2763 333 2764 337
rect 2758 332 2764 333
rect 2910 337 2916 338
rect 2910 333 2911 337
rect 2915 333 2916 337
rect 2910 332 2916 333
rect 3062 337 3068 338
rect 3062 333 3063 337
rect 3067 333 3068 337
rect 3062 332 3068 333
rect 2760 311 2762 332
rect 2912 311 2914 332
rect 3064 311 3066 332
rect 2759 310 2763 311
rect 2759 305 2763 306
rect 2911 310 2915 311
rect 2911 305 2915 306
rect 2919 310 2923 311
rect 2919 305 2923 306
rect 3063 310 3067 311
rect 3063 305 3067 306
rect 3087 310 3091 311
rect 3087 305 3091 306
rect 2760 288 2762 305
rect 2920 288 2922 305
rect 3088 288 3090 305
rect 2758 287 2764 288
rect 2758 283 2759 287
rect 2763 283 2764 287
rect 2758 282 2764 283
rect 2918 287 2924 288
rect 2918 283 2919 287
rect 2923 283 2924 287
rect 2918 282 2924 283
rect 3086 287 3092 288
rect 3086 283 3087 287
rect 3091 283 3092 287
rect 3086 282 3092 283
rect 3168 280 3170 366
rect 3224 357 3226 373
rect 3222 356 3228 357
rect 3222 352 3223 356
rect 3227 352 3228 356
rect 3222 351 3228 352
rect 3222 337 3228 338
rect 3222 333 3223 337
rect 3227 333 3228 337
rect 3222 332 3228 333
rect 3224 311 3226 332
rect 3223 310 3227 311
rect 3223 305 3227 306
rect 3255 310 3259 311
rect 3255 305 3259 306
rect 3256 288 3258 305
rect 3254 287 3260 288
rect 3254 283 3255 287
rect 3259 283 3260 287
rect 3254 282 3260 283
rect 3166 279 3172 280
rect 2830 275 2836 276
rect 2830 271 2831 275
rect 2835 271 2836 275
rect 2830 270 2836 271
rect 2990 275 2996 276
rect 2990 271 2991 275
rect 2995 271 2996 275
rect 3166 275 3167 279
rect 3171 275 3172 279
rect 3166 274 3172 275
rect 2990 270 2996 271
rect 2758 268 2764 269
rect 2758 264 2759 268
rect 2763 264 2764 268
rect 2758 263 2764 264
rect 2678 251 2684 252
rect 2678 247 2679 251
rect 2683 247 2684 251
rect 2678 246 2684 247
rect 2760 243 2762 263
rect 2832 252 2834 270
rect 2918 268 2924 269
rect 2918 264 2919 268
rect 2923 264 2924 268
rect 2918 263 2924 264
rect 2814 251 2820 252
rect 2814 247 2815 251
rect 2819 247 2820 251
rect 2814 246 2820 247
rect 2830 251 2836 252
rect 2830 247 2831 251
rect 2835 247 2836 251
rect 2830 246 2836 247
rect 2679 242 2683 243
rect 2679 237 2683 238
rect 2759 242 2763 243
rect 2759 237 2763 238
rect 2590 235 2596 236
rect 2590 231 2591 235
rect 2595 231 2596 235
rect 2590 230 2596 231
rect 2670 235 2676 236
rect 2670 231 2671 235
rect 2675 231 2676 235
rect 2670 230 2676 231
rect 2350 220 2356 221
rect 2350 216 2351 220
rect 2355 216 2356 220
rect 2350 215 2356 216
rect 2510 220 2516 221
rect 2510 216 2511 220
rect 2515 216 2516 220
rect 2510 215 2516 216
rect 2592 212 2594 230
rect 2680 221 2682 237
rect 2678 220 2684 221
rect 2678 216 2679 220
rect 2683 216 2684 220
rect 2678 215 2684 216
rect 2816 212 2818 246
rect 2920 243 2922 263
rect 2992 252 2994 270
rect 3086 268 3092 269
rect 3086 264 3087 268
rect 3091 264 3092 268
rect 3086 263 3092 264
rect 3254 268 3260 269
rect 3254 264 3255 268
rect 3259 264 3260 268
rect 3254 263 3260 264
rect 2990 251 2996 252
rect 2990 247 2991 251
rect 2995 247 2996 251
rect 2990 246 2996 247
rect 3088 243 3090 263
rect 3256 243 3258 263
rect 3336 252 3338 406
rect 3366 404 3372 405
rect 3366 400 3367 404
rect 3371 400 3372 404
rect 3462 403 3463 407
rect 3467 403 3468 407
rect 3462 402 3468 403
rect 3366 399 3372 400
rect 3368 379 3370 399
rect 3430 387 3436 388
rect 3430 383 3431 387
rect 3435 383 3436 387
rect 3430 382 3436 383
rect 3367 378 3371 379
rect 3367 373 3371 374
rect 3368 357 3370 373
rect 3366 356 3372 357
rect 3366 352 3367 356
rect 3371 352 3372 356
rect 3366 351 3372 352
rect 3432 348 3434 382
rect 3464 379 3466 402
rect 3463 378 3467 379
rect 3463 373 3467 374
rect 3438 371 3444 372
rect 3438 367 3439 371
rect 3443 367 3444 371
rect 3438 366 3444 367
rect 3430 347 3436 348
rect 3430 343 3431 347
rect 3435 343 3436 347
rect 3430 342 3436 343
rect 3366 337 3372 338
rect 3366 333 3367 337
rect 3371 333 3372 337
rect 3366 332 3372 333
rect 3368 311 3370 332
rect 3367 310 3371 311
rect 3367 305 3371 306
rect 3334 251 3340 252
rect 3334 247 3335 251
rect 3339 247 3340 251
rect 3334 246 3340 247
rect 2847 242 2851 243
rect 2847 237 2851 238
rect 2919 242 2923 243
rect 2919 237 2923 238
rect 3023 242 3027 243
rect 3023 237 3027 238
rect 3087 242 3091 243
rect 3087 237 3091 238
rect 3207 242 3211 243
rect 3207 237 3211 238
rect 3255 242 3259 243
rect 3255 237 3259 238
rect 3367 242 3371 243
rect 3367 237 3371 238
rect 2848 221 2850 237
rect 2926 235 2932 236
rect 2926 231 2927 235
rect 2931 231 2932 235
rect 2926 230 2932 231
rect 2846 220 2852 221
rect 2846 216 2847 220
rect 2851 216 2852 220
rect 2846 215 2852 216
rect 2928 212 2930 230
rect 3024 221 3026 237
rect 3126 235 3132 236
rect 3126 231 3127 235
rect 3131 231 3132 235
rect 3126 230 3132 231
rect 3022 220 3028 221
rect 3022 216 3023 220
rect 3027 216 3028 220
rect 3022 215 3028 216
rect 2270 211 2276 212
rect 2270 207 2271 211
rect 2275 207 2276 211
rect 2270 206 2276 207
rect 2322 211 2328 212
rect 2322 207 2323 211
rect 2327 207 2328 211
rect 2322 206 2328 207
rect 2454 211 2460 212
rect 2454 207 2455 211
rect 2459 207 2460 211
rect 2454 206 2460 207
rect 2590 211 2596 212
rect 2590 207 2591 211
rect 2595 207 2596 211
rect 2590 206 2596 207
rect 2814 211 2820 212
rect 2814 207 2815 211
rect 2819 207 2820 211
rect 2814 206 2820 207
rect 2926 211 2932 212
rect 2926 207 2927 211
rect 2931 207 2932 211
rect 2926 206 2932 207
rect 2350 201 2356 202
rect 2350 197 2351 201
rect 2355 197 2356 201
rect 2350 196 2356 197
rect 2352 159 2354 196
rect 2279 158 2283 159
rect 2279 153 2283 154
rect 2351 158 2355 159
rect 2351 153 2355 154
rect 2399 158 2403 159
rect 2399 153 2403 154
rect 2280 136 2282 153
rect 2400 136 2402 153
rect 2278 135 2284 136
rect 2278 131 2279 135
rect 2283 131 2284 135
rect 2278 130 2284 131
rect 2398 135 2404 136
rect 2398 131 2399 135
rect 2403 131 2404 135
rect 2398 130 2404 131
rect 2238 127 2244 128
rect 1902 123 1908 124
rect 1766 120 1772 121
rect 1406 119 1412 120
rect 1406 115 1407 119
rect 1411 115 1412 119
rect 1406 114 1412 115
rect 1494 119 1500 120
rect 1494 115 1495 119
rect 1499 115 1500 119
rect 1494 114 1500 115
rect 1582 119 1588 120
rect 1582 115 1583 119
rect 1587 115 1588 119
rect 1582 114 1588 115
rect 1670 119 1676 120
rect 1670 115 1671 119
rect 1675 115 1676 119
rect 1766 116 1767 120
rect 1771 116 1772 120
rect 1766 115 1772 116
rect 1806 119 1812 120
rect 1806 115 1807 119
rect 1811 115 1812 119
rect 1902 119 1903 123
rect 1907 119 1908 123
rect 1902 118 1908 119
rect 1990 123 1996 124
rect 1990 119 1991 123
rect 1995 119 1996 123
rect 1990 118 1996 119
rect 2110 123 2116 124
rect 2110 119 2111 123
rect 2115 119 2116 123
rect 2110 118 2116 119
rect 2230 123 2236 124
rect 2230 119 2231 123
rect 2235 119 2236 123
rect 2238 123 2239 127
rect 2243 123 2244 127
rect 2238 122 2244 123
rect 2230 118 2236 119
rect 1670 114 1676 115
rect 1806 114 1812 115
rect 1830 116 1836 117
rect 1478 107 1484 108
rect 1478 103 1479 107
rect 1483 103 1484 107
rect 1478 102 1484 103
rect 1566 107 1572 108
rect 1566 103 1567 107
rect 1571 103 1572 107
rect 1566 102 1572 103
rect 1654 107 1660 108
rect 1654 103 1655 107
rect 1659 103 1660 107
rect 1654 102 1660 103
rect 1766 103 1772 104
rect 1406 100 1412 101
rect 1406 96 1407 100
rect 1411 96 1412 100
rect 1406 95 1412 96
rect 1399 92 1403 93
rect 1399 87 1403 88
rect 1382 83 1388 84
rect 1382 79 1383 83
rect 1387 79 1388 83
rect 1408 79 1410 95
rect 1480 84 1482 102
rect 1494 100 1500 101
rect 1494 96 1495 100
rect 1499 96 1500 100
rect 1494 95 1500 96
rect 1478 83 1484 84
rect 1478 79 1479 83
rect 1483 79 1484 83
rect 1496 79 1498 95
rect 1568 84 1570 102
rect 1582 100 1588 101
rect 1582 96 1583 100
rect 1587 96 1588 100
rect 1582 95 1588 96
rect 1566 83 1572 84
rect 1566 79 1567 83
rect 1571 79 1572 83
rect 1584 79 1586 95
rect 1656 84 1658 102
rect 1670 100 1676 101
rect 1670 96 1671 100
rect 1675 96 1676 100
rect 1766 99 1767 103
rect 1771 99 1772 103
rect 1766 98 1772 99
rect 1670 95 1676 96
rect 1654 83 1660 84
rect 1654 79 1655 83
rect 1659 79 1660 83
rect 1672 79 1674 95
rect 1768 79 1770 98
rect 1808 95 1810 114
rect 1830 112 1831 116
rect 1835 112 1836 116
rect 1830 111 1836 112
rect 1832 95 1834 111
rect 1904 100 1906 118
rect 1918 116 1924 117
rect 1918 112 1919 116
rect 1923 112 1924 116
rect 1918 111 1924 112
rect 1902 99 1908 100
rect 1902 95 1903 99
rect 1907 95 1908 99
rect 1920 95 1922 111
rect 1992 100 1994 118
rect 2038 116 2044 117
rect 2038 112 2039 116
rect 2043 112 2044 116
rect 2038 111 2044 112
rect 1990 99 1996 100
rect 1990 95 1991 99
rect 1995 95 1996 99
rect 2040 95 2042 111
rect 2112 100 2114 118
rect 2158 116 2164 117
rect 2158 112 2159 116
rect 2163 112 2164 116
rect 2158 111 2164 112
rect 2110 99 2116 100
rect 2110 95 2111 99
rect 2115 95 2116 99
rect 2160 95 2162 111
rect 2232 100 2234 118
rect 2278 116 2284 117
rect 2278 112 2279 116
rect 2283 112 2284 116
rect 2278 111 2284 112
rect 2398 116 2404 117
rect 2398 112 2399 116
rect 2403 112 2404 116
rect 2398 111 2404 112
rect 2230 99 2236 100
rect 2230 95 2231 99
rect 2235 95 2236 99
rect 2280 95 2282 111
rect 2400 95 2402 111
rect 2456 100 2458 206
rect 2510 201 2516 202
rect 2510 197 2511 201
rect 2515 197 2516 201
rect 2510 196 2516 197
rect 2678 201 2684 202
rect 2678 197 2679 201
rect 2683 197 2684 201
rect 2678 196 2684 197
rect 2846 201 2852 202
rect 2846 197 2847 201
rect 2851 197 2852 201
rect 2846 196 2852 197
rect 3022 201 3028 202
rect 3022 197 3023 201
rect 3027 197 3028 201
rect 3022 196 3028 197
rect 2512 159 2514 196
rect 2680 159 2682 196
rect 2848 159 2850 196
rect 3024 159 3026 196
rect 2511 158 2515 159
rect 2511 153 2515 154
rect 2623 158 2627 159
rect 2623 153 2627 154
rect 2679 158 2683 159
rect 2679 153 2683 154
rect 2735 158 2739 159
rect 2735 153 2739 154
rect 2839 158 2843 159
rect 2839 153 2843 154
rect 2847 158 2851 159
rect 2847 153 2851 154
rect 2943 158 2947 159
rect 2943 153 2947 154
rect 3023 158 3027 159
rect 3023 153 3027 154
rect 3055 158 3059 159
rect 3055 153 3059 154
rect 2512 136 2514 153
rect 2624 136 2626 153
rect 2736 136 2738 153
rect 2840 136 2842 153
rect 2944 136 2946 153
rect 3056 136 3058 153
rect 2510 135 2516 136
rect 2510 131 2511 135
rect 2515 131 2516 135
rect 2510 130 2516 131
rect 2622 135 2628 136
rect 2622 131 2623 135
rect 2627 131 2628 135
rect 2622 130 2628 131
rect 2734 135 2740 136
rect 2734 131 2735 135
rect 2739 131 2740 135
rect 2734 130 2740 131
rect 2838 135 2844 136
rect 2838 131 2839 135
rect 2843 131 2844 135
rect 2838 130 2844 131
rect 2942 135 2948 136
rect 2942 131 2943 135
rect 2947 131 2948 135
rect 2942 130 2948 131
rect 3054 135 3060 136
rect 3054 131 3055 135
rect 3059 131 3060 135
rect 3054 130 3060 131
rect 3128 128 3130 230
rect 3208 221 3210 237
rect 3368 221 3370 237
rect 3430 235 3436 236
rect 3430 231 3431 235
rect 3435 231 3436 235
rect 3430 230 3436 231
rect 3206 220 3212 221
rect 3206 216 3207 220
rect 3211 216 3212 220
rect 3206 215 3212 216
rect 3366 220 3372 221
rect 3366 216 3367 220
rect 3371 216 3372 220
rect 3366 215 3372 216
rect 3270 211 3276 212
rect 3270 207 3271 211
rect 3275 207 3276 211
rect 3270 206 3276 207
rect 3206 201 3212 202
rect 3206 197 3207 201
rect 3211 197 3212 201
rect 3206 196 3212 197
rect 3208 159 3210 196
rect 3167 158 3171 159
rect 3167 153 3171 154
rect 3207 158 3211 159
rect 3207 153 3211 154
rect 3168 136 3170 153
rect 3166 135 3172 136
rect 3166 131 3167 135
rect 3171 131 3172 135
rect 3166 130 3172 131
rect 3126 127 3132 128
rect 2470 123 2476 124
rect 2470 119 2471 123
rect 2475 119 2476 123
rect 2470 118 2476 119
rect 2582 123 2588 124
rect 2582 119 2583 123
rect 2587 119 2588 123
rect 2582 118 2588 119
rect 2694 123 2700 124
rect 2694 119 2695 123
rect 2699 119 2700 123
rect 2694 118 2700 119
rect 2806 123 2812 124
rect 2806 119 2807 123
rect 2811 119 2812 123
rect 2806 118 2812 119
rect 2910 123 2916 124
rect 2910 119 2911 123
rect 2915 119 2916 123
rect 2910 118 2916 119
rect 3014 123 3020 124
rect 3014 119 3015 123
rect 3019 119 3020 123
rect 3126 123 3127 127
rect 3131 123 3132 127
rect 3126 122 3132 123
rect 3014 118 3020 119
rect 2472 100 2474 118
rect 2510 116 2516 117
rect 2510 112 2511 116
rect 2515 112 2516 116
rect 2510 111 2516 112
rect 2454 99 2460 100
rect 2454 95 2455 99
rect 2459 95 2460 99
rect 1807 94 1811 95
rect 1807 89 1811 90
rect 1831 94 1835 95
rect 1902 94 1908 95
rect 1919 94 1923 95
rect 1990 94 1996 95
rect 2039 94 2043 95
rect 2110 94 2116 95
rect 2159 94 2163 95
rect 2230 94 2236 95
rect 2279 94 2283 95
rect 1831 89 1835 90
rect 1919 89 1923 90
rect 2039 89 2043 90
rect 2159 89 2163 90
rect 2279 89 2283 90
rect 2399 94 2403 95
rect 2454 94 2460 95
rect 2470 99 2476 100
rect 2470 95 2471 99
rect 2475 95 2476 99
rect 2512 95 2514 111
rect 2584 100 2586 118
rect 2622 116 2628 117
rect 2622 112 2623 116
rect 2627 112 2628 116
rect 2622 111 2628 112
rect 2582 99 2588 100
rect 2582 95 2583 99
rect 2587 95 2588 99
rect 2624 95 2626 111
rect 2696 100 2698 118
rect 2734 116 2740 117
rect 2734 112 2735 116
rect 2739 112 2740 116
rect 2734 111 2740 112
rect 2694 99 2700 100
rect 2694 95 2695 99
rect 2699 95 2700 99
rect 2736 95 2738 111
rect 2808 100 2810 118
rect 2838 116 2844 117
rect 2838 112 2839 116
rect 2843 112 2844 116
rect 2838 111 2844 112
rect 2806 99 2812 100
rect 2806 95 2807 99
rect 2811 95 2812 99
rect 2840 95 2842 111
rect 2912 100 2914 118
rect 2942 116 2948 117
rect 2942 112 2943 116
rect 2947 112 2948 116
rect 2942 111 2948 112
rect 2910 99 2916 100
rect 2910 95 2911 99
rect 2915 95 2916 99
rect 2944 95 2946 111
rect 3016 100 3018 118
rect 3054 116 3060 117
rect 3054 112 3055 116
rect 3059 112 3060 116
rect 3054 111 3060 112
rect 3166 116 3172 117
rect 3166 112 3167 116
rect 3171 112 3172 116
rect 3166 111 3172 112
rect 3014 99 3020 100
rect 3014 95 3015 99
rect 3019 95 3020 99
rect 3056 95 3058 111
rect 3168 95 3170 111
rect 3272 100 3274 206
rect 3366 201 3372 202
rect 3366 197 3367 201
rect 3371 197 3372 201
rect 3366 196 3372 197
rect 3368 159 3370 196
rect 3279 158 3283 159
rect 3279 153 3283 154
rect 3367 158 3371 159
rect 3367 153 3371 154
rect 3280 136 3282 153
rect 3368 136 3370 153
rect 3278 135 3284 136
rect 3278 131 3279 135
rect 3283 131 3284 135
rect 3278 130 3284 131
rect 3366 135 3372 136
rect 3366 131 3367 135
rect 3371 131 3372 135
rect 3432 132 3434 230
rect 3440 212 3442 366
rect 3464 354 3466 373
rect 3462 353 3468 354
rect 3462 349 3463 353
rect 3467 349 3468 353
rect 3462 348 3468 349
rect 3462 336 3468 337
rect 3462 332 3463 336
rect 3467 332 3468 336
rect 3462 331 3468 332
rect 3464 311 3466 331
rect 3463 310 3467 311
rect 3463 305 3467 306
rect 3464 289 3466 305
rect 3462 288 3468 289
rect 3462 284 3463 288
rect 3467 284 3468 288
rect 3462 283 3468 284
rect 3462 271 3468 272
rect 3462 267 3463 271
rect 3467 267 3468 271
rect 3462 266 3468 267
rect 3464 243 3466 266
rect 3463 242 3467 243
rect 3463 237 3467 238
rect 3464 218 3466 237
rect 3462 217 3468 218
rect 3462 213 3463 217
rect 3467 213 3468 217
rect 3462 212 3468 213
rect 3438 211 3444 212
rect 3438 207 3439 211
rect 3443 207 3444 211
rect 3438 206 3444 207
rect 3462 200 3468 201
rect 3462 196 3463 200
rect 3467 196 3468 200
rect 3462 195 3468 196
rect 3464 159 3466 195
rect 3463 158 3467 159
rect 3463 153 3467 154
rect 3464 137 3466 153
rect 3462 136 3468 137
rect 3462 132 3463 136
rect 3467 132 3468 136
rect 3366 130 3372 131
rect 3430 131 3436 132
rect 3462 131 3468 132
rect 3430 127 3431 131
rect 3435 127 3436 131
rect 3430 126 3436 127
rect 3350 123 3356 124
rect 3350 119 3351 123
rect 3355 119 3356 123
rect 3350 118 3356 119
rect 3462 119 3468 120
rect 3278 116 3284 117
rect 3278 112 3279 116
rect 3283 112 3284 116
rect 3278 111 3284 112
rect 3270 99 3276 100
rect 3270 95 3271 99
rect 3275 95 3276 99
rect 3280 95 3282 111
rect 3352 100 3354 118
rect 3366 116 3372 117
rect 3366 112 3367 116
rect 3371 112 3372 116
rect 3462 115 3463 119
rect 3467 115 3468 119
rect 3462 114 3468 115
rect 3366 111 3372 112
rect 3350 99 3356 100
rect 3350 95 3351 99
rect 3355 95 3356 99
rect 3368 95 3370 111
rect 3464 95 3466 114
rect 2470 94 2476 95
rect 2511 94 2515 95
rect 2582 94 2588 95
rect 2623 94 2627 95
rect 2694 94 2700 95
rect 2735 94 2739 95
rect 2806 94 2812 95
rect 2839 94 2843 95
rect 2910 94 2916 95
rect 2943 94 2947 95
rect 3014 94 3020 95
rect 3055 94 3059 95
rect 2399 89 2403 90
rect 2511 89 2515 90
rect 2623 89 2627 90
rect 2735 89 2739 90
rect 2839 89 2843 90
rect 2943 89 2947 90
rect 3055 89 3059 90
rect 3167 94 3171 95
rect 3270 94 3276 95
rect 3279 94 3283 95
rect 3350 94 3356 95
rect 3367 94 3371 95
rect 3167 89 3171 90
rect 3279 89 3283 90
rect 3367 89 3371 90
rect 3463 94 3467 95
rect 3463 89 3467 90
rect 918 78 924 79
rect 943 78 947 79
rect 1014 78 1020 79
rect 1031 78 1035 79
rect 1102 78 1108 79
rect 1119 78 1123 79
rect 1190 78 1196 79
rect 1215 78 1219 79
rect 1286 78 1292 79
rect 1311 78 1315 79
rect 1382 78 1388 79
rect 1407 78 1411 79
rect 1478 78 1484 79
rect 1495 78 1499 79
rect 1566 78 1572 79
rect 1583 78 1587 79
rect 1654 78 1660 79
rect 1671 78 1675 79
rect 847 73 851 74
rect 943 73 947 74
rect 1031 73 1035 74
rect 1119 73 1123 74
rect 1215 73 1219 74
rect 1311 73 1315 74
rect 1407 73 1411 74
rect 1495 73 1499 74
rect 1583 73 1587 74
rect 1671 73 1675 74
rect 1767 78 1771 79
rect 1767 73 1771 74
<< m4c >>
rect 1807 3518 1811 3522
rect 2007 3518 2011 3522
rect 2239 3518 2243 3522
rect 2455 3518 2459 3522
rect 2655 3518 2659 3522
rect 2855 3518 2859 3522
rect 3047 3518 3051 3522
rect 3247 3518 3251 3522
rect 3463 3518 3467 3522
rect 111 3482 115 3486
rect 455 3482 459 3486
rect 543 3482 547 3486
rect 631 3482 635 3486
rect 719 3482 723 3486
rect 807 3482 811 3486
rect 895 3482 899 3486
rect 983 3482 987 3486
rect 1071 3482 1075 3486
rect 1159 3482 1163 3486
rect 1767 3482 1771 3486
rect 111 3418 115 3422
rect 415 3418 419 3422
rect 455 3418 459 3422
rect 503 3418 507 3422
rect 543 3418 547 3422
rect 591 3418 595 3422
rect 1807 3454 1811 3458
rect 1831 3454 1835 3458
rect 1943 3454 1947 3458
rect 2007 3454 2011 3458
rect 2079 3454 2083 3458
rect 2215 3454 2219 3458
rect 2239 3454 2243 3458
rect 2351 3454 2355 3458
rect 631 3418 635 3422
rect 679 3418 683 3422
rect 719 3418 723 3422
rect 767 3418 771 3422
rect 807 3418 811 3422
rect 855 3418 859 3422
rect 895 3418 899 3422
rect 943 3418 947 3422
rect 983 3418 987 3422
rect 1031 3418 1035 3422
rect 1071 3418 1075 3422
rect 1119 3418 1123 3422
rect 1159 3418 1163 3422
rect 1207 3418 1211 3422
rect 1303 3418 1307 3422
rect 1767 3418 1771 3422
rect 111 3350 115 3354
rect 399 3350 403 3354
rect 415 3350 419 3354
rect 495 3350 499 3354
rect 503 3350 507 3354
rect 591 3350 595 3354
rect 599 3350 603 3354
rect 679 3350 683 3354
rect 703 3350 707 3354
rect 767 3350 771 3354
rect 807 3350 811 3354
rect 855 3350 859 3354
rect 911 3350 915 3354
rect 943 3350 947 3354
rect 1015 3350 1019 3354
rect 1031 3350 1035 3354
rect 1119 3350 1123 3354
rect 1207 3350 1211 3354
rect 1223 3350 1227 3354
rect 1807 3382 1811 3386
rect 1831 3382 1835 3386
rect 1943 3382 1947 3386
rect 1951 3382 1955 3386
rect 2079 3382 2083 3386
rect 2095 3382 2099 3386
rect 2455 3454 2459 3458
rect 2479 3454 2483 3458
rect 2599 3454 2603 3458
rect 2655 3454 2659 3458
rect 2719 3454 2723 3458
rect 2847 3454 2851 3458
rect 2855 3454 2859 3458
rect 2975 3454 2979 3458
rect 3047 3454 3051 3458
rect 3247 3454 3251 3458
rect 3463 3454 3467 3458
rect 2215 3382 2219 3386
rect 2239 3382 2243 3386
rect 1303 3350 1307 3354
rect 1327 3350 1331 3354
rect 1767 3350 1771 3354
rect 111 3282 115 3286
rect 383 3282 387 3286
rect 399 3282 403 3286
rect 495 3282 499 3286
rect 599 3282 603 3286
rect 607 3282 611 3286
rect 703 3282 707 3286
rect 727 3282 731 3286
rect 807 3282 811 3286
rect 847 3282 851 3286
rect 1807 3310 1811 3314
rect 911 3282 915 3286
rect 967 3282 971 3286
rect 1015 3282 1019 3286
rect 1087 3282 1091 3286
rect 1119 3282 1123 3286
rect 1207 3282 1211 3286
rect 1223 3282 1227 3286
rect 1327 3282 1331 3286
rect 1335 3282 1339 3286
rect 111 3214 115 3218
rect 303 3214 307 3218
rect 383 3214 387 3218
rect 423 3214 427 3218
rect 495 3214 499 3218
rect 543 3214 547 3218
rect 111 3138 115 3142
rect 175 3138 179 3142
rect 303 3138 307 3142
rect 319 3138 323 3142
rect 423 3138 427 3142
rect 471 3138 475 3142
rect 607 3214 611 3218
rect 671 3214 675 3218
rect 727 3214 731 3218
rect 799 3214 803 3218
rect 847 3214 851 3218
rect 927 3214 931 3218
rect 967 3214 971 3218
rect 1831 3310 1835 3314
rect 1767 3282 1771 3286
rect 2351 3382 2355 3386
rect 2383 3382 2387 3386
rect 2479 3382 2483 3386
rect 2519 3382 2523 3386
rect 2599 3382 2603 3386
rect 2647 3382 2651 3386
rect 2719 3382 2723 3386
rect 2775 3382 2779 3386
rect 2847 3382 2851 3386
rect 2903 3382 2907 3386
rect 2975 3382 2979 3386
rect 3039 3382 3043 3386
rect 3463 3382 3467 3386
rect 1951 3310 1955 3314
rect 1975 3310 1979 3314
rect 2095 3310 2099 3314
rect 2151 3310 2155 3314
rect 2239 3310 2243 3314
rect 2335 3310 2339 3314
rect 2383 3310 2387 3314
rect 1807 3238 1811 3242
rect 1831 3238 1835 3242
rect 1975 3238 1979 3242
rect 2031 3238 2035 3242
rect 1055 3214 1059 3218
rect 1087 3214 1091 3218
rect 1175 3214 1179 3218
rect 1207 3214 1211 3218
rect 1303 3214 1307 3218
rect 1335 3214 1339 3218
rect 1431 3214 1435 3218
rect 1767 3214 1771 3218
rect 2511 3310 2515 3314
rect 2519 3310 2523 3314
rect 2647 3310 2651 3314
rect 2679 3310 2683 3314
rect 2775 3310 2779 3314
rect 2831 3310 2835 3314
rect 2903 3310 2907 3314
rect 2975 3310 2979 3314
rect 3039 3310 3043 3314
rect 3111 3310 3115 3314
rect 3247 3310 3251 3314
rect 3367 3310 3371 3314
rect 3463 3310 3467 3314
rect 2151 3238 2155 3242
rect 2247 3238 2251 3242
rect 543 3138 547 3142
rect 623 3138 627 3142
rect 671 3138 675 3142
rect 775 3138 779 3142
rect 799 3138 803 3142
rect 919 3138 923 3142
rect 927 3138 931 3142
rect 1055 3138 1059 3142
rect 1063 3138 1067 3142
rect 1175 3138 1179 3142
rect 1199 3138 1203 3142
rect 2335 3238 2339 3242
rect 2455 3238 2459 3242
rect 2511 3238 2515 3242
rect 2655 3238 2659 3242
rect 2679 3238 2683 3242
rect 2831 3238 2835 3242
rect 2839 3238 2843 3242
rect 2975 3238 2979 3242
rect 3023 3238 3027 3242
rect 3111 3238 3115 3242
rect 3207 3238 3211 3242
rect 3247 3238 3251 3242
rect 3367 3238 3371 3242
rect 3463 3238 3467 3242
rect 1807 3174 1811 3178
rect 1831 3174 1835 3178
rect 1839 3174 1843 3178
rect 2031 3174 2035 3178
rect 2223 3174 2227 3178
rect 2247 3174 2251 3178
rect 2407 3174 2411 3178
rect 2455 3174 2459 3178
rect 2575 3174 2579 3178
rect 1303 3138 1307 3142
rect 1343 3138 1347 3142
rect 1431 3138 1435 3142
rect 1487 3138 1491 3142
rect 1767 3138 1771 3142
rect 111 3066 115 3070
rect 135 3066 139 3070
rect 175 3066 179 3070
rect 263 3066 267 3070
rect 319 3066 323 3070
rect 111 2998 115 3002
rect 135 2998 139 3002
rect 263 2998 267 3002
rect 327 2998 331 3002
rect 431 3066 435 3070
rect 471 3066 475 3070
rect 607 3066 611 3070
rect 623 3066 627 3070
rect 775 3066 779 3070
rect 791 3066 795 3070
rect 919 3066 923 3070
rect 967 3066 971 3070
rect 1063 3066 1067 3070
rect 1143 3066 1147 3070
rect 1199 3066 1203 3070
rect 1327 3066 1331 3070
rect 1343 3066 1347 3070
rect 1487 3066 1491 3070
rect 1511 3066 1515 3070
rect 1807 3106 1811 3110
rect 1839 3106 1843 3110
rect 1935 3106 1939 3110
rect 2031 3106 2035 3110
rect 2055 3106 2059 3110
rect 2175 3106 2179 3110
rect 2223 3106 2227 3110
rect 2655 3174 2659 3178
rect 2735 3174 2739 3178
rect 2839 3174 2843 3178
rect 2879 3174 2883 3178
rect 3007 3174 3011 3178
rect 3023 3174 3027 3178
rect 2303 3106 2307 3110
rect 2407 3106 2411 3110
rect 2431 3106 2435 3110
rect 1767 3066 1771 3070
rect 1807 3034 1811 3038
rect 1935 3034 1939 3038
rect 431 2998 435 3002
rect 535 2998 539 3002
rect 607 2998 611 3002
rect 735 2998 739 3002
rect 791 2998 795 3002
rect 927 2998 931 3002
rect 967 2998 971 3002
rect 2023 3034 2027 3038
rect 2055 3034 2059 3038
rect 2127 3034 2131 3038
rect 2175 3034 2179 3038
rect 2231 3034 2235 3038
rect 2303 3034 2307 3038
rect 2335 3034 2339 3038
rect 1103 2998 1107 3002
rect 1143 2998 1147 3002
rect 1279 2998 1283 3002
rect 1327 2998 1331 3002
rect 1447 2998 1451 3002
rect 1511 2998 1515 3002
rect 1623 2998 1627 3002
rect 1767 2998 1771 3002
rect 111 2926 115 2930
rect 135 2926 139 2930
rect 263 2926 267 2930
rect 327 2926 331 2930
rect 431 2926 435 2930
rect 535 2926 539 2930
rect 607 2926 611 2930
rect 735 2926 739 2930
rect 783 2926 787 2930
rect 927 2926 931 2930
rect 951 2926 955 2930
rect 1103 2926 1107 2930
rect 1111 2926 1115 2930
rect 1271 2926 1275 2930
rect 1279 2926 1283 2930
rect 1431 2926 1435 2930
rect 1447 2926 1451 2930
rect 1591 2926 1595 2930
rect 1623 2926 1627 2930
rect 1807 2970 1811 2974
rect 2023 2970 2027 2974
rect 2055 2970 2059 2974
rect 2127 2970 2131 2974
rect 2567 3106 2571 3110
rect 2575 3106 2579 3110
rect 2719 3106 2723 3110
rect 2735 3106 2739 3110
rect 2871 3106 2875 3110
rect 2879 3106 2883 3110
rect 3135 3174 3139 3178
rect 3207 3174 3211 3178
rect 3263 3174 3267 3178
rect 3367 3174 3371 3178
rect 3007 3106 3011 3110
rect 3031 3106 3035 3110
rect 3135 3106 3139 3110
rect 3199 3106 3203 3110
rect 3263 3106 3267 3110
rect 3463 3174 3467 3178
rect 3367 3106 3371 3110
rect 3463 3106 3467 3110
rect 2431 3034 2435 3038
rect 2439 3034 2443 3038
rect 2543 3034 2547 3038
rect 2567 3034 2571 3038
rect 2647 3034 2651 3038
rect 2719 3034 2723 3038
rect 2759 3034 2763 3038
rect 2143 2970 2147 2974
rect 2231 2970 2235 2974
rect 2319 2970 2323 2974
rect 2335 2970 2339 2974
rect 1767 2926 1771 2930
rect 1807 2898 1811 2902
rect 2055 2898 2059 2902
rect 2071 2898 2075 2902
rect 2143 2898 2147 2902
rect 2175 2898 2179 2902
rect 2231 2898 2235 2902
rect 111 2858 115 2862
rect 135 2858 139 2862
rect 255 2858 259 2862
rect 263 2858 267 2862
rect 407 2858 411 2862
rect 431 2858 435 2862
rect 567 2858 571 2862
rect 607 2858 611 2862
rect 727 2858 731 2862
rect 783 2858 787 2862
rect 879 2858 883 2862
rect 951 2858 955 2862
rect 1023 2858 1027 2862
rect 1111 2858 1115 2862
rect 1167 2858 1171 2862
rect 1271 2858 1275 2862
rect 1311 2858 1315 2862
rect 1431 2858 1435 2862
rect 111 2786 115 2790
rect 135 2786 139 2790
rect 255 2786 259 2790
rect 287 2786 291 2790
rect 391 2786 395 2790
rect 407 2786 411 2790
rect 503 2786 507 2790
rect 567 2786 571 2790
rect 623 2786 627 2790
rect 727 2786 731 2790
rect 743 2786 747 2790
rect 855 2786 859 2790
rect 879 2786 883 2790
rect 967 2786 971 2790
rect 1023 2786 1027 2790
rect 1079 2786 1083 2790
rect 1167 2786 1171 2790
rect 1199 2786 1203 2790
rect 1463 2858 1467 2862
rect 1591 2858 1595 2862
rect 1767 2858 1771 2862
rect 1807 2830 1811 2834
rect 1983 2830 1987 2834
rect 2271 2898 2275 2902
rect 2319 2898 2323 2902
rect 2367 2898 2371 2902
rect 2407 2970 2411 2974
rect 2439 2970 2443 2974
rect 2495 2970 2499 2974
rect 2543 2970 2547 2974
rect 2583 2970 2587 2974
rect 2647 2970 2651 2974
rect 2871 3034 2875 3038
rect 3031 3034 3035 3038
rect 3199 3034 3203 3038
rect 3367 3034 3371 3038
rect 3463 3034 3467 3038
rect 2671 2970 2675 2974
rect 2759 2970 2763 2974
rect 2847 2970 2851 2974
rect 3463 2970 3467 2974
rect 2407 2898 2411 2902
rect 2471 2898 2475 2902
rect 2495 2898 2499 2902
rect 2575 2898 2579 2902
rect 2583 2898 2587 2902
rect 2671 2898 2675 2902
rect 2679 2898 2683 2902
rect 2759 2898 2763 2902
rect 2783 2898 2787 2902
rect 2847 2898 2851 2902
rect 2071 2830 2075 2834
rect 2111 2830 2115 2834
rect 2175 2830 2179 2834
rect 2239 2830 2243 2834
rect 2271 2830 2275 2834
rect 2367 2830 2371 2834
rect 1311 2786 1315 2790
rect 1319 2786 1323 2790
rect 1463 2786 1467 2790
rect 1767 2786 1771 2790
rect 1807 2762 1811 2766
rect 1887 2762 1891 2766
rect 1983 2762 1987 2766
rect 2031 2762 2035 2766
rect 2111 2762 2115 2766
rect 2183 2762 2187 2766
rect 2239 2762 2243 2766
rect 111 2718 115 2722
rect 287 2718 291 2722
rect 391 2718 395 2722
rect 479 2718 483 2722
rect 503 2718 507 2722
rect 567 2718 571 2722
rect 623 2718 627 2722
rect 655 2718 659 2722
rect 743 2718 747 2722
rect 831 2718 835 2722
rect 855 2718 859 2722
rect 919 2718 923 2722
rect 967 2718 971 2722
rect 1007 2718 1011 2722
rect 1079 2718 1083 2722
rect 1095 2718 1099 2722
rect 1183 2718 1187 2722
rect 111 2646 115 2650
rect 471 2646 475 2650
rect 479 2646 483 2650
rect 559 2646 563 2650
rect 567 2646 571 2650
rect 647 2646 651 2650
rect 655 2646 659 2650
rect 735 2646 739 2650
rect 743 2646 747 2650
rect 823 2646 827 2650
rect 831 2646 835 2650
rect 111 2570 115 2574
rect 223 2570 227 2574
rect 311 2570 315 2574
rect 407 2570 411 2574
rect 471 2570 475 2574
rect 503 2570 507 2574
rect 911 2646 915 2650
rect 919 2646 923 2650
rect 999 2646 1003 2650
rect 1007 2646 1011 2650
rect 1199 2718 1203 2722
rect 1319 2718 1323 2722
rect 1767 2718 1771 2722
rect 1807 2698 1811 2702
rect 1831 2698 1835 2702
rect 1887 2698 1891 2702
rect 2471 2830 2475 2834
rect 2487 2830 2491 2834
rect 3463 2898 3467 2902
rect 2575 2830 2579 2834
rect 2607 2830 2611 2834
rect 2679 2830 2683 2834
rect 2719 2830 2723 2834
rect 2783 2830 2787 2834
rect 2839 2830 2843 2834
rect 2959 2830 2963 2834
rect 3463 2830 3467 2834
rect 2335 2762 2339 2766
rect 2367 2762 2371 2766
rect 2479 2762 2483 2766
rect 2487 2762 2491 2766
rect 2607 2762 2611 2766
rect 2623 2762 2627 2766
rect 2719 2762 2723 2766
rect 2767 2762 2771 2766
rect 2839 2762 2843 2766
rect 2911 2762 2915 2766
rect 2959 2762 2963 2766
rect 3055 2762 3059 2766
rect 3463 2762 3467 2766
rect 2023 2698 2027 2702
rect 2031 2698 2035 2702
rect 2183 2698 2187 2702
rect 2231 2698 2235 2702
rect 2335 2698 2339 2702
rect 2431 2698 2435 2702
rect 2479 2698 2483 2702
rect 1087 2646 1091 2650
rect 1095 2646 1099 2650
rect 1183 2646 1187 2650
rect 1767 2646 1771 2650
rect 1807 2630 1811 2634
rect 1831 2630 1835 2634
rect 1999 2630 2003 2634
rect 2023 2630 2027 2634
rect 2183 2630 2187 2634
rect 2231 2630 2235 2634
rect 559 2570 563 2574
rect 591 2570 595 2574
rect 647 2570 651 2574
rect 679 2570 683 2574
rect 735 2570 739 2574
rect 767 2570 771 2574
rect 823 2570 827 2574
rect 111 2506 115 2510
rect 135 2506 139 2510
rect 223 2506 227 2510
rect 247 2506 251 2510
rect 311 2506 315 2510
rect 111 2426 115 2430
rect 135 2426 139 2430
rect 391 2506 395 2510
rect 407 2506 411 2510
rect 503 2506 507 2510
rect 543 2506 547 2510
rect 591 2506 595 2510
rect 679 2506 683 2510
rect 695 2506 699 2510
rect 767 2506 771 2510
rect 855 2570 859 2574
rect 911 2570 915 2574
rect 943 2570 947 2574
rect 999 2570 1003 2574
rect 1031 2570 1035 2574
rect 1087 2570 1091 2574
rect 1119 2570 1123 2574
rect 1215 2570 1219 2574
rect 1311 2570 1315 2574
rect 1407 2570 1411 2574
rect 1495 2570 1499 2574
rect 1583 2570 1587 2574
rect 1671 2570 1675 2574
rect 1767 2570 1771 2574
rect 839 2506 843 2510
rect 855 2506 859 2510
rect 943 2506 947 2510
rect 975 2506 979 2510
rect 1031 2506 1035 2510
rect 1103 2506 1107 2510
rect 1119 2506 1123 2510
rect 1215 2506 1219 2510
rect 1231 2506 1235 2510
rect 1311 2506 1315 2510
rect 1351 2506 1355 2510
rect 239 2426 243 2430
rect 247 2426 251 2430
rect 391 2426 395 2430
rect 543 2426 547 2430
rect 551 2426 555 2430
rect 695 2426 699 2430
rect 719 2426 723 2430
rect 839 2426 843 2430
rect 895 2426 899 2430
rect 975 2426 979 2430
rect 111 2354 115 2358
rect 135 2354 139 2358
rect 239 2354 243 2358
rect 375 2354 379 2358
rect 391 2354 395 2358
rect 479 2354 483 2358
rect 551 2354 555 2358
rect 599 2354 603 2358
rect 719 2354 723 2358
rect 847 2354 851 2358
rect 895 2354 899 2358
rect 1063 2426 1067 2430
rect 1103 2426 1107 2430
rect 1231 2426 1235 2430
rect 1239 2426 1243 2430
rect 1407 2506 1411 2510
rect 1463 2506 1467 2510
rect 1495 2506 1499 2510
rect 1575 2506 1579 2510
rect 1583 2506 1587 2510
rect 2359 2630 2363 2634
rect 2615 2698 2619 2702
rect 2623 2698 2627 2702
rect 2767 2698 2771 2702
rect 2783 2698 2787 2702
rect 2911 2698 2915 2702
rect 2943 2698 2947 2702
rect 3055 2698 3059 2702
rect 3095 2698 3099 2702
rect 3239 2698 3243 2702
rect 3367 2698 3371 2702
rect 3463 2698 3467 2702
rect 2431 2630 2435 2634
rect 2519 2630 2523 2634
rect 2615 2630 2619 2634
rect 2671 2630 2675 2634
rect 2783 2630 2787 2634
rect 2807 2630 2811 2634
rect 2927 2630 2931 2634
rect 2943 2630 2947 2634
rect 3047 2630 3051 2634
rect 3095 2630 3099 2634
rect 3159 2630 3163 2634
rect 3239 2630 3243 2634
rect 3271 2630 3275 2634
rect 1807 2558 1811 2562
rect 1831 2558 1835 2562
rect 1999 2558 2003 2562
rect 2183 2558 2187 2562
rect 2207 2558 2211 2562
rect 1671 2506 1675 2510
rect 1767 2506 1771 2510
rect 1807 2478 1811 2482
rect 2015 2478 2019 2482
rect 2359 2558 2363 2562
rect 2519 2558 2523 2562
rect 2671 2558 2675 2562
rect 2799 2558 2803 2562
rect 2807 2558 2811 2562
rect 3367 2630 3371 2634
rect 3463 2630 3467 2634
rect 2927 2558 2931 2562
rect 3047 2558 3051 2562
rect 3159 2558 3163 2562
rect 3271 2558 3275 2562
rect 3367 2558 3371 2562
rect 3463 2558 3467 2562
rect 2199 2478 2203 2482
rect 2207 2478 2211 2482
rect 2367 2478 2371 2482
rect 2527 2478 2531 2482
rect 2671 2478 2675 2482
rect 2799 2478 2803 2482
rect 2807 2478 2811 2482
rect 2927 2478 2931 2482
rect 3047 2478 3051 2482
rect 3159 2478 3163 2482
rect 3271 2478 3275 2482
rect 3367 2478 3371 2482
rect 1351 2426 1355 2430
rect 1415 2426 1419 2430
rect 1463 2426 1467 2430
rect 1575 2426 1579 2430
rect 1591 2426 1595 2430
rect 1671 2426 1675 2430
rect 1767 2426 1771 2430
rect 975 2354 979 2358
rect 1063 2354 1067 2358
rect 1103 2354 1107 2358
rect 1239 2354 1243 2358
rect 1375 2354 1379 2358
rect 1415 2354 1419 2358
rect 1511 2354 1515 2358
rect 1591 2354 1595 2358
rect 1807 2410 1811 2414
rect 1839 2410 1843 2414
rect 2007 2410 2011 2414
rect 2015 2410 2019 2414
rect 2183 2410 2187 2414
rect 2199 2410 2203 2414
rect 2367 2410 2371 2414
rect 1767 2354 1771 2358
rect 1807 2346 1811 2350
rect 1839 2346 1843 2350
rect 1887 2346 1891 2350
rect 2527 2410 2531 2414
rect 2559 2410 2563 2414
rect 3463 2478 3467 2482
rect 2671 2410 2675 2414
rect 2759 2410 2763 2414
rect 2807 2410 2811 2414
rect 2927 2410 2931 2414
rect 2967 2410 2971 2414
rect 3047 2410 3051 2414
rect 3159 2410 3163 2414
rect 3175 2410 3179 2414
rect 3271 2410 3275 2414
rect 3367 2410 3371 2414
rect 3463 2410 3467 2414
rect 2007 2346 2011 2350
rect 2015 2346 2019 2350
rect 2151 2346 2155 2350
rect 2183 2346 2187 2350
rect 2303 2346 2307 2350
rect 2367 2346 2371 2350
rect 2463 2346 2467 2350
rect 2559 2346 2563 2350
rect 2647 2346 2651 2350
rect 2759 2346 2763 2350
rect 2839 2346 2843 2350
rect 2967 2346 2971 2350
rect 3047 2346 3051 2350
rect 3175 2346 3179 2350
rect 3255 2346 3259 2350
rect 3367 2346 3371 2350
rect 111 2282 115 2286
rect 375 2282 379 2286
rect 479 2282 483 2286
rect 575 2282 579 2286
rect 599 2282 603 2286
rect 663 2282 667 2286
rect 719 2282 723 2286
rect 759 2282 763 2286
rect 847 2282 851 2286
rect 863 2282 867 2286
rect 967 2282 971 2286
rect 975 2282 979 2286
rect 1079 2282 1083 2286
rect 1103 2282 1107 2286
rect 111 2218 115 2222
rect 439 2218 443 2222
rect 527 2218 531 2222
rect 575 2218 579 2222
rect 615 2218 619 2222
rect 663 2218 667 2222
rect 703 2218 707 2222
rect 111 2138 115 2142
rect 303 2138 307 2142
rect 407 2138 411 2142
rect 439 2138 443 2142
rect 519 2138 523 2142
rect 527 2138 531 2142
rect 111 2074 115 2078
rect 255 2074 259 2078
rect 303 2074 307 2078
rect 759 2218 763 2222
rect 791 2218 795 2222
rect 1191 2282 1195 2286
rect 1239 2282 1243 2286
rect 1303 2282 1307 2286
rect 1375 2282 1379 2286
rect 1415 2282 1419 2286
rect 1511 2282 1515 2286
rect 1767 2282 1771 2286
rect 1807 2278 1811 2282
rect 1887 2278 1891 2282
rect 2015 2278 2019 2282
rect 2039 2278 2043 2282
rect 2135 2278 2139 2282
rect 2151 2278 2155 2282
rect 863 2218 867 2222
rect 879 2218 883 2222
rect 967 2218 971 2222
rect 1055 2218 1059 2222
rect 1079 2218 1083 2222
rect 1143 2218 1147 2222
rect 1191 2218 1195 2222
rect 1231 2218 1235 2222
rect 1303 2218 1307 2222
rect 1319 2218 1323 2222
rect 1415 2218 1419 2222
rect 1767 2218 1771 2222
rect 2239 2278 2243 2282
rect 2303 2278 2307 2282
rect 2343 2278 2347 2282
rect 2463 2278 2467 2282
rect 2591 2278 2595 2282
rect 2647 2278 2651 2282
rect 2735 2278 2739 2282
rect 2839 2278 2843 2282
rect 2887 2278 2891 2282
rect 3047 2278 3051 2282
rect 3215 2278 3219 2282
rect 3255 2278 3259 2282
rect 1807 2202 1811 2206
rect 2039 2202 2043 2206
rect 2135 2202 2139 2206
rect 2183 2202 2187 2206
rect 2239 2202 2243 2206
rect 2279 2202 2283 2206
rect 2343 2202 2347 2206
rect 2383 2202 2387 2206
rect 2463 2202 2467 2206
rect 2495 2202 2499 2206
rect 2591 2202 2595 2206
rect 2607 2202 2611 2206
rect 2719 2202 2723 2206
rect 2735 2202 2739 2206
rect 2839 2202 2843 2206
rect 2887 2202 2891 2206
rect 2967 2202 2971 2206
rect 3367 2278 3371 2282
rect 3463 2346 3467 2350
rect 3463 2278 3467 2282
rect 3047 2202 3051 2206
rect 3103 2202 3107 2206
rect 3215 2202 3219 2206
rect 3247 2202 3251 2206
rect 615 2138 619 2142
rect 631 2138 635 2142
rect 703 2138 707 2142
rect 743 2138 747 2142
rect 791 2138 795 2142
rect 863 2138 867 2142
rect 879 2138 883 2142
rect 967 2138 971 2142
rect 983 2138 987 2142
rect 1055 2138 1059 2142
rect 1143 2138 1147 2142
rect 1231 2138 1235 2142
rect 1319 2138 1323 2142
rect 1767 2138 1771 2142
rect 375 2074 379 2078
rect 407 2074 411 2078
rect 495 2074 499 2078
rect 519 2074 523 2078
rect 615 2074 619 2078
rect 631 2074 635 2078
rect 727 2074 731 2078
rect 743 2074 747 2078
rect 831 2074 835 2078
rect 863 2074 867 2078
rect 935 2074 939 2078
rect 983 2074 987 2078
rect 1807 2130 1811 2134
rect 2135 2130 2139 2134
rect 2183 2130 2187 2134
rect 2255 2130 2259 2134
rect 2279 2130 2283 2134
rect 2383 2130 2387 2134
rect 2495 2130 2499 2134
rect 2519 2130 2523 2134
rect 2607 2130 2611 2134
rect 2655 2130 2659 2134
rect 1039 2074 1043 2078
rect 1143 2074 1147 2078
rect 1255 2074 1259 2078
rect 1767 2074 1771 2078
rect 1807 2058 1811 2062
rect 2135 2058 2139 2062
rect 111 2010 115 2014
rect 255 2010 259 2014
rect 359 2010 363 2014
rect 375 2010 379 2014
rect 487 2010 491 2014
rect 495 2010 499 2014
rect 615 2010 619 2014
rect 623 2010 627 2014
rect 727 2010 731 2014
rect 759 2010 763 2014
rect 111 1946 115 1950
rect 359 1946 363 1950
rect 447 1946 451 1950
rect 487 1946 491 1950
rect 575 1946 579 1950
rect 623 1946 627 1950
rect 2719 2130 2723 2134
rect 2783 2130 2787 2134
rect 2839 2130 2843 2134
rect 2911 2130 2915 2134
rect 2967 2130 2971 2134
rect 3031 2130 3035 2134
rect 3103 2130 3107 2134
rect 3151 2130 3155 2134
rect 3247 2130 3251 2134
rect 3271 2130 3275 2134
rect 3367 2202 3371 2206
rect 3463 2202 3467 2206
rect 3367 2130 3371 2134
rect 2247 2058 2251 2062
rect 2255 2058 2259 2062
rect 2383 2058 2387 2062
rect 2415 2058 2419 2062
rect 2519 2058 2523 2062
rect 2575 2058 2579 2062
rect 2655 2058 2659 2062
rect 2727 2058 2731 2062
rect 2783 2058 2787 2062
rect 2871 2058 2875 2062
rect 2911 2058 2915 2062
rect 3007 2058 3011 2062
rect 3031 2058 3035 2062
rect 3135 2058 3139 2062
rect 3151 2058 3155 2062
rect 3263 2058 3267 2062
rect 3271 2058 3275 2062
rect 831 2010 835 2014
rect 895 2010 899 2014
rect 935 2010 939 2014
rect 1023 2010 1027 2014
rect 1039 2010 1043 2014
rect 1143 2010 1147 2014
rect 1151 2010 1155 2014
rect 1255 2010 1259 2014
rect 1271 2010 1275 2014
rect 1399 2010 1403 2014
rect 1527 2010 1531 2014
rect 1767 2010 1771 2014
rect 711 1946 715 1950
rect 759 1946 763 1950
rect 847 1946 851 1950
rect 895 1946 899 1950
rect 111 1882 115 1886
rect 447 1882 451 1886
rect 559 1882 563 1886
rect 575 1882 579 1886
rect 695 1882 699 1886
rect 711 1882 715 1886
rect 831 1882 835 1886
rect 847 1882 851 1886
rect 983 1946 987 1950
rect 1023 1946 1027 1950
rect 1119 1946 1123 1950
rect 1151 1946 1155 1950
rect 1255 1946 1259 1950
rect 1271 1946 1275 1950
rect 1383 1946 1387 1950
rect 1399 1946 1403 1950
rect 1519 1946 1523 1950
rect 1527 1946 1531 1950
rect 1807 1978 1811 1982
rect 1831 1978 1835 1982
rect 1919 1978 1923 1982
rect 2047 1978 2051 1982
rect 2183 1978 2187 1982
rect 2247 1978 2251 1982
rect 2327 1978 2331 1982
rect 2415 1978 2419 1982
rect 2471 1978 2475 1982
rect 1655 1946 1659 1950
rect 1767 1946 1771 1950
rect 959 1882 963 1886
rect 983 1882 987 1886
rect 1079 1882 1083 1886
rect 1119 1882 1123 1886
rect 1199 1882 1203 1886
rect 1255 1882 1259 1886
rect 1327 1882 1331 1886
rect 1383 1882 1387 1886
rect 111 1810 115 1814
rect 135 1810 139 1814
rect 223 1810 227 1814
rect 311 1810 315 1814
rect 407 1810 411 1814
rect 527 1810 531 1814
rect 559 1810 563 1814
rect 655 1810 659 1814
rect 695 1810 699 1814
rect 799 1810 803 1814
rect 831 1810 835 1814
rect 943 1810 947 1814
rect 959 1810 963 1814
rect 1079 1810 1083 1814
rect 1087 1810 1091 1814
rect 1807 1910 1811 1914
rect 1831 1910 1835 1914
rect 1919 1910 1923 1914
rect 2039 1910 2043 1914
rect 2047 1910 2051 1914
rect 2167 1910 2171 1914
rect 2183 1910 2187 1914
rect 2303 1910 2307 1914
rect 2327 1910 2331 1914
rect 1455 1882 1459 1886
rect 1519 1882 1523 1886
rect 1655 1882 1659 1886
rect 1767 1882 1771 1886
rect 1807 1842 1811 1846
rect 1831 1842 1835 1846
rect 1199 1810 1203 1814
rect 1239 1810 1243 1814
rect 1327 1810 1331 1814
rect 1391 1810 1395 1814
rect 1455 1810 1459 1814
rect 1543 1810 1547 1814
rect 1671 1810 1675 1814
rect 1767 1810 1771 1814
rect 111 1734 115 1738
rect 135 1734 139 1738
rect 223 1734 227 1738
rect 247 1734 251 1738
rect 311 1734 315 1738
rect 399 1734 403 1738
rect 407 1734 411 1738
rect 527 1734 531 1738
rect 567 1734 571 1738
rect 655 1734 659 1738
rect 751 1734 755 1738
rect 799 1734 803 1738
rect 935 1734 939 1738
rect 943 1734 947 1738
rect 111 1666 115 1670
rect 135 1666 139 1670
rect 191 1666 195 1670
rect 247 1666 251 1670
rect 295 1666 299 1670
rect 399 1666 403 1670
rect 407 1666 411 1670
rect 1087 1734 1091 1738
rect 1119 1734 1123 1738
rect 1239 1734 1243 1738
rect 1311 1734 1315 1738
rect 535 1666 539 1670
rect 567 1666 571 1670
rect 687 1666 691 1670
rect 111 1598 115 1602
rect 191 1598 195 1602
rect 295 1598 299 1602
rect 327 1598 331 1602
rect 407 1598 411 1602
rect 431 1598 435 1602
rect 535 1598 539 1602
rect 543 1598 547 1602
rect 111 1530 115 1534
rect 223 1530 227 1534
rect 327 1530 331 1534
rect 343 1530 347 1534
rect 431 1530 435 1534
rect 751 1666 755 1670
rect 855 1666 859 1670
rect 935 1666 939 1670
rect 1039 1666 1043 1670
rect 1119 1666 1123 1670
rect 1919 1842 1923 1846
rect 1959 1842 1963 1846
rect 2039 1842 2043 1846
rect 2575 1978 2579 1982
rect 2615 1978 2619 1982
rect 2727 1978 2731 1982
rect 2751 1978 2755 1982
rect 2871 1978 2875 1982
rect 2887 1978 2891 1982
rect 3007 1978 3011 1982
rect 3031 1978 3035 1982
rect 3135 1978 3139 1982
rect 3175 1978 3179 1982
rect 3263 1978 3267 1982
rect 3319 1978 3323 1982
rect 2455 1910 2459 1914
rect 2471 1910 2475 1914
rect 3367 2058 3371 2062
rect 3367 1978 3371 1982
rect 2615 1910 2619 1914
rect 2751 1910 2755 1914
rect 2791 1910 2795 1914
rect 2887 1910 2891 1914
rect 2983 1910 2987 1914
rect 3031 1910 3035 1914
rect 3175 1910 3179 1914
rect 2111 1842 2115 1846
rect 2167 1842 2171 1846
rect 2255 1842 2259 1846
rect 2303 1842 2307 1846
rect 2407 1842 2411 1846
rect 1807 1766 1811 1770
rect 1831 1766 1835 1770
rect 1879 1766 1883 1770
rect 1959 1766 1963 1770
rect 2015 1766 2019 1770
rect 2111 1766 2115 1770
rect 2151 1766 2155 1770
rect 2255 1766 2259 1770
rect 2303 1766 2307 1770
rect 1391 1734 1395 1738
rect 1503 1734 1507 1738
rect 1543 1734 1547 1738
rect 1671 1734 1675 1738
rect 1767 1734 1771 1738
rect 1231 1666 1235 1670
rect 1311 1666 1315 1670
rect 1431 1666 1435 1670
rect 1503 1666 1507 1670
rect 1639 1666 1643 1670
rect 1671 1666 1675 1670
rect 671 1598 675 1602
rect 687 1598 691 1602
rect 815 1598 819 1602
rect 855 1598 859 1602
rect 967 1598 971 1602
rect 1039 1598 1043 1602
rect 1119 1598 1123 1602
rect 1231 1598 1235 1602
rect 1279 1598 1283 1602
rect 1431 1598 1435 1602
rect 1439 1598 1443 1602
rect 471 1530 475 1534
rect 543 1530 547 1534
rect 607 1530 611 1534
rect 671 1530 675 1534
rect 751 1530 755 1534
rect 111 1458 115 1462
rect 135 1458 139 1462
rect 223 1458 227 1462
rect 303 1458 307 1462
rect 343 1458 347 1462
rect 471 1458 475 1462
rect 111 1390 115 1394
rect 135 1390 139 1394
rect 279 1390 283 1394
rect 303 1390 307 1394
rect 815 1530 819 1534
rect 895 1530 899 1534
rect 967 1530 971 1534
rect 1047 1530 1051 1534
rect 1119 1530 1123 1534
rect 1807 1694 1811 1698
rect 1831 1694 1835 1698
rect 1879 1694 1883 1698
rect 1935 1694 1939 1698
rect 2015 1694 2019 1698
rect 2063 1694 2067 1698
rect 2151 1694 2155 1698
rect 2183 1694 2187 1698
rect 1767 1666 1771 1670
rect 2455 1842 2459 1846
rect 2567 1842 2571 1846
rect 2615 1842 2619 1846
rect 2743 1842 2747 1846
rect 2791 1842 2795 1846
rect 2935 1842 2939 1846
rect 2983 1842 2987 1846
rect 3183 1910 3187 1914
rect 3319 1910 3323 1914
rect 3367 1910 3371 1914
rect 3135 1842 3139 1846
rect 3183 1842 3187 1846
rect 3343 1842 3347 1846
rect 3367 1842 3371 1846
rect 2407 1766 2411 1770
rect 2479 1766 2483 1770
rect 2567 1766 2571 1770
rect 2687 1766 2691 1770
rect 2743 1766 2747 1770
rect 2911 1766 2915 1770
rect 2303 1694 2307 1698
rect 2311 1694 2315 1698
rect 1807 1622 1811 1626
rect 1831 1622 1835 1626
rect 1607 1598 1611 1602
rect 1639 1598 1643 1602
rect 1767 1598 1771 1602
rect 2439 1694 2443 1698
rect 2479 1694 2483 1698
rect 2575 1694 2579 1698
rect 2687 1694 2691 1698
rect 2727 1694 2731 1698
rect 2935 1766 2939 1770
rect 3135 1766 3139 1770
rect 3151 1766 3155 1770
rect 2887 1694 2891 1698
rect 2911 1694 2915 1698
rect 3047 1694 3051 1698
rect 3151 1694 3155 1698
rect 3215 1694 3219 1698
rect 1935 1622 1939 1626
rect 1943 1622 1947 1626
rect 2063 1622 2067 1626
rect 2087 1622 2091 1626
rect 2183 1622 2187 1626
rect 2231 1622 2235 1626
rect 2311 1622 2315 1626
rect 2367 1622 2371 1626
rect 1199 1530 1203 1534
rect 1279 1530 1283 1534
rect 1351 1530 1355 1534
rect 1807 1550 1811 1554
rect 1831 1550 1835 1554
rect 1839 1550 1843 1554
rect 1943 1550 1947 1554
rect 1991 1550 1995 1554
rect 2087 1550 2091 1554
rect 2151 1550 2155 1554
rect 2231 1550 2235 1554
rect 1439 1530 1443 1534
rect 1503 1530 1507 1534
rect 1607 1530 1611 1534
rect 1767 1530 1771 1534
rect 2439 1622 2443 1626
rect 2503 1622 2507 1626
rect 2575 1622 2579 1626
rect 2639 1622 2643 1626
rect 2727 1622 2731 1626
rect 2767 1622 2771 1626
rect 2887 1622 2891 1626
rect 2895 1622 2899 1626
rect 3015 1622 3019 1626
rect 3047 1622 3051 1626
rect 2303 1550 2307 1554
rect 2367 1550 2371 1554
rect 607 1458 611 1462
rect 631 1458 635 1462
rect 751 1458 755 1462
rect 783 1458 787 1462
rect 895 1458 899 1462
rect 927 1458 931 1462
rect 447 1390 451 1394
rect 471 1390 475 1394
rect 607 1390 611 1394
rect 631 1390 635 1394
rect 759 1390 763 1394
rect 783 1390 787 1394
rect 111 1322 115 1326
rect 135 1322 139 1326
rect 903 1390 907 1394
rect 927 1390 931 1394
rect 1047 1458 1051 1462
rect 1063 1458 1067 1462
rect 1199 1458 1203 1462
rect 1335 1458 1339 1462
rect 1351 1458 1355 1462
rect 1471 1458 1475 1462
rect 1503 1458 1507 1462
rect 1807 1478 1811 1482
rect 1839 1478 1843 1482
rect 1767 1458 1771 1462
rect 2455 1550 2459 1554
rect 2503 1550 2507 1554
rect 3135 1622 3139 1626
rect 3463 2130 3467 2134
rect 3463 2058 3467 2062
rect 3463 1978 3467 1982
rect 3463 1910 3467 1914
rect 3343 1766 3347 1770
rect 3367 1766 3371 1770
rect 3367 1694 3371 1698
rect 3463 1842 3467 1846
rect 3463 1766 3467 1770
rect 3463 1694 3467 1698
rect 3215 1622 3219 1626
rect 3263 1622 3267 1626
rect 3367 1622 3371 1626
rect 3463 1622 3467 1626
rect 2599 1550 2603 1554
rect 2639 1550 2643 1554
rect 2735 1550 2739 1554
rect 2767 1550 2771 1554
rect 2871 1550 2875 1554
rect 2895 1550 2899 1554
rect 3007 1550 3011 1554
rect 3015 1550 3019 1554
rect 3135 1550 3139 1554
rect 3143 1550 3147 1554
rect 3263 1550 3267 1554
rect 3367 1550 3371 1554
rect 3463 1550 3467 1554
rect 1943 1478 1947 1482
rect 1991 1478 1995 1482
rect 2055 1478 2059 1482
rect 2151 1478 2155 1482
rect 2191 1478 2195 1482
rect 2303 1478 2307 1482
rect 2335 1478 2339 1482
rect 2455 1478 2459 1482
rect 2479 1478 2483 1482
rect 1031 1390 1035 1394
rect 1063 1390 1067 1394
rect 1159 1390 1163 1394
rect 1199 1390 1203 1394
rect 1807 1406 1811 1410
rect 1943 1406 1947 1410
rect 2055 1406 2059 1410
rect 2095 1406 2099 1410
rect 2191 1406 2195 1410
rect 2199 1406 2203 1410
rect 2319 1406 2323 1410
rect 2335 1406 2339 1410
rect 1287 1390 1291 1394
rect 1335 1390 1339 1394
rect 1415 1390 1419 1394
rect 1471 1390 1475 1394
rect 1767 1390 1771 1394
rect 2599 1478 2603 1482
rect 2631 1478 2635 1482
rect 2735 1478 2739 1482
rect 2783 1478 2787 1482
rect 2871 1478 2875 1482
rect 2935 1478 2939 1482
rect 3007 1478 3011 1482
rect 3087 1478 3091 1482
rect 3143 1478 3147 1482
rect 2455 1406 2459 1410
rect 2479 1406 2483 1410
rect 2599 1406 2603 1410
rect 2631 1406 2635 1410
rect 279 1322 283 1326
rect 439 1322 443 1326
rect 447 1322 451 1326
rect 583 1322 587 1326
rect 607 1322 611 1326
rect 719 1322 723 1326
rect 759 1322 763 1326
rect 847 1322 851 1326
rect 903 1322 907 1326
rect 967 1322 971 1326
rect 1031 1322 1035 1326
rect 1079 1322 1083 1326
rect 1159 1322 1163 1326
rect 1191 1322 1195 1326
rect 111 1254 115 1258
rect 135 1254 139 1258
rect 239 1254 243 1258
rect 279 1254 283 1258
rect 367 1254 371 1258
rect 439 1254 443 1258
rect 495 1254 499 1258
rect 583 1254 587 1258
rect 615 1254 619 1258
rect 1287 1322 1291 1326
rect 1311 1322 1315 1326
rect 2743 1406 2747 1410
rect 2783 1406 2787 1410
rect 3239 1478 3243 1482
rect 3463 1478 3467 1482
rect 2887 1406 2891 1410
rect 2935 1406 2939 1410
rect 3031 1406 3035 1410
rect 3087 1406 3091 1410
rect 3175 1406 3179 1410
rect 3239 1406 3243 1410
rect 3327 1406 3331 1410
rect 3463 1406 3467 1410
rect 1807 1338 1811 1342
rect 2095 1338 2099 1342
rect 2103 1338 2107 1342
rect 2199 1338 2203 1342
rect 2239 1338 2243 1342
rect 2319 1338 2323 1342
rect 2383 1338 2387 1342
rect 2455 1338 2459 1342
rect 2535 1338 2539 1342
rect 2599 1338 2603 1342
rect 1415 1322 1419 1326
rect 1767 1322 1771 1326
rect 719 1254 723 1258
rect 735 1254 739 1258
rect 847 1254 851 1258
rect 959 1254 963 1258
rect 967 1254 971 1258
rect 111 1186 115 1190
rect 135 1186 139 1190
rect 239 1186 243 1190
rect 367 1186 371 1190
rect 375 1186 379 1190
rect 495 1186 499 1190
rect 511 1186 515 1190
rect 615 1186 619 1190
rect 111 1118 115 1122
rect 135 1118 139 1122
rect 1807 1274 1811 1278
rect 1935 1274 1939 1278
rect 2063 1274 2067 1278
rect 2103 1274 2107 1278
rect 2199 1274 2203 1278
rect 2239 1274 2243 1278
rect 1071 1254 1075 1258
rect 1079 1254 1083 1258
rect 1191 1254 1195 1258
rect 1311 1254 1315 1258
rect 1767 1254 1771 1258
rect 2687 1338 2691 1342
rect 2743 1338 2747 1342
rect 2839 1338 2843 1342
rect 2887 1338 2891 1342
rect 2991 1338 2995 1342
rect 3031 1338 3035 1342
rect 3143 1338 3147 1342
rect 3175 1338 3179 1342
rect 3303 1338 3307 1342
rect 3327 1338 3331 1342
rect 2343 1274 2347 1278
rect 2383 1274 2387 1278
rect 2495 1274 2499 1278
rect 2535 1274 2539 1278
rect 2655 1274 2659 1278
rect 2687 1274 2691 1278
rect 1807 1210 1811 1214
rect 1831 1210 1835 1214
rect 1935 1210 1939 1214
rect 2063 1210 2067 1214
rect 2079 1210 2083 1214
rect 2199 1210 2203 1214
rect 2231 1210 2235 1214
rect 655 1186 659 1190
rect 735 1186 739 1190
rect 791 1186 795 1190
rect 847 1186 851 1190
rect 927 1186 931 1190
rect 959 1186 963 1190
rect 1063 1186 1067 1190
rect 1071 1186 1075 1190
rect 1191 1186 1195 1190
rect 1199 1186 1203 1190
rect 1335 1186 1339 1190
rect 1767 1186 1771 1190
rect 191 1118 195 1122
rect 239 1118 243 1122
rect 335 1118 339 1122
rect 375 1118 379 1122
rect 495 1118 499 1122
rect 511 1118 515 1122
rect 655 1118 659 1122
rect 791 1118 795 1122
rect 815 1118 819 1122
rect 927 1118 931 1122
rect 967 1118 971 1122
rect 1063 1118 1067 1122
rect 1119 1118 1123 1122
rect 1199 1118 1203 1122
rect 1263 1118 1267 1122
rect 111 1046 115 1050
rect 191 1046 195 1050
rect 327 1046 331 1050
rect 335 1046 339 1050
rect 463 1046 467 1050
rect 495 1046 499 1050
rect 607 1046 611 1050
rect 655 1046 659 1050
rect 1807 1134 1811 1138
rect 1831 1134 1835 1138
rect 1863 1134 1867 1138
rect 1335 1118 1339 1122
rect 1407 1118 1411 1122
rect 1559 1118 1563 1122
rect 1767 1118 1771 1122
rect 2343 1210 2347 1214
rect 2391 1210 2395 1214
rect 2495 1210 2499 1214
rect 2543 1210 2547 1214
rect 2815 1274 2819 1278
rect 2839 1274 2843 1278
rect 2975 1274 2979 1278
rect 2991 1274 2995 1278
rect 3463 1338 3467 1342
rect 3143 1274 3147 1278
rect 3303 1274 3307 1278
rect 3463 1274 3467 1278
rect 2655 1210 2659 1214
rect 2695 1210 2699 1214
rect 2815 1210 2819 1214
rect 2847 1210 2851 1214
rect 2975 1210 2979 1214
rect 2999 1210 3003 1214
rect 3143 1210 3147 1214
rect 3159 1210 3163 1214
rect 3463 1210 3467 1214
rect 1935 1134 1939 1138
rect 1983 1134 1987 1138
rect 2079 1134 2083 1138
rect 2111 1134 2115 1138
rect 2231 1134 2235 1138
rect 2247 1134 2251 1138
rect 2383 1134 2387 1138
rect 2391 1134 2395 1138
rect 2511 1134 2515 1138
rect 2543 1134 2547 1138
rect 1807 1062 1811 1066
rect 1863 1062 1867 1066
rect 1983 1062 1987 1066
rect 2103 1062 2107 1066
rect 2111 1062 2115 1066
rect 2191 1062 2195 1066
rect 767 1046 771 1050
rect 815 1046 819 1050
rect 927 1046 931 1050
rect 967 1046 971 1050
rect 1079 1046 1083 1050
rect 1119 1046 1123 1050
rect 1231 1046 1235 1050
rect 1263 1046 1267 1050
rect 1383 1046 1387 1050
rect 1407 1046 1411 1050
rect 1535 1046 1539 1050
rect 1559 1046 1563 1050
rect 1671 1046 1675 1050
rect 1767 1046 1771 1050
rect 111 978 115 982
rect 327 978 331 982
rect 463 978 467 982
rect 471 978 475 982
rect 567 978 571 982
rect 607 978 611 982
rect 671 978 675 982
rect 767 978 771 982
rect 783 978 787 982
rect 887 978 891 982
rect 927 978 931 982
rect 991 978 995 982
rect 111 910 115 914
rect 471 910 475 914
rect 1079 978 1083 982
rect 1095 978 1099 982
rect 1199 978 1203 982
rect 1231 978 1235 982
rect 1295 978 1299 982
rect 1383 978 1387 982
rect 1391 978 1395 982
rect 2247 1062 2251 1066
rect 2279 1062 2283 1066
rect 2367 1062 2371 1066
rect 2383 1062 2387 1066
rect 2455 1062 2459 1066
rect 2511 1062 2515 1066
rect 2543 1062 2547 1066
rect 1487 978 1491 982
rect 1535 978 1539 982
rect 1583 978 1587 982
rect 567 910 571 914
rect 607 910 611 914
rect 671 910 675 914
rect 695 910 699 914
rect 783 910 787 914
rect 791 910 795 914
rect 887 910 891 914
rect 895 910 899 914
rect 991 910 995 914
rect 999 910 1003 914
rect 1807 998 1811 1002
rect 2103 998 2107 1002
rect 2191 998 2195 1002
rect 2279 998 2283 1002
rect 2311 998 2315 1002
rect 2367 998 2371 1002
rect 2407 998 2411 1002
rect 2455 998 2459 1002
rect 1671 978 1675 982
rect 1767 978 1771 982
rect 2639 1134 2643 1138
rect 2695 1134 2699 1138
rect 2759 1134 2763 1138
rect 2847 1134 2851 1138
rect 2871 1134 2875 1138
rect 2975 1134 2979 1138
rect 2999 1134 3003 1138
rect 3079 1134 3083 1138
rect 3159 1134 3163 1138
rect 3183 1134 3187 1138
rect 3279 1134 3283 1138
rect 3367 1134 3371 1138
rect 3463 1134 3467 1138
rect 2631 1062 2635 1066
rect 2639 1062 2643 1066
rect 2719 1062 2723 1066
rect 2759 1062 2763 1066
rect 2807 1062 2811 1066
rect 2871 1062 2875 1066
rect 2975 1062 2979 1066
rect 3079 1062 3083 1066
rect 3183 1062 3187 1066
rect 3279 1062 3283 1066
rect 3367 1062 3371 1066
rect 2511 998 2515 1002
rect 2543 998 2547 1002
rect 2623 998 2627 1002
rect 2631 998 2635 1002
rect 2719 998 2723 1002
rect 2751 998 2755 1002
rect 2807 998 2811 1002
rect 1807 922 1811 926
rect 1831 922 1835 926
rect 1983 922 1987 926
rect 2151 922 2155 926
rect 1095 910 1099 914
rect 1111 910 1115 914
rect 1199 910 1203 914
rect 1223 910 1227 914
rect 1295 910 1299 914
rect 1343 910 1347 914
rect 111 842 115 846
rect 519 842 523 846
rect 607 842 611 846
rect 615 842 619 846
rect 695 842 699 846
rect 719 842 723 846
rect 791 842 795 846
rect 831 842 835 846
rect 895 842 899 846
rect 951 842 955 846
rect 999 842 1003 846
rect 1391 910 1395 914
rect 1463 910 1467 914
rect 1487 910 1491 914
rect 1583 910 1587 914
rect 1671 910 1675 914
rect 1767 910 1771 914
rect 1071 842 1075 846
rect 1111 842 1115 846
rect 1191 842 1195 846
rect 111 774 115 778
rect 383 774 387 778
rect 471 774 475 778
rect 519 774 523 778
rect 575 774 579 778
rect 615 774 619 778
rect 679 774 683 778
rect 719 774 723 778
rect 791 774 795 778
rect 111 702 115 706
rect 247 702 251 706
rect 343 702 347 706
rect 383 702 387 706
rect 455 702 459 706
rect 471 702 475 706
rect 567 702 571 706
rect 575 702 579 706
rect 831 774 835 778
rect 911 774 915 778
rect 951 774 955 778
rect 1031 774 1035 778
rect 1071 774 1075 778
rect 1223 842 1227 846
rect 1311 842 1315 846
rect 1343 842 1347 846
rect 1431 842 1435 846
rect 1463 842 1467 846
rect 1559 842 1563 846
rect 1583 842 1587 846
rect 1807 854 1811 858
rect 1831 854 1835 858
rect 1767 842 1771 846
rect 1159 774 1163 778
rect 1191 774 1195 778
rect 1959 854 1963 858
rect 1983 854 1987 858
rect 2895 998 2899 1002
rect 3055 998 3059 1002
rect 3223 998 3227 1002
rect 3367 998 3371 1002
rect 3463 1062 3467 1066
rect 3463 998 3467 1002
rect 2311 922 2315 926
rect 2327 922 2331 926
rect 2407 922 2411 926
rect 2511 922 2515 926
rect 2519 922 2523 926
rect 2623 922 2627 926
rect 2719 922 2723 926
rect 2751 922 2755 926
rect 2895 922 2899 926
rect 2935 922 2939 926
rect 3055 922 3059 926
rect 3159 922 3163 926
rect 3223 922 3227 926
rect 3367 922 3371 926
rect 3463 922 3467 926
rect 2087 854 2091 858
rect 2151 854 2155 858
rect 2207 854 2211 858
rect 2327 854 2331 858
rect 1807 786 1811 790
rect 1831 786 1835 790
rect 1879 786 1883 790
rect 1959 786 1963 790
rect 2015 786 2019 790
rect 1287 774 1291 778
rect 1311 774 1315 778
rect 1415 774 1419 778
rect 1431 774 1435 778
rect 1559 774 1563 778
rect 1767 774 1771 778
rect 2087 786 2091 790
rect 2151 786 2155 790
rect 2207 786 2211 790
rect 2463 854 2467 858
rect 2519 854 2523 858
rect 2615 854 2619 858
rect 2719 854 2723 858
rect 2791 854 2795 858
rect 2935 854 2939 858
rect 2983 854 2987 858
rect 3159 854 3163 858
rect 3183 854 3187 858
rect 3367 854 3371 858
rect 3463 854 3467 858
rect 2287 786 2291 790
rect 2327 786 2331 790
rect 2423 786 2427 790
rect 2463 786 2467 790
rect 2559 786 2563 790
rect 2615 786 2619 790
rect 2711 786 2715 790
rect 2791 786 2795 790
rect 2871 786 2875 790
rect 2983 786 2987 790
rect 3039 786 3043 790
rect 3183 786 3187 790
rect 3215 786 3219 790
rect 3367 786 3371 790
rect 679 702 683 706
rect 695 702 699 706
rect 791 702 795 706
rect 831 702 835 706
rect 911 702 915 706
rect 983 702 987 706
rect 111 634 115 638
rect 135 634 139 638
rect 231 634 235 638
rect 247 634 251 638
rect 343 634 347 638
rect 359 634 363 638
rect 455 634 459 638
rect 487 634 491 638
rect 567 634 571 638
rect 623 634 627 638
rect 695 634 699 638
rect 767 634 771 638
rect 111 566 115 570
rect 135 566 139 570
rect 1807 718 1811 722
rect 1831 718 1835 722
rect 1879 718 1883 722
rect 1951 718 1955 722
rect 1031 702 1035 706
rect 1151 702 1155 706
rect 1159 702 1163 706
rect 1287 702 1291 706
rect 1327 702 1331 706
rect 1415 702 1419 706
rect 1511 702 1515 706
rect 1671 702 1675 706
rect 1767 702 1771 706
rect 831 634 835 638
rect 911 634 915 638
rect 983 634 987 638
rect 1055 634 1059 638
rect 1151 634 1155 638
rect 1207 634 1211 638
rect 231 566 235 570
rect 247 566 251 570
rect 359 566 363 570
rect 407 566 411 570
rect 487 566 491 570
rect 583 566 587 570
rect 623 566 627 570
rect 767 566 771 570
rect 911 566 915 570
rect 951 566 955 570
rect 111 498 115 502
rect 135 498 139 502
rect 247 498 251 502
rect 399 498 403 502
rect 407 498 411 502
rect 567 498 571 502
rect 583 498 587 502
rect 1055 566 1059 570
rect 1327 634 1331 638
rect 1367 634 1371 638
rect 1511 634 1515 638
rect 1527 634 1531 638
rect 1671 634 1675 638
rect 2015 718 2019 722
rect 2103 718 2107 722
rect 2151 718 2155 722
rect 2263 718 2267 722
rect 2287 718 2291 722
rect 2415 718 2419 722
rect 2423 718 2427 722
rect 3463 786 3467 790
rect 2559 718 2563 722
rect 2567 718 2571 722
rect 2711 718 2715 722
rect 2719 718 2723 722
rect 2871 718 2875 722
rect 2879 718 2883 722
rect 3039 718 3043 722
rect 3199 718 3203 722
rect 3215 718 3219 722
rect 1807 654 1811 658
rect 1831 654 1835 658
rect 1951 654 1955 658
rect 1975 654 1979 658
rect 2103 654 2107 658
rect 1767 634 1771 638
rect 1135 566 1139 570
rect 1207 566 1211 570
rect 1319 566 1323 570
rect 1367 566 1371 570
rect 1807 582 1811 586
rect 1895 582 1899 586
rect 1503 566 1507 570
rect 1527 566 1531 570
rect 1671 566 1675 570
rect 1767 566 1771 570
rect 2239 654 2243 658
rect 2263 654 2267 658
rect 2415 654 2419 658
rect 2479 654 2483 658
rect 2567 654 2571 658
rect 1975 582 1979 586
rect 2015 582 2019 586
rect 2143 582 2147 586
rect 2239 582 2243 586
rect 2279 582 2283 586
rect 2423 582 2427 586
rect 2479 582 2483 586
rect 2567 582 2571 586
rect 735 498 739 502
rect 767 498 771 502
rect 903 498 907 502
rect 951 498 955 502
rect 1063 498 1067 502
rect 1135 498 1139 502
rect 1223 498 1227 502
rect 1319 498 1323 502
rect 1375 498 1379 502
rect 1503 498 1507 502
rect 1527 498 1531 502
rect 1671 498 1675 502
rect 111 430 115 434
rect 247 430 251 434
rect 399 430 403 434
rect 519 430 523 434
rect 567 430 571 434
rect 615 430 619 434
rect 719 430 723 434
rect 735 430 739 434
rect 823 430 827 434
rect 903 430 907 434
rect 927 430 931 434
rect 1807 514 1811 518
rect 1895 514 1899 518
rect 2015 514 2019 518
rect 2135 514 2139 518
rect 2143 514 2147 518
rect 2239 514 2243 518
rect 1767 498 1771 502
rect 2279 514 2283 518
rect 2359 514 2363 518
rect 2423 514 2427 518
rect 2687 654 2691 658
rect 2719 654 2723 658
rect 2879 654 2883 658
rect 2687 582 2691 586
rect 2719 582 2723 586
rect 3039 654 3043 658
rect 3055 654 3059 658
rect 3367 718 3371 722
rect 3199 654 3203 658
rect 3223 654 3227 658
rect 3367 654 3371 658
rect 2871 582 2875 586
rect 2879 582 2883 586
rect 3031 582 3035 586
rect 3055 582 3059 586
rect 2487 514 2491 518
rect 2567 514 2571 518
rect 2615 514 2619 518
rect 2719 514 2723 518
rect 2751 514 2755 518
rect 1023 430 1027 434
rect 1063 430 1067 434
rect 1127 430 1131 434
rect 1223 430 1227 434
rect 1231 430 1235 434
rect 111 362 115 366
rect 471 362 475 366
rect 519 362 523 366
rect 559 362 563 366
rect 615 362 619 366
rect 647 362 651 366
rect 719 362 723 366
rect 735 362 739 366
rect 823 362 827 366
rect 111 294 115 298
rect 279 294 283 298
rect 367 294 371 298
rect 463 294 467 298
rect 471 294 475 298
rect 559 294 563 298
rect 911 362 915 366
rect 927 362 931 366
rect 999 362 1003 366
rect 1023 362 1027 366
rect 1087 362 1091 366
rect 1127 362 1131 366
rect 1175 362 1179 366
rect 1807 442 1811 446
rect 2135 442 2139 446
rect 2239 442 2243 446
rect 2335 442 2339 446
rect 2359 442 2363 446
rect 2447 442 2451 446
rect 2487 442 2491 446
rect 2559 442 2563 446
rect 2615 442 2619 446
rect 1335 430 1339 434
rect 1375 430 1379 434
rect 1439 430 1443 434
rect 1527 430 1531 434
rect 1671 430 1675 434
rect 1767 430 1771 434
rect 2871 514 2875 518
rect 2879 514 2883 518
rect 3007 514 3011 518
rect 3031 514 3035 518
rect 3135 514 3139 518
rect 2679 442 2683 446
rect 2751 442 2755 446
rect 2799 442 2803 446
rect 2879 442 2883 446
rect 2911 442 2915 446
rect 3007 442 3011 446
rect 3023 442 3027 446
rect 3199 582 3203 586
rect 3223 582 3227 586
rect 3367 582 3371 586
rect 3463 718 3467 722
rect 3463 654 3467 658
rect 3463 582 3467 586
rect 3199 514 3203 518
rect 3263 514 3267 518
rect 3367 514 3371 518
rect 3463 514 3467 518
rect 3135 442 3139 446
rect 3143 442 3147 446
rect 3263 442 3267 446
rect 1807 374 1811 378
rect 2063 374 2067 378
rect 2151 374 2155 378
rect 2239 374 2243 378
rect 2247 374 2251 378
rect 2335 374 2339 378
rect 2359 374 2363 378
rect 2447 374 2451 378
rect 1231 362 1235 366
rect 1263 362 1267 366
rect 1335 362 1339 366
rect 1439 362 1443 366
rect 1767 362 1771 366
rect 647 294 651 298
rect 655 294 659 298
rect 735 294 739 298
rect 751 294 755 298
rect 823 294 827 298
rect 847 294 851 298
rect 1807 306 1811 310
rect 1927 306 1931 310
rect 2039 306 2043 310
rect 2063 306 2067 310
rect 2151 306 2155 310
rect 2167 306 2171 310
rect 2247 306 2251 310
rect 2303 306 2307 310
rect 2359 306 2363 310
rect 911 294 915 298
rect 943 294 947 298
rect 999 294 1003 298
rect 1047 294 1051 298
rect 1087 294 1091 298
rect 1151 294 1155 298
rect 1175 294 1179 298
rect 1263 294 1267 298
rect 1767 294 1771 298
rect 2479 374 2483 378
rect 2559 374 2563 378
rect 2615 374 2619 378
rect 2679 374 2683 378
rect 2759 374 2763 378
rect 2799 374 2803 378
rect 2911 374 2915 378
rect 3367 442 3371 446
rect 3463 442 3467 446
rect 3023 374 3027 378
rect 3063 374 3067 378
rect 3143 374 3147 378
rect 3223 374 3227 378
rect 3263 374 3267 378
rect 2447 306 2451 310
rect 2479 306 2483 310
rect 2599 306 2603 310
rect 2615 306 2619 310
rect 1807 238 1811 242
rect 1831 238 1835 242
rect 1927 238 1931 242
rect 2039 238 2043 242
rect 2055 238 2059 242
rect 2167 238 2171 242
rect 2199 238 2203 242
rect 2303 238 2307 242
rect 2351 238 2355 242
rect 111 226 115 230
rect 167 226 171 230
rect 279 226 283 230
rect 343 226 347 230
rect 367 226 371 230
rect 463 226 467 230
rect 511 226 515 230
rect 559 226 563 230
rect 655 226 659 230
rect 679 226 683 230
rect 751 226 755 230
rect 839 226 843 230
rect 847 226 851 230
rect 943 226 947 230
rect 991 226 995 230
rect 1047 226 1051 230
rect 1135 226 1139 230
rect 1151 226 1155 230
rect 1279 226 1283 230
rect 1431 226 1435 230
rect 1767 226 1771 230
rect 231 160 235 164
rect 743 160 747 164
rect 111 138 115 142
rect 135 138 139 142
rect 167 138 171 142
rect 223 138 227 142
rect 311 138 315 142
rect 343 138 347 142
rect 399 138 403 142
rect 487 138 491 142
rect 511 138 515 142
rect 575 138 579 142
rect 663 138 667 142
rect 679 138 683 142
rect 751 138 755 142
rect 839 138 843 142
rect 847 138 851 142
rect 943 138 947 142
rect 991 138 995 142
rect 1031 138 1035 142
rect 1119 138 1123 142
rect 1135 138 1139 142
rect 1215 138 1219 142
rect 1279 138 1283 142
rect 1311 138 1315 142
rect 903 88 907 92
rect 111 74 115 78
rect 135 74 139 78
rect 223 74 227 78
rect 311 74 315 78
rect 399 74 403 78
rect 487 74 491 78
rect 575 74 579 78
rect 663 74 667 78
rect 751 74 755 78
rect 1807 154 1811 158
rect 1831 154 1835 158
rect 1919 154 1923 158
rect 1927 154 1931 158
rect 2039 154 2043 158
rect 2055 154 2059 158
rect 2159 154 2163 158
rect 2199 154 2203 158
rect 1407 138 1411 142
rect 1431 138 1435 142
rect 1495 138 1499 142
rect 1583 138 1587 142
rect 1671 138 1675 142
rect 1767 138 1771 142
rect 2447 238 2451 242
rect 2511 238 2515 242
rect 2599 238 2603 242
rect 2759 306 2763 310
rect 2911 306 2915 310
rect 2919 306 2923 310
rect 3063 306 3067 310
rect 3087 306 3091 310
rect 3223 306 3227 310
rect 3255 306 3259 310
rect 2679 238 2683 242
rect 2759 238 2763 242
rect 3367 374 3371 378
rect 3463 374 3467 378
rect 3367 306 3371 310
rect 2847 238 2851 242
rect 2919 238 2923 242
rect 3023 238 3027 242
rect 3087 238 3091 242
rect 3207 238 3211 242
rect 3255 238 3259 242
rect 3367 238 3371 242
rect 2279 154 2283 158
rect 2351 154 2355 158
rect 2399 154 2403 158
rect 1399 88 1403 92
rect 2511 154 2515 158
rect 2623 154 2627 158
rect 2679 154 2683 158
rect 2735 154 2739 158
rect 2839 154 2843 158
rect 2847 154 2851 158
rect 2943 154 2947 158
rect 3023 154 3027 158
rect 3055 154 3059 158
rect 3167 154 3171 158
rect 3207 154 3211 158
rect 1807 90 1811 94
rect 1831 90 1835 94
rect 1919 90 1923 94
rect 2039 90 2043 94
rect 2159 90 2163 94
rect 2279 90 2283 94
rect 3279 154 3283 158
rect 3367 154 3371 158
rect 3463 306 3467 310
rect 3463 238 3467 242
rect 3463 154 3467 158
rect 2399 90 2403 94
rect 2511 90 2515 94
rect 2623 90 2627 94
rect 2735 90 2739 94
rect 2839 90 2843 94
rect 2943 90 2947 94
rect 3055 90 3059 94
rect 3167 90 3171 94
rect 3279 90 3283 94
rect 3367 90 3371 94
rect 3463 90 3467 94
rect 847 74 851 78
rect 943 74 947 78
rect 1031 74 1035 78
rect 1119 74 1123 78
rect 1215 74 1219 78
rect 1311 74 1315 78
rect 1407 74 1411 78
rect 1495 74 1499 78
rect 1583 74 1587 78
rect 1671 74 1675 78
rect 1767 74 1771 78
<< m4 >>
rect 1790 3517 1791 3523
rect 1797 3522 3499 3523
rect 1797 3518 1807 3522
rect 1811 3518 2007 3522
rect 2011 3518 2239 3522
rect 2243 3518 2455 3522
rect 2459 3518 2655 3522
rect 2659 3518 2855 3522
rect 2859 3518 3047 3522
rect 3051 3518 3247 3522
rect 3251 3518 3463 3522
rect 3467 3518 3499 3522
rect 1797 3517 3499 3518
rect 3505 3517 3506 3523
rect 96 3481 97 3487
rect 103 3486 1791 3487
rect 103 3482 111 3486
rect 115 3482 455 3486
rect 459 3482 543 3486
rect 547 3482 631 3486
rect 635 3482 719 3486
rect 723 3482 807 3486
rect 811 3482 895 3486
rect 899 3482 983 3486
rect 987 3482 1071 3486
rect 1075 3482 1159 3486
rect 1163 3482 1767 3486
rect 1771 3482 1791 3486
rect 103 3481 1791 3482
rect 1797 3481 1798 3487
rect 1778 3453 1779 3459
rect 1785 3458 3487 3459
rect 1785 3454 1807 3458
rect 1811 3454 1831 3458
rect 1835 3454 1943 3458
rect 1947 3454 2007 3458
rect 2011 3454 2079 3458
rect 2083 3454 2215 3458
rect 2219 3454 2239 3458
rect 2243 3454 2351 3458
rect 2355 3454 2455 3458
rect 2459 3454 2479 3458
rect 2483 3454 2599 3458
rect 2603 3454 2655 3458
rect 2659 3454 2719 3458
rect 2723 3454 2847 3458
rect 2851 3454 2855 3458
rect 2859 3454 2975 3458
rect 2979 3454 3047 3458
rect 3051 3454 3247 3458
rect 3251 3454 3463 3458
rect 3467 3454 3487 3458
rect 1785 3453 3487 3454
rect 3493 3453 3494 3459
rect 84 3417 85 3423
rect 91 3422 1779 3423
rect 91 3418 111 3422
rect 115 3418 415 3422
rect 419 3418 455 3422
rect 459 3418 503 3422
rect 507 3418 543 3422
rect 547 3418 591 3422
rect 595 3418 631 3422
rect 635 3418 679 3422
rect 683 3418 719 3422
rect 723 3418 767 3422
rect 771 3418 807 3422
rect 811 3418 855 3422
rect 859 3418 895 3422
rect 899 3418 943 3422
rect 947 3418 983 3422
rect 987 3418 1031 3422
rect 1035 3418 1071 3422
rect 1075 3418 1119 3422
rect 1123 3418 1159 3422
rect 1163 3418 1207 3422
rect 1211 3418 1303 3422
rect 1307 3418 1767 3422
rect 1771 3418 1779 3422
rect 91 3417 1779 3418
rect 1785 3417 1786 3423
rect 1790 3381 1791 3387
rect 1797 3386 3499 3387
rect 1797 3382 1807 3386
rect 1811 3382 1831 3386
rect 1835 3382 1943 3386
rect 1947 3382 1951 3386
rect 1955 3382 2079 3386
rect 2083 3382 2095 3386
rect 2099 3382 2215 3386
rect 2219 3382 2239 3386
rect 2243 3382 2351 3386
rect 2355 3382 2383 3386
rect 2387 3382 2479 3386
rect 2483 3382 2519 3386
rect 2523 3382 2599 3386
rect 2603 3382 2647 3386
rect 2651 3382 2719 3386
rect 2723 3382 2775 3386
rect 2779 3382 2847 3386
rect 2851 3382 2903 3386
rect 2907 3382 2975 3386
rect 2979 3382 3039 3386
rect 3043 3382 3463 3386
rect 3467 3382 3499 3386
rect 1797 3381 3499 3382
rect 3505 3381 3506 3387
rect 96 3349 97 3355
rect 103 3354 1791 3355
rect 103 3350 111 3354
rect 115 3350 399 3354
rect 403 3350 415 3354
rect 419 3350 495 3354
rect 499 3350 503 3354
rect 507 3350 591 3354
rect 595 3350 599 3354
rect 603 3350 679 3354
rect 683 3350 703 3354
rect 707 3350 767 3354
rect 771 3350 807 3354
rect 811 3350 855 3354
rect 859 3350 911 3354
rect 915 3350 943 3354
rect 947 3350 1015 3354
rect 1019 3350 1031 3354
rect 1035 3350 1119 3354
rect 1123 3350 1207 3354
rect 1211 3350 1223 3354
rect 1227 3350 1303 3354
rect 1307 3350 1327 3354
rect 1331 3350 1767 3354
rect 1771 3350 1791 3354
rect 103 3349 1791 3350
rect 1797 3349 1798 3355
rect 1778 3309 1779 3315
rect 1785 3314 3487 3315
rect 1785 3310 1807 3314
rect 1811 3310 1831 3314
rect 1835 3310 1951 3314
rect 1955 3310 1975 3314
rect 1979 3310 2095 3314
rect 2099 3310 2151 3314
rect 2155 3310 2239 3314
rect 2243 3310 2335 3314
rect 2339 3310 2383 3314
rect 2387 3310 2511 3314
rect 2515 3310 2519 3314
rect 2523 3310 2647 3314
rect 2651 3310 2679 3314
rect 2683 3310 2775 3314
rect 2779 3310 2831 3314
rect 2835 3310 2903 3314
rect 2907 3310 2975 3314
rect 2979 3310 3039 3314
rect 3043 3310 3111 3314
rect 3115 3310 3247 3314
rect 3251 3310 3367 3314
rect 3371 3310 3463 3314
rect 3467 3310 3487 3314
rect 1785 3309 3487 3310
rect 3493 3309 3494 3315
rect 84 3281 85 3287
rect 91 3286 1779 3287
rect 91 3282 111 3286
rect 115 3282 383 3286
rect 387 3282 399 3286
rect 403 3282 495 3286
rect 499 3282 599 3286
rect 603 3282 607 3286
rect 611 3282 703 3286
rect 707 3282 727 3286
rect 731 3282 807 3286
rect 811 3282 847 3286
rect 851 3282 911 3286
rect 915 3282 967 3286
rect 971 3282 1015 3286
rect 1019 3282 1087 3286
rect 1091 3282 1119 3286
rect 1123 3282 1207 3286
rect 1211 3282 1223 3286
rect 1227 3282 1327 3286
rect 1331 3282 1335 3286
rect 1339 3282 1767 3286
rect 1771 3282 1779 3286
rect 91 3281 1779 3282
rect 1785 3281 1786 3287
rect 1790 3237 1791 3243
rect 1797 3242 3499 3243
rect 1797 3238 1807 3242
rect 1811 3238 1831 3242
rect 1835 3238 1975 3242
rect 1979 3238 2031 3242
rect 2035 3238 2151 3242
rect 2155 3238 2247 3242
rect 2251 3238 2335 3242
rect 2339 3238 2455 3242
rect 2459 3238 2511 3242
rect 2515 3238 2655 3242
rect 2659 3238 2679 3242
rect 2683 3238 2831 3242
rect 2835 3238 2839 3242
rect 2843 3238 2975 3242
rect 2979 3238 3023 3242
rect 3027 3238 3111 3242
rect 3115 3238 3207 3242
rect 3211 3238 3247 3242
rect 3251 3238 3367 3242
rect 3371 3238 3463 3242
rect 3467 3238 3499 3242
rect 1797 3237 3499 3238
rect 3505 3237 3506 3243
rect 96 3213 97 3219
rect 103 3218 1791 3219
rect 103 3214 111 3218
rect 115 3214 303 3218
rect 307 3214 383 3218
rect 387 3214 423 3218
rect 427 3214 495 3218
rect 499 3214 543 3218
rect 547 3214 607 3218
rect 611 3214 671 3218
rect 675 3214 727 3218
rect 731 3214 799 3218
rect 803 3214 847 3218
rect 851 3214 927 3218
rect 931 3214 967 3218
rect 971 3214 1055 3218
rect 1059 3214 1087 3218
rect 1091 3214 1175 3218
rect 1179 3214 1207 3218
rect 1211 3214 1303 3218
rect 1307 3214 1335 3218
rect 1339 3214 1431 3218
rect 1435 3214 1767 3218
rect 1771 3214 1791 3218
rect 103 3213 1791 3214
rect 1797 3213 1798 3219
rect 1778 3173 1779 3179
rect 1785 3178 3487 3179
rect 1785 3174 1807 3178
rect 1811 3174 1831 3178
rect 1835 3174 1839 3178
rect 1843 3174 2031 3178
rect 2035 3174 2223 3178
rect 2227 3174 2247 3178
rect 2251 3174 2407 3178
rect 2411 3174 2455 3178
rect 2459 3174 2575 3178
rect 2579 3174 2655 3178
rect 2659 3174 2735 3178
rect 2739 3174 2839 3178
rect 2843 3174 2879 3178
rect 2883 3174 3007 3178
rect 3011 3174 3023 3178
rect 3027 3174 3135 3178
rect 3139 3174 3207 3178
rect 3211 3174 3263 3178
rect 3267 3174 3367 3178
rect 3371 3174 3463 3178
rect 3467 3174 3487 3178
rect 1785 3173 3487 3174
rect 3493 3173 3494 3179
rect 84 3137 85 3143
rect 91 3142 1779 3143
rect 91 3138 111 3142
rect 115 3138 175 3142
rect 179 3138 303 3142
rect 307 3138 319 3142
rect 323 3138 423 3142
rect 427 3138 471 3142
rect 475 3138 543 3142
rect 547 3138 623 3142
rect 627 3138 671 3142
rect 675 3138 775 3142
rect 779 3138 799 3142
rect 803 3138 919 3142
rect 923 3138 927 3142
rect 931 3138 1055 3142
rect 1059 3138 1063 3142
rect 1067 3138 1175 3142
rect 1179 3138 1199 3142
rect 1203 3138 1303 3142
rect 1307 3138 1343 3142
rect 1347 3138 1431 3142
rect 1435 3138 1487 3142
rect 1491 3138 1767 3142
rect 1771 3138 1779 3142
rect 91 3137 1779 3138
rect 1785 3137 1786 3143
rect 1790 3105 1791 3111
rect 1797 3110 3499 3111
rect 1797 3106 1807 3110
rect 1811 3106 1839 3110
rect 1843 3106 1935 3110
rect 1939 3106 2031 3110
rect 2035 3106 2055 3110
rect 2059 3106 2175 3110
rect 2179 3106 2223 3110
rect 2227 3106 2303 3110
rect 2307 3106 2407 3110
rect 2411 3106 2431 3110
rect 2435 3106 2567 3110
rect 2571 3106 2575 3110
rect 2579 3106 2719 3110
rect 2723 3106 2735 3110
rect 2739 3106 2871 3110
rect 2875 3106 2879 3110
rect 2883 3106 3007 3110
rect 3011 3106 3031 3110
rect 3035 3106 3135 3110
rect 3139 3106 3199 3110
rect 3203 3106 3263 3110
rect 3267 3106 3367 3110
rect 3371 3106 3463 3110
rect 3467 3106 3499 3110
rect 1797 3105 3499 3106
rect 3505 3105 3506 3111
rect 96 3065 97 3071
rect 103 3070 1791 3071
rect 103 3066 111 3070
rect 115 3066 135 3070
rect 139 3066 175 3070
rect 179 3066 263 3070
rect 267 3066 319 3070
rect 323 3066 431 3070
rect 435 3066 471 3070
rect 475 3066 607 3070
rect 611 3066 623 3070
rect 627 3066 775 3070
rect 779 3066 791 3070
rect 795 3066 919 3070
rect 923 3066 967 3070
rect 971 3066 1063 3070
rect 1067 3066 1143 3070
rect 1147 3066 1199 3070
rect 1203 3066 1327 3070
rect 1331 3066 1343 3070
rect 1347 3066 1487 3070
rect 1491 3066 1511 3070
rect 1515 3066 1767 3070
rect 1771 3066 1791 3070
rect 103 3065 1791 3066
rect 1797 3065 1798 3071
rect 1778 3033 1779 3039
rect 1785 3038 3487 3039
rect 1785 3034 1807 3038
rect 1811 3034 1935 3038
rect 1939 3034 2023 3038
rect 2027 3034 2055 3038
rect 2059 3034 2127 3038
rect 2131 3034 2175 3038
rect 2179 3034 2231 3038
rect 2235 3034 2303 3038
rect 2307 3034 2335 3038
rect 2339 3034 2431 3038
rect 2435 3034 2439 3038
rect 2443 3034 2543 3038
rect 2547 3034 2567 3038
rect 2571 3034 2647 3038
rect 2651 3034 2719 3038
rect 2723 3034 2759 3038
rect 2763 3034 2871 3038
rect 2875 3034 3031 3038
rect 3035 3034 3199 3038
rect 3203 3034 3367 3038
rect 3371 3034 3463 3038
rect 3467 3034 3487 3038
rect 1785 3033 3487 3034
rect 3493 3033 3494 3039
rect 84 2997 85 3003
rect 91 3002 1779 3003
rect 91 2998 111 3002
rect 115 2998 135 3002
rect 139 2998 263 3002
rect 267 2998 327 3002
rect 331 2998 431 3002
rect 435 2998 535 3002
rect 539 2998 607 3002
rect 611 2998 735 3002
rect 739 2998 791 3002
rect 795 2998 927 3002
rect 931 2998 967 3002
rect 971 2998 1103 3002
rect 1107 2998 1143 3002
rect 1147 2998 1279 3002
rect 1283 2998 1327 3002
rect 1331 2998 1447 3002
rect 1451 2998 1511 3002
rect 1515 2998 1623 3002
rect 1627 2998 1767 3002
rect 1771 2998 1779 3002
rect 91 2997 1779 2998
rect 1785 2997 1786 3003
rect 1790 2969 1791 2975
rect 1797 2974 3499 2975
rect 1797 2970 1807 2974
rect 1811 2970 2023 2974
rect 2027 2970 2055 2974
rect 2059 2970 2127 2974
rect 2131 2970 2143 2974
rect 2147 2970 2231 2974
rect 2235 2970 2319 2974
rect 2323 2970 2335 2974
rect 2339 2970 2407 2974
rect 2411 2970 2439 2974
rect 2443 2970 2495 2974
rect 2499 2970 2543 2974
rect 2547 2970 2583 2974
rect 2587 2970 2647 2974
rect 2651 2970 2671 2974
rect 2675 2970 2759 2974
rect 2763 2970 2847 2974
rect 2851 2970 3463 2974
rect 3467 2970 3499 2974
rect 1797 2969 3499 2970
rect 3505 2969 3506 2975
rect 96 2925 97 2931
rect 103 2930 1791 2931
rect 103 2926 111 2930
rect 115 2926 135 2930
rect 139 2926 263 2930
rect 267 2926 327 2930
rect 331 2926 431 2930
rect 435 2926 535 2930
rect 539 2926 607 2930
rect 611 2926 735 2930
rect 739 2926 783 2930
rect 787 2926 927 2930
rect 931 2926 951 2930
rect 955 2926 1103 2930
rect 1107 2926 1111 2930
rect 1115 2926 1271 2930
rect 1275 2926 1279 2930
rect 1283 2926 1431 2930
rect 1435 2926 1447 2930
rect 1451 2926 1591 2930
rect 1595 2926 1623 2930
rect 1627 2926 1767 2930
rect 1771 2926 1791 2930
rect 103 2925 1791 2926
rect 1797 2925 1798 2931
rect 1778 2897 1779 2903
rect 1785 2902 3487 2903
rect 1785 2898 1807 2902
rect 1811 2898 2055 2902
rect 2059 2898 2071 2902
rect 2075 2898 2143 2902
rect 2147 2898 2175 2902
rect 2179 2898 2231 2902
rect 2235 2898 2271 2902
rect 2275 2898 2319 2902
rect 2323 2898 2367 2902
rect 2371 2898 2407 2902
rect 2411 2898 2471 2902
rect 2475 2898 2495 2902
rect 2499 2898 2575 2902
rect 2579 2898 2583 2902
rect 2587 2898 2671 2902
rect 2675 2898 2679 2902
rect 2683 2898 2759 2902
rect 2763 2898 2783 2902
rect 2787 2898 2847 2902
rect 2851 2898 3463 2902
rect 3467 2898 3487 2902
rect 1785 2897 3487 2898
rect 3493 2897 3494 2903
rect 84 2857 85 2863
rect 91 2862 1779 2863
rect 91 2858 111 2862
rect 115 2858 135 2862
rect 139 2858 255 2862
rect 259 2858 263 2862
rect 267 2858 407 2862
rect 411 2858 431 2862
rect 435 2858 567 2862
rect 571 2858 607 2862
rect 611 2858 727 2862
rect 731 2858 783 2862
rect 787 2858 879 2862
rect 883 2858 951 2862
rect 955 2858 1023 2862
rect 1027 2858 1111 2862
rect 1115 2858 1167 2862
rect 1171 2858 1271 2862
rect 1275 2858 1311 2862
rect 1315 2858 1431 2862
rect 1435 2858 1463 2862
rect 1467 2858 1591 2862
rect 1595 2858 1767 2862
rect 1771 2858 1779 2862
rect 91 2857 1779 2858
rect 1785 2857 1786 2863
rect 1790 2829 1791 2835
rect 1797 2834 3499 2835
rect 1797 2830 1807 2834
rect 1811 2830 1983 2834
rect 1987 2830 2071 2834
rect 2075 2830 2111 2834
rect 2115 2830 2175 2834
rect 2179 2830 2239 2834
rect 2243 2830 2271 2834
rect 2275 2830 2367 2834
rect 2371 2830 2471 2834
rect 2475 2830 2487 2834
rect 2491 2830 2575 2834
rect 2579 2830 2607 2834
rect 2611 2830 2679 2834
rect 2683 2830 2719 2834
rect 2723 2830 2783 2834
rect 2787 2830 2839 2834
rect 2843 2830 2959 2834
rect 2963 2830 3463 2834
rect 3467 2830 3499 2834
rect 1797 2829 3499 2830
rect 3505 2829 3506 2835
rect 96 2785 97 2791
rect 103 2790 1791 2791
rect 103 2786 111 2790
rect 115 2786 135 2790
rect 139 2786 255 2790
rect 259 2786 287 2790
rect 291 2786 391 2790
rect 395 2786 407 2790
rect 411 2786 503 2790
rect 507 2786 567 2790
rect 571 2786 623 2790
rect 627 2786 727 2790
rect 731 2786 743 2790
rect 747 2786 855 2790
rect 859 2786 879 2790
rect 883 2786 967 2790
rect 971 2786 1023 2790
rect 1027 2786 1079 2790
rect 1083 2786 1167 2790
rect 1171 2786 1199 2790
rect 1203 2786 1311 2790
rect 1315 2786 1319 2790
rect 1323 2786 1463 2790
rect 1467 2786 1767 2790
rect 1771 2786 1791 2790
rect 103 2785 1791 2786
rect 1797 2785 1798 2791
rect 1778 2761 1779 2767
rect 1785 2766 3487 2767
rect 1785 2762 1807 2766
rect 1811 2762 1887 2766
rect 1891 2762 1983 2766
rect 1987 2762 2031 2766
rect 2035 2762 2111 2766
rect 2115 2762 2183 2766
rect 2187 2762 2239 2766
rect 2243 2762 2335 2766
rect 2339 2762 2367 2766
rect 2371 2762 2479 2766
rect 2483 2762 2487 2766
rect 2491 2762 2607 2766
rect 2611 2762 2623 2766
rect 2627 2762 2719 2766
rect 2723 2762 2767 2766
rect 2771 2762 2839 2766
rect 2843 2762 2911 2766
rect 2915 2762 2959 2766
rect 2963 2762 3055 2766
rect 3059 2762 3463 2766
rect 3467 2762 3487 2766
rect 1785 2761 3487 2762
rect 3493 2761 3494 2767
rect 84 2717 85 2723
rect 91 2722 1779 2723
rect 91 2718 111 2722
rect 115 2718 287 2722
rect 291 2718 391 2722
rect 395 2718 479 2722
rect 483 2718 503 2722
rect 507 2718 567 2722
rect 571 2718 623 2722
rect 627 2718 655 2722
rect 659 2718 743 2722
rect 747 2718 831 2722
rect 835 2718 855 2722
rect 859 2718 919 2722
rect 923 2718 967 2722
rect 971 2718 1007 2722
rect 1011 2718 1079 2722
rect 1083 2718 1095 2722
rect 1099 2718 1183 2722
rect 1187 2718 1199 2722
rect 1203 2718 1319 2722
rect 1323 2718 1767 2722
rect 1771 2718 1779 2722
rect 91 2717 1779 2718
rect 1785 2717 1786 2723
rect 1790 2697 1791 2703
rect 1797 2702 3499 2703
rect 1797 2698 1807 2702
rect 1811 2698 1831 2702
rect 1835 2698 1887 2702
rect 1891 2698 2023 2702
rect 2027 2698 2031 2702
rect 2035 2698 2183 2702
rect 2187 2698 2231 2702
rect 2235 2698 2335 2702
rect 2339 2698 2431 2702
rect 2435 2698 2479 2702
rect 2483 2698 2615 2702
rect 2619 2698 2623 2702
rect 2627 2698 2767 2702
rect 2771 2698 2783 2702
rect 2787 2698 2911 2702
rect 2915 2698 2943 2702
rect 2947 2698 3055 2702
rect 3059 2698 3095 2702
rect 3099 2698 3239 2702
rect 3243 2698 3367 2702
rect 3371 2698 3463 2702
rect 3467 2698 3499 2702
rect 1797 2697 3499 2698
rect 3505 2697 3506 2703
rect 96 2645 97 2651
rect 103 2650 1791 2651
rect 103 2646 111 2650
rect 115 2646 471 2650
rect 475 2646 479 2650
rect 483 2646 559 2650
rect 563 2646 567 2650
rect 571 2646 647 2650
rect 651 2646 655 2650
rect 659 2646 735 2650
rect 739 2646 743 2650
rect 747 2646 823 2650
rect 827 2646 831 2650
rect 835 2646 911 2650
rect 915 2646 919 2650
rect 923 2646 999 2650
rect 1003 2646 1007 2650
rect 1011 2646 1087 2650
rect 1091 2646 1095 2650
rect 1099 2646 1183 2650
rect 1187 2646 1767 2650
rect 1771 2646 1791 2650
rect 103 2645 1791 2646
rect 1797 2645 1798 2651
rect 1778 2629 1779 2635
rect 1785 2634 3487 2635
rect 1785 2630 1807 2634
rect 1811 2630 1831 2634
rect 1835 2630 1999 2634
rect 2003 2630 2023 2634
rect 2027 2630 2183 2634
rect 2187 2630 2231 2634
rect 2235 2630 2359 2634
rect 2363 2630 2431 2634
rect 2435 2630 2519 2634
rect 2523 2630 2615 2634
rect 2619 2630 2671 2634
rect 2675 2630 2783 2634
rect 2787 2630 2807 2634
rect 2811 2630 2927 2634
rect 2931 2630 2943 2634
rect 2947 2630 3047 2634
rect 3051 2630 3095 2634
rect 3099 2630 3159 2634
rect 3163 2630 3239 2634
rect 3243 2630 3271 2634
rect 3275 2630 3367 2634
rect 3371 2630 3463 2634
rect 3467 2630 3487 2634
rect 1785 2629 3487 2630
rect 3493 2629 3494 2635
rect 84 2569 85 2575
rect 91 2574 1779 2575
rect 91 2570 111 2574
rect 115 2570 223 2574
rect 227 2570 311 2574
rect 315 2570 407 2574
rect 411 2570 471 2574
rect 475 2570 503 2574
rect 507 2570 559 2574
rect 563 2570 591 2574
rect 595 2570 647 2574
rect 651 2570 679 2574
rect 683 2570 735 2574
rect 739 2570 767 2574
rect 771 2570 823 2574
rect 827 2570 855 2574
rect 859 2570 911 2574
rect 915 2570 943 2574
rect 947 2570 999 2574
rect 1003 2570 1031 2574
rect 1035 2570 1087 2574
rect 1091 2570 1119 2574
rect 1123 2570 1215 2574
rect 1219 2570 1311 2574
rect 1315 2570 1407 2574
rect 1411 2570 1495 2574
rect 1499 2570 1583 2574
rect 1587 2570 1671 2574
rect 1675 2570 1767 2574
rect 1771 2570 1779 2574
rect 91 2569 1779 2570
rect 1785 2569 1786 2575
rect 1790 2557 1791 2563
rect 1797 2562 3499 2563
rect 1797 2558 1807 2562
rect 1811 2558 1831 2562
rect 1835 2558 1999 2562
rect 2003 2558 2183 2562
rect 2187 2558 2207 2562
rect 2211 2558 2359 2562
rect 2363 2558 2519 2562
rect 2523 2558 2671 2562
rect 2675 2558 2799 2562
rect 2803 2558 2807 2562
rect 2811 2558 2927 2562
rect 2931 2558 3047 2562
rect 3051 2558 3159 2562
rect 3163 2558 3271 2562
rect 3275 2558 3367 2562
rect 3371 2558 3463 2562
rect 3467 2558 3499 2562
rect 1797 2557 3499 2558
rect 3505 2557 3506 2563
rect 96 2505 97 2511
rect 103 2510 1791 2511
rect 103 2506 111 2510
rect 115 2506 135 2510
rect 139 2506 223 2510
rect 227 2506 247 2510
rect 251 2506 311 2510
rect 315 2506 391 2510
rect 395 2506 407 2510
rect 411 2506 503 2510
rect 507 2506 543 2510
rect 547 2506 591 2510
rect 595 2506 679 2510
rect 683 2506 695 2510
rect 699 2506 767 2510
rect 771 2506 839 2510
rect 843 2506 855 2510
rect 859 2506 943 2510
rect 947 2506 975 2510
rect 979 2506 1031 2510
rect 1035 2506 1103 2510
rect 1107 2506 1119 2510
rect 1123 2506 1215 2510
rect 1219 2506 1231 2510
rect 1235 2506 1311 2510
rect 1315 2506 1351 2510
rect 1355 2506 1407 2510
rect 1411 2506 1463 2510
rect 1467 2506 1495 2510
rect 1499 2506 1575 2510
rect 1579 2506 1583 2510
rect 1587 2506 1671 2510
rect 1675 2506 1767 2510
rect 1771 2506 1791 2510
rect 103 2505 1791 2506
rect 1797 2505 1798 2511
rect 1778 2477 1779 2483
rect 1785 2482 3487 2483
rect 1785 2478 1807 2482
rect 1811 2478 2015 2482
rect 2019 2478 2199 2482
rect 2203 2478 2207 2482
rect 2211 2478 2367 2482
rect 2371 2478 2527 2482
rect 2531 2478 2671 2482
rect 2675 2478 2799 2482
rect 2803 2478 2807 2482
rect 2811 2478 2927 2482
rect 2931 2478 3047 2482
rect 3051 2478 3159 2482
rect 3163 2478 3271 2482
rect 3275 2478 3367 2482
rect 3371 2478 3463 2482
rect 3467 2478 3487 2482
rect 1785 2477 3487 2478
rect 3493 2477 3494 2483
rect 84 2425 85 2431
rect 91 2430 1779 2431
rect 91 2426 111 2430
rect 115 2426 135 2430
rect 139 2426 239 2430
rect 243 2426 247 2430
rect 251 2426 391 2430
rect 395 2426 543 2430
rect 547 2426 551 2430
rect 555 2426 695 2430
rect 699 2426 719 2430
rect 723 2426 839 2430
rect 843 2426 895 2430
rect 899 2426 975 2430
rect 979 2426 1063 2430
rect 1067 2426 1103 2430
rect 1107 2426 1231 2430
rect 1235 2426 1239 2430
rect 1243 2426 1351 2430
rect 1355 2426 1415 2430
rect 1419 2426 1463 2430
rect 1467 2426 1575 2430
rect 1579 2426 1591 2430
rect 1595 2426 1671 2430
rect 1675 2426 1767 2430
rect 1771 2426 1779 2430
rect 91 2425 1779 2426
rect 1785 2425 1786 2431
rect 1790 2409 1791 2415
rect 1797 2414 3499 2415
rect 1797 2410 1807 2414
rect 1811 2410 1839 2414
rect 1843 2410 2007 2414
rect 2011 2410 2015 2414
rect 2019 2410 2183 2414
rect 2187 2410 2199 2414
rect 2203 2410 2367 2414
rect 2371 2410 2527 2414
rect 2531 2410 2559 2414
rect 2563 2410 2671 2414
rect 2675 2410 2759 2414
rect 2763 2410 2807 2414
rect 2811 2410 2927 2414
rect 2931 2410 2967 2414
rect 2971 2410 3047 2414
rect 3051 2410 3159 2414
rect 3163 2410 3175 2414
rect 3179 2410 3271 2414
rect 3275 2410 3367 2414
rect 3371 2410 3463 2414
rect 3467 2410 3499 2414
rect 1797 2409 3499 2410
rect 3505 2409 3506 2415
rect 1778 2363 1779 2369
rect 1785 2363 1810 2369
rect 96 2353 97 2359
rect 103 2358 1791 2359
rect 103 2354 111 2358
rect 115 2354 135 2358
rect 139 2354 239 2358
rect 243 2354 375 2358
rect 379 2354 391 2358
rect 395 2354 479 2358
rect 483 2354 551 2358
rect 555 2354 599 2358
rect 603 2354 719 2358
rect 723 2354 847 2358
rect 851 2354 895 2358
rect 899 2354 975 2358
rect 979 2354 1063 2358
rect 1067 2354 1103 2358
rect 1107 2354 1239 2358
rect 1243 2354 1375 2358
rect 1379 2354 1415 2358
rect 1419 2354 1511 2358
rect 1515 2354 1591 2358
rect 1595 2354 1767 2358
rect 1771 2354 1791 2358
rect 103 2353 1791 2354
rect 1797 2353 1798 2359
rect 1804 2351 1810 2363
rect 1804 2350 3487 2351
rect 1804 2346 1807 2350
rect 1811 2346 1839 2350
rect 1843 2346 1887 2350
rect 1891 2346 2007 2350
rect 2011 2346 2015 2350
rect 2019 2346 2151 2350
rect 2155 2346 2183 2350
rect 2187 2346 2303 2350
rect 2307 2346 2367 2350
rect 2371 2346 2463 2350
rect 2467 2346 2559 2350
rect 2563 2346 2647 2350
rect 2651 2346 2759 2350
rect 2763 2346 2839 2350
rect 2843 2346 2967 2350
rect 2971 2346 3047 2350
rect 3051 2346 3175 2350
rect 3179 2346 3255 2350
rect 3259 2346 3367 2350
rect 3371 2346 3463 2350
rect 3467 2346 3487 2350
rect 1804 2345 3487 2346
rect 3493 2345 3494 2351
rect 84 2281 85 2287
rect 91 2286 1779 2287
rect 91 2282 111 2286
rect 115 2282 375 2286
rect 379 2282 479 2286
rect 483 2282 575 2286
rect 579 2282 599 2286
rect 603 2282 663 2286
rect 667 2282 719 2286
rect 723 2282 759 2286
rect 763 2282 847 2286
rect 851 2282 863 2286
rect 867 2282 967 2286
rect 971 2282 975 2286
rect 979 2282 1079 2286
rect 1083 2282 1103 2286
rect 1107 2282 1191 2286
rect 1195 2282 1239 2286
rect 1243 2282 1303 2286
rect 1307 2282 1375 2286
rect 1379 2282 1415 2286
rect 1419 2282 1511 2286
rect 1515 2282 1767 2286
rect 1771 2282 1779 2286
rect 91 2281 1779 2282
rect 1785 2281 1786 2287
rect 1790 2277 1791 2283
rect 1797 2282 3499 2283
rect 1797 2278 1807 2282
rect 1811 2278 1887 2282
rect 1891 2278 2015 2282
rect 2019 2278 2039 2282
rect 2043 2278 2135 2282
rect 2139 2278 2151 2282
rect 2155 2278 2239 2282
rect 2243 2278 2303 2282
rect 2307 2278 2343 2282
rect 2347 2278 2463 2282
rect 2467 2278 2591 2282
rect 2595 2278 2647 2282
rect 2651 2278 2735 2282
rect 2739 2278 2839 2282
rect 2843 2278 2887 2282
rect 2891 2278 3047 2282
rect 3051 2278 3215 2282
rect 3219 2278 3255 2282
rect 3259 2278 3367 2282
rect 3371 2278 3463 2282
rect 3467 2278 3499 2282
rect 1797 2277 3499 2278
rect 3505 2277 3506 2283
rect 96 2217 97 2223
rect 103 2222 1791 2223
rect 103 2218 111 2222
rect 115 2218 439 2222
rect 443 2218 527 2222
rect 531 2218 575 2222
rect 579 2218 615 2222
rect 619 2218 663 2222
rect 667 2218 703 2222
rect 707 2218 759 2222
rect 763 2218 791 2222
rect 795 2218 863 2222
rect 867 2218 879 2222
rect 883 2218 967 2222
rect 971 2218 1055 2222
rect 1059 2218 1079 2222
rect 1083 2218 1143 2222
rect 1147 2218 1191 2222
rect 1195 2218 1231 2222
rect 1235 2218 1303 2222
rect 1307 2218 1319 2222
rect 1323 2218 1415 2222
rect 1419 2218 1767 2222
rect 1771 2218 1791 2222
rect 103 2217 1791 2218
rect 1797 2217 1798 2223
rect 1778 2201 1779 2207
rect 1785 2206 3487 2207
rect 1785 2202 1807 2206
rect 1811 2202 2039 2206
rect 2043 2202 2135 2206
rect 2139 2202 2183 2206
rect 2187 2202 2239 2206
rect 2243 2202 2279 2206
rect 2283 2202 2343 2206
rect 2347 2202 2383 2206
rect 2387 2202 2463 2206
rect 2467 2202 2495 2206
rect 2499 2202 2591 2206
rect 2595 2202 2607 2206
rect 2611 2202 2719 2206
rect 2723 2202 2735 2206
rect 2739 2202 2839 2206
rect 2843 2202 2887 2206
rect 2891 2202 2967 2206
rect 2971 2202 3047 2206
rect 3051 2202 3103 2206
rect 3107 2202 3215 2206
rect 3219 2202 3247 2206
rect 3251 2202 3367 2206
rect 3371 2202 3463 2206
rect 3467 2202 3487 2206
rect 1785 2201 3487 2202
rect 3493 2201 3494 2207
rect 84 2137 85 2143
rect 91 2142 1779 2143
rect 91 2138 111 2142
rect 115 2138 303 2142
rect 307 2138 407 2142
rect 411 2138 439 2142
rect 443 2138 519 2142
rect 523 2138 527 2142
rect 531 2138 615 2142
rect 619 2138 631 2142
rect 635 2138 703 2142
rect 707 2138 743 2142
rect 747 2138 791 2142
rect 795 2138 863 2142
rect 867 2138 879 2142
rect 883 2138 967 2142
rect 971 2138 983 2142
rect 987 2138 1055 2142
rect 1059 2138 1143 2142
rect 1147 2138 1231 2142
rect 1235 2138 1319 2142
rect 1323 2138 1767 2142
rect 1771 2138 1779 2142
rect 91 2137 1779 2138
rect 1785 2137 1786 2143
rect 1790 2129 1791 2135
rect 1797 2134 3499 2135
rect 1797 2130 1807 2134
rect 1811 2130 2135 2134
rect 2139 2130 2183 2134
rect 2187 2130 2255 2134
rect 2259 2130 2279 2134
rect 2283 2130 2383 2134
rect 2387 2130 2495 2134
rect 2499 2130 2519 2134
rect 2523 2130 2607 2134
rect 2611 2130 2655 2134
rect 2659 2130 2719 2134
rect 2723 2130 2783 2134
rect 2787 2130 2839 2134
rect 2843 2130 2911 2134
rect 2915 2130 2967 2134
rect 2971 2130 3031 2134
rect 3035 2130 3103 2134
rect 3107 2130 3151 2134
rect 3155 2130 3247 2134
rect 3251 2130 3271 2134
rect 3275 2130 3367 2134
rect 3371 2130 3463 2134
rect 3467 2130 3499 2134
rect 1797 2129 3499 2130
rect 3505 2129 3506 2135
rect 96 2073 97 2079
rect 103 2078 1791 2079
rect 103 2074 111 2078
rect 115 2074 255 2078
rect 259 2074 303 2078
rect 307 2074 375 2078
rect 379 2074 407 2078
rect 411 2074 495 2078
rect 499 2074 519 2078
rect 523 2074 615 2078
rect 619 2074 631 2078
rect 635 2074 727 2078
rect 731 2074 743 2078
rect 747 2074 831 2078
rect 835 2074 863 2078
rect 867 2074 935 2078
rect 939 2074 983 2078
rect 987 2074 1039 2078
rect 1043 2074 1143 2078
rect 1147 2074 1255 2078
rect 1259 2074 1767 2078
rect 1771 2074 1791 2078
rect 103 2073 1791 2074
rect 1797 2073 1798 2079
rect 1778 2057 1779 2063
rect 1785 2062 3487 2063
rect 1785 2058 1807 2062
rect 1811 2058 2135 2062
rect 2139 2058 2247 2062
rect 2251 2058 2255 2062
rect 2259 2058 2383 2062
rect 2387 2058 2415 2062
rect 2419 2058 2519 2062
rect 2523 2058 2575 2062
rect 2579 2058 2655 2062
rect 2659 2058 2727 2062
rect 2731 2058 2783 2062
rect 2787 2058 2871 2062
rect 2875 2058 2911 2062
rect 2915 2058 3007 2062
rect 3011 2058 3031 2062
rect 3035 2058 3135 2062
rect 3139 2058 3151 2062
rect 3155 2058 3263 2062
rect 3267 2058 3271 2062
rect 3275 2058 3367 2062
rect 3371 2058 3463 2062
rect 3467 2058 3487 2062
rect 1785 2057 3487 2058
rect 3493 2057 3494 2063
rect 84 2009 85 2015
rect 91 2014 1779 2015
rect 91 2010 111 2014
rect 115 2010 255 2014
rect 259 2010 359 2014
rect 363 2010 375 2014
rect 379 2010 487 2014
rect 491 2010 495 2014
rect 499 2010 615 2014
rect 619 2010 623 2014
rect 627 2010 727 2014
rect 731 2010 759 2014
rect 763 2010 831 2014
rect 835 2010 895 2014
rect 899 2010 935 2014
rect 939 2010 1023 2014
rect 1027 2010 1039 2014
rect 1043 2010 1143 2014
rect 1147 2010 1151 2014
rect 1155 2010 1255 2014
rect 1259 2010 1271 2014
rect 1275 2010 1399 2014
rect 1403 2010 1527 2014
rect 1531 2010 1767 2014
rect 1771 2010 1779 2014
rect 91 2009 1779 2010
rect 1785 2009 1786 2015
rect 1790 1977 1791 1983
rect 1797 1982 3499 1983
rect 1797 1978 1807 1982
rect 1811 1978 1831 1982
rect 1835 1978 1919 1982
rect 1923 1978 2047 1982
rect 2051 1978 2183 1982
rect 2187 1978 2247 1982
rect 2251 1978 2327 1982
rect 2331 1978 2415 1982
rect 2419 1978 2471 1982
rect 2475 1978 2575 1982
rect 2579 1978 2615 1982
rect 2619 1978 2727 1982
rect 2731 1978 2751 1982
rect 2755 1978 2871 1982
rect 2875 1978 2887 1982
rect 2891 1978 3007 1982
rect 3011 1978 3031 1982
rect 3035 1978 3135 1982
rect 3139 1978 3175 1982
rect 3179 1978 3263 1982
rect 3267 1978 3319 1982
rect 3323 1978 3367 1982
rect 3371 1978 3463 1982
rect 3467 1978 3499 1982
rect 1797 1977 3499 1978
rect 3505 1977 3506 1983
rect 96 1945 97 1951
rect 103 1950 1791 1951
rect 103 1946 111 1950
rect 115 1946 359 1950
rect 363 1946 447 1950
rect 451 1946 487 1950
rect 491 1946 575 1950
rect 579 1946 623 1950
rect 627 1946 711 1950
rect 715 1946 759 1950
rect 763 1946 847 1950
rect 851 1946 895 1950
rect 899 1946 983 1950
rect 987 1946 1023 1950
rect 1027 1946 1119 1950
rect 1123 1946 1151 1950
rect 1155 1946 1255 1950
rect 1259 1946 1271 1950
rect 1275 1946 1383 1950
rect 1387 1946 1399 1950
rect 1403 1946 1519 1950
rect 1523 1946 1527 1950
rect 1531 1946 1655 1950
rect 1659 1946 1767 1950
rect 1771 1946 1791 1950
rect 103 1945 1791 1946
rect 1797 1945 1798 1951
rect 1778 1909 1779 1915
rect 1785 1914 3487 1915
rect 1785 1910 1807 1914
rect 1811 1910 1831 1914
rect 1835 1910 1919 1914
rect 1923 1910 2039 1914
rect 2043 1910 2047 1914
rect 2051 1910 2167 1914
rect 2171 1910 2183 1914
rect 2187 1910 2303 1914
rect 2307 1910 2327 1914
rect 2331 1910 2455 1914
rect 2459 1910 2471 1914
rect 2475 1910 2615 1914
rect 2619 1910 2751 1914
rect 2755 1910 2791 1914
rect 2795 1910 2887 1914
rect 2891 1910 2983 1914
rect 2987 1910 3031 1914
rect 3035 1910 3175 1914
rect 3179 1910 3183 1914
rect 3187 1910 3319 1914
rect 3323 1910 3367 1914
rect 3371 1910 3463 1914
rect 3467 1910 3487 1914
rect 1785 1909 3487 1910
rect 3493 1909 3494 1915
rect 84 1881 85 1887
rect 91 1886 1779 1887
rect 91 1882 111 1886
rect 115 1882 447 1886
rect 451 1882 559 1886
rect 563 1882 575 1886
rect 579 1882 695 1886
rect 699 1882 711 1886
rect 715 1882 831 1886
rect 835 1882 847 1886
rect 851 1882 959 1886
rect 963 1882 983 1886
rect 987 1882 1079 1886
rect 1083 1882 1119 1886
rect 1123 1882 1199 1886
rect 1203 1882 1255 1886
rect 1259 1882 1327 1886
rect 1331 1882 1383 1886
rect 1387 1882 1455 1886
rect 1459 1882 1519 1886
rect 1523 1882 1655 1886
rect 1659 1882 1767 1886
rect 1771 1882 1779 1886
rect 91 1881 1779 1882
rect 1785 1881 1786 1887
rect 1790 1841 1791 1847
rect 1797 1846 3499 1847
rect 1797 1842 1807 1846
rect 1811 1842 1831 1846
rect 1835 1842 1919 1846
rect 1923 1842 1959 1846
rect 1963 1842 2039 1846
rect 2043 1842 2111 1846
rect 2115 1842 2167 1846
rect 2171 1842 2255 1846
rect 2259 1842 2303 1846
rect 2307 1842 2407 1846
rect 2411 1842 2455 1846
rect 2459 1842 2567 1846
rect 2571 1842 2615 1846
rect 2619 1842 2743 1846
rect 2747 1842 2791 1846
rect 2795 1842 2935 1846
rect 2939 1842 2983 1846
rect 2987 1842 3135 1846
rect 3139 1842 3183 1846
rect 3187 1842 3343 1846
rect 3347 1842 3367 1846
rect 3371 1842 3463 1846
rect 3467 1842 3499 1846
rect 1797 1841 3499 1842
rect 3505 1841 3506 1847
rect 96 1809 97 1815
rect 103 1814 1791 1815
rect 103 1810 111 1814
rect 115 1810 135 1814
rect 139 1810 223 1814
rect 227 1810 311 1814
rect 315 1810 407 1814
rect 411 1810 527 1814
rect 531 1810 559 1814
rect 563 1810 655 1814
rect 659 1810 695 1814
rect 699 1810 799 1814
rect 803 1810 831 1814
rect 835 1810 943 1814
rect 947 1810 959 1814
rect 963 1810 1079 1814
rect 1083 1810 1087 1814
rect 1091 1810 1199 1814
rect 1203 1810 1239 1814
rect 1243 1810 1327 1814
rect 1331 1810 1391 1814
rect 1395 1810 1455 1814
rect 1459 1810 1543 1814
rect 1547 1810 1671 1814
rect 1675 1810 1767 1814
rect 1771 1810 1791 1814
rect 103 1809 1791 1810
rect 1797 1809 1798 1815
rect 1778 1765 1779 1771
rect 1785 1770 3487 1771
rect 1785 1766 1807 1770
rect 1811 1766 1831 1770
rect 1835 1766 1879 1770
rect 1883 1766 1959 1770
rect 1963 1766 2015 1770
rect 2019 1766 2111 1770
rect 2115 1766 2151 1770
rect 2155 1766 2255 1770
rect 2259 1766 2303 1770
rect 2307 1766 2407 1770
rect 2411 1766 2479 1770
rect 2483 1766 2567 1770
rect 2571 1766 2687 1770
rect 2691 1766 2743 1770
rect 2747 1766 2911 1770
rect 2915 1766 2935 1770
rect 2939 1766 3135 1770
rect 3139 1766 3151 1770
rect 3155 1766 3343 1770
rect 3347 1766 3367 1770
rect 3371 1766 3463 1770
rect 3467 1766 3487 1770
rect 1785 1765 3487 1766
rect 3493 1765 3494 1771
rect 84 1733 85 1739
rect 91 1738 1779 1739
rect 91 1734 111 1738
rect 115 1734 135 1738
rect 139 1734 223 1738
rect 227 1734 247 1738
rect 251 1734 311 1738
rect 315 1734 399 1738
rect 403 1734 407 1738
rect 411 1734 527 1738
rect 531 1734 567 1738
rect 571 1734 655 1738
rect 659 1734 751 1738
rect 755 1734 799 1738
rect 803 1734 935 1738
rect 939 1734 943 1738
rect 947 1734 1087 1738
rect 1091 1734 1119 1738
rect 1123 1734 1239 1738
rect 1243 1734 1311 1738
rect 1315 1734 1391 1738
rect 1395 1734 1503 1738
rect 1507 1734 1543 1738
rect 1547 1734 1671 1738
rect 1675 1734 1767 1738
rect 1771 1734 1779 1738
rect 91 1733 1779 1734
rect 1785 1733 1786 1739
rect 1790 1693 1791 1699
rect 1797 1698 3499 1699
rect 1797 1694 1807 1698
rect 1811 1694 1831 1698
rect 1835 1694 1879 1698
rect 1883 1694 1935 1698
rect 1939 1694 2015 1698
rect 2019 1694 2063 1698
rect 2067 1694 2151 1698
rect 2155 1694 2183 1698
rect 2187 1694 2303 1698
rect 2307 1694 2311 1698
rect 2315 1694 2439 1698
rect 2443 1694 2479 1698
rect 2483 1694 2575 1698
rect 2579 1694 2687 1698
rect 2691 1694 2727 1698
rect 2731 1694 2887 1698
rect 2891 1694 2911 1698
rect 2915 1694 3047 1698
rect 3051 1694 3151 1698
rect 3155 1694 3215 1698
rect 3219 1694 3367 1698
rect 3371 1694 3463 1698
rect 3467 1694 3499 1698
rect 1797 1693 3499 1694
rect 3505 1693 3506 1699
rect 96 1665 97 1671
rect 103 1670 1791 1671
rect 103 1666 111 1670
rect 115 1666 135 1670
rect 139 1666 191 1670
rect 195 1666 247 1670
rect 251 1666 295 1670
rect 299 1666 399 1670
rect 403 1666 407 1670
rect 411 1666 535 1670
rect 539 1666 567 1670
rect 571 1666 687 1670
rect 691 1666 751 1670
rect 755 1666 855 1670
rect 859 1666 935 1670
rect 939 1666 1039 1670
rect 1043 1666 1119 1670
rect 1123 1666 1231 1670
rect 1235 1666 1311 1670
rect 1315 1666 1431 1670
rect 1435 1666 1503 1670
rect 1507 1666 1639 1670
rect 1643 1666 1671 1670
rect 1675 1666 1767 1670
rect 1771 1666 1791 1670
rect 103 1665 1791 1666
rect 1797 1665 1798 1671
rect 1778 1621 1779 1627
rect 1785 1626 3487 1627
rect 1785 1622 1807 1626
rect 1811 1622 1831 1626
rect 1835 1622 1935 1626
rect 1939 1622 1943 1626
rect 1947 1622 2063 1626
rect 2067 1622 2087 1626
rect 2091 1622 2183 1626
rect 2187 1622 2231 1626
rect 2235 1622 2311 1626
rect 2315 1622 2367 1626
rect 2371 1622 2439 1626
rect 2443 1622 2503 1626
rect 2507 1622 2575 1626
rect 2579 1622 2639 1626
rect 2643 1622 2727 1626
rect 2731 1622 2767 1626
rect 2771 1622 2887 1626
rect 2891 1622 2895 1626
rect 2899 1622 3015 1626
rect 3019 1622 3047 1626
rect 3051 1622 3135 1626
rect 3139 1622 3215 1626
rect 3219 1622 3263 1626
rect 3267 1622 3367 1626
rect 3371 1622 3463 1626
rect 3467 1622 3487 1626
rect 1785 1621 3487 1622
rect 3493 1621 3494 1627
rect 84 1597 85 1603
rect 91 1602 1779 1603
rect 91 1598 111 1602
rect 115 1598 191 1602
rect 195 1598 295 1602
rect 299 1598 327 1602
rect 331 1598 407 1602
rect 411 1598 431 1602
rect 435 1598 535 1602
rect 539 1598 543 1602
rect 547 1598 671 1602
rect 675 1598 687 1602
rect 691 1598 815 1602
rect 819 1598 855 1602
rect 859 1598 967 1602
rect 971 1598 1039 1602
rect 1043 1598 1119 1602
rect 1123 1598 1231 1602
rect 1235 1598 1279 1602
rect 1283 1598 1431 1602
rect 1435 1598 1439 1602
rect 1443 1598 1607 1602
rect 1611 1598 1639 1602
rect 1643 1598 1767 1602
rect 1771 1598 1779 1602
rect 91 1597 1779 1598
rect 1785 1597 1786 1603
rect 1790 1549 1791 1555
rect 1797 1554 3499 1555
rect 1797 1550 1807 1554
rect 1811 1550 1831 1554
rect 1835 1550 1839 1554
rect 1843 1550 1943 1554
rect 1947 1550 1991 1554
rect 1995 1550 2087 1554
rect 2091 1550 2151 1554
rect 2155 1550 2231 1554
rect 2235 1550 2303 1554
rect 2307 1550 2367 1554
rect 2371 1550 2455 1554
rect 2459 1550 2503 1554
rect 2507 1550 2599 1554
rect 2603 1550 2639 1554
rect 2643 1550 2735 1554
rect 2739 1550 2767 1554
rect 2771 1550 2871 1554
rect 2875 1550 2895 1554
rect 2899 1550 3007 1554
rect 3011 1550 3015 1554
rect 3019 1550 3135 1554
rect 3139 1550 3143 1554
rect 3147 1550 3263 1554
rect 3267 1550 3367 1554
rect 3371 1550 3463 1554
rect 3467 1550 3499 1554
rect 1797 1549 3499 1550
rect 3505 1549 3506 1555
rect 96 1529 97 1535
rect 103 1534 1791 1535
rect 103 1530 111 1534
rect 115 1530 223 1534
rect 227 1530 327 1534
rect 331 1530 343 1534
rect 347 1530 431 1534
rect 435 1530 471 1534
rect 475 1530 543 1534
rect 547 1530 607 1534
rect 611 1530 671 1534
rect 675 1530 751 1534
rect 755 1530 815 1534
rect 819 1530 895 1534
rect 899 1530 967 1534
rect 971 1530 1047 1534
rect 1051 1530 1119 1534
rect 1123 1530 1199 1534
rect 1203 1530 1279 1534
rect 1283 1530 1351 1534
rect 1355 1530 1439 1534
rect 1443 1530 1503 1534
rect 1507 1530 1607 1534
rect 1611 1530 1767 1534
rect 1771 1530 1791 1534
rect 103 1529 1791 1530
rect 1797 1529 1798 1535
rect 1778 1477 1779 1483
rect 1785 1482 3487 1483
rect 1785 1478 1807 1482
rect 1811 1478 1839 1482
rect 1843 1478 1943 1482
rect 1947 1478 1991 1482
rect 1995 1478 2055 1482
rect 2059 1478 2151 1482
rect 2155 1478 2191 1482
rect 2195 1478 2303 1482
rect 2307 1478 2335 1482
rect 2339 1478 2455 1482
rect 2459 1478 2479 1482
rect 2483 1478 2599 1482
rect 2603 1478 2631 1482
rect 2635 1478 2735 1482
rect 2739 1478 2783 1482
rect 2787 1478 2871 1482
rect 2875 1478 2935 1482
rect 2939 1478 3007 1482
rect 3011 1478 3087 1482
rect 3091 1478 3143 1482
rect 3147 1478 3239 1482
rect 3243 1478 3463 1482
rect 3467 1478 3487 1482
rect 1785 1477 3487 1478
rect 3493 1477 3494 1483
rect 84 1457 85 1463
rect 91 1462 1779 1463
rect 91 1458 111 1462
rect 115 1458 135 1462
rect 139 1458 223 1462
rect 227 1458 303 1462
rect 307 1458 343 1462
rect 347 1458 471 1462
rect 475 1458 607 1462
rect 611 1458 631 1462
rect 635 1458 751 1462
rect 755 1458 783 1462
rect 787 1458 895 1462
rect 899 1458 927 1462
rect 931 1458 1047 1462
rect 1051 1458 1063 1462
rect 1067 1458 1199 1462
rect 1203 1458 1335 1462
rect 1339 1458 1351 1462
rect 1355 1458 1471 1462
rect 1475 1458 1503 1462
rect 1507 1458 1767 1462
rect 1771 1458 1779 1462
rect 91 1457 1779 1458
rect 1785 1457 1786 1463
rect 1790 1405 1791 1411
rect 1797 1410 3499 1411
rect 1797 1406 1807 1410
rect 1811 1406 1943 1410
rect 1947 1406 2055 1410
rect 2059 1406 2095 1410
rect 2099 1406 2191 1410
rect 2195 1406 2199 1410
rect 2203 1406 2319 1410
rect 2323 1406 2335 1410
rect 2339 1406 2455 1410
rect 2459 1406 2479 1410
rect 2483 1406 2599 1410
rect 2603 1406 2631 1410
rect 2635 1406 2743 1410
rect 2747 1406 2783 1410
rect 2787 1406 2887 1410
rect 2891 1406 2935 1410
rect 2939 1406 3031 1410
rect 3035 1406 3087 1410
rect 3091 1406 3175 1410
rect 3179 1406 3239 1410
rect 3243 1406 3327 1410
rect 3331 1406 3463 1410
rect 3467 1406 3499 1410
rect 1797 1405 3499 1406
rect 3505 1405 3506 1411
rect 96 1389 97 1395
rect 103 1394 1791 1395
rect 103 1390 111 1394
rect 115 1390 135 1394
rect 139 1390 279 1394
rect 283 1390 303 1394
rect 307 1390 447 1394
rect 451 1390 471 1394
rect 475 1390 607 1394
rect 611 1390 631 1394
rect 635 1390 759 1394
rect 763 1390 783 1394
rect 787 1390 903 1394
rect 907 1390 927 1394
rect 931 1390 1031 1394
rect 1035 1390 1063 1394
rect 1067 1390 1159 1394
rect 1163 1390 1199 1394
rect 1203 1390 1287 1394
rect 1291 1390 1335 1394
rect 1339 1390 1415 1394
rect 1419 1390 1471 1394
rect 1475 1390 1767 1394
rect 1771 1390 1791 1394
rect 103 1389 1791 1390
rect 1797 1389 1798 1395
rect 1778 1337 1779 1343
rect 1785 1342 3487 1343
rect 1785 1338 1807 1342
rect 1811 1338 2095 1342
rect 2099 1338 2103 1342
rect 2107 1338 2199 1342
rect 2203 1338 2239 1342
rect 2243 1338 2319 1342
rect 2323 1338 2383 1342
rect 2387 1338 2455 1342
rect 2459 1338 2535 1342
rect 2539 1338 2599 1342
rect 2603 1338 2687 1342
rect 2691 1338 2743 1342
rect 2747 1338 2839 1342
rect 2843 1338 2887 1342
rect 2891 1338 2991 1342
rect 2995 1338 3031 1342
rect 3035 1338 3143 1342
rect 3147 1338 3175 1342
rect 3179 1338 3303 1342
rect 3307 1338 3327 1342
rect 3331 1338 3463 1342
rect 3467 1338 3487 1342
rect 1785 1337 3487 1338
rect 3493 1337 3494 1343
rect 84 1321 85 1327
rect 91 1326 1779 1327
rect 91 1322 111 1326
rect 115 1322 135 1326
rect 139 1322 279 1326
rect 283 1322 439 1326
rect 443 1322 447 1326
rect 451 1322 583 1326
rect 587 1322 607 1326
rect 611 1322 719 1326
rect 723 1322 759 1326
rect 763 1322 847 1326
rect 851 1322 903 1326
rect 907 1322 967 1326
rect 971 1322 1031 1326
rect 1035 1322 1079 1326
rect 1083 1322 1159 1326
rect 1163 1322 1191 1326
rect 1195 1322 1287 1326
rect 1291 1322 1311 1326
rect 1315 1322 1415 1326
rect 1419 1322 1767 1326
rect 1771 1322 1779 1326
rect 91 1321 1779 1322
rect 1785 1321 1786 1327
rect 1790 1273 1791 1279
rect 1797 1278 3499 1279
rect 1797 1274 1807 1278
rect 1811 1274 1935 1278
rect 1939 1274 2063 1278
rect 2067 1274 2103 1278
rect 2107 1274 2199 1278
rect 2203 1274 2239 1278
rect 2243 1274 2343 1278
rect 2347 1274 2383 1278
rect 2387 1274 2495 1278
rect 2499 1274 2535 1278
rect 2539 1274 2655 1278
rect 2659 1274 2687 1278
rect 2691 1274 2815 1278
rect 2819 1274 2839 1278
rect 2843 1274 2975 1278
rect 2979 1274 2991 1278
rect 2995 1274 3143 1278
rect 3147 1274 3303 1278
rect 3307 1274 3463 1278
rect 3467 1274 3499 1278
rect 1797 1273 3499 1274
rect 3505 1273 3506 1279
rect 96 1253 97 1259
rect 103 1258 1791 1259
rect 103 1254 111 1258
rect 115 1254 135 1258
rect 139 1254 239 1258
rect 243 1254 279 1258
rect 283 1254 367 1258
rect 371 1254 439 1258
rect 443 1254 495 1258
rect 499 1254 583 1258
rect 587 1254 615 1258
rect 619 1254 719 1258
rect 723 1254 735 1258
rect 739 1254 847 1258
rect 851 1254 959 1258
rect 963 1254 967 1258
rect 971 1254 1071 1258
rect 1075 1254 1079 1258
rect 1083 1254 1191 1258
rect 1195 1254 1311 1258
rect 1315 1254 1767 1258
rect 1771 1254 1791 1258
rect 103 1253 1791 1254
rect 1797 1253 1798 1259
rect 1778 1209 1779 1215
rect 1785 1214 3487 1215
rect 1785 1210 1807 1214
rect 1811 1210 1831 1214
rect 1835 1210 1935 1214
rect 1939 1210 2063 1214
rect 2067 1210 2079 1214
rect 2083 1210 2199 1214
rect 2203 1210 2231 1214
rect 2235 1210 2343 1214
rect 2347 1210 2391 1214
rect 2395 1210 2495 1214
rect 2499 1210 2543 1214
rect 2547 1210 2655 1214
rect 2659 1210 2695 1214
rect 2699 1210 2815 1214
rect 2819 1210 2847 1214
rect 2851 1210 2975 1214
rect 2979 1210 2999 1214
rect 3003 1210 3143 1214
rect 3147 1210 3159 1214
rect 3163 1210 3463 1214
rect 3467 1210 3487 1214
rect 1785 1209 3487 1210
rect 3493 1209 3494 1215
rect 84 1185 85 1191
rect 91 1190 1779 1191
rect 91 1186 111 1190
rect 115 1186 135 1190
rect 139 1186 239 1190
rect 243 1186 367 1190
rect 371 1186 375 1190
rect 379 1186 495 1190
rect 499 1186 511 1190
rect 515 1186 615 1190
rect 619 1186 655 1190
rect 659 1186 735 1190
rect 739 1186 791 1190
rect 795 1186 847 1190
rect 851 1186 927 1190
rect 931 1186 959 1190
rect 963 1186 1063 1190
rect 1067 1186 1071 1190
rect 1075 1186 1191 1190
rect 1195 1186 1199 1190
rect 1203 1186 1335 1190
rect 1339 1186 1767 1190
rect 1771 1186 1779 1190
rect 91 1185 1779 1186
rect 1785 1185 1786 1191
rect 1790 1133 1791 1139
rect 1797 1138 3499 1139
rect 1797 1134 1807 1138
rect 1811 1134 1831 1138
rect 1835 1134 1863 1138
rect 1867 1134 1935 1138
rect 1939 1134 1983 1138
rect 1987 1134 2079 1138
rect 2083 1134 2111 1138
rect 2115 1134 2231 1138
rect 2235 1134 2247 1138
rect 2251 1134 2383 1138
rect 2387 1134 2391 1138
rect 2395 1134 2511 1138
rect 2515 1134 2543 1138
rect 2547 1134 2639 1138
rect 2643 1134 2695 1138
rect 2699 1134 2759 1138
rect 2763 1134 2847 1138
rect 2851 1134 2871 1138
rect 2875 1134 2975 1138
rect 2979 1134 2999 1138
rect 3003 1134 3079 1138
rect 3083 1134 3159 1138
rect 3163 1134 3183 1138
rect 3187 1134 3279 1138
rect 3283 1134 3367 1138
rect 3371 1134 3463 1138
rect 3467 1134 3499 1138
rect 1797 1133 3499 1134
rect 3505 1133 3506 1139
rect 96 1117 97 1123
rect 103 1122 1791 1123
rect 103 1118 111 1122
rect 115 1118 135 1122
rect 139 1118 191 1122
rect 195 1118 239 1122
rect 243 1118 335 1122
rect 339 1118 375 1122
rect 379 1118 495 1122
rect 499 1118 511 1122
rect 515 1118 655 1122
rect 659 1118 791 1122
rect 795 1118 815 1122
rect 819 1118 927 1122
rect 931 1118 967 1122
rect 971 1118 1063 1122
rect 1067 1118 1119 1122
rect 1123 1118 1199 1122
rect 1203 1118 1263 1122
rect 1267 1118 1335 1122
rect 1339 1118 1407 1122
rect 1411 1118 1559 1122
rect 1563 1118 1767 1122
rect 1771 1118 1791 1122
rect 103 1117 1791 1118
rect 1797 1117 1798 1123
rect 1778 1061 1779 1067
rect 1785 1066 3487 1067
rect 1785 1062 1807 1066
rect 1811 1062 1863 1066
rect 1867 1062 1983 1066
rect 1987 1062 2103 1066
rect 2107 1062 2111 1066
rect 2115 1062 2191 1066
rect 2195 1062 2247 1066
rect 2251 1062 2279 1066
rect 2283 1062 2367 1066
rect 2371 1062 2383 1066
rect 2387 1062 2455 1066
rect 2459 1062 2511 1066
rect 2515 1062 2543 1066
rect 2547 1062 2631 1066
rect 2635 1062 2639 1066
rect 2643 1062 2719 1066
rect 2723 1062 2759 1066
rect 2763 1062 2807 1066
rect 2811 1062 2871 1066
rect 2875 1062 2975 1066
rect 2979 1062 3079 1066
rect 3083 1062 3183 1066
rect 3187 1062 3279 1066
rect 3283 1062 3367 1066
rect 3371 1062 3463 1066
rect 3467 1062 3487 1066
rect 1785 1061 3487 1062
rect 3493 1061 3494 1067
rect 84 1045 85 1051
rect 91 1050 1779 1051
rect 91 1046 111 1050
rect 115 1046 191 1050
rect 195 1046 327 1050
rect 331 1046 335 1050
rect 339 1046 463 1050
rect 467 1046 495 1050
rect 499 1046 607 1050
rect 611 1046 655 1050
rect 659 1046 767 1050
rect 771 1046 815 1050
rect 819 1046 927 1050
rect 931 1046 967 1050
rect 971 1046 1079 1050
rect 1083 1046 1119 1050
rect 1123 1046 1231 1050
rect 1235 1046 1263 1050
rect 1267 1046 1383 1050
rect 1387 1046 1407 1050
rect 1411 1046 1535 1050
rect 1539 1046 1559 1050
rect 1563 1046 1671 1050
rect 1675 1046 1767 1050
rect 1771 1046 1779 1050
rect 91 1045 1779 1046
rect 1785 1045 1786 1051
rect 1790 997 1791 1003
rect 1797 1002 3499 1003
rect 1797 998 1807 1002
rect 1811 998 2103 1002
rect 2107 998 2191 1002
rect 2195 998 2279 1002
rect 2283 998 2311 1002
rect 2315 998 2367 1002
rect 2371 998 2407 1002
rect 2411 998 2455 1002
rect 2459 998 2511 1002
rect 2515 998 2543 1002
rect 2547 998 2623 1002
rect 2627 998 2631 1002
rect 2635 998 2719 1002
rect 2723 998 2751 1002
rect 2755 998 2807 1002
rect 2811 998 2895 1002
rect 2899 998 3055 1002
rect 3059 998 3223 1002
rect 3227 998 3367 1002
rect 3371 998 3463 1002
rect 3467 998 3499 1002
rect 1797 997 3499 998
rect 3505 997 3506 1003
rect 96 977 97 983
rect 103 982 1791 983
rect 103 978 111 982
rect 115 978 327 982
rect 331 978 463 982
rect 467 978 471 982
rect 475 978 567 982
rect 571 978 607 982
rect 611 978 671 982
rect 675 978 767 982
rect 771 978 783 982
rect 787 978 887 982
rect 891 978 927 982
rect 931 978 991 982
rect 995 978 1079 982
rect 1083 978 1095 982
rect 1099 978 1199 982
rect 1203 978 1231 982
rect 1235 978 1295 982
rect 1299 978 1383 982
rect 1387 978 1391 982
rect 1395 978 1487 982
rect 1491 978 1535 982
rect 1539 978 1583 982
rect 1587 978 1671 982
rect 1675 978 1767 982
rect 1771 978 1791 982
rect 103 977 1791 978
rect 1797 977 1798 983
rect 1778 921 1779 927
rect 1785 926 3487 927
rect 1785 922 1807 926
rect 1811 922 1831 926
rect 1835 922 1983 926
rect 1987 922 2151 926
rect 2155 922 2311 926
rect 2315 922 2327 926
rect 2331 922 2407 926
rect 2411 922 2511 926
rect 2515 922 2519 926
rect 2523 922 2623 926
rect 2627 922 2719 926
rect 2723 922 2751 926
rect 2755 922 2895 926
rect 2899 922 2935 926
rect 2939 922 3055 926
rect 3059 922 3159 926
rect 3163 922 3223 926
rect 3227 922 3367 926
rect 3371 922 3463 926
rect 3467 922 3487 926
rect 1785 921 3487 922
rect 3493 921 3494 927
rect 84 909 85 915
rect 91 914 1779 915
rect 91 910 111 914
rect 115 910 471 914
rect 475 910 567 914
rect 571 910 607 914
rect 611 910 671 914
rect 675 910 695 914
rect 699 910 783 914
rect 787 910 791 914
rect 795 910 887 914
rect 891 910 895 914
rect 899 910 991 914
rect 995 910 999 914
rect 1003 910 1095 914
rect 1099 910 1111 914
rect 1115 910 1199 914
rect 1203 910 1223 914
rect 1227 910 1295 914
rect 1299 910 1343 914
rect 1347 910 1391 914
rect 1395 910 1463 914
rect 1467 910 1487 914
rect 1491 910 1583 914
rect 1587 910 1671 914
rect 1675 910 1767 914
rect 1771 910 1779 914
rect 91 909 1779 910
rect 1785 909 1786 915
rect 1790 853 1791 859
rect 1797 858 3499 859
rect 1797 854 1807 858
rect 1811 854 1831 858
rect 1835 854 1959 858
rect 1963 854 1983 858
rect 1987 854 2087 858
rect 2091 854 2151 858
rect 2155 854 2207 858
rect 2211 854 2327 858
rect 2331 854 2463 858
rect 2467 854 2519 858
rect 2523 854 2615 858
rect 2619 854 2719 858
rect 2723 854 2791 858
rect 2795 854 2935 858
rect 2939 854 2983 858
rect 2987 854 3159 858
rect 3163 854 3183 858
rect 3187 854 3367 858
rect 3371 854 3463 858
rect 3467 854 3499 858
rect 1797 853 3499 854
rect 3505 853 3506 859
rect 96 841 97 847
rect 103 846 1791 847
rect 103 842 111 846
rect 115 842 519 846
rect 523 842 607 846
rect 611 842 615 846
rect 619 842 695 846
rect 699 842 719 846
rect 723 842 791 846
rect 795 842 831 846
rect 835 842 895 846
rect 899 842 951 846
rect 955 842 999 846
rect 1003 842 1071 846
rect 1075 842 1111 846
rect 1115 842 1191 846
rect 1195 842 1223 846
rect 1227 842 1311 846
rect 1315 842 1343 846
rect 1347 842 1431 846
rect 1435 842 1463 846
rect 1467 842 1559 846
rect 1563 842 1583 846
rect 1587 842 1767 846
rect 1771 842 1791 846
rect 103 841 1791 842
rect 1797 841 1798 847
rect 1778 785 1779 791
rect 1785 790 3487 791
rect 1785 786 1807 790
rect 1811 786 1831 790
rect 1835 786 1879 790
rect 1883 786 1959 790
rect 1963 786 2015 790
rect 2019 786 2087 790
rect 2091 786 2151 790
rect 2155 786 2207 790
rect 2211 786 2287 790
rect 2291 786 2327 790
rect 2331 786 2423 790
rect 2427 786 2463 790
rect 2467 786 2559 790
rect 2563 786 2615 790
rect 2619 786 2711 790
rect 2715 786 2791 790
rect 2795 786 2871 790
rect 2875 786 2983 790
rect 2987 786 3039 790
rect 3043 786 3183 790
rect 3187 786 3215 790
rect 3219 786 3367 790
rect 3371 786 3463 790
rect 3467 786 3487 790
rect 1785 785 3487 786
rect 3493 785 3494 791
rect 84 773 85 779
rect 91 778 1779 779
rect 91 774 111 778
rect 115 774 383 778
rect 387 774 471 778
rect 475 774 519 778
rect 523 774 575 778
rect 579 774 615 778
rect 619 774 679 778
rect 683 774 719 778
rect 723 774 791 778
rect 795 774 831 778
rect 835 774 911 778
rect 915 774 951 778
rect 955 774 1031 778
rect 1035 774 1071 778
rect 1075 774 1159 778
rect 1163 774 1191 778
rect 1195 774 1287 778
rect 1291 774 1311 778
rect 1315 774 1415 778
rect 1419 774 1431 778
rect 1435 774 1559 778
rect 1563 774 1767 778
rect 1771 774 1779 778
rect 91 773 1779 774
rect 1785 773 1786 779
rect 1790 717 1791 723
rect 1797 722 3499 723
rect 1797 718 1807 722
rect 1811 718 1831 722
rect 1835 718 1879 722
rect 1883 718 1951 722
rect 1955 718 2015 722
rect 2019 718 2103 722
rect 2107 718 2151 722
rect 2155 718 2263 722
rect 2267 718 2287 722
rect 2291 718 2415 722
rect 2419 718 2423 722
rect 2427 718 2559 722
rect 2563 718 2567 722
rect 2571 718 2711 722
rect 2715 718 2719 722
rect 2723 718 2871 722
rect 2875 718 2879 722
rect 2883 718 3039 722
rect 3043 718 3199 722
rect 3203 718 3215 722
rect 3219 718 3367 722
rect 3371 718 3463 722
rect 3467 718 3499 722
rect 1797 717 3499 718
rect 3505 717 3506 723
rect 96 701 97 707
rect 103 706 1791 707
rect 103 702 111 706
rect 115 702 247 706
rect 251 702 343 706
rect 347 702 383 706
rect 387 702 455 706
rect 459 702 471 706
rect 475 702 567 706
rect 571 702 575 706
rect 579 702 679 706
rect 683 702 695 706
rect 699 702 791 706
rect 795 702 831 706
rect 835 702 911 706
rect 915 702 983 706
rect 987 702 1031 706
rect 1035 702 1151 706
rect 1155 702 1159 706
rect 1163 702 1287 706
rect 1291 702 1327 706
rect 1331 702 1415 706
rect 1419 702 1511 706
rect 1515 702 1671 706
rect 1675 702 1767 706
rect 1771 702 1791 706
rect 103 701 1791 702
rect 1797 701 1798 707
rect 1778 653 1779 659
rect 1785 658 3487 659
rect 1785 654 1807 658
rect 1811 654 1831 658
rect 1835 654 1951 658
rect 1955 654 1975 658
rect 1979 654 2103 658
rect 2107 654 2239 658
rect 2243 654 2263 658
rect 2267 654 2415 658
rect 2419 654 2479 658
rect 2483 654 2567 658
rect 2571 654 2687 658
rect 2691 654 2719 658
rect 2723 654 2879 658
rect 2883 654 3039 658
rect 3043 654 3055 658
rect 3059 654 3199 658
rect 3203 654 3223 658
rect 3227 654 3367 658
rect 3371 654 3463 658
rect 3467 654 3487 658
rect 1785 653 3487 654
rect 3493 653 3494 659
rect 84 633 85 639
rect 91 638 1779 639
rect 91 634 111 638
rect 115 634 135 638
rect 139 634 231 638
rect 235 634 247 638
rect 251 634 343 638
rect 347 634 359 638
rect 363 634 455 638
rect 459 634 487 638
rect 491 634 567 638
rect 571 634 623 638
rect 627 634 695 638
rect 699 634 767 638
rect 771 634 831 638
rect 835 634 911 638
rect 915 634 983 638
rect 987 634 1055 638
rect 1059 634 1151 638
rect 1155 634 1207 638
rect 1211 634 1327 638
rect 1331 634 1367 638
rect 1371 634 1511 638
rect 1515 634 1527 638
rect 1531 634 1671 638
rect 1675 634 1767 638
rect 1771 634 1779 638
rect 91 633 1779 634
rect 1785 633 1786 639
rect 1790 581 1791 587
rect 1797 586 3499 587
rect 1797 582 1807 586
rect 1811 582 1895 586
rect 1899 582 1975 586
rect 1979 582 2015 586
rect 2019 582 2143 586
rect 2147 582 2239 586
rect 2243 582 2279 586
rect 2283 582 2423 586
rect 2427 582 2479 586
rect 2483 582 2567 586
rect 2571 582 2687 586
rect 2691 582 2719 586
rect 2723 582 2871 586
rect 2875 582 2879 586
rect 2883 582 3031 586
rect 3035 582 3055 586
rect 3059 582 3199 586
rect 3203 582 3223 586
rect 3227 582 3367 586
rect 3371 582 3463 586
rect 3467 582 3499 586
rect 1797 581 3499 582
rect 3505 581 3506 587
rect 96 565 97 571
rect 103 570 1791 571
rect 103 566 111 570
rect 115 566 135 570
rect 139 566 231 570
rect 235 566 247 570
rect 251 566 359 570
rect 363 566 407 570
rect 411 566 487 570
rect 491 566 583 570
rect 587 566 623 570
rect 627 566 767 570
rect 771 566 911 570
rect 915 566 951 570
rect 955 566 1055 570
rect 1059 566 1135 570
rect 1139 566 1207 570
rect 1211 566 1319 570
rect 1323 566 1367 570
rect 1371 566 1503 570
rect 1507 566 1527 570
rect 1531 566 1671 570
rect 1675 566 1767 570
rect 1771 566 1791 570
rect 103 565 1791 566
rect 1797 565 1798 571
rect 1778 513 1779 519
rect 1785 518 3487 519
rect 1785 514 1807 518
rect 1811 514 1895 518
rect 1899 514 2015 518
rect 2019 514 2135 518
rect 2139 514 2143 518
rect 2147 514 2239 518
rect 2243 514 2279 518
rect 2283 514 2359 518
rect 2363 514 2423 518
rect 2427 514 2487 518
rect 2491 514 2567 518
rect 2571 514 2615 518
rect 2619 514 2719 518
rect 2723 514 2751 518
rect 2755 514 2871 518
rect 2875 514 2879 518
rect 2883 514 3007 518
rect 3011 514 3031 518
rect 3035 514 3135 518
rect 3139 514 3199 518
rect 3203 514 3263 518
rect 3267 514 3367 518
rect 3371 514 3463 518
rect 3467 514 3487 518
rect 1785 513 3487 514
rect 3493 513 3494 519
rect 84 497 85 503
rect 91 502 1779 503
rect 91 498 111 502
rect 115 498 135 502
rect 139 498 247 502
rect 251 498 399 502
rect 403 498 407 502
rect 411 498 567 502
rect 571 498 583 502
rect 587 498 735 502
rect 739 498 767 502
rect 771 498 903 502
rect 907 498 951 502
rect 955 498 1063 502
rect 1067 498 1135 502
rect 1139 498 1223 502
rect 1227 498 1319 502
rect 1323 498 1375 502
rect 1379 498 1503 502
rect 1507 498 1527 502
rect 1531 498 1671 502
rect 1675 498 1767 502
rect 1771 498 1779 502
rect 91 497 1779 498
rect 1785 497 1786 503
rect 1790 441 1791 447
rect 1797 446 3499 447
rect 1797 442 1807 446
rect 1811 442 2135 446
rect 2139 442 2239 446
rect 2243 442 2335 446
rect 2339 442 2359 446
rect 2363 442 2447 446
rect 2451 442 2487 446
rect 2491 442 2559 446
rect 2563 442 2615 446
rect 2619 442 2679 446
rect 2683 442 2751 446
rect 2755 442 2799 446
rect 2803 442 2879 446
rect 2883 442 2911 446
rect 2915 442 3007 446
rect 3011 442 3023 446
rect 3027 442 3135 446
rect 3139 442 3143 446
rect 3147 442 3263 446
rect 3267 442 3367 446
rect 3371 442 3463 446
rect 3467 442 3499 446
rect 1797 441 3499 442
rect 3505 441 3506 447
rect 96 429 97 435
rect 103 434 1791 435
rect 103 430 111 434
rect 115 430 247 434
rect 251 430 399 434
rect 403 430 519 434
rect 523 430 567 434
rect 571 430 615 434
rect 619 430 719 434
rect 723 430 735 434
rect 739 430 823 434
rect 827 430 903 434
rect 907 430 927 434
rect 931 430 1023 434
rect 1027 430 1063 434
rect 1067 430 1127 434
rect 1131 430 1223 434
rect 1227 430 1231 434
rect 1235 430 1335 434
rect 1339 430 1375 434
rect 1379 430 1439 434
rect 1443 430 1527 434
rect 1531 430 1671 434
rect 1675 430 1767 434
rect 1771 430 1791 434
rect 103 429 1791 430
rect 1797 429 1798 435
rect 1778 373 1779 379
rect 1785 378 3487 379
rect 1785 374 1807 378
rect 1811 374 2063 378
rect 2067 374 2151 378
rect 2155 374 2239 378
rect 2243 374 2247 378
rect 2251 374 2335 378
rect 2339 374 2359 378
rect 2363 374 2447 378
rect 2451 374 2479 378
rect 2483 374 2559 378
rect 2563 374 2615 378
rect 2619 374 2679 378
rect 2683 374 2759 378
rect 2763 374 2799 378
rect 2803 374 2911 378
rect 2915 374 3023 378
rect 3027 374 3063 378
rect 3067 374 3143 378
rect 3147 374 3223 378
rect 3227 374 3263 378
rect 3267 374 3367 378
rect 3371 374 3463 378
rect 3467 374 3487 378
rect 1785 373 3487 374
rect 3493 373 3494 379
rect 84 361 85 367
rect 91 366 1779 367
rect 91 362 111 366
rect 115 362 471 366
rect 475 362 519 366
rect 523 362 559 366
rect 563 362 615 366
rect 619 362 647 366
rect 651 362 719 366
rect 723 362 735 366
rect 739 362 823 366
rect 827 362 911 366
rect 915 362 927 366
rect 931 362 999 366
rect 1003 362 1023 366
rect 1027 362 1087 366
rect 1091 362 1127 366
rect 1131 362 1175 366
rect 1179 362 1231 366
rect 1235 362 1263 366
rect 1267 362 1335 366
rect 1339 362 1439 366
rect 1443 362 1767 366
rect 1771 362 1779 366
rect 91 361 1779 362
rect 1785 361 1786 367
rect 1790 305 1791 311
rect 1797 310 3499 311
rect 1797 306 1807 310
rect 1811 306 1927 310
rect 1931 306 2039 310
rect 2043 306 2063 310
rect 2067 306 2151 310
rect 2155 306 2167 310
rect 2171 306 2247 310
rect 2251 306 2303 310
rect 2307 306 2359 310
rect 2363 306 2447 310
rect 2451 306 2479 310
rect 2483 306 2599 310
rect 2603 306 2615 310
rect 2619 306 2759 310
rect 2763 306 2911 310
rect 2915 306 2919 310
rect 2923 306 3063 310
rect 3067 306 3087 310
rect 3091 306 3223 310
rect 3227 306 3255 310
rect 3259 306 3367 310
rect 3371 306 3463 310
rect 3467 306 3499 310
rect 1797 305 3499 306
rect 3505 305 3506 311
rect 96 293 97 299
rect 103 298 1791 299
rect 103 294 111 298
rect 115 294 279 298
rect 283 294 367 298
rect 371 294 463 298
rect 467 294 471 298
rect 475 294 559 298
rect 563 294 647 298
rect 651 294 655 298
rect 659 294 735 298
rect 739 294 751 298
rect 755 294 823 298
rect 827 294 847 298
rect 851 294 911 298
rect 915 294 943 298
rect 947 294 999 298
rect 1003 294 1047 298
rect 1051 294 1087 298
rect 1091 294 1151 298
rect 1155 294 1175 298
rect 1179 294 1263 298
rect 1267 294 1767 298
rect 1771 294 1791 298
rect 103 293 1791 294
rect 1797 293 1798 299
rect 1778 237 1779 243
rect 1785 242 3487 243
rect 1785 238 1807 242
rect 1811 238 1831 242
rect 1835 238 1927 242
rect 1931 238 2039 242
rect 2043 238 2055 242
rect 2059 238 2167 242
rect 2171 238 2199 242
rect 2203 238 2303 242
rect 2307 238 2351 242
rect 2355 238 2447 242
rect 2451 238 2511 242
rect 2515 238 2599 242
rect 2603 238 2679 242
rect 2683 238 2759 242
rect 2763 238 2847 242
rect 2851 238 2919 242
rect 2923 238 3023 242
rect 3027 238 3087 242
rect 3091 238 3207 242
rect 3211 238 3255 242
rect 3259 238 3367 242
rect 3371 238 3463 242
rect 3467 238 3487 242
rect 1785 237 3487 238
rect 3493 237 3494 243
rect 84 225 85 231
rect 91 230 1779 231
rect 91 226 111 230
rect 115 226 167 230
rect 171 226 279 230
rect 283 226 343 230
rect 347 226 367 230
rect 371 226 463 230
rect 467 226 511 230
rect 515 226 559 230
rect 563 226 655 230
rect 659 226 679 230
rect 683 226 751 230
rect 755 226 839 230
rect 843 226 847 230
rect 851 226 943 230
rect 947 226 991 230
rect 995 226 1047 230
rect 1051 226 1135 230
rect 1139 226 1151 230
rect 1155 226 1279 230
rect 1283 226 1431 230
rect 1435 226 1767 230
rect 1771 226 1779 230
rect 91 225 1779 226
rect 1785 225 1786 231
rect 230 164 236 165
rect 742 164 748 165
rect 230 160 231 164
rect 235 160 743 164
rect 747 160 748 164
rect 230 159 236 160
rect 742 159 748 160
rect 1790 153 1791 159
rect 1797 158 3499 159
rect 1797 154 1807 158
rect 1811 154 1831 158
rect 1835 154 1919 158
rect 1923 154 1927 158
rect 1931 154 2039 158
rect 2043 154 2055 158
rect 2059 154 2159 158
rect 2163 154 2199 158
rect 2203 154 2279 158
rect 2283 154 2351 158
rect 2355 154 2399 158
rect 2403 154 2511 158
rect 2515 154 2623 158
rect 2627 154 2679 158
rect 2683 154 2735 158
rect 2739 154 2839 158
rect 2843 154 2847 158
rect 2851 154 2943 158
rect 2947 154 3023 158
rect 3027 154 3055 158
rect 3059 154 3167 158
rect 3171 154 3207 158
rect 3211 154 3279 158
rect 3283 154 3367 158
rect 3371 154 3463 158
rect 3467 154 3499 158
rect 1797 153 3499 154
rect 3505 153 3506 159
rect 96 137 97 143
rect 103 142 1791 143
rect 103 138 111 142
rect 115 138 135 142
rect 139 138 167 142
rect 171 138 223 142
rect 227 138 311 142
rect 315 138 343 142
rect 347 138 399 142
rect 403 138 487 142
rect 491 138 511 142
rect 515 138 575 142
rect 579 138 663 142
rect 667 138 679 142
rect 683 138 751 142
rect 755 138 839 142
rect 843 138 847 142
rect 851 138 943 142
rect 947 138 991 142
rect 995 138 1031 142
rect 1035 138 1119 142
rect 1123 138 1135 142
rect 1139 138 1215 142
rect 1219 138 1279 142
rect 1283 138 1311 142
rect 1315 138 1407 142
rect 1411 138 1431 142
rect 1435 138 1495 142
rect 1499 138 1583 142
rect 1587 138 1671 142
rect 1675 138 1767 142
rect 1771 138 1791 142
rect 103 137 1791 138
rect 1797 137 1798 143
rect 902 92 908 93
rect 1398 92 1404 93
rect 902 88 903 92
rect 907 88 1399 92
rect 1403 88 1404 92
rect 1778 89 1779 95
rect 1785 94 3487 95
rect 1785 90 1807 94
rect 1811 90 1831 94
rect 1835 90 1919 94
rect 1923 90 2039 94
rect 2043 90 2159 94
rect 2163 90 2279 94
rect 2283 90 2399 94
rect 2403 90 2511 94
rect 2515 90 2623 94
rect 2627 90 2735 94
rect 2739 90 2839 94
rect 2843 90 2943 94
rect 2947 90 3055 94
rect 3059 90 3167 94
rect 3171 90 3279 94
rect 3283 90 3367 94
rect 3371 90 3463 94
rect 3467 90 3487 94
rect 1785 89 3487 90
rect 3493 89 3494 95
rect 902 87 908 88
rect 1398 87 1404 88
rect 84 73 85 79
rect 91 78 1779 79
rect 91 74 111 78
rect 115 74 135 78
rect 139 74 223 78
rect 227 74 311 78
rect 315 74 399 78
rect 403 74 487 78
rect 491 74 575 78
rect 579 74 663 78
rect 667 74 751 78
rect 755 74 847 78
rect 851 74 943 78
rect 947 74 1031 78
rect 1035 74 1119 78
rect 1123 74 1215 78
rect 1219 74 1311 78
rect 1315 74 1407 78
rect 1411 74 1495 78
rect 1499 74 1583 78
rect 1587 74 1671 78
rect 1675 74 1767 78
rect 1771 74 1779 78
rect 91 73 1779 74
rect 1785 73 1786 79
<< m5c >>
rect 1791 3517 1797 3523
rect 3499 3517 3505 3523
rect 97 3481 103 3487
rect 1791 3481 1797 3487
rect 1779 3453 1785 3459
rect 3487 3453 3493 3459
rect 85 3417 91 3423
rect 1779 3417 1785 3423
rect 1791 3381 1797 3387
rect 3499 3381 3505 3387
rect 97 3349 103 3355
rect 1791 3349 1797 3355
rect 1779 3309 1785 3315
rect 3487 3309 3493 3315
rect 85 3281 91 3287
rect 1779 3281 1785 3287
rect 1791 3237 1797 3243
rect 3499 3237 3505 3243
rect 97 3213 103 3219
rect 1791 3213 1797 3219
rect 1779 3173 1785 3179
rect 3487 3173 3493 3179
rect 85 3137 91 3143
rect 1779 3137 1785 3143
rect 1791 3105 1797 3111
rect 3499 3105 3505 3111
rect 97 3065 103 3071
rect 1791 3065 1797 3071
rect 1779 3033 1785 3039
rect 3487 3033 3493 3039
rect 85 2997 91 3003
rect 1779 2997 1785 3003
rect 1791 2969 1797 2975
rect 3499 2969 3505 2975
rect 97 2925 103 2931
rect 1791 2925 1797 2931
rect 1779 2897 1785 2903
rect 3487 2897 3493 2903
rect 85 2857 91 2863
rect 1779 2857 1785 2863
rect 1791 2829 1797 2835
rect 3499 2829 3505 2835
rect 97 2785 103 2791
rect 1791 2785 1797 2791
rect 1779 2761 1785 2767
rect 3487 2761 3493 2767
rect 85 2717 91 2723
rect 1779 2717 1785 2723
rect 1791 2697 1797 2703
rect 3499 2697 3505 2703
rect 97 2645 103 2651
rect 1791 2645 1797 2651
rect 1779 2629 1785 2635
rect 3487 2629 3493 2635
rect 85 2569 91 2575
rect 1779 2569 1785 2575
rect 1791 2557 1797 2563
rect 3499 2557 3505 2563
rect 97 2505 103 2511
rect 1791 2505 1797 2511
rect 1779 2477 1785 2483
rect 3487 2477 3493 2483
rect 85 2425 91 2431
rect 1779 2425 1785 2431
rect 1791 2409 1797 2415
rect 3499 2409 3505 2415
rect 1779 2363 1785 2369
rect 97 2353 103 2359
rect 1791 2353 1797 2359
rect 3487 2345 3493 2351
rect 85 2281 91 2287
rect 1779 2281 1785 2287
rect 1791 2277 1797 2283
rect 3499 2277 3505 2283
rect 97 2217 103 2223
rect 1791 2217 1797 2223
rect 1779 2201 1785 2207
rect 3487 2201 3493 2207
rect 85 2137 91 2143
rect 1779 2137 1785 2143
rect 1791 2129 1797 2135
rect 3499 2129 3505 2135
rect 97 2073 103 2079
rect 1791 2073 1797 2079
rect 1779 2057 1785 2063
rect 3487 2057 3493 2063
rect 85 2009 91 2015
rect 1779 2009 1785 2015
rect 1791 1977 1797 1983
rect 3499 1977 3505 1983
rect 97 1945 103 1951
rect 1791 1945 1797 1951
rect 1779 1909 1785 1915
rect 3487 1909 3493 1915
rect 85 1881 91 1887
rect 1779 1881 1785 1887
rect 1791 1841 1797 1847
rect 3499 1841 3505 1847
rect 97 1809 103 1815
rect 1791 1809 1797 1815
rect 1779 1765 1785 1771
rect 3487 1765 3493 1771
rect 85 1733 91 1739
rect 1779 1733 1785 1739
rect 1791 1693 1797 1699
rect 3499 1693 3505 1699
rect 97 1665 103 1671
rect 1791 1665 1797 1671
rect 1779 1621 1785 1627
rect 3487 1621 3493 1627
rect 85 1597 91 1603
rect 1779 1597 1785 1603
rect 1791 1549 1797 1555
rect 3499 1549 3505 1555
rect 97 1529 103 1535
rect 1791 1529 1797 1535
rect 1779 1477 1785 1483
rect 3487 1477 3493 1483
rect 85 1457 91 1463
rect 1779 1457 1785 1463
rect 1791 1405 1797 1411
rect 3499 1405 3505 1411
rect 97 1389 103 1395
rect 1791 1389 1797 1395
rect 1779 1337 1785 1343
rect 3487 1337 3493 1343
rect 85 1321 91 1327
rect 1779 1321 1785 1327
rect 1791 1273 1797 1279
rect 3499 1273 3505 1279
rect 97 1253 103 1259
rect 1791 1253 1797 1259
rect 1779 1209 1785 1215
rect 3487 1209 3493 1215
rect 85 1185 91 1191
rect 1779 1185 1785 1191
rect 1791 1133 1797 1139
rect 3499 1133 3505 1139
rect 97 1117 103 1123
rect 1791 1117 1797 1123
rect 1779 1061 1785 1067
rect 3487 1061 3493 1067
rect 85 1045 91 1051
rect 1779 1045 1785 1051
rect 1791 997 1797 1003
rect 3499 997 3505 1003
rect 97 977 103 983
rect 1791 977 1797 983
rect 1779 921 1785 927
rect 3487 921 3493 927
rect 85 909 91 915
rect 1779 909 1785 915
rect 1791 853 1797 859
rect 3499 853 3505 859
rect 97 841 103 847
rect 1791 841 1797 847
rect 1779 785 1785 791
rect 3487 785 3493 791
rect 85 773 91 779
rect 1779 773 1785 779
rect 1791 717 1797 723
rect 3499 717 3505 723
rect 97 701 103 707
rect 1791 701 1797 707
rect 1779 653 1785 659
rect 3487 653 3493 659
rect 85 633 91 639
rect 1779 633 1785 639
rect 1791 581 1797 587
rect 3499 581 3505 587
rect 97 565 103 571
rect 1791 565 1797 571
rect 1779 513 1785 519
rect 3487 513 3493 519
rect 85 497 91 503
rect 1779 497 1785 503
rect 1791 441 1797 447
rect 3499 441 3505 447
rect 97 429 103 435
rect 1791 429 1797 435
rect 1779 373 1785 379
rect 3487 373 3493 379
rect 85 361 91 367
rect 1779 361 1785 367
rect 1791 305 1797 311
rect 3499 305 3505 311
rect 97 293 103 299
rect 1791 293 1797 299
rect 1779 237 1785 243
rect 3487 237 3493 243
rect 85 225 91 231
rect 1779 225 1785 231
rect 1791 153 1797 159
rect 3499 153 3505 159
rect 97 137 103 143
rect 1791 137 1797 143
rect 1779 89 1785 95
rect 3487 89 3493 95
rect 85 73 91 79
rect 1779 73 1785 79
<< m5 >>
rect 84 3423 92 3528
rect 84 3417 85 3423
rect 91 3417 92 3423
rect 84 3287 92 3417
rect 84 3281 85 3287
rect 91 3281 92 3287
rect 84 3143 92 3281
rect 84 3137 85 3143
rect 91 3137 92 3143
rect 84 3003 92 3137
rect 84 2997 85 3003
rect 91 2997 92 3003
rect 84 2863 92 2997
rect 84 2857 85 2863
rect 91 2857 92 2863
rect 84 2723 92 2857
rect 84 2717 85 2723
rect 91 2717 92 2723
rect 84 2575 92 2717
rect 84 2569 85 2575
rect 91 2569 92 2575
rect 84 2431 92 2569
rect 84 2425 85 2431
rect 91 2425 92 2431
rect 84 2287 92 2425
rect 84 2281 85 2287
rect 91 2281 92 2287
rect 84 2143 92 2281
rect 84 2137 85 2143
rect 91 2137 92 2143
rect 84 2015 92 2137
rect 84 2009 85 2015
rect 91 2009 92 2015
rect 84 1887 92 2009
rect 84 1881 85 1887
rect 91 1881 92 1887
rect 84 1739 92 1881
rect 84 1733 85 1739
rect 91 1733 92 1739
rect 84 1603 92 1733
rect 84 1597 85 1603
rect 91 1597 92 1603
rect 84 1463 92 1597
rect 84 1457 85 1463
rect 91 1457 92 1463
rect 84 1327 92 1457
rect 84 1321 85 1327
rect 91 1321 92 1327
rect 84 1191 92 1321
rect 84 1185 85 1191
rect 91 1185 92 1191
rect 84 1051 92 1185
rect 84 1045 85 1051
rect 91 1045 92 1051
rect 84 915 92 1045
rect 84 909 85 915
rect 91 909 92 915
rect 84 779 92 909
rect 84 773 85 779
rect 91 773 92 779
rect 84 639 92 773
rect 84 633 85 639
rect 91 633 92 639
rect 84 503 92 633
rect 84 497 85 503
rect 91 497 92 503
rect 84 367 92 497
rect 84 361 85 367
rect 91 361 92 367
rect 84 231 92 361
rect 84 225 85 231
rect 91 225 92 231
rect 84 79 92 225
rect 84 73 85 79
rect 91 73 92 79
rect 84 72 92 73
rect 96 3487 104 3528
rect 96 3481 97 3487
rect 103 3481 104 3487
rect 96 3355 104 3481
rect 96 3349 97 3355
rect 103 3349 104 3355
rect 96 3219 104 3349
rect 96 3213 97 3219
rect 103 3213 104 3219
rect 96 3071 104 3213
rect 96 3065 97 3071
rect 103 3065 104 3071
rect 96 2931 104 3065
rect 96 2925 97 2931
rect 103 2925 104 2931
rect 96 2791 104 2925
rect 96 2785 97 2791
rect 103 2785 104 2791
rect 96 2651 104 2785
rect 96 2645 97 2651
rect 103 2645 104 2651
rect 96 2511 104 2645
rect 96 2505 97 2511
rect 103 2505 104 2511
rect 96 2359 104 2505
rect 96 2353 97 2359
rect 103 2353 104 2359
rect 96 2223 104 2353
rect 96 2217 97 2223
rect 103 2217 104 2223
rect 96 2079 104 2217
rect 96 2073 97 2079
rect 103 2073 104 2079
rect 96 1951 104 2073
rect 96 1945 97 1951
rect 103 1945 104 1951
rect 96 1815 104 1945
rect 96 1809 97 1815
rect 103 1809 104 1815
rect 96 1671 104 1809
rect 96 1665 97 1671
rect 103 1665 104 1671
rect 96 1535 104 1665
rect 96 1529 97 1535
rect 103 1529 104 1535
rect 96 1395 104 1529
rect 96 1389 97 1395
rect 103 1389 104 1395
rect 96 1259 104 1389
rect 96 1253 97 1259
rect 103 1253 104 1259
rect 96 1123 104 1253
rect 96 1117 97 1123
rect 103 1117 104 1123
rect 96 983 104 1117
rect 96 977 97 983
rect 103 977 104 983
rect 96 847 104 977
rect 96 841 97 847
rect 103 841 104 847
rect 96 707 104 841
rect 96 701 97 707
rect 103 701 104 707
rect 96 571 104 701
rect 96 565 97 571
rect 103 565 104 571
rect 96 435 104 565
rect 96 429 97 435
rect 103 429 104 435
rect 96 299 104 429
rect 96 293 97 299
rect 103 293 104 299
rect 96 143 104 293
rect 96 137 97 143
rect 103 137 104 143
rect 96 72 104 137
rect 1778 3459 1786 3528
rect 1778 3453 1779 3459
rect 1785 3453 1786 3459
rect 1778 3423 1786 3453
rect 1778 3417 1779 3423
rect 1785 3417 1786 3423
rect 1778 3315 1786 3417
rect 1778 3309 1779 3315
rect 1785 3309 1786 3315
rect 1778 3287 1786 3309
rect 1778 3281 1779 3287
rect 1785 3281 1786 3287
rect 1778 3179 1786 3281
rect 1778 3173 1779 3179
rect 1785 3173 1786 3179
rect 1778 3143 1786 3173
rect 1778 3137 1779 3143
rect 1785 3137 1786 3143
rect 1778 3039 1786 3137
rect 1778 3033 1779 3039
rect 1785 3033 1786 3039
rect 1778 3003 1786 3033
rect 1778 2997 1779 3003
rect 1785 2997 1786 3003
rect 1778 2903 1786 2997
rect 1778 2897 1779 2903
rect 1785 2897 1786 2903
rect 1778 2863 1786 2897
rect 1778 2857 1779 2863
rect 1785 2857 1786 2863
rect 1778 2767 1786 2857
rect 1778 2761 1779 2767
rect 1785 2761 1786 2767
rect 1778 2723 1786 2761
rect 1778 2717 1779 2723
rect 1785 2717 1786 2723
rect 1778 2635 1786 2717
rect 1778 2629 1779 2635
rect 1785 2629 1786 2635
rect 1778 2575 1786 2629
rect 1778 2569 1779 2575
rect 1785 2569 1786 2575
rect 1778 2483 1786 2569
rect 1778 2477 1779 2483
rect 1785 2477 1786 2483
rect 1778 2431 1786 2477
rect 1778 2425 1779 2431
rect 1785 2425 1786 2431
rect 1778 2369 1786 2425
rect 1778 2363 1779 2369
rect 1785 2363 1786 2369
rect 1778 2287 1786 2363
rect 1778 2281 1779 2287
rect 1785 2281 1786 2287
rect 1778 2207 1786 2281
rect 1778 2201 1779 2207
rect 1785 2201 1786 2207
rect 1778 2143 1786 2201
rect 1778 2137 1779 2143
rect 1785 2137 1786 2143
rect 1778 2063 1786 2137
rect 1778 2057 1779 2063
rect 1785 2057 1786 2063
rect 1778 2015 1786 2057
rect 1778 2009 1779 2015
rect 1785 2009 1786 2015
rect 1778 1915 1786 2009
rect 1778 1909 1779 1915
rect 1785 1909 1786 1915
rect 1778 1887 1786 1909
rect 1778 1881 1779 1887
rect 1785 1881 1786 1887
rect 1778 1771 1786 1881
rect 1778 1765 1779 1771
rect 1785 1765 1786 1771
rect 1778 1739 1786 1765
rect 1778 1733 1779 1739
rect 1785 1733 1786 1739
rect 1778 1627 1786 1733
rect 1778 1621 1779 1627
rect 1785 1621 1786 1627
rect 1778 1603 1786 1621
rect 1778 1597 1779 1603
rect 1785 1597 1786 1603
rect 1778 1483 1786 1597
rect 1778 1477 1779 1483
rect 1785 1477 1786 1483
rect 1778 1463 1786 1477
rect 1778 1457 1779 1463
rect 1785 1457 1786 1463
rect 1778 1343 1786 1457
rect 1778 1337 1779 1343
rect 1785 1337 1786 1343
rect 1778 1327 1786 1337
rect 1778 1321 1779 1327
rect 1785 1321 1786 1327
rect 1778 1215 1786 1321
rect 1778 1209 1779 1215
rect 1785 1209 1786 1215
rect 1778 1191 1786 1209
rect 1778 1185 1779 1191
rect 1785 1185 1786 1191
rect 1778 1067 1786 1185
rect 1778 1061 1779 1067
rect 1785 1061 1786 1067
rect 1778 1051 1786 1061
rect 1778 1045 1779 1051
rect 1785 1045 1786 1051
rect 1778 927 1786 1045
rect 1778 921 1779 927
rect 1785 921 1786 927
rect 1778 915 1786 921
rect 1778 909 1779 915
rect 1785 909 1786 915
rect 1778 791 1786 909
rect 1778 785 1779 791
rect 1785 785 1786 791
rect 1778 779 1786 785
rect 1778 773 1779 779
rect 1785 773 1786 779
rect 1778 659 1786 773
rect 1778 653 1779 659
rect 1785 653 1786 659
rect 1778 639 1786 653
rect 1778 633 1779 639
rect 1785 633 1786 639
rect 1778 519 1786 633
rect 1778 513 1779 519
rect 1785 513 1786 519
rect 1778 503 1786 513
rect 1778 497 1779 503
rect 1785 497 1786 503
rect 1778 379 1786 497
rect 1778 373 1779 379
rect 1785 373 1786 379
rect 1778 367 1786 373
rect 1778 361 1779 367
rect 1785 361 1786 367
rect 1778 243 1786 361
rect 1778 237 1779 243
rect 1785 237 1786 243
rect 1778 231 1786 237
rect 1778 225 1779 231
rect 1785 225 1786 231
rect 1778 95 1786 225
rect 1778 89 1779 95
rect 1785 89 1786 95
rect 1778 79 1786 89
rect 1778 73 1779 79
rect 1785 73 1786 79
rect 1778 72 1786 73
rect 1790 3523 1798 3528
rect 1790 3517 1791 3523
rect 1797 3517 1798 3523
rect 1790 3487 1798 3517
rect 1790 3481 1791 3487
rect 1797 3481 1798 3487
rect 1790 3387 1798 3481
rect 1790 3381 1791 3387
rect 1797 3381 1798 3387
rect 1790 3355 1798 3381
rect 1790 3349 1791 3355
rect 1797 3349 1798 3355
rect 1790 3243 1798 3349
rect 1790 3237 1791 3243
rect 1797 3237 1798 3243
rect 1790 3219 1798 3237
rect 1790 3213 1791 3219
rect 1797 3213 1798 3219
rect 1790 3111 1798 3213
rect 1790 3105 1791 3111
rect 1797 3105 1798 3111
rect 1790 3071 1798 3105
rect 1790 3065 1791 3071
rect 1797 3065 1798 3071
rect 1790 2975 1798 3065
rect 1790 2969 1791 2975
rect 1797 2969 1798 2975
rect 1790 2931 1798 2969
rect 1790 2925 1791 2931
rect 1797 2925 1798 2931
rect 1790 2835 1798 2925
rect 1790 2829 1791 2835
rect 1797 2829 1798 2835
rect 1790 2791 1798 2829
rect 1790 2785 1791 2791
rect 1797 2785 1798 2791
rect 1790 2703 1798 2785
rect 1790 2697 1791 2703
rect 1797 2697 1798 2703
rect 1790 2651 1798 2697
rect 1790 2645 1791 2651
rect 1797 2645 1798 2651
rect 1790 2563 1798 2645
rect 1790 2557 1791 2563
rect 1797 2557 1798 2563
rect 1790 2511 1798 2557
rect 1790 2505 1791 2511
rect 1797 2505 1798 2511
rect 1790 2415 1798 2505
rect 1790 2409 1791 2415
rect 1797 2409 1798 2415
rect 1790 2359 1798 2409
rect 1790 2353 1791 2359
rect 1797 2353 1798 2359
rect 1790 2283 1798 2353
rect 1790 2277 1791 2283
rect 1797 2277 1798 2283
rect 1790 2223 1798 2277
rect 1790 2217 1791 2223
rect 1797 2217 1798 2223
rect 1790 2135 1798 2217
rect 1790 2129 1791 2135
rect 1797 2129 1798 2135
rect 1790 2079 1798 2129
rect 1790 2073 1791 2079
rect 1797 2073 1798 2079
rect 1790 1983 1798 2073
rect 1790 1977 1791 1983
rect 1797 1977 1798 1983
rect 1790 1951 1798 1977
rect 1790 1945 1791 1951
rect 1797 1945 1798 1951
rect 1790 1847 1798 1945
rect 1790 1841 1791 1847
rect 1797 1841 1798 1847
rect 1790 1815 1798 1841
rect 1790 1809 1791 1815
rect 1797 1809 1798 1815
rect 1790 1699 1798 1809
rect 1790 1693 1791 1699
rect 1797 1693 1798 1699
rect 1790 1671 1798 1693
rect 1790 1665 1791 1671
rect 1797 1665 1798 1671
rect 1790 1555 1798 1665
rect 1790 1549 1791 1555
rect 1797 1549 1798 1555
rect 1790 1535 1798 1549
rect 1790 1529 1791 1535
rect 1797 1529 1798 1535
rect 1790 1411 1798 1529
rect 1790 1405 1791 1411
rect 1797 1405 1798 1411
rect 1790 1395 1798 1405
rect 1790 1389 1791 1395
rect 1797 1389 1798 1395
rect 1790 1279 1798 1389
rect 1790 1273 1791 1279
rect 1797 1273 1798 1279
rect 1790 1259 1798 1273
rect 1790 1253 1791 1259
rect 1797 1253 1798 1259
rect 1790 1139 1798 1253
rect 1790 1133 1791 1139
rect 1797 1133 1798 1139
rect 1790 1123 1798 1133
rect 1790 1117 1791 1123
rect 1797 1117 1798 1123
rect 1790 1003 1798 1117
rect 1790 997 1791 1003
rect 1797 997 1798 1003
rect 1790 983 1798 997
rect 1790 977 1791 983
rect 1797 977 1798 983
rect 1790 859 1798 977
rect 1790 853 1791 859
rect 1797 853 1798 859
rect 1790 847 1798 853
rect 1790 841 1791 847
rect 1797 841 1798 847
rect 1790 723 1798 841
rect 1790 717 1791 723
rect 1797 717 1798 723
rect 1790 707 1798 717
rect 1790 701 1791 707
rect 1797 701 1798 707
rect 1790 587 1798 701
rect 1790 581 1791 587
rect 1797 581 1798 587
rect 1790 571 1798 581
rect 1790 565 1791 571
rect 1797 565 1798 571
rect 1790 447 1798 565
rect 1790 441 1791 447
rect 1797 441 1798 447
rect 1790 435 1798 441
rect 1790 429 1791 435
rect 1797 429 1798 435
rect 1790 311 1798 429
rect 1790 305 1791 311
rect 1797 305 1798 311
rect 1790 299 1798 305
rect 1790 293 1791 299
rect 1797 293 1798 299
rect 1790 159 1798 293
rect 1790 153 1791 159
rect 1797 153 1798 159
rect 1790 143 1798 153
rect 1790 137 1791 143
rect 1797 137 1798 143
rect 1790 72 1798 137
rect 3486 3459 3494 3528
rect 3486 3453 3487 3459
rect 3493 3453 3494 3459
rect 3486 3315 3494 3453
rect 3486 3309 3487 3315
rect 3493 3309 3494 3315
rect 3486 3179 3494 3309
rect 3486 3173 3487 3179
rect 3493 3173 3494 3179
rect 3486 3039 3494 3173
rect 3486 3033 3487 3039
rect 3493 3033 3494 3039
rect 3486 2903 3494 3033
rect 3486 2897 3487 2903
rect 3493 2897 3494 2903
rect 3486 2767 3494 2897
rect 3486 2761 3487 2767
rect 3493 2761 3494 2767
rect 3486 2635 3494 2761
rect 3486 2629 3487 2635
rect 3493 2629 3494 2635
rect 3486 2483 3494 2629
rect 3486 2477 3487 2483
rect 3493 2477 3494 2483
rect 3486 2351 3494 2477
rect 3486 2345 3487 2351
rect 3493 2345 3494 2351
rect 3486 2207 3494 2345
rect 3486 2201 3487 2207
rect 3493 2201 3494 2207
rect 3486 2063 3494 2201
rect 3486 2057 3487 2063
rect 3493 2057 3494 2063
rect 3486 1915 3494 2057
rect 3486 1909 3487 1915
rect 3493 1909 3494 1915
rect 3486 1771 3494 1909
rect 3486 1765 3487 1771
rect 3493 1765 3494 1771
rect 3486 1627 3494 1765
rect 3486 1621 3487 1627
rect 3493 1621 3494 1627
rect 3486 1483 3494 1621
rect 3486 1477 3487 1483
rect 3493 1477 3494 1483
rect 3486 1343 3494 1477
rect 3486 1337 3487 1343
rect 3493 1337 3494 1343
rect 3486 1215 3494 1337
rect 3486 1209 3487 1215
rect 3493 1209 3494 1215
rect 3486 1067 3494 1209
rect 3486 1061 3487 1067
rect 3493 1061 3494 1067
rect 3486 927 3494 1061
rect 3486 921 3487 927
rect 3493 921 3494 927
rect 3486 791 3494 921
rect 3486 785 3487 791
rect 3493 785 3494 791
rect 3486 659 3494 785
rect 3486 653 3487 659
rect 3493 653 3494 659
rect 3486 519 3494 653
rect 3486 513 3487 519
rect 3493 513 3494 519
rect 3486 379 3494 513
rect 3486 373 3487 379
rect 3493 373 3494 379
rect 3486 243 3494 373
rect 3486 237 3487 243
rect 3493 237 3494 243
rect 3486 95 3494 237
rect 3486 89 3487 95
rect 3493 89 3494 95
rect 3486 72 3494 89
rect 3498 3523 3506 3528
rect 3498 3517 3499 3523
rect 3505 3517 3506 3523
rect 3498 3387 3506 3517
rect 3498 3381 3499 3387
rect 3505 3381 3506 3387
rect 3498 3243 3506 3381
rect 3498 3237 3499 3243
rect 3505 3237 3506 3243
rect 3498 3111 3506 3237
rect 3498 3105 3499 3111
rect 3505 3105 3506 3111
rect 3498 2975 3506 3105
rect 3498 2969 3499 2975
rect 3505 2969 3506 2975
rect 3498 2835 3506 2969
rect 3498 2829 3499 2835
rect 3505 2829 3506 2835
rect 3498 2703 3506 2829
rect 3498 2697 3499 2703
rect 3505 2697 3506 2703
rect 3498 2563 3506 2697
rect 3498 2557 3499 2563
rect 3505 2557 3506 2563
rect 3498 2415 3506 2557
rect 3498 2409 3499 2415
rect 3505 2409 3506 2415
rect 3498 2283 3506 2409
rect 3498 2277 3499 2283
rect 3505 2277 3506 2283
rect 3498 2135 3506 2277
rect 3498 2129 3499 2135
rect 3505 2129 3506 2135
rect 3498 1983 3506 2129
rect 3498 1977 3499 1983
rect 3505 1977 3506 1983
rect 3498 1847 3506 1977
rect 3498 1841 3499 1847
rect 3505 1841 3506 1847
rect 3498 1699 3506 1841
rect 3498 1693 3499 1699
rect 3505 1693 3506 1699
rect 3498 1555 3506 1693
rect 3498 1549 3499 1555
rect 3505 1549 3506 1555
rect 3498 1411 3506 1549
rect 3498 1405 3499 1411
rect 3505 1405 3506 1411
rect 3498 1279 3506 1405
rect 3498 1273 3499 1279
rect 3505 1273 3506 1279
rect 3498 1139 3506 1273
rect 3498 1133 3499 1139
rect 3505 1133 3506 1139
rect 3498 1003 3506 1133
rect 3498 997 3499 1003
rect 3505 997 3506 1003
rect 3498 859 3506 997
rect 3498 853 3499 859
rect 3505 853 3506 859
rect 3498 723 3506 853
rect 3498 717 3499 723
rect 3505 717 3506 723
rect 3498 587 3506 717
rect 3498 581 3499 587
rect 3505 581 3506 587
rect 3498 447 3506 581
rect 3498 441 3499 447
rect 3505 441 3506 447
rect 3498 311 3506 441
rect 3498 305 3499 311
rect 3505 305 3506 311
rect 3498 159 3506 305
rect 3498 153 3499 159
rect 3505 153 3506 159
rect 3498 72 3506 153
use circuitwell  npwells
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use circuitppnp  ppnps
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use welltap_svt  __well_tap__195
timestamp 1731220329
transform 1 0 3456 0 1 3476
box 7 3 12 24
use welltap_svt  __well_tap__194
timestamp 1731220329
transform 1 0 1800 0 1 3476
box 7 3 12 24
use welltap_svt  __well_tap__193
timestamp 1731220329
transform 1 0 3456 0 -1 3436
box 7 3 12 24
use welltap_svt  __well_tap__192
timestamp 1731220329
transform 1 0 1800 0 -1 3436
box 7 3 12 24
use welltap_svt  __well_tap__191
timestamp 1731220329
transform 1 0 3456 0 1 3340
box 7 3 12 24
use welltap_svt  __well_tap__190
timestamp 1731220329
transform 1 0 1800 0 1 3340
box 7 3 12 24
use welltap_svt  __well_tap__189
timestamp 1731220329
transform 1 0 3456 0 -1 3292
box 7 3 12 24
use welltap_svt  __well_tap__188
timestamp 1731220329
transform 1 0 1800 0 -1 3292
box 7 3 12 24
use welltap_svt  __well_tap__187
timestamp 1731220329
transform 1 0 3456 0 1 3196
box 7 3 12 24
use welltap_svt  __well_tap__186
timestamp 1731220329
transform 1 0 1800 0 1 3196
box 7 3 12 24
use welltap_svt  __well_tap__185
timestamp 1731220329
transform 1 0 3456 0 -1 3156
box 7 3 12 24
use welltap_svt  __well_tap__184
timestamp 1731220329
transform 1 0 1800 0 -1 3156
box 7 3 12 24
use welltap_svt  __well_tap__183
timestamp 1731220329
transform 1 0 3456 0 1 3064
box 7 3 12 24
use welltap_svt  __well_tap__182
timestamp 1731220329
transform 1 0 1800 0 1 3064
box 7 3 12 24
use welltap_svt  __well_tap__181
timestamp 1731220329
transform 1 0 3456 0 -1 3016
box 7 3 12 24
use welltap_svt  __well_tap__180
timestamp 1731220329
transform 1 0 1800 0 -1 3016
box 7 3 12 24
use welltap_svt  __well_tap__179
timestamp 1731220329
transform 1 0 3456 0 1 2928
box 7 3 12 24
use welltap_svt  __well_tap__178
timestamp 1731220329
transform 1 0 1800 0 1 2928
box 7 3 12 24
use welltap_svt  __well_tap__177
timestamp 1731220329
transform 1 0 3456 0 -1 2880
box 7 3 12 24
use welltap_svt  __well_tap__176
timestamp 1731220329
transform 1 0 1800 0 -1 2880
box 7 3 12 24
use welltap_svt  __well_tap__175
timestamp 1731220329
transform 1 0 3456 0 1 2788
box 7 3 12 24
use welltap_svt  __well_tap__174
timestamp 1731220329
transform 1 0 1800 0 1 2788
box 7 3 12 24
use welltap_svt  __well_tap__173
timestamp 1731220329
transform 1 0 3456 0 -1 2744
box 7 3 12 24
use welltap_svt  __well_tap__172
timestamp 1731220329
transform 1 0 1800 0 -1 2744
box 7 3 12 24
use welltap_svt  __well_tap__171
timestamp 1731220329
transform 1 0 3456 0 1 2656
box 7 3 12 24
use welltap_svt  __well_tap__170
timestamp 1731220329
transform 1 0 1800 0 1 2656
box 7 3 12 24
use welltap_svt  __well_tap__169
timestamp 1731220329
transform 1 0 3456 0 -1 2612
box 7 3 12 24
use welltap_svt  __well_tap__168
timestamp 1731220329
transform 1 0 1800 0 -1 2612
box 7 3 12 24
use welltap_svt  __well_tap__167
timestamp 1731220329
transform 1 0 3456 0 1 2516
box 7 3 12 24
use welltap_svt  __well_tap__166
timestamp 1731220329
transform 1 0 1800 0 1 2516
box 7 3 12 24
use welltap_svt  __well_tap__165
timestamp 1731220329
transform 1 0 3456 0 -1 2460
box 7 3 12 24
use welltap_svt  __well_tap__164
timestamp 1731220329
transform 1 0 1800 0 -1 2460
box 7 3 12 24
use welltap_svt  __well_tap__163
timestamp 1731220329
transform 1 0 3456 0 1 2368
box 7 3 12 24
use welltap_svt  __well_tap__162
timestamp 1731220329
transform 1 0 1800 0 1 2368
box 7 3 12 24
use welltap_svt  __well_tap__161
timestamp 1731220329
transform 1 0 3456 0 -1 2328
box 7 3 12 24
use welltap_svt  __well_tap__160
timestamp 1731220329
transform 1 0 1800 0 -1 2328
box 7 3 12 24
use welltap_svt  __well_tap__159
timestamp 1731220329
transform 1 0 3456 0 1 2236
box 7 3 12 24
use welltap_svt  __well_tap__158
timestamp 1731220329
transform 1 0 1800 0 1 2236
box 7 3 12 24
use welltap_svt  __well_tap__157
timestamp 1731220329
transform 1 0 3456 0 -1 2184
box 7 3 12 24
use welltap_svt  __well_tap__156
timestamp 1731220329
transform 1 0 1800 0 -1 2184
box 7 3 12 24
use welltap_svt  __well_tap__155
timestamp 1731220329
transform 1 0 3456 0 1 2088
box 7 3 12 24
use welltap_svt  __well_tap__154
timestamp 1731220329
transform 1 0 1800 0 1 2088
box 7 3 12 24
use welltap_svt  __well_tap__153
timestamp 1731220329
transform 1 0 3456 0 -1 2040
box 7 3 12 24
use welltap_svt  __well_tap__152
timestamp 1731220329
transform 1 0 1800 0 -1 2040
box 7 3 12 24
use welltap_svt  __well_tap__151
timestamp 1731220329
transform 1 0 3456 0 1 1936
box 7 3 12 24
use welltap_svt  __well_tap__150
timestamp 1731220329
transform 1 0 1800 0 1 1936
box 7 3 12 24
use welltap_svt  __well_tap__149
timestamp 1731220329
transform 1 0 3456 0 -1 1892
box 7 3 12 24
use welltap_svt  __well_tap__148
timestamp 1731220329
transform 1 0 1800 0 -1 1892
box 7 3 12 24
use welltap_svt  __well_tap__147
timestamp 1731220329
transform 1 0 3456 0 1 1800
box 7 3 12 24
use welltap_svt  __well_tap__146
timestamp 1731220329
transform 1 0 1800 0 1 1800
box 7 3 12 24
use welltap_svt  __well_tap__145
timestamp 1731220329
transform 1 0 3456 0 -1 1748
box 7 3 12 24
use welltap_svt  __well_tap__144
timestamp 1731220329
transform 1 0 1800 0 -1 1748
box 7 3 12 24
use welltap_svt  __well_tap__143
timestamp 1731220329
transform 1 0 3456 0 1 1652
box 7 3 12 24
use welltap_svt  __well_tap__142
timestamp 1731220329
transform 1 0 1800 0 1 1652
box 7 3 12 24
use welltap_svt  __well_tap__141
timestamp 1731220329
transform 1 0 3456 0 -1 1604
box 7 3 12 24
use welltap_svt  __well_tap__140
timestamp 1731220329
transform 1 0 1800 0 -1 1604
box 7 3 12 24
use welltap_svt  __well_tap__139
timestamp 1731220329
transform 1 0 3456 0 1 1508
box 7 3 12 24
use welltap_svt  __well_tap__138
timestamp 1731220329
transform 1 0 1800 0 1 1508
box 7 3 12 24
use welltap_svt  __well_tap__137
timestamp 1731220329
transform 1 0 3456 0 -1 1460
box 7 3 12 24
use welltap_svt  __well_tap__136
timestamp 1731220329
transform 1 0 1800 0 -1 1460
box 7 3 12 24
use welltap_svt  __well_tap__135
timestamp 1731220329
transform 1 0 3456 0 1 1364
box 7 3 12 24
use welltap_svt  __well_tap__134
timestamp 1731220329
transform 1 0 1800 0 1 1364
box 7 3 12 24
use welltap_svt  __well_tap__133
timestamp 1731220329
transform 1 0 3456 0 -1 1320
box 7 3 12 24
use welltap_svt  __well_tap__132
timestamp 1731220329
transform 1 0 1800 0 -1 1320
box 7 3 12 24
use welltap_svt  __well_tap__131
timestamp 1731220329
transform 1 0 3456 0 1 1232
box 7 3 12 24
use welltap_svt  __well_tap__130
timestamp 1731220329
transform 1 0 1800 0 1 1232
box 7 3 12 24
use welltap_svt  __well_tap__129
timestamp 1731220329
transform 1 0 3456 0 -1 1192
box 7 3 12 24
use welltap_svt  __well_tap__128
timestamp 1731220329
transform 1 0 1800 0 -1 1192
box 7 3 12 24
use welltap_svt  __well_tap__127
timestamp 1731220329
transform 1 0 3456 0 1 1092
box 7 3 12 24
use welltap_svt  __well_tap__126
timestamp 1731220329
transform 1 0 1800 0 1 1092
box 7 3 12 24
use welltap_svt  __well_tap__125
timestamp 1731220329
transform 1 0 3456 0 -1 1044
box 7 3 12 24
use welltap_svt  __well_tap__124
timestamp 1731220329
transform 1 0 1800 0 -1 1044
box 7 3 12 24
use welltap_svt  __well_tap__123
timestamp 1731220329
transform 1 0 3456 0 1 956
box 7 3 12 24
use welltap_svt  __well_tap__122
timestamp 1731220329
transform 1 0 1800 0 1 956
box 7 3 12 24
use welltap_svt  __well_tap__121
timestamp 1731220329
transform 1 0 3456 0 -1 904
box 7 3 12 24
use welltap_svt  __well_tap__120
timestamp 1731220329
transform 1 0 1800 0 -1 904
box 7 3 12 24
use welltap_svt  __well_tap__119
timestamp 1731220329
transform 1 0 3456 0 1 812
box 7 3 12 24
use welltap_svt  __well_tap__118
timestamp 1731220329
transform 1 0 1800 0 1 812
box 7 3 12 24
use welltap_svt  __well_tap__117
timestamp 1731220329
transform 1 0 3456 0 -1 768
box 7 3 12 24
use welltap_svt  __well_tap__116
timestamp 1731220329
transform 1 0 1800 0 -1 768
box 7 3 12 24
use welltap_svt  __well_tap__115
timestamp 1731220329
transform 1 0 3456 0 1 676
box 7 3 12 24
use welltap_svt  __well_tap__114
timestamp 1731220329
transform 1 0 1800 0 1 676
box 7 3 12 24
use welltap_svt  __well_tap__113
timestamp 1731220329
transform 1 0 3456 0 -1 636
box 7 3 12 24
use welltap_svt  __well_tap__112
timestamp 1731220329
transform 1 0 1800 0 -1 636
box 7 3 12 24
use welltap_svt  __well_tap__111
timestamp 1731220329
transform 1 0 3456 0 1 540
box 7 3 12 24
use welltap_svt  __well_tap__110
timestamp 1731220329
transform 1 0 1800 0 1 540
box 7 3 12 24
use welltap_svt  __well_tap__109
timestamp 1731220329
transform 1 0 3456 0 -1 496
box 7 3 12 24
use welltap_svt  __well_tap__108
timestamp 1731220329
transform 1 0 1800 0 -1 496
box 7 3 12 24
use welltap_svt  __well_tap__107
timestamp 1731220329
transform 1 0 3456 0 1 400
box 7 3 12 24
use welltap_svt  __well_tap__106
timestamp 1731220329
transform 1 0 1800 0 1 400
box 7 3 12 24
use welltap_svt  __well_tap__105
timestamp 1731220329
transform 1 0 3456 0 -1 356
box 7 3 12 24
use welltap_svt  __well_tap__104
timestamp 1731220329
transform 1 0 1800 0 -1 356
box 7 3 12 24
use welltap_svt  __well_tap__103
timestamp 1731220329
transform 1 0 3456 0 1 264
box 7 3 12 24
use welltap_svt  __well_tap__102
timestamp 1731220329
transform 1 0 1800 0 1 264
box 7 3 12 24
use welltap_svt  __well_tap__101
timestamp 1731220329
transform 1 0 3456 0 -1 220
box 7 3 12 24
use welltap_svt  __well_tap__100
timestamp 1731220329
transform 1 0 1800 0 -1 220
box 7 3 12 24
use welltap_svt  __well_tap__99
timestamp 1731220329
transform 1 0 3456 0 1 112
box 7 3 12 24
use welltap_svt  __well_tap__98
timestamp 1731220329
transform 1 0 1800 0 1 112
box 7 3 12 24
use welltap_svt  __well_tap__97
timestamp 1731220329
transform 1 0 1760 0 1 3440
box 7 3 12 24
use welltap_svt  __well_tap__96
timestamp 1731220329
transform 1 0 104 0 1 3440
box 7 3 12 24
use welltap_svt  __well_tap__95
timestamp 1731220329
transform 1 0 1760 0 -1 3400
box 7 3 12 24
use welltap_svt  __well_tap__94
timestamp 1731220329
transform 1 0 104 0 -1 3400
box 7 3 12 24
use welltap_svt  __well_tap__93
timestamp 1731220329
transform 1 0 1760 0 1 3308
box 7 3 12 24
use welltap_svt  __well_tap__92
timestamp 1731220329
transform 1 0 104 0 1 3308
box 7 3 12 24
use welltap_svt  __well_tap__91
timestamp 1731220329
transform 1 0 1760 0 -1 3264
box 7 3 12 24
use welltap_svt  __well_tap__90
timestamp 1731220329
transform 1 0 104 0 -1 3264
box 7 3 12 24
use welltap_svt  __well_tap__89
timestamp 1731220329
transform 1 0 1760 0 1 3172
box 7 3 12 24
use welltap_svt  __well_tap__88
timestamp 1731220329
transform 1 0 104 0 1 3172
box 7 3 12 24
use welltap_svt  __well_tap__87
timestamp 1731220329
transform 1 0 1760 0 -1 3120
box 7 3 12 24
use welltap_svt  __well_tap__86
timestamp 1731220329
transform 1 0 104 0 -1 3120
box 7 3 12 24
use welltap_svt  __well_tap__85
timestamp 1731220329
transform 1 0 1760 0 1 3024
box 7 3 12 24
use welltap_svt  __well_tap__84
timestamp 1731220329
transform 1 0 104 0 1 3024
box 7 3 12 24
use welltap_svt  __well_tap__83
timestamp 1731220329
transform 1 0 1760 0 -1 2980
box 7 3 12 24
use welltap_svt  __well_tap__82
timestamp 1731220329
transform 1 0 104 0 -1 2980
box 7 3 12 24
use welltap_svt  __well_tap__81
timestamp 1731220329
transform 1 0 1760 0 1 2884
box 7 3 12 24
use welltap_svt  __well_tap__80
timestamp 1731220329
transform 1 0 104 0 1 2884
box 7 3 12 24
use welltap_svt  __well_tap__79
timestamp 1731220329
transform 1 0 1760 0 -1 2840
box 7 3 12 24
use welltap_svt  __well_tap__78
timestamp 1731220329
transform 1 0 104 0 -1 2840
box 7 3 12 24
use welltap_svt  __well_tap__77
timestamp 1731220329
transform 1 0 1760 0 1 2744
box 7 3 12 24
use welltap_svt  __well_tap__76
timestamp 1731220329
transform 1 0 104 0 1 2744
box 7 3 12 24
use welltap_svt  __well_tap__75
timestamp 1731220329
transform 1 0 1760 0 -1 2700
box 7 3 12 24
use welltap_svt  __well_tap__74
timestamp 1731220329
transform 1 0 104 0 -1 2700
box 7 3 12 24
use welltap_svt  __well_tap__73
timestamp 1731220329
transform 1 0 1760 0 1 2604
box 7 3 12 24
use welltap_svt  __well_tap__72
timestamp 1731220329
transform 1 0 104 0 1 2604
box 7 3 12 24
use welltap_svt  __well_tap__71
timestamp 1731220329
transform 1 0 1760 0 -1 2552
box 7 3 12 24
use welltap_svt  __well_tap__70
timestamp 1731220329
transform 1 0 104 0 -1 2552
box 7 3 12 24
use welltap_svt  __well_tap__69
timestamp 1731220329
transform 1 0 1760 0 1 2464
box 7 3 12 24
use welltap_svt  __well_tap__68
timestamp 1731220329
transform 1 0 104 0 1 2464
box 7 3 12 24
use welltap_svt  __well_tap__67
timestamp 1731220329
transform 1 0 1760 0 -1 2408
box 7 3 12 24
use welltap_svt  __well_tap__66
timestamp 1731220329
transform 1 0 104 0 -1 2408
box 7 3 12 24
use welltap_svt  __well_tap__65
timestamp 1731220329
transform 1 0 1760 0 1 2312
box 7 3 12 24
use welltap_svt  __well_tap__64
timestamp 1731220329
transform 1 0 104 0 1 2312
box 7 3 12 24
use welltap_svt  __well_tap__63
timestamp 1731220329
transform 1 0 1760 0 -1 2264
box 7 3 12 24
use welltap_svt  __well_tap__62
timestamp 1731220329
transform 1 0 104 0 -1 2264
box 7 3 12 24
use welltap_svt  __well_tap__61
timestamp 1731220329
transform 1 0 1760 0 1 2176
box 7 3 12 24
use welltap_svt  __well_tap__60
timestamp 1731220329
transform 1 0 104 0 1 2176
box 7 3 12 24
use welltap_svt  __well_tap__59
timestamp 1731220329
transform 1 0 1760 0 -1 2120
box 7 3 12 24
use welltap_svt  __well_tap__58
timestamp 1731220329
transform 1 0 104 0 -1 2120
box 7 3 12 24
use welltap_svt  __well_tap__57
timestamp 1731220329
transform 1 0 1760 0 1 2032
box 7 3 12 24
use welltap_svt  __well_tap__56
timestamp 1731220329
transform 1 0 104 0 1 2032
box 7 3 12 24
use welltap_svt  __well_tap__55
timestamp 1731220329
transform 1 0 1760 0 -1 1992
box 7 3 12 24
use welltap_svt  __well_tap__54
timestamp 1731220329
transform 1 0 104 0 -1 1992
box 7 3 12 24
use welltap_svt  __well_tap__53
timestamp 1731220329
transform 1 0 1760 0 1 1904
box 7 3 12 24
use welltap_svt  __well_tap__52
timestamp 1731220329
transform 1 0 104 0 1 1904
box 7 3 12 24
use welltap_svt  __well_tap__51
timestamp 1731220329
transform 1 0 1760 0 -1 1864
box 7 3 12 24
use welltap_svt  __well_tap__50
timestamp 1731220329
transform 1 0 104 0 -1 1864
box 7 3 12 24
use welltap_svt  __well_tap__49
timestamp 1731220329
transform 1 0 1760 0 1 1768
box 7 3 12 24
use welltap_svt  __well_tap__48
timestamp 1731220329
transform 1 0 104 0 1 1768
box 7 3 12 24
use welltap_svt  __well_tap__47
timestamp 1731220329
transform 1 0 1760 0 -1 1716
box 7 3 12 24
use welltap_svt  __well_tap__46
timestamp 1731220329
transform 1 0 104 0 -1 1716
box 7 3 12 24
use welltap_svt  __well_tap__45
timestamp 1731220329
transform 1 0 1760 0 1 1624
box 7 3 12 24
use welltap_svt  __well_tap__44
timestamp 1731220329
transform 1 0 104 0 1 1624
box 7 3 12 24
use welltap_svt  __well_tap__43
timestamp 1731220329
transform 1 0 1760 0 -1 1580
box 7 3 12 24
use welltap_svt  __well_tap__42
timestamp 1731220329
transform 1 0 104 0 -1 1580
box 7 3 12 24
use welltap_svt  __well_tap__41
timestamp 1731220329
transform 1 0 1760 0 1 1488
box 7 3 12 24
use welltap_svt  __well_tap__40
timestamp 1731220329
transform 1 0 104 0 1 1488
box 7 3 12 24
use welltap_svt  __well_tap__39
timestamp 1731220329
transform 1 0 1760 0 -1 1440
box 7 3 12 24
use welltap_svt  __well_tap__38
timestamp 1731220329
transform 1 0 104 0 -1 1440
box 7 3 12 24
use welltap_svt  __well_tap__37
timestamp 1731220329
transform 1 0 1760 0 1 1348
box 7 3 12 24
use welltap_svt  __well_tap__36
timestamp 1731220329
transform 1 0 104 0 1 1348
box 7 3 12 24
use welltap_svt  __well_tap__35
timestamp 1731220329
transform 1 0 1760 0 -1 1304
box 7 3 12 24
use welltap_svt  __well_tap__34
timestamp 1731220329
transform 1 0 104 0 -1 1304
box 7 3 12 24
use welltap_svt  __well_tap__33
timestamp 1731220329
transform 1 0 1760 0 1 1212
box 7 3 12 24
use welltap_svt  __well_tap__32
timestamp 1731220329
transform 1 0 104 0 1 1212
box 7 3 12 24
use welltap_svt  __well_tap__31
timestamp 1731220329
transform 1 0 1760 0 -1 1168
box 7 3 12 24
use welltap_svt  __well_tap__30
timestamp 1731220329
transform 1 0 104 0 -1 1168
box 7 3 12 24
use welltap_svt  __well_tap__29
timestamp 1731220329
transform 1 0 1760 0 1 1076
box 7 3 12 24
use welltap_svt  __well_tap__28
timestamp 1731220329
transform 1 0 104 0 1 1076
box 7 3 12 24
use welltap_svt  __well_tap__27
timestamp 1731220329
transform 1 0 1760 0 -1 1028
box 7 3 12 24
use welltap_svt  __well_tap__26
timestamp 1731220329
transform 1 0 104 0 -1 1028
box 7 3 12 24
use welltap_svt  __well_tap__25
timestamp 1731220329
transform 1 0 1760 0 1 936
box 7 3 12 24
use welltap_svt  __well_tap__24
timestamp 1731220329
transform 1 0 104 0 1 936
box 7 3 12 24
use welltap_svt  __well_tap__23
timestamp 1731220329
transform 1 0 1760 0 -1 892
box 7 3 12 24
use welltap_svt  __well_tap__22
timestamp 1731220329
transform 1 0 104 0 -1 892
box 7 3 12 24
use welltap_svt  __well_tap__21
timestamp 1731220329
transform 1 0 1760 0 1 800
box 7 3 12 24
use welltap_svt  __well_tap__20
timestamp 1731220329
transform 1 0 104 0 1 800
box 7 3 12 24
use welltap_svt  __well_tap__19
timestamp 1731220329
transform 1 0 1760 0 -1 756
box 7 3 12 24
use welltap_svt  __well_tap__18
timestamp 1731220329
transform 1 0 104 0 -1 756
box 7 3 12 24
use welltap_svt  __well_tap__17
timestamp 1731220329
transform 1 0 1760 0 1 660
box 7 3 12 24
use welltap_svt  __well_tap__16
timestamp 1731220329
transform 1 0 104 0 1 660
box 7 3 12 24
use welltap_svt  __well_tap__15
timestamp 1731220329
transform 1 0 1760 0 -1 616
box 7 3 12 24
use welltap_svt  __well_tap__14
timestamp 1731220329
transform 1 0 104 0 -1 616
box 7 3 12 24
use welltap_svt  __well_tap__13
timestamp 1731220329
transform 1 0 1760 0 1 524
box 7 3 12 24
use welltap_svt  __well_tap__12
timestamp 1731220329
transform 1 0 104 0 1 524
box 7 3 12 24
use welltap_svt  __well_tap__11
timestamp 1731220329
transform 1 0 1760 0 -1 480
box 7 3 12 24
use welltap_svt  __well_tap__10
timestamp 1731220329
transform 1 0 104 0 -1 480
box 7 3 12 24
use welltap_svt  __well_tap__9
timestamp 1731220329
transform 1 0 1760 0 1 388
box 7 3 12 24
use welltap_svt  __well_tap__8
timestamp 1731220329
transform 1 0 104 0 1 388
box 7 3 12 24
use welltap_svt  __well_tap__7
timestamp 1731220329
transform 1 0 1760 0 -1 344
box 7 3 12 24
use welltap_svt  __well_tap__6
timestamp 1731220329
transform 1 0 104 0 -1 344
box 7 3 12 24
use welltap_svt  __well_tap__5
timestamp 1731220329
transform 1 0 1760 0 1 252
box 7 3 12 24
use welltap_svt  __well_tap__4
timestamp 1731220329
transform 1 0 104 0 1 252
box 7 3 12 24
use welltap_svt  __well_tap__3
timestamp 1731220329
transform 1 0 1760 0 -1 208
box 7 3 12 24
use welltap_svt  __well_tap__2
timestamp 1731220329
transform 1 0 104 0 -1 208
box 7 3 12 24
use welltap_svt  __well_tap__1
timestamp 1731220329
transform 1 0 1760 0 1 96
box 7 3 12 24
use welltap_svt  __well_tap__0
timestamp 1731220329
transform 1 0 104 0 1 96
box 7 3 12 24
use _0_0cell_0_0gcelem2x0  tst_5999_6
timestamp 1731220329
transform 1 0 3240 0 1 3456
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5998_6
timestamp 1731220329
transform 1 0 3040 0 1 3456
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5997_6
timestamp 1731220329
transform 1 0 2848 0 1 3456
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5996_6
timestamp 1731220329
transform 1 0 2648 0 1 3456
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5995_6
timestamp 1731220329
transform 1 0 2968 0 -1 3456
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5994_6
timestamp 1731220329
transform 1 0 2840 0 -1 3456
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5993_6
timestamp 1731220329
transform 1 0 2712 0 -1 3456
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5992_6
timestamp 1731220329
transform 1 0 2592 0 -1 3456
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5991_6
timestamp 1731220329
transform 1 0 2472 0 -1 3456
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5990_6
timestamp 1731220329
transform 1 0 2512 0 1 3320
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5989_6
timestamp 1731220329
transform 1 0 2640 0 1 3320
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5988_6
timestamp 1731220329
transform 1 0 2768 0 1 3320
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5987_6
timestamp 1731220329
transform 1 0 3032 0 1 3320
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5986_6
timestamp 1731220329
transform 1 0 2896 0 1 3320
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5985_6
timestamp 1731220329
transform 1 0 2824 0 -1 3312
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5984_6
timestamp 1731220329
transform 1 0 2672 0 -1 3312
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5983_6
timestamp 1731220329
transform 1 0 2968 0 -1 3312
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5982_6
timestamp 1731220329
transform 1 0 3104 0 -1 3312
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5981_6
timestamp 1731220329
transform 1 0 3240 0 -1 3312
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5980_6
timestamp 1731220329
transform 1 0 3360 0 -1 3312
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5979_6
timestamp 1731220329
transform 1 0 3360 0 1 3176
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5978_6
timestamp 1731220329
transform 1 0 3360 0 -1 3176
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5977_6
timestamp 1731220329
transform 1 0 3256 0 -1 3176
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5976_6
timestamp 1731220329
transform 1 0 3360 0 1 3044
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5975_6
timestamp 1731220329
transform 1 0 3192 0 1 3044
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5974_6
timestamp 1731220329
transform 1 0 3128 0 -1 3176
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5973_6
timestamp 1731220329
transform 1 0 3000 0 -1 3176
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5972_6
timestamp 1731220329
transform 1 0 3200 0 1 3176
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5971_6
timestamp 1731220329
transform 1 0 3016 0 1 3176
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5970_6
timestamp 1731220329
transform 1 0 2832 0 1 3176
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5969_6
timestamp 1731220329
transform 1 0 2648 0 1 3176
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5968_6
timestamp 1731220329
transform 1 0 2568 0 -1 3176
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5967_6
timestamp 1731220329
transform 1 0 2728 0 -1 3176
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5966_6
timestamp 1731220329
transform 1 0 2872 0 -1 3176
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5965_6
timestamp 1731220329
transform 1 0 3024 0 1 3044
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5964_6
timestamp 1731220329
transform 1 0 2864 0 1 3044
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5963_6
timestamp 1731220329
transform 1 0 2712 0 1 3044
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5962_6
timestamp 1731220329
transform 1 0 2560 0 1 3044
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5961_6
timestamp 1731220329
transform 1 0 2752 0 -1 3036
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5960_6
timestamp 1731220329
transform 1 0 2640 0 -1 3036
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5959_6
timestamp 1731220329
transform 1 0 2536 0 -1 3036
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5958_6
timestamp 1731220329
transform 1 0 2432 0 -1 3036
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5957_6
timestamp 1731220329
transform 1 0 2664 0 1 2908
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5956_6
timestamp 1731220329
transform 1 0 2576 0 1 2908
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5955_6
timestamp 1731220329
transform 1 0 2488 0 1 2908
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5954_6
timestamp 1731220329
transform 1 0 2400 0 1 2908
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5953_6
timestamp 1731220329
transform 1 0 2224 0 1 2908
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5952_6
timestamp 1731220329
transform 1 0 2752 0 1 2908
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5951_6
timestamp 1731220329
transform 1 0 2840 0 1 2908
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5950_6
timestamp 1731220329
transform 1 0 2776 0 -1 2900
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5949_6
timestamp 1731220329
transform 1 0 2672 0 -1 2900
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5948_6
timestamp 1731220329
transform 1 0 2568 0 -1 2900
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5947_6
timestamp 1731220329
transform 1 0 2464 0 -1 2900
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5946_6
timestamp 1731220329
transform 1 0 2480 0 1 2768
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5945_6
timestamp 1731220329
transform 1 0 2600 0 1 2768
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5944_6
timestamp 1731220329
transform 1 0 2712 0 1 2768
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5943_6
timestamp 1731220329
transform 1 0 2952 0 1 2768
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5942_6
timestamp 1731220329
transform 1 0 2832 0 1 2768
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5941_6
timestamp 1731220329
transform 1 0 2760 0 -1 2764
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5940_6
timestamp 1731220329
transform 1 0 2616 0 -1 2764
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5939_6
timestamp 1731220329
transform 1 0 2904 0 -1 2764
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5938_6
timestamp 1731220329
transform 1 0 3048 0 -1 2764
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5937_6
timestamp 1731220329
transform 1 0 3088 0 1 2636
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5936_6
timestamp 1731220329
transform 1 0 2936 0 1 2636
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5935_6
timestamp 1731220329
transform 1 0 2776 0 1 2636
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5934_6
timestamp 1731220329
transform 1 0 2608 0 1 2636
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5933_6
timestamp 1731220329
transform 1 0 2512 0 -1 2632
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5932_6
timestamp 1731220329
transform 1 0 2664 0 -1 2632
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5931_6
timestamp 1731220329
transform 1 0 2800 0 -1 2632
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5930_6
timestamp 1731220329
transform 1 0 2920 0 -1 2632
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5929_6
timestamp 1731220329
transform 1 0 3040 0 -1 2632
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5928_6
timestamp 1731220329
transform 1 0 3152 0 -1 2632
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5927_6
timestamp 1731220329
transform 1 0 3264 0 -1 2632
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5926_6
timestamp 1731220329
transform 1 0 3232 0 1 2636
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5925_6
timestamp 1731220329
transform 1 0 3360 0 1 2636
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5924_6
timestamp 1731220329
transform 1 0 3360 0 -1 2632
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5923_6
timestamp 1731220329
transform 1 0 2792 0 1 2496
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5922_6
timestamp 1731220329
transform 1 0 3360 0 1 2496
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5921_6
timestamp 1731220329
transform 1 0 3360 0 -1 2480
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5920_6
timestamp 1731220329
transform 1 0 3360 0 1 2348
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5919_6
timestamp 1731220329
transform 1 0 3360 0 1 2216
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5918_6
timestamp 1731220329
transform 1 0 3360 0 -1 2204
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5917_6
timestamp 1731220329
transform 1 0 3360 0 -1 2060
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5916_6
timestamp 1731220329
transform 1 0 3360 0 -1 1912
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5915_6
timestamp 1731220329
transform 1 0 3360 0 -1 1768
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5914_6
timestamp 1731220329
transform 1 0 3360 0 1 1632
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5913_6
timestamp 1731220329
transform 1 0 3360 0 -1 1624
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5912_6
timestamp 1731220329
transform 1 0 3256 0 -1 1624
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5911_6
timestamp 1731220329
transform 1 0 3128 0 -1 1624
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5910_6
timestamp 1731220329
transform 1 0 3208 0 1 1632
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5909_6
timestamp 1731220329
transform 1 0 3336 0 1 1780
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5908_6
timestamp 1731220329
transform 1 0 3312 0 1 1916
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5907_6
timestamp 1731220329
transform 1 0 3360 0 1 2068
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5906_6
timestamp 1731220329
transform 1 0 3208 0 1 2216
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5905_6
timestamp 1731220329
transform 1 0 3248 0 -1 2348
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5904_6
timestamp 1731220329
transform 1 0 3168 0 1 2348
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5903_6
timestamp 1731220329
transform 1 0 3264 0 -1 2480
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5902_6
timestamp 1731220329
transform 1 0 3152 0 -1 2480
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5901_6
timestamp 1731220329
transform 1 0 3040 0 -1 2480
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5900_6
timestamp 1731220329
transform 1 0 2920 0 -1 2480
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5899_6
timestamp 1731220329
transform 1 0 2800 0 -1 2480
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5898_6
timestamp 1731220329
transform 1 0 2664 0 -1 2480
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5897_6
timestamp 1731220329
transform 1 0 2520 0 -1 2480
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5896_6
timestamp 1731220329
transform 1 0 2552 0 1 2348
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5895_6
timestamp 1731220329
transform 1 0 2752 0 1 2348
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5894_6
timestamp 1731220329
transform 1 0 2960 0 1 2348
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5893_6
timestamp 1731220329
transform 1 0 3040 0 -1 2348
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5892_6
timestamp 1731220329
transform 1 0 2832 0 -1 2348
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5891_6
timestamp 1731220329
transform 1 0 2640 0 -1 2348
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5890_6
timestamp 1731220329
transform 1 0 2456 0 -1 2348
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5889_6
timestamp 1731220329
transform 1 0 2584 0 1 2216
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5888_6
timestamp 1731220329
transform 1 0 2728 0 1 2216
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5887_6
timestamp 1731220329
transform 1 0 2880 0 1 2216
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5886_6
timestamp 1731220329
transform 1 0 3040 0 1 2216
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5885_6
timestamp 1731220329
transform 1 0 2960 0 -1 2204
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5884_6
timestamp 1731220329
transform 1 0 2832 0 -1 2204
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5883_6
timestamp 1731220329
transform 1 0 2712 0 -1 2204
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5882_6
timestamp 1731220329
transform 1 0 3240 0 -1 2204
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5881_6
timestamp 1731220329
transform 1 0 3096 0 -1 2204
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5880_6
timestamp 1731220329
transform 1 0 3024 0 1 2068
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5879_6
timestamp 1731220329
transform 1 0 2904 0 1 2068
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5878_6
timestamp 1731220329
transform 1 0 2776 0 1 2068
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5877_6
timestamp 1731220329
transform 1 0 3144 0 1 2068
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5876_6
timestamp 1731220329
transform 1 0 3264 0 1 2068
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5875_6
timestamp 1731220329
transform 1 0 3256 0 -1 2060
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5874_6
timestamp 1731220329
transform 1 0 3128 0 -1 2060
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5873_6
timestamp 1731220329
transform 1 0 3000 0 -1 2060
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5872_6
timestamp 1731220329
transform 1 0 2864 0 -1 2060
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5871_6
timestamp 1731220329
transform 1 0 2720 0 -1 2060
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5870_6
timestamp 1731220329
transform 1 0 3168 0 1 1916
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5869_6
timestamp 1731220329
transform 1 0 3024 0 1 1916
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5868_6
timestamp 1731220329
transform 1 0 2880 0 1 1916
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5867_6
timestamp 1731220329
transform 1 0 2744 0 1 1916
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5866_6
timestamp 1731220329
transform 1 0 2608 0 1 1916
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5865_6
timestamp 1731220329
transform 1 0 3176 0 -1 1912
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5864_6
timestamp 1731220329
transform 1 0 2976 0 -1 1912
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5863_6
timestamp 1731220329
transform 1 0 2784 0 -1 1912
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5862_6
timestamp 1731220329
transform 1 0 2608 0 -1 1912
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5861_6
timestamp 1731220329
transform 1 0 3128 0 1 1780
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5860_6
timestamp 1731220329
transform 1 0 2928 0 1 1780
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5859_6
timestamp 1731220329
transform 1 0 2736 0 1 1780
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5858_6
timestamp 1731220329
transform 1 0 2560 0 1 1780
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5857_6
timestamp 1731220329
transform 1 0 2400 0 1 1780
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5856_6
timestamp 1731220329
transform 1 0 2472 0 -1 1768
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5855_6
timestamp 1731220329
transform 1 0 2680 0 -1 1768
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5854_6
timestamp 1731220329
transform 1 0 3144 0 -1 1768
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5853_6
timestamp 1731220329
transform 1 0 2904 0 -1 1768
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5852_6
timestamp 1731220329
transform 1 0 2720 0 1 1632
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5851_6
timestamp 1731220329
transform 1 0 2568 0 1 1632
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5850_6
timestamp 1731220329
transform 1 0 2432 0 1 1632
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5849_6
timestamp 1731220329
transform 1 0 2880 0 1 1632
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5848_6
timestamp 1731220329
transform 1 0 3040 0 1 1632
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5847_6
timestamp 1731220329
transform 1 0 3008 0 -1 1624
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5846_6
timestamp 1731220329
transform 1 0 2888 0 -1 1624
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5845_6
timestamp 1731220329
transform 1 0 2760 0 -1 1624
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5844_6
timestamp 1731220329
transform 1 0 2632 0 -1 1624
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5843_6
timestamp 1731220329
transform 1 0 2496 0 -1 1624
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5842_6
timestamp 1731220329
transform 1 0 2592 0 1 1488
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5841_6
timestamp 1731220329
transform 1 0 2728 0 1 1488
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5840_6
timestamp 1731220329
transform 1 0 2864 0 1 1488
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5839_6
timestamp 1731220329
transform 1 0 3000 0 1 1488
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5838_6
timestamp 1731220329
transform 1 0 3136 0 1 1488
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5837_6
timestamp 1731220329
transform 1 0 3232 0 -1 1480
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5836_6
timestamp 1731220329
transform 1 0 3080 0 -1 1480
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5835_6
timestamp 1731220329
transform 1 0 2928 0 -1 1480
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5834_6
timestamp 1731220329
transform 1 0 2776 0 -1 1480
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5833_6
timestamp 1731220329
transform 1 0 2880 0 1 1344
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5832_6
timestamp 1731220329
transform 1 0 3024 0 1 1344
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5831_6
timestamp 1731220329
transform 1 0 3168 0 1 1344
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5830_6
timestamp 1731220329
transform 1 0 3320 0 1 1344
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5829_6
timestamp 1731220329
transform 1 0 3296 0 -1 1340
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5828_6
timestamp 1731220329
transform 1 0 3136 0 -1 1340
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5827_6
timestamp 1731220329
transform 1 0 2984 0 -1 1340
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5826_6
timestamp 1731220329
transform 1 0 2832 0 -1 1340
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5825_6
timestamp 1731220329
transform 1 0 3136 0 1 1212
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5824_6
timestamp 1731220329
transform 1 0 2968 0 1 1212
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5823_6
timestamp 1731220329
transform 1 0 2808 0 1 1212
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5822_6
timestamp 1731220329
transform 1 0 2688 0 -1 1212
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5821_6
timestamp 1731220329
transform 1 0 2840 0 -1 1212
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5820_6
timestamp 1731220329
transform 1 0 3152 0 -1 1212
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5819_6
timestamp 1731220329
transform 1 0 2992 0 -1 1212
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5818_6
timestamp 1731220329
transform 1 0 2864 0 1 1072
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5817_6
timestamp 1731220329
transform 1 0 2752 0 1 1072
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5816_6
timestamp 1731220329
transform 1 0 2632 0 1 1072
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5815_6
timestamp 1731220329
transform 1 0 2968 0 1 1072
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5814_6
timestamp 1731220329
transform 1 0 3072 0 1 1072
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5813_6
timestamp 1731220329
transform 1 0 3176 0 1 1072
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5812_6
timestamp 1731220329
transform 1 0 3272 0 1 1072
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5811_6
timestamp 1731220329
transform 1 0 3360 0 1 1072
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5810_6
timestamp 1731220329
transform 1 0 3360 0 1 936
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5809_6
timestamp 1731220329
transform 1 0 3360 0 -1 924
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5808_6
timestamp 1731220329
transform 1 0 3360 0 1 792
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5807_6
timestamp 1731220329
transform 1 0 3360 0 -1 788
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5806_6
timestamp 1731220329
transform 1 0 3360 0 -1 656
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5805_6
timestamp 1731220329
transform 1 0 3360 0 1 520
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5804_6
timestamp 1731220329
transform 1 0 3360 0 -1 516
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5803_6
timestamp 1731220329
transform 1 0 3360 0 1 380
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5802_6
timestamp 1731220329
transform 1 0 3360 0 -1 376
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5801_6
timestamp 1731220329
transform 1 0 3360 0 -1 240
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5800_6
timestamp 1731220329
transform 1 0 3360 0 1 92
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5799_6
timestamp 1731220329
transform 1 0 3272 0 1 92
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5798_6
timestamp 1731220329
transform 1 0 3160 0 1 92
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5797_6
timestamp 1731220329
transform 1 0 3200 0 -1 240
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5796_6
timestamp 1731220329
transform 1 0 3248 0 1 244
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5795_6
timestamp 1731220329
transform 1 0 3256 0 1 380
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5794_6
timestamp 1731220329
transform 1 0 3256 0 -1 516
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5793_6
timestamp 1731220329
transform 1 0 3128 0 -1 516
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5792_6
timestamp 1731220329
transform 1 0 3216 0 -1 656
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5791_6
timestamp 1731220329
transform 1 0 3048 0 -1 656
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5790_6
timestamp 1731220329
transform 1 0 3032 0 1 656
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5789_6
timestamp 1731220329
transform 1 0 2872 0 -1 656
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5788_6
timestamp 1731220329
transform 1 0 2680 0 -1 656
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5787_6
timestamp 1731220329
transform 1 0 2472 0 -1 656
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5786_6
timestamp 1731220329
transform 1 0 2864 0 1 520
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5785_6
timestamp 1731220329
transform 1 0 3192 0 1 520
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5784_6
timestamp 1731220329
transform 1 0 3024 0 1 520
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5783_6
timestamp 1731220329
transform 1 0 3000 0 -1 516
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5782_6
timestamp 1731220329
transform 1 0 2872 0 -1 516
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5781_6
timestamp 1731220329
transform 1 0 3136 0 1 380
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5780_6
timestamp 1731220329
transform 1 0 3016 0 1 380
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5779_6
timestamp 1731220329
transform 1 0 2904 0 1 380
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5778_6
timestamp 1731220329
transform 1 0 2904 0 -1 376
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5777_6
timestamp 1731220329
transform 1 0 3056 0 -1 376
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5776_6
timestamp 1731220329
transform 1 0 3216 0 -1 376
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5775_6
timestamp 1731220329
transform 1 0 3080 0 1 244
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5774_6
timestamp 1731220329
transform 1 0 2912 0 1 244
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5773_6
timestamp 1731220329
transform 1 0 2752 0 1 244
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5772_6
timestamp 1731220329
transform 1 0 2840 0 -1 240
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5771_6
timestamp 1731220329
transform 1 0 3016 0 -1 240
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5770_6
timestamp 1731220329
transform 1 0 3048 0 1 92
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5769_6
timestamp 1731220329
transform 1 0 2936 0 1 92
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5768_6
timestamp 1731220329
transform 1 0 2832 0 1 92
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5767_6
timestamp 1731220329
transform 1 0 2728 0 1 92
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5766_6
timestamp 1731220329
transform 1 0 2616 0 1 92
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5765_6
timestamp 1731220329
transform 1 0 2504 0 1 92
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5764_6
timestamp 1731220329
transform 1 0 2392 0 1 92
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5763_6
timestamp 1731220329
transform 1 0 2504 0 -1 240
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5762_6
timestamp 1731220329
transform 1 0 2672 0 -1 240
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5761_6
timestamp 1731220329
transform 1 0 2592 0 1 244
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5760_6
timestamp 1731220329
transform 1 0 2608 0 -1 376
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5759_6
timestamp 1731220329
transform 1 0 2752 0 -1 376
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5758_6
timestamp 1731220329
transform 1 0 2792 0 1 380
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5757_6
timestamp 1731220329
transform 1 0 2744 0 -1 516
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5756_6
timestamp 1731220329
transform 1 0 2712 0 1 520
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5755_6
timestamp 1731220329
transform 1 0 2560 0 1 520
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5754_6
timestamp 1731220329
transform 1 0 2560 0 1 656
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5753_6
timestamp 1731220329
transform 1 0 2712 0 1 656
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5752_6
timestamp 1731220329
transform 1 0 2872 0 1 656
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5751_6
timestamp 1731220329
transform 1 0 3192 0 1 656
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5750_6
timestamp 1731220329
transform 1 0 3208 0 -1 788
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5749_6
timestamp 1731220329
transform 1 0 3032 0 -1 788
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5748_6
timestamp 1731220329
transform 1 0 2864 0 -1 788
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5747_6
timestamp 1731220329
transform 1 0 2704 0 -1 788
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5746_6
timestamp 1731220329
transform 1 0 2552 0 -1 788
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5745_6
timestamp 1731220329
transform 1 0 3176 0 1 792
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5744_6
timestamp 1731220329
transform 1 0 2976 0 1 792
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5743_6
timestamp 1731220329
transform 1 0 2784 0 1 792
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5742_6
timestamp 1731220329
transform 1 0 2608 0 1 792
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5741_6
timestamp 1731220329
transform 1 0 2456 0 1 792
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5740_6
timestamp 1731220329
transform 1 0 2320 0 -1 924
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5739_6
timestamp 1731220329
transform 1 0 2512 0 -1 924
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5738_6
timestamp 1731220329
transform 1 0 2712 0 -1 924
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5737_6
timestamp 1731220329
transform 1 0 3152 0 -1 924
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5736_6
timestamp 1731220329
transform 1 0 2928 0 -1 924
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5735_6
timestamp 1731220329
transform 1 0 2744 0 1 936
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5734_6
timestamp 1731220329
transform 1 0 2616 0 1 936
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5733_6
timestamp 1731220329
transform 1 0 3216 0 1 936
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5732_6
timestamp 1731220329
transform 1 0 3048 0 1 936
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5731_6
timestamp 1731220329
transform 1 0 2888 0 1 936
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5730_6
timestamp 1731220329
transform 1 0 2800 0 -1 1064
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5729_6
timestamp 1731220329
transform 1 0 2712 0 -1 1064
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5728_6
timestamp 1731220329
transform 1 0 2624 0 -1 1064
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5727_6
timestamp 1731220329
transform 1 0 2536 0 -1 1064
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5726_6
timestamp 1731220329
transform 1 0 2504 0 1 1072
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5725_6
timestamp 1731220329
transform 1 0 2536 0 -1 1212
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5724_6
timestamp 1731220329
transform 1 0 2488 0 1 1212
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5723_6
timestamp 1731220329
transform 1 0 2648 0 1 1212
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5722_6
timestamp 1731220329
transform 1 0 2680 0 -1 1340
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5721_6
timestamp 1731220329
transform 1 0 2736 0 1 1344
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5720_6
timestamp 1731220329
transform 1 0 2624 0 -1 1480
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5719_6
timestamp 1731220329
transform 1 0 2448 0 1 1488
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5718_6
timestamp 1731220329
transform 1 0 2360 0 -1 1624
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5717_6
timestamp 1731220329
transform 1 0 2304 0 1 1632
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5716_6
timestamp 1731220329
transform 1 0 2296 0 -1 1768
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5715_6
timestamp 1731220329
transform 1 0 2248 0 1 1780
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5714_6
timestamp 1731220329
transform 1 0 2448 0 -1 1912
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5713_6
timestamp 1731220329
transform 1 0 2464 0 1 1916
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5712_6
timestamp 1731220329
transform 1 0 2568 0 -1 2060
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5711_6
timestamp 1731220329
transform 1 0 2408 0 -1 2060
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5710_6
timestamp 1731220329
transform 1 0 2240 0 -1 2060
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5709_6
timestamp 1731220329
transform 1 0 2128 0 1 2068
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5708_6
timestamp 1731220329
transform 1 0 2248 0 1 2068
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5707_6
timestamp 1731220329
transform 1 0 2376 0 1 2068
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5706_6
timestamp 1731220329
transform 1 0 2512 0 1 2068
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5705_6
timestamp 1731220329
transform 1 0 2648 0 1 2068
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5704_6
timestamp 1731220329
transform 1 0 2600 0 -1 2204
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5703_6
timestamp 1731220329
transform 1 0 2488 0 -1 2204
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5702_6
timestamp 1731220329
transform 1 0 2376 0 -1 2204
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5701_6
timestamp 1731220329
transform 1 0 2272 0 -1 2204
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5700_6
timestamp 1731220329
transform 1 0 2176 0 -1 2204
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5699_6
timestamp 1731220329
transform 1 0 2456 0 1 2216
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5698_6
timestamp 1731220329
transform 1 0 2336 0 1 2216
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5697_6
timestamp 1731220329
transform 1 0 2232 0 1 2216
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5696_6
timestamp 1731220329
transform 1 0 2128 0 1 2216
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5695_6
timestamp 1731220329
transform 1 0 2032 0 1 2216
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5694_6
timestamp 1731220329
transform 1 0 2296 0 -1 2348
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5693_6
timestamp 1731220329
transform 1 0 2144 0 -1 2348
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5692_6
timestamp 1731220329
transform 1 0 2008 0 -1 2348
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5691_6
timestamp 1731220329
transform 1 0 1880 0 -1 2348
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5690_6
timestamp 1731220329
transform 1 0 1832 0 1 2348
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5689_6
timestamp 1731220329
transform 1 0 2000 0 1 2348
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5688_6
timestamp 1731220329
transform 1 0 2176 0 1 2348
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5687_6
timestamp 1731220329
transform 1 0 2360 0 1 2348
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5686_6
timestamp 1731220329
transform 1 0 2360 0 -1 2480
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5685_6
timestamp 1731220329
transform 1 0 2192 0 -1 2480
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5684_6
timestamp 1731220329
transform 1 0 2008 0 -1 2480
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5683_6
timestamp 1731220329
transform 1 0 2200 0 1 2496
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5682_6
timestamp 1731220329
transform 1 0 2352 0 -1 2632
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5681_6
timestamp 1731220329
transform 1 0 2424 0 1 2636
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5680_6
timestamp 1731220329
transform 1 0 2472 0 -1 2764
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5679_6
timestamp 1731220329
transform 1 0 2328 0 -1 2764
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5678_6
timestamp 1731220329
transform 1 0 2360 0 1 2768
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5677_6
timestamp 1731220329
transform 1 0 2360 0 -1 2900
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5676_6
timestamp 1731220329
transform 1 0 2312 0 1 2908
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5675_6
timestamp 1731220329
transform 1 0 2328 0 -1 3036
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5674_6
timestamp 1731220329
transform 1 0 2296 0 1 3044
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5673_6
timestamp 1731220329
transform 1 0 2424 0 1 3044
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5672_6
timestamp 1731220329
transform 1 0 2400 0 -1 3176
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5671_6
timestamp 1731220329
transform 1 0 2448 0 1 3176
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5670_6
timestamp 1731220329
transform 1 0 2240 0 1 3176
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5669_6
timestamp 1731220329
transform 1 0 2328 0 -1 3312
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5668_6
timestamp 1731220329
transform 1 0 2504 0 -1 3312
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5667_6
timestamp 1731220329
transform 1 0 2376 0 1 3320
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5666_6
timestamp 1731220329
transform 1 0 2232 0 1 3320
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5665_6
timestamp 1731220329
transform 1 0 2208 0 -1 3456
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5664_6
timestamp 1731220329
transform 1 0 2344 0 -1 3456
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5663_6
timestamp 1731220329
transform 1 0 2448 0 1 3456
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5662_6
timestamp 1731220329
transform 1 0 2232 0 1 3456
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5661_6
timestamp 1731220329
transform 1 0 2000 0 1 3456
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5660_6
timestamp 1731220329
transform 1 0 1936 0 -1 3456
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5659_6
timestamp 1731220329
transform 1 0 1824 0 -1 3456
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5658_6
timestamp 1731220329
transform 1 0 2072 0 -1 3456
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5657_6
timestamp 1731220329
transform 1 0 2088 0 1 3320
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5656_6
timestamp 1731220329
transform 1 0 1944 0 1 3320
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5655_6
timestamp 1731220329
transform 1 0 1824 0 1 3320
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5654_6
timestamp 1731220329
transform 1 0 1824 0 -1 3312
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5653_6
timestamp 1731220329
transform 1 0 1968 0 -1 3312
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5652_6
timestamp 1731220329
transform 1 0 2144 0 -1 3312
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5651_6
timestamp 1731220329
transform 1 0 2024 0 1 3176
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5650_6
timestamp 1731220329
transform 1 0 1824 0 1 3176
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5649_6
timestamp 1731220329
transform 1 0 1832 0 -1 3176
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5648_6
timestamp 1731220329
transform 1 0 2024 0 -1 3176
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5647_6
timestamp 1731220329
transform 1 0 2216 0 -1 3176
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5646_6
timestamp 1731220329
transform 1 0 2168 0 1 3044
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5645_6
timestamp 1731220329
transform 1 0 2048 0 1 3044
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5644_6
timestamp 1731220329
transform 1 0 1928 0 1 3044
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5643_6
timestamp 1731220329
transform 1 0 2016 0 -1 3036
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5642_6
timestamp 1731220329
transform 1 0 2224 0 -1 3036
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5641_6
timestamp 1731220329
transform 1 0 2120 0 -1 3036
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5640_6
timestamp 1731220329
transform 1 0 2048 0 1 2908
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5639_6
timestamp 1731220329
transform 1 0 2136 0 1 2908
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5638_6
timestamp 1731220329
transform 1 0 2264 0 -1 2900
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5637_6
timestamp 1731220329
transform 1 0 2168 0 -1 2900
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5636_6
timestamp 1731220329
transform 1 0 2064 0 -1 2900
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5635_6
timestamp 1731220329
transform 1 0 1976 0 1 2768
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5634_6
timestamp 1731220329
transform 1 0 2104 0 1 2768
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5633_6
timestamp 1731220329
transform 1 0 2232 0 1 2768
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5632_6
timestamp 1731220329
transform 1 0 2176 0 -1 2764
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5631_6
timestamp 1731220329
transform 1 0 2024 0 -1 2764
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5630_6
timestamp 1731220329
transform 1 0 1880 0 -1 2764
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5629_6
timestamp 1731220329
transform 1 0 1824 0 1 2636
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5628_6
timestamp 1731220329
transform 1 0 2016 0 1 2636
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5627_6
timestamp 1731220329
transform 1 0 2224 0 1 2636
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5626_6
timestamp 1731220329
transform 1 0 2176 0 -1 2632
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5625_6
timestamp 1731220329
transform 1 0 1992 0 -1 2632
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5624_6
timestamp 1731220329
transform 1 0 1824 0 -1 2632
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5623_6
timestamp 1731220329
transform 1 0 1664 0 -1 2572
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5622_6
timestamp 1731220329
transform 1 0 1576 0 -1 2572
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5621_6
timestamp 1731220329
transform 1 0 1488 0 -1 2572
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5620_6
timestamp 1731220329
transform 1 0 1400 0 -1 2572
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5619_6
timestamp 1731220329
transform 1 0 1664 0 1 2444
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5618_6
timestamp 1731220329
transform 1 0 1568 0 1 2444
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5617_6
timestamp 1731220329
transform 1 0 1456 0 1 2444
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5616_6
timestamp 1731220329
transform 1 0 1304 0 -1 2572
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5615_6
timestamp 1731220329
transform 1 0 1208 0 -1 2572
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5614_6
timestamp 1731220329
transform 1 0 1112 0 -1 2572
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5613_6
timestamp 1731220329
transform 1 0 1024 0 -1 2572
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5612_6
timestamp 1731220329
transform 1 0 936 0 -1 2572
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5611_6
timestamp 1731220329
transform 1 0 848 0 -1 2572
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5610_6
timestamp 1731220329
transform 1 0 1096 0 1 2444
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5609_6
timestamp 1731220329
transform 1 0 1224 0 1 2444
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5608_6
timestamp 1731220329
transform 1 0 1344 0 1 2444
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5607_6
timestamp 1731220329
transform 1 0 1232 0 -1 2428
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5606_6
timestamp 1731220329
transform 1 0 1408 0 -1 2428
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5605_6
timestamp 1731220329
transform 1 0 1584 0 -1 2428
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5604_6
timestamp 1731220329
transform 1 0 1504 0 1 2292
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5603_6
timestamp 1731220329
transform 1 0 1368 0 1 2292
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5602_6
timestamp 1731220329
transform 1 0 1232 0 1 2292
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5601_6
timestamp 1731220329
transform 1 0 1184 0 -1 2284
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5600_6
timestamp 1731220329
transform 1 0 1296 0 -1 2284
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5599_6
timestamp 1731220329
transform 1 0 1408 0 -1 2284
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5598_6
timestamp 1731220329
transform 1 0 1312 0 1 2156
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5597_6
timestamp 1731220329
transform 1 0 1224 0 1 2156
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5596_6
timestamp 1731220329
transform 1 0 1136 0 1 2156
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5595_6
timestamp 1731220329
transform 1 0 1048 0 1 2156
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5594_6
timestamp 1731220329
transform 1 0 960 0 1 2156
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5593_6
timestamp 1731220329
transform 1 0 872 0 1 2156
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5592_6
timestamp 1731220329
transform 1 0 656 0 -1 2284
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5591_6
timestamp 1731220329
transform 1 0 568 0 -1 2284
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5590_6
timestamp 1731220329
transform 1 0 712 0 1 2292
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5589_6
timestamp 1731220329
transform 1 0 592 0 1 2292
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5588_6
timestamp 1731220329
transform 1 0 472 0 1 2292
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5587_6
timestamp 1731220329
transform 1 0 368 0 1 2292
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5586_6
timestamp 1731220329
transform 1 0 712 0 -1 2428
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5585_6
timestamp 1731220329
transform 1 0 544 0 -1 2428
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5584_6
timestamp 1731220329
transform 1 0 384 0 -1 2428
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5583_6
timestamp 1731220329
transform 1 0 232 0 -1 2428
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5582_6
timestamp 1731220329
transform 1 0 128 0 -1 2428
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5581_6
timestamp 1731220329
transform 1 0 128 0 1 2444
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5580_6
timestamp 1731220329
transform 1 0 240 0 1 2444
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5579_6
timestamp 1731220329
transform 1 0 688 0 1 2444
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5578_6
timestamp 1731220329
transform 1 0 536 0 1 2444
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5577_6
timestamp 1731220329
transform 1 0 384 0 1 2444
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5576_6
timestamp 1731220329
transform 1 0 304 0 -1 2572
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5575_6
timestamp 1731220329
transform 1 0 216 0 -1 2572
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5574_6
timestamp 1731220329
transform 1 0 400 0 -1 2572
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5573_6
timestamp 1731220329
transform 1 0 584 0 -1 2572
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5572_6
timestamp 1731220329
transform 1 0 496 0 -1 2572
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5571_6
timestamp 1731220329
transform 1 0 464 0 1 2584
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5570_6
timestamp 1731220329
transform 1 0 552 0 1 2584
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5569_6
timestamp 1731220329
transform 1 0 640 0 1 2584
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5568_6
timestamp 1731220329
transform 1 0 728 0 1 2584
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5567_6
timestamp 1731220329
transform 1 0 816 0 1 2584
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5566_6
timestamp 1731220329
transform 1 0 824 0 -1 2720
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5565_6
timestamp 1731220329
transform 1 0 736 0 -1 2720
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5564_6
timestamp 1731220329
transform 1 0 648 0 -1 2720
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5563_6
timestamp 1731220329
transform 1 0 560 0 -1 2720
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5562_6
timestamp 1731220329
transform 1 0 472 0 -1 2720
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5561_6
timestamp 1731220329
transform 1 0 736 0 1 2724
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5560_6
timestamp 1731220329
transform 1 0 616 0 1 2724
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5559_6
timestamp 1731220329
transform 1 0 496 0 1 2724
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5558_6
timestamp 1731220329
transform 1 0 384 0 1 2724
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5557_6
timestamp 1731220329
transform 1 0 280 0 1 2724
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5556_6
timestamp 1731220329
transform 1 0 720 0 -1 2860
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5555_6
timestamp 1731220329
transform 1 0 560 0 -1 2860
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5554_6
timestamp 1731220329
transform 1 0 400 0 -1 2860
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5553_6
timestamp 1731220329
transform 1 0 248 0 -1 2860
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5552_6
timestamp 1731220329
transform 1 0 128 0 -1 2860
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5551_6
timestamp 1731220329
transform 1 0 776 0 1 2864
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5550_6
timestamp 1731220329
transform 1 0 600 0 1 2864
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5549_6
timestamp 1731220329
transform 1 0 424 0 1 2864
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5548_6
timestamp 1731220329
transform 1 0 256 0 1 2864
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5547_6
timestamp 1731220329
transform 1 0 128 0 1 2864
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5546_6
timestamp 1731220329
transform 1 0 128 0 -1 3000
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5545_6
timestamp 1731220329
transform 1 0 728 0 -1 3000
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5544_6
timestamp 1731220329
transform 1 0 528 0 -1 3000
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5543_6
timestamp 1731220329
transform 1 0 320 0 -1 3000
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5542_6
timestamp 1731220329
transform 1 0 256 0 1 3004
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5541_6
timestamp 1731220329
transform 1 0 128 0 1 3004
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5540_6
timestamp 1731220329
transform 1 0 784 0 1 3004
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5539_6
timestamp 1731220329
transform 1 0 600 0 1 3004
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5538_6
timestamp 1731220329
transform 1 0 424 0 1 3004
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5537_6
timestamp 1731220329
transform 1 0 312 0 -1 3140
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5536_6
timestamp 1731220329
transform 1 0 168 0 -1 3140
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5535_6
timestamp 1731220329
transform 1 0 768 0 -1 3140
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5534_6
timestamp 1731220329
transform 1 0 616 0 -1 3140
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5533_6
timestamp 1731220329
transform 1 0 464 0 -1 3140
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5532_6
timestamp 1731220329
transform 1 0 416 0 1 3152
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5531_6
timestamp 1731220329
transform 1 0 296 0 1 3152
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5530_6
timestamp 1731220329
transform 1 0 792 0 1 3152
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5529_6
timestamp 1731220329
transform 1 0 664 0 1 3152
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5528_6
timestamp 1731220329
transform 1 0 536 0 1 3152
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5527_6
timestamp 1731220329
transform 1 0 488 0 -1 3284
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5526_6
timestamp 1731220329
transform 1 0 376 0 -1 3284
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5525_6
timestamp 1731220329
transform 1 0 600 0 -1 3284
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5524_6
timestamp 1731220329
transform 1 0 720 0 -1 3284
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5523_6
timestamp 1731220329
transform 1 0 840 0 -1 3284
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5522_6
timestamp 1731220329
transform 1 0 800 0 1 3288
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5521_6
timestamp 1731220329
transform 1 0 696 0 1 3288
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5520_6
timestamp 1731220329
transform 1 0 592 0 1 3288
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5519_6
timestamp 1731220329
transform 1 0 488 0 1 3288
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5518_6
timestamp 1731220329
transform 1 0 392 0 1 3288
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5517_6
timestamp 1731220329
transform 1 0 408 0 -1 3420
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5516_6
timestamp 1731220329
transform 1 0 496 0 -1 3420
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5515_6
timestamp 1731220329
transform 1 0 760 0 -1 3420
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5514_6
timestamp 1731220329
transform 1 0 672 0 -1 3420
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5513_6
timestamp 1731220329
transform 1 0 584 0 -1 3420
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5512_6
timestamp 1731220329
transform 1 0 536 0 1 3420
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5511_6
timestamp 1731220329
transform 1 0 448 0 1 3420
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5510_6
timestamp 1731220329
transform 1 0 624 0 1 3420
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5509_6
timestamp 1731220329
transform 1 0 712 0 1 3420
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5508_6
timestamp 1731220329
transform 1 0 800 0 1 3420
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5507_6
timestamp 1731220329
transform 1 0 888 0 1 3420
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5506_6
timestamp 1731220329
transform 1 0 976 0 1 3420
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5505_6
timestamp 1731220329
transform 1 0 1152 0 1 3420
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5504_6
timestamp 1731220329
transform 1 0 1064 0 1 3420
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5503_6
timestamp 1731220329
transform 1 0 1024 0 -1 3420
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5502_6
timestamp 1731220329
transform 1 0 936 0 -1 3420
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5501_6
timestamp 1731220329
transform 1 0 848 0 -1 3420
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5500_6
timestamp 1731220329
transform 1 0 1112 0 -1 3420
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5499_6
timestamp 1731220329
transform 1 0 1296 0 -1 3420
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5498_6
timestamp 1731220329
transform 1 0 1200 0 -1 3420
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5497_6
timestamp 1731220329
transform 1 0 1112 0 1 3288
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5496_6
timestamp 1731220329
transform 1 0 1008 0 1 3288
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5495_6
timestamp 1731220329
transform 1 0 904 0 1 3288
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5494_6
timestamp 1731220329
transform 1 0 1216 0 1 3288
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5493_6
timestamp 1731220329
transform 1 0 1320 0 1 3288
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5492_6
timestamp 1731220329
transform 1 0 1328 0 -1 3284
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5491_6
timestamp 1731220329
transform 1 0 1200 0 -1 3284
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5490_6
timestamp 1731220329
transform 1 0 1080 0 -1 3284
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5489_6
timestamp 1731220329
transform 1 0 960 0 -1 3284
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5488_6
timestamp 1731220329
transform 1 0 920 0 1 3152
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5487_6
timestamp 1731220329
transform 1 0 1048 0 1 3152
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5486_6
timestamp 1731220329
transform 1 0 1168 0 1 3152
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5485_6
timestamp 1731220329
transform 1 0 1424 0 1 3152
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5484_6
timestamp 1731220329
transform 1 0 1296 0 1 3152
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5483_6
timestamp 1731220329
transform 1 0 1192 0 -1 3140
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5482_6
timestamp 1731220329
transform 1 0 1056 0 -1 3140
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5481_6
timestamp 1731220329
transform 1 0 912 0 -1 3140
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5480_6
timestamp 1731220329
transform 1 0 1336 0 -1 3140
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5479_6
timestamp 1731220329
transform 1 0 1480 0 -1 3140
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5478_6
timestamp 1731220329
transform 1 0 1504 0 1 3004
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5477_6
timestamp 1731220329
transform 1 0 1320 0 1 3004
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5476_6
timestamp 1731220329
transform 1 0 1136 0 1 3004
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5475_6
timestamp 1731220329
transform 1 0 960 0 1 3004
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5474_6
timestamp 1731220329
transform 1 0 920 0 -1 3000
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5473_6
timestamp 1731220329
transform 1 0 1096 0 -1 3000
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5472_6
timestamp 1731220329
transform 1 0 1272 0 -1 3000
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5471_6
timestamp 1731220329
transform 1 0 1440 0 -1 3000
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5470_6
timestamp 1731220329
transform 1 0 1616 0 -1 3000
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5469_6
timestamp 1731220329
transform 1 0 1584 0 1 2864
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5468_6
timestamp 1731220329
transform 1 0 1424 0 1 2864
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5467_6
timestamp 1731220329
transform 1 0 1264 0 1 2864
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5466_6
timestamp 1731220329
transform 1 0 1104 0 1 2864
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5465_6
timestamp 1731220329
transform 1 0 944 0 1 2864
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5464_6
timestamp 1731220329
transform 1 0 1456 0 -1 2860
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5463_6
timestamp 1731220329
transform 1 0 1304 0 -1 2860
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5462_6
timestamp 1731220329
transform 1 0 1160 0 -1 2860
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5461_6
timestamp 1731220329
transform 1 0 1016 0 -1 2860
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5460_6
timestamp 1731220329
transform 1 0 872 0 -1 2860
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5459_6
timestamp 1731220329
transform 1 0 1312 0 1 2724
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5458_6
timestamp 1731220329
transform 1 0 1192 0 1 2724
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5457_6
timestamp 1731220329
transform 1 0 1072 0 1 2724
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5456_6
timestamp 1731220329
transform 1 0 960 0 1 2724
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5455_6
timestamp 1731220329
transform 1 0 848 0 1 2724
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5454_6
timestamp 1731220329
transform 1 0 1176 0 -1 2720
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5453_6
timestamp 1731220329
transform 1 0 1088 0 -1 2720
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5452_6
timestamp 1731220329
transform 1 0 1000 0 -1 2720
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5451_6
timestamp 1731220329
transform 1 0 912 0 -1 2720
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5450_6
timestamp 1731220329
transform 1 0 1080 0 1 2584
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5449_6
timestamp 1731220329
transform 1 0 992 0 1 2584
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5448_6
timestamp 1731220329
transform 1 0 904 0 1 2584
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5447_6
timestamp 1731220329
transform 1 0 760 0 -1 2572
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5446_6
timestamp 1731220329
transform 1 0 672 0 -1 2572
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5445_6
timestamp 1731220329
transform 1 0 832 0 1 2444
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5444_6
timestamp 1731220329
transform 1 0 968 0 1 2444
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5443_6
timestamp 1731220329
transform 1 0 1056 0 -1 2428
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5442_6
timestamp 1731220329
transform 1 0 888 0 -1 2428
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5441_6
timestamp 1731220329
transform 1 0 840 0 1 2292
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5440_6
timestamp 1731220329
transform 1 0 968 0 1 2292
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5439_6
timestamp 1731220329
transform 1 0 1096 0 1 2292
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5438_6
timestamp 1731220329
transform 1 0 1072 0 -1 2284
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5437_6
timestamp 1731220329
transform 1 0 960 0 -1 2284
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5436_6
timestamp 1731220329
transform 1 0 856 0 -1 2284
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5435_6
timestamp 1731220329
transform 1 0 752 0 -1 2284
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5434_6
timestamp 1731220329
transform 1 0 784 0 1 2156
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5433_6
timestamp 1731220329
transform 1 0 696 0 1 2156
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5432_6
timestamp 1731220329
transform 1 0 608 0 1 2156
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5431_6
timestamp 1731220329
transform 1 0 520 0 1 2156
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5430_6
timestamp 1731220329
transform 1 0 432 0 1 2156
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5429_6
timestamp 1731220329
transform 1 0 624 0 -1 2140
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5428_6
timestamp 1731220329
transform 1 0 512 0 -1 2140
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5427_6
timestamp 1731220329
transform 1 0 400 0 -1 2140
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5426_6
timestamp 1731220329
transform 1 0 296 0 -1 2140
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5425_6
timestamp 1731220329
transform 1 0 248 0 1 2012
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5424_6
timestamp 1731220329
transform 1 0 368 0 1 2012
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5423_6
timestamp 1731220329
transform 1 0 488 0 1 2012
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5422_6
timestamp 1731220329
transform 1 0 480 0 -1 2012
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5421_6
timestamp 1731220329
transform 1 0 352 0 -1 2012
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5420_6
timestamp 1731220329
transform 1 0 616 0 -1 2012
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5419_6
timestamp 1731220329
transform 1 0 704 0 1 1884
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5418_6
timestamp 1731220329
transform 1 0 568 0 1 1884
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5417_6
timestamp 1731220329
transform 1 0 440 0 1 1884
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5416_6
timestamp 1731220329
transform 1 0 552 0 -1 1884
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5415_6
timestamp 1731220329
transform 1 0 688 0 -1 1884
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5414_6
timestamp 1731220329
transform 1 0 824 0 -1 1884
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5413_6
timestamp 1731220329
transform 1 0 840 0 1 1884
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5412_6
timestamp 1731220329
transform 1 0 976 0 1 1884
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5411_6
timestamp 1731220329
transform 1 0 888 0 -1 2012
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5410_6
timestamp 1731220329
transform 1 0 752 0 -1 2012
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5409_6
timestamp 1731220329
transform 1 0 720 0 1 2012
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5408_6
timestamp 1731220329
transform 1 0 608 0 1 2012
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5407_6
timestamp 1731220329
transform 1 0 736 0 -1 2140
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5406_6
timestamp 1731220329
transform 1 0 856 0 -1 2140
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5405_6
timestamp 1731220329
transform 1 0 976 0 -1 2140
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5404_6
timestamp 1731220329
transform 1 0 928 0 1 2012
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5403_6
timestamp 1731220329
transform 1 0 824 0 1 2012
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5402_6
timestamp 1731220329
transform 1 0 1032 0 1 2012
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5401_6
timestamp 1731220329
transform 1 0 1136 0 1 2012
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5400_6
timestamp 1731220329
transform 1 0 1248 0 1 2012
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5399_6
timestamp 1731220329
transform 1 0 1144 0 -1 2012
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5398_6
timestamp 1731220329
transform 1 0 1016 0 -1 2012
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5397_6
timestamp 1731220329
transform 1 0 1264 0 -1 2012
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5396_6
timestamp 1731220329
transform 1 0 1392 0 -1 2012
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5395_6
timestamp 1731220329
transform 1 0 1520 0 -1 2012
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5394_6
timestamp 1731220329
transform 1 0 1648 0 1 1884
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5393_6
timestamp 1731220329
transform 1 0 1512 0 1 1884
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5392_6
timestamp 1731220329
transform 1 0 1376 0 1 1884
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5391_6
timestamp 1731220329
transform 1 0 1248 0 1 1884
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5390_6
timestamp 1731220329
transform 1 0 1112 0 1 1884
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5389_6
timestamp 1731220329
transform 1 0 1448 0 -1 1884
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5388_6
timestamp 1731220329
transform 1 0 1320 0 -1 1884
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5387_6
timestamp 1731220329
transform 1 0 1192 0 -1 1884
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5386_6
timestamp 1731220329
transform 1 0 1072 0 -1 1884
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5385_6
timestamp 1731220329
transform 1 0 952 0 -1 1884
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5384_6
timestamp 1731220329
transform 1 0 1232 0 1 1748
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5383_6
timestamp 1731220329
transform 1 0 1080 0 1 1748
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5382_6
timestamp 1731220329
transform 1 0 936 0 1 1748
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5381_6
timestamp 1731220329
transform 1 0 928 0 -1 1736
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5380_6
timestamp 1731220329
transform 1 0 1112 0 -1 1736
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5379_6
timestamp 1731220329
transform 1 0 1224 0 1 1604
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5378_6
timestamp 1731220329
transform 1 0 1032 0 1 1604
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5377_6
timestamp 1731220329
transform 1 0 848 0 1 1604
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5376_6
timestamp 1731220329
transform 1 0 960 0 -1 1600
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5375_6
timestamp 1731220329
transform 1 0 1112 0 -1 1600
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5374_6
timestamp 1731220329
transform 1 0 1192 0 1 1468
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5373_6
timestamp 1731220329
transform 1 0 1040 0 1 1468
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5372_6
timestamp 1731220329
transform 1 0 888 0 1 1468
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5371_6
timestamp 1731220329
transform 1 0 1056 0 -1 1460
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5370_6
timestamp 1731220329
transform 1 0 920 0 -1 1460
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5369_6
timestamp 1731220329
transform 1 0 896 0 1 1328
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5368_6
timestamp 1731220329
transform 1 0 1024 0 1 1328
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5367_6
timestamp 1731220329
transform 1 0 1152 0 1 1328
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5366_6
timestamp 1731220329
transform 1 0 1184 0 -1 1324
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5365_6
timestamp 1731220329
transform 1 0 1304 0 -1 1324
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5364_6
timestamp 1731220329
transform 1 0 1408 0 1 1328
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5363_6
timestamp 1731220329
transform 1 0 1280 0 1 1328
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5362_6
timestamp 1731220329
transform 1 0 1192 0 -1 1460
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5361_6
timestamp 1731220329
transform 1 0 1328 0 -1 1460
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5360_6
timestamp 1731220329
transform 1 0 1464 0 -1 1460
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5359_6
timestamp 1731220329
transform 1 0 1496 0 1 1468
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5358_6
timestamp 1731220329
transform 1 0 1344 0 1 1468
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5357_6
timestamp 1731220329
transform 1 0 1272 0 -1 1600
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5356_6
timestamp 1731220329
transform 1 0 1600 0 -1 1600
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5355_6
timestamp 1731220329
transform 1 0 1432 0 -1 1600
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5354_6
timestamp 1731220329
transform 1 0 1424 0 1 1604
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5353_6
timestamp 1731220329
transform 1 0 1632 0 1 1604
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5352_6
timestamp 1731220329
transform 1 0 1664 0 -1 1736
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5351_6
timestamp 1731220329
transform 1 0 1496 0 -1 1736
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5350_6
timestamp 1731220329
transform 1 0 1304 0 -1 1736
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5349_6
timestamp 1731220329
transform 1 0 1384 0 1 1748
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5348_6
timestamp 1731220329
transform 1 0 1536 0 1 1748
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5347_6
timestamp 1731220329
transform 1 0 1664 0 1 1748
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5346_6
timestamp 1731220329
transform 1 0 1824 0 1 1780
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5345_6
timestamp 1731220329
transform 1 0 1824 0 -1 1912
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5344_6
timestamp 1731220329
transform 1 0 1912 0 -1 1912
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5343_6
timestamp 1731220329
transform 1 0 1824 0 1 1916
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5342_6
timestamp 1731220329
transform 1 0 1912 0 1 1916
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5341_6
timestamp 1731220329
transform 1 0 2040 0 1 1916
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5340_6
timestamp 1731220329
transform 1 0 2176 0 1 1916
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5339_6
timestamp 1731220329
transform 1 0 2320 0 1 1916
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5338_6
timestamp 1731220329
transform 1 0 2296 0 -1 1912
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5337_6
timestamp 1731220329
transform 1 0 2160 0 -1 1912
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5336_6
timestamp 1731220329
transform 1 0 2032 0 -1 1912
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5335_6
timestamp 1731220329
transform 1 0 2104 0 1 1780
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5334_6
timestamp 1731220329
transform 1 0 1952 0 1 1780
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5333_6
timestamp 1731220329
transform 1 0 1872 0 -1 1768
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5332_6
timestamp 1731220329
transform 1 0 2008 0 -1 1768
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5331_6
timestamp 1731220329
transform 1 0 2144 0 -1 1768
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5330_6
timestamp 1731220329
transform 1 0 2176 0 1 1632
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5329_6
timestamp 1731220329
transform 1 0 2056 0 1 1632
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5328_6
timestamp 1731220329
transform 1 0 1928 0 1 1632
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5327_6
timestamp 1731220329
transform 1 0 1824 0 1 1632
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5326_6
timestamp 1731220329
transform 1 0 1824 0 -1 1624
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5325_6
timestamp 1731220329
transform 1 0 1936 0 -1 1624
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5324_6
timestamp 1731220329
transform 1 0 2080 0 -1 1624
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5323_6
timestamp 1731220329
transform 1 0 2224 0 -1 1624
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5322_6
timestamp 1731220329
transform 1 0 2296 0 1 1488
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5321_6
timestamp 1731220329
transform 1 0 2144 0 1 1488
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5320_6
timestamp 1731220329
transform 1 0 1984 0 1 1488
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5319_6
timestamp 1731220329
transform 1 0 1832 0 1 1488
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5318_6
timestamp 1731220329
transform 1 0 1936 0 -1 1480
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5317_6
timestamp 1731220329
transform 1 0 2048 0 -1 1480
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5316_6
timestamp 1731220329
transform 1 0 2184 0 -1 1480
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5315_6
timestamp 1731220329
transform 1 0 2472 0 -1 1480
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5314_6
timestamp 1731220329
transform 1 0 2328 0 -1 1480
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5313_6
timestamp 1731220329
transform 1 0 2312 0 1 1344
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5312_6
timestamp 1731220329
transform 1 0 2192 0 1 1344
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5311_6
timestamp 1731220329
transform 1 0 2088 0 1 1344
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5310_6
timestamp 1731220329
transform 1 0 2448 0 1 1344
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5309_6
timestamp 1731220329
transform 1 0 2592 0 1 1344
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5308_6
timestamp 1731220329
transform 1 0 2528 0 -1 1340
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5307_6
timestamp 1731220329
transform 1 0 2376 0 -1 1340
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5306_6
timestamp 1731220329
transform 1 0 2232 0 -1 1340
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5305_6
timestamp 1731220329
transform 1 0 2096 0 -1 1340
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5304_6
timestamp 1731220329
transform 1 0 2336 0 1 1212
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5303_6
timestamp 1731220329
transform 1 0 2192 0 1 1212
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5302_6
timestamp 1731220329
transform 1 0 2056 0 1 1212
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5301_6
timestamp 1731220329
transform 1 0 1928 0 1 1212
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5300_6
timestamp 1731220329
transform 1 0 2384 0 -1 1212
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5299_6
timestamp 1731220329
transform 1 0 2224 0 -1 1212
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5298_6
timestamp 1731220329
transform 1 0 2072 0 -1 1212
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5297_6
timestamp 1731220329
transform 1 0 1928 0 -1 1212
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5296_6
timestamp 1731220329
transform 1 0 1824 0 -1 1212
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5295_6
timestamp 1731220329
transform 1 0 1856 0 1 1072
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5294_6
timestamp 1731220329
transform 1 0 1976 0 1 1072
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5293_6
timestamp 1731220329
transform 1 0 2104 0 1 1072
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5292_6
timestamp 1731220329
transform 1 0 2240 0 1 1072
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5291_6
timestamp 1731220329
transform 1 0 2376 0 1 1072
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5290_6
timestamp 1731220329
transform 1 0 2272 0 -1 1064
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5289_6
timestamp 1731220329
transform 1 0 2184 0 -1 1064
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5288_6
timestamp 1731220329
transform 1 0 2096 0 -1 1064
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5287_6
timestamp 1731220329
transform 1 0 2360 0 -1 1064
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5286_6
timestamp 1731220329
transform 1 0 2448 0 -1 1064
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5285_6
timestamp 1731220329
transform 1 0 2504 0 1 936
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5284_6
timestamp 1731220329
transform 1 0 2400 0 1 936
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5283_6
timestamp 1731220329
transform 1 0 2304 0 1 936
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5282_6
timestamp 1731220329
transform 1 0 2144 0 -1 924
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5281_6
timestamp 1731220329
transform 1 0 1976 0 -1 924
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5280_6
timestamp 1731220329
transform 1 0 2080 0 1 792
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5279_6
timestamp 1731220329
transform 1 0 2320 0 1 792
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5278_6
timestamp 1731220329
transform 1 0 2200 0 1 792
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5277_6
timestamp 1731220329
transform 1 0 2144 0 -1 788
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5276_6
timestamp 1731220329
transform 1 0 2280 0 -1 788
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5275_6
timestamp 1731220329
transform 1 0 2416 0 -1 788
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5274_6
timestamp 1731220329
transform 1 0 2408 0 1 656
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5273_6
timestamp 1731220329
transform 1 0 2256 0 1 656
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5272_6
timestamp 1731220329
transform 1 0 2096 0 1 656
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5271_6
timestamp 1731220329
transform 1 0 2232 0 -1 656
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5270_6
timestamp 1731220329
transform 1 0 1968 0 -1 656
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5269_6
timestamp 1731220329
transform 1 0 1888 0 1 520
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5268_6
timestamp 1731220329
transform 1 0 2008 0 1 520
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5267_6
timestamp 1731220329
transform 1 0 2136 0 1 520
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5266_6
timestamp 1731220329
transform 1 0 2272 0 1 520
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5265_6
timestamp 1731220329
transform 1 0 2416 0 1 520
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5264_6
timestamp 1731220329
transform 1 0 2352 0 -1 516
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5263_6
timestamp 1731220329
transform 1 0 2232 0 -1 516
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5262_6
timestamp 1731220329
transform 1 0 2128 0 -1 516
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5261_6
timestamp 1731220329
transform 1 0 2480 0 -1 516
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5260_6
timestamp 1731220329
transform 1 0 2608 0 -1 516
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5259_6
timestamp 1731220329
transform 1 0 2672 0 1 380
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5258_6
timestamp 1731220329
transform 1 0 2552 0 1 380
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5257_6
timestamp 1731220329
transform 1 0 2440 0 1 380
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5256_6
timestamp 1731220329
transform 1 0 2328 0 1 380
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5255_6
timestamp 1731220329
transform 1 0 2232 0 1 380
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5254_6
timestamp 1731220329
transform 1 0 2472 0 -1 376
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5253_6
timestamp 1731220329
transform 1 0 2352 0 -1 376
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5252_6
timestamp 1731220329
transform 1 0 2240 0 -1 376
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5251_6
timestamp 1731220329
transform 1 0 2144 0 -1 376
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5250_6
timestamp 1731220329
transform 1 0 2056 0 -1 376
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5249_6
timestamp 1731220329
transform 1 0 2440 0 1 244
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5248_6
timestamp 1731220329
transform 1 0 2296 0 1 244
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5247_6
timestamp 1731220329
transform 1 0 2160 0 1 244
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5246_6
timestamp 1731220329
transform 1 0 2032 0 1 244
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5245_6
timestamp 1731220329
transform 1 0 1920 0 1 244
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5244_6
timestamp 1731220329
transform 1 0 2344 0 -1 240
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5243_6
timestamp 1731220329
transform 1 0 2192 0 -1 240
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5242_6
timestamp 1731220329
transform 1 0 2048 0 -1 240
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5241_6
timestamp 1731220329
transform 1 0 1920 0 -1 240
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5240_6
timestamp 1731220329
transform 1 0 1824 0 -1 240
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5239_6
timestamp 1731220329
transform 1 0 2272 0 1 92
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5238_6
timestamp 1731220329
transform 1 0 2152 0 1 92
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5237_6
timestamp 1731220329
transform 1 0 2032 0 1 92
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5236_6
timestamp 1731220329
transform 1 0 1912 0 1 92
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5235_6
timestamp 1731220329
transform 1 0 1824 0 1 92
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5234_6
timestamp 1731220329
transform 1 0 1664 0 1 76
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5233_6
timestamp 1731220329
transform 1 0 1576 0 1 76
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5232_6
timestamp 1731220329
transform 1 0 1488 0 1 76
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5231_6
timestamp 1731220329
transform 1 0 1400 0 1 76
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5230_6
timestamp 1731220329
transform 1 0 1304 0 1 76
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5229_6
timestamp 1731220329
transform 1 0 1208 0 1 76
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5228_6
timestamp 1731220329
transform 1 0 1112 0 1 76
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5227_6
timestamp 1731220329
transform 1 0 1024 0 1 76
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5226_6
timestamp 1731220329
transform 1 0 936 0 1 76
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5225_6
timestamp 1731220329
transform 1 0 840 0 1 76
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5224_6
timestamp 1731220329
transform 1 0 1424 0 -1 228
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5223_6
timestamp 1731220329
transform 1 0 1272 0 -1 228
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5222_6
timestamp 1731220329
transform 1 0 1128 0 -1 228
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5221_6
timestamp 1731220329
transform 1 0 984 0 -1 228
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5220_6
timestamp 1731220329
transform 1 0 832 0 -1 228
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5219_6
timestamp 1731220329
transform 1 0 1144 0 1 232
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5218_6
timestamp 1731220329
transform 1 0 1040 0 1 232
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5217_6
timestamp 1731220329
transform 1 0 936 0 1 232
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5216_6
timestamp 1731220329
transform 1 0 840 0 1 232
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5215_6
timestamp 1731220329
transform 1 0 744 0 1 232
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5214_6
timestamp 1731220329
transform 1 0 904 0 -1 364
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5213_6
timestamp 1731220329
transform 1 0 992 0 -1 364
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5212_6
timestamp 1731220329
transform 1 0 1080 0 -1 364
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5211_6
timestamp 1731220329
transform 1 0 1256 0 -1 364
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5210_6
timestamp 1731220329
transform 1 0 1168 0 -1 364
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5209_6
timestamp 1731220329
transform 1 0 1120 0 1 368
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5208_6
timestamp 1731220329
transform 1 0 1016 0 1 368
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5207_6
timestamp 1731220329
transform 1 0 1224 0 1 368
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5206_6
timestamp 1731220329
transform 1 0 1432 0 1 368
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5205_6
timestamp 1731220329
transform 1 0 1328 0 1 368
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5204_6
timestamp 1731220329
transform 1 0 1216 0 -1 500
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5203_6
timestamp 1731220329
transform 1 0 1056 0 -1 500
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5202_6
timestamp 1731220329
transform 1 0 1368 0 -1 500
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5201_6
timestamp 1731220329
transform 1 0 1520 0 -1 500
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5200_6
timestamp 1731220329
transform 1 0 1664 0 -1 500
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5199_6
timestamp 1731220329
transform 1 0 1664 0 1 504
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5198_6
timestamp 1731220329
transform 1 0 1496 0 1 504
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5197_6
timestamp 1731220329
transform 1 0 1312 0 1 504
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5196_6
timestamp 1731220329
transform 1 0 1520 0 -1 636
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5195_6
timestamp 1731220329
transform 1 0 1664 0 -1 636
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5194_6
timestamp 1731220329
transform 1 0 1664 0 1 640
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5193_6
timestamp 1731220329
transform 1 0 1824 0 1 656
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5192_6
timestamp 1731220329
transform 1 0 1944 0 1 656
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5191_6
timestamp 1731220329
transform 1 0 1872 0 -1 788
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5190_6
timestamp 1731220329
transform 1 0 2008 0 -1 788
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5189_6
timestamp 1731220329
transform 1 0 1952 0 1 792
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5188_6
timestamp 1731220329
transform 1 0 1824 0 1 792
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5187_6
timestamp 1731220329
transform 1 0 1824 0 -1 924
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5186_6
timestamp 1731220329
transform 1 0 1664 0 1 916
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5185_6
timestamp 1731220329
transform 1 0 1576 0 1 916
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5184_6
timestamp 1731220329
transform 1 0 1480 0 1 916
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5183_6
timestamp 1731220329
transform 1 0 1664 0 -1 1048
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5182_6
timestamp 1731220329
transform 1 0 1528 0 -1 1048
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5181_6
timestamp 1731220329
transform 1 0 1376 0 -1 1048
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5180_6
timestamp 1731220329
transform 1 0 1384 0 1 916
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5179_6
timestamp 1731220329
transform 1 0 1288 0 1 916
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5178_6
timestamp 1731220329
transform 1 0 1192 0 1 916
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5177_6
timestamp 1731220329
transform 1 0 1088 0 1 916
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5176_6
timestamp 1731220329
transform 1 0 1336 0 -1 912
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5175_6
timestamp 1731220329
transform 1 0 1456 0 -1 912
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5174_6
timestamp 1731220329
transform 1 0 1576 0 -1 912
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5173_6
timestamp 1731220329
transform 1 0 1552 0 1 780
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5172_6
timestamp 1731220329
transform 1 0 1424 0 1 780
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5171_6
timestamp 1731220329
transform 1 0 1304 0 1 780
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5170_6
timestamp 1731220329
transform 1 0 1184 0 1 780
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5169_6
timestamp 1731220329
transform 1 0 1152 0 -1 776
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5168_6
timestamp 1731220329
transform 1 0 1280 0 -1 776
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5167_6
timestamp 1731220329
transform 1 0 1408 0 -1 776
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5166_6
timestamp 1731220329
transform 1 0 1504 0 1 640
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5165_6
timestamp 1731220329
transform 1 0 1320 0 1 640
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5164_6
timestamp 1731220329
transform 1 0 1144 0 1 640
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5163_6
timestamp 1731220329
transform 1 0 1360 0 -1 636
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5162_6
timestamp 1731220329
transform 1 0 1200 0 -1 636
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5161_6
timestamp 1731220329
transform 1 0 1048 0 -1 636
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5160_6
timestamp 1731220329
transform 1 0 1128 0 1 504
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5159_6
timestamp 1731220329
transform 1 0 944 0 1 504
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5158_6
timestamp 1731220329
transform 1 0 904 0 -1 636
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5157_6
timestamp 1731220329
transform 1 0 760 0 -1 636
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5156_6
timestamp 1731220329
transform 1 0 824 0 1 640
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5155_6
timestamp 1731220329
transform 1 0 976 0 1 640
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5154_6
timestamp 1731220329
transform 1 0 904 0 -1 776
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5153_6
timestamp 1731220329
transform 1 0 1024 0 -1 776
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5152_6
timestamp 1731220329
transform 1 0 1064 0 1 780
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5151_6
timestamp 1731220329
transform 1 0 1216 0 -1 912
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5150_6
timestamp 1731220329
transform 1 0 1104 0 -1 912
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5149_6
timestamp 1731220329
transform 1 0 984 0 1 916
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5148_6
timestamp 1731220329
transform 1 0 1072 0 -1 1048
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5147_6
timestamp 1731220329
transform 1 0 1224 0 -1 1048
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5146_6
timestamp 1731220329
transform 1 0 1552 0 1 1056
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5145_6
timestamp 1731220329
transform 1 0 1400 0 1 1056
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5144_6
timestamp 1731220329
transform 1 0 1256 0 1 1056
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5143_6
timestamp 1731220329
transform 1 0 1112 0 1 1056
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5142_6
timestamp 1731220329
transform 1 0 960 0 1 1056
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5141_6
timestamp 1731220329
transform 1 0 1328 0 -1 1188
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5140_6
timestamp 1731220329
transform 1 0 1192 0 -1 1188
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5139_6
timestamp 1731220329
transform 1 0 1056 0 -1 1188
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5138_6
timestamp 1731220329
transform 1 0 920 0 -1 1188
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5137_6
timestamp 1731220329
transform 1 0 784 0 -1 1188
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5136_6
timestamp 1731220329
transform 1 0 1184 0 1 1192
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5135_6
timestamp 1731220329
transform 1 0 1064 0 1 1192
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5134_6
timestamp 1731220329
transform 1 0 952 0 1 1192
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5133_6
timestamp 1731220329
transform 1 0 840 0 1 1192
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5132_6
timestamp 1731220329
transform 1 0 728 0 1 1192
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5131_6
timestamp 1731220329
transform 1 0 1072 0 -1 1324
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5130_6
timestamp 1731220329
transform 1 0 960 0 -1 1324
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5129_6
timestamp 1731220329
transform 1 0 840 0 -1 1324
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5128_6
timestamp 1731220329
transform 1 0 712 0 -1 1324
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5127_6
timestamp 1731220329
transform 1 0 608 0 1 1192
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5126_6
timestamp 1731220329
transform 1 0 576 0 -1 1324
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5125_6
timestamp 1731220329
transform 1 0 432 0 -1 1324
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5124_6
timestamp 1731220329
transform 1 0 272 0 -1 1324
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5123_6
timestamp 1731220329
transform 1 0 600 0 1 1328
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5122_6
timestamp 1731220329
transform 1 0 752 0 1 1328
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5121_6
timestamp 1731220329
transform 1 0 776 0 -1 1460
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5120_6
timestamp 1731220329
transform 1 0 624 0 -1 1460
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5119_6
timestamp 1731220329
transform 1 0 464 0 -1 1460
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5118_6
timestamp 1731220329
transform 1 0 600 0 1 1468
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5117_6
timestamp 1731220329
transform 1 0 744 0 1 1468
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5116_6
timestamp 1731220329
transform 1 0 808 0 -1 1600
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5115_6
timestamp 1731220329
transform 1 0 664 0 -1 1600
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5114_6
timestamp 1731220329
transform 1 0 536 0 -1 1600
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5113_6
timestamp 1731220329
transform 1 0 528 0 1 1604
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5112_6
timestamp 1731220329
transform 1 0 680 0 1 1604
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5111_6
timestamp 1731220329
transform 1 0 560 0 -1 1736
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5110_6
timestamp 1731220329
transform 1 0 744 0 -1 1736
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5109_6
timestamp 1731220329
transform 1 0 792 0 1 1748
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5108_6
timestamp 1731220329
transform 1 0 648 0 1 1748
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5107_6
timestamp 1731220329
transform 1 0 520 0 1 1748
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5106_6
timestamp 1731220329
transform 1 0 400 0 1 1748
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5105_6
timestamp 1731220329
transform 1 0 304 0 1 1748
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5104_6
timestamp 1731220329
transform 1 0 216 0 1 1748
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5103_6
timestamp 1731220329
transform 1 0 128 0 1 1748
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5102_6
timestamp 1731220329
transform 1 0 128 0 -1 1736
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5101_6
timestamp 1731220329
transform 1 0 240 0 -1 1736
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5100_6
timestamp 1731220329
transform 1 0 392 0 -1 1736
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_599_6
timestamp 1731220329
transform 1 0 400 0 1 1604
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_598_6
timestamp 1731220329
transform 1 0 288 0 1 1604
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_597_6
timestamp 1731220329
transform 1 0 184 0 1 1604
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_596_6
timestamp 1731220329
transform 1 0 320 0 -1 1600
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_595_6
timestamp 1731220329
transform 1 0 424 0 -1 1600
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_594_6
timestamp 1731220329
transform 1 0 464 0 1 1468
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_593_6
timestamp 1731220329
transform 1 0 336 0 1 1468
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_592_6
timestamp 1731220329
transform 1 0 216 0 1 1468
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_591_6
timestamp 1731220329
transform 1 0 128 0 -1 1460
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_590_6
timestamp 1731220329
transform 1 0 296 0 -1 1460
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_589_6
timestamp 1731220329
transform 1 0 440 0 1 1328
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_588_6
timestamp 1731220329
transform 1 0 272 0 1 1328
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_587_6
timestamp 1731220329
transform 1 0 128 0 1 1328
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_586_6
timestamp 1731220329
transform 1 0 128 0 -1 1324
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_585_6
timestamp 1731220329
transform 1 0 128 0 1 1192
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_584_6
timestamp 1731220329
transform 1 0 232 0 1 1192
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_583_6
timestamp 1731220329
transform 1 0 360 0 1 1192
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_582_6
timestamp 1731220329
transform 1 0 488 0 1 1192
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_581_6
timestamp 1731220329
transform 1 0 648 0 -1 1188
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_580_6
timestamp 1731220329
transform 1 0 504 0 -1 1188
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_579_6
timestamp 1731220329
transform 1 0 368 0 -1 1188
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_578_6
timestamp 1731220329
transform 1 0 232 0 -1 1188
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_577_6
timestamp 1731220329
transform 1 0 128 0 -1 1188
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_576_6
timestamp 1731220329
transform 1 0 184 0 1 1056
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_575_6
timestamp 1731220329
transform 1 0 328 0 1 1056
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_574_6
timestamp 1731220329
transform 1 0 488 0 1 1056
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_573_6
timestamp 1731220329
transform 1 0 808 0 1 1056
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_572_6
timestamp 1731220329
transform 1 0 648 0 1 1056
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_571_6
timestamp 1731220329
transform 1 0 600 0 -1 1048
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_570_6
timestamp 1731220329
transform 1 0 456 0 -1 1048
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_569_6
timestamp 1731220329
transform 1 0 320 0 -1 1048
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_568_6
timestamp 1731220329
transform 1 0 760 0 -1 1048
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_567_6
timestamp 1731220329
transform 1 0 920 0 -1 1048
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_566_6
timestamp 1731220329
transform 1 0 880 0 1 916
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_565_6
timestamp 1731220329
transform 1 0 776 0 1 916
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_564_6
timestamp 1731220329
transform 1 0 664 0 1 916
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_563_6
timestamp 1731220329
transform 1 0 560 0 1 916
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_562_6
timestamp 1731220329
transform 1 0 464 0 1 916
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_561_6
timestamp 1731220329
transform 1 0 600 0 -1 912
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_560_6
timestamp 1731220329
transform 1 0 688 0 -1 912
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_559_6
timestamp 1731220329
transform 1 0 784 0 -1 912
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_558_6
timestamp 1731220329
transform 1 0 888 0 -1 912
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_557_6
timestamp 1731220329
transform 1 0 992 0 -1 912
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_556_6
timestamp 1731220329
transform 1 0 944 0 1 780
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_555_6
timestamp 1731220329
transform 1 0 824 0 1 780
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_554_6
timestamp 1731220329
transform 1 0 712 0 1 780
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_553_6
timestamp 1731220329
transform 1 0 608 0 1 780
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_552_6
timestamp 1731220329
transform 1 0 512 0 1 780
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_551_6
timestamp 1731220329
transform 1 0 784 0 -1 776
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_550_6
timestamp 1731220329
transform 1 0 672 0 -1 776
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_549_6
timestamp 1731220329
transform 1 0 568 0 -1 776
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_548_6
timestamp 1731220329
transform 1 0 464 0 -1 776
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_547_6
timestamp 1731220329
transform 1 0 376 0 -1 776
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_546_6
timestamp 1731220329
transform 1 0 688 0 1 640
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_545_6
timestamp 1731220329
transform 1 0 560 0 1 640
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_544_6
timestamp 1731220329
transform 1 0 448 0 1 640
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_543_6
timestamp 1731220329
transform 1 0 336 0 1 640
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_542_6
timestamp 1731220329
transform 1 0 240 0 1 640
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_541_6
timestamp 1731220329
transform 1 0 616 0 -1 636
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_540_6
timestamp 1731220329
transform 1 0 480 0 -1 636
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_539_6
timestamp 1731220329
transform 1 0 352 0 -1 636
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_538_6
timestamp 1731220329
transform 1 0 224 0 -1 636
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_537_6
timestamp 1731220329
transform 1 0 128 0 -1 636
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_536_6
timestamp 1731220329
transform 1 0 128 0 1 504
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_535_6
timestamp 1731220329
transform 1 0 240 0 1 504
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_534_6
timestamp 1731220329
transform 1 0 400 0 1 504
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_533_6
timestamp 1731220329
transform 1 0 760 0 1 504
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_532_6
timestamp 1731220329
transform 1 0 576 0 1 504
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_531_6
timestamp 1731220329
transform 1 0 560 0 -1 500
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_530_6
timestamp 1731220329
transform 1 0 392 0 -1 500
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_529_6
timestamp 1731220329
transform 1 0 240 0 -1 500
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_528_6
timestamp 1731220329
transform 1 0 728 0 -1 500
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_527_6
timestamp 1731220329
transform 1 0 896 0 -1 500
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_526_6
timestamp 1731220329
transform 1 0 920 0 1 368
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_525_6
timestamp 1731220329
transform 1 0 712 0 1 368
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_524_6
timestamp 1731220329
transform 1 0 608 0 1 368
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_523_6
timestamp 1731220329
transform 1 0 512 0 1 368
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_522_6
timestamp 1731220329
transform 1 0 816 0 1 368
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_521_6
timestamp 1731220329
transform 1 0 816 0 -1 364
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_520_6
timestamp 1731220329
transform 1 0 728 0 -1 364
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_519_6
timestamp 1731220329
transform 1 0 640 0 -1 364
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_518_6
timestamp 1731220329
transform 1 0 552 0 -1 364
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_517_6
timestamp 1731220329
transform 1 0 464 0 -1 364
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_516_6
timestamp 1731220329
transform 1 0 648 0 1 232
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_515_6
timestamp 1731220329
transform 1 0 552 0 1 232
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_514_6
timestamp 1731220329
transform 1 0 456 0 1 232
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_513_6
timestamp 1731220329
transform 1 0 360 0 1 232
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_512_6
timestamp 1731220329
transform 1 0 272 0 1 232
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_511_6
timestamp 1731220329
transform 1 0 672 0 -1 228
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_510_6
timestamp 1731220329
transform 1 0 504 0 -1 228
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_59_6
timestamp 1731220329
transform 1 0 336 0 -1 228
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_58_6
timestamp 1731220329
transform 1 0 160 0 -1 228
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_57_6
timestamp 1731220329
transform 1 0 744 0 1 76
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_56_6
timestamp 1731220329
transform 1 0 656 0 1 76
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_55_6
timestamp 1731220329
transform 1 0 568 0 1 76
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_54_6
timestamp 1731220329
transform 1 0 480 0 1 76
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_53_6
timestamp 1731220329
transform 1 0 392 0 1 76
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_52_6
timestamp 1731220329
transform 1 0 304 0 1 76
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_51_6
timestamp 1731220329
transform 1 0 216 0 1 76
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_50_6
timestamp 1731220329
transform 1 0 128 0 1 76
box 8 4 84 60
<< end >>
