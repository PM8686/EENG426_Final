magic
tech sky130l
timestamp 1730743719
<< m1 >>
rect 616 635 620 675
rect 344 563 348 583
rect 200 423 204 437
rect 248 343 252 379
rect 552 307 556 321
rect 264 163 268 227
<< m2c >>
rect 288 769 292 773
rect 376 769 380 773
rect 472 769 476 773
rect 568 769 572 773
rect 648 769 652 773
rect 111 753 115 757
rect 295 752 299 756
rect 304 751 308 755
rect 383 752 387 756
rect 392 751 396 755
rect 479 752 483 756
rect 488 751 492 755
rect 575 752 579 756
rect 655 752 659 756
rect 687 753 691 757
rect 111 735 115 739
rect 687 735 691 739
rect 584 731 588 735
rect 111 709 115 713
rect 344 711 348 715
rect 664 711 668 715
rect 687 709 691 713
rect 111 691 115 695
rect 215 692 219 696
rect 224 691 228 695
rect 255 692 259 696
rect 264 691 268 695
rect 295 692 299 696
rect 304 691 308 695
rect 335 692 339 696
rect 375 692 379 696
rect 384 691 388 695
rect 423 692 427 696
rect 432 691 436 695
rect 479 692 483 696
rect 488 691 492 695
rect 543 692 547 696
rect 552 691 556 695
rect 607 692 611 696
rect 616 691 620 695
rect 655 692 659 696
rect 687 691 691 695
rect 208 675 212 679
rect 248 675 252 679
rect 288 675 292 679
rect 328 675 332 679
rect 368 675 372 679
rect 416 675 420 679
rect 472 675 476 679
rect 536 675 540 679
rect 600 675 604 679
rect 616 675 620 679
rect 648 675 652 679
rect 168 661 172 665
rect 224 661 228 665
rect 288 661 292 665
rect 360 661 364 665
rect 432 661 436 665
rect 512 661 516 665
rect 592 661 596 665
rect 111 645 115 649
rect 175 644 179 648
rect 184 643 188 647
rect 231 644 235 648
rect 240 643 244 647
rect 295 644 299 648
rect 304 643 308 647
rect 367 644 371 648
rect 439 644 443 648
rect 519 644 523 648
rect 599 644 603 648
rect 648 661 652 665
rect 655 644 659 648
rect 687 645 691 649
rect 608 631 612 635
rect 616 631 620 635
rect 111 627 115 631
rect 687 627 691 631
rect 376 623 380 627
rect 448 623 452 627
rect 528 623 532 627
rect 664 623 668 627
rect 111 593 115 597
rect 224 595 228 599
rect 320 595 324 599
rect 664 595 668 599
rect 687 593 691 597
rect 264 583 268 587
rect 344 583 348 587
rect 376 583 380 587
rect 440 583 444 587
rect 111 575 115 579
rect 215 576 219 580
rect 255 576 259 580
rect 311 576 315 580
rect 367 576 371 580
rect 431 576 435 580
rect 503 576 507 580
rect 512 575 516 579
rect 583 576 587 580
rect 592 575 596 579
rect 655 576 659 580
rect 687 575 691 579
rect 208 559 212 563
rect 248 559 252 563
rect 304 559 308 563
rect 344 559 348 563
rect 360 559 364 563
rect 424 559 428 563
rect 496 559 500 563
rect 576 559 580 563
rect 648 559 652 563
rect 320 545 324 549
rect 360 545 364 549
rect 400 545 404 549
rect 448 545 452 549
rect 496 545 500 549
rect 552 545 556 549
rect 608 545 612 549
rect 648 545 652 549
rect 111 529 115 533
rect 327 528 331 532
rect 336 527 340 531
rect 367 528 371 532
rect 376 527 380 531
rect 407 528 411 532
rect 416 527 420 531
rect 455 528 459 532
rect 503 528 507 532
rect 512 527 516 531
rect 559 528 563 532
rect 615 528 619 532
rect 624 527 628 531
rect 655 528 659 532
rect 687 529 691 533
rect 111 511 115 515
rect 687 511 691 515
rect 464 507 468 511
rect 568 507 572 511
rect 664 507 668 511
rect 111 485 115 489
rect 536 487 540 491
rect 664 487 668 491
rect 687 485 691 489
rect 111 467 115 471
rect 271 468 275 472
rect 280 467 284 471
rect 311 468 315 472
rect 320 467 324 471
rect 351 468 355 472
rect 360 467 364 471
rect 407 468 411 472
rect 416 467 420 471
rect 463 468 467 472
rect 472 467 476 471
rect 527 468 531 472
rect 599 468 603 472
rect 608 467 612 471
rect 655 468 659 472
rect 687 467 691 471
rect 264 451 268 455
rect 304 451 308 455
rect 344 451 348 455
rect 400 451 404 455
rect 456 451 460 455
rect 520 451 524 455
rect 592 451 596 455
rect 648 451 652 455
rect 168 437 172 441
rect 200 437 204 441
rect 216 437 220 441
rect 272 437 276 441
rect 336 437 340 441
rect 408 437 412 441
rect 488 437 492 441
rect 576 437 580 441
rect 648 437 652 441
rect 111 421 115 425
rect 175 420 179 424
rect 184 419 188 423
rect 200 419 204 423
rect 223 420 227 424
rect 232 419 236 423
rect 279 420 283 424
rect 288 419 292 423
rect 343 420 347 424
rect 352 419 356 423
rect 415 420 419 424
rect 424 419 428 423
rect 495 420 499 424
rect 504 419 508 423
rect 583 420 587 424
rect 655 420 659 424
rect 664 419 668 423
rect 687 421 691 425
rect 111 403 115 407
rect 687 403 691 407
rect 592 399 596 403
rect 248 379 252 383
rect 111 373 115 377
rect 200 375 204 379
rect 240 363 244 367
rect 111 355 115 359
rect 151 356 155 360
rect 160 355 164 359
rect 191 356 195 360
rect 231 356 235 360
rect 304 375 308 379
rect 664 375 668 379
rect 687 373 691 377
rect 440 363 444 367
rect 295 356 299 360
rect 359 356 363 360
rect 368 355 372 359
rect 431 356 435 360
rect 511 356 515 360
rect 520 355 524 359
rect 591 356 595 360
rect 600 355 604 359
rect 655 356 659 360
rect 687 355 691 359
rect 144 339 148 343
rect 184 339 188 343
rect 224 339 228 343
rect 248 339 252 343
rect 288 339 292 343
rect 352 339 356 343
rect 424 339 428 343
rect 504 339 508 343
rect 584 339 588 343
rect 648 339 652 343
rect 248 321 252 325
rect 288 321 292 325
rect 328 321 332 325
rect 376 321 380 325
rect 424 321 428 325
rect 472 321 476 325
rect 520 321 524 325
rect 552 321 556 325
rect 568 321 572 325
rect 608 321 612 325
rect 648 321 652 325
rect 111 305 115 309
rect 255 304 259 308
rect 264 303 268 307
rect 295 304 299 308
rect 304 303 308 307
rect 335 304 339 308
rect 344 303 348 307
rect 383 304 387 308
rect 431 304 435 308
rect 440 303 444 307
rect 479 304 483 308
rect 488 303 492 307
rect 527 304 531 308
rect 536 303 540 307
rect 552 303 556 307
rect 575 304 579 308
rect 615 304 619 308
rect 655 304 659 308
rect 687 305 691 309
rect 111 287 115 291
rect 687 287 691 291
rect 392 283 396 287
rect 584 283 588 287
rect 624 283 628 287
rect 664 283 668 287
rect 111 261 115 265
rect 664 263 668 267
rect 464 259 468 263
rect 687 261 691 265
rect 111 243 115 247
rect 255 244 259 248
rect 264 243 268 247
rect 295 244 299 248
rect 304 243 308 247
rect 335 244 339 248
rect 344 243 348 247
rect 375 244 379 248
rect 384 243 388 247
rect 415 244 419 248
rect 424 243 428 247
rect 455 244 459 248
rect 495 244 499 248
rect 504 243 508 247
rect 535 244 539 248
rect 544 243 548 247
rect 575 244 579 248
rect 584 243 588 247
rect 615 244 619 248
rect 624 243 628 247
rect 655 244 659 248
rect 687 243 691 247
rect 248 227 252 231
rect 264 227 268 231
rect 288 227 292 231
rect 328 227 332 231
rect 368 227 372 231
rect 408 227 412 231
rect 448 227 452 231
rect 488 227 492 231
rect 528 227 532 231
rect 568 227 572 231
rect 608 227 612 231
rect 648 227 652 231
rect 200 201 204 205
rect 240 201 244 205
rect 111 185 115 189
rect 207 184 211 188
rect 216 183 220 187
rect 247 184 251 188
rect 111 167 115 171
rect 256 167 260 171
rect 280 201 284 205
rect 320 201 324 205
rect 360 201 364 205
rect 400 201 404 205
rect 287 184 291 188
rect 296 183 300 187
rect 327 184 331 188
rect 336 183 340 187
rect 367 184 371 188
rect 376 183 380 187
rect 407 184 411 188
rect 687 185 691 189
rect 687 167 691 171
rect 416 163 420 167
rect 264 159 268 163
rect 111 125 115 129
rect 480 127 484 131
rect 687 125 691 129
rect 111 107 115 111
rect 151 108 155 112
rect 160 107 164 111
rect 191 108 195 112
rect 200 107 204 111
rect 231 108 235 112
rect 240 107 244 111
rect 271 108 275 112
rect 280 107 284 111
rect 311 108 315 112
rect 320 107 324 111
rect 351 108 355 112
rect 360 107 364 111
rect 391 108 395 112
rect 400 107 404 111
rect 431 108 435 112
rect 440 107 444 111
rect 471 108 475 112
rect 687 107 691 111
rect 184 91 188 95
rect 224 91 228 95
rect 264 91 268 95
rect 304 91 308 95
rect 344 91 348 95
rect 384 91 388 95
rect 424 91 428 95
rect 464 91 468 95
<< m2 >>
rect 287 773 293 774
rect 287 769 288 773
rect 292 772 293 773
rect 374 773 381 774
rect 292 770 306 772
rect 342 771 348 772
rect 342 770 343 771
rect 292 769 293 770
rect 287 768 293 769
rect 304 768 343 770
rect 342 767 343 768
rect 347 767 348 771
rect 374 769 375 773
rect 380 769 381 773
rect 374 768 381 769
rect 454 773 460 774
rect 454 769 455 773
rect 459 772 460 773
rect 471 773 477 774
rect 471 772 472 773
rect 459 770 472 772
rect 459 769 460 770
rect 454 768 460 769
rect 471 769 472 770
rect 476 769 477 773
rect 471 768 477 769
rect 550 773 556 774
rect 550 769 551 773
rect 555 772 556 773
rect 567 773 573 774
rect 567 772 568 773
rect 555 770 568 772
rect 555 769 556 770
rect 550 768 556 769
rect 567 769 568 770
rect 572 769 573 773
rect 567 768 573 769
rect 647 773 653 774
rect 647 769 648 773
rect 652 772 653 773
rect 662 773 668 774
rect 662 772 663 773
rect 652 770 663 772
rect 652 769 653 770
rect 647 768 653 769
rect 662 769 663 770
rect 667 769 668 773
rect 662 768 668 769
rect 342 766 348 767
rect 110 757 116 758
rect 686 757 692 758
rect 110 753 111 757
rect 115 753 116 757
rect 110 752 116 753
rect 294 756 300 757
rect 382 756 388 757
rect 478 756 484 757
rect 574 756 580 757
rect 294 752 295 756
rect 299 752 300 756
rect 294 751 300 752
rect 303 755 309 756
rect 303 751 304 755
rect 308 754 309 755
rect 374 755 380 756
rect 374 754 375 755
rect 308 752 375 754
rect 308 751 309 752
rect 303 750 309 751
rect 374 751 375 752
rect 379 751 380 755
rect 382 752 383 756
rect 387 752 388 756
rect 382 751 388 752
rect 391 755 397 756
rect 391 751 392 755
rect 396 754 397 755
rect 454 755 460 756
rect 454 754 455 755
rect 396 752 455 754
rect 396 751 397 752
rect 374 750 380 751
rect 391 750 397 751
rect 454 751 455 752
rect 459 751 460 755
rect 478 752 479 756
rect 483 752 484 756
rect 478 751 484 752
rect 487 755 493 756
rect 487 751 488 755
rect 492 754 493 755
rect 550 755 556 756
rect 550 754 551 755
rect 492 752 551 754
rect 492 751 493 752
rect 454 750 460 751
rect 487 750 493 751
rect 550 751 551 752
rect 555 751 556 755
rect 574 752 575 756
rect 579 752 580 756
rect 574 751 580 752
rect 654 756 660 757
rect 654 752 655 756
rect 659 752 660 756
rect 686 753 687 757
rect 691 753 692 757
rect 686 752 692 753
rect 654 751 660 752
rect 550 750 556 751
rect 278 741 284 742
rect 110 739 116 740
rect 110 735 111 739
rect 115 735 116 739
rect 278 737 279 741
rect 283 737 284 741
rect 278 736 284 737
rect 366 741 372 742
rect 366 737 367 741
rect 371 737 372 741
rect 366 736 372 737
rect 462 741 468 742
rect 462 737 463 741
rect 467 737 468 741
rect 462 736 468 737
rect 558 741 564 742
rect 558 737 559 741
rect 563 737 564 741
rect 558 736 564 737
rect 638 741 644 742
rect 638 737 639 741
rect 643 737 644 741
rect 638 736 644 737
rect 686 739 692 740
rect 110 734 116 735
rect 390 735 396 736
rect 390 731 391 735
rect 395 734 396 735
rect 583 735 589 736
rect 583 734 584 735
rect 395 732 584 734
rect 395 731 396 732
rect 390 730 396 731
rect 583 731 584 732
rect 588 731 589 735
rect 686 735 687 739
rect 691 735 692 739
rect 686 734 692 735
rect 583 730 589 731
rect 342 715 349 716
rect 110 713 116 714
rect 110 709 111 713
rect 115 709 116 713
rect 110 708 116 709
rect 198 711 204 712
rect 198 707 199 711
rect 203 707 204 711
rect 198 706 204 707
rect 238 711 244 712
rect 238 707 239 711
rect 243 707 244 711
rect 238 706 244 707
rect 278 711 284 712
rect 278 707 279 711
rect 283 707 284 711
rect 278 706 284 707
rect 318 711 324 712
rect 318 707 319 711
rect 323 707 324 711
rect 342 711 343 715
rect 348 711 349 715
rect 662 715 669 716
rect 342 710 349 711
rect 358 711 364 712
rect 318 706 324 707
rect 358 707 359 711
rect 363 707 364 711
rect 358 706 364 707
rect 406 711 412 712
rect 406 707 407 711
rect 411 707 412 711
rect 406 706 412 707
rect 462 711 468 712
rect 462 707 463 711
rect 467 707 468 711
rect 462 706 468 707
rect 526 711 532 712
rect 526 707 527 711
rect 531 707 532 711
rect 526 706 532 707
rect 590 711 596 712
rect 590 707 591 711
rect 595 707 596 711
rect 590 706 596 707
rect 638 711 644 712
rect 638 707 639 711
rect 643 707 644 711
rect 662 711 663 715
rect 668 711 669 715
rect 662 710 669 711
rect 686 713 692 714
rect 686 709 687 713
rect 691 709 692 713
rect 686 708 692 709
rect 638 706 644 707
rect 214 696 220 697
rect 254 696 260 697
rect 294 696 300 697
rect 334 696 340 697
rect 110 695 116 696
rect 110 691 111 695
rect 115 691 116 695
rect 214 692 215 696
rect 219 692 220 696
rect 214 691 220 692
rect 223 695 229 696
rect 223 691 224 695
rect 228 694 229 695
rect 228 692 238 694
rect 228 691 229 692
rect 110 690 116 691
rect 223 690 229 691
rect 207 679 213 680
rect 207 675 208 679
rect 212 678 213 679
rect 222 679 228 680
rect 222 678 223 679
rect 212 676 223 678
rect 212 675 213 676
rect 207 674 213 675
rect 222 675 223 676
rect 227 675 228 679
rect 236 678 238 692
rect 254 692 255 696
rect 259 692 260 696
rect 254 691 260 692
rect 263 695 269 696
rect 263 691 264 695
rect 268 694 269 695
rect 268 692 278 694
rect 268 691 269 692
rect 263 690 269 691
rect 247 679 253 680
rect 247 678 248 679
rect 236 676 248 678
rect 222 674 228 675
rect 247 675 248 676
rect 252 675 253 679
rect 276 678 278 692
rect 294 692 295 696
rect 299 692 300 696
rect 294 691 300 692
rect 303 695 309 696
rect 303 691 304 695
rect 308 694 309 695
rect 308 692 314 694
rect 308 691 309 692
rect 303 690 309 691
rect 287 679 293 680
rect 287 678 288 679
rect 276 676 288 678
rect 247 674 253 675
rect 287 675 288 676
rect 292 675 293 679
rect 312 678 314 692
rect 334 692 335 696
rect 339 692 340 696
rect 334 691 340 692
rect 374 696 380 697
rect 422 696 428 697
rect 478 696 484 697
rect 542 696 548 697
rect 606 696 612 697
rect 654 696 660 697
rect 374 692 375 696
rect 379 692 380 696
rect 374 691 380 692
rect 383 695 389 696
rect 383 691 384 695
rect 388 694 389 695
rect 388 692 402 694
rect 388 691 389 692
rect 383 690 389 691
rect 327 679 333 680
rect 327 678 328 679
rect 312 676 328 678
rect 287 674 293 675
rect 327 675 328 676
rect 332 675 333 679
rect 327 674 333 675
rect 367 679 373 680
rect 367 675 368 679
rect 372 678 373 679
rect 390 679 396 680
rect 390 678 391 679
rect 372 676 391 678
rect 372 675 373 676
rect 367 674 373 675
rect 390 675 391 676
rect 395 675 396 679
rect 400 678 402 692
rect 422 692 423 696
rect 427 692 428 696
rect 422 691 428 692
rect 431 695 437 696
rect 431 691 432 695
rect 436 694 437 695
rect 436 692 454 694
rect 436 691 437 692
rect 431 690 437 691
rect 415 679 421 680
rect 415 678 416 679
rect 400 676 416 678
rect 390 674 396 675
rect 415 675 416 676
rect 420 675 421 679
rect 452 678 454 692
rect 478 692 479 696
rect 483 692 484 696
rect 478 691 484 692
rect 487 695 493 696
rect 487 691 488 695
rect 492 694 493 695
rect 492 692 514 694
rect 492 691 493 692
rect 487 690 493 691
rect 471 679 477 680
rect 471 678 472 679
rect 452 676 472 678
rect 415 674 421 675
rect 471 675 472 676
rect 476 675 477 679
rect 512 678 514 692
rect 542 692 543 696
rect 547 692 548 696
rect 542 691 548 692
rect 550 695 557 696
rect 550 691 551 695
rect 556 691 557 695
rect 606 692 607 696
rect 611 692 612 696
rect 606 691 612 692
rect 615 695 621 696
rect 615 691 616 695
rect 620 694 621 695
rect 620 692 634 694
rect 620 691 621 692
rect 550 690 557 691
rect 615 690 621 691
rect 535 679 541 680
rect 535 678 536 679
rect 512 676 536 678
rect 471 674 477 675
rect 535 675 536 676
rect 540 675 541 679
rect 535 674 541 675
rect 599 679 605 680
rect 599 675 600 679
rect 604 678 605 679
rect 615 679 621 680
rect 615 678 616 679
rect 604 676 616 678
rect 604 675 605 676
rect 599 674 605 675
rect 615 675 616 676
rect 620 675 621 679
rect 632 678 634 692
rect 654 692 655 696
rect 659 692 660 696
rect 654 691 660 692
rect 686 695 692 696
rect 686 691 687 695
rect 691 691 692 695
rect 686 690 692 691
rect 647 679 653 680
rect 647 678 648 679
rect 632 676 648 678
rect 615 674 621 675
rect 647 675 648 676
rect 652 675 653 679
rect 647 674 653 675
rect 502 667 508 668
rect 502 666 503 667
rect 167 665 173 666
rect 167 661 168 665
rect 172 664 173 665
rect 186 665 192 666
rect 186 664 187 665
rect 172 662 187 664
rect 172 661 173 662
rect 167 660 173 661
rect 186 661 187 662
rect 191 661 192 665
rect 186 660 192 661
rect 206 665 212 666
rect 206 661 207 665
rect 211 664 212 665
rect 223 665 229 666
rect 223 664 224 665
rect 211 662 224 664
rect 211 661 212 662
rect 206 660 212 661
rect 223 661 224 662
rect 228 661 229 665
rect 223 660 229 661
rect 270 665 276 666
rect 270 661 271 665
rect 275 664 276 665
rect 287 665 293 666
rect 287 664 288 665
rect 275 662 288 664
rect 275 661 276 662
rect 270 660 276 661
rect 287 661 288 662
rect 292 661 293 665
rect 287 660 293 661
rect 358 665 365 666
rect 358 661 359 665
rect 364 661 365 665
rect 358 660 365 661
rect 431 665 437 666
rect 431 661 432 665
rect 436 664 437 665
rect 456 664 503 666
rect 436 662 458 664
rect 502 663 503 664
rect 507 663 508 667
rect 550 667 556 668
rect 550 666 551 667
rect 502 662 508 663
rect 511 665 517 666
rect 436 661 437 662
rect 431 660 437 661
rect 511 661 512 665
rect 516 664 517 665
rect 532 664 551 666
rect 516 662 534 664
rect 550 663 551 664
rect 555 663 556 667
rect 550 662 556 663
rect 591 665 597 666
rect 516 661 517 662
rect 511 660 517 661
rect 591 661 592 665
rect 596 662 597 665
rect 647 665 653 666
rect 630 663 636 664
rect 630 662 631 663
rect 596 661 631 662
rect 591 660 631 661
rect 630 659 631 660
rect 635 659 636 663
rect 647 661 648 665
rect 652 664 653 665
rect 662 665 668 666
rect 662 664 663 665
rect 652 662 663 664
rect 652 661 653 662
rect 647 660 653 661
rect 662 661 663 662
rect 667 661 668 665
rect 662 660 668 661
rect 630 658 636 659
rect 110 649 116 650
rect 686 649 692 650
rect 110 645 111 649
rect 115 645 116 649
rect 110 644 116 645
rect 174 648 180 649
rect 230 648 236 649
rect 294 648 300 649
rect 366 648 372 649
rect 174 644 175 648
rect 179 644 180 648
rect 174 643 180 644
rect 183 647 189 648
rect 183 643 184 647
rect 188 646 189 647
rect 206 647 212 648
rect 206 646 207 647
rect 188 644 207 646
rect 188 643 189 644
rect 183 642 189 643
rect 206 643 207 644
rect 211 643 212 647
rect 230 644 231 648
rect 235 644 236 648
rect 230 643 236 644
rect 239 647 245 648
rect 239 643 240 647
rect 244 646 245 647
rect 270 647 276 648
rect 270 646 271 647
rect 244 644 271 646
rect 244 643 245 644
rect 206 642 212 643
rect 239 642 245 643
rect 270 643 271 644
rect 275 643 276 647
rect 294 644 295 648
rect 299 644 300 648
rect 294 643 300 644
rect 303 647 309 648
rect 303 643 304 647
rect 308 646 309 647
rect 358 647 364 648
rect 358 646 359 647
rect 308 644 359 646
rect 308 643 309 644
rect 270 642 276 643
rect 303 642 309 643
rect 358 643 359 644
rect 363 643 364 647
rect 366 644 367 648
rect 371 644 372 648
rect 366 643 372 644
rect 438 648 444 649
rect 438 644 439 648
rect 443 644 444 648
rect 438 643 444 644
rect 518 648 524 649
rect 518 644 519 648
rect 523 644 524 648
rect 518 643 524 644
rect 598 648 604 649
rect 598 644 599 648
rect 603 644 604 648
rect 598 643 604 644
rect 654 648 660 649
rect 654 644 655 648
rect 659 644 660 648
rect 686 645 687 649
rect 691 645 692 649
rect 686 644 692 645
rect 654 643 660 644
rect 358 642 364 643
rect 607 635 613 636
rect 158 633 164 634
rect 110 631 116 632
rect 110 627 111 631
rect 115 627 116 631
rect 158 629 159 633
rect 163 629 164 633
rect 158 628 164 629
rect 214 633 220 634
rect 214 629 215 633
rect 219 629 220 633
rect 214 628 220 629
rect 278 633 284 634
rect 278 629 279 633
rect 283 629 284 633
rect 278 628 284 629
rect 350 633 356 634
rect 350 629 351 633
rect 355 629 356 633
rect 350 628 356 629
rect 422 633 428 634
rect 422 629 423 633
rect 427 629 428 633
rect 422 628 428 629
rect 502 633 508 634
rect 502 629 503 633
rect 507 629 508 633
rect 502 628 508 629
rect 582 633 588 634
rect 582 629 583 633
rect 587 629 588 633
rect 607 631 608 635
rect 612 634 613 635
rect 615 635 621 636
rect 615 634 616 635
rect 612 632 616 634
rect 612 631 613 632
rect 607 630 613 631
rect 615 631 616 632
rect 620 631 621 635
rect 615 630 621 631
rect 638 633 644 634
rect 582 628 588 629
rect 638 629 639 633
rect 643 629 644 633
rect 638 628 644 629
rect 686 631 692 632
rect 110 626 116 627
rect 222 627 228 628
rect 222 623 223 627
rect 227 626 228 627
rect 375 627 381 628
rect 375 626 376 627
rect 227 624 376 626
rect 227 623 228 624
rect 222 622 228 623
rect 375 623 376 624
rect 380 623 381 627
rect 375 622 381 623
rect 447 627 453 628
rect 447 623 448 627
rect 452 626 453 627
rect 494 627 500 628
rect 494 626 495 627
rect 452 624 495 626
rect 452 623 453 624
rect 447 622 453 623
rect 494 623 495 624
rect 499 623 500 627
rect 494 622 500 623
rect 510 627 516 628
rect 510 623 511 627
rect 515 626 516 627
rect 527 627 533 628
rect 527 626 528 627
rect 515 624 528 626
rect 515 623 516 624
rect 510 622 516 623
rect 527 623 528 624
rect 532 623 533 627
rect 527 622 533 623
rect 630 627 636 628
rect 630 623 631 627
rect 635 626 636 627
rect 663 627 669 628
rect 663 626 664 627
rect 635 624 664 626
rect 635 623 636 624
rect 630 622 636 623
rect 663 623 664 624
rect 668 623 669 627
rect 686 627 687 631
rect 691 627 692 631
rect 686 626 692 627
rect 663 622 669 623
rect 186 603 192 604
rect 186 599 187 603
rect 191 602 192 603
rect 262 603 268 604
rect 191 600 210 602
rect 191 599 192 600
rect 186 598 192 599
rect 208 598 210 600
rect 223 599 229 600
rect 223 598 224 599
rect 110 597 116 598
rect 110 593 111 597
rect 115 593 116 597
rect 208 596 224 598
rect 110 592 116 593
rect 198 595 204 596
rect 198 591 199 595
rect 203 591 204 595
rect 223 595 224 596
rect 228 595 229 599
rect 262 599 263 603
rect 267 602 268 603
rect 267 600 321 602
rect 267 599 268 600
rect 262 598 268 599
rect 319 599 325 600
rect 223 594 229 595
rect 238 595 244 596
rect 198 590 204 591
rect 238 591 239 595
rect 243 591 244 595
rect 238 590 244 591
rect 294 595 300 596
rect 294 591 295 595
rect 299 591 300 595
rect 319 595 320 599
rect 324 595 325 599
rect 662 599 669 600
rect 319 594 325 595
rect 350 595 356 596
rect 294 590 300 591
rect 350 591 351 595
rect 355 591 356 595
rect 350 590 356 591
rect 414 595 420 596
rect 414 591 415 595
rect 419 591 420 595
rect 414 590 420 591
rect 486 595 492 596
rect 486 591 487 595
rect 491 591 492 595
rect 486 590 492 591
rect 566 595 572 596
rect 566 591 567 595
rect 571 591 572 595
rect 566 590 572 591
rect 638 595 644 596
rect 638 591 639 595
rect 643 591 644 595
rect 662 595 663 599
rect 668 595 669 599
rect 662 594 669 595
rect 686 597 692 598
rect 686 593 687 597
rect 691 593 692 597
rect 686 592 692 593
rect 638 590 644 591
rect 222 587 228 588
rect 222 583 223 587
rect 227 586 228 587
rect 263 587 269 588
rect 263 586 264 587
rect 227 584 264 586
rect 227 583 228 584
rect 222 582 228 583
rect 263 583 264 584
rect 268 583 269 587
rect 263 582 269 583
rect 343 587 349 588
rect 343 583 344 587
rect 348 586 349 587
rect 375 587 381 588
rect 375 586 376 587
rect 348 584 376 586
rect 348 583 349 584
rect 343 582 349 583
rect 375 583 376 584
rect 380 583 381 587
rect 375 582 381 583
rect 402 587 408 588
rect 402 583 403 587
rect 407 586 408 587
rect 439 587 445 588
rect 439 586 440 587
rect 407 584 440 586
rect 407 583 408 584
rect 402 582 408 583
rect 439 583 440 584
rect 444 583 445 587
rect 439 582 445 583
rect 214 580 220 581
rect 110 579 116 580
rect 110 575 111 579
rect 115 575 116 579
rect 214 576 215 580
rect 219 576 220 580
rect 214 575 220 576
rect 254 580 260 581
rect 254 576 255 580
rect 259 576 260 580
rect 254 575 260 576
rect 310 580 316 581
rect 310 576 311 580
rect 315 576 316 580
rect 310 575 316 576
rect 366 580 372 581
rect 366 576 367 580
rect 371 576 372 580
rect 366 575 372 576
rect 430 580 436 581
rect 430 576 431 580
rect 435 576 436 580
rect 430 575 436 576
rect 502 580 508 581
rect 582 580 588 581
rect 654 580 660 581
rect 502 576 503 580
rect 507 576 508 580
rect 502 575 508 576
rect 511 579 517 580
rect 511 575 512 579
rect 516 578 517 579
rect 516 576 546 578
rect 516 575 517 576
rect 110 574 116 575
rect 511 574 517 575
rect 207 563 213 564
rect 207 559 208 563
rect 212 562 213 563
rect 222 563 228 564
rect 222 562 223 563
rect 212 560 223 562
rect 212 559 213 560
rect 207 558 213 559
rect 222 559 223 560
rect 227 559 228 563
rect 222 558 228 559
rect 247 563 253 564
rect 247 559 248 563
rect 252 562 253 563
rect 262 563 268 564
rect 262 562 263 563
rect 252 560 263 562
rect 252 559 253 560
rect 247 558 253 559
rect 262 559 263 560
rect 267 559 268 563
rect 262 558 268 559
rect 303 563 309 564
rect 303 559 304 563
rect 308 562 309 563
rect 343 563 349 564
rect 343 562 344 563
rect 308 560 344 562
rect 308 559 309 560
rect 303 558 309 559
rect 343 559 344 560
rect 348 559 349 563
rect 343 558 349 559
rect 359 563 365 564
rect 359 559 360 563
rect 364 562 365 563
rect 402 563 408 564
rect 402 562 403 563
rect 364 560 403 562
rect 364 559 365 560
rect 359 558 365 559
rect 402 559 403 560
rect 407 559 408 563
rect 402 558 408 559
rect 418 563 429 564
rect 418 559 419 563
rect 423 559 424 563
rect 428 559 429 563
rect 418 558 429 559
rect 494 563 501 564
rect 494 559 495 563
rect 500 559 501 563
rect 544 562 546 576
rect 582 576 583 580
rect 587 576 588 580
rect 582 575 588 576
rect 590 579 597 580
rect 590 575 591 579
rect 596 575 597 579
rect 654 576 655 580
rect 659 576 660 580
rect 654 575 660 576
rect 686 579 692 580
rect 686 575 687 579
rect 691 575 692 579
rect 590 574 597 575
rect 686 574 692 575
rect 575 563 581 564
rect 575 562 576 563
rect 544 560 576 562
rect 494 558 501 559
rect 575 559 576 560
rect 580 559 581 563
rect 575 558 581 559
rect 626 563 632 564
rect 626 559 627 563
rect 631 562 632 563
rect 647 563 653 564
rect 647 562 648 563
rect 631 560 648 562
rect 631 559 632 560
rect 626 558 632 559
rect 647 559 648 560
rect 652 559 653 563
rect 647 558 653 559
rect 510 555 516 556
rect 510 554 511 555
rect 472 552 511 554
rect 319 549 325 550
rect 319 545 320 549
rect 324 548 325 549
rect 338 549 344 550
rect 338 548 339 549
rect 324 546 339 548
rect 324 545 325 546
rect 319 544 325 545
rect 338 545 339 546
rect 343 545 344 549
rect 338 544 344 545
rect 346 549 352 550
rect 346 545 347 549
rect 351 548 352 549
rect 359 549 365 550
rect 359 548 360 549
rect 351 546 360 548
rect 351 545 352 546
rect 346 544 352 545
rect 359 545 360 546
rect 364 545 365 549
rect 359 544 365 545
rect 386 549 392 550
rect 386 545 387 549
rect 391 548 392 549
rect 399 549 405 550
rect 399 548 400 549
rect 391 546 400 548
rect 391 545 392 546
rect 386 544 392 545
rect 399 545 400 546
rect 404 545 405 549
rect 399 544 405 545
rect 447 549 453 550
rect 447 545 448 549
rect 452 548 453 549
rect 472 548 474 552
rect 510 551 511 552
rect 515 551 516 555
rect 510 550 516 551
rect 590 551 596 552
rect 590 550 591 551
rect 452 546 474 548
rect 495 549 501 550
rect 452 545 453 546
rect 447 544 453 545
rect 495 545 496 549
rect 500 548 501 549
rect 551 549 591 550
rect 500 546 522 548
rect 534 547 540 548
rect 534 546 535 547
rect 500 545 501 546
rect 495 544 501 545
rect 520 544 535 546
rect 534 543 535 544
rect 539 543 540 547
rect 551 545 552 549
rect 556 548 591 549
rect 556 545 557 548
rect 590 547 591 548
rect 595 547 596 551
rect 590 546 596 547
rect 606 549 613 550
rect 551 544 557 545
rect 606 545 607 549
rect 612 545 613 549
rect 606 544 613 545
rect 647 549 653 550
rect 647 545 648 549
rect 652 548 653 549
rect 662 549 668 550
rect 662 548 663 549
rect 652 546 663 548
rect 652 545 653 546
rect 647 544 653 545
rect 662 545 663 546
rect 667 545 668 549
rect 662 544 668 545
rect 534 542 540 543
rect 110 533 116 534
rect 686 533 692 534
rect 110 529 111 533
rect 115 529 116 533
rect 110 528 116 529
rect 326 532 332 533
rect 366 532 372 533
rect 406 532 412 533
rect 454 532 460 533
rect 326 528 327 532
rect 331 528 332 532
rect 326 527 332 528
rect 335 531 341 532
rect 335 527 336 531
rect 340 530 341 531
rect 346 531 352 532
rect 346 530 347 531
rect 340 528 347 530
rect 340 527 341 528
rect 335 526 341 527
rect 346 527 347 528
rect 351 527 352 531
rect 366 528 367 532
rect 371 528 372 532
rect 366 527 372 528
rect 375 531 381 532
rect 375 527 376 531
rect 380 530 381 531
rect 386 531 392 532
rect 386 530 387 531
rect 380 528 387 530
rect 380 527 381 528
rect 346 526 352 527
rect 375 526 381 527
rect 386 527 387 528
rect 391 527 392 531
rect 406 528 407 532
rect 411 528 412 532
rect 406 527 412 528
rect 415 531 424 532
rect 415 527 416 531
rect 423 527 424 531
rect 454 528 455 532
rect 459 528 460 532
rect 454 527 460 528
rect 502 532 508 533
rect 558 532 564 533
rect 502 528 503 532
rect 507 528 508 532
rect 502 527 508 528
rect 510 531 517 532
rect 510 527 511 531
rect 516 527 517 531
rect 558 528 559 532
rect 563 528 564 532
rect 558 527 564 528
rect 614 532 620 533
rect 654 532 660 533
rect 614 528 615 532
rect 619 528 620 532
rect 614 527 620 528
rect 623 531 632 532
rect 623 527 624 531
rect 631 527 632 531
rect 654 528 655 532
rect 659 528 660 532
rect 686 529 687 533
rect 691 529 692 533
rect 686 528 692 529
rect 654 527 660 528
rect 386 526 392 527
rect 415 526 424 527
rect 510 526 517 527
rect 623 526 632 527
rect 310 517 316 518
rect 110 515 116 516
rect 110 511 111 515
rect 115 511 116 515
rect 310 513 311 517
rect 315 513 316 517
rect 310 512 316 513
rect 350 517 356 518
rect 350 513 351 517
rect 355 513 356 517
rect 350 512 356 513
rect 390 517 396 518
rect 390 513 391 517
rect 395 513 396 517
rect 390 512 396 513
rect 438 517 444 518
rect 438 513 439 517
rect 443 513 444 517
rect 438 512 444 513
rect 486 517 492 518
rect 486 513 487 517
rect 491 513 492 517
rect 486 512 492 513
rect 542 517 548 518
rect 542 513 543 517
rect 547 513 548 517
rect 542 512 548 513
rect 598 517 604 518
rect 598 513 599 517
rect 603 513 604 517
rect 598 512 604 513
rect 638 517 644 518
rect 638 513 639 517
rect 643 513 644 517
rect 638 512 644 513
rect 686 515 692 516
rect 110 510 116 511
rect 338 511 344 512
rect 338 507 339 511
rect 343 510 344 511
rect 463 511 469 512
rect 463 510 464 511
rect 343 508 464 510
rect 343 507 344 508
rect 338 506 344 507
rect 463 507 464 508
rect 468 507 469 511
rect 463 506 469 507
rect 567 511 573 512
rect 567 507 568 511
rect 572 510 573 511
rect 590 511 596 512
rect 590 510 591 511
rect 572 508 591 510
rect 572 507 573 508
rect 567 506 573 507
rect 590 507 591 508
rect 595 507 596 511
rect 590 506 596 507
rect 606 511 612 512
rect 606 507 607 511
rect 611 510 612 511
rect 663 511 669 512
rect 663 510 664 511
rect 611 508 664 510
rect 611 507 612 508
rect 606 506 612 507
rect 663 507 664 508
rect 668 507 669 511
rect 686 511 687 515
rect 691 511 692 515
rect 686 510 692 511
rect 663 506 669 507
rect 534 491 541 492
rect 110 489 116 490
rect 110 485 111 489
rect 115 485 116 489
rect 110 484 116 485
rect 254 487 260 488
rect 254 483 255 487
rect 259 483 260 487
rect 254 482 260 483
rect 294 487 300 488
rect 294 483 295 487
rect 299 483 300 487
rect 294 482 300 483
rect 334 487 340 488
rect 334 483 335 487
rect 339 483 340 487
rect 334 482 340 483
rect 390 487 396 488
rect 390 483 391 487
rect 395 483 396 487
rect 390 482 396 483
rect 446 487 452 488
rect 446 483 447 487
rect 451 483 452 487
rect 446 482 452 483
rect 510 487 516 488
rect 510 483 511 487
rect 515 483 516 487
rect 534 487 535 491
rect 540 487 541 491
rect 662 491 669 492
rect 534 486 541 487
rect 582 487 588 488
rect 510 482 516 483
rect 582 483 583 487
rect 587 483 588 487
rect 582 482 588 483
rect 638 487 644 488
rect 638 483 639 487
rect 643 483 644 487
rect 662 487 663 491
rect 668 487 669 491
rect 662 486 669 487
rect 686 489 692 490
rect 686 485 687 489
rect 691 485 692 489
rect 686 484 692 485
rect 638 482 644 483
rect 270 472 276 473
rect 310 472 316 473
rect 350 472 356 473
rect 406 472 412 473
rect 462 472 468 473
rect 526 472 532 473
rect 110 471 116 472
rect 110 467 111 471
rect 115 467 116 471
rect 270 468 271 472
rect 275 468 276 472
rect 270 467 276 468
rect 279 471 285 472
rect 279 467 280 471
rect 284 470 285 471
rect 284 468 294 470
rect 284 467 285 468
rect 110 466 116 467
rect 279 466 285 467
rect 263 455 269 456
rect 263 451 264 455
rect 268 451 269 455
rect 292 454 294 468
rect 310 468 311 472
rect 315 468 316 472
rect 310 467 316 468
rect 319 471 325 472
rect 319 467 320 471
rect 324 470 325 471
rect 324 468 334 470
rect 324 467 325 468
rect 319 466 325 467
rect 303 455 309 456
rect 303 454 304 455
rect 292 452 304 454
rect 263 450 269 451
rect 303 451 304 452
rect 308 451 309 455
rect 332 454 334 468
rect 350 468 351 472
rect 355 468 356 472
rect 350 467 356 468
rect 359 471 365 472
rect 359 467 360 471
rect 364 470 365 471
rect 364 468 382 470
rect 364 467 365 468
rect 359 466 365 467
rect 343 455 349 456
rect 343 454 344 455
rect 332 452 344 454
rect 303 450 309 451
rect 343 451 344 452
rect 348 451 349 455
rect 380 454 382 468
rect 406 468 407 472
rect 411 468 412 472
rect 406 467 412 468
rect 415 471 421 472
rect 415 467 416 471
rect 420 470 421 471
rect 420 468 438 470
rect 420 467 421 468
rect 415 466 421 467
rect 399 455 405 456
rect 399 454 400 455
rect 380 452 400 454
rect 343 450 349 451
rect 399 451 400 452
rect 404 451 405 455
rect 436 454 438 468
rect 462 468 463 472
rect 467 468 468 472
rect 462 467 468 468
rect 471 471 477 472
rect 471 467 472 471
rect 476 470 477 471
rect 476 468 498 470
rect 476 467 477 468
rect 471 466 477 467
rect 455 455 461 456
rect 455 454 456 455
rect 436 452 456 454
rect 399 450 405 451
rect 455 451 456 452
rect 460 451 461 455
rect 496 454 498 468
rect 526 468 527 472
rect 531 468 532 472
rect 526 467 532 468
rect 598 472 604 473
rect 654 472 660 473
rect 598 468 599 472
rect 603 468 604 472
rect 598 467 604 468
rect 606 471 613 472
rect 606 467 607 471
rect 612 467 613 471
rect 654 468 655 472
rect 659 468 660 472
rect 654 467 660 468
rect 686 471 692 472
rect 686 467 687 471
rect 691 467 692 471
rect 606 466 613 467
rect 686 466 692 467
rect 519 455 525 456
rect 519 454 520 455
rect 496 452 520 454
rect 455 450 461 451
rect 519 451 520 452
rect 524 451 525 455
rect 519 450 525 451
rect 590 455 597 456
rect 590 451 591 455
rect 596 451 597 455
rect 590 450 597 451
rect 647 455 653 456
rect 647 451 648 455
rect 652 454 653 455
rect 662 455 668 456
rect 662 454 663 455
rect 652 452 663 454
rect 652 451 653 452
rect 647 450 653 451
rect 662 451 663 452
rect 667 451 668 455
rect 662 450 668 451
rect 265 446 267 450
rect 502 447 508 448
rect 502 446 503 447
rect 265 444 503 446
rect 502 443 503 444
rect 507 443 508 447
rect 502 442 508 443
rect 606 443 612 444
rect 606 442 607 443
rect 167 441 173 442
rect 167 437 168 441
rect 172 440 173 441
rect 182 441 188 442
rect 182 440 183 441
rect 172 438 183 440
rect 172 437 173 438
rect 167 436 173 437
rect 182 437 183 438
rect 187 437 188 441
rect 182 436 188 437
rect 199 441 205 442
rect 199 437 200 441
rect 204 440 205 441
rect 215 441 221 442
rect 215 440 216 441
rect 204 438 216 440
rect 204 437 205 438
rect 199 436 205 437
rect 215 437 216 438
rect 220 437 221 441
rect 215 436 221 437
rect 254 441 260 442
rect 254 437 255 441
rect 259 440 260 441
rect 271 441 277 442
rect 271 440 272 441
rect 259 438 272 440
rect 259 437 260 438
rect 254 436 260 437
rect 271 437 272 438
rect 276 437 277 441
rect 271 436 277 437
rect 334 441 341 442
rect 334 437 335 441
rect 340 437 341 441
rect 334 436 341 437
rect 390 441 396 442
rect 390 437 391 441
rect 395 440 396 441
rect 407 441 413 442
rect 407 440 408 441
rect 395 438 408 440
rect 395 437 396 438
rect 390 436 396 437
rect 407 437 408 438
rect 412 437 413 441
rect 407 436 413 437
rect 470 441 476 442
rect 470 437 471 441
rect 475 440 476 441
rect 487 441 493 442
rect 487 440 488 441
rect 475 438 488 440
rect 475 437 476 438
rect 470 436 476 437
rect 487 437 488 438
rect 492 437 493 441
rect 487 436 493 437
rect 575 441 581 442
rect 575 437 576 441
rect 580 440 581 441
rect 592 440 607 442
rect 580 438 594 440
rect 606 439 607 440
rect 611 439 612 443
rect 606 438 612 439
rect 646 441 653 442
rect 580 437 581 438
rect 575 436 581 437
rect 646 437 647 441
rect 652 437 653 441
rect 646 436 653 437
rect 110 425 116 426
rect 686 425 692 426
rect 110 421 111 425
rect 115 421 116 425
rect 110 420 116 421
rect 174 424 180 425
rect 222 424 228 425
rect 278 424 284 425
rect 342 424 348 425
rect 414 424 420 425
rect 494 424 500 425
rect 582 424 588 425
rect 174 420 175 424
rect 179 420 180 424
rect 174 419 180 420
rect 183 423 189 424
rect 183 419 184 423
rect 188 422 189 423
rect 199 423 205 424
rect 199 422 200 423
rect 188 420 200 422
rect 188 419 189 420
rect 183 418 189 419
rect 199 419 200 420
rect 204 419 205 423
rect 222 420 223 424
rect 227 420 228 424
rect 222 419 228 420
rect 231 423 237 424
rect 231 419 232 423
rect 236 422 237 423
rect 254 423 260 424
rect 254 422 255 423
rect 236 420 255 422
rect 236 419 237 420
rect 199 418 205 419
rect 231 418 237 419
rect 254 419 255 420
rect 259 419 260 423
rect 278 420 279 424
rect 283 420 284 424
rect 278 419 284 420
rect 287 423 293 424
rect 287 419 288 423
rect 292 422 293 423
rect 334 423 340 424
rect 334 422 335 423
rect 292 420 335 422
rect 292 419 293 420
rect 254 418 260 419
rect 287 418 293 419
rect 334 419 335 420
rect 339 419 340 423
rect 342 420 343 424
rect 347 420 348 424
rect 342 419 348 420
rect 351 423 357 424
rect 351 419 352 423
rect 356 422 357 423
rect 390 423 396 424
rect 390 422 391 423
rect 356 420 391 422
rect 356 419 357 420
rect 334 418 340 419
rect 351 418 357 419
rect 390 419 391 420
rect 395 419 396 423
rect 414 420 415 424
rect 419 420 420 424
rect 414 419 420 420
rect 423 423 429 424
rect 423 419 424 423
rect 428 422 429 423
rect 470 423 476 424
rect 470 422 471 423
rect 428 420 471 422
rect 428 419 429 420
rect 390 418 396 419
rect 423 418 429 419
rect 470 419 471 420
rect 475 419 476 423
rect 494 420 495 424
rect 499 420 500 424
rect 494 419 500 420
rect 502 423 509 424
rect 502 419 503 423
rect 508 419 509 423
rect 582 420 583 424
rect 587 420 588 424
rect 582 419 588 420
rect 654 424 660 425
rect 654 420 655 424
rect 659 420 660 424
rect 654 419 660 420
rect 662 423 669 424
rect 662 419 663 423
rect 668 419 669 423
rect 686 421 687 425
rect 691 421 692 425
rect 686 420 692 421
rect 470 418 476 419
rect 502 418 509 419
rect 662 418 669 419
rect 158 409 164 410
rect 110 407 116 408
rect 110 403 111 407
rect 115 403 116 407
rect 158 405 159 409
rect 163 405 164 409
rect 158 404 164 405
rect 206 409 212 410
rect 206 405 207 409
rect 211 405 212 409
rect 206 404 212 405
rect 262 409 268 410
rect 262 405 263 409
rect 267 405 268 409
rect 262 404 268 405
rect 326 409 332 410
rect 326 405 327 409
rect 331 405 332 409
rect 326 404 332 405
rect 398 409 404 410
rect 398 405 399 409
rect 403 405 404 409
rect 398 404 404 405
rect 478 409 484 410
rect 478 405 479 409
rect 483 405 484 409
rect 478 404 484 405
rect 566 409 572 410
rect 566 405 567 409
rect 571 405 572 409
rect 566 404 572 405
rect 638 409 644 410
rect 638 405 639 409
rect 643 405 644 409
rect 638 404 644 405
rect 686 407 692 408
rect 110 402 116 403
rect 546 403 552 404
rect 546 399 547 403
rect 551 402 552 403
rect 591 403 597 404
rect 591 402 592 403
rect 551 400 592 402
rect 551 399 552 400
rect 546 398 552 399
rect 591 399 592 400
rect 596 399 597 403
rect 686 403 687 407
rect 691 403 692 407
rect 686 402 692 403
rect 591 398 597 399
rect 182 383 188 384
rect 182 379 183 383
rect 187 379 188 383
rect 247 383 253 384
rect 182 378 188 379
rect 199 379 205 380
rect 199 378 200 379
rect 110 377 116 378
rect 110 373 111 377
rect 115 373 116 377
rect 184 376 200 378
rect 110 372 116 373
rect 134 375 140 376
rect 134 371 135 375
rect 139 371 140 375
rect 134 370 140 371
rect 174 375 180 376
rect 174 371 175 375
rect 179 371 180 375
rect 199 375 200 376
rect 204 375 205 379
rect 247 379 248 383
rect 252 382 253 383
rect 646 383 652 384
rect 252 380 307 382
rect 252 379 253 380
rect 247 378 253 379
rect 303 379 309 380
rect 199 374 205 375
rect 214 375 220 376
rect 174 370 180 371
rect 214 371 215 375
rect 219 371 220 375
rect 214 370 220 371
rect 278 375 284 376
rect 278 371 279 375
rect 283 371 284 375
rect 303 375 304 379
rect 308 375 309 379
rect 646 379 647 383
rect 651 382 652 383
rect 651 380 667 382
rect 651 379 652 380
rect 646 378 652 379
rect 663 379 669 380
rect 303 374 309 375
rect 342 375 348 376
rect 278 370 284 371
rect 342 371 343 375
rect 347 371 348 375
rect 342 370 348 371
rect 414 375 420 376
rect 414 371 415 375
rect 419 371 420 375
rect 414 370 420 371
rect 494 375 500 376
rect 494 371 495 375
rect 499 371 500 375
rect 494 370 500 371
rect 574 375 580 376
rect 574 371 575 375
rect 579 371 580 375
rect 574 370 580 371
rect 638 375 644 376
rect 638 371 639 375
rect 643 371 644 375
rect 663 375 664 379
rect 668 375 669 379
rect 663 374 669 375
rect 686 377 692 378
rect 686 373 687 377
rect 691 373 692 377
rect 686 372 692 373
rect 638 370 644 371
rect 158 367 164 368
rect 158 363 159 367
rect 163 366 164 367
rect 239 367 245 368
rect 239 366 240 367
rect 163 364 240 366
rect 163 363 164 364
rect 158 362 164 363
rect 239 363 240 364
rect 244 363 245 367
rect 239 362 245 363
rect 302 367 308 368
rect 302 363 303 367
rect 307 366 308 367
rect 439 367 445 368
rect 439 366 440 367
rect 307 364 440 366
rect 307 363 308 364
rect 302 362 308 363
rect 439 363 440 364
rect 444 363 445 367
rect 439 362 445 363
rect 150 360 156 361
rect 190 360 196 361
rect 110 359 116 360
rect 110 355 111 359
rect 115 355 116 359
rect 150 356 151 360
rect 155 356 156 360
rect 150 355 156 356
rect 159 359 165 360
rect 159 355 160 359
rect 164 358 165 359
rect 164 356 174 358
rect 164 355 165 356
rect 110 354 116 355
rect 159 354 165 355
rect 143 343 149 344
rect 143 339 144 343
rect 148 342 149 343
rect 158 343 164 344
rect 158 342 159 343
rect 148 340 159 342
rect 148 339 149 340
rect 143 338 149 339
rect 158 339 159 340
rect 163 339 164 343
rect 172 342 174 356
rect 190 356 191 360
rect 195 356 196 360
rect 190 355 196 356
rect 230 360 236 361
rect 230 356 231 360
rect 235 356 236 360
rect 230 355 236 356
rect 294 360 300 361
rect 294 356 295 360
rect 299 356 300 360
rect 294 355 300 356
rect 358 360 364 361
rect 430 360 436 361
rect 358 356 359 360
rect 363 356 364 360
rect 358 355 364 356
rect 367 359 373 360
rect 367 355 368 359
rect 372 358 373 359
rect 372 356 398 358
rect 372 355 373 356
rect 367 354 373 355
rect 183 343 189 344
rect 183 342 184 343
rect 172 340 184 342
rect 158 338 164 339
rect 183 339 184 340
rect 188 339 189 343
rect 183 338 189 339
rect 223 343 229 344
rect 223 339 224 343
rect 228 342 229 343
rect 247 343 253 344
rect 247 342 248 343
rect 228 340 248 342
rect 228 339 229 340
rect 223 338 229 339
rect 247 339 248 340
rect 252 339 253 343
rect 247 338 253 339
rect 287 343 293 344
rect 287 339 288 343
rect 292 342 293 343
rect 302 343 308 344
rect 302 342 303 343
rect 292 340 303 342
rect 292 339 293 340
rect 287 338 293 339
rect 302 339 303 340
rect 307 339 308 343
rect 302 338 308 339
rect 346 343 357 344
rect 346 339 347 343
rect 351 339 352 343
rect 356 339 357 343
rect 396 342 398 356
rect 430 356 431 360
rect 435 356 436 360
rect 430 355 436 356
rect 510 360 516 361
rect 590 360 596 361
rect 654 360 660 361
rect 510 356 511 360
rect 515 356 516 360
rect 510 355 516 356
rect 518 359 525 360
rect 518 355 519 359
rect 524 355 525 359
rect 590 356 591 360
rect 595 356 596 360
rect 590 355 596 356
rect 599 359 605 360
rect 599 355 600 359
rect 604 358 605 359
rect 604 356 626 358
rect 604 355 605 356
rect 518 354 525 355
rect 599 354 605 355
rect 423 343 429 344
rect 423 342 424 343
rect 396 340 424 342
rect 346 338 357 339
rect 423 339 424 340
rect 428 339 429 343
rect 423 338 429 339
rect 503 343 509 344
rect 503 339 504 343
rect 508 342 509 343
rect 546 343 552 344
rect 546 342 547 343
rect 508 340 547 342
rect 508 339 509 340
rect 503 338 509 339
rect 546 339 547 340
rect 551 339 552 343
rect 546 338 552 339
rect 583 343 589 344
rect 583 339 584 343
rect 588 342 589 343
rect 606 343 612 344
rect 606 342 607 343
rect 588 340 607 342
rect 588 339 589 340
rect 583 338 589 339
rect 606 339 607 340
rect 611 339 612 343
rect 624 342 626 356
rect 654 356 655 360
rect 659 356 660 360
rect 654 355 660 356
rect 686 359 692 360
rect 686 355 687 359
rect 691 355 692 359
rect 686 354 692 355
rect 647 343 653 344
rect 647 342 648 343
rect 624 340 648 342
rect 606 338 612 339
rect 647 339 648 340
rect 652 339 653 343
rect 647 338 653 339
rect 438 331 444 332
rect 438 330 439 331
rect 400 328 439 330
rect 314 327 320 328
rect 247 325 253 326
rect 247 321 248 325
rect 252 324 253 325
rect 266 325 272 326
rect 266 324 267 325
rect 252 322 267 324
rect 252 321 253 322
rect 247 320 253 321
rect 266 321 267 322
rect 271 321 272 325
rect 266 320 272 321
rect 274 325 280 326
rect 274 321 275 325
rect 279 324 280 325
rect 287 325 293 326
rect 287 324 288 325
rect 279 322 288 324
rect 279 321 280 322
rect 274 320 280 321
rect 287 321 288 322
rect 292 321 293 325
rect 314 323 315 327
rect 319 326 320 327
rect 319 324 321 326
rect 327 325 333 326
rect 327 324 328 325
rect 319 323 328 324
rect 314 322 328 323
rect 287 320 293 321
rect 327 321 328 322
rect 332 321 333 325
rect 327 320 333 321
rect 375 325 381 326
rect 375 321 376 325
rect 380 324 381 325
rect 400 324 402 328
rect 438 327 439 328
rect 443 327 444 331
rect 486 331 492 332
rect 486 330 487 331
rect 438 326 444 327
rect 448 328 487 330
rect 380 322 402 324
rect 423 325 429 326
rect 380 321 381 322
rect 375 320 381 321
rect 423 321 424 325
rect 428 324 429 325
rect 448 324 450 328
rect 486 327 487 328
rect 491 327 492 331
rect 486 326 492 327
rect 428 322 450 324
rect 470 325 477 326
rect 428 321 429 322
rect 423 320 429 321
rect 470 321 471 325
rect 476 321 477 325
rect 470 320 477 321
rect 518 325 525 326
rect 518 321 519 325
rect 524 321 525 325
rect 518 320 525 321
rect 551 325 557 326
rect 551 321 552 325
rect 556 324 557 325
rect 567 325 573 326
rect 567 324 568 325
rect 556 322 568 324
rect 556 321 557 322
rect 551 320 557 321
rect 567 321 568 322
rect 572 321 573 325
rect 567 320 573 321
rect 607 325 613 326
rect 607 321 608 325
rect 612 324 613 325
rect 626 325 632 326
rect 626 324 627 325
rect 612 322 627 324
rect 612 321 613 322
rect 607 320 613 321
rect 626 321 627 322
rect 631 321 632 325
rect 626 320 632 321
rect 647 325 653 326
rect 647 321 648 325
rect 652 324 653 325
rect 662 325 668 326
rect 662 324 663 325
rect 652 322 663 324
rect 652 321 653 322
rect 647 320 653 321
rect 662 321 663 322
rect 667 321 668 325
rect 662 320 668 321
rect 110 309 116 310
rect 686 309 692 310
rect 110 305 111 309
rect 115 305 116 309
rect 110 304 116 305
rect 254 308 260 309
rect 294 308 300 309
rect 334 308 340 309
rect 382 308 388 309
rect 254 304 255 308
rect 259 304 260 308
rect 254 303 260 304
rect 263 307 269 308
rect 263 303 264 307
rect 268 306 269 307
rect 274 307 280 308
rect 274 306 275 307
rect 268 304 275 306
rect 268 303 269 304
rect 263 302 269 303
rect 274 303 275 304
rect 279 303 280 307
rect 294 304 295 308
rect 299 304 300 308
rect 294 303 300 304
rect 303 307 309 308
rect 303 303 304 307
rect 308 306 309 307
rect 314 307 320 308
rect 314 306 315 307
rect 308 304 315 306
rect 308 303 309 304
rect 274 302 280 303
rect 303 302 309 303
rect 314 303 315 304
rect 319 303 320 307
rect 334 304 335 308
rect 339 304 340 308
rect 334 303 340 304
rect 343 307 352 308
rect 343 303 344 307
rect 351 303 352 307
rect 382 304 383 308
rect 387 304 388 308
rect 382 303 388 304
rect 430 308 436 309
rect 478 308 484 309
rect 526 308 532 309
rect 574 308 580 309
rect 430 304 431 308
rect 435 304 436 308
rect 430 303 436 304
rect 438 307 445 308
rect 438 303 439 307
rect 444 303 445 307
rect 478 304 479 308
rect 483 304 484 308
rect 478 303 484 304
rect 486 307 493 308
rect 486 303 487 307
rect 492 303 493 307
rect 526 304 527 308
rect 531 304 532 308
rect 526 303 532 304
rect 535 307 541 308
rect 535 303 536 307
rect 540 306 541 307
rect 551 307 557 308
rect 551 306 552 307
rect 540 304 552 306
rect 540 303 541 304
rect 314 302 320 303
rect 343 302 352 303
rect 438 302 445 303
rect 486 302 493 303
rect 535 302 541 303
rect 551 303 552 304
rect 556 303 557 307
rect 574 304 575 308
rect 579 304 580 308
rect 574 303 580 304
rect 614 308 620 309
rect 614 304 615 308
rect 619 304 620 308
rect 614 303 620 304
rect 654 308 660 309
rect 654 304 655 308
rect 659 304 660 308
rect 686 305 687 309
rect 691 305 692 309
rect 686 304 692 305
rect 654 303 660 304
rect 551 302 557 303
rect 626 295 632 296
rect 238 293 244 294
rect 110 291 116 292
rect 110 287 111 291
rect 115 287 116 291
rect 238 289 239 293
rect 243 289 244 293
rect 238 288 244 289
rect 278 293 284 294
rect 278 289 279 293
rect 283 289 284 293
rect 278 288 284 289
rect 318 293 324 294
rect 318 289 319 293
rect 323 289 324 293
rect 318 288 324 289
rect 366 293 372 294
rect 366 289 367 293
rect 371 289 372 293
rect 366 288 372 289
rect 414 293 420 294
rect 414 289 415 293
rect 419 289 420 293
rect 414 288 420 289
rect 462 293 468 294
rect 462 289 463 293
rect 467 289 468 293
rect 462 288 468 289
rect 510 293 516 294
rect 510 289 511 293
rect 515 289 516 293
rect 510 288 516 289
rect 558 293 564 294
rect 558 289 559 293
rect 563 289 564 293
rect 558 288 564 289
rect 598 293 604 294
rect 598 289 599 293
rect 603 289 604 293
rect 626 291 627 295
rect 631 294 632 295
rect 631 291 634 294
rect 626 290 634 291
rect 598 288 604 289
rect 110 286 116 287
rect 266 287 272 288
rect 266 283 267 287
rect 271 286 272 287
rect 391 287 397 288
rect 391 286 392 287
rect 271 284 392 286
rect 271 283 272 284
rect 266 282 272 283
rect 391 283 392 284
rect 396 283 397 287
rect 391 282 397 283
rect 502 287 508 288
rect 502 283 503 287
rect 507 286 508 287
rect 583 287 589 288
rect 583 286 584 287
rect 507 284 584 286
rect 507 283 508 284
rect 502 282 508 283
rect 583 283 584 284
rect 588 283 589 287
rect 583 282 589 283
rect 606 287 612 288
rect 606 283 607 287
rect 611 286 612 287
rect 623 287 629 288
rect 623 286 624 287
rect 611 284 624 286
rect 611 283 612 284
rect 606 282 612 283
rect 623 283 624 284
rect 628 283 629 287
rect 632 286 634 290
rect 638 293 644 294
rect 638 289 639 293
rect 643 289 644 293
rect 638 288 644 289
rect 686 291 692 292
rect 663 287 669 288
rect 663 286 664 287
rect 632 284 664 286
rect 623 282 629 283
rect 663 283 664 284
rect 668 283 669 287
rect 686 287 687 291
rect 691 287 692 291
rect 686 286 692 287
rect 663 282 669 283
rect 662 267 669 268
rect 110 265 116 266
rect 110 261 111 265
rect 115 261 116 265
rect 110 260 116 261
rect 238 263 244 264
rect 238 259 239 263
rect 243 259 244 263
rect 238 258 244 259
rect 278 263 284 264
rect 278 259 279 263
rect 283 259 284 263
rect 278 258 284 259
rect 318 263 324 264
rect 318 259 319 263
rect 323 259 324 263
rect 318 258 324 259
rect 358 263 364 264
rect 358 259 359 263
rect 363 259 364 263
rect 358 258 364 259
rect 398 263 404 264
rect 398 259 399 263
rect 403 259 404 263
rect 398 258 404 259
rect 438 263 444 264
rect 438 259 439 263
rect 443 259 444 263
rect 438 258 444 259
rect 462 263 469 264
rect 462 259 463 263
rect 468 259 469 263
rect 462 258 469 259
rect 478 263 484 264
rect 478 259 479 263
rect 483 259 484 263
rect 478 258 484 259
rect 518 263 524 264
rect 518 259 519 263
rect 523 259 524 263
rect 518 258 524 259
rect 558 263 564 264
rect 558 259 559 263
rect 563 259 564 263
rect 558 258 564 259
rect 598 263 604 264
rect 598 259 599 263
rect 603 259 604 263
rect 598 258 604 259
rect 638 263 644 264
rect 638 259 639 263
rect 643 259 644 263
rect 662 263 663 267
rect 668 263 669 267
rect 662 262 669 263
rect 686 265 692 266
rect 686 261 687 265
rect 691 261 692 265
rect 686 260 692 261
rect 638 258 644 259
rect 254 248 260 249
rect 294 248 300 249
rect 334 248 340 249
rect 374 248 380 249
rect 414 248 420 249
rect 454 248 460 249
rect 110 247 116 248
rect 110 243 111 247
rect 115 243 116 247
rect 254 244 255 248
rect 259 244 260 248
rect 254 243 260 244
rect 263 247 269 248
rect 263 243 264 247
rect 268 246 269 247
rect 268 244 278 246
rect 268 243 269 244
rect 110 242 116 243
rect 263 242 269 243
rect 247 231 253 232
rect 247 227 248 231
rect 252 230 253 231
rect 263 231 269 232
rect 263 230 264 231
rect 252 228 264 230
rect 252 227 253 228
rect 247 226 253 227
rect 263 227 264 228
rect 268 227 269 231
rect 276 230 278 244
rect 294 244 295 248
rect 299 244 300 248
rect 294 243 300 244
rect 303 247 309 248
rect 303 243 304 247
rect 308 246 309 247
rect 308 244 314 246
rect 308 243 309 244
rect 303 242 309 243
rect 287 231 293 232
rect 287 230 288 231
rect 276 228 288 230
rect 263 226 269 227
rect 287 227 288 228
rect 292 227 293 231
rect 312 230 314 244
rect 334 244 335 248
rect 339 244 340 248
rect 334 243 340 244
rect 343 247 349 248
rect 343 243 344 247
rect 348 246 349 247
rect 348 244 358 246
rect 348 243 349 244
rect 343 242 349 243
rect 327 231 333 232
rect 327 230 328 231
rect 312 228 328 230
rect 287 226 293 227
rect 327 227 328 228
rect 332 227 333 231
rect 356 230 358 244
rect 374 244 375 248
rect 379 244 380 248
rect 374 243 380 244
rect 383 247 389 248
rect 383 243 384 247
rect 388 246 389 247
rect 388 244 398 246
rect 388 243 389 244
rect 383 242 389 243
rect 367 231 373 232
rect 367 230 368 231
rect 356 228 368 230
rect 327 226 333 227
rect 367 227 368 228
rect 372 227 373 231
rect 396 230 398 244
rect 414 244 415 248
rect 419 244 420 248
rect 414 243 420 244
rect 423 247 429 248
rect 423 243 424 247
rect 428 246 429 247
rect 428 244 438 246
rect 428 243 429 244
rect 423 242 429 243
rect 407 231 413 232
rect 407 230 408 231
rect 396 228 408 230
rect 367 226 373 227
rect 407 227 408 228
rect 412 227 413 231
rect 436 230 438 244
rect 454 244 455 248
rect 459 244 460 248
rect 454 243 460 244
rect 494 248 500 249
rect 534 248 540 249
rect 574 248 580 249
rect 614 248 620 249
rect 654 248 660 249
rect 494 244 495 248
rect 499 244 500 248
rect 494 243 500 244
rect 503 247 509 248
rect 503 243 504 247
rect 508 246 509 247
rect 508 244 518 246
rect 508 243 509 244
rect 503 242 509 243
rect 447 231 453 232
rect 447 230 448 231
rect 436 228 448 230
rect 407 226 413 227
rect 447 227 448 228
rect 452 227 453 231
rect 447 226 453 227
rect 487 231 493 232
rect 487 227 488 231
rect 492 230 493 231
rect 502 231 508 232
rect 502 230 503 231
rect 492 228 503 230
rect 492 227 493 228
rect 487 226 493 227
rect 502 227 503 228
rect 507 227 508 231
rect 516 230 518 244
rect 534 244 535 248
rect 539 244 540 248
rect 534 243 540 244
rect 543 247 549 248
rect 543 243 544 247
rect 548 246 549 247
rect 548 244 558 246
rect 548 243 549 244
rect 543 242 549 243
rect 527 231 533 232
rect 527 230 528 231
rect 516 228 528 230
rect 502 226 508 227
rect 527 227 528 228
rect 532 227 533 231
rect 556 230 558 244
rect 574 244 575 248
rect 579 244 580 248
rect 574 243 580 244
rect 583 247 589 248
rect 583 243 584 247
rect 588 246 589 247
rect 588 244 598 246
rect 588 243 589 244
rect 583 242 589 243
rect 567 231 573 232
rect 567 230 568 231
rect 556 228 568 230
rect 527 226 533 227
rect 567 227 568 228
rect 572 227 573 231
rect 596 230 598 244
rect 614 244 615 248
rect 619 244 620 248
rect 614 243 620 244
rect 623 247 629 248
rect 623 243 624 247
rect 628 246 629 247
rect 628 244 638 246
rect 628 243 629 244
rect 623 242 629 243
rect 607 231 613 232
rect 607 230 608 231
rect 596 228 608 230
rect 567 226 573 227
rect 607 227 608 228
rect 612 227 613 231
rect 636 230 638 244
rect 654 244 655 248
rect 659 244 660 248
rect 654 243 660 244
rect 686 247 692 248
rect 686 243 687 247
rect 691 243 692 247
rect 686 242 692 243
rect 647 231 653 232
rect 647 230 648 231
rect 636 228 648 230
rect 607 226 613 227
rect 647 227 648 228
rect 652 227 653 231
rect 647 226 653 227
rect 198 205 205 206
rect 198 201 199 205
rect 204 201 205 205
rect 198 200 205 201
rect 226 205 232 206
rect 226 201 227 205
rect 231 204 232 205
rect 239 205 245 206
rect 239 204 240 205
rect 231 202 240 204
rect 231 201 232 202
rect 226 200 232 201
rect 239 201 240 202
rect 244 201 245 205
rect 239 200 245 201
rect 262 205 268 206
rect 262 201 263 205
rect 267 204 268 205
rect 279 205 285 206
rect 279 204 280 205
rect 267 202 280 204
rect 267 201 268 202
rect 262 200 268 201
rect 279 201 280 202
rect 284 201 285 205
rect 319 205 325 206
rect 319 202 320 205
rect 279 200 285 201
rect 308 201 320 202
rect 324 201 325 205
rect 308 200 325 201
rect 346 205 352 206
rect 346 201 347 205
rect 351 204 352 205
rect 359 205 365 206
rect 359 204 360 205
rect 351 202 360 204
rect 351 201 352 202
rect 346 200 352 201
rect 359 201 360 202
rect 364 201 365 205
rect 359 200 365 201
rect 386 205 392 206
rect 386 201 387 205
rect 391 204 392 205
rect 399 205 405 206
rect 399 204 400 205
rect 391 202 400 204
rect 391 201 392 202
rect 386 200 392 201
rect 399 201 400 202
rect 404 201 405 205
rect 399 200 405 201
rect 110 189 116 190
rect 110 185 111 189
rect 115 185 116 189
rect 110 184 116 185
rect 206 188 212 189
rect 246 188 252 189
rect 206 184 207 188
rect 211 184 212 188
rect 206 183 212 184
rect 215 187 221 188
rect 215 183 216 187
rect 220 186 221 187
rect 226 187 232 188
rect 226 186 227 187
rect 220 184 227 186
rect 220 183 221 184
rect 215 182 221 183
rect 226 183 227 184
rect 231 183 232 187
rect 246 184 247 188
rect 251 184 252 188
rect 246 183 252 184
rect 286 188 292 189
rect 286 184 287 188
rect 291 184 292 188
rect 286 183 292 184
rect 295 187 301 188
rect 295 183 296 187
rect 300 186 301 187
rect 308 186 310 200
rect 686 189 692 190
rect 300 184 310 186
rect 326 188 332 189
rect 366 188 372 189
rect 406 188 412 189
rect 326 184 327 188
rect 331 184 332 188
rect 300 183 301 184
rect 326 183 332 184
rect 335 187 341 188
rect 335 183 336 187
rect 340 186 341 187
rect 346 187 352 188
rect 346 186 347 187
rect 340 184 347 186
rect 340 183 341 184
rect 226 182 232 183
rect 295 182 301 183
rect 335 182 341 183
rect 346 183 347 184
rect 351 183 352 187
rect 366 184 367 188
rect 371 184 372 188
rect 366 183 372 184
rect 375 187 381 188
rect 375 183 376 187
rect 380 186 381 187
rect 386 187 392 188
rect 386 186 387 187
rect 380 184 387 186
rect 380 183 381 184
rect 346 182 352 183
rect 375 182 381 183
rect 386 183 387 184
rect 391 183 392 187
rect 406 184 407 188
rect 411 184 412 188
rect 686 185 687 189
rect 691 185 692 189
rect 686 184 692 185
rect 406 183 412 184
rect 386 182 392 183
rect 190 173 196 174
rect 110 171 116 172
rect 110 167 111 171
rect 115 167 116 171
rect 190 169 191 173
rect 195 169 196 173
rect 190 168 196 169
rect 230 173 236 174
rect 230 169 231 173
rect 235 169 236 173
rect 270 173 276 174
rect 230 168 236 169
rect 254 171 261 172
rect 110 166 116 167
rect 254 167 255 171
rect 260 167 261 171
rect 270 169 271 173
rect 275 169 276 173
rect 270 168 276 169
rect 310 173 316 174
rect 310 169 311 173
rect 315 169 316 173
rect 310 168 316 169
rect 350 173 356 174
rect 350 169 351 173
rect 355 169 356 173
rect 350 168 356 169
rect 390 173 396 174
rect 390 169 391 173
rect 395 169 396 173
rect 390 168 396 169
rect 686 171 692 172
rect 254 166 261 167
rect 415 167 421 168
rect 415 166 416 167
rect 319 164 416 166
rect 263 163 269 164
rect 263 159 264 163
rect 268 162 269 163
rect 319 162 321 164
rect 415 163 416 164
rect 420 163 421 167
rect 686 167 687 171
rect 691 167 692 171
rect 686 166 692 167
rect 415 162 421 163
rect 268 160 321 162
rect 268 159 269 160
rect 263 158 269 159
rect 198 135 204 136
rect 198 131 199 135
rect 203 134 204 135
rect 203 132 466 134
rect 203 131 204 132
rect 198 130 204 131
rect 464 130 466 132
rect 479 131 485 132
rect 479 130 480 131
rect 110 129 116 130
rect 110 125 111 129
rect 115 125 116 129
rect 464 128 480 130
rect 110 124 116 125
rect 134 127 140 128
rect 134 123 135 127
rect 139 123 140 127
rect 134 122 140 123
rect 174 127 180 128
rect 174 123 175 127
rect 179 123 180 127
rect 174 122 180 123
rect 214 127 220 128
rect 214 123 215 127
rect 219 123 220 127
rect 214 122 220 123
rect 254 127 260 128
rect 254 123 255 127
rect 259 123 260 127
rect 254 122 260 123
rect 294 127 300 128
rect 294 123 295 127
rect 299 123 300 127
rect 294 122 300 123
rect 334 127 340 128
rect 334 123 335 127
rect 339 123 340 127
rect 334 122 340 123
rect 374 127 380 128
rect 374 123 375 127
rect 379 123 380 127
rect 374 122 380 123
rect 414 127 420 128
rect 414 123 415 127
rect 419 123 420 127
rect 414 122 420 123
rect 454 127 460 128
rect 454 123 455 127
rect 459 123 460 127
rect 479 127 480 128
rect 484 127 485 131
rect 479 126 485 127
rect 686 129 692 130
rect 686 125 687 129
rect 691 125 692 129
rect 686 124 692 125
rect 454 122 460 123
rect 150 112 156 113
rect 190 112 196 113
rect 230 112 236 113
rect 270 112 276 113
rect 310 112 316 113
rect 350 112 356 113
rect 390 112 396 113
rect 430 112 436 113
rect 470 112 476 113
rect 110 111 116 112
rect 110 107 111 111
rect 115 107 116 111
rect 150 108 151 112
rect 155 108 156 112
rect 150 107 156 108
rect 159 111 165 112
rect 159 107 160 111
rect 164 110 165 111
rect 164 108 174 110
rect 164 107 165 108
rect 110 106 116 107
rect 159 106 165 107
rect 172 94 174 108
rect 190 108 191 112
rect 195 108 196 112
rect 190 107 196 108
rect 199 111 205 112
rect 199 107 200 111
rect 204 110 205 111
rect 204 108 214 110
rect 204 107 205 108
rect 199 106 205 107
rect 183 95 189 96
rect 183 94 184 95
rect 172 92 184 94
rect 183 91 184 92
rect 188 91 189 95
rect 212 94 214 108
rect 230 108 231 112
rect 235 108 236 112
rect 230 107 236 108
rect 239 111 245 112
rect 239 107 240 111
rect 244 110 245 111
rect 244 108 254 110
rect 244 107 245 108
rect 239 106 245 107
rect 223 95 229 96
rect 223 94 224 95
rect 212 92 224 94
rect 183 90 189 91
rect 223 91 224 92
rect 228 91 229 95
rect 252 94 254 108
rect 270 108 271 112
rect 275 108 276 112
rect 270 107 276 108
rect 279 111 285 112
rect 279 107 280 111
rect 284 110 285 111
rect 284 108 294 110
rect 284 107 285 108
rect 279 106 285 107
rect 263 95 269 96
rect 263 94 264 95
rect 252 92 264 94
rect 223 90 229 91
rect 263 91 264 92
rect 268 91 269 95
rect 292 94 294 108
rect 310 108 311 112
rect 315 108 316 112
rect 310 107 316 108
rect 319 111 325 112
rect 319 107 320 111
rect 324 110 325 111
rect 324 108 334 110
rect 324 107 325 108
rect 319 106 325 107
rect 303 95 309 96
rect 303 94 304 95
rect 292 92 304 94
rect 263 90 269 91
rect 303 91 304 92
rect 308 91 309 95
rect 332 94 334 108
rect 350 108 351 112
rect 355 108 356 112
rect 350 107 356 108
rect 359 111 365 112
rect 359 107 360 111
rect 364 110 365 111
rect 364 108 374 110
rect 364 107 365 108
rect 359 106 365 107
rect 343 95 349 96
rect 343 94 344 95
rect 332 92 344 94
rect 303 90 309 91
rect 343 91 344 92
rect 348 91 349 95
rect 372 94 374 108
rect 390 108 391 112
rect 395 108 396 112
rect 390 107 396 108
rect 399 111 405 112
rect 399 107 400 111
rect 404 110 405 111
rect 404 108 414 110
rect 404 107 405 108
rect 399 106 405 107
rect 383 95 389 96
rect 383 94 384 95
rect 372 92 384 94
rect 343 90 349 91
rect 383 91 384 92
rect 388 91 389 95
rect 412 94 414 108
rect 430 108 431 112
rect 435 108 436 112
rect 430 107 436 108
rect 439 111 445 112
rect 439 107 440 111
rect 444 110 445 111
rect 444 108 454 110
rect 444 107 445 108
rect 439 106 445 107
rect 423 95 429 96
rect 423 94 424 95
rect 412 92 424 94
rect 383 90 389 91
rect 423 91 424 92
rect 428 91 429 95
rect 452 94 454 108
rect 470 108 471 112
rect 475 108 476 112
rect 470 107 476 108
rect 686 111 692 112
rect 686 107 687 111
rect 691 107 692 111
rect 686 106 692 107
rect 463 95 469 96
rect 463 94 464 95
rect 452 92 464 94
rect 423 90 429 91
rect 463 91 464 92
rect 468 91 469 95
rect 463 90 469 91
<< m3c >>
rect 343 767 347 771
rect 375 769 376 773
rect 376 769 379 773
rect 455 769 459 773
rect 551 769 555 773
rect 663 769 667 773
rect 111 753 115 757
rect 295 752 299 756
rect 375 751 379 755
rect 383 752 387 756
rect 455 751 459 755
rect 479 752 483 756
rect 551 751 555 755
rect 575 752 579 756
rect 655 752 659 756
rect 687 753 691 757
rect 111 735 115 739
rect 279 737 283 741
rect 367 737 371 741
rect 463 737 467 741
rect 559 737 563 741
rect 639 737 643 741
rect 391 731 395 735
rect 687 735 691 739
rect 111 709 115 713
rect 199 707 203 711
rect 239 707 243 711
rect 279 707 283 711
rect 319 707 323 711
rect 343 711 344 715
rect 344 711 347 715
rect 359 707 363 711
rect 407 707 411 711
rect 463 707 467 711
rect 527 707 531 711
rect 591 707 595 711
rect 639 707 643 711
rect 663 711 664 715
rect 664 711 667 715
rect 687 709 691 713
rect 111 691 115 695
rect 215 692 219 696
rect 223 675 227 679
rect 255 692 259 696
rect 295 692 299 696
rect 335 692 339 696
rect 375 692 379 696
rect 391 675 395 679
rect 423 692 427 696
rect 479 692 483 696
rect 543 692 547 696
rect 551 691 552 695
rect 552 691 555 695
rect 607 692 611 696
rect 655 692 659 696
rect 687 691 691 695
rect 187 661 191 665
rect 207 661 211 665
rect 271 661 275 665
rect 359 661 360 665
rect 360 661 363 665
rect 503 663 507 667
rect 551 663 555 667
rect 631 659 635 663
rect 663 661 667 665
rect 111 645 115 649
rect 175 644 179 648
rect 207 643 211 647
rect 231 644 235 648
rect 271 643 275 647
rect 295 644 299 648
rect 359 643 363 647
rect 367 644 371 648
rect 439 644 443 648
rect 519 644 523 648
rect 599 644 603 648
rect 655 644 659 648
rect 687 645 691 649
rect 111 627 115 631
rect 159 629 163 633
rect 215 629 219 633
rect 279 629 283 633
rect 351 629 355 633
rect 423 629 427 633
rect 503 629 507 633
rect 583 629 587 633
rect 639 629 643 633
rect 223 623 227 627
rect 495 623 499 627
rect 511 623 515 627
rect 631 623 635 627
rect 687 627 691 631
rect 187 599 191 603
rect 111 593 115 597
rect 199 591 203 595
rect 263 599 267 603
rect 239 591 243 595
rect 295 591 299 595
rect 351 591 355 595
rect 415 591 419 595
rect 487 591 491 595
rect 567 591 571 595
rect 639 591 643 595
rect 663 595 664 599
rect 664 595 667 599
rect 687 593 691 597
rect 223 583 227 587
rect 403 583 407 587
rect 111 575 115 579
rect 215 576 219 580
rect 255 576 259 580
rect 311 576 315 580
rect 367 576 371 580
rect 431 576 435 580
rect 503 576 507 580
rect 223 559 227 563
rect 263 559 267 563
rect 403 559 407 563
rect 419 559 423 563
rect 495 559 496 563
rect 496 559 499 563
rect 583 576 587 580
rect 591 575 592 579
rect 592 575 595 579
rect 655 576 659 580
rect 687 575 691 579
rect 627 559 631 563
rect 339 545 343 549
rect 347 545 351 549
rect 387 545 391 549
rect 511 551 515 555
rect 535 543 539 547
rect 591 547 595 551
rect 607 545 608 549
rect 608 545 611 549
rect 663 545 667 549
rect 111 529 115 533
rect 327 528 331 532
rect 347 527 351 531
rect 367 528 371 532
rect 387 527 391 531
rect 407 528 411 532
rect 419 527 420 531
rect 420 527 423 531
rect 455 528 459 532
rect 503 528 507 532
rect 511 527 512 531
rect 512 527 515 531
rect 559 528 563 532
rect 615 528 619 532
rect 627 527 628 531
rect 628 527 631 531
rect 655 528 659 532
rect 687 529 691 533
rect 111 511 115 515
rect 311 513 315 517
rect 351 513 355 517
rect 391 513 395 517
rect 439 513 443 517
rect 487 513 491 517
rect 543 513 547 517
rect 599 513 603 517
rect 639 513 643 517
rect 339 507 343 511
rect 591 507 595 511
rect 607 507 611 511
rect 687 511 691 515
rect 111 485 115 489
rect 255 483 259 487
rect 295 483 299 487
rect 335 483 339 487
rect 391 483 395 487
rect 447 483 451 487
rect 511 483 515 487
rect 535 487 536 491
rect 536 487 539 491
rect 583 483 587 487
rect 639 483 643 487
rect 663 487 664 491
rect 664 487 667 491
rect 687 485 691 489
rect 111 467 115 471
rect 271 468 275 472
rect 311 468 315 472
rect 351 468 355 472
rect 407 468 411 472
rect 463 468 467 472
rect 527 468 531 472
rect 599 468 603 472
rect 607 467 608 471
rect 608 467 611 471
rect 655 468 659 472
rect 687 467 691 471
rect 591 451 592 455
rect 592 451 595 455
rect 663 451 667 455
rect 503 443 507 447
rect 183 437 187 441
rect 255 437 259 441
rect 335 437 336 441
rect 336 437 339 441
rect 391 437 395 441
rect 471 437 475 441
rect 607 439 611 443
rect 647 437 648 441
rect 648 437 651 441
rect 111 421 115 425
rect 175 420 179 424
rect 223 420 227 424
rect 255 419 259 423
rect 279 420 283 424
rect 335 419 339 423
rect 343 420 347 424
rect 391 419 395 423
rect 415 420 419 424
rect 471 419 475 423
rect 495 420 499 424
rect 503 419 504 423
rect 504 419 507 423
rect 583 420 587 424
rect 655 420 659 424
rect 663 419 664 423
rect 664 419 667 423
rect 687 421 691 425
rect 111 403 115 407
rect 159 405 163 409
rect 207 405 211 409
rect 263 405 267 409
rect 327 405 331 409
rect 399 405 403 409
rect 479 405 483 409
rect 567 405 571 409
rect 639 405 643 409
rect 547 399 551 403
rect 687 403 691 407
rect 183 379 187 383
rect 111 373 115 377
rect 135 371 139 375
rect 175 371 179 375
rect 215 371 219 375
rect 279 371 283 375
rect 647 379 651 383
rect 343 371 347 375
rect 415 371 419 375
rect 495 371 499 375
rect 575 371 579 375
rect 639 371 643 375
rect 687 373 691 377
rect 159 363 163 367
rect 303 363 307 367
rect 111 355 115 359
rect 151 356 155 360
rect 159 339 163 343
rect 191 356 195 360
rect 231 356 235 360
rect 295 356 299 360
rect 359 356 363 360
rect 303 339 307 343
rect 347 339 351 343
rect 431 356 435 360
rect 511 356 515 360
rect 519 355 520 359
rect 520 355 523 359
rect 591 356 595 360
rect 547 339 551 343
rect 607 339 611 343
rect 655 356 659 360
rect 687 355 691 359
rect 267 321 271 325
rect 275 321 279 325
rect 315 323 319 327
rect 439 327 443 331
rect 487 327 491 331
rect 471 321 472 325
rect 472 321 475 325
rect 519 321 520 325
rect 520 321 523 325
rect 627 321 631 325
rect 663 321 667 325
rect 111 305 115 309
rect 255 304 259 308
rect 275 303 279 307
rect 295 304 299 308
rect 315 303 319 307
rect 335 304 339 308
rect 347 303 348 307
rect 348 303 351 307
rect 383 304 387 308
rect 431 304 435 308
rect 439 303 440 307
rect 440 303 443 307
rect 479 304 483 308
rect 487 303 488 307
rect 488 303 491 307
rect 527 304 531 308
rect 575 304 579 308
rect 615 304 619 308
rect 655 304 659 308
rect 687 305 691 309
rect 111 287 115 291
rect 239 289 243 293
rect 279 289 283 293
rect 319 289 323 293
rect 367 289 371 293
rect 415 289 419 293
rect 463 289 467 293
rect 511 289 515 293
rect 559 289 563 293
rect 599 289 603 293
rect 627 291 631 295
rect 267 283 271 287
rect 503 283 507 287
rect 607 283 611 287
rect 639 289 643 293
rect 687 287 691 291
rect 111 261 115 265
rect 239 259 243 263
rect 279 259 283 263
rect 319 259 323 263
rect 359 259 363 263
rect 399 259 403 263
rect 439 259 443 263
rect 463 259 464 263
rect 464 259 467 263
rect 479 259 483 263
rect 519 259 523 263
rect 559 259 563 263
rect 599 259 603 263
rect 639 259 643 263
rect 663 263 664 267
rect 664 263 667 267
rect 687 261 691 265
rect 111 243 115 247
rect 255 244 259 248
rect 295 244 299 248
rect 335 244 339 248
rect 375 244 379 248
rect 415 244 419 248
rect 455 244 459 248
rect 495 244 499 248
rect 503 227 507 231
rect 535 244 539 248
rect 575 244 579 248
rect 615 244 619 248
rect 655 244 659 248
rect 687 243 691 247
rect 199 201 200 205
rect 200 201 203 205
rect 227 201 231 205
rect 263 201 267 205
rect 347 201 351 205
rect 387 201 391 205
rect 111 185 115 189
rect 207 184 211 188
rect 227 183 231 187
rect 247 184 251 188
rect 287 184 291 188
rect 327 184 331 188
rect 347 183 351 187
rect 367 184 371 188
rect 387 183 391 187
rect 407 184 411 188
rect 687 185 691 189
rect 111 167 115 171
rect 191 169 195 173
rect 231 169 235 173
rect 255 167 256 171
rect 256 167 259 171
rect 271 169 275 173
rect 311 169 315 173
rect 351 169 355 173
rect 391 169 395 173
rect 687 167 691 171
rect 199 131 203 135
rect 111 125 115 129
rect 135 123 139 127
rect 175 123 179 127
rect 215 123 219 127
rect 255 123 259 127
rect 295 123 299 127
rect 335 123 339 127
rect 375 123 379 127
rect 415 123 419 127
rect 455 123 459 127
rect 687 125 691 129
rect 111 107 115 111
rect 151 108 155 112
rect 191 108 195 112
rect 231 108 235 112
rect 271 108 275 112
rect 311 108 315 112
rect 351 108 355 112
rect 391 108 395 112
rect 431 108 435 112
rect 471 108 475 112
rect 687 107 691 111
<< m3 >>
rect 111 778 115 779
rect 111 773 115 774
rect 295 778 299 779
rect 383 778 387 779
rect 479 778 483 779
rect 575 778 579 779
rect 295 773 299 774
rect 374 773 380 774
rect 383 773 387 774
rect 454 773 460 774
rect 479 773 483 774
rect 550 773 556 774
rect 575 773 579 774
rect 655 778 659 779
rect 687 778 691 779
rect 655 773 659 774
rect 662 773 668 774
rect 687 773 691 774
rect 112 758 114 773
rect 110 757 116 758
rect 296 757 298 773
rect 342 771 348 772
rect 342 767 343 771
rect 347 767 348 771
rect 374 769 375 773
rect 379 769 380 773
rect 374 768 380 769
rect 342 766 348 767
rect 110 753 111 757
rect 115 753 116 757
rect 110 752 116 753
rect 294 756 300 757
rect 294 752 295 756
rect 299 752 300 756
rect 294 751 300 752
rect 278 741 284 742
rect 110 739 116 740
rect 110 735 111 739
rect 115 735 116 739
rect 278 737 279 741
rect 283 737 284 741
rect 278 736 284 737
rect 110 734 116 735
rect 112 727 114 734
rect 280 727 282 736
rect 111 726 115 727
rect 111 721 115 722
rect 199 726 203 727
rect 199 721 203 722
rect 239 726 243 727
rect 239 721 243 722
rect 279 726 283 727
rect 279 721 283 722
rect 319 726 323 727
rect 319 721 323 722
rect 112 714 114 721
rect 110 713 116 714
rect 110 709 111 713
rect 115 709 116 713
rect 200 712 202 721
rect 240 712 242 721
rect 280 712 282 721
rect 320 712 322 721
rect 344 716 346 766
rect 376 756 378 768
rect 384 757 386 773
rect 454 769 455 773
rect 459 769 460 773
rect 454 768 460 769
rect 382 756 388 757
rect 456 756 458 768
rect 480 757 482 773
rect 550 769 551 773
rect 555 769 556 773
rect 550 768 556 769
rect 478 756 484 757
rect 552 756 554 768
rect 576 757 578 773
rect 656 757 658 773
rect 662 769 663 773
rect 667 769 668 773
rect 662 768 668 769
rect 574 756 580 757
rect 374 755 380 756
rect 374 751 375 755
rect 379 751 380 755
rect 382 752 383 756
rect 387 752 388 756
rect 382 751 388 752
rect 454 755 460 756
rect 454 751 455 755
rect 459 751 460 755
rect 478 752 479 756
rect 483 752 484 756
rect 478 751 484 752
rect 550 755 556 756
rect 550 751 551 755
rect 555 751 556 755
rect 574 752 575 756
rect 579 752 580 756
rect 574 751 580 752
rect 654 756 660 757
rect 654 752 655 756
rect 659 752 660 756
rect 654 751 660 752
rect 374 750 380 751
rect 454 750 460 751
rect 550 750 556 751
rect 366 741 372 742
rect 366 737 367 741
rect 371 737 372 741
rect 366 736 372 737
rect 462 741 468 742
rect 462 737 463 741
rect 467 737 468 741
rect 462 736 468 737
rect 558 741 564 742
rect 558 737 559 741
rect 563 737 564 741
rect 558 736 564 737
rect 638 741 644 742
rect 638 737 639 741
rect 643 737 644 741
rect 638 736 644 737
rect 368 727 370 736
rect 390 735 396 736
rect 390 731 391 735
rect 395 731 396 735
rect 390 730 396 731
rect 359 726 363 727
rect 359 721 363 722
rect 367 726 371 727
rect 367 721 371 722
rect 342 715 348 716
rect 110 708 116 709
rect 198 711 204 712
rect 198 707 199 711
rect 203 707 204 711
rect 198 706 204 707
rect 238 711 244 712
rect 238 707 239 711
rect 243 707 244 711
rect 238 706 244 707
rect 278 711 284 712
rect 278 707 279 711
rect 283 707 284 711
rect 278 706 284 707
rect 318 711 324 712
rect 318 707 319 711
rect 323 707 324 711
rect 342 711 343 715
rect 347 711 348 715
rect 360 712 362 721
rect 342 710 348 711
rect 358 711 364 712
rect 318 706 324 707
rect 358 707 359 711
rect 363 707 364 711
rect 358 706 364 707
rect 214 696 220 697
rect 110 695 116 696
rect 110 691 111 695
rect 115 691 116 695
rect 214 692 215 696
rect 219 692 220 696
rect 214 691 220 692
rect 254 696 260 697
rect 254 692 255 696
rect 259 692 260 696
rect 254 691 260 692
rect 294 696 300 697
rect 294 692 295 696
rect 299 692 300 696
rect 294 691 300 692
rect 334 696 340 697
rect 334 692 335 696
rect 339 692 340 696
rect 334 691 340 692
rect 374 696 380 697
rect 374 692 375 696
rect 379 692 380 696
rect 374 691 380 692
rect 110 690 116 691
rect 112 671 114 690
rect 216 671 218 691
rect 222 679 228 680
rect 222 675 223 679
rect 227 675 228 679
rect 222 674 228 675
rect 111 670 115 671
rect 111 665 115 666
rect 175 670 179 671
rect 215 670 219 671
rect 175 665 179 666
rect 186 665 192 666
rect 112 650 114 665
rect 110 649 116 650
rect 176 649 178 665
rect 186 661 187 665
rect 191 661 192 665
rect 186 660 192 661
rect 206 665 212 666
rect 215 665 219 666
rect 206 661 207 665
rect 211 661 212 665
rect 206 660 212 661
rect 110 645 111 649
rect 115 645 116 649
rect 110 644 116 645
rect 174 648 180 649
rect 174 644 175 648
rect 179 644 180 648
rect 174 643 180 644
rect 158 633 164 634
rect 110 631 116 632
rect 110 627 111 631
rect 115 627 116 631
rect 158 629 159 633
rect 163 629 164 633
rect 158 628 164 629
rect 110 626 116 627
rect 112 611 114 626
rect 160 611 162 628
rect 111 610 115 611
rect 111 605 115 606
rect 159 610 163 611
rect 159 605 163 606
rect 112 598 114 605
rect 188 604 190 660
rect 208 648 210 660
rect 206 647 212 648
rect 206 643 207 647
rect 211 643 212 647
rect 206 642 212 643
rect 214 633 220 634
rect 214 629 215 633
rect 219 629 220 633
rect 214 628 220 629
rect 224 628 226 674
rect 256 671 258 691
rect 296 671 298 691
rect 336 671 338 691
rect 376 671 378 691
rect 392 680 394 730
rect 464 727 466 736
rect 560 727 562 736
rect 640 727 642 736
rect 407 726 411 727
rect 407 721 411 722
rect 463 726 467 727
rect 463 721 467 722
rect 527 726 531 727
rect 527 721 531 722
rect 559 726 563 727
rect 559 721 563 722
rect 591 726 595 727
rect 591 721 595 722
rect 639 726 643 727
rect 639 721 643 722
rect 408 712 410 721
rect 464 712 466 721
rect 528 712 530 721
rect 592 712 594 721
rect 640 712 642 721
rect 664 716 666 768
rect 688 758 690 773
rect 686 757 692 758
rect 686 753 687 757
rect 691 753 692 757
rect 686 752 692 753
rect 686 739 692 740
rect 686 735 687 739
rect 691 735 692 739
rect 686 734 692 735
rect 688 727 690 734
rect 687 726 691 727
rect 687 721 691 722
rect 662 715 668 716
rect 406 711 412 712
rect 406 707 407 711
rect 411 707 412 711
rect 406 706 412 707
rect 462 711 468 712
rect 462 707 463 711
rect 467 707 468 711
rect 462 706 468 707
rect 526 711 532 712
rect 526 707 527 711
rect 531 707 532 711
rect 526 706 532 707
rect 590 711 596 712
rect 590 707 591 711
rect 595 707 596 711
rect 590 706 596 707
rect 638 711 644 712
rect 638 707 639 711
rect 643 707 644 711
rect 662 711 663 715
rect 667 711 668 715
rect 688 714 690 721
rect 662 710 668 711
rect 686 713 692 714
rect 686 709 687 713
rect 691 709 692 713
rect 686 708 692 709
rect 638 706 644 707
rect 422 696 428 697
rect 422 692 423 696
rect 427 692 428 696
rect 422 691 428 692
rect 478 696 484 697
rect 478 692 479 696
rect 483 692 484 696
rect 478 691 484 692
rect 542 696 548 697
rect 606 696 612 697
rect 542 692 543 696
rect 547 692 548 696
rect 542 691 548 692
rect 550 695 556 696
rect 550 691 551 695
rect 555 691 556 695
rect 606 692 607 696
rect 611 692 612 696
rect 606 691 612 692
rect 654 696 660 697
rect 654 692 655 696
rect 659 692 660 696
rect 654 691 660 692
rect 686 695 692 696
rect 686 691 687 695
rect 691 691 692 695
rect 390 679 396 680
rect 390 675 391 679
rect 395 675 396 679
rect 390 674 396 675
rect 424 671 426 691
rect 480 671 482 691
rect 544 671 546 691
rect 550 690 556 691
rect 231 670 235 671
rect 231 665 235 666
rect 255 670 259 671
rect 295 670 299 671
rect 255 665 259 666
rect 270 665 276 666
rect 295 665 299 666
rect 335 670 339 671
rect 367 670 371 671
rect 335 665 339 666
rect 358 665 364 666
rect 367 665 371 666
rect 375 670 379 671
rect 375 665 379 666
rect 423 670 427 671
rect 423 665 427 666
rect 439 670 443 671
rect 439 665 443 666
rect 479 670 483 671
rect 519 670 523 671
rect 479 665 483 666
rect 502 667 508 668
rect 232 649 234 665
rect 270 661 271 665
rect 275 661 276 665
rect 270 660 276 661
rect 230 648 236 649
rect 272 648 274 660
rect 296 649 298 665
rect 358 661 359 665
rect 363 661 364 665
rect 358 660 364 661
rect 294 648 300 649
rect 360 648 362 660
rect 368 649 370 665
rect 440 649 442 665
rect 502 663 503 667
rect 507 663 508 667
rect 519 665 523 666
rect 543 670 547 671
rect 552 668 554 690
rect 608 671 610 691
rect 656 671 658 691
rect 686 690 692 691
rect 688 671 690 690
rect 599 670 603 671
rect 543 665 547 666
rect 550 667 556 668
rect 502 662 508 663
rect 504 651 506 662
rect 504 649 514 651
rect 520 649 522 665
rect 550 663 551 667
rect 555 663 556 667
rect 599 665 603 666
rect 607 670 611 671
rect 607 665 611 666
rect 655 670 659 671
rect 687 670 691 671
rect 655 665 659 666
rect 662 665 668 666
rect 687 665 691 666
rect 550 662 556 663
rect 600 649 602 665
rect 630 663 636 664
rect 630 659 631 663
rect 635 659 636 663
rect 630 658 636 659
rect 366 648 372 649
rect 230 644 231 648
rect 235 644 236 648
rect 230 643 236 644
rect 270 647 276 648
rect 270 643 271 647
rect 275 643 276 647
rect 294 644 295 648
rect 299 644 300 648
rect 294 643 300 644
rect 358 647 364 648
rect 358 643 359 647
rect 363 643 364 647
rect 366 644 367 648
rect 371 644 372 648
rect 366 643 372 644
rect 438 648 444 649
rect 438 644 439 648
rect 443 644 444 648
rect 438 643 444 644
rect 270 642 276 643
rect 358 642 364 643
rect 278 633 284 634
rect 278 629 279 633
rect 283 629 284 633
rect 278 628 284 629
rect 350 633 356 634
rect 350 629 351 633
rect 355 629 356 633
rect 350 628 356 629
rect 422 633 428 634
rect 422 629 423 633
rect 427 629 428 633
rect 422 628 428 629
rect 502 633 508 634
rect 502 629 503 633
rect 507 629 508 633
rect 502 628 508 629
rect 512 628 514 649
rect 518 648 524 649
rect 518 644 519 648
rect 523 644 524 648
rect 518 643 524 644
rect 598 648 604 649
rect 598 644 599 648
rect 603 644 604 648
rect 598 643 604 644
rect 582 633 588 634
rect 582 629 583 633
rect 587 629 588 633
rect 582 628 588 629
rect 632 628 634 658
rect 656 649 658 665
rect 662 661 663 665
rect 667 661 668 665
rect 662 660 668 661
rect 654 648 660 649
rect 654 644 655 648
rect 659 644 660 648
rect 654 643 660 644
rect 638 633 644 634
rect 638 629 639 633
rect 643 629 644 633
rect 638 628 644 629
rect 216 611 218 628
rect 222 627 228 628
rect 222 623 223 627
rect 227 623 228 627
rect 222 622 228 623
rect 280 611 282 628
rect 352 611 354 628
rect 424 611 426 628
rect 494 627 500 628
rect 494 623 495 627
rect 499 623 500 627
rect 494 622 500 623
rect 199 610 203 611
rect 199 605 203 606
rect 215 610 219 611
rect 215 605 219 606
rect 239 610 243 611
rect 239 605 243 606
rect 279 610 283 611
rect 279 605 283 606
rect 295 610 299 611
rect 295 605 299 606
rect 351 610 355 611
rect 351 605 355 606
rect 415 610 419 611
rect 415 605 419 606
rect 423 610 427 611
rect 423 605 427 606
rect 487 610 491 611
rect 487 605 491 606
rect 186 603 192 604
rect 186 599 187 603
rect 191 599 192 603
rect 186 598 192 599
rect 110 597 116 598
rect 110 593 111 597
rect 115 593 116 597
rect 200 596 202 605
rect 240 596 242 605
rect 262 603 268 604
rect 262 599 263 603
rect 267 599 268 603
rect 262 598 268 599
rect 110 592 116 593
rect 198 595 204 596
rect 198 591 199 595
rect 203 591 204 595
rect 198 590 204 591
rect 238 595 244 596
rect 238 591 239 595
rect 243 591 244 595
rect 238 590 244 591
rect 222 587 228 588
rect 222 583 223 587
rect 227 583 228 587
rect 222 582 228 583
rect 214 580 220 581
rect 110 579 116 580
rect 110 575 111 579
rect 115 575 116 579
rect 214 576 215 580
rect 219 576 220 580
rect 214 575 220 576
rect 110 574 116 575
rect 112 555 114 574
rect 216 555 218 575
rect 224 564 226 582
rect 254 580 260 581
rect 254 576 255 580
rect 259 576 260 580
rect 254 575 260 576
rect 222 563 228 564
rect 222 559 223 563
rect 227 559 228 563
rect 222 558 228 559
rect 256 555 258 575
rect 264 564 266 598
rect 296 596 298 605
rect 352 596 354 605
rect 416 596 418 605
rect 488 596 490 605
rect 294 595 300 596
rect 294 591 295 595
rect 299 591 300 595
rect 294 590 300 591
rect 350 595 356 596
rect 350 591 351 595
rect 355 591 356 595
rect 350 590 356 591
rect 414 595 420 596
rect 414 591 415 595
rect 419 591 420 595
rect 414 590 420 591
rect 486 595 492 596
rect 486 591 487 595
rect 491 591 492 595
rect 486 590 492 591
rect 402 587 408 588
rect 402 583 403 587
rect 407 583 408 587
rect 402 582 408 583
rect 310 580 316 581
rect 310 576 311 580
rect 315 576 316 580
rect 310 575 316 576
rect 366 580 372 581
rect 366 576 367 580
rect 371 576 372 580
rect 366 575 372 576
rect 262 563 268 564
rect 262 559 263 563
rect 267 559 268 563
rect 262 558 268 559
rect 312 555 314 575
rect 368 555 370 575
rect 404 564 406 582
rect 430 580 436 581
rect 430 576 431 580
rect 435 576 436 580
rect 430 575 436 576
rect 402 563 408 564
rect 402 559 403 563
rect 407 559 408 563
rect 402 558 408 559
rect 418 563 424 564
rect 418 559 419 563
rect 423 559 424 563
rect 418 558 424 559
rect 111 554 115 555
rect 111 549 115 550
rect 215 554 219 555
rect 215 549 219 550
rect 255 554 259 555
rect 255 549 259 550
rect 311 554 315 555
rect 311 549 315 550
rect 327 554 331 555
rect 367 554 371 555
rect 407 554 411 555
rect 327 549 331 550
rect 338 549 344 550
rect 112 534 114 549
rect 110 533 116 534
rect 328 533 330 549
rect 338 545 339 549
rect 343 545 344 549
rect 338 544 344 545
rect 346 549 352 550
rect 367 549 371 550
rect 386 549 392 550
rect 407 549 411 550
rect 346 545 347 549
rect 351 545 352 549
rect 346 544 352 545
rect 110 529 111 533
rect 115 529 116 533
rect 110 528 116 529
rect 326 532 332 533
rect 326 528 327 532
rect 331 528 332 532
rect 326 527 332 528
rect 310 517 316 518
rect 110 515 116 516
rect 110 511 111 515
rect 115 511 116 515
rect 310 513 311 517
rect 315 513 316 517
rect 310 512 316 513
rect 340 512 342 544
rect 348 532 350 544
rect 368 533 370 549
rect 386 545 387 549
rect 391 545 392 549
rect 386 544 392 545
rect 366 532 372 533
rect 388 532 390 544
rect 408 533 410 549
rect 406 532 412 533
rect 420 532 422 558
rect 432 555 434 575
rect 496 564 498 622
rect 504 611 506 628
rect 510 627 516 628
rect 510 623 511 627
rect 515 623 516 627
rect 510 622 516 623
rect 584 611 586 628
rect 630 627 636 628
rect 630 623 631 627
rect 635 623 636 627
rect 630 622 636 623
rect 640 611 642 628
rect 503 610 507 611
rect 503 605 507 606
rect 567 610 571 611
rect 567 605 571 606
rect 583 610 587 611
rect 583 605 587 606
rect 639 610 643 611
rect 639 605 643 606
rect 568 596 570 605
rect 640 596 642 605
rect 664 600 666 660
rect 688 650 690 665
rect 686 649 692 650
rect 686 645 687 649
rect 691 645 692 649
rect 686 644 692 645
rect 686 631 692 632
rect 686 627 687 631
rect 691 627 692 631
rect 686 626 692 627
rect 688 611 690 626
rect 687 610 691 611
rect 687 605 691 606
rect 662 599 668 600
rect 566 595 572 596
rect 566 591 567 595
rect 571 591 572 595
rect 566 590 572 591
rect 638 595 644 596
rect 638 591 639 595
rect 643 591 644 595
rect 662 595 663 599
rect 667 595 668 599
rect 688 598 690 605
rect 662 594 668 595
rect 686 597 692 598
rect 686 593 687 597
rect 691 593 692 597
rect 686 592 692 593
rect 638 590 644 591
rect 502 580 508 581
rect 502 576 503 580
rect 507 576 508 580
rect 502 575 508 576
rect 582 580 588 581
rect 654 580 660 581
rect 582 576 583 580
rect 587 576 588 580
rect 582 575 588 576
rect 590 579 596 580
rect 590 575 591 579
rect 595 575 596 579
rect 654 576 655 580
rect 659 576 660 580
rect 654 575 660 576
rect 686 579 692 580
rect 686 575 687 579
rect 691 575 692 579
rect 494 563 500 564
rect 494 559 495 563
rect 499 559 500 563
rect 494 558 500 559
rect 504 555 506 575
rect 510 555 516 556
rect 584 555 586 575
rect 590 574 596 575
rect 431 554 435 555
rect 431 549 435 550
rect 455 554 459 555
rect 455 549 459 550
rect 503 554 507 555
rect 510 551 511 555
rect 515 551 516 555
rect 510 550 516 551
rect 559 554 563 555
rect 503 549 507 550
rect 456 533 458 549
rect 504 533 506 549
rect 454 532 460 533
rect 346 531 352 532
rect 346 527 347 531
rect 351 527 352 531
rect 366 528 367 532
rect 371 528 372 532
rect 366 527 372 528
rect 386 531 392 532
rect 386 527 387 531
rect 391 527 392 531
rect 406 528 407 532
rect 411 528 412 532
rect 406 527 412 528
rect 418 531 424 532
rect 418 527 419 531
rect 423 527 424 531
rect 454 528 455 532
rect 459 528 460 532
rect 454 527 460 528
rect 502 532 508 533
rect 512 532 514 550
rect 559 549 563 550
rect 583 554 587 555
rect 592 552 594 574
rect 626 563 632 564
rect 626 559 627 563
rect 631 559 632 563
rect 626 558 632 559
rect 615 554 619 555
rect 583 549 587 550
rect 590 551 596 552
rect 534 547 540 548
rect 534 543 535 547
rect 539 543 540 547
rect 534 542 540 543
rect 502 528 503 532
rect 507 528 508 532
rect 502 527 508 528
rect 510 531 516 532
rect 510 527 511 531
rect 515 527 516 531
rect 346 526 352 527
rect 386 526 392 527
rect 418 526 424 527
rect 510 526 516 527
rect 350 517 356 518
rect 350 513 351 517
rect 355 513 356 517
rect 350 512 356 513
rect 390 517 396 518
rect 390 513 391 517
rect 395 513 396 517
rect 390 512 396 513
rect 438 517 444 518
rect 438 513 439 517
rect 443 513 444 517
rect 438 512 444 513
rect 486 517 492 518
rect 486 513 487 517
rect 491 513 492 517
rect 486 512 492 513
rect 110 510 116 511
rect 112 503 114 510
rect 312 503 314 512
rect 338 511 344 512
rect 338 507 339 511
rect 343 507 344 511
rect 338 506 344 507
rect 352 503 354 512
rect 392 503 394 512
rect 440 503 442 512
rect 488 503 490 512
rect 111 502 115 503
rect 111 497 115 498
rect 255 502 259 503
rect 255 497 259 498
rect 295 502 299 503
rect 295 497 299 498
rect 311 502 315 503
rect 311 497 315 498
rect 335 502 339 503
rect 335 497 339 498
rect 351 502 355 503
rect 351 497 355 498
rect 391 502 395 503
rect 391 497 395 498
rect 439 502 443 503
rect 439 497 443 498
rect 447 502 451 503
rect 447 497 451 498
rect 487 502 491 503
rect 487 497 491 498
rect 511 502 515 503
rect 511 497 515 498
rect 112 490 114 497
rect 110 489 116 490
rect 110 485 111 489
rect 115 485 116 489
rect 256 488 258 497
rect 296 488 298 497
rect 336 488 338 497
rect 392 488 394 497
rect 448 488 450 497
rect 512 488 514 497
rect 536 492 538 542
rect 560 533 562 549
rect 590 547 591 551
rect 595 547 596 551
rect 590 546 596 547
rect 606 549 612 550
rect 615 549 619 550
rect 606 545 607 549
rect 611 545 612 549
rect 606 544 612 545
rect 558 532 564 533
rect 558 528 559 532
rect 563 528 564 532
rect 558 527 564 528
rect 542 517 548 518
rect 542 513 543 517
rect 547 513 548 517
rect 542 512 548 513
rect 598 517 604 518
rect 598 513 599 517
rect 603 513 604 517
rect 598 512 604 513
rect 608 512 610 544
rect 616 533 618 549
rect 614 532 620 533
rect 628 532 630 558
rect 656 555 658 575
rect 686 574 692 575
rect 688 555 690 574
rect 655 554 659 555
rect 687 554 691 555
rect 655 549 659 550
rect 662 549 668 550
rect 687 549 691 550
rect 656 533 658 549
rect 662 545 663 549
rect 667 545 668 549
rect 662 544 668 545
rect 654 532 660 533
rect 614 528 615 532
rect 619 528 620 532
rect 614 527 620 528
rect 626 531 632 532
rect 626 527 627 531
rect 631 527 632 531
rect 654 528 655 532
rect 659 528 660 532
rect 654 527 660 528
rect 626 526 632 527
rect 638 517 644 518
rect 638 513 639 517
rect 643 513 644 517
rect 638 512 644 513
rect 544 503 546 512
rect 590 511 596 512
rect 590 507 591 511
rect 595 507 596 511
rect 590 506 596 507
rect 543 502 547 503
rect 543 497 547 498
rect 583 502 587 503
rect 583 497 587 498
rect 534 491 540 492
rect 110 484 116 485
rect 254 487 260 488
rect 254 483 255 487
rect 259 483 260 487
rect 254 482 260 483
rect 294 487 300 488
rect 294 483 295 487
rect 299 483 300 487
rect 294 482 300 483
rect 334 487 340 488
rect 334 483 335 487
rect 339 483 340 487
rect 334 482 340 483
rect 390 487 396 488
rect 390 483 391 487
rect 395 483 396 487
rect 390 482 396 483
rect 446 487 452 488
rect 446 483 447 487
rect 451 483 452 487
rect 446 482 452 483
rect 510 487 516 488
rect 510 483 511 487
rect 515 483 516 487
rect 534 487 535 491
rect 539 487 540 491
rect 584 488 586 497
rect 534 486 540 487
rect 582 487 588 488
rect 510 482 516 483
rect 582 483 583 487
rect 587 483 588 487
rect 582 482 588 483
rect 270 472 276 473
rect 110 471 116 472
rect 110 467 111 471
rect 115 467 116 471
rect 270 468 271 472
rect 275 468 276 472
rect 270 467 276 468
rect 310 472 316 473
rect 310 468 311 472
rect 315 468 316 472
rect 310 467 316 468
rect 350 472 356 473
rect 350 468 351 472
rect 355 468 356 472
rect 350 467 356 468
rect 406 472 412 473
rect 406 468 407 472
rect 411 468 412 472
rect 406 467 412 468
rect 462 472 468 473
rect 462 468 463 472
rect 467 468 468 472
rect 462 467 468 468
rect 526 472 532 473
rect 526 468 527 472
rect 531 468 532 472
rect 526 467 532 468
rect 110 466 116 467
rect 112 447 114 466
rect 272 447 274 467
rect 312 447 314 467
rect 352 447 354 467
rect 408 447 410 467
rect 464 447 466 467
rect 502 447 508 448
rect 528 447 530 467
rect 592 456 594 506
rect 600 503 602 512
rect 606 511 612 512
rect 606 507 607 511
rect 611 507 612 511
rect 606 506 612 507
rect 640 503 642 512
rect 599 502 603 503
rect 599 497 603 498
rect 639 502 643 503
rect 639 497 643 498
rect 640 488 642 497
rect 664 492 666 544
rect 688 534 690 549
rect 686 533 692 534
rect 686 529 687 533
rect 691 529 692 533
rect 686 528 692 529
rect 686 515 692 516
rect 686 511 687 515
rect 691 511 692 515
rect 686 510 692 511
rect 688 503 690 510
rect 687 502 691 503
rect 687 497 691 498
rect 662 491 668 492
rect 638 487 644 488
rect 638 483 639 487
rect 643 483 644 487
rect 662 487 663 491
rect 667 487 668 491
rect 688 490 690 497
rect 662 486 668 487
rect 686 489 692 490
rect 686 485 687 489
rect 691 485 692 489
rect 686 484 692 485
rect 638 482 644 483
rect 598 472 604 473
rect 654 472 660 473
rect 598 468 599 472
rect 603 468 604 472
rect 598 467 604 468
rect 606 471 612 472
rect 606 467 607 471
rect 611 467 612 471
rect 654 468 655 472
rect 659 468 660 472
rect 654 467 660 468
rect 686 471 692 472
rect 686 467 687 471
rect 691 467 692 471
rect 590 455 596 456
rect 590 451 591 455
rect 595 451 596 455
rect 590 450 596 451
rect 600 447 602 467
rect 606 466 612 467
rect 111 446 115 447
rect 111 441 115 442
rect 175 446 179 447
rect 223 446 227 447
rect 271 446 275 447
rect 175 441 179 442
rect 182 441 188 442
rect 223 441 227 442
rect 254 441 260 442
rect 271 441 275 442
rect 279 446 283 447
rect 279 441 283 442
rect 311 446 315 447
rect 343 446 347 447
rect 311 441 315 442
rect 334 441 340 442
rect 343 441 347 442
rect 351 446 355 447
rect 407 446 411 447
rect 351 441 355 442
rect 390 441 396 442
rect 407 441 411 442
rect 415 446 419 447
rect 415 441 419 442
rect 463 446 467 447
rect 495 446 499 447
rect 502 443 503 447
rect 507 443 508 447
rect 502 442 508 443
rect 527 446 531 447
rect 463 441 467 442
rect 470 441 476 442
rect 495 441 499 442
rect 112 426 114 441
rect 110 425 116 426
rect 176 425 178 441
rect 182 437 183 441
rect 187 437 188 441
rect 182 436 188 437
rect 110 421 111 425
rect 115 421 116 425
rect 110 420 116 421
rect 174 424 180 425
rect 174 420 175 424
rect 179 420 180 424
rect 174 419 180 420
rect 158 409 164 410
rect 110 407 116 408
rect 110 403 111 407
rect 115 403 116 407
rect 158 405 159 409
rect 163 405 164 409
rect 158 404 164 405
rect 110 402 116 403
rect 112 391 114 402
rect 160 391 162 404
rect 111 390 115 391
rect 111 385 115 386
rect 135 390 139 391
rect 135 385 139 386
rect 159 390 163 391
rect 159 385 163 386
rect 175 390 179 391
rect 175 385 179 386
rect 112 378 114 385
rect 110 377 116 378
rect 110 373 111 377
rect 115 373 116 377
rect 136 376 138 385
rect 176 376 178 385
rect 184 384 186 436
rect 224 425 226 441
rect 254 437 255 441
rect 259 437 260 441
rect 254 436 260 437
rect 222 424 228 425
rect 256 424 258 436
rect 280 425 282 441
rect 334 437 335 441
rect 339 437 340 441
rect 334 436 340 437
rect 278 424 284 425
rect 336 424 338 436
rect 344 425 346 441
rect 390 437 391 441
rect 395 437 396 441
rect 390 436 396 437
rect 342 424 348 425
rect 392 424 394 436
rect 416 425 418 441
rect 470 437 471 441
rect 475 437 476 441
rect 470 436 476 437
rect 414 424 420 425
rect 472 424 474 436
rect 496 425 498 441
rect 494 424 500 425
rect 504 424 506 442
rect 527 441 531 442
rect 583 446 587 447
rect 583 441 587 442
rect 599 446 603 447
rect 608 444 610 466
rect 656 447 658 467
rect 686 466 692 467
rect 662 455 668 456
rect 662 451 663 455
rect 667 451 668 455
rect 662 450 668 451
rect 655 446 659 447
rect 599 441 603 442
rect 606 443 612 444
rect 584 425 586 441
rect 606 439 607 443
rect 611 439 612 443
rect 606 438 612 439
rect 646 441 652 442
rect 655 441 659 442
rect 646 437 647 441
rect 651 437 652 441
rect 646 436 652 437
rect 582 424 588 425
rect 222 420 223 424
rect 227 420 228 424
rect 222 419 228 420
rect 254 423 260 424
rect 254 419 255 423
rect 259 419 260 423
rect 278 420 279 424
rect 283 420 284 424
rect 278 419 284 420
rect 334 423 340 424
rect 334 419 335 423
rect 339 419 340 423
rect 342 420 343 424
rect 347 420 348 424
rect 342 419 348 420
rect 390 423 396 424
rect 390 419 391 423
rect 395 419 396 423
rect 414 420 415 424
rect 419 420 420 424
rect 414 419 420 420
rect 470 423 476 424
rect 470 419 471 423
rect 475 419 476 423
rect 494 420 495 424
rect 499 420 500 424
rect 494 419 500 420
rect 502 423 508 424
rect 502 419 503 423
rect 507 419 508 423
rect 582 420 583 424
rect 587 420 588 424
rect 582 419 588 420
rect 254 418 260 419
rect 334 418 340 419
rect 390 418 396 419
rect 470 418 476 419
rect 502 418 508 419
rect 206 409 212 410
rect 206 405 207 409
rect 211 405 212 409
rect 206 404 212 405
rect 262 409 268 410
rect 262 405 263 409
rect 267 405 268 409
rect 262 404 268 405
rect 326 409 332 410
rect 326 405 327 409
rect 331 405 332 409
rect 326 404 332 405
rect 398 409 404 410
rect 398 405 399 409
rect 403 405 404 409
rect 398 404 404 405
rect 478 409 484 410
rect 478 405 479 409
rect 483 405 484 409
rect 478 404 484 405
rect 566 409 572 410
rect 566 405 567 409
rect 571 405 572 409
rect 566 404 572 405
rect 638 409 644 410
rect 638 405 639 409
rect 643 405 644 409
rect 638 404 644 405
rect 208 391 210 404
rect 264 391 266 404
rect 328 391 330 404
rect 400 391 402 404
rect 480 391 482 404
rect 546 403 552 404
rect 546 399 547 403
rect 551 399 552 403
rect 546 398 552 399
rect 207 390 211 391
rect 207 385 211 386
rect 215 390 219 391
rect 215 385 219 386
rect 263 390 267 391
rect 263 385 267 386
rect 279 390 283 391
rect 279 385 283 386
rect 327 390 331 391
rect 327 385 331 386
rect 343 390 347 391
rect 343 385 347 386
rect 399 390 403 391
rect 399 385 403 386
rect 415 390 419 391
rect 415 385 419 386
rect 479 390 483 391
rect 479 385 483 386
rect 495 390 499 391
rect 495 385 499 386
rect 182 383 188 384
rect 182 379 183 383
rect 187 379 188 383
rect 182 378 188 379
rect 216 376 218 385
rect 280 376 282 385
rect 344 376 346 385
rect 416 376 418 385
rect 496 376 498 385
rect 110 372 116 373
rect 134 375 140 376
rect 134 371 135 375
rect 139 371 140 375
rect 134 370 140 371
rect 174 375 180 376
rect 174 371 175 375
rect 179 371 180 375
rect 174 370 180 371
rect 214 375 220 376
rect 214 371 215 375
rect 219 371 220 375
rect 214 370 220 371
rect 278 375 284 376
rect 278 371 279 375
rect 283 371 284 375
rect 278 370 284 371
rect 342 375 348 376
rect 342 371 343 375
rect 347 371 348 375
rect 342 370 348 371
rect 414 375 420 376
rect 414 371 415 375
rect 419 371 420 375
rect 414 370 420 371
rect 494 375 500 376
rect 494 371 495 375
rect 499 371 500 375
rect 494 370 500 371
rect 158 367 164 368
rect 158 363 159 367
rect 163 363 164 367
rect 158 362 164 363
rect 302 367 308 368
rect 302 363 303 367
rect 307 363 308 367
rect 302 362 308 363
rect 150 360 156 361
rect 110 359 116 360
rect 110 355 111 359
rect 115 355 116 359
rect 150 356 151 360
rect 155 356 156 360
rect 150 355 156 356
rect 110 354 116 355
rect 112 331 114 354
rect 152 331 154 355
rect 160 344 162 362
rect 190 360 196 361
rect 190 356 191 360
rect 195 356 196 360
rect 190 355 196 356
rect 230 360 236 361
rect 230 356 231 360
rect 235 356 236 360
rect 230 355 236 356
rect 294 360 300 361
rect 294 356 295 360
rect 299 356 300 360
rect 294 355 300 356
rect 158 343 164 344
rect 158 339 159 343
rect 163 339 164 343
rect 158 338 164 339
rect 192 331 194 355
rect 232 331 234 355
rect 296 331 298 355
rect 304 344 306 362
rect 358 360 364 361
rect 358 356 359 360
rect 363 356 364 360
rect 358 355 364 356
rect 430 360 436 361
rect 430 356 431 360
rect 435 356 436 360
rect 430 355 436 356
rect 510 360 516 361
rect 510 356 511 360
rect 515 356 516 360
rect 510 355 516 356
rect 518 359 524 360
rect 518 355 519 359
rect 523 355 524 359
rect 302 343 308 344
rect 302 339 303 343
rect 307 339 308 343
rect 302 338 308 339
rect 346 343 352 344
rect 346 339 347 343
rect 351 339 352 343
rect 346 338 352 339
rect 111 330 115 331
rect 111 325 115 326
rect 151 330 155 331
rect 151 325 155 326
rect 191 330 195 331
rect 191 325 195 326
rect 231 330 235 331
rect 231 325 235 326
rect 255 330 259 331
rect 295 330 299 331
rect 335 330 339 331
rect 255 325 259 326
rect 266 325 272 326
rect 112 310 114 325
rect 110 309 116 310
rect 256 309 258 325
rect 266 321 267 325
rect 271 321 272 325
rect 266 320 272 321
rect 274 325 280 326
rect 295 325 299 326
rect 314 327 320 328
rect 274 321 275 325
rect 279 321 280 325
rect 274 320 280 321
rect 110 305 111 309
rect 115 305 116 309
rect 110 304 116 305
rect 254 308 260 309
rect 254 304 255 308
rect 259 304 260 308
rect 254 303 260 304
rect 238 293 244 294
rect 110 291 116 292
rect 110 287 111 291
rect 115 287 116 291
rect 238 289 239 293
rect 243 289 244 293
rect 238 288 244 289
rect 268 288 270 320
rect 276 308 278 320
rect 296 309 298 325
rect 314 323 315 327
rect 319 323 320 327
rect 335 325 339 326
rect 314 322 320 323
rect 294 308 300 309
rect 316 308 318 322
rect 336 309 338 325
rect 334 308 340 309
rect 348 308 350 338
rect 360 331 362 355
rect 432 331 434 355
rect 438 331 444 332
rect 486 331 492 332
rect 512 331 514 355
rect 518 354 524 355
rect 359 330 363 331
rect 359 325 363 326
rect 383 330 387 331
rect 383 325 387 326
rect 431 330 435 331
rect 438 327 439 331
rect 443 327 444 331
rect 438 326 444 327
rect 479 330 483 331
rect 486 327 487 331
rect 491 327 492 331
rect 486 326 492 327
rect 511 330 515 331
rect 520 326 522 354
rect 548 344 550 398
rect 568 391 570 404
rect 640 391 642 404
rect 567 390 571 391
rect 567 385 571 386
rect 575 390 579 391
rect 575 385 579 386
rect 639 390 643 391
rect 639 385 643 386
rect 576 376 578 385
rect 640 376 642 385
rect 648 384 650 436
rect 656 425 658 441
rect 654 424 660 425
rect 664 424 666 450
rect 688 447 690 466
rect 687 446 691 447
rect 687 441 691 442
rect 688 426 690 441
rect 686 425 692 426
rect 654 420 655 424
rect 659 420 660 424
rect 654 419 660 420
rect 662 423 668 424
rect 662 419 663 423
rect 667 419 668 423
rect 686 421 687 425
rect 691 421 692 425
rect 686 420 692 421
rect 662 418 668 419
rect 686 407 692 408
rect 686 403 687 407
rect 691 403 692 407
rect 686 402 692 403
rect 688 391 690 402
rect 687 390 691 391
rect 687 385 691 386
rect 646 383 652 384
rect 646 379 647 383
rect 651 379 652 383
rect 646 378 652 379
rect 688 378 690 385
rect 686 377 692 378
rect 574 375 580 376
rect 574 371 575 375
rect 579 371 580 375
rect 574 370 580 371
rect 638 375 644 376
rect 638 371 639 375
rect 643 371 644 375
rect 686 373 687 377
rect 691 373 692 377
rect 686 372 692 373
rect 638 370 644 371
rect 590 360 596 361
rect 590 356 591 360
rect 595 356 596 360
rect 590 355 596 356
rect 654 360 660 361
rect 654 356 655 360
rect 659 356 660 360
rect 654 355 660 356
rect 686 359 692 360
rect 686 355 687 359
rect 691 355 692 359
rect 546 343 552 344
rect 546 339 547 343
rect 551 339 552 343
rect 546 338 552 339
rect 592 331 594 355
rect 606 343 612 344
rect 606 339 607 343
rect 611 339 612 343
rect 606 338 612 339
rect 527 330 531 331
rect 431 325 435 326
rect 384 309 386 325
rect 432 309 434 325
rect 382 308 388 309
rect 274 307 280 308
rect 274 303 275 307
rect 279 303 280 307
rect 294 304 295 308
rect 299 304 300 308
rect 294 303 300 304
rect 314 307 320 308
rect 314 303 315 307
rect 319 303 320 307
rect 334 304 335 308
rect 339 304 340 308
rect 334 303 340 304
rect 346 307 352 308
rect 346 303 347 307
rect 351 303 352 307
rect 382 304 383 308
rect 387 304 388 308
rect 382 303 388 304
rect 430 308 436 309
rect 440 308 442 326
rect 470 325 476 326
rect 479 325 483 326
rect 470 321 471 325
rect 475 321 476 325
rect 470 320 476 321
rect 430 304 431 308
rect 435 304 436 308
rect 430 303 436 304
rect 438 307 444 308
rect 438 303 439 307
rect 443 303 444 307
rect 274 302 280 303
rect 314 302 320 303
rect 346 302 352 303
rect 438 302 444 303
rect 278 293 284 294
rect 278 289 279 293
rect 283 289 284 293
rect 278 288 284 289
rect 318 293 324 294
rect 318 289 319 293
rect 323 289 324 293
rect 318 288 324 289
rect 366 293 372 294
rect 366 289 367 293
rect 371 289 372 293
rect 366 288 372 289
rect 414 293 420 294
rect 414 289 415 293
rect 419 289 420 293
rect 414 288 420 289
rect 462 293 468 294
rect 462 289 463 293
rect 467 289 468 293
rect 462 288 468 289
rect 110 286 116 287
rect 112 279 114 286
rect 240 279 242 288
rect 266 287 272 288
rect 266 283 267 287
rect 271 283 272 287
rect 266 282 272 283
rect 280 279 282 288
rect 320 279 322 288
rect 368 279 370 288
rect 416 279 418 288
rect 464 279 466 288
rect 111 278 115 279
rect 111 273 115 274
rect 239 278 243 279
rect 239 273 243 274
rect 279 278 283 279
rect 279 273 283 274
rect 319 278 323 279
rect 319 273 323 274
rect 359 278 363 279
rect 359 273 363 274
rect 367 278 371 279
rect 367 273 371 274
rect 399 278 403 279
rect 399 273 403 274
rect 415 278 419 279
rect 415 273 419 274
rect 439 278 443 279
rect 439 273 443 274
rect 463 278 467 279
rect 463 273 467 274
rect 112 266 114 273
rect 110 265 116 266
rect 110 261 111 265
rect 115 261 116 265
rect 240 264 242 273
rect 280 264 282 273
rect 320 264 322 273
rect 360 264 362 273
rect 400 264 402 273
rect 440 264 442 273
rect 472 266 474 320
rect 480 309 482 325
rect 478 308 484 309
rect 488 308 490 326
rect 511 325 515 326
rect 518 325 524 326
rect 527 325 531 326
rect 575 330 579 331
rect 575 325 579 326
rect 591 330 595 331
rect 591 325 595 326
rect 518 321 519 325
rect 523 321 524 325
rect 518 320 524 321
rect 528 309 530 325
rect 576 309 578 325
rect 526 308 532 309
rect 478 304 479 308
rect 483 304 484 308
rect 478 303 484 304
rect 486 307 492 308
rect 486 303 487 307
rect 491 303 492 307
rect 526 304 527 308
rect 531 304 532 308
rect 526 303 532 304
rect 574 308 580 309
rect 574 304 575 308
rect 579 304 580 308
rect 574 303 580 304
rect 486 302 492 303
rect 510 293 516 294
rect 510 289 511 293
rect 515 289 516 293
rect 510 288 516 289
rect 558 293 564 294
rect 558 289 559 293
rect 563 289 564 293
rect 558 288 564 289
rect 598 293 604 294
rect 598 289 599 293
rect 603 289 604 293
rect 598 288 604 289
rect 608 288 610 338
rect 656 331 658 355
rect 686 354 692 355
rect 688 331 690 354
rect 615 330 619 331
rect 655 330 659 331
rect 687 330 691 331
rect 615 325 619 326
rect 626 325 632 326
rect 655 325 659 326
rect 662 325 668 326
rect 687 325 691 326
rect 616 309 618 325
rect 626 321 627 325
rect 631 321 632 325
rect 626 320 632 321
rect 614 308 620 309
rect 614 304 615 308
rect 619 304 620 308
rect 614 303 620 304
rect 628 296 630 320
rect 656 309 658 325
rect 662 321 663 325
rect 667 321 668 325
rect 662 320 668 321
rect 654 308 660 309
rect 654 304 655 308
rect 659 304 660 308
rect 654 303 660 304
rect 626 295 632 296
rect 626 291 627 295
rect 631 291 632 295
rect 626 290 632 291
rect 638 293 644 294
rect 638 289 639 293
rect 643 289 644 293
rect 638 288 644 289
rect 502 287 508 288
rect 502 283 503 287
rect 507 283 508 287
rect 502 282 508 283
rect 479 278 483 279
rect 479 273 483 274
rect 464 264 474 266
rect 480 264 482 273
rect 110 260 116 261
rect 238 263 244 264
rect 238 259 239 263
rect 243 259 244 263
rect 238 258 244 259
rect 278 263 284 264
rect 278 259 279 263
rect 283 259 284 263
rect 278 258 284 259
rect 318 263 324 264
rect 318 259 319 263
rect 323 259 324 263
rect 318 258 324 259
rect 358 263 364 264
rect 358 259 359 263
rect 363 259 364 263
rect 358 258 364 259
rect 398 263 404 264
rect 398 259 399 263
rect 403 259 404 263
rect 398 258 404 259
rect 438 263 444 264
rect 438 259 439 263
rect 443 259 444 263
rect 438 258 444 259
rect 462 263 468 264
rect 462 259 463 263
rect 467 259 468 263
rect 462 258 468 259
rect 478 263 484 264
rect 478 259 479 263
rect 483 259 484 263
rect 478 258 484 259
rect 254 248 260 249
rect 110 247 116 248
rect 110 243 111 247
rect 115 243 116 247
rect 254 244 255 248
rect 259 244 260 248
rect 254 243 260 244
rect 294 248 300 249
rect 294 244 295 248
rect 299 244 300 248
rect 294 243 300 244
rect 334 248 340 249
rect 334 244 335 248
rect 339 244 340 248
rect 334 243 340 244
rect 374 248 380 249
rect 374 244 375 248
rect 379 244 380 248
rect 374 243 380 244
rect 414 248 420 249
rect 414 244 415 248
rect 419 244 420 248
rect 414 243 420 244
rect 454 248 460 249
rect 454 244 455 248
rect 459 244 460 248
rect 454 243 460 244
rect 494 248 500 249
rect 494 244 495 248
rect 499 244 500 248
rect 494 243 500 244
rect 110 242 116 243
rect 112 211 114 242
rect 256 211 258 243
rect 296 211 298 243
rect 336 211 338 243
rect 376 211 378 243
rect 416 211 418 243
rect 456 211 458 243
rect 496 211 498 243
rect 504 232 506 282
rect 512 279 514 288
rect 560 279 562 288
rect 600 279 602 288
rect 606 287 612 288
rect 606 283 607 287
rect 611 283 612 287
rect 606 282 612 283
rect 640 279 642 288
rect 511 278 515 279
rect 511 273 515 274
rect 519 278 523 279
rect 519 273 523 274
rect 559 278 563 279
rect 559 273 563 274
rect 599 278 603 279
rect 599 273 603 274
rect 639 278 643 279
rect 639 273 643 274
rect 520 264 522 273
rect 560 264 562 273
rect 600 264 602 273
rect 640 264 642 273
rect 664 268 666 320
rect 688 310 690 325
rect 686 309 692 310
rect 686 305 687 309
rect 691 305 692 309
rect 686 304 692 305
rect 686 291 692 292
rect 686 287 687 291
rect 691 287 692 291
rect 686 286 692 287
rect 688 279 690 286
rect 687 278 691 279
rect 687 273 691 274
rect 662 267 668 268
rect 518 263 524 264
rect 518 259 519 263
rect 523 259 524 263
rect 518 258 524 259
rect 558 263 564 264
rect 558 259 559 263
rect 563 259 564 263
rect 558 258 564 259
rect 598 263 604 264
rect 598 259 599 263
rect 603 259 604 263
rect 598 258 604 259
rect 638 263 644 264
rect 638 259 639 263
rect 643 259 644 263
rect 662 263 663 267
rect 667 263 668 267
rect 688 266 690 273
rect 662 262 668 263
rect 686 265 692 266
rect 686 261 687 265
rect 691 261 692 265
rect 686 260 692 261
rect 638 258 644 259
rect 534 248 540 249
rect 534 244 535 248
rect 539 244 540 248
rect 534 243 540 244
rect 574 248 580 249
rect 574 244 575 248
rect 579 244 580 248
rect 574 243 580 244
rect 614 248 620 249
rect 614 244 615 248
rect 619 244 620 248
rect 614 243 620 244
rect 654 248 660 249
rect 654 244 655 248
rect 659 244 660 248
rect 654 243 660 244
rect 686 247 692 248
rect 686 243 687 247
rect 691 243 692 247
rect 502 231 508 232
rect 502 227 503 231
rect 507 227 508 231
rect 502 226 508 227
rect 536 211 538 243
rect 576 211 578 243
rect 616 211 618 243
rect 656 211 658 243
rect 686 242 692 243
rect 688 211 690 242
rect 111 210 115 211
rect 207 210 211 211
rect 247 210 251 211
rect 111 205 115 206
rect 198 205 204 206
rect 207 205 211 206
rect 226 205 232 206
rect 247 205 251 206
rect 255 210 259 211
rect 287 210 291 211
rect 255 205 259 206
rect 262 205 268 206
rect 287 205 291 206
rect 295 210 299 211
rect 295 205 299 206
rect 327 210 331 211
rect 327 205 331 206
rect 335 210 339 211
rect 367 210 371 211
rect 335 205 339 206
rect 346 205 352 206
rect 367 205 371 206
rect 375 210 379 211
rect 407 210 411 211
rect 375 205 379 206
rect 386 205 392 206
rect 407 205 411 206
rect 415 210 419 211
rect 415 205 419 206
rect 455 210 459 211
rect 455 205 459 206
rect 495 210 499 211
rect 495 205 499 206
rect 535 210 539 211
rect 535 205 539 206
rect 575 210 579 211
rect 575 205 579 206
rect 615 210 619 211
rect 615 205 619 206
rect 655 210 659 211
rect 655 205 659 206
rect 687 210 691 211
rect 687 205 691 206
rect 112 190 114 205
rect 198 201 199 205
rect 203 201 204 205
rect 198 200 204 201
rect 110 189 116 190
rect 110 185 111 189
rect 115 185 116 189
rect 110 184 116 185
rect 190 173 196 174
rect 110 171 116 172
rect 110 167 111 171
rect 115 167 116 171
rect 190 169 191 173
rect 195 169 196 173
rect 190 168 196 169
rect 110 166 116 167
rect 112 143 114 166
rect 192 143 194 168
rect 111 142 115 143
rect 111 137 115 138
rect 135 142 139 143
rect 135 137 139 138
rect 175 142 179 143
rect 175 137 179 138
rect 191 142 195 143
rect 191 137 195 138
rect 112 130 114 137
rect 110 129 116 130
rect 110 125 111 129
rect 115 125 116 129
rect 136 128 138 137
rect 176 128 178 137
rect 200 136 202 200
rect 208 189 210 205
rect 226 201 227 205
rect 231 201 232 205
rect 226 200 232 201
rect 206 188 212 189
rect 228 188 230 200
rect 248 189 250 205
rect 262 201 263 205
rect 267 201 268 205
rect 262 200 268 201
rect 246 188 252 189
rect 206 184 207 188
rect 211 184 212 188
rect 206 183 212 184
rect 226 187 232 188
rect 226 183 227 187
rect 231 183 232 187
rect 246 184 247 188
rect 251 184 252 188
rect 264 187 266 200
rect 288 189 290 205
rect 328 189 330 205
rect 346 201 347 205
rect 351 201 352 205
rect 346 200 352 201
rect 246 183 252 184
rect 256 185 266 187
rect 286 188 292 189
rect 226 182 232 183
rect 230 173 236 174
rect 230 169 231 173
rect 235 169 236 173
rect 256 172 258 185
rect 286 184 287 188
rect 291 184 292 188
rect 286 183 292 184
rect 326 188 332 189
rect 348 188 350 200
rect 368 189 370 205
rect 386 201 387 205
rect 391 201 392 205
rect 386 200 392 201
rect 366 188 372 189
rect 388 188 390 200
rect 408 189 410 205
rect 688 190 690 205
rect 686 189 692 190
rect 406 188 412 189
rect 326 184 327 188
rect 331 184 332 188
rect 326 183 332 184
rect 346 187 352 188
rect 346 183 347 187
rect 351 183 352 187
rect 366 184 367 188
rect 371 184 372 188
rect 366 183 372 184
rect 386 187 392 188
rect 386 183 387 187
rect 391 183 392 187
rect 406 184 407 188
rect 411 184 412 188
rect 686 185 687 189
rect 691 185 692 189
rect 686 184 692 185
rect 406 183 412 184
rect 346 182 352 183
rect 386 182 392 183
rect 270 173 276 174
rect 230 168 236 169
rect 254 171 260 172
rect 232 143 234 168
rect 254 167 255 171
rect 259 167 260 171
rect 270 169 271 173
rect 275 169 276 173
rect 270 168 276 169
rect 310 173 316 174
rect 310 169 311 173
rect 315 169 316 173
rect 310 168 316 169
rect 350 173 356 174
rect 350 169 351 173
rect 355 169 356 173
rect 350 168 356 169
rect 390 173 396 174
rect 390 169 391 173
rect 395 169 396 173
rect 390 168 396 169
rect 686 171 692 172
rect 254 166 260 167
rect 272 143 274 168
rect 312 143 314 168
rect 352 143 354 168
rect 392 143 394 168
rect 686 167 687 171
rect 691 167 692 171
rect 686 166 692 167
rect 688 143 690 166
rect 215 142 219 143
rect 215 137 219 138
rect 231 142 235 143
rect 231 137 235 138
rect 255 142 259 143
rect 255 137 259 138
rect 271 142 275 143
rect 271 137 275 138
rect 295 142 299 143
rect 295 137 299 138
rect 311 142 315 143
rect 311 137 315 138
rect 335 142 339 143
rect 335 137 339 138
rect 351 142 355 143
rect 351 137 355 138
rect 375 142 379 143
rect 375 137 379 138
rect 391 142 395 143
rect 391 137 395 138
rect 415 142 419 143
rect 415 137 419 138
rect 455 142 459 143
rect 455 137 459 138
rect 687 142 691 143
rect 687 137 691 138
rect 198 135 204 136
rect 198 131 199 135
rect 203 131 204 135
rect 198 130 204 131
rect 216 128 218 137
rect 256 128 258 137
rect 296 128 298 137
rect 336 128 338 137
rect 376 128 378 137
rect 416 128 418 137
rect 456 128 458 137
rect 688 130 690 137
rect 686 129 692 130
rect 110 124 116 125
rect 134 127 140 128
rect 134 123 135 127
rect 139 123 140 127
rect 134 122 140 123
rect 174 127 180 128
rect 174 123 175 127
rect 179 123 180 127
rect 174 122 180 123
rect 214 127 220 128
rect 214 123 215 127
rect 219 123 220 127
rect 214 122 220 123
rect 254 127 260 128
rect 254 123 255 127
rect 259 123 260 127
rect 254 122 260 123
rect 294 127 300 128
rect 294 123 295 127
rect 299 123 300 127
rect 294 122 300 123
rect 334 127 340 128
rect 334 123 335 127
rect 339 123 340 127
rect 334 122 340 123
rect 374 127 380 128
rect 374 123 375 127
rect 379 123 380 127
rect 374 122 380 123
rect 414 127 420 128
rect 414 123 415 127
rect 419 123 420 127
rect 414 122 420 123
rect 454 127 460 128
rect 454 123 455 127
rect 459 123 460 127
rect 686 125 687 129
rect 691 125 692 129
rect 686 124 692 125
rect 454 122 460 123
rect 150 112 156 113
rect 110 111 116 112
rect 110 107 111 111
rect 115 107 116 111
rect 150 108 151 112
rect 155 108 156 112
rect 150 107 156 108
rect 190 112 196 113
rect 190 108 191 112
rect 195 108 196 112
rect 190 107 196 108
rect 230 112 236 113
rect 230 108 231 112
rect 235 108 236 112
rect 230 107 236 108
rect 270 112 276 113
rect 270 108 271 112
rect 275 108 276 112
rect 270 107 276 108
rect 310 112 316 113
rect 310 108 311 112
rect 315 108 316 112
rect 310 107 316 108
rect 350 112 356 113
rect 350 108 351 112
rect 355 108 356 112
rect 350 107 356 108
rect 390 112 396 113
rect 390 108 391 112
rect 395 108 396 112
rect 390 107 396 108
rect 430 112 436 113
rect 430 108 431 112
rect 435 108 436 112
rect 430 107 436 108
rect 470 112 476 113
rect 470 108 471 112
rect 475 108 476 112
rect 470 107 476 108
rect 686 111 692 112
rect 686 107 687 111
rect 691 107 692 111
rect 110 106 116 107
rect 112 91 114 106
rect 152 91 154 107
rect 192 91 194 107
rect 232 91 234 107
rect 272 91 274 107
rect 312 91 314 107
rect 352 91 354 107
rect 392 91 394 107
rect 432 91 434 107
rect 472 91 474 107
rect 686 106 692 107
rect 688 91 690 106
rect 111 90 115 91
rect 111 85 115 86
rect 151 90 155 91
rect 151 85 155 86
rect 191 90 195 91
rect 191 85 195 86
rect 231 90 235 91
rect 231 85 235 86
rect 271 90 275 91
rect 271 85 275 86
rect 311 90 315 91
rect 311 85 315 86
rect 351 90 355 91
rect 351 85 355 86
rect 391 90 395 91
rect 391 85 395 86
rect 431 90 435 91
rect 431 85 435 86
rect 471 90 475 91
rect 471 85 475 86
rect 687 90 691 91
rect 687 85 691 86
<< m4c >>
rect 111 774 115 778
rect 295 774 299 778
rect 383 774 387 778
rect 479 774 483 778
rect 575 774 579 778
rect 655 774 659 778
rect 687 774 691 778
rect 111 722 115 726
rect 199 722 203 726
rect 239 722 243 726
rect 279 722 283 726
rect 319 722 323 726
rect 359 722 363 726
rect 367 722 371 726
rect 111 666 115 670
rect 175 666 179 670
rect 215 666 219 670
rect 111 606 115 610
rect 159 606 163 610
rect 407 722 411 726
rect 463 722 467 726
rect 527 722 531 726
rect 559 722 563 726
rect 591 722 595 726
rect 639 722 643 726
rect 687 722 691 726
rect 231 666 235 670
rect 255 666 259 670
rect 295 666 299 670
rect 335 666 339 670
rect 367 666 371 670
rect 375 666 379 670
rect 423 666 427 670
rect 439 666 443 670
rect 479 666 483 670
rect 519 666 523 670
rect 543 666 547 670
rect 599 666 603 670
rect 607 666 611 670
rect 655 666 659 670
rect 687 666 691 670
rect 199 606 203 610
rect 215 606 219 610
rect 239 606 243 610
rect 279 606 283 610
rect 295 606 299 610
rect 351 606 355 610
rect 415 606 419 610
rect 423 606 427 610
rect 487 606 491 610
rect 111 550 115 554
rect 215 550 219 554
rect 255 550 259 554
rect 311 550 315 554
rect 327 550 331 554
rect 367 550 371 554
rect 407 550 411 554
rect 503 606 507 610
rect 567 606 571 610
rect 583 606 587 610
rect 639 606 643 610
rect 687 606 691 610
rect 431 550 435 554
rect 455 550 459 554
rect 503 550 507 554
rect 559 550 563 554
rect 583 550 587 554
rect 111 498 115 502
rect 255 498 259 502
rect 295 498 299 502
rect 311 498 315 502
rect 335 498 339 502
rect 351 498 355 502
rect 391 498 395 502
rect 439 498 443 502
rect 447 498 451 502
rect 487 498 491 502
rect 511 498 515 502
rect 615 550 619 554
rect 655 550 659 554
rect 687 550 691 554
rect 543 498 547 502
rect 583 498 587 502
rect 599 498 603 502
rect 639 498 643 502
rect 687 498 691 502
rect 111 442 115 446
rect 175 442 179 446
rect 223 442 227 446
rect 271 442 275 446
rect 279 442 283 446
rect 311 442 315 446
rect 343 442 347 446
rect 351 442 355 446
rect 407 442 411 446
rect 415 442 419 446
rect 463 442 467 446
rect 495 442 499 446
rect 527 442 531 446
rect 111 386 115 390
rect 135 386 139 390
rect 159 386 163 390
rect 175 386 179 390
rect 583 442 587 446
rect 599 442 603 446
rect 655 442 659 446
rect 207 386 211 390
rect 215 386 219 390
rect 263 386 267 390
rect 279 386 283 390
rect 327 386 331 390
rect 343 386 347 390
rect 399 386 403 390
rect 415 386 419 390
rect 479 386 483 390
rect 495 386 499 390
rect 111 326 115 330
rect 151 326 155 330
rect 191 326 195 330
rect 231 326 235 330
rect 255 326 259 330
rect 295 326 299 330
rect 335 326 339 330
rect 359 326 363 330
rect 383 326 387 330
rect 431 326 435 330
rect 479 326 483 330
rect 511 326 515 330
rect 567 386 571 390
rect 575 386 579 390
rect 639 386 643 390
rect 687 442 691 446
rect 687 386 691 390
rect 527 326 531 330
rect 111 274 115 278
rect 239 274 243 278
rect 279 274 283 278
rect 319 274 323 278
rect 359 274 363 278
rect 367 274 371 278
rect 399 274 403 278
rect 415 274 419 278
rect 439 274 443 278
rect 463 274 467 278
rect 575 326 579 330
rect 591 326 595 330
rect 615 326 619 330
rect 655 326 659 330
rect 687 326 691 330
rect 479 274 483 278
rect 511 274 515 278
rect 519 274 523 278
rect 559 274 563 278
rect 599 274 603 278
rect 639 274 643 278
rect 687 274 691 278
rect 111 206 115 210
rect 207 206 211 210
rect 247 206 251 210
rect 255 206 259 210
rect 287 206 291 210
rect 295 206 299 210
rect 327 206 331 210
rect 335 206 339 210
rect 367 206 371 210
rect 375 206 379 210
rect 407 206 411 210
rect 415 206 419 210
rect 455 206 459 210
rect 495 206 499 210
rect 535 206 539 210
rect 575 206 579 210
rect 615 206 619 210
rect 655 206 659 210
rect 687 206 691 210
rect 111 138 115 142
rect 135 138 139 142
rect 175 138 179 142
rect 191 138 195 142
rect 215 138 219 142
rect 231 138 235 142
rect 255 138 259 142
rect 271 138 275 142
rect 295 138 299 142
rect 311 138 315 142
rect 335 138 339 142
rect 351 138 355 142
rect 375 138 379 142
rect 391 138 395 142
rect 415 138 419 142
rect 455 138 459 142
rect 687 138 691 142
rect 111 86 115 90
rect 151 86 155 90
rect 191 86 195 90
rect 231 86 235 90
rect 271 86 275 90
rect 311 86 315 90
rect 351 86 355 90
rect 391 86 395 90
rect 431 86 435 90
rect 471 86 475 90
rect 687 86 691 90
<< m4 >>
rect 84 773 85 779
rect 91 778 711 779
rect 91 774 111 778
rect 115 774 295 778
rect 299 774 383 778
rect 387 774 479 778
rect 483 774 575 778
rect 579 774 655 778
rect 659 774 687 778
rect 691 774 711 778
rect 91 773 711 774
rect 717 773 718 779
rect 96 721 97 727
rect 103 726 723 727
rect 103 722 111 726
rect 115 722 199 726
rect 203 722 239 726
rect 243 722 279 726
rect 283 722 319 726
rect 323 722 359 726
rect 363 722 367 726
rect 371 722 407 726
rect 411 722 463 726
rect 467 722 527 726
rect 531 722 559 726
rect 563 722 591 726
rect 595 722 639 726
rect 643 722 687 726
rect 691 722 723 726
rect 103 721 723 722
rect 729 721 730 727
rect 84 665 85 671
rect 91 670 711 671
rect 91 666 111 670
rect 115 666 175 670
rect 179 666 215 670
rect 219 666 231 670
rect 235 666 255 670
rect 259 666 295 670
rect 299 666 335 670
rect 339 666 367 670
rect 371 666 375 670
rect 379 666 423 670
rect 427 666 439 670
rect 443 666 479 670
rect 483 666 519 670
rect 523 666 543 670
rect 547 666 599 670
rect 603 666 607 670
rect 611 666 655 670
rect 659 666 687 670
rect 691 666 711 670
rect 91 665 711 666
rect 717 665 718 671
rect 96 605 97 611
rect 103 610 723 611
rect 103 606 111 610
rect 115 606 159 610
rect 163 606 199 610
rect 203 606 215 610
rect 219 606 239 610
rect 243 606 279 610
rect 283 606 295 610
rect 299 606 351 610
rect 355 606 415 610
rect 419 606 423 610
rect 427 606 487 610
rect 491 606 503 610
rect 507 606 567 610
rect 571 606 583 610
rect 587 606 639 610
rect 643 606 687 610
rect 691 606 723 610
rect 103 605 723 606
rect 729 605 730 611
rect 84 549 85 555
rect 91 554 711 555
rect 91 550 111 554
rect 115 550 215 554
rect 219 550 255 554
rect 259 550 311 554
rect 315 550 327 554
rect 331 550 367 554
rect 371 550 407 554
rect 411 550 431 554
rect 435 550 455 554
rect 459 550 503 554
rect 507 550 559 554
rect 563 550 583 554
rect 587 550 615 554
rect 619 550 655 554
rect 659 550 687 554
rect 691 550 711 554
rect 91 549 711 550
rect 717 549 718 555
rect 96 497 97 503
rect 103 502 723 503
rect 103 498 111 502
rect 115 498 255 502
rect 259 498 295 502
rect 299 498 311 502
rect 315 498 335 502
rect 339 498 351 502
rect 355 498 391 502
rect 395 498 439 502
rect 443 498 447 502
rect 451 498 487 502
rect 491 498 511 502
rect 515 498 543 502
rect 547 498 583 502
rect 587 498 599 502
rect 603 498 639 502
rect 643 498 687 502
rect 691 498 723 502
rect 103 497 723 498
rect 729 497 730 503
rect 84 441 85 447
rect 91 446 711 447
rect 91 442 111 446
rect 115 442 175 446
rect 179 442 223 446
rect 227 442 271 446
rect 275 442 279 446
rect 283 442 311 446
rect 315 442 343 446
rect 347 442 351 446
rect 355 442 407 446
rect 411 442 415 446
rect 419 442 463 446
rect 467 442 495 446
rect 499 442 527 446
rect 531 442 583 446
rect 587 442 599 446
rect 603 442 655 446
rect 659 442 687 446
rect 691 442 711 446
rect 91 441 711 442
rect 717 441 718 447
rect 96 385 97 391
rect 103 390 723 391
rect 103 386 111 390
rect 115 386 135 390
rect 139 386 159 390
rect 163 386 175 390
rect 179 386 207 390
rect 211 386 215 390
rect 219 386 263 390
rect 267 386 279 390
rect 283 386 327 390
rect 331 386 343 390
rect 347 386 399 390
rect 403 386 415 390
rect 419 386 479 390
rect 483 386 495 390
rect 499 386 567 390
rect 571 386 575 390
rect 579 386 639 390
rect 643 386 687 390
rect 691 386 723 390
rect 103 385 723 386
rect 729 385 730 391
rect 84 325 85 331
rect 91 330 711 331
rect 91 326 111 330
rect 115 326 151 330
rect 155 326 191 330
rect 195 326 231 330
rect 235 326 255 330
rect 259 326 295 330
rect 299 326 335 330
rect 339 326 359 330
rect 363 326 383 330
rect 387 326 431 330
rect 435 326 479 330
rect 483 326 511 330
rect 515 326 527 330
rect 531 326 575 330
rect 579 326 591 330
rect 595 326 615 330
rect 619 326 655 330
rect 659 326 687 330
rect 691 326 711 330
rect 91 325 711 326
rect 717 325 718 331
rect 96 273 97 279
rect 103 278 723 279
rect 103 274 111 278
rect 115 274 239 278
rect 243 274 279 278
rect 283 274 319 278
rect 323 274 359 278
rect 363 274 367 278
rect 371 274 399 278
rect 403 274 415 278
rect 419 274 439 278
rect 443 274 463 278
rect 467 274 479 278
rect 483 274 511 278
rect 515 274 519 278
rect 523 274 559 278
rect 563 274 599 278
rect 603 274 639 278
rect 643 274 687 278
rect 691 274 723 278
rect 103 273 723 274
rect 729 273 730 279
rect 84 205 85 211
rect 91 210 711 211
rect 91 206 111 210
rect 115 206 207 210
rect 211 206 247 210
rect 251 206 255 210
rect 259 206 287 210
rect 291 206 295 210
rect 299 206 327 210
rect 331 206 335 210
rect 339 206 367 210
rect 371 206 375 210
rect 379 206 407 210
rect 411 206 415 210
rect 419 206 455 210
rect 459 206 495 210
rect 499 206 535 210
rect 539 206 575 210
rect 579 206 615 210
rect 619 206 655 210
rect 659 206 687 210
rect 691 206 711 210
rect 91 205 711 206
rect 717 205 718 211
rect 96 137 97 143
rect 103 142 723 143
rect 103 138 111 142
rect 115 138 135 142
rect 139 138 175 142
rect 179 138 191 142
rect 195 138 215 142
rect 219 138 231 142
rect 235 138 255 142
rect 259 138 271 142
rect 275 138 295 142
rect 299 138 311 142
rect 315 138 335 142
rect 339 138 351 142
rect 355 138 375 142
rect 379 138 391 142
rect 395 138 415 142
rect 419 138 455 142
rect 459 138 687 142
rect 691 138 723 142
rect 103 137 723 138
rect 729 137 730 143
rect 84 85 85 91
rect 91 90 711 91
rect 91 86 111 90
rect 115 86 151 90
rect 155 86 191 90
rect 195 86 231 90
rect 235 86 271 90
rect 275 86 311 90
rect 315 86 351 90
rect 355 86 391 90
rect 395 86 431 90
rect 435 86 471 90
rect 475 86 687 90
rect 691 86 711 90
rect 91 85 711 86
rect 717 85 718 91
<< m5c >>
rect 85 773 91 779
rect 711 773 717 779
rect 97 721 103 727
rect 723 721 729 727
rect 85 665 91 671
rect 711 665 717 671
rect 97 605 103 611
rect 723 605 729 611
rect 85 549 91 555
rect 711 549 717 555
rect 97 497 103 503
rect 723 497 729 503
rect 85 441 91 447
rect 711 441 717 447
rect 97 385 103 391
rect 723 385 729 391
rect 85 325 91 331
rect 711 325 717 331
rect 97 273 103 279
rect 723 273 729 279
rect 85 205 91 211
rect 711 205 717 211
rect 97 137 103 143
rect 723 137 729 143
rect 85 85 91 91
rect 711 85 717 91
<< m5 >>
rect 84 779 92 792
rect 84 773 85 779
rect 91 773 92 779
rect 84 671 92 773
rect 84 665 85 671
rect 91 665 92 671
rect 84 555 92 665
rect 84 549 85 555
rect 91 549 92 555
rect 84 447 92 549
rect 84 441 85 447
rect 91 441 92 447
rect 84 331 92 441
rect 84 325 85 331
rect 91 325 92 331
rect 84 211 92 325
rect 84 205 85 211
rect 91 205 92 211
rect 84 91 92 205
rect 84 85 85 91
rect 91 85 92 91
rect 84 72 92 85
rect 96 727 104 792
rect 96 721 97 727
rect 103 721 104 727
rect 96 611 104 721
rect 96 605 97 611
rect 103 605 104 611
rect 96 503 104 605
rect 96 497 97 503
rect 103 497 104 503
rect 96 391 104 497
rect 96 385 97 391
rect 103 385 104 391
rect 96 279 104 385
rect 96 273 97 279
rect 103 273 104 279
rect 96 143 104 273
rect 96 137 97 143
rect 103 137 104 143
rect 96 72 104 137
rect 710 779 718 792
rect 710 773 711 779
rect 717 773 718 779
rect 710 671 718 773
rect 710 665 711 671
rect 717 665 718 671
rect 710 555 718 665
rect 710 549 711 555
rect 717 549 718 555
rect 710 447 718 549
rect 710 441 711 447
rect 717 441 718 447
rect 710 331 718 441
rect 710 325 711 331
rect 717 325 718 331
rect 710 211 718 325
rect 710 205 711 211
rect 717 205 718 211
rect 710 91 718 205
rect 710 85 711 91
rect 717 85 718 91
rect 710 72 718 85
rect 722 727 730 792
rect 722 721 723 727
rect 729 721 730 727
rect 722 611 730 721
rect 722 605 723 611
rect 729 605 730 611
rect 722 503 730 605
rect 722 497 723 503
rect 729 497 730 503
rect 722 391 730 497
rect 722 385 723 391
rect 729 385 730 391
rect 722 279 730 385
rect 722 273 723 279
rect 729 273 730 279
rect 722 143 730 273
rect 722 137 723 143
rect 729 137 730 143
rect 722 72 730 137
use circuitppnp  ppnps
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use circuitwell  npwells
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use circuitppnp  ppnps
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use circuitwell  npwells
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use circuitppnp  ppnps
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use circuitwell  npwells
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use _0_0std_0_0cells_0_0AND2X1  and_50_6
timestamp 1730743719
transform 1 0 128 0 1 88
box 8 4 36 49
use welltap_svt  __well_tap__0
timestamp 1730743719
transform 1 0 104 0 1 104
box 8 4 12 24
use _0_0std_0_0cells_0_0AND2X1  and_50_6
timestamp 1730743719
transform 1 0 128 0 1 88
box 8 4 36 49
use welltap_svt  __well_tap__0
timestamp 1730743719
transform 1 0 104 0 1 104
box 8 4 12 24
use _0_0std_0_0cells_0_0AND2X1  and_50_6
timestamp 1730743719
transform 1 0 128 0 1 88
box 8 4 36 49
use welltap_svt  __well_tap__0
timestamp 1730743719
transform 1 0 104 0 1 104
box 8 4 12 24
use _0_0std_0_0cells_0_0AND2X1  and_51_6
timestamp 1730743719
transform 1 0 168 0 1 88
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_51_6
timestamp 1730743719
transform 1 0 168 0 1 88
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_51_6
timestamp 1730743719
transform 1 0 168 0 1 88
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_52_6
timestamp 1730743719
transform 1 0 208 0 1 88
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_52_6
timestamp 1730743719
transform 1 0 208 0 1 88
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_52_6
timestamp 1730743719
transform 1 0 208 0 1 88
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_53_6
timestamp 1730743719
transform 1 0 248 0 1 88
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_53_6
timestamp 1730743719
transform 1 0 248 0 1 88
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_53_6
timestamp 1730743719
transform 1 0 248 0 1 88
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_54_6
timestamp 1730743719
transform 1 0 288 0 1 88
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_54_6
timestamp 1730743719
transform 1 0 288 0 1 88
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_54_6
timestamp 1730743719
transform 1 0 288 0 1 88
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_55_6
timestamp 1730743719
transform 1 0 328 0 1 88
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_55_6
timestamp 1730743719
transform 1 0 328 0 1 88
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_55_6
timestamp 1730743719
transform 1 0 328 0 1 88
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_56_6
timestamp 1730743719
transform 1 0 368 0 1 88
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_56_6
timestamp 1730743719
transform 1 0 368 0 1 88
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_56_6
timestamp 1730743719
transform 1 0 368 0 1 88
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_57_6
timestamp 1730743719
transform 1 0 408 0 1 88
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_57_6
timestamp 1730743719
transform 1 0 408 0 1 88
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_57_6
timestamp 1730743719
transform 1 0 408 0 1 88
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_58_6
timestamp 1730743719
transform 1 0 448 0 1 88
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_58_6
timestamp 1730743719
transform 1 0 448 0 1 88
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_58_6
timestamp 1730743719
transform 1 0 448 0 1 88
box 8 4 36 49
use welltap_svt  __well_tap__1
timestamp 1730743719
transform 1 0 680 0 1 104
box 8 4 12 24
use welltap_svt  __well_tap__1
timestamp 1730743719
transform 1 0 680 0 1 104
box 8 4 12 24
use welltap_svt  __well_tap__1
timestamp 1730743719
transform 1 0 680 0 1 104
box 8 4 12 24
use _0_0std_0_0cells_0_0AND2X1  and_59_6
timestamp 1730743719
transform 1 0 184 0 -1 208
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_59_6
timestamp 1730743719
transform 1 0 184 0 -1 208
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_59_6
timestamp 1730743719
transform 1 0 184 0 -1 208
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_510_6
timestamp 1730743719
transform 1 0 224 0 -1 208
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_510_6
timestamp 1730743719
transform 1 0 224 0 -1 208
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_510_6
timestamp 1730743719
transform 1 0 224 0 -1 208
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_511_6
timestamp 1730743719
transform 1 0 264 0 -1 208
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_511_6
timestamp 1730743719
transform 1 0 264 0 -1 208
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_511_6
timestamp 1730743719
transform 1 0 264 0 -1 208
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_512_6
timestamp 1730743719
transform 1 0 304 0 -1 208
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_512_6
timestamp 1730743719
transform 1 0 304 0 -1 208
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_512_6
timestamp 1730743719
transform 1 0 304 0 -1 208
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_513_6
timestamp 1730743719
transform 1 0 344 0 -1 208
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_513_6
timestamp 1730743719
transform 1 0 344 0 -1 208
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_513_6
timestamp 1730743719
transform 1 0 344 0 -1 208
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_514_6
timestamp 1730743719
transform 1 0 384 0 -1 208
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_514_6
timestamp 1730743719
transform 1 0 384 0 -1 208
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_514_6
timestamp 1730743719
transform 1 0 384 0 -1 208
box 8 4 36 49
use welltap_svt  __well_tap__2
timestamp 1730743719
transform 1 0 104 0 -1 192
box 8 4 12 24
use welltap_svt  __well_tap__2
timestamp 1730743719
transform 1 0 104 0 -1 192
box 8 4 12 24
use welltap_svt  __well_tap__2
timestamp 1730743719
transform 1 0 104 0 -1 192
box 8 4 12 24
use welltap_svt  __well_tap__3
timestamp 1730743719
transform 1 0 680 0 -1 192
box 8 4 12 24
use welltap_svt  __well_tap__3
timestamp 1730743719
transform 1 0 680 0 -1 192
box 8 4 12 24
use welltap_svt  __well_tap__3
timestamp 1730743719
transform 1 0 680 0 -1 192
box 8 4 12 24
use welltap_svt  __well_tap__4
timestamp 1730743719
transform 1 0 104 0 1 240
box 8 4 12 24
use welltap_svt  __well_tap__4
timestamp 1730743719
transform 1 0 104 0 1 240
box 8 4 12 24
use welltap_svt  __well_tap__4
timestamp 1730743719
transform 1 0 104 0 1 240
box 8 4 12 24
use _0_0std_0_0cells_0_0AND2X1  and_515_6
timestamp 1730743719
transform 1 0 232 0 1 224
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_515_6
timestamp 1730743719
transform 1 0 232 0 1 224
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_515_6
timestamp 1730743719
transform 1 0 232 0 1 224
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_516_6
timestamp 1730743719
transform 1 0 272 0 1 224
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_516_6
timestamp 1730743719
transform 1 0 272 0 1 224
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_516_6
timestamp 1730743719
transform 1 0 272 0 1 224
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_517_6
timestamp 1730743719
transform 1 0 312 0 1 224
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_517_6
timestamp 1730743719
transform 1 0 312 0 1 224
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_517_6
timestamp 1730743719
transform 1 0 312 0 1 224
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_518_6
timestamp 1730743719
transform 1 0 352 0 1 224
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_518_6
timestamp 1730743719
transform 1 0 352 0 1 224
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_518_6
timestamp 1730743719
transform 1 0 352 0 1 224
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_519_6
timestamp 1730743719
transform 1 0 392 0 1 224
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_519_6
timestamp 1730743719
transform 1 0 392 0 1 224
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_519_6
timestamp 1730743719
transform 1 0 392 0 1 224
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_520_6
timestamp 1730743719
transform 1 0 432 0 1 224
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_520_6
timestamp 1730743719
transform 1 0 432 0 1 224
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_520_6
timestamp 1730743719
transform 1 0 432 0 1 224
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_581_6
timestamp 1730743719
transform 1 0 472 0 1 224
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_581_6
timestamp 1730743719
transform 1 0 472 0 1 224
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_581_6
timestamp 1730743719
transform 1 0 472 0 1 224
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_582_6
timestamp 1730743719
transform 1 0 512 0 1 224
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_582_6
timestamp 1730743719
transform 1 0 512 0 1 224
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_582_6
timestamp 1730743719
transform 1 0 512 0 1 224
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_583_6
timestamp 1730743719
transform 1 0 552 0 1 224
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_583_6
timestamp 1730743719
transform 1 0 552 0 1 224
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_583_6
timestamp 1730743719
transform 1 0 552 0 1 224
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_584_6
timestamp 1730743719
transform 1 0 592 0 1 224
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_584_6
timestamp 1730743719
transform 1 0 592 0 1 224
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_584_6
timestamp 1730743719
transform 1 0 592 0 1 224
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_585_6
timestamp 1730743719
transform 1 0 632 0 1 224
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_585_6
timestamp 1730743719
transform 1 0 632 0 1 224
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_585_6
timestamp 1730743719
transform 1 0 632 0 1 224
box 8 4 36 49
use welltap_svt  __well_tap__5
timestamp 1730743719
transform 1 0 680 0 1 240
box 8 4 12 24
use welltap_svt  __well_tap__5
timestamp 1730743719
transform 1 0 680 0 1 240
box 8 4 12 24
use welltap_svt  __well_tap__5
timestamp 1730743719
transform 1 0 680 0 1 240
box 8 4 12 24
use welltap_svt  __well_tap__6
timestamp 1730743719
transform 1 0 104 0 -1 312
box 8 4 12 24
use welltap_svt  __well_tap__6
timestamp 1730743719
transform 1 0 104 0 -1 312
box 8 4 12 24
use welltap_svt  __well_tap__6
timestamp 1730743719
transform 1 0 104 0 -1 312
box 8 4 12 24
use _0_0std_0_0cells_0_0AND2X1  and_524_6
timestamp 1730743719
transform 1 0 232 0 -1 328
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_524_6
timestamp 1730743719
transform 1 0 232 0 -1 328
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_524_6
timestamp 1730743719
transform 1 0 232 0 -1 328
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_525_6
timestamp 1730743719
transform 1 0 272 0 -1 328
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_525_6
timestamp 1730743719
transform 1 0 272 0 -1 328
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_525_6
timestamp 1730743719
transform 1 0 272 0 -1 328
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_526_6
timestamp 1730743719
transform 1 0 312 0 -1 328
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_526_6
timestamp 1730743719
transform 1 0 312 0 -1 328
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_526_6
timestamp 1730743719
transform 1 0 312 0 -1 328
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_523_6
timestamp 1730743719
transform 1 0 360 0 -1 328
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_523_6
timestamp 1730743719
transform 1 0 360 0 -1 328
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_523_6
timestamp 1730743719
transform 1 0 360 0 -1 328
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_522_6
timestamp 1730743719
transform 1 0 408 0 -1 328
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_522_6
timestamp 1730743719
transform 1 0 408 0 -1 328
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_522_6
timestamp 1730743719
transform 1 0 408 0 -1 328
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_521_6
timestamp 1730743719
transform 1 0 456 0 -1 328
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_521_6
timestamp 1730743719
transform 1 0 456 0 -1 328
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_521_6
timestamp 1730743719
transform 1 0 456 0 -1 328
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_579_6
timestamp 1730743719
transform 1 0 504 0 -1 328
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_579_6
timestamp 1730743719
transform 1 0 504 0 -1 328
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_579_6
timestamp 1730743719
transform 1 0 504 0 -1 328
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_580_6
timestamp 1730743719
transform 1 0 552 0 -1 328
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_580_6
timestamp 1730743719
transform 1 0 552 0 -1 328
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_580_6
timestamp 1730743719
transform 1 0 552 0 -1 328
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_587_6
timestamp 1730743719
transform 1 0 592 0 -1 328
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_587_6
timestamp 1730743719
transform 1 0 592 0 -1 328
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_587_6
timestamp 1730743719
transform 1 0 592 0 -1 328
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_586_6
timestamp 1730743719
transform 1 0 632 0 -1 328
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_586_6
timestamp 1730743719
transform 1 0 632 0 -1 328
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_586_6
timestamp 1730743719
transform 1 0 632 0 -1 328
box 8 4 36 49
use welltap_svt  __well_tap__7
timestamp 1730743719
transform 1 0 680 0 -1 312
box 8 4 12 24
use welltap_svt  __well_tap__7
timestamp 1730743719
transform 1 0 680 0 -1 312
box 8 4 12 24
use welltap_svt  __well_tap__7
timestamp 1730743719
transform 1 0 680 0 -1 312
box 8 4 12 24
use _0_0std_0_0cells_0_0AND2X1  and_531_6
timestamp 1730743719
transform 1 0 128 0 1 336
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_531_6
timestamp 1730743719
transform 1 0 128 0 1 336
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_531_6
timestamp 1730743719
transform 1 0 128 0 1 336
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_532_6
timestamp 1730743719
transform 1 0 168 0 1 336
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_532_6
timestamp 1730743719
transform 1 0 168 0 1 336
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_532_6
timestamp 1730743719
transform 1 0 168 0 1 336
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_530_6
timestamp 1730743719
transform 1 0 208 0 1 336
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_530_6
timestamp 1730743719
transform 1 0 208 0 1 336
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_530_6
timestamp 1730743719
transform 1 0 208 0 1 336
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_529_6
timestamp 1730743719
transform 1 0 272 0 1 336
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_529_6
timestamp 1730743719
transform 1 0 272 0 1 336
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_529_6
timestamp 1730743719
transform 1 0 272 0 1 336
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_527_6
timestamp 1730743719
transform 1 0 336 0 1 336
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_527_6
timestamp 1730743719
transform 1 0 336 0 1 336
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_527_6
timestamp 1730743719
transform 1 0 336 0 1 336
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_528_6
timestamp 1730743719
transform 1 0 408 0 1 336
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_528_6
timestamp 1730743719
transform 1 0 408 0 1 336
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_528_6
timestamp 1730743719
transform 1 0 408 0 1 336
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_578_6
timestamp 1730743719
transform 1 0 488 0 1 336
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_578_6
timestamp 1730743719
transform 1 0 488 0 1 336
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_578_6
timestamp 1730743719
transform 1 0 488 0 1 336
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_588_6
timestamp 1730743719
transform 1 0 568 0 1 336
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_588_6
timestamp 1730743719
transform 1 0 568 0 1 336
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_588_6
timestamp 1730743719
transform 1 0 568 0 1 336
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_589_6
timestamp 1730743719
transform 1 0 632 0 1 336
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_589_6
timestamp 1730743719
transform 1 0 632 0 1 336
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_589_6
timestamp 1730743719
transform 1 0 632 0 1 336
box 8 4 36 49
use welltap_svt  __well_tap__8
timestamp 1730743719
transform 1 0 104 0 1 352
box 8 4 12 24
use welltap_svt  __well_tap__8
timestamp 1730743719
transform 1 0 104 0 1 352
box 8 4 12 24
use welltap_svt  __well_tap__8
timestamp 1730743719
transform 1 0 104 0 1 352
box 8 4 12 24
use welltap_svt  __well_tap__9
timestamp 1730743719
transform 1 0 680 0 1 352
box 8 4 12 24
use welltap_svt  __well_tap__9
timestamp 1730743719
transform 1 0 680 0 1 352
box 8 4 12 24
use welltap_svt  __well_tap__9
timestamp 1730743719
transform 1 0 680 0 1 352
box 8 4 12 24
use welltap_svt  __well_tap__10
timestamp 1730743719
transform 1 0 104 0 -1 428
box 8 4 12 24
use welltap_svt  __well_tap__10
timestamp 1730743719
transform 1 0 104 0 -1 428
box 8 4 12 24
use welltap_svt  __well_tap__10
timestamp 1730743719
transform 1 0 104 0 -1 428
box 8 4 12 24
use _0_0std_0_0cells_0_0AND2X1  and_533_6
timestamp 1730743719
transform 1 0 152 0 -1 444
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_533_6
timestamp 1730743719
transform 1 0 152 0 -1 444
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_533_6
timestamp 1730743719
transform 1 0 152 0 -1 444
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_534_6
timestamp 1730743719
transform 1 0 200 0 -1 444
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_534_6
timestamp 1730743719
transform 1 0 200 0 -1 444
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_534_6
timestamp 1730743719
transform 1 0 200 0 -1 444
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_535_6
timestamp 1730743719
transform 1 0 256 0 -1 444
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_535_6
timestamp 1730743719
transform 1 0 256 0 -1 444
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_535_6
timestamp 1730743719
transform 1 0 256 0 -1 444
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_536_6
timestamp 1730743719
transform 1 0 320 0 -1 444
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_536_6
timestamp 1730743719
transform 1 0 320 0 -1 444
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_536_6
timestamp 1730743719
transform 1 0 320 0 -1 444
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_537_6
timestamp 1730743719
transform 1 0 392 0 -1 444
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_537_6
timestamp 1730743719
transform 1 0 392 0 -1 444
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_537_6
timestamp 1730743719
transform 1 0 392 0 -1 444
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_538_6
timestamp 1730743719
transform 1 0 472 0 -1 444
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_538_6
timestamp 1730743719
transform 1 0 472 0 -1 444
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_538_6
timestamp 1730743719
transform 1 0 472 0 -1 444
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_577_6
timestamp 1730743719
transform 1 0 560 0 -1 444
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_577_6
timestamp 1730743719
transform 1 0 560 0 -1 444
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_577_6
timestamp 1730743719
transform 1 0 560 0 -1 444
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_590_6
timestamp 1730743719
transform 1 0 632 0 -1 444
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_590_6
timestamp 1730743719
transform 1 0 632 0 -1 444
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_590_6
timestamp 1730743719
transform 1 0 632 0 -1 444
box 8 4 36 49
use welltap_svt  __well_tap__11
timestamp 1730743719
transform 1 0 680 0 -1 428
box 8 4 12 24
use welltap_svt  __well_tap__11
timestamp 1730743719
transform 1 0 680 0 -1 428
box 8 4 12 24
use welltap_svt  __well_tap__11
timestamp 1730743719
transform 1 0 680 0 -1 428
box 8 4 12 24
use welltap_svt  __well_tap__12
timestamp 1730743719
transform 1 0 104 0 1 464
box 8 4 12 24
use welltap_svt  __well_tap__12
timestamp 1730743719
transform 1 0 104 0 1 464
box 8 4 12 24
use welltap_svt  __well_tap__12
timestamp 1730743719
transform 1 0 104 0 1 464
box 8 4 12 24
use _0_0std_0_0cells_0_0AND2X1  and_539_6
timestamp 1730743719
transform 1 0 248 0 1 448
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_539_6
timestamp 1730743719
transform 1 0 248 0 1 448
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_539_6
timestamp 1730743719
transform 1 0 248 0 1 448
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_540_6
timestamp 1730743719
transform 1 0 288 0 1 448
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_540_6
timestamp 1730743719
transform 1 0 288 0 1 448
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_540_6
timestamp 1730743719
transform 1 0 288 0 1 448
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_541_6
timestamp 1730743719
transform 1 0 328 0 1 448
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_541_6
timestamp 1730743719
transform 1 0 328 0 1 448
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_541_6
timestamp 1730743719
transform 1 0 328 0 1 448
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_542_6
timestamp 1730743719
transform 1 0 384 0 1 448
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_542_6
timestamp 1730743719
transform 1 0 384 0 1 448
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_542_6
timestamp 1730743719
transform 1 0 384 0 1 448
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_543_6
timestamp 1730743719
transform 1 0 440 0 1 448
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_543_6
timestamp 1730743719
transform 1 0 440 0 1 448
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_543_6
timestamp 1730743719
transform 1 0 440 0 1 448
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_544_6
timestamp 1730743719
transform 1 0 504 0 1 448
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_544_6
timestamp 1730743719
transform 1 0 504 0 1 448
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_544_6
timestamp 1730743719
transform 1 0 504 0 1 448
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_576_6
timestamp 1730743719
transform 1 0 576 0 1 448
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_576_6
timestamp 1730743719
transform 1 0 576 0 1 448
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_576_6
timestamp 1730743719
transform 1 0 576 0 1 448
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_591_6
timestamp 1730743719
transform 1 0 632 0 1 448
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_591_6
timestamp 1730743719
transform 1 0 632 0 1 448
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_591_6
timestamp 1730743719
transform 1 0 632 0 1 448
box 8 4 36 49
use welltap_svt  __well_tap__13
timestamp 1730743719
transform 1 0 680 0 1 464
box 8 4 12 24
use welltap_svt  __well_tap__13
timestamp 1730743719
transform 1 0 680 0 1 464
box 8 4 12 24
use welltap_svt  __well_tap__13
timestamp 1730743719
transform 1 0 680 0 1 464
box 8 4 12 24
use welltap_svt  __well_tap__14
timestamp 1730743719
transform 1 0 104 0 -1 536
box 8 4 12 24
use welltap_svt  __well_tap__14
timestamp 1730743719
transform 1 0 104 0 -1 536
box 8 4 12 24
use welltap_svt  __well_tap__14
timestamp 1730743719
transform 1 0 104 0 -1 536
box 8 4 12 24
use _0_0std_0_0cells_0_0AND2X1  and_547_6
timestamp 1730743719
transform 1 0 304 0 -1 552
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_547_6
timestamp 1730743719
transform 1 0 304 0 -1 552
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_547_6
timestamp 1730743719
transform 1 0 304 0 -1 552
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_548_6
timestamp 1730743719
transform 1 0 344 0 -1 552
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_548_6
timestamp 1730743719
transform 1 0 344 0 -1 552
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_548_6
timestamp 1730743719
transform 1 0 344 0 -1 552
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_549_6
timestamp 1730743719
transform 1 0 384 0 -1 552
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_549_6
timestamp 1730743719
transform 1 0 384 0 -1 552
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_549_6
timestamp 1730743719
transform 1 0 384 0 -1 552
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_546_6
timestamp 1730743719
transform 1 0 432 0 -1 552
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_546_6
timestamp 1730743719
transform 1 0 432 0 -1 552
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_546_6
timestamp 1730743719
transform 1 0 432 0 -1 552
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_545_6
timestamp 1730743719
transform 1 0 480 0 -1 552
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_545_6
timestamp 1730743719
transform 1 0 480 0 -1 552
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_545_6
timestamp 1730743719
transform 1 0 480 0 -1 552
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_575_6
timestamp 1730743719
transform 1 0 536 0 -1 552
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_575_6
timestamp 1730743719
transform 1 0 536 0 -1 552
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_575_6
timestamp 1730743719
transform 1 0 536 0 -1 552
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_593_6
timestamp 1730743719
transform 1 0 592 0 -1 552
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_593_6
timestamp 1730743719
transform 1 0 592 0 -1 552
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_593_6
timestamp 1730743719
transform 1 0 592 0 -1 552
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_592_6
timestamp 1730743719
transform 1 0 632 0 -1 552
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_592_6
timestamp 1730743719
transform 1 0 632 0 -1 552
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_592_6
timestamp 1730743719
transform 1 0 632 0 -1 552
box 8 4 36 49
use welltap_svt  __well_tap__15
timestamp 1730743719
transform 1 0 680 0 -1 536
box 8 4 12 24
use welltap_svt  __well_tap__15
timestamp 1730743719
transform 1 0 680 0 -1 536
box 8 4 12 24
use welltap_svt  __well_tap__15
timestamp 1730743719
transform 1 0 680 0 -1 536
box 8 4 12 24
use welltap_svt  __well_tap__16
timestamp 1730743719
transform 1 0 104 0 1 572
box 8 4 12 24
use welltap_svt  __well_tap__16
timestamp 1730743719
transform 1 0 104 0 1 572
box 8 4 12 24
use welltap_svt  __well_tap__16
timestamp 1730743719
transform 1 0 104 0 1 572
box 8 4 12 24
use _0_0std_0_0cells_0_0AND2X1  and_554_6
timestamp 1730743719
transform 1 0 192 0 1 556
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_554_6
timestamp 1730743719
transform 1 0 192 0 1 556
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_554_6
timestamp 1730743719
transform 1 0 192 0 1 556
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_553_6
timestamp 1730743719
transform 1 0 232 0 1 556
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_553_6
timestamp 1730743719
transform 1 0 232 0 1 556
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_553_6
timestamp 1730743719
transform 1 0 232 0 1 556
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_552_6
timestamp 1730743719
transform 1 0 288 0 1 556
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_552_6
timestamp 1730743719
transform 1 0 288 0 1 556
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_552_6
timestamp 1730743719
transform 1 0 288 0 1 556
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_551_6
timestamp 1730743719
transform 1 0 344 0 1 556
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_551_6
timestamp 1730743719
transform 1 0 344 0 1 556
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_551_6
timestamp 1730743719
transform 1 0 344 0 1 556
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_550_6
timestamp 1730743719
transform 1 0 408 0 1 556
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_550_6
timestamp 1730743719
transform 1 0 408 0 1 556
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_550_6
timestamp 1730743719
transform 1 0 408 0 1 556
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_573_6
timestamp 1730743719
transform 1 0 480 0 1 556
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_573_6
timestamp 1730743719
transform 1 0 480 0 1 556
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_573_6
timestamp 1730743719
transform 1 0 480 0 1 556
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_574_6
timestamp 1730743719
transform 1 0 560 0 1 556
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_574_6
timestamp 1730743719
transform 1 0 560 0 1 556
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_574_6
timestamp 1730743719
transform 1 0 560 0 1 556
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_594_6
timestamp 1730743719
transform 1 0 632 0 1 556
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_594_6
timestamp 1730743719
transform 1 0 632 0 1 556
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_594_6
timestamp 1730743719
transform 1 0 632 0 1 556
box 8 4 36 49
use welltap_svt  __well_tap__17
timestamp 1730743719
transform 1 0 680 0 1 572
box 8 4 12 24
use welltap_svt  __well_tap__17
timestamp 1730743719
transform 1 0 680 0 1 572
box 8 4 12 24
use welltap_svt  __well_tap__17
timestamp 1730743719
transform 1 0 680 0 1 572
box 8 4 12 24
use _0_0std_0_0cells_0_0AND2X1  and_555_6
timestamp 1730743719
transform 1 0 152 0 -1 668
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_555_6
timestamp 1730743719
transform 1 0 152 0 -1 668
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_555_6
timestamp 1730743719
transform 1 0 152 0 -1 668
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_556_6
timestamp 1730743719
transform 1 0 208 0 -1 668
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_556_6
timestamp 1730743719
transform 1 0 208 0 -1 668
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_556_6
timestamp 1730743719
transform 1 0 208 0 -1 668
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_557_6
timestamp 1730743719
transform 1 0 272 0 -1 668
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_557_6
timestamp 1730743719
transform 1 0 272 0 -1 668
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_557_6
timestamp 1730743719
transform 1 0 272 0 -1 668
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_558_6
timestamp 1730743719
transform 1 0 344 0 -1 668
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_558_6
timestamp 1730743719
transform 1 0 344 0 -1 668
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_558_6
timestamp 1730743719
transform 1 0 344 0 -1 668
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_572_6
timestamp 1730743719
transform 1 0 416 0 -1 668
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_572_6
timestamp 1730743719
transform 1 0 416 0 -1 668
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_572_6
timestamp 1730743719
transform 1 0 416 0 -1 668
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_571_6
timestamp 1730743719
transform 1 0 496 0 -1 668
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_571_6
timestamp 1730743719
transform 1 0 496 0 -1 668
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_571_6
timestamp 1730743719
transform 1 0 496 0 -1 668
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_596_6
timestamp 1730743719
transform 1 0 576 0 -1 668
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_596_6
timestamp 1730743719
transform 1 0 576 0 -1 668
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_596_6
timestamp 1730743719
transform 1 0 576 0 -1 668
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_595_6
timestamp 1730743719
transform 1 0 632 0 -1 668
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_595_6
timestamp 1730743719
transform 1 0 632 0 -1 668
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_595_6
timestamp 1730743719
transform 1 0 632 0 -1 668
box 8 4 36 49
use welltap_svt  __well_tap__18
timestamp 1730743719
transform 1 0 104 0 -1 652
box 8 4 12 24
use welltap_svt  __well_tap__18
timestamp 1730743719
transform 1 0 104 0 -1 652
box 8 4 12 24
use welltap_svt  __well_tap__18
timestamp 1730743719
transform 1 0 104 0 -1 652
box 8 4 12 24
use welltap_svt  __well_tap__19
timestamp 1730743719
transform 1 0 680 0 -1 652
box 8 4 12 24
use welltap_svt  __well_tap__19
timestamp 1730743719
transform 1 0 680 0 -1 652
box 8 4 12 24
use welltap_svt  __well_tap__19
timestamp 1730743719
transform 1 0 680 0 -1 652
box 8 4 12 24
use welltap_svt  __well_tap__20
timestamp 1730743719
transform 1 0 104 0 1 688
box 8 4 12 24
use welltap_svt  __well_tap__20
timestamp 1730743719
transform 1 0 104 0 1 688
box 8 4 12 24
use welltap_svt  __well_tap__20
timestamp 1730743719
transform 1 0 104 0 1 688
box 8 4 12 24
use _0_0std_0_0cells_0_0AND2X1  and_559_6
timestamp 1730743719
transform 1 0 192 0 1 672
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_559_6
timestamp 1730743719
transform 1 0 192 0 1 672
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_559_6
timestamp 1730743719
transform 1 0 192 0 1 672
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_560_6
timestamp 1730743719
transform 1 0 232 0 1 672
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_560_6
timestamp 1730743719
transform 1 0 232 0 1 672
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_560_6
timestamp 1730743719
transform 1 0 232 0 1 672
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_561_6
timestamp 1730743719
transform 1 0 272 0 1 672
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_561_6
timestamp 1730743719
transform 1 0 272 0 1 672
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_561_6
timestamp 1730743719
transform 1 0 272 0 1 672
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_562_6
timestamp 1730743719
transform 1 0 312 0 1 672
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_562_6
timestamp 1730743719
transform 1 0 312 0 1 672
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_562_6
timestamp 1730743719
transform 1 0 312 0 1 672
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_567_6
timestamp 1730743719
transform 1 0 352 0 1 672
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_567_6
timestamp 1730743719
transform 1 0 352 0 1 672
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_567_6
timestamp 1730743719
transform 1 0 352 0 1 672
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_568_6
timestamp 1730743719
transform 1 0 400 0 1 672
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_568_6
timestamp 1730743719
transform 1 0 400 0 1 672
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_568_6
timestamp 1730743719
transform 1 0 400 0 1 672
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_569_6
timestamp 1730743719
transform 1 0 456 0 1 672
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_569_6
timestamp 1730743719
transform 1 0 456 0 1 672
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_569_6
timestamp 1730743719
transform 1 0 456 0 1 672
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_570_6
timestamp 1730743719
transform 1 0 520 0 1 672
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_570_6
timestamp 1730743719
transform 1 0 520 0 1 672
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_570_6
timestamp 1730743719
transform 1 0 520 0 1 672
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_597_6
timestamp 1730743719
transform 1 0 584 0 1 672
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_597_6
timestamp 1730743719
transform 1 0 584 0 1 672
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_597_6
timestamp 1730743719
transform 1 0 584 0 1 672
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_598_6
timestamp 1730743719
transform 1 0 632 0 1 672
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_598_6
timestamp 1730743719
transform 1 0 632 0 1 672
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_598_6
timestamp 1730743719
transform 1 0 632 0 1 672
box 8 4 36 49
use welltap_svt  __well_tap__21
timestamp 1730743719
transform 1 0 680 0 1 688
box 8 4 12 24
use welltap_svt  __well_tap__21
timestamp 1730743719
transform 1 0 680 0 1 688
box 8 4 12 24
use welltap_svt  __well_tap__21
timestamp 1730743719
transform 1 0 680 0 1 688
box 8 4 12 24
use welltap_svt  __well_tap__22
timestamp 1730743719
transform 1 0 104 0 -1 760
box 8 4 12 24
use welltap_svt  __well_tap__22
timestamp 1730743719
transform 1 0 104 0 -1 760
box 8 4 12 24
use welltap_svt  __well_tap__22
timestamp 1730743719
transform 1 0 104 0 -1 760
box 8 4 12 24
use _0_0std_0_0cells_0_0AND2X1  and_563_6
timestamp 1730743719
transform 1 0 272 0 -1 776
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_563_6
timestamp 1730743719
transform 1 0 272 0 -1 776
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_563_6
timestamp 1730743719
transform 1 0 272 0 -1 776
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_564_6
timestamp 1730743719
transform 1 0 360 0 -1 776
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_564_6
timestamp 1730743719
transform 1 0 360 0 -1 776
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_564_6
timestamp 1730743719
transform 1 0 360 0 -1 776
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_565_6
timestamp 1730743719
transform 1 0 456 0 -1 776
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_565_6
timestamp 1730743719
transform 1 0 456 0 -1 776
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_565_6
timestamp 1730743719
transform 1 0 456 0 -1 776
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_566_6
timestamp 1730743719
transform 1 0 552 0 -1 776
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_566_6
timestamp 1730743719
transform 1 0 552 0 -1 776
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_566_6
timestamp 1730743719
transform 1 0 552 0 -1 776
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_599_6
timestamp 1730743719
transform 1 0 632 0 -1 776
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_599_6
timestamp 1730743719
transform 1 0 632 0 -1 776
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_599_6
timestamp 1730743719
transform 1 0 632 0 -1 776
box 8 4 36 49
use welltap_svt  __well_tap__23
timestamp 1730743719
transform 1 0 680 0 -1 760
box 8 4 12 24
use welltap_svt  __well_tap__23
timestamp 1730743719
transform 1 0 680 0 -1 760
box 8 4 12 24
use welltap_svt  __well_tap__23
timestamp 1730743719
transform 1 0 680 0 -1 760
box 8 4 12 24
<< end >>
